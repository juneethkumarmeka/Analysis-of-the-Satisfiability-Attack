module basic_3000_30000_3500_60_levels_10xor_7(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999,N_25000,N_25001,N_25002,N_25003,N_25004,N_25005,N_25006,N_25007,N_25008,N_25009,N_25010,N_25011,N_25012,N_25013,N_25014,N_25015,N_25016,N_25017,N_25018,N_25019,N_25020,N_25021,N_25022,N_25023,N_25024,N_25025,N_25026,N_25027,N_25028,N_25029,N_25030,N_25031,N_25032,N_25033,N_25034,N_25035,N_25036,N_25037,N_25038,N_25039,N_25040,N_25041,N_25042,N_25043,N_25044,N_25045,N_25046,N_25047,N_25048,N_25049,N_25050,N_25051,N_25052,N_25053,N_25054,N_25055,N_25056,N_25057,N_25058,N_25059,N_25060,N_25061,N_25062,N_25063,N_25064,N_25065,N_25066,N_25067,N_25068,N_25069,N_25070,N_25071,N_25072,N_25073,N_25074,N_25075,N_25076,N_25077,N_25078,N_25079,N_25080,N_25081,N_25082,N_25083,N_25084,N_25085,N_25086,N_25087,N_25088,N_25089,N_25090,N_25091,N_25092,N_25093,N_25094,N_25095,N_25096,N_25097,N_25098,N_25099,N_25100,N_25101,N_25102,N_25103,N_25104,N_25105,N_25106,N_25107,N_25108,N_25109,N_25110,N_25111,N_25112,N_25113,N_25114,N_25115,N_25116,N_25117,N_25118,N_25119,N_25120,N_25121,N_25122,N_25123,N_25124,N_25125,N_25126,N_25127,N_25128,N_25129,N_25130,N_25131,N_25132,N_25133,N_25134,N_25135,N_25136,N_25137,N_25138,N_25139,N_25140,N_25141,N_25142,N_25143,N_25144,N_25145,N_25146,N_25147,N_25148,N_25149,N_25150,N_25151,N_25152,N_25153,N_25154,N_25155,N_25156,N_25157,N_25158,N_25159,N_25160,N_25161,N_25162,N_25163,N_25164,N_25165,N_25166,N_25167,N_25168,N_25169,N_25170,N_25171,N_25172,N_25173,N_25174,N_25175,N_25176,N_25177,N_25178,N_25179,N_25180,N_25181,N_25182,N_25183,N_25184,N_25185,N_25186,N_25187,N_25188,N_25189,N_25190,N_25191,N_25192,N_25193,N_25194,N_25195,N_25196,N_25197,N_25198,N_25199,N_25200,N_25201,N_25202,N_25203,N_25204,N_25205,N_25206,N_25207,N_25208,N_25209,N_25210,N_25211,N_25212,N_25213,N_25214,N_25215,N_25216,N_25217,N_25218,N_25219,N_25220,N_25221,N_25222,N_25223,N_25224,N_25225,N_25226,N_25227,N_25228,N_25229,N_25230,N_25231,N_25232,N_25233,N_25234,N_25235,N_25236,N_25237,N_25238,N_25239,N_25240,N_25241,N_25242,N_25243,N_25244,N_25245,N_25246,N_25247,N_25248,N_25249,N_25250,N_25251,N_25252,N_25253,N_25254,N_25255,N_25256,N_25257,N_25258,N_25259,N_25260,N_25261,N_25262,N_25263,N_25264,N_25265,N_25266,N_25267,N_25268,N_25269,N_25270,N_25271,N_25272,N_25273,N_25274,N_25275,N_25276,N_25277,N_25278,N_25279,N_25280,N_25281,N_25282,N_25283,N_25284,N_25285,N_25286,N_25287,N_25288,N_25289,N_25290,N_25291,N_25292,N_25293,N_25294,N_25295,N_25296,N_25297,N_25298,N_25299,N_25300,N_25301,N_25302,N_25303,N_25304,N_25305,N_25306,N_25307,N_25308,N_25309,N_25310,N_25311,N_25312,N_25313,N_25314,N_25315,N_25316,N_25317,N_25318,N_25319,N_25320,N_25321,N_25322,N_25323,N_25324,N_25325,N_25326,N_25327,N_25328,N_25329,N_25330,N_25331,N_25332,N_25333,N_25334,N_25335,N_25336,N_25337,N_25338,N_25339,N_25340,N_25341,N_25342,N_25343,N_25344,N_25345,N_25346,N_25347,N_25348,N_25349,N_25350,N_25351,N_25352,N_25353,N_25354,N_25355,N_25356,N_25357,N_25358,N_25359,N_25360,N_25361,N_25362,N_25363,N_25364,N_25365,N_25366,N_25367,N_25368,N_25369,N_25370,N_25371,N_25372,N_25373,N_25374,N_25375,N_25376,N_25377,N_25378,N_25379,N_25380,N_25381,N_25382,N_25383,N_25384,N_25385,N_25386,N_25387,N_25388,N_25389,N_25390,N_25391,N_25392,N_25393,N_25394,N_25395,N_25396,N_25397,N_25398,N_25399,N_25400,N_25401,N_25402,N_25403,N_25404,N_25405,N_25406,N_25407,N_25408,N_25409,N_25410,N_25411,N_25412,N_25413,N_25414,N_25415,N_25416,N_25417,N_25418,N_25419,N_25420,N_25421,N_25422,N_25423,N_25424,N_25425,N_25426,N_25427,N_25428,N_25429,N_25430,N_25431,N_25432,N_25433,N_25434,N_25435,N_25436,N_25437,N_25438,N_25439,N_25440,N_25441,N_25442,N_25443,N_25444,N_25445,N_25446,N_25447,N_25448,N_25449,N_25450,N_25451,N_25452,N_25453,N_25454,N_25455,N_25456,N_25457,N_25458,N_25459,N_25460,N_25461,N_25462,N_25463,N_25464,N_25465,N_25466,N_25467,N_25468,N_25469,N_25470,N_25471,N_25472,N_25473,N_25474,N_25475,N_25476,N_25477,N_25478,N_25479,N_25480,N_25481,N_25482,N_25483,N_25484,N_25485,N_25486,N_25487,N_25488,N_25489,N_25490,N_25491,N_25492,N_25493,N_25494,N_25495,N_25496,N_25497,N_25498,N_25499,N_25500,N_25501,N_25502,N_25503,N_25504,N_25505,N_25506,N_25507,N_25508,N_25509,N_25510,N_25511,N_25512,N_25513,N_25514,N_25515,N_25516,N_25517,N_25518,N_25519,N_25520,N_25521,N_25522,N_25523,N_25524,N_25525,N_25526,N_25527,N_25528,N_25529,N_25530,N_25531,N_25532,N_25533,N_25534,N_25535,N_25536,N_25537,N_25538,N_25539,N_25540,N_25541,N_25542,N_25543,N_25544,N_25545,N_25546,N_25547,N_25548,N_25549,N_25550,N_25551,N_25552,N_25553,N_25554,N_25555,N_25556,N_25557,N_25558,N_25559,N_25560,N_25561,N_25562,N_25563,N_25564,N_25565,N_25566,N_25567,N_25568,N_25569,N_25570,N_25571,N_25572,N_25573,N_25574,N_25575,N_25576,N_25577,N_25578,N_25579,N_25580,N_25581,N_25582,N_25583,N_25584,N_25585,N_25586,N_25587,N_25588,N_25589,N_25590,N_25591,N_25592,N_25593,N_25594,N_25595,N_25596,N_25597,N_25598,N_25599,N_25600,N_25601,N_25602,N_25603,N_25604,N_25605,N_25606,N_25607,N_25608,N_25609,N_25610,N_25611,N_25612,N_25613,N_25614,N_25615,N_25616,N_25617,N_25618,N_25619,N_25620,N_25621,N_25622,N_25623,N_25624,N_25625,N_25626,N_25627,N_25628,N_25629,N_25630,N_25631,N_25632,N_25633,N_25634,N_25635,N_25636,N_25637,N_25638,N_25639,N_25640,N_25641,N_25642,N_25643,N_25644,N_25645,N_25646,N_25647,N_25648,N_25649,N_25650,N_25651,N_25652,N_25653,N_25654,N_25655,N_25656,N_25657,N_25658,N_25659,N_25660,N_25661,N_25662,N_25663,N_25664,N_25665,N_25666,N_25667,N_25668,N_25669,N_25670,N_25671,N_25672,N_25673,N_25674,N_25675,N_25676,N_25677,N_25678,N_25679,N_25680,N_25681,N_25682,N_25683,N_25684,N_25685,N_25686,N_25687,N_25688,N_25689,N_25690,N_25691,N_25692,N_25693,N_25694,N_25695,N_25696,N_25697,N_25698,N_25699,N_25700,N_25701,N_25702,N_25703,N_25704,N_25705,N_25706,N_25707,N_25708,N_25709,N_25710,N_25711,N_25712,N_25713,N_25714,N_25715,N_25716,N_25717,N_25718,N_25719,N_25720,N_25721,N_25722,N_25723,N_25724,N_25725,N_25726,N_25727,N_25728,N_25729,N_25730,N_25731,N_25732,N_25733,N_25734,N_25735,N_25736,N_25737,N_25738,N_25739,N_25740,N_25741,N_25742,N_25743,N_25744,N_25745,N_25746,N_25747,N_25748,N_25749,N_25750,N_25751,N_25752,N_25753,N_25754,N_25755,N_25756,N_25757,N_25758,N_25759,N_25760,N_25761,N_25762,N_25763,N_25764,N_25765,N_25766,N_25767,N_25768,N_25769,N_25770,N_25771,N_25772,N_25773,N_25774,N_25775,N_25776,N_25777,N_25778,N_25779,N_25780,N_25781,N_25782,N_25783,N_25784,N_25785,N_25786,N_25787,N_25788,N_25789,N_25790,N_25791,N_25792,N_25793,N_25794,N_25795,N_25796,N_25797,N_25798,N_25799,N_25800,N_25801,N_25802,N_25803,N_25804,N_25805,N_25806,N_25807,N_25808,N_25809,N_25810,N_25811,N_25812,N_25813,N_25814,N_25815,N_25816,N_25817,N_25818,N_25819,N_25820,N_25821,N_25822,N_25823,N_25824,N_25825,N_25826,N_25827,N_25828,N_25829,N_25830,N_25831,N_25832,N_25833,N_25834,N_25835,N_25836,N_25837,N_25838,N_25839,N_25840,N_25841,N_25842,N_25843,N_25844,N_25845,N_25846,N_25847,N_25848,N_25849,N_25850,N_25851,N_25852,N_25853,N_25854,N_25855,N_25856,N_25857,N_25858,N_25859,N_25860,N_25861,N_25862,N_25863,N_25864,N_25865,N_25866,N_25867,N_25868,N_25869,N_25870,N_25871,N_25872,N_25873,N_25874,N_25875,N_25876,N_25877,N_25878,N_25879,N_25880,N_25881,N_25882,N_25883,N_25884,N_25885,N_25886,N_25887,N_25888,N_25889,N_25890,N_25891,N_25892,N_25893,N_25894,N_25895,N_25896,N_25897,N_25898,N_25899,N_25900,N_25901,N_25902,N_25903,N_25904,N_25905,N_25906,N_25907,N_25908,N_25909,N_25910,N_25911,N_25912,N_25913,N_25914,N_25915,N_25916,N_25917,N_25918,N_25919,N_25920,N_25921,N_25922,N_25923,N_25924,N_25925,N_25926,N_25927,N_25928,N_25929,N_25930,N_25931,N_25932,N_25933,N_25934,N_25935,N_25936,N_25937,N_25938,N_25939,N_25940,N_25941,N_25942,N_25943,N_25944,N_25945,N_25946,N_25947,N_25948,N_25949,N_25950,N_25951,N_25952,N_25953,N_25954,N_25955,N_25956,N_25957,N_25958,N_25959,N_25960,N_25961,N_25962,N_25963,N_25964,N_25965,N_25966,N_25967,N_25968,N_25969,N_25970,N_25971,N_25972,N_25973,N_25974,N_25975,N_25976,N_25977,N_25978,N_25979,N_25980,N_25981,N_25982,N_25983,N_25984,N_25985,N_25986,N_25987,N_25988,N_25989,N_25990,N_25991,N_25992,N_25993,N_25994,N_25995,N_25996,N_25997,N_25998,N_25999,N_26000,N_26001,N_26002,N_26003,N_26004,N_26005,N_26006,N_26007,N_26008,N_26009,N_26010,N_26011,N_26012,N_26013,N_26014,N_26015,N_26016,N_26017,N_26018,N_26019,N_26020,N_26021,N_26022,N_26023,N_26024,N_26025,N_26026,N_26027,N_26028,N_26029,N_26030,N_26031,N_26032,N_26033,N_26034,N_26035,N_26036,N_26037,N_26038,N_26039,N_26040,N_26041,N_26042,N_26043,N_26044,N_26045,N_26046,N_26047,N_26048,N_26049,N_26050,N_26051,N_26052,N_26053,N_26054,N_26055,N_26056,N_26057,N_26058,N_26059,N_26060,N_26061,N_26062,N_26063,N_26064,N_26065,N_26066,N_26067,N_26068,N_26069,N_26070,N_26071,N_26072,N_26073,N_26074,N_26075,N_26076,N_26077,N_26078,N_26079,N_26080,N_26081,N_26082,N_26083,N_26084,N_26085,N_26086,N_26087,N_26088,N_26089,N_26090,N_26091,N_26092,N_26093,N_26094,N_26095,N_26096,N_26097,N_26098,N_26099,N_26100,N_26101,N_26102,N_26103,N_26104,N_26105,N_26106,N_26107,N_26108,N_26109,N_26110,N_26111,N_26112,N_26113,N_26114,N_26115,N_26116,N_26117,N_26118,N_26119,N_26120,N_26121,N_26122,N_26123,N_26124,N_26125,N_26126,N_26127,N_26128,N_26129,N_26130,N_26131,N_26132,N_26133,N_26134,N_26135,N_26136,N_26137,N_26138,N_26139,N_26140,N_26141,N_26142,N_26143,N_26144,N_26145,N_26146,N_26147,N_26148,N_26149,N_26150,N_26151,N_26152,N_26153,N_26154,N_26155,N_26156,N_26157,N_26158,N_26159,N_26160,N_26161,N_26162,N_26163,N_26164,N_26165,N_26166,N_26167,N_26168,N_26169,N_26170,N_26171,N_26172,N_26173,N_26174,N_26175,N_26176,N_26177,N_26178,N_26179,N_26180,N_26181,N_26182,N_26183,N_26184,N_26185,N_26186,N_26187,N_26188,N_26189,N_26190,N_26191,N_26192,N_26193,N_26194,N_26195,N_26196,N_26197,N_26198,N_26199,N_26200,N_26201,N_26202,N_26203,N_26204,N_26205,N_26206,N_26207,N_26208,N_26209,N_26210,N_26211,N_26212,N_26213,N_26214,N_26215,N_26216,N_26217,N_26218,N_26219,N_26220,N_26221,N_26222,N_26223,N_26224,N_26225,N_26226,N_26227,N_26228,N_26229,N_26230,N_26231,N_26232,N_26233,N_26234,N_26235,N_26236,N_26237,N_26238,N_26239,N_26240,N_26241,N_26242,N_26243,N_26244,N_26245,N_26246,N_26247,N_26248,N_26249,N_26250,N_26251,N_26252,N_26253,N_26254,N_26255,N_26256,N_26257,N_26258,N_26259,N_26260,N_26261,N_26262,N_26263,N_26264,N_26265,N_26266,N_26267,N_26268,N_26269,N_26270,N_26271,N_26272,N_26273,N_26274,N_26275,N_26276,N_26277,N_26278,N_26279,N_26280,N_26281,N_26282,N_26283,N_26284,N_26285,N_26286,N_26287,N_26288,N_26289,N_26290,N_26291,N_26292,N_26293,N_26294,N_26295,N_26296,N_26297,N_26298,N_26299,N_26300,N_26301,N_26302,N_26303,N_26304,N_26305,N_26306,N_26307,N_26308,N_26309,N_26310,N_26311,N_26312,N_26313,N_26314,N_26315,N_26316,N_26317,N_26318,N_26319,N_26320,N_26321,N_26322,N_26323,N_26324,N_26325,N_26326,N_26327,N_26328,N_26329,N_26330,N_26331,N_26332,N_26333,N_26334,N_26335,N_26336,N_26337,N_26338,N_26339,N_26340,N_26341,N_26342,N_26343,N_26344,N_26345,N_26346,N_26347,N_26348,N_26349,N_26350,N_26351,N_26352,N_26353,N_26354,N_26355,N_26356,N_26357,N_26358,N_26359,N_26360,N_26361,N_26362,N_26363,N_26364,N_26365,N_26366,N_26367,N_26368,N_26369,N_26370,N_26371,N_26372,N_26373,N_26374,N_26375,N_26376,N_26377,N_26378,N_26379,N_26380,N_26381,N_26382,N_26383,N_26384,N_26385,N_26386,N_26387,N_26388,N_26389,N_26390,N_26391,N_26392,N_26393,N_26394,N_26395,N_26396,N_26397,N_26398,N_26399,N_26400,N_26401,N_26402,N_26403,N_26404,N_26405,N_26406,N_26407,N_26408,N_26409,N_26410,N_26411,N_26412,N_26413,N_26414,N_26415,N_26416,N_26417,N_26418,N_26419,N_26420,N_26421,N_26422,N_26423,N_26424,N_26425,N_26426,N_26427,N_26428,N_26429,N_26430,N_26431,N_26432,N_26433,N_26434,N_26435,N_26436,N_26437,N_26438,N_26439,N_26440,N_26441,N_26442,N_26443,N_26444,N_26445,N_26446,N_26447,N_26448,N_26449,N_26450,N_26451,N_26452,N_26453,N_26454,N_26455,N_26456,N_26457,N_26458,N_26459,N_26460,N_26461,N_26462,N_26463,N_26464,N_26465,N_26466,N_26467,N_26468,N_26469,N_26470,N_26471,N_26472,N_26473,N_26474,N_26475,N_26476,N_26477,N_26478,N_26479,N_26480,N_26481,N_26482,N_26483,N_26484,N_26485,N_26486,N_26487,N_26488,N_26489,N_26490,N_26491,N_26492,N_26493,N_26494,N_26495,N_26496,N_26497,N_26498,N_26499,N_26500,N_26501,N_26502,N_26503,N_26504,N_26505,N_26506,N_26507,N_26508,N_26509,N_26510,N_26511,N_26512,N_26513,N_26514,N_26515,N_26516,N_26517,N_26518,N_26519,N_26520,N_26521,N_26522,N_26523,N_26524,N_26525,N_26526,N_26527,N_26528,N_26529,N_26530,N_26531,N_26532,N_26533,N_26534,N_26535,N_26536,N_26537,N_26538,N_26539,N_26540,N_26541,N_26542,N_26543,N_26544,N_26545,N_26546,N_26547,N_26548,N_26549,N_26550,N_26551,N_26552,N_26553,N_26554,N_26555,N_26556,N_26557,N_26558,N_26559,N_26560,N_26561,N_26562,N_26563,N_26564,N_26565,N_26566,N_26567,N_26568,N_26569,N_26570,N_26571,N_26572,N_26573,N_26574,N_26575,N_26576,N_26577,N_26578,N_26579,N_26580,N_26581,N_26582,N_26583,N_26584,N_26585,N_26586,N_26587,N_26588,N_26589,N_26590,N_26591,N_26592,N_26593,N_26594,N_26595,N_26596,N_26597,N_26598,N_26599,N_26600,N_26601,N_26602,N_26603,N_26604,N_26605,N_26606,N_26607,N_26608,N_26609,N_26610,N_26611,N_26612,N_26613,N_26614,N_26615,N_26616,N_26617,N_26618,N_26619,N_26620,N_26621,N_26622,N_26623,N_26624,N_26625,N_26626,N_26627,N_26628,N_26629,N_26630,N_26631,N_26632,N_26633,N_26634,N_26635,N_26636,N_26637,N_26638,N_26639,N_26640,N_26641,N_26642,N_26643,N_26644,N_26645,N_26646,N_26647,N_26648,N_26649,N_26650,N_26651,N_26652,N_26653,N_26654,N_26655,N_26656,N_26657,N_26658,N_26659,N_26660,N_26661,N_26662,N_26663,N_26664,N_26665,N_26666,N_26667,N_26668,N_26669,N_26670,N_26671,N_26672,N_26673,N_26674,N_26675,N_26676,N_26677,N_26678,N_26679,N_26680,N_26681,N_26682,N_26683,N_26684,N_26685,N_26686,N_26687,N_26688,N_26689,N_26690,N_26691,N_26692,N_26693,N_26694,N_26695,N_26696,N_26697,N_26698,N_26699,N_26700,N_26701,N_26702,N_26703,N_26704,N_26705,N_26706,N_26707,N_26708,N_26709,N_26710,N_26711,N_26712,N_26713,N_26714,N_26715,N_26716,N_26717,N_26718,N_26719,N_26720,N_26721,N_26722,N_26723,N_26724,N_26725,N_26726,N_26727,N_26728,N_26729,N_26730,N_26731,N_26732,N_26733,N_26734,N_26735,N_26736,N_26737,N_26738,N_26739,N_26740,N_26741,N_26742,N_26743,N_26744,N_26745,N_26746,N_26747,N_26748,N_26749,N_26750,N_26751,N_26752,N_26753,N_26754,N_26755,N_26756,N_26757,N_26758,N_26759,N_26760,N_26761,N_26762,N_26763,N_26764,N_26765,N_26766,N_26767,N_26768,N_26769,N_26770,N_26771,N_26772,N_26773,N_26774,N_26775,N_26776,N_26777,N_26778,N_26779,N_26780,N_26781,N_26782,N_26783,N_26784,N_26785,N_26786,N_26787,N_26788,N_26789,N_26790,N_26791,N_26792,N_26793,N_26794,N_26795,N_26796,N_26797,N_26798,N_26799,N_26800,N_26801,N_26802,N_26803,N_26804,N_26805,N_26806,N_26807,N_26808,N_26809,N_26810,N_26811,N_26812,N_26813,N_26814,N_26815,N_26816,N_26817,N_26818,N_26819,N_26820,N_26821,N_26822,N_26823,N_26824,N_26825,N_26826,N_26827,N_26828,N_26829,N_26830,N_26831,N_26832,N_26833,N_26834,N_26835,N_26836,N_26837,N_26838,N_26839,N_26840,N_26841,N_26842,N_26843,N_26844,N_26845,N_26846,N_26847,N_26848,N_26849,N_26850,N_26851,N_26852,N_26853,N_26854,N_26855,N_26856,N_26857,N_26858,N_26859,N_26860,N_26861,N_26862,N_26863,N_26864,N_26865,N_26866,N_26867,N_26868,N_26869,N_26870,N_26871,N_26872,N_26873,N_26874,N_26875,N_26876,N_26877,N_26878,N_26879,N_26880,N_26881,N_26882,N_26883,N_26884,N_26885,N_26886,N_26887,N_26888,N_26889,N_26890,N_26891,N_26892,N_26893,N_26894,N_26895,N_26896,N_26897,N_26898,N_26899,N_26900,N_26901,N_26902,N_26903,N_26904,N_26905,N_26906,N_26907,N_26908,N_26909,N_26910,N_26911,N_26912,N_26913,N_26914,N_26915,N_26916,N_26917,N_26918,N_26919,N_26920,N_26921,N_26922,N_26923,N_26924,N_26925,N_26926,N_26927,N_26928,N_26929,N_26930,N_26931,N_26932,N_26933,N_26934,N_26935,N_26936,N_26937,N_26938,N_26939,N_26940,N_26941,N_26942,N_26943,N_26944,N_26945,N_26946,N_26947,N_26948,N_26949,N_26950,N_26951,N_26952,N_26953,N_26954,N_26955,N_26956,N_26957,N_26958,N_26959,N_26960,N_26961,N_26962,N_26963,N_26964,N_26965,N_26966,N_26967,N_26968,N_26969,N_26970,N_26971,N_26972,N_26973,N_26974,N_26975,N_26976,N_26977,N_26978,N_26979,N_26980,N_26981,N_26982,N_26983,N_26984,N_26985,N_26986,N_26987,N_26988,N_26989,N_26990,N_26991,N_26992,N_26993,N_26994,N_26995,N_26996,N_26997,N_26998,N_26999,N_27000,N_27001,N_27002,N_27003,N_27004,N_27005,N_27006,N_27007,N_27008,N_27009,N_27010,N_27011,N_27012,N_27013,N_27014,N_27015,N_27016,N_27017,N_27018,N_27019,N_27020,N_27021,N_27022,N_27023,N_27024,N_27025,N_27026,N_27027,N_27028,N_27029,N_27030,N_27031,N_27032,N_27033,N_27034,N_27035,N_27036,N_27037,N_27038,N_27039,N_27040,N_27041,N_27042,N_27043,N_27044,N_27045,N_27046,N_27047,N_27048,N_27049,N_27050,N_27051,N_27052,N_27053,N_27054,N_27055,N_27056,N_27057,N_27058,N_27059,N_27060,N_27061,N_27062,N_27063,N_27064,N_27065,N_27066,N_27067,N_27068,N_27069,N_27070,N_27071,N_27072,N_27073,N_27074,N_27075,N_27076,N_27077,N_27078,N_27079,N_27080,N_27081,N_27082,N_27083,N_27084,N_27085,N_27086,N_27087,N_27088,N_27089,N_27090,N_27091,N_27092,N_27093,N_27094,N_27095,N_27096,N_27097,N_27098,N_27099,N_27100,N_27101,N_27102,N_27103,N_27104,N_27105,N_27106,N_27107,N_27108,N_27109,N_27110,N_27111,N_27112,N_27113,N_27114,N_27115,N_27116,N_27117,N_27118,N_27119,N_27120,N_27121,N_27122,N_27123,N_27124,N_27125,N_27126,N_27127,N_27128,N_27129,N_27130,N_27131,N_27132,N_27133,N_27134,N_27135,N_27136,N_27137,N_27138,N_27139,N_27140,N_27141,N_27142,N_27143,N_27144,N_27145,N_27146,N_27147,N_27148,N_27149,N_27150,N_27151,N_27152,N_27153,N_27154,N_27155,N_27156,N_27157,N_27158,N_27159,N_27160,N_27161,N_27162,N_27163,N_27164,N_27165,N_27166,N_27167,N_27168,N_27169,N_27170,N_27171,N_27172,N_27173,N_27174,N_27175,N_27176,N_27177,N_27178,N_27179,N_27180,N_27181,N_27182,N_27183,N_27184,N_27185,N_27186,N_27187,N_27188,N_27189,N_27190,N_27191,N_27192,N_27193,N_27194,N_27195,N_27196,N_27197,N_27198,N_27199,N_27200,N_27201,N_27202,N_27203,N_27204,N_27205,N_27206,N_27207,N_27208,N_27209,N_27210,N_27211,N_27212,N_27213,N_27214,N_27215,N_27216,N_27217,N_27218,N_27219,N_27220,N_27221,N_27222,N_27223,N_27224,N_27225,N_27226,N_27227,N_27228,N_27229,N_27230,N_27231,N_27232,N_27233,N_27234,N_27235,N_27236,N_27237,N_27238,N_27239,N_27240,N_27241,N_27242,N_27243,N_27244,N_27245,N_27246,N_27247,N_27248,N_27249,N_27250,N_27251,N_27252,N_27253,N_27254,N_27255,N_27256,N_27257,N_27258,N_27259,N_27260,N_27261,N_27262,N_27263,N_27264,N_27265,N_27266,N_27267,N_27268,N_27269,N_27270,N_27271,N_27272,N_27273,N_27274,N_27275,N_27276,N_27277,N_27278,N_27279,N_27280,N_27281,N_27282,N_27283,N_27284,N_27285,N_27286,N_27287,N_27288,N_27289,N_27290,N_27291,N_27292,N_27293,N_27294,N_27295,N_27296,N_27297,N_27298,N_27299,N_27300,N_27301,N_27302,N_27303,N_27304,N_27305,N_27306,N_27307,N_27308,N_27309,N_27310,N_27311,N_27312,N_27313,N_27314,N_27315,N_27316,N_27317,N_27318,N_27319,N_27320,N_27321,N_27322,N_27323,N_27324,N_27325,N_27326,N_27327,N_27328,N_27329,N_27330,N_27331,N_27332,N_27333,N_27334,N_27335,N_27336,N_27337,N_27338,N_27339,N_27340,N_27341,N_27342,N_27343,N_27344,N_27345,N_27346,N_27347,N_27348,N_27349,N_27350,N_27351,N_27352,N_27353,N_27354,N_27355,N_27356,N_27357,N_27358,N_27359,N_27360,N_27361,N_27362,N_27363,N_27364,N_27365,N_27366,N_27367,N_27368,N_27369,N_27370,N_27371,N_27372,N_27373,N_27374,N_27375,N_27376,N_27377,N_27378,N_27379,N_27380,N_27381,N_27382,N_27383,N_27384,N_27385,N_27386,N_27387,N_27388,N_27389,N_27390,N_27391,N_27392,N_27393,N_27394,N_27395,N_27396,N_27397,N_27398,N_27399,N_27400,N_27401,N_27402,N_27403,N_27404,N_27405,N_27406,N_27407,N_27408,N_27409,N_27410,N_27411,N_27412,N_27413,N_27414,N_27415,N_27416,N_27417,N_27418,N_27419,N_27420,N_27421,N_27422,N_27423,N_27424,N_27425,N_27426,N_27427,N_27428,N_27429,N_27430,N_27431,N_27432,N_27433,N_27434,N_27435,N_27436,N_27437,N_27438,N_27439,N_27440,N_27441,N_27442,N_27443,N_27444,N_27445,N_27446,N_27447,N_27448,N_27449,N_27450,N_27451,N_27452,N_27453,N_27454,N_27455,N_27456,N_27457,N_27458,N_27459,N_27460,N_27461,N_27462,N_27463,N_27464,N_27465,N_27466,N_27467,N_27468,N_27469,N_27470,N_27471,N_27472,N_27473,N_27474,N_27475,N_27476,N_27477,N_27478,N_27479,N_27480,N_27481,N_27482,N_27483,N_27484,N_27485,N_27486,N_27487,N_27488,N_27489,N_27490,N_27491,N_27492,N_27493,N_27494,N_27495,N_27496,N_27497,N_27498,N_27499,N_27500,N_27501,N_27502,N_27503,N_27504,N_27505,N_27506,N_27507,N_27508,N_27509,N_27510,N_27511,N_27512,N_27513,N_27514,N_27515,N_27516,N_27517,N_27518,N_27519,N_27520,N_27521,N_27522,N_27523,N_27524,N_27525,N_27526,N_27527,N_27528,N_27529,N_27530,N_27531,N_27532,N_27533,N_27534,N_27535,N_27536,N_27537,N_27538,N_27539,N_27540,N_27541,N_27542,N_27543,N_27544,N_27545,N_27546,N_27547,N_27548,N_27549,N_27550,N_27551,N_27552,N_27553,N_27554,N_27555,N_27556,N_27557,N_27558,N_27559,N_27560,N_27561,N_27562,N_27563,N_27564,N_27565,N_27566,N_27567,N_27568,N_27569,N_27570,N_27571,N_27572,N_27573,N_27574,N_27575,N_27576,N_27577,N_27578,N_27579,N_27580,N_27581,N_27582,N_27583,N_27584,N_27585,N_27586,N_27587,N_27588,N_27589,N_27590,N_27591,N_27592,N_27593,N_27594,N_27595,N_27596,N_27597,N_27598,N_27599,N_27600,N_27601,N_27602,N_27603,N_27604,N_27605,N_27606,N_27607,N_27608,N_27609,N_27610,N_27611,N_27612,N_27613,N_27614,N_27615,N_27616,N_27617,N_27618,N_27619,N_27620,N_27621,N_27622,N_27623,N_27624,N_27625,N_27626,N_27627,N_27628,N_27629,N_27630,N_27631,N_27632,N_27633,N_27634,N_27635,N_27636,N_27637,N_27638,N_27639,N_27640,N_27641,N_27642,N_27643,N_27644,N_27645,N_27646,N_27647,N_27648,N_27649,N_27650,N_27651,N_27652,N_27653,N_27654,N_27655,N_27656,N_27657,N_27658,N_27659,N_27660,N_27661,N_27662,N_27663,N_27664,N_27665,N_27666,N_27667,N_27668,N_27669,N_27670,N_27671,N_27672,N_27673,N_27674,N_27675,N_27676,N_27677,N_27678,N_27679,N_27680,N_27681,N_27682,N_27683,N_27684,N_27685,N_27686,N_27687,N_27688,N_27689,N_27690,N_27691,N_27692,N_27693,N_27694,N_27695,N_27696,N_27697,N_27698,N_27699,N_27700,N_27701,N_27702,N_27703,N_27704,N_27705,N_27706,N_27707,N_27708,N_27709,N_27710,N_27711,N_27712,N_27713,N_27714,N_27715,N_27716,N_27717,N_27718,N_27719,N_27720,N_27721,N_27722,N_27723,N_27724,N_27725,N_27726,N_27727,N_27728,N_27729,N_27730,N_27731,N_27732,N_27733,N_27734,N_27735,N_27736,N_27737,N_27738,N_27739,N_27740,N_27741,N_27742,N_27743,N_27744,N_27745,N_27746,N_27747,N_27748,N_27749,N_27750,N_27751,N_27752,N_27753,N_27754,N_27755,N_27756,N_27757,N_27758,N_27759,N_27760,N_27761,N_27762,N_27763,N_27764,N_27765,N_27766,N_27767,N_27768,N_27769,N_27770,N_27771,N_27772,N_27773,N_27774,N_27775,N_27776,N_27777,N_27778,N_27779,N_27780,N_27781,N_27782,N_27783,N_27784,N_27785,N_27786,N_27787,N_27788,N_27789,N_27790,N_27791,N_27792,N_27793,N_27794,N_27795,N_27796,N_27797,N_27798,N_27799,N_27800,N_27801,N_27802,N_27803,N_27804,N_27805,N_27806,N_27807,N_27808,N_27809,N_27810,N_27811,N_27812,N_27813,N_27814,N_27815,N_27816,N_27817,N_27818,N_27819,N_27820,N_27821,N_27822,N_27823,N_27824,N_27825,N_27826,N_27827,N_27828,N_27829,N_27830,N_27831,N_27832,N_27833,N_27834,N_27835,N_27836,N_27837,N_27838,N_27839,N_27840,N_27841,N_27842,N_27843,N_27844,N_27845,N_27846,N_27847,N_27848,N_27849,N_27850,N_27851,N_27852,N_27853,N_27854,N_27855,N_27856,N_27857,N_27858,N_27859,N_27860,N_27861,N_27862,N_27863,N_27864,N_27865,N_27866,N_27867,N_27868,N_27869,N_27870,N_27871,N_27872,N_27873,N_27874,N_27875,N_27876,N_27877,N_27878,N_27879,N_27880,N_27881,N_27882,N_27883,N_27884,N_27885,N_27886,N_27887,N_27888,N_27889,N_27890,N_27891,N_27892,N_27893,N_27894,N_27895,N_27896,N_27897,N_27898,N_27899,N_27900,N_27901,N_27902,N_27903,N_27904,N_27905,N_27906,N_27907,N_27908,N_27909,N_27910,N_27911,N_27912,N_27913,N_27914,N_27915,N_27916,N_27917,N_27918,N_27919,N_27920,N_27921,N_27922,N_27923,N_27924,N_27925,N_27926,N_27927,N_27928,N_27929,N_27930,N_27931,N_27932,N_27933,N_27934,N_27935,N_27936,N_27937,N_27938,N_27939,N_27940,N_27941,N_27942,N_27943,N_27944,N_27945,N_27946,N_27947,N_27948,N_27949,N_27950,N_27951,N_27952,N_27953,N_27954,N_27955,N_27956,N_27957,N_27958,N_27959,N_27960,N_27961,N_27962,N_27963,N_27964,N_27965,N_27966,N_27967,N_27968,N_27969,N_27970,N_27971,N_27972,N_27973,N_27974,N_27975,N_27976,N_27977,N_27978,N_27979,N_27980,N_27981,N_27982,N_27983,N_27984,N_27985,N_27986,N_27987,N_27988,N_27989,N_27990,N_27991,N_27992,N_27993,N_27994,N_27995,N_27996,N_27997,N_27998,N_27999,N_28000,N_28001,N_28002,N_28003,N_28004,N_28005,N_28006,N_28007,N_28008,N_28009,N_28010,N_28011,N_28012,N_28013,N_28014,N_28015,N_28016,N_28017,N_28018,N_28019,N_28020,N_28021,N_28022,N_28023,N_28024,N_28025,N_28026,N_28027,N_28028,N_28029,N_28030,N_28031,N_28032,N_28033,N_28034,N_28035,N_28036,N_28037,N_28038,N_28039,N_28040,N_28041,N_28042,N_28043,N_28044,N_28045,N_28046,N_28047,N_28048,N_28049,N_28050,N_28051,N_28052,N_28053,N_28054,N_28055,N_28056,N_28057,N_28058,N_28059,N_28060,N_28061,N_28062,N_28063,N_28064,N_28065,N_28066,N_28067,N_28068,N_28069,N_28070,N_28071,N_28072,N_28073,N_28074,N_28075,N_28076,N_28077,N_28078,N_28079,N_28080,N_28081,N_28082,N_28083,N_28084,N_28085,N_28086,N_28087,N_28088,N_28089,N_28090,N_28091,N_28092,N_28093,N_28094,N_28095,N_28096,N_28097,N_28098,N_28099,N_28100,N_28101,N_28102,N_28103,N_28104,N_28105,N_28106,N_28107,N_28108,N_28109,N_28110,N_28111,N_28112,N_28113,N_28114,N_28115,N_28116,N_28117,N_28118,N_28119,N_28120,N_28121,N_28122,N_28123,N_28124,N_28125,N_28126,N_28127,N_28128,N_28129,N_28130,N_28131,N_28132,N_28133,N_28134,N_28135,N_28136,N_28137,N_28138,N_28139,N_28140,N_28141,N_28142,N_28143,N_28144,N_28145,N_28146,N_28147,N_28148,N_28149,N_28150,N_28151,N_28152,N_28153,N_28154,N_28155,N_28156,N_28157,N_28158,N_28159,N_28160,N_28161,N_28162,N_28163,N_28164,N_28165,N_28166,N_28167,N_28168,N_28169,N_28170,N_28171,N_28172,N_28173,N_28174,N_28175,N_28176,N_28177,N_28178,N_28179,N_28180,N_28181,N_28182,N_28183,N_28184,N_28185,N_28186,N_28187,N_28188,N_28189,N_28190,N_28191,N_28192,N_28193,N_28194,N_28195,N_28196,N_28197,N_28198,N_28199,N_28200,N_28201,N_28202,N_28203,N_28204,N_28205,N_28206,N_28207,N_28208,N_28209,N_28210,N_28211,N_28212,N_28213,N_28214,N_28215,N_28216,N_28217,N_28218,N_28219,N_28220,N_28221,N_28222,N_28223,N_28224,N_28225,N_28226,N_28227,N_28228,N_28229,N_28230,N_28231,N_28232,N_28233,N_28234,N_28235,N_28236,N_28237,N_28238,N_28239,N_28240,N_28241,N_28242,N_28243,N_28244,N_28245,N_28246,N_28247,N_28248,N_28249,N_28250,N_28251,N_28252,N_28253,N_28254,N_28255,N_28256,N_28257,N_28258,N_28259,N_28260,N_28261,N_28262,N_28263,N_28264,N_28265,N_28266,N_28267,N_28268,N_28269,N_28270,N_28271,N_28272,N_28273,N_28274,N_28275,N_28276,N_28277,N_28278,N_28279,N_28280,N_28281,N_28282,N_28283,N_28284,N_28285,N_28286,N_28287,N_28288,N_28289,N_28290,N_28291,N_28292,N_28293,N_28294,N_28295,N_28296,N_28297,N_28298,N_28299,N_28300,N_28301,N_28302,N_28303,N_28304,N_28305,N_28306,N_28307,N_28308,N_28309,N_28310,N_28311,N_28312,N_28313,N_28314,N_28315,N_28316,N_28317,N_28318,N_28319,N_28320,N_28321,N_28322,N_28323,N_28324,N_28325,N_28326,N_28327,N_28328,N_28329,N_28330,N_28331,N_28332,N_28333,N_28334,N_28335,N_28336,N_28337,N_28338,N_28339,N_28340,N_28341,N_28342,N_28343,N_28344,N_28345,N_28346,N_28347,N_28348,N_28349,N_28350,N_28351,N_28352,N_28353,N_28354,N_28355,N_28356,N_28357,N_28358,N_28359,N_28360,N_28361,N_28362,N_28363,N_28364,N_28365,N_28366,N_28367,N_28368,N_28369,N_28370,N_28371,N_28372,N_28373,N_28374,N_28375,N_28376,N_28377,N_28378,N_28379,N_28380,N_28381,N_28382,N_28383,N_28384,N_28385,N_28386,N_28387,N_28388,N_28389,N_28390,N_28391,N_28392,N_28393,N_28394,N_28395,N_28396,N_28397,N_28398,N_28399,N_28400,N_28401,N_28402,N_28403,N_28404,N_28405,N_28406,N_28407,N_28408,N_28409,N_28410,N_28411,N_28412,N_28413,N_28414,N_28415,N_28416,N_28417,N_28418,N_28419,N_28420,N_28421,N_28422,N_28423,N_28424,N_28425,N_28426,N_28427,N_28428,N_28429,N_28430,N_28431,N_28432,N_28433,N_28434,N_28435,N_28436,N_28437,N_28438,N_28439,N_28440,N_28441,N_28442,N_28443,N_28444,N_28445,N_28446,N_28447,N_28448,N_28449,N_28450,N_28451,N_28452,N_28453,N_28454,N_28455,N_28456,N_28457,N_28458,N_28459,N_28460,N_28461,N_28462,N_28463,N_28464,N_28465,N_28466,N_28467,N_28468,N_28469,N_28470,N_28471,N_28472,N_28473,N_28474,N_28475,N_28476,N_28477,N_28478,N_28479,N_28480,N_28481,N_28482,N_28483,N_28484,N_28485,N_28486,N_28487,N_28488,N_28489,N_28490,N_28491,N_28492,N_28493,N_28494,N_28495,N_28496,N_28497,N_28498,N_28499,N_28500,N_28501,N_28502,N_28503,N_28504,N_28505,N_28506,N_28507,N_28508,N_28509,N_28510,N_28511,N_28512,N_28513,N_28514,N_28515,N_28516,N_28517,N_28518,N_28519,N_28520,N_28521,N_28522,N_28523,N_28524,N_28525,N_28526,N_28527,N_28528,N_28529,N_28530,N_28531,N_28532,N_28533,N_28534,N_28535,N_28536,N_28537,N_28538,N_28539,N_28540,N_28541,N_28542,N_28543,N_28544,N_28545,N_28546,N_28547,N_28548,N_28549,N_28550,N_28551,N_28552,N_28553,N_28554,N_28555,N_28556,N_28557,N_28558,N_28559,N_28560,N_28561,N_28562,N_28563,N_28564,N_28565,N_28566,N_28567,N_28568,N_28569,N_28570,N_28571,N_28572,N_28573,N_28574,N_28575,N_28576,N_28577,N_28578,N_28579,N_28580,N_28581,N_28582,N_28583,N_28584,N_28585,N_28586,N_28587,N_28588,N_28589,N_28590,N_28591,N_28592,N_28593,N_28594,N_28595,N_28596,N_28597,N_28598,N_28599,N_28600,N_28601,N_28602,N_28603,N_28604,N_28605,N_28606,N_28607,N_28608,N_28609,N_28610,N_28611,N_28612,N_28613,N_28614,N_28615,N_28616,N_28617,N_28618,N_28619,N_28620,N_28621,N_28622,N_28623,N_28624,N_28625,N_28626,N_28627,N_28628,N_28629,N_28630,N_28631,N_28632,N_28633,N_28634,N_28635,N_28636,N_28637,N_28638,N_28639,N_28640,N_28641,N_28642,N_28643,N_28644,N_28645,N_28646,N_28647,N_28648,N_28649,N_28650,N_28651,N_28652,N_28653,N_28654,N_28655,N_28656,N_28657,N_28658,N_28659,N_28660,N_28661,N_28662,N_28663,N_28664,N_28665,N_28666,N_28667,N_28668,N_28669,N_28670,N_28671,N_28672,N_28673,N_28674,N_28675,N_28676,N_28677,N_28678,N_28679,N_28680,N_28681,N_28682,N_28683,N_28684,N_28685,N_28686,N_28687,N_28688,N_28689,N_28690,N_28691,N_28692,N_28693,N_28694,N_28695,N_28696,N_28697,N_28698,N_28699,N_28700,N_28701,N_28702,N_28703,N_28704,N_28705,N_28706,N_28707,N_28708,N_28709,N_28710,N_28711,N_28712,N_28713,N_28714,N_28715,N_28716,N_28717,N_28718,N_28719,N_28720,N_28721,N_28722,N_28723,N_28724,N_28725,N_28726,N_28727,N_28728,N_28729,N_28730,N_28731,N_28732,N_28733,N_28734,N_28735,N_28736,N_28737,N_28738,N_28739,N_28740,N_28741,N_28742,N_28743,N_28744,N_28745,N_28746,N_28747,N_28748,N_28749,N_28750,N_28751,N_28752,N_28753,N_28754,N_28755,N_28756,N_28757,N_28758,N_28759,N_28760,N_28761,N_28762,N_28763,N_28764,N_28765,N_28766,N_28767,N_28768,N_28769,N_28770,N_28771,N_28772,N_28773,N_28774,N_28775,N_28776,N_28777,N_28778,N_28779,N_28780,N_28781,N_28782,N_28783,N_28784,N_28785,N_28786,N_28787,N_28788,N_28789,N_28790,N_28791,N_28792,N_28793,N_28794,N_28795,N_28796,N_28797,N_28798,N_28799,N_28800,N_28801,N_28802,N_28803,N_28804,N_28805,N_28806,N_28807,N_28808,N_28809,N_28810,N_28811,N_28812,N_28813,N_28814,N_28815,N_28816,N_28817,N_28818,N_28819,N_28820,N_28821,N_28822,N_28823,N_28824,N_28825,N_28826,N_28827,N_28828,N_28829,N_28830,N_28831,N_28832,N_28833,N_28834,N_28835,N_28836,N_28837,N_28838,N_28839,N_28840,N_28841,N_28842,N_28843,N_28844,N_28845,N_28846,N_28847,N_28848,N_28849,N_28850,N_28851,N_28852,N_28853,N_28854,N_28855,N_28856,N_28857,N_28858,N_28859,N_28860,N_28861,N_28862,N_28863,N_28864,N_28865,N_28866,N_28867,N_28868,N_28869,N_28870,N_28871,N_28872,N_28873,N_28874,N_28875,N_28876,N_28877,N_28878,N_28879,N_28880,N_28881,N_28882,N_28883,N_28884,N_28885,N_28886,N_28887,N_28888,N_28889,N_28890,N_28891,N_28892,N_28893,N_28894,N_28895,N_28896,N_28897,N_28898,N_28899,N_28900,N_28901,N_28902,N_28903,N_28904,N_28905,N_28906,N_28907,N_28908,N_28909,N_28910,N_28911,N_28912,N_28913,N_28914,N_28915,N_28916,N_28917,N_28918,N_28919,N_28920,N_28921,N_28922,N_28923,N_28924,N_28925,N_28926,N_28927,N_28928,N_28929,N_28930,N_28931,N_28932,N_28933,N_28934,N_28935,N_28936,N_28937,N_28938,N_28939,N_28940,N_28941,N_28942,N_28943,N_28944,N_28945,N_28946,N_28947,N_28948,N_28949,N_28950,N_28951,N_28952,N_28953,N_28954,N_28955,N_28956,N_28957,N_28958,N_28959,N_28960,N_28961,N_28962,N_28963,N_28964,N_28965,N_28966,N_28967,N_28968,N_28969,N_28970,N_28971,N_28972,N_28973,N_28974,N_28975,N_28976,N_28977,N_28978,N_28979,N_28980,N_28981,N_28982,N_28983,N_28984,N_28985,N_28986,N_28987,N_28988,N_28989,N_28990,N_28991,N_28992,N_28993,N_28994,N_28995,N_28996,N_28997,N_28998,N_28999,N_29000,N_29001,N_29002,N_29003,N_29004,N_29005,N_29006,N_29007,N_29008,N_29009,N_29010,N_29011,N_29012,N_29013,N_29014,N_29015,N_29016,N_29017,N_29018,N_29019,N_29020,N_29021,N_29022,N_29023,N_29024,N_29025,N_29026,N_29027,N_29028,N_29029,N_29030,N_29031,N_29032,N_29033,N_29034,N_29035,N_29036,N_29037,N_29038,N_29039,N_29040,N_29041,N_29042,N_29043,N_29044,N_29045,N_29046,N_29047,N_29048,N_29049,N_29050,N_29051,N_29052,N_29053,N_29054,N_29055,N_29056,N_29057,N_29058,N_29059,N_29060,N_29061,N_29062,N_29063,N_29064,N_29065,N_29066,N_29067,N_29068,N_29069,N_29070,N_29071,N_29072,N_29073,N_29074,N_29075,N_29076,N_29077,N_29078,N_29079,N_29080,N_29081,N_29082,N_29083,N_29084,N_29085,N_29086,N_29087,N_29088,N_29089,N_29090,N_29091,N_29092,N_29093,N_29094,N_29095,N_29096,N_29097,N_29098,N_29099,N_29100,N_29101,N_29102,N_29103,N_29104,N_29105,N_29106,N_29107,N_29108,N_29109,N_29110,N_29111,N_29112,N_29113,N_29114,N_29115,N_29116,N_29117,N_29118,N_29119,N_29120,N_29121,N_29122,N_29123,N_29124,N_29125,N_29126,N_29127,N_29128,N_29129,N_29130,N_29131,N_29132,N_29133,N_29134,N_29135,N_29136,N_29137,N_29138,N_29139,N_29140,N_29141,N_29142,N_29143,N_29144,N_29145,N_29146,N_29147,N_29148,N_29149,N_29150,N_29151,N_29152,N_29153,N_29154,N_29155,N_29156,N_29157,N_29158,N_29159,N_29160,N_29161,N_29162,N_29163,N_29164,N_29165,N_29166,N_29167,N_29168,N_29169,N_29170,N_29171,N_29172,N_29173,N_29174,N_29175,N_29176,N_29177,N_29178,N_29179,N_29180,N_29181,N_29182,N_29183,N_29184,N_29185,N_29186,N_29187,N_29188,N_29189,N_29190,N_29191,N_29192,N_29193,N_29194,N_29195,N_29196,N_29197,N_29198,N_29199,N_29200,N_29201,N_29202,N_29203,N_29204,N_29205,N_29206,N_29207,N_29208,N_29209,N_29210,N_29211,N_29212,N_29213,N_29214,N_29215,N_29216,N_29217,N_29218,N_29219,N_29220,N_29221,N_29222,N_29223,N_29224,N_29225,N_29226,N_29227,N_29228,N_29229,N_29230,N_29231,N_29232,N_29233,N_29234,N_29235,N_29236,N_29237,N_29238,N_29239,N_29240,N_29241,N_29242,N_29243,N_29244,N_29245,N_29246,N_29247,N_29248,N_29249,N_29250,N_29251,N_29252,N_29253,N_29254,N_29255,N_29256,N_29257,N_29258,N_29259,N_29260,N_29261,N_29262,N_29263,N_29264,N_29265,N_29266,N_29267,N_29268,N_29269,N_29270,N_29271,N_29272,N_29273,N_29274,N_29275,N_29276,N_29277,N_29278,N_29279,N_29280,N_29281,N_29282,N_29283,N_29284,N_29285,N_29286,N_29287,N_29288,N_29289,N_29290,N_29291,N_29292,N_29293,N_29294,N_29295,N_29296,N_29297,N_29298,N_29299,N_29300,N_29301,N_29302,N_29303,N_29304,N_29305,N_29306,N_29307,N_29308,N_29309,N_29310,N_29311,N_29312,N_29313,N_29314,N_29315,N_29316,N_29317,N_29318,N_29319,N_29320,N_29321,N_29322,N_29323,N_29324,N_29325,N_29326,N_29327,N_29328,N_29329,N_29330,N_29331,N_29332,N_29333,N_29334,N_29335,N_29336,N_29337,N_29338,N_29339,N_29340,N_29341,N_29342,N_29343,N_29344,N_29345,N_29346,N_29347,N_29348,N_29349,N_29350,N_29351,N_29352,N_29353,N_29354,N_29355,N_29356,N_29357,N_29358,N_29359,N_29360,N_29361,N_29362,N_29363,N_29364,N_29365,N_29366,N_29367,N_29368,N_29369,N_29370,N_29371,N_29372,N_29373,N_29374,N_29375,N_29376,N_29377,N_29378,N_29379,N_29380,N_29381,N_29382,N_29383,N_29384,N_29385,N_29386,N_29387,N_29388,N_29389,N_29390,N_29391,N_29392,N_29393,N_29394,N_29395,N_29396,N_29397,N_29398,N_29399,N_29400,N_29401,N_29402,N_29403,N_29404,N_29405,N_29406,N_29407,N_29408,N_29409,N_29410,N_29411,N_29412,N_29413,N_29414,N_29415,N_29416,N_29417,N_29418,N_29419,N_29420,N_29421,N_29422,N_29423,N_29424,N_29425,N_29426,N_29427,N_29428,N_29429,N_29430,N_29431,N_29432,N_29433,N_29434,N_29435,N_29436,N_29437,N_29438,N_29439,N_29440,N_29441,N_29442,N_29443,N_29444,N_29445,N_29446,N_29447,N_29448,N_29449,N_29450,N_29451,N_29452,N_29453,N_29454,N_29455,N_29456,N_29457,N_29458,N_29459,N_29460,N_29461,N_29462,N_29463,N_29464,N_29465,N_29466,N_29467,N_29468,N_29469,N_29470,N_29471,N_29472,N_29473,N_29474,N_29475,N_29476,N_29477,N_29478,N_29479,N_29480,N_29481,N_29482,N_29483,N_29484,N_29485,N_29486,N_29487,N_29488,N_29489,N_29490,N_29491,N_29492,N_29493,N_29494,N_29495,N_29496,N_29497,N_29498,N_29499,N_29500,N_29501,N_29502,N_29503,N_29504,N_29505,N_29506,N_29507,N_29508,N_29509,N_29510,N_29511,N_29512,N_29513,N_29514,N_29515,N_29516,N_29517,N_29518,N_29519,N_29520,N_29521,N_29522,N_29523,N_29524,N_29525,N_29526,N_29527,N_29528,N_29529,N_29530,N_29531,N_29532,N_29533,N_29534,N_29535,N_29536,N_29537,N_29538,N_29539,N_29540,N_29541,N_29542,N_29543,N_29544,N_29545,N_29546,N_29547,N_29548,N_29549,N_29550,N_29551,N_29552,N_29553,N_29554,N_29555,N_29556,N_29557,N_29558,N_29559,N_29560,N_29561,N_29562,N_29563,N_29564,N_29565,N_29566,N_29567,N_29568,N_29569,N_29570,N_29571,N_29572,N_29573,N_29574,N_29575,N_29576,N_29577,N_29578,N_29579,N_29580,N_29581,N_29582,N_29583,N_29584,N_29585,N_29586,N_29587,N_29588,N_29589,N_29590,N_29591,N_29592,N_29593,N_29594,N_29595,N_29596,N_29597,N_29598,N_29599,N_29600,N_29601,N_29602,N_29603,N_29604,N_29605,N_29606,N_29607,N_29608,N_29609,N_29610,N_29611,N_29612,N_29613,N_29614,N_29615,N_29616,N_29617,N_29618,N_29619,N_29620,N_29621,N_29622,N_29623,N_29624,N_29625,N_29626,N_29627,N_29628,N_29629,N_29630,N_29631,N_29632,N_29633,N_29634,N_29635,N_29636,N_29637,N_29638,N_29639,N_29640,N_29641,N_29642,N_29643,N_29644,N_29645,N_29646,N_29647,N_29648,N_29649,N_29650,N_29651,N_29652,N_29653,N_29654,N_29655,N_29656,N_29657,N_29658,N_29659,N_29660,N_29661,N_29662,N_29663,N_29664,N_29665,N_29666,N_29667,N_29668,N_29669,N_29670,N_29671,N_29672,N_29673,N_29674,N_29675,N_29676,N_29677,N_29678,N_29679,N_29680,N_29681,N_29682,N_29683,N_29684,N_29685,N_29686,N_29687,N_29688,N_29689,N_29690,N_29691,N_29692,N_29693,N_29694,N_29695,N_29696,N_29697,N_29698,N_29699,N_29700,N_29701,N_29702,N_29703,N_29704,N_29705,N_29706,N_29707,N_29708,N_29709,N_29710,N_29711,N_29712,N_29713,N_29714,N_29715,N_29716,N_29717,N_29718,N_29719,N_29720,N_29721,N_29722,N_29723,N_29724,N_29725,N_29726,N_29727,N_29728,N_29729,N_29730,N_29731,N_29732,N_29733,N_29734,N_29735,N_29736,N_29737,N_29738,N_29739,N_29740,N_29741,N_29742,N_29743,N_29744,N_29745,N_29746,N_29747,N_29748,N_29749,N_29750,N_29751,N_29752,N_29753,N_29754,N_29755,N_29756,N_29757,N_29758,N_29759,N_29760,N_29761,N_29762,N_29763,N_29764,N_29765,N_29766,N_29767,N_29768,N_29769,N_29770,N_29771,N_29772,N_29773,N_29774,N_29775,N_29776,N_29777,N_29778,N_29779,N_29780,N_29781,N_29782,N_29783,N_29784,N_29785,N_29786,N_29787,N_29788,N_29789,N_29790,N_29791,N_29792,N_29793,N_29794,N_29795,N_29796,N_29797,N_29798,N_29799,N_29800,N_29801,N_29802,N_29803,N_29804,N_29805,N_29806,N_29807,N_29808,N_29809,N_29810,N_29811,N_29812,N_29813,N_29814,N_29815,N_29816,N_29817,N_29818,N_29819,N_29820,N_29821,N_29822,N_29823,N_29824,N_29825,N_29826,N_29827,N_29828,N_29829,N_29830,N_29831,N_29832,N_29833,N_29834,N_29835,N_29836,N_29837,N_29838,N_29839,N_29840,N_29841,N_29842,N_29843,N_29844,N_29845,N_29846,N_29847,N_29848,N_29849,N_29850,N_29851,N_29852,N_29853,N_29854,N_29855,N_29856,N_29857,N_29858,N_29859,N_29860,N_29861,N_29862,N_29863,N_29864,N_29865,N_29866,N_29867,N_29868,N_29869,N_29870,N_29871,N_29872,N_29873,N_29874,N_29875,N_29876,N_29877,N_29878,N_29879,N_29880,N_29881,N_29882,N_29883,N_29884,N_29885,N_29886,N_29887,N_29888,N_29889,N_29890,N_29891,N_29892,N_29893,N_29894,N_29895,N_29896,N_29897,N_29898,N_29899,N_29900,N_29901,N_29902,N_29903,N_29904,N_29905,N_29906,N_29907,N_29908,N_29909,N_29910,N_29911,N_29912,N_29913,N_29914,N_29915,N_29916,N_29917,N_29918,N_29919,N_29920,N_29921,N_29922,N_29923,N_29924,N_29925,N_29926,N_29927,N_29928,N_29929,N_29930,N_29931,N_29932,N_29933,N_29934,N_29935,N_29936,N_29937,N_29938,N_29939,N_29940,N_29941,N_29942,N_29943,N_29944,N_29945,N_29946,N_29947,N_29948,N_29949,N_29950,N_29951,N_29952,N_29953,N_29954,N_29955,N_29956,N_29957,N_29958,N_29959,N_29960,N_29961,N_29962,N_29963,N_29964,N_29965,N_29966,N_29967,N_29968,N_29969,N_29970,N_29971,N_29972,N_29973,N_29974,N_29975,N_29976,N_29977,N_29978,N_29979,N_29980,N_29981,N_29982,N_29983,N_29984,N_29985,N_29986,N_29987,N_29988,N_29989,N_29990,N_29991,N_29992,N_29993,N_29994,N_29995,N_29996,N_29997,N_29998,N_29999;
nand U0 (N_0,In_883,In_539);
nand U1 (N_1,In_2268,In_2422);
xnor U2 (N_2,In_1232,In_546);
or U3 (N_3,In_379,In_863);
nand U4 (N_4,In_2486,In_669);
xnor U5 (N_5,In_467,In_1723);
xnor U6 (N_6,In_268,In_2820);
and U7 (N_7,In_2765,In_400);
or U8 (N_8,In_493,In_2750);
nand U9 (N_9,In_1687,In_181);
or U10 (N_10,In_413,In_341);
and U11 (N_11,In_874,In_2383);
and U12 (N_12,In_1424,In_621);
nor U13 (N_13,In_1043,In_1944);
nand U14 (N_14,In_208,In_2842);
or U15 (N_15,In_2870,In_497);
or U16 (N_16,In_2535,In_2651);
or U17 (N_17,In_1906,In_2231);
nor U18 (N_18,In_1725,In_943);
and U19 (N_19,In_584,In_1600);
or U20 (N_20,In_1006,In_1577);
or U21 (N_21,In_1486,In_24);
or U22 (N_22,In_1970,In_76);
nand U23 (N_23,In_2304,In_2663);
nand U24 (N_24,In_897,In_2796);
xor U25 (N_25,In_123,In_1870);
or U26 (N_26,In_423,In_372);
and U27 (N_27,In_622,In_1613);
nor U28 (N_28,In_1416,In_2472);
or U29 (N_29,In_2114,In_248);
xnor U30 (N_30,In_2584,In_14);
nor U31 (N_31,In_2794,In_8);
or U32 (N_32,In_1352,In_762);
nand U33 (N_33,In_1058,In_798);
nor U34 (N_34,In_211,In_1088);
or U35 (N_35,In_2825,In_2060);
nor U36 (N_36,In_905,In_2602);
nand U37 (N_37,In_1858,In_752);
nand U38 (N_38,In_2484,In_1897);
or U39 (N_39,In_418,In_837);
nor U40 (N_40,In_1543,In_2139);
nand U41 (N_41,In_2416,In_2840);
and U42 (N_42,In_2993,In_1339);
xor U43 (N_43,In_280,In_1143);
and U44 (N_44,In_957,In_1489);
nor U45 (N_45,In_647,In_1718);
or U46 (N_46,In_1239,In_1810);
xnor U47 (N_47,In_1535,In_242);
xor U48 (N_48,In_911,In_2297);
and U49 (N_49,In_2145,In_2889);
nor U50 (N_50,In_1082,In_2434);
xnor U51 (N_51,In_2021,In_1555);
nor U52 (N_52,In_756,In_187);
nand U53 (N_53,In_2996,In_755);
and U54 (N_54,In_2051,In_1634);
nor U55 (N_55,In_1010,In_1562);
xor U56 (N_56,In_558,In_54);
nor U57 (N_57,In_742,In_816);
and U58 (N_58,In_2625,In_2182);
nand U59 (N_59,In_2927,In_2401);
xor U60 (N_60,In_1198,In_1672);
and U61 (N_61,In_70,In_2864);
xnor U62 (N_62,In_1698,In_1031);
nor U63 (N_63,In_1981,In_2575);
and U64 (N_64,In_420,In_1520);
nor U65 (N_65,In_1961,In_679);
xnor U66 (N_66,In_488,In_1479);
or U67 (N_67,In_1952,In_2705);
nand U68 (N_68,In_1709,In_946);
nor U69 (N_69,In_1265,In_968);
or U70 (N_70,In_2862,In_2379);
and U71 (N_71,In_78,In_2546);
or U72 (N_72,In_2679,In_2184);
nor U73 (N_73,In_1472,In_1840);
nor U74 (N_74,In_250,In_1697);
xor U75 (N_75,In_2099,In_786);
and U76 (N_76,In_1115,In_2799);
and U77 (N_77,In_514,In_2874);
xnor U78 (N_78,In_2487,In_655);
nor U79 (N_79,In_430,In_599);
nand U80 (N_80,In_274,In_2450);
nand U81 (N_81,In_1392,In_2776);
nand U82 (N_82,In_2746,In_486);
nor U83 (N_83,In_1298,In_1151);
and U84 (N_84,In_363,In_543);
nand U85 (N_85,In_1550,In_1735);
or U86 (N_86,In_2078,In_1018);
nand U87 (N_87,In_2210,In_2042);
or U88 (N_88,In_1774,In_1051);
and U89 (N_89,In_2667,In_2312);
xnor U90 (N_90,In_1074,In_1131);
nor U91 (N_91,In_2220,In_1533);
and U92 (N_92,In_2175,In_2665);
and U93 (N_93,In_1238,In_650);
and U94 (N_94,In_983,In_595);
and U95 (N_95,In_2859,In_1386);
or U96 (N_96,In_1935,In_2744);
or U97 (N_97,In_2346,In_2565);
nor U98 (N_98,In_2218,In_1077);
nand U99 (N_99,In_2463,In_1449);
nor U100 (N_100,In_240,In_2160);
xnor U101 (N_101,In_2639,In_690);
or U102 (N_102,In_577,In_2208);
and U103 (N_103,In_585,In_1327);
and U104 (N_104,In_1004,In_1693);
nor U105 (N_105,In_1427,In_2691);
nor U106 (N_106,In_900,In_2000);
and U107 (N_107,In_1442,In_619);
and U108 (N_108,In_2465,In_990);
nor U109 (N_109,In_2038,In_2787);
nor U110 (N_110,In_1569,In_698);
xor U111 (N_111,In_1932,In_2154);
xnor U112 (N_112,In_1263,In_2480);
nor U113 (N_113,In_1734,In_1595);
and U114 (N_114,In_1341,In_1225);
or U115 (N_115,In_589,In_1450);
nor U116 (N_116,In_2935,In_1623);
or U117 (N_117,In_1355,In_2683);
nor U118 (N_118,In_2396,In_2795);
nand U119 (N_119,In_1590,In_1170);
and U120 (N_120,In_2543,In_1605);
nor U121 (N_121,In_176,In_1256);
xnor U122 (N_122,In_2556,In_228);
xnor U123 (N_123,In_727,In_263);
nand U124 (N_124,In_1254,In_2590);
or U125 (N_125,In_1181,In_116);
or U126 (N_126,In_106,In_399);
or U127 (N_127,In_2557,In_457);
xnor U128 (N_128,In_1173,In_2479);
nand U129 (N_129,In_1506,In_2293);
or U130 (N_130,In_197,In_1525);
xnor U131 (N_131,In_2646,In_1586);
and U132 (N_132,In_2959,In_2939);
nor U133 (N_133,In_2421,In_866);
and U134 (N_134,In_1731,In_719);
nand U135 (N_135,In_1856,In_454);
xnor U136 (N_136,In_1484,In_2295);
and U137 (N_137,In_358,In_2248);
and U138 (N_138,In_328,In_1237);
or U139 (N_139,In_829,In_2868);
nor U140 (N_140,In_1843,In_1946);
and U141 (N_141,In_233,In_1596);
and U142 (N_142,In_2934,In_2355);
nand U143 (N_143,In_1971,In_2497);
nand U144 (N_144,In_1191,In_2132);
or U145 (N_145,In_2867,In_1368);
or U146 (N_146,In_1124,In_1868);
or U147 (N_147,In_2211,In_1408);
xor U148 (N_148,In_537,In_1350);
and U149 (N_149,In_2599,In_805);
xnor U150 (N_150,In_1656,In_2332);
nor U151 (N_151,In_2455,In_80);
xor U152 (N_152,In_823,In_2014);
nor U153 (N_153,In_1787,In_2334);
nand U154 (N_154,In_1455,In_1948);
xor U155 (N_155,In_1029,In_1854);
or U156 (N_156,In_1065,In_88);
or U157 (N_157,In_620,In_1813);
nand U158 (N_158,In_2398,In_583);
nor U159 (N_159,In_230,In_2013);
and U160 (N_160,In_136,In_804);
xnor U161 (N_161,In_27,In_1460);
or U162 (N_162,In_2901,In_1193);
nand U163 (N_163,In_521,In_1013);
and U164 (N_164,In_2707,In_1876);
or U165 (N_165,In_933,In_2107);
nand U166 (N_166,In_442,In_353);
or U167 (N_167,In_383,In_2659);
or U168 (N_168,In_12,In_1487);
nor U169 (N_169,In_2294,In_434);
nand U170 (N_170,In_62,In_1554);
nand U171 (N_171,In_167,In_2884);
nand U172 (N_172,In_1669,In_1997);
and U173 (N_173,In_1273,In_177);
nand U174 (N_174,In_641,In_17);
and U175 (N_175,In_1844,In_2485);
nand U176 (N_176,In_2680,In_182);
nor U177 (N_177,In_2101,In_1281);
xor U178 (N_178,In_2581,In_1675);
and U179 (N_179,In_2923,In_2843);
nand U180 (N_180,In_1502,In_1199);
or U181 (N_181,In_580,In_879);
or U182 (N_182,In_672,In_979);
nand U183 (N_183,In_1452,In_374);
xnor U184 (N_184,In_2028,In_544);
or U185 (N_185,In_1429,In_474);
nand U186 (N_186,In_1098,In_724);
nand U187 (N_187,In_212,In_485);
and U188 (N_188,In_186,In_225);
nor U189 (N_189,In_2756,In_936);
nand U190 (N_190,In_601,In_2399);
or U191 (N_191,In_1433,In_157);
xor U192 (N_192,In_1766,In_404);
and U193 (N_193,In_2635,In_1169);
nor U194 (N_194,In_627,In_787);
nor U195 (N_195,In_1523,In_1793);
nand U196 (N_196,In_711,In_1838);
or U197 (N_197,In_376,In_728);
nor U198 (N_198,In_2306,In_1706);
nor U199 (N_199,In_1957,In_1207);
or U200 (N_200,In_2991,In_1791);
or U201 (N_201,In_1304,In_291);
nor U202 (N_202,In_2394,In_1602);
or U203 (N_203,In_2637,In_209);
nand U204 (N_204,In_2035,In_677);
or U205 (N_205,In_2405,In_576);
and U206 (N_206,In_624,In_1309);
nor U207 (N_207,In_2029,In_2922);
and U208 (N_208,In_2109,In_2273);
nor U209 (N_209,In_2549,In_403);
and U210 (N_210,In_648,In_2092);
nand U211 (N_211,In_2104,In_1837);
and U212 (N_212,In_2747,In_644);
and U213 (N_213,In_1365,In_1943);
nand U214 (N_214,In_820,In_1756);
xor U215 (N_215,In_143,In_825);
or U216 (N_216,In_1260,In_381);
nor U217 (N_217,In_2678,In_30);
nand U218 (N_218,In_2327,In_1319);
or U219 (N_219,In_2841,In_1641);
or U220 (N_220,In_1741,In_2652);
or U221 (N_221,In_315,In_875);
nand U222 (N_222,In_2685,In_155);
or U223 (N_223,In_2284,In_2658);
nand U224 (N_224,In_1026,In_2677);
nand U225 (N_225,In_984,In_2246);
xnor U226 (N_226,In_960,In_963);
or U227 (N_227,In_952,In_1720);
xor U228 (N_228,In_135,In_708);
nor U229 (N_229,In_1839,In_1528);
or U230 (N_230,In_2681,In_587);
nand U231 (N_231,In_2880,In_1089);
nand U232 (N_232,In_1768,In_1348);
and U233 (N_233,In_1616,In_1511);
xnor U234 (N_234,In_759,In_2987);
and U235 (N_235,In_1405,In_1308);
or U236 (N_236,In_2969,In_1855);
nand U237 (N_237,In_44,In_562);
or U238 (N_238,In_16,In_2122);
and U239 (N_239,In_1120,In_331);
or U240 (N_240,In_1829,In_226);
and U241 (N_241,In_1123,In_1517);
nor U242 (N_242,In_2505,In_1568);
nor U243 (N_243,In_1537,In_2283);
nor U244 (N_244,In_516,In_1476);
xnor U245 (N_245,In_1188,In_777);
xnor U246 (N_246,In_34,In_1174);
xor U247 (N_247,In_1885,In_1908);
nor U248 (N_248,In_2568,In_2482);
and U249 (N_249,In_929,In_1257);
and U250 (N_250,In_718,In_2168);
and U251 (N_251,In_2238,In_1028);
and U252 (N_252,In_1708,In_2279);
xnor U253 (N_253,In_552,In_1775);
nand U254 (N_254,In_1160,In_2261);
and U255 (N_255,In_2162,In_678);
xor U256 (N_256,In_2203,In_792);
and U257 (N_257,In_1510,In_2826);
nand U258 (N_258,In_2061,In_2081);
and U259 (N_259,In_2320,In_2457);
nand U260 (N_260,In_801,In_1445);
nand U261 (N_261,In_2858,In_466);
or U262 (N_262,In_2117,In_687);
nand U263 (N_263,In_1584,In_2588);
xor U264 (N_264,In_958,In_163);
and U265 (N_265,In_1384,In_1134);
and U266 (N_266,In_462,In_389);
nor U267 (N_267,In_2266,In_239);
and U268 (N_268,In_244,In_2366);
or U269 (N_269,In_1048,In_2442);
and U270 (N_270,In_2003,In_2286);
nand U271 (N_271,In_661,In_1473);
nand U272 (N_272,In_2740,In_2302);
and U273 (N_273,In_2587,In_204);
or U274 (N_274,In_2098,In_85);
nand U275 (N_275,In_2962,In_1094);
and U276 (N_276,In_317,In_2566);
and U277 (N_277,In_2687,In_579);
and U278 (N_278,In_1955,In_2360);
nand U279 (N_279,In_1575,In_956);
or U280 (N_280,In_858,In_1333);
nand U281 (N_281,In_1694,In_2361);
xor U282 (N_282,In_1719,In_2538);
and U283 (N_283,In_2447,In_667);
or U284 (N_284,In_1567,In_219);
and U285 (N_285,In_1748,In_818);
xor U286 (N_286,In_723,In_1607);
or U287 (N_287,In_1608,In_1390);
and U288 (N_288,In_651,In_2020);
or U289 (N_289,In_169,In_1326);
xnor U290 (N_290,In_64,In_789);
and U291 (N_291,In_2812,In_1905);
nor U292 (N_292,In_1385,In_588);
nand U293 (N_293,In_2749,In_1673);
xnor U294 (N_294,In_2780,In_977);
or U295 (N_295,In_2140,In_1772);
or U296 (N_296,In_2885,In_2941);
nand U297 (N_297,In_939,In_2569);
or U298 (N_298,In_2965,In_32);
nand U299 (N_299,In_194,In_2328);
xor U300 (N_300,In_2159,In_784);
and U301 (N_301,In_1356,In_2836);
or U302 (N_302,In_937,In_1682);
and U303 (N_303,In_782,In_284);
and U304 (N_304,In_2783,In_2633);
nor U305 (N_305,In_709,In_2449);
nand U306 (N_306,In_1823,In_1132);
xnor U307 (N_307,In_140,In_1372);
and U308 (N_308,In_1846,In_1996);
xor U309 (N_309,In_1990,In_1165);
nor U310 (N_310,In_2483,In_1505);
and U311 (N_311,In_2904,In_498);
xnor U312 (N_312,In_2298,In_1627);
nor U313 (N_313,In_1729,In_2269);
xor U314 (N_314,In_112,In_2490);
or U315 (N_315,In_1526,In_691);
nor U316 (N_316,In_2108,In_247);
nor U317 (N_317,In_326,In_2477);
or U318 (N_318,In_995,In_355);
nor U319 (N_319,In_1796,In_1979);
nor U320 (N_320,In_1660,In_2015);
xnor U321 (N_321,In_2164,In_1338);
nor U322 (N_322,In_2254,In_2044);
nor U323 (N_323,In_2761,In_571);
nor U324 (N_324,In_1745,In_1508);
and U325 (N_325,In_2392,In_2771);
xor U326 (N_326,In_1572,In_2630);
or U327 (N_327,In_53,In_2572);
and U328 (N_328,In_1847,In_1030);
or U329 (N_329,In_1114,In_2811);
and U330 (N_330,In_556,In_22);
xor U331 (N_331,In_2614,In_561);
or U332 (N_332,In_2915,In_2900);
nand U333 (N_333,In_2171,In_2460);
nand U334 (N_334,In_1492,In_2032);
xnor U335 (N_335,In_2834,In_2785);
and U336 (N_336,In_1500,In_2609);
and U337 (N_337,In_1037,In_2781);
or U338 (N_338,In_151,In_1993);
nand U339 (N_339,In_468,In_1444);
and U340 (N_340,In_477,In_1279);
nor U341 (N_341,In_1481,In_2324);
and U342 (N_342,In_668,In_2069);
or U343 (N_343,In_2031,In_1202);
nor U344 (N_344,In_100,In_427);
nand U345 (N_345,In_1084,In_124);
nand U346 (N_346,In_1685,In_987);
or U347 (N_347,In_908,In_1597);
and U348 (N_348,In_103,In_2290);
or U349 (N_349,In_2561,In_2340);
and U350 (N_350,In_1253,In_722);
nor U351 (N_351,In_249,In_2608);
nor U352 (N_352,In_361,In_2512);
or U353 (N_353,In_2919,In_1069);
nor U354 (N_354,In_1918,In_127);
nand U355 (N_355,In_1835,In_594);
and U356 (N_356,In_2628,In_121);
nand U357 (N_357,In_452,In_200);
or U358 (N_358,In_1924,In_2530);
nand U359 (N_359,In_2045,In_2767);
or U360 (N_360,In_780,In_1559);
or U361 (N_361,In_1285,In_1397);
and U362 (N_362,In_689,In_1085);
and U363 (N_363,In_1293,In_1755);
and U364 (N_364,In_2562,In_1681);
nand U365 (N_365,In_94,In_405);
or U366 (N_366,In_3,In_417);
or U367 (N_367,In_414,In_227);
xnor U368 (N_368,In_1371,In_2196);
or U369 (N_369,In_2296,In_2773);
and U370 (N_370,In_508,In_702);
or U371 (N_371,In_241,In_881);
or U372 (N_372,In_1967,In_749);
nor U373 (N_373,In_659,In_581);
nand U374 (N_374,In_61,In_1210);
xnor U375 (N_375,In_1512,In_63);
or U376 (N_376,In_1610,In_2194);
xnor U377 (N_377,In_2034,In_1278);
nor U378 (N_378,In_2696,In_694);
or U379 (N_379,In_2445,In_710);
xnor U380 (N_380,In_2520,In_258);
xnor U381 (N_381,In_447,In_443);
xor U382 (N_382,In_653,In_596);
and U383 (N_383,In_2626,In_1644);
or U384 (N_384,In_134,In_2262);
nor U385 (N_385,In_2611,In_2470);
and U386 (N_386,In_2318,In_378);
xnor U387 (N_387,In_923,In_1176);
and U388 (N_388,In_2305,In_1332);
xnor U389 (N_389,In_2661,In_1343);
or U390 (N_390,In_2300,In_2133);
xnor U391 (N_391,In_604,In_2775);
nor U392 (N_392,In_2289,In_736);
or U393 (N_393,In_517,In_991);
and U394 (N_394,In_2339,In_1154);
nand U395 (N_395,In_2085,In_1035);
nor U396 (N_396,In_2183,In_269);
xnor U397 (N_397,In_25,In_2977);
nand U398 (N_398,In_2471,In_0);
or U399 (N_399,In_388,In_1201);
nor U400 (N_400,In_2720,In_2370);
and U401 (N_401,In_2835,In_1626);
nor U402 (N_402,In_2664,In_769);
nand U403 (N_403,In_1336,In_645);
xnor U404 (N_404,In_2105,In_1376);
or U405 (N_405,In_686,In_115);
nor U406 (N_406,In_1757,In_348);
xor U407 (N_407,In_2067,In_868);
or U408 (N_408,In_1515,In_2205);
or U409 (N_409,In_2423,In_629);
nor U410 (N_410,In_1782,In_2070);
nor U411 (N_411,In_2854,In_1142);
or U412 (N_412,In_6,In_191);
or U413 (N_413,In_1378,In_438);
nor U414 (N_414,In_2121,In_1387);
nand U415 (N_415,In_2754,In_766);
or U416 (N_416,In_2944,In_2335);
nor U417 (N_417,In_1138,In_440);
and U418 (N_418,In_1654,In_2219);
and U419 (N_419,In_1162,In_453);
and U420 (N_420,In_126,In_2610);
nor U421 (N_421,In_19,In_981);
xor U422 (N_422,In_2350,In_1581);
nand U423 (N_423,In_2452,In_1631);
xnor U424 (N_424,In_2188,In_2976);
or U425 (N_425,In_1779,In_1036);
nand U426 (N_426,In_843,In_1803);
and U427 (N_427,In_301,In_2973);
nor U428 (N_428,In_1300,In_2506);
nand U429 (N_429,In_2225,In_1916);
or U430 (N_430,In_1556,In_2563);
and U431 (N_431,In_2136,In_887);
nand U432 (N_432,In_2451,In_2612);
nand U433 (N_433,In_2997,In_2703);
and U434 (N_434,In_2752,In_273);
nor U435 (N_435,In_207,In_1262);
nor U436 (N_436,In_2251,In_410);
nand U437 (N_437,In_2719,In_2525);
nor U438 (N_438,In_2547,In_29);
nand U439 (N_439,In_873,In_696);
nor U440 (N_440,In_1310,In_2012);
nor U441 (N_441,In_202,In_2230);
and U442 (N_442,In_2435,In_2365);
xor U443 (N_443,In_2558,In_1765);
xnor U444 (N_444,In_2786,In_168);
xor U445 (N_445,In_429,In_2141);
xor U446 (N_446,In_2528,In_1686);
xor U447 (N_447,In_479,In_2242);
nand U448 (N_448,In_1195,In_2699);
or U449 (N_449,In_253,In_145);
xor U450 (N_450,In_2185,In_1877);
xnor U451 (N_451,In_628,In_449);
xnor U452 (N_452,In_132,In_743);
nor U453 (N_453,In_254,In_1743);
or U454 (N_454,In_1157,In_2701);
nand U455 (N_455,In_93,In_1324);
or U456 (N_456,In_520,In_1313);
nor U457 (N_457,In_2272,In_1244);
xnor U458 (N_458,In_2533,In_2545);
or U459 (N_459,In_1534,In_2966);
nor U460 (N_460,In_1842,In_2426);
nor U461 (N_461,In_573,In_2010);
xnor U462 (N_462,In_2291,In_643);
and U463 (N_463,In_1377,In_1561);
nor U464 (N_464,In_2734,In_1714);
nor U465 (N_465,In_2878,In_433);
and U466 (N_466,In_1146,In_1153);
xor U467 (N_467,In_892,In_1183);
or U468 (N_468,In_1306,In_1367);
and U469 (N_469,In_1546,In_862);
nor U470 (N_470,In_934,In_2191);
nand U471 (N_471,In_2409,In_2598);
and U472 (N_472,In_1620,In_1532);
and U473 (N_473,In_854,In_1495);
xor U474 (N_474,In_1073,In_1678);
xor U475 (N_475,In_2552,In_1934);
nand U476 (N_476,In_119,In_1483);
xnor U477 (N_477,In_1192,In_1354);
xor U478 (N_478,In_1507,In_1108);
and U479 (N_479,In_1099,In_2413);
xor U480 (N_480,In_2936,In_407);
nor U481 (N_481,In_65,In_338);
or U482 (N_482,In_1362,In_2810);
xnor U483 (N_483,In_701,In_2855);
xnor U484 (N_484,In_60,In_2515);
xor U485 (N_485,In_179,In_1812);
nand U486 (N_486,In_992,In_783);
nand U487 (N_487,In_1117,In_2690);
xnor U488 (N_488,In_424,In_138);
and U489 (N_489,In_2689,In_2055);
xor U490 (N_490,In_278,In_2620);
and U491 (N_491,In_1804,In_1025);
and U492 (N_492,In_534,In_482);
xnor U493 (N_493,In_349,In_1374);
nor U494 (N_494,In_1078,In_551);
nor U495 (N_495,In_794,In_2321);
xor U496 (N_496,In_20,In_831);
nand U497 (N_497,In_1914,In_2240);
and U498 (N_498,In_1217,In_512);
nand U499 (N_499,In_464,In_1054);
xor U500 (N_500,N_89,In_2621);
xor U501 (N_501,In_275,In_1439);
or U502 (N_502,In_2738,In_791);
and U503 (N_503,N_299,In_1499);
and U504 (N_504,In_907,In_847);
or U505 (N_505,In_1468,In_1055);
xor U506 (N_506,N_151,In_2745);
and U507 (N_507,In_1821,In_1235);
and U508 (N_508,In_2403,In_1825);
or U509 (N_509,In_2653,In_529);
nor U510 (N_510,N_168,In_2865);
xor U511 (N_511,In_2427,N_120);
nand U512 (N_512,In_803,In_120);
nand U513 (N_513,In_951,In_2271);
or U514 (N_514,N_49,In_332);
nor U515 (N_515,N_294,N_321);
and U516 (N_516,In_1539,In_2597);
xor U517 (N_517,N_156,N_436);
or U518 (N_518,N_426,In_768);
nand U519 (N_519,In_300,In_2096);
and U520 (N_520,N_478,In_1156);
and U521 (N_521,In_1629,In_2961);
nor U522 (N_522,In_685,In_193);
xnor U523 (N_523,In_210,In_1248);
nor U524 (N_524,In_2510,In_2500);
nand U525 (N_525,In_2195,In_55);
xnor U526 (N_526,In_2057,In_848);
nand U527 (N_527,In_928,N_131);
or U528 (N_528,In_90,In_2983);
xor U529 (N_529,In_58,In_2702);
nor U530 (N_530,In_1635,In_1251);
or U531 (N_531,In_1822,In_2116);
or U532 (N_532,In_704,In_2287);
and U533 (N_533,In_1815,In_1771);
and U534 (N_534,In_830,In_616);
nand U535 (N_535,In_445,In_1962);
nor U536 (N_536,In_190,In_2369);
or U537 (N_537,In_1353,In_352);
or U538 (N_538,In_2106,In_2071);
or U539 (N_539,In_2235,N_15);
and U540 (N_540,N_261,N_477);
and U541 (N_541,In_2424,N_468);
and U542 (N_542,N_486,N_334);
nor U543 (N_543,In_377,In_1925);
and U544 (N_544,In_969,In_634);
nor U545 (N_545,In_1466,In_1419);
and U546 (N_546,N_354,In_1360);
xnor U547 (N_547,In_2004,In_1802);
and U548 (N_548,In_428,In_500);
nor U549 (N_549,In_2234,In_2682);
xnor U550 (N_550,In_1865,In_139);
or U551 (N_551,In_2946,In_2036);
or U552 (N_552,In_633,In_256);
xnor U553 (N_553,In_184,In_1583);
xor U554 (N_554,In_156,In_199);
nor U555 (N_555,In_86,N_200);
and U556 (N_556,In_2669,In_384);
nand U557 (N_557,In_1521,In_2319);
nor U558 (N_558,N_377,In_370);
nor U559 (N_559,N_458,In_754);
nand U560 (N_560,In_1942,In_1215);
nand U561 (N_561,In_625,In_1783);
and U562 (N_562,In_2250,In_1987);
or U563 (N_563,In_2649,N_355);
and U564 (N_564,In_2419,In_684);
and U565 (N_565,In_2763,In_1598);
or U566 (N_566,In_1194,In_259);
or U567 (N_567,N_254,N_116);
and U568 (N_568,In_1513,In_2894);
nand U569 (N_569,In_510,In_2536);
and U570 (N_570,In_1242,In_2064);
nor U571 (N_571,In_114,N_253);
or U572 (N_572,N_337,In_1977);
and U573 (N_573,In_860,In_470);
nand U574 (N_574,In_1409,N_66);
and U575 (N_575,In_891,N_136);
xnor U576 (N_576,In_2807,In_2115);
nor U577 (N_577,N_446,In_2458);
nor U578 (N_578,N_3,In_2087);
xor U579 (N_579,In_2925,N_218);
or U580 (N_580,N_245,N_194);
nor U581 (N_581,N_98,In_2493);
nand U582 (N_582,In_1860,In_901);
and U583 (N_583,In_2345,In_1083);
nor U584 (N_584,In_1063,In_906);
or U585 (N_585,In_1224,N_118);
nor U586 (N_586,In_72,In_1022);
and U587 (N_587,In_554,In_1648);
nor U588 (N_588,In_255,In_896);
and U589 (N_589,In_1529,In_2349);
nand U590 (N_590,In_42,In_95);
nor U591 (N_591,In_1992,In_1410);
xnor U592 (N_592,N_224,In_2876);
nand U593 (N_593,In_597,In_1882);
xnor U594 (N_594,In_1894,In_2544);
and U595 (N_595,In_1266,In_2461);
xnor U596 (N_596,In_1928,N_431);
nor U597 (N_597,In_1403,In_175);
xnor U598 (N_598,In_2241,N_52);
nor U599 (N_599,In_1430,In_380);
xor U600 (N_600,In_2352,In_2692);
nor U601 (N_601,In_1845,N_128);
or U602 (N_602,In_1570,In_1394);
nor U603 (N_603,In_1465,In_266);
nor U604 (N_604,N_217,N_225);
nor U605 (N_605,In_771,In_2624);
nand U606 (N_606,In_2887,In_2006);
nor U607 (N_607,In_344,In_1436);
nor U608 (N_608,In_1323,In_2337);
or U609 (N_609,In_2088,In_737);
nor U610 (N_610,N_357,N_155);
or U611 (N_611,In_2638,In_133);
xnor U612 (N_612,N_306,In_834);
xnor U613 (N_613,In_994,In_288);
and U614 (N_614,In_1895,In_2607);
and U615 (N_615,N_130,In_2429);
or U616 (N_616,In_2888,In_721);
and U617 (N_617,In_1703,In_1347);
nor U618 (N_618,In_2524,In_2722);
and U619 (N_619,In_183,In_2079);
or U620 (N_620,In_2930,In_304);
xnor U621 (N_621,In_2198,In_945);
or U622 (N_622,N_343,In_2260);
nor U623 (N_623,N_432,In_2438);
and U624 (N_624,In_638,N_315);
and U625 (N_625,In_1320,In_2743);
and U626 (N_626,In_1695,In_2605);
and U627 (N_627,In_469,In_828);
or U628 (N_628,In_231,N_308);
or U629 (N_629,In_2972,In_2489);
or U630 (N_630,In_800,In_1956);
nor U631 (N_631,In_1621,In_2281);
and U632 (N_632,In_2292,In_335);
nor U633 (N_633,In_1276,In_1884);
or U634 (N_634,In_1639,In_744);
xnor U635 (N_635,In_2189,In_2778);
xnor U636 (N_636,In_1968,In_1663);
and U637 (N_637,In_1064,In_1042);
and U638 (N_638,In_2947,In_826);
nor U639 (N_639,In_1459,In_2072);
nand U640 (N_640,In_1302,In_2772);
nor U641 (N_641,In_2094,In_674);
xor U642 (N_642,In_2984,N_192);
or U643 (N_643,In_1363,In_997);
nand U644 (N_644,In_333,N_67);
and U645 (N_645,N_380,In_2267);
nand U646 (N_646,In_1361,In_195);
or U647 (N_647,In_2571,N_262);
nand U648 (N_648,In_2886,In_2697);
and U649 (N_649,In_1417,N_25);
and U650 (N_650,In_2918,In_1679);
xor U651 (N_651,In_2131,N_496);
and U652 (N_652,In_327,In_639);
xor U653 (N_653,In_444,In_745);
nand U654 (N_654,In_2908,In_998);
nand U655 (N_655,N_366,In_476);
nand U656 (N_656,In_1172,In_2570);
and U657 (N_657,In_1612,In_1880);
or U658 (N_658,In_2706,N_102);
xnor U659 (N_659,In_2950,N_23);
and U660 (N_660,In_913,In_1951);
nor U661 (N_661,In_2668,In_215);
nand U662 (N_662,In_1402,In_851);
or U663 (N_663,N_148,In_1834);
and U664 (N_664,In_2049,In_40);
nor U665 (N_665,In_671,In_1456);
and U666 (N_666,N_454,In_137);
or U667 (N_667,N_46,In_652);
xnor U668 (N_668,N_85,In_1305);
nand U669 (N_669,In_2343,N_345);
xnor U670 (N_670,In_2798,In_1231);
xor U671 (N_671,N_384,In_1830);
nor U672 (N_672,N_179,In_764);
and U673 (N_673,In_1190,In_122);
xor U674 (N_674,In_1715,In_2943);
and U675 (N_675,In_2808,In_2736);
and U676 (N_676,In_2671,N_169);
nand U677 (N_677,In_56,N_167);
nor U678 (N_678,N_140,In_2002);
and U679 (N_679,N_427,In_2619);
xnor U680 (N_680,In_1662,In_2232);
nor U681 (N_681,In_2209,In_1874);
or U682 (N_682,N_138,In_2187);
and U683 (N_683,In_2929,In_141);
nand U684 (N_684,In_2542,In_525);
xnor U685 (N_685,In_1959,In_2879);
and U686 (N_686,In_2911,In_173);
xnor U687 (N_687,In_2481,N_100);
and U688 (N_688,In_885,N_434);
xor U689 (N_689,N_406,In_92);
nor U690 (N_690,In_2285,N_215);
nor U691 (N_691,N_170,In_1746);
or U692 (N_692,In_2567,In_2440);
xnor U693 (N_693,In_2730,In_1008);
nor U694 (N_694,In_1593,In_229);
nor U695 (N_695,In_841,In_2165);
xnor U696 (N_696,In_1448,In_2555);
nand U697 (N_697,N_103,In_1701);
nor U698 (N_698,In_695,In_1057);
nor U699 (N_699,In_1121,In_739);
nor U700 (N_700,In_2553,In_2666);
or U701 (N_701,In_1617,N_448);
xnor U702 (N_702,N_257,N_227);
and U703 (N_703,In_2980,N_74);
nand U704 (N_704,In_1711,In_1047);
xnor U705 (N_705,In_1949,In_1118);
xnor U706 (N_706,In_2532,In_626);
or U707 (N_707,N_92,In_1294);
xnor U708 (N_708,In_2243,In_1817);
or U709 (N_709,In_1015,In_1137);
xor U710 (N_710,In_125,N_247);
and U711 (N_711,In_1184,In_2397);
nand U712 (N_712,In_509,In_970);
nor U713 (N_713,In_2388,In_2153);
nand U714 (N_714,In_2877,In_1125);
and U715 (N_715,In_82,In_1808);
and U716 (N_716,In_2527,In_1475);
nor U717 (N_717,In_1382,In_1680);
xor U718 (N_718,N_236,In_2945);
and U719 (N_719,In_761,In_2149);
xor U720 (N_720,In_2577,In_357);
xnor U721 (N_721,N_183,In_2274);
nand U722 (N_722,In_2456,In_528);
and U723 (N_723,N_444,In_1328);
nor U724 (N_724,In_1886,In_523);
nand U725 (N_725,In_1609,In_334);
nor U726 (N_726,In_809,In_1632);
nor U727 (N_727,In_1241,In_2475);
nor U728 (N_728,In_555,In_2406);
nor U729 (N_729,In_2540,In_2647);
and U730 (N_730,In_1234,In_2642);
xor U731 (N_731,In_1790,In_1989);
nand U732 (N_732,N_125,In_2953);
xnor U733 (N_733,N_490,In_1530);
or U734 (N_734,In_1288,In_1721);
nand U735 (N_735,In_1464,In_2871);
xnor U736 (N_736,In_1040,N_199);
and U737 (N_737,In_1828,In_910);
nand U738 (N_738,N_87,In_1689);
or U739 (N_739,N_346,In_2790);
nor U740 (N_740,In_959,In_2508);
nor U741 (N_741,N_229,N_175);
nor U742 (N_742,In_770,In_69);
or U743 (N_743,In_307,In_2342);
xnor U744 (N_744,In_2819,In_2716);
and U745 (N_745,In_2522,In_395);
nand U746 (N_746,N_383,N_86);
xor U747 (N_747,In_757,In_2338);
xor U748 (N_748,In_1930,N_212);
nor U749 (N_749,In_271,In_499);
or U750 (N_750,In_1767,In_1197);
nand U751 (N_751,In_2464,In_31);
xor U752 (N_752,In_1152,In_1426);
or U753 (N_753,In_1491,In_1863);
and U754 (N_754,In_1862,In_1751);
nor U755 (N_755,N_72,N_1);
or U756 (N_756,N_437,In_2823);
xor U757 (N_757,In_2382,N_99);
and U758 (N_758,N_272,In_775);
nand U759 (N_759,In_2933,In_1220);
or U760 (N_760,In_463,In_2018);
and U761 (N_761,In_1007,In_1140);
or U762 (N_762,In_2112,In_1655);
nor U763 (N_763,In_2981,In_682);
xor U764 (N_764,In_1522,In_1833);
and U765 (N_765,In_1133,In_2123);
or U766 (N_766,In_1696,In_257);
xnor U767 (N_767,In_1806,In_832);
xor U768 (N_768,In_2412,In_864);
nor U769 (N_769,In_1096,In_1518);
xor U770 (N_770,In_2120,N_484);
nand U771 (N_771,N_325,In_1155);
nor U772 (N_772,In_1691,In_1312);
or U773 (N_773,In_2709,In_1226);
or U774 (N_774,In_2102,In_819);
or U775 (N_775,N_145,In_1400);
nor U776 (N_776,In_2845,In_1204);
nor U777 (N_777,N_195,In_1003);
or U778 (N_778,In_2662,In_1318);
nor U779 (N_779,In_1728,In_1831);
or U780 (N_780,In_435,In_2921);
and U781 (N_781,In_2124,N_126);
and U782 (N_782,In_1297,In_2755);
nand U783 (N_783,In_2978,In_437);
and U784 (N_784,In_2554,In_2033);
xor U785 (N_785,In_2968,In_1167);
and U786 (N_786,In_1773,In_919);
and U787 (N_787,N_230,In_631);
and U788 (N_788,In_912,N_54);
and U789 (N_789,In_986,In_615);
nor U790 (N_790,N_365,In_1322);
or U791 (N_791,In_2573,N_360);
or U792 (N_792,In_646,In_1650);
nand U793 (N_793,In_1212,In_113);
nand U794 (N_794,In_950,In_882);
and U795 (N_795,In_2322,In_776);
or U796 (N_796,In_2462,In_217);
nand U797 (N_797,In_1582,In_101);
or U798 (N_798,N_356,N_470);
xnor U799 (N_799,In_2129,In_2167);
and U800 (N_800,In_1814,N_240);
nor U801 (N_801,In_846,In_39);
or U802 (N_802,N_48,In_2916);
and U803 (N_803,In_2158,In_2068);
and U804 (N_804,In_1425,In_2444);
nand U805 (N_805,In_1984,In_166);
or U806 (N_806,N_320,N_163);
nor U807 (N_807,N_259,In_1750);
nor U808 (N_808,In_415,N_266);
and U809 (N_809,In_2062,In_2155);
xor U810 (N_810,N_488,In_2430);
xnor U811 (N_811,In_2970,In_808);
nor U812 (N_812,In_147,In_1255);
nor U813 (N_813,In_1280,In_1872);
and U814 (N_814,In_2791,In_2368);
nor U815 (N_815,In_2084,In_2377);
nand U816 (N_816,In_1820,N_71);
or U817 (N_817,In_1447,In_2711);
or U818 (N_818,In_1451,N_107);
and U819 (N_819,In_1800,In_2008);
nand U820 (N_820,In_339,In_1075);
nor U821 (N_821,N_425,In_471);
xnor U822 (N_822,N_137,In_2513);
nand U823 (N_823,In_48,In_856);
nand U824 (N_824,In_28,In_1861);
nor U825 (N_825,In_2309,N_361);
and U826 (N_826,In_2509,In_2178);
nand U827 (N_827,In_975,In_2618);
nor U828 (N_828,In_2769,In_1936);
xnor U829 (N_829,N_302,N_497);
or U830 (N_830,In_366,In_289);
nor U831 (N_831,In_2491,In_1275);
nor U832 (N_832,In_1614,N_322);
or U833 (N_833,N_364,In_716);
nand U834 (N_834,In_2906,In_2849);
nor U835 (N_835,In_2710,In_1072);
nor U836 (N_836,In_1141,In_41);
xor U837 (N_837,In_2134,In_1722);
and U838 (N_838,In_2860,In_2244);
or U839 (N_839,In_490,N_378);
nand U840 (N_840,In_2645,In_2259);
nand U841 (N_841,In_460,In_2764);
nor U842 (N_842,N_221,In_1739);
xnor U843 (N_843,In_385,In_2063);
xnor U844 (N_844,In_2731,In_2170);
nor U845 (N_845,In_111,In_1001);
and U846 (N_846,In_1090,In_973);
xor U847 (N_847,In_441,In_2579);
xor U848 (N_848,In_267,N_207);
nor U849 (N_849,In_1653,In_1816);
xnor U850 (N_850,In_1482,In_2214);
xnor U851 (N_851,In_1527,N_150);
and U852 (N_852,In_2019,In_1881);
nand U853 (N_853,In_396,In_1818);
nand U854 (N_854,In_222,N_237);
nor U855 (N_855,In_916,In_1911);
and U856 (N_856,In_1295,In_1878);
nor U857 (N_857,In_2420,In_1763);
xor U858 (N_858,In_2,In_386);
nand U859 (N_859,In_1222,In_2725);
xnor U860 (N_860,In_2931,N_187);
xor U861 (N_861,In_1578,In_732);
nand U862 (N_862,In_419,N_55);
or U863 (N_863,In_2529,In_375);
and U864 (N_864,In_649,In_286);
xnor U865 (N_865,N_326,In_2174);
nand U866 (N_866,In_1041,In_246);
or U867 (N_867,In_822,In_1164);
and U868 (N_868,In_1432,N_115);
and U869 (N_869,In_2822,In_515);
or U870 (N_870,In_746,In_2837);
nor U871 (N_871,In_37,In_2400);
nand U872 (N_872,In_329,N_491);
nor U873 (N_873,In_2957,In_1890);
nor U874 (N_874,In_675,N_290);
xnor U875 (N_875,In_224,In_402);
nor U876 (N_876,N_347,In_1434);
nor U877 (N_877,In_310,In_71);
nor U878 (N_878,In_2848,In_2616);
nand U879 (N_879,N_117,In_1712);
or U880 (N_880,In_1849,N_295);
xnor U881 (N_881,N_430,In_2110);
nand U882 (N_882,In_2125,In_533);
or U883 (N_883,In_2237,In_1736);
nand U884 (N_884,In_1317,In_43);
xnor U885 (N_885,N_61,In_1461);
xnor U886 (N_886,In_2631,In_2788);
nand U887 (N_887,In_1267,In_2829);
and U888 (N_888,N_39,In_1875);
or U889 (N_889,In_1428,In_1699);
nor U890 (N_890,In_1292,In_697);
xor U891 (N_891,In_2404,In_1401);
or U892 (N_892,In_213,In_7);
nand U893 (N_893,In_2082,In_2792);
xnor U894 (N_894,In_45,In_316);
nor U895 (N_895,N_463,In_741);
xor U896 (N_896,In_360,In_1548);
nand U897 (N_897,In_2362,In_2721);
or U898 (N_898,In_270,N_44);
and U899 (N_899,In_1732,In_1684);
nand U900 (N_900,In_564,In_2770);
or U901 (N_901,In_2833,In_1150);
and U902 (N_902,In_346,In_681);
or U903 (N_903,In_1642,In_221);
nand U904 (N_904,In_1045,N_202);
nor U905 (N_905,In_2896,In_1891);
nor U906 (N_906,N_42,In_609);
and U907 (N_907,In_642,In_2824);
or U908 (N_908,N_231,N_127);
or U909 (N_909,In_2774,In_884);
and U910 (N_910,In_2417,In_861);
nor U911 (N_911,In_412,N_190);
nor U912 (N_912,In_1446,N_439);
or U913 (N_913,In_2821,In_1435);
and U914 (N_914,In_2344,In_237);
and U915 (N_915,In_1549,In_1116);
or U916 (N_916,In_2228,In_390);
or U917 (N_917,In_921,In_1185);
nand U918 (N_918,In_1247,In_369);
nor U919 (N_919,N_41,In_773);
and U920 (N_920,N_392,In_2265);
and U921 (N_921,In_2437,In_2054);
and U922 (N_922,In_281,In_1805);
or U923 (N_923,In_726,In_1200);
and U924 (N_924,In_1252,In_59);
nor U925 (N_925,In_351,N_165);
xnor U926 (N_926,In_2233,In_2902);
nand U927 (N_927,N_402,In_607);
xnor U928 (N_928,In_1175,In_611);
nand U929 (N_929,N_88,In_557);
nor U930 (N_930,In_2733,In_1538);
nand U931 (N_931,In_2560,In_1463);
nor U932 (N_932,In_2166,In_2757);
and U933 (N_933,In_976,In_2518);
and U934 (N_934,In_522,In_1126);
or U935 (N_935,In_953,In_899);
nand U936 (N_936,In_2359,In_2698);
or U937 (N_937,In_2037,In_662);
nand U938 (N_938,In_1211,In_1603);
and U939 (N_939,In_1033,In_1848);
nand U940 (N_940,N_313,In_276);
and U941 (N_941,In_1396,N_59);
xor U942 (N_942,N_182,In_1781);
and U943 (N_943,N_58,In_153);
nand U944 (N_944,N_95,In_2592);
nor U945 (N_945,N_288,In_343);
nand U946 (N_946,In_2111,In_102);
xnor U947 (N_947,In_2391,N_435);
nand U948 (N_948,In_760,In_2151);
and U949 (N_949,In_1647,In_2156);
and U950 (N_950,In_2938,N_374);
or U951 (N_951,In_323,N_219);
nor U952 (N_952,In_2816,In_1415);
xnor U953 (N_953,In_944,N_451);
and U954 (N_954,In_2963,In_2007);
or U955 (N_955,In_87,In_2378);
or U956 (N_956,In_1315,In_2436);
xnor U957 (N_957,In_1758,N_271);
nand U958 (N_958,In_630,In_245);
xnor U959 (N_959,In_1139,In_104);
xor U960 (N_960,In_2866,N_493);
and U961 (N_961,In_2143,In_2531);
or U962 (N_962,In_1277,N_289);
and U963 (N_963,N_312,In_196);
nand U964 (N_964,In_2910,In_542);
or U965 (N_965,In_2955,In_1182);
nand U966 (N_966,N_319,In_2844);
nor U967 (N_967,In_1261,N_278);
nand U968 (N_968,In_382,In_778);
or U969 (N_969,In_2395,In_2053);
nand U970 (N_970,In_836,In_720);
nor U971 (N_971,In_2541,In_1661);
or U972 (N_972,In_2718,In_2999);
or U973 (N_973,N_388,In_1780);
xor U974 (N_974,N_396,N_363);
nor U975 (N_975,In_1062,In_2314);
nand U976 (N_976,In_2909,N_197);
nor U977 (N_977,In_109,In_13);
nand U978 (N_978,In_66,In_572);
xor U979 (N_979,In_1467,In_2025);
or U980 (N_980,In_1611,In_2142);
xnor U981 (N_981,N_393,In_793);
or U982 (N_982,In_785,In_320);
xor U983 (N_983,N_394,In_2591);
and U984 (N_984,In_293,N_164);
nand U985 (N_985,In_1664,In_364);
and U986 (N_986,In_2411,N_21);
or U987 (N_987,In_1504,In_1462);
or U988 (N_988,In_569,In_635);
nor U989 (N_989,In_1488,N_17);
and U990 (N_990,In_2768,In_898);
and U991 (N_991,In_940,In_2074);
and U992 (N_992,In_797,N_47);
or U993 (N_993,N_327,In_170);
or U994 (N_994,In_264,In_1913);
xnor U995 (N_995,In_2050,In_965);
and U996 (N_996,In_663,In_610);
nand U997 (N_997,In_2065,In_2043);
nand U998 (N_998,In_2459,In_1334);
xnor U999 (N_999,In_971,In_2086);
nand U1000 (N_1000,N_275,N_825);
or U1001 (N_1001,N_403,In_2223);
nor U1002 (N_1002,In_1591,In_593);
nor U1003 (N_1003,In_220,In_1344);
xor U1004 (N_1004,N_833,N_466);
xnor U1005 (N_1005,In_2971,In_1423);
nor U1006 (N_1006,In_833,In_252);
xnor U1007 (N_1007,In_2083,In_1437);
and U1008 (N_1008,In_2723,In_1494);
nor U1009 (N_1009,In_842,In_850);
xnor U1010 (N_1010,In_36,In_894);
and U1011 (N_1011,In_1346,N_241);
and U1012 (N_1012,In_2766,N_421);
xnor U1013 (N_1013,In_692,In_1019);
nand U1014 (N_1014,In_2347,N_538);
and U1015 (N_1015,In_172,In_2627);
nand U1016 (N_1016,N_869,In_654);
or U1017 (N_1017,In_2027,In_1643);
nand U1018 (N_1018,N_996,In_504);
nand U1019 (N_1019,In_1379,N_595);
nor U1020 (N_1020,N_416,N_832);
xor U1021 (N_1021,In_2920,In_2875);
nor U1022 (N_1022,In_15,In_2367);
nand U1023 (N_1023,N_296,N_968);
and U1024 (N_1024,N_691,In_2190);
and U1025 (N_1025,N_703,In_1187);
and U1026 (N_1026,In_47,In_2891);
or U1027 (N_1027,In_262,In_2478);
nor U1028 (N_1028,N_369,N_371);
nand U1029 (N_1029,In_2636,N_234);
xor U1030 (N_1030,In_2869,N_279);
nor U1031 (N_1031,N_688,In_549);
nor U1032 (N_1032,In_1588,In_670);
or U1033 (N_1033,In_2899,In_2372);
or U1034 (N_1034,N_153,In_806);
and U1035 (N_1035,In_1727,In_1027);
and U1036 (N_1036,In_446,N_82);
nor U1037 (N_1037,In_2517,In_853);
and U1038 (N_1038,N_452,In_1713);
xnor U1039 (N_1039,N_805,N_958);
and U1040 (N_1040,In_260,N_729);
nor U1041 (N_1041,N_983,N_63);
nor U1042 (N_1042,In_1303,In_2937);
and U1043 (N_1043,In_548,N_348);
nand U1044 (N_1044,N_238,In_1046);
xnor U1045 (N_1045,N_856,In_1585);
nand U1046 (N_1046,In_1784,In_356);
nand U1047 (N_1047,N_379,In_2494);
and U1048 (N_1048,In_1485,In_73);
nor U1049 (N_1049,N_176,In_1002);
nor U1050 (N_1050,In_2717,N_579);
nor U1051 (N_1051,In_1391,In_2307);
or U1052 (N_1052,N_594,In_1633);
and U1053 (N_1053,N_846,N_113);
nand U1054 (N_1054,N_526,In_23);
nand U1055 (N_1055,N_847,In_292);
nand U1056 (N_1056,In_2439,In_857);
xor U1057 (N_1057,In_2895,N_722);
nand U1058 (N_1058,N_62,In_2161);
nor U1059 (N_1059,N_791,N_18);
nor U1060 (N_1060,In_312,N_709);
nor U1061 (N_1061,In_130,In_2655);
nand U1062 (N_1062,In_2942,In_733);
or U1063 (N_1063,N_502,In_340);
nand U1064 (N_1064,N_536,In_2024);
xnor U1065 (N_1065,In_1982,In_2654);
nand U1066 (N_1066,In_67,N_11);
and U1067 (N_1067,N_500,In_203);
nand U1068 (N_1068,In_368,In_2928);
xor U1069 (N_1069,In_2476,In_2215);
xnor U1070 (N_1070,In_144,N_649);
and U1071 (N_1071,In_2351,N_521);
or U1072 (N_1072,In_1864,N_510);
or U1073 (N_1073,N_419,N_90);
or U1074 (N_1074,N_755,In_2075);
nor U1075 (N_1075,N_157,N_527);
xor U1076 (N_1076,In_1412,In_2726);
and U1077 (N_1077,In_656,In_2559);
nand U1078 (N_1078,In_2303,N_263);
and U1079 (N_1079,In_1726,In_1707);
nand U1080 (N_1080,In_387,In_1092);
nor U1081 (N_1081,In_1340,In_1544);
or U1082 (N_1082,N_789,In_2735);
nor U1083 (N_1083,In_1826,N_111);
or U1084 (N_1084,N_965,N_817);
xor U1085 (N_1085,In_2009,In_501);
and U1086 (N_1086,N_511,In_2389);
nand U1087 (N_1087,N_146,In_779);
and U1088 (N_1088,N_376,In_715);
nor U1089 (N_1089,N_945,N_152);
or U1090 (N_1090,N_756,N_820);
nand U1091 (N_1091,N_555,In_302);
nor U1092 (N_1092,N_710,In_1624);
or U1093 (N_1093,In_1744,In_1671);
and U1094 (N_1094,In_1514,In_397);
or U1095 (N_1095,N_777,In_680);
or U1096 (N_1096,In_904,In_827);
or U1097 (N_1097,In_1945,N_273);
xnor U1098 (N_1098,N_911,In_391);
nand U1099 (N_1099,In_2989,N_571);
and U1100 (N_1100,N_411,In_535);
nor U1101 (N_1101,N_973,In_1869);
nor U1102 (N_1102,N_404,In_2052);
and U1103 (N_1103,N_635,N_778);
nor U1104 (N_1104,In_1221,In_1);
and U1105 (N_1105,In_1272,In_734);
xor U1106 (N_1106,In_938,In_1061);
and U1107 (N_1107,In_1388,N_246);
nand U1108 (N_1108,In_1710,In_810);
or U1109 (N_1109,N_871,N_455);
xor U1110 (N_1110,In_2255,In_545);
nand U1111 (N_1111,In_840,N_947);
nor U1112 (N_1112,N_483,N_387);
xor U1113 (N_1113,In_730,In_313);
and U1114 (N_1114,N_12,In_297);
and U1115 (N_1115,In_282,In_519);
nor U1116 (N_1116,N_700,N_577);
xnor U1117 (N_1117,In_2473,In_1792);
xnor U1118 (N_1118,N_801,In_2954);
xnor U1119 (N_1119,In_1923,N_904);
and U1120 (N_1120,In_673,In_2407);
or U1121 (N_1121,N_792,In_159);
and U1122 (N_1122,N_5,In_2022);
nor U1123 (N_1123,N_912,In_472);
nor U1124 (N_1124,N_554,In_1674);
nand U1125 (N_1125,In_1366,N_556);
nor U1126 (N_1126,In_636,In_524);
nor U1127 (N_1127,N_839,N_819);
or U1128 (N_1128,N_6,In_2148);
and U1129 (N_1129,N_878,N_808);
nand U1130 (N_1130,In_2496,In_1974);
or U1131 (N_1131,In_1690,N_858);
or U1132 (N_1132,In_2138,N_32);
or U1133 (N_1133,In_1564,In_1651);
xor U1134 (N_1134,In_640,In_1068);
nand U1135 (N_1135,In_2348,In_2511);
nand U1136 (N_1136,In_2466,In_2245);
nor U1137 (N_1137,In_2615,N_821);
nand U1138 (N_1138,N_276,In_243);
nor U1139 (N_1139,N_665,In_632);
xor U1140 (N_1140,N_13,In_174);
or U1141 (N_1141,In_455,N_180);
nor U1142 (N_1142,In_2313,In_459);
or U1143 (N_1143,In_1853,N_260);
nor U1144 (N_1144,N_617,N_142);
or U1145 (N_1145,In_1670,In_2550);
xnor U1146 (N_1146,In_2325,In_688);
or U1147 (N_1147,In_1166,N_723);
nand U1148 (N_1148,In_2596,In_1186);
or U1149 (N_1149,In_2729,In_527);
and U1150 (N_1150,In_1630,N_204);
and U1151 (N_1151,In_1592,In_1103);
nand U1152 (N_1152,N_781,N_966);
nor U1153 (N_1153,N_865,N_797);
and U1154 (N_1154,In_2163,In_2595);
nand U1155 (N_1155,In_350,N_336);
xnor U1156 (N_1156,N_761,N_794);
nor U1157 (N_1157,In_2782,In_2830);
nor U1158 (N_1158,N_872,In_272);
and U1159 (N_1159,In_1364,N_413);
nor U1160 (N_1160,In_1819,N_563);
nor U1161 (N_1161,N_20,In_2172);
xor U1162 (N_1162,In_1794,N_964);
nor U1163 (N_1163,In_1851,N_34);
or U1164 (N_1164,In_10,In_345);
xor U1165 (N_1165,In_1329,N_311);
and U1166 (N_1166,In_2317,N_952);
or U1167 (N_1167,In_1941,In_1668);
nor U1168 (N_1168,N_70,In_1411);
or U1169 (N_1169,In_160,N_351);
xnor U1170 (N_1170,In_1677,In_261);
nor U1171 (N_1171,N_350,In_394);
or U1172 (N_1172,N_43,In_2213);
nor U1173 (N_1173,N_621,In_2576);
nor U1174 (N_1174,In_1938,In_406);
nand U1175 (N_1175,N_559,In_1753);
xnor U1176 (N_1176,In_1050,In_2224);
or U1177 (N_1177,In_1776,In_2186);
nor U1178 (N_1178,N_768,In_2192);
or U1179 (N_1179,N_757,In_2857);
and U1180 (N_1180,In_623,In_2872);
or U1181 (N_1181,N_735,N_990);
xnor U1182 (N_1182,N_711,In_1705);
xor U1183 (N_1183,In_1973,N_837);
nor U1184 (N_1184,N_506,In_774);
nand U1185 (N_1185,N_920,In_1223);
or U1186 (N_1186,N_372,In_1922);
and U1187 (N_1187,In_2640,In_1381);
nand U1188 (N_1188,In_1738,In_373);
xor U1189 (N_1189,N_84,N_677);
xor U1190 (N_1190,N_765,N_779);
and U1191 (N_1191,N_891,N_309);
or U1192 (N_1192,N_704,In_2995);
and U1193 (N_1193,In_964,N_575);
or U1194 (N_1194,In_2514,N_424);
xor U1195 (N_1195,In_2385,N_134);
nand U1196 (N_1196,In_1087,In_83);
and U1197 (N_1197,N_701,N_683);
and U1198 (N_1198,N_693,In_290);
nor U1199 (N_1199,N_73,N_407);
and U1200 (N_1200,N_739,In_336);
nand U1201 (N_1201,N_277,In_2041);
and U1202 (N_1202,In_1307,In_978);
nand U1203 (N_1203,N_876,In_570);
nand U1204 (N_1204,In_966,In_799);
or U1205 (N_1205,In_2748,N_890);
xnor U1206 (N_1206,N_518,In_1100);
or U1207 (N_1207,N_798,In_1516);
and U1208 (N_1208,In_890,N_589);
and U1209 (N_1209,In_617,N_612);
and U1210 (N_1210,N_251,In_815);
nor U1211 (N_1211,In_2898,N_606);
and U1212 (N_1212,In_559,In_2089);
xnor U1213 (N_1213,In_1245,In_2393);
nor U1214 (N_1214,N_694,In_325);
xor U1215 (N_1215,In_1929,N_626);
nor U1216 (N_1216,In_188,N_208);
and U1217 (N_1217,In_2093,In_1888);
or U1218 (N_1218,In_1163,N_987);
nor U1219 (N_1219,N_608,N_969);
xor U1220 (N_1220,In_980,N_531);
and U1221 (N_1221,In_299,In_1259);
nand U1222 (N_1222,In_309,In_1902);
and U1223 (N_1223,In_1144,In_2622);
and U1224 (N_1224,N_504,N_93);
and U1225 (N_1225,N_80,In_2913);
or U1226 (N_1226,In_748,N_897);
or U1227 (N_1227,N_60,N_702);
nand U1228 (N_1228,N_913,In_1966);
xor U1229 (N_1229,N_409,In_2091);
nand U1230 (N_1230,In_2492,N_109);
or U1231 (N_1231,N_879,N_135);
nor U1232 (N_1232,N_487,In_1898);
nor U1233 (N_1233,In_314,N_827);
nor U1234 (N_1234,In_2657,N_853);
xor U1235 (N_1235,In_878,In_1540);
xnor U1236 (N_1236,In_2390,In_712);
xnor U1237 (N_1237,In_1056,In_2252);
and U1238 (N_1238,N_859,N_746);
and U1239 (N_1239,N_473,In_2805);
nor U1240 (N_1240,N_737,In_2594);
and U1241 (N_1241,N_866,N_508);
nand U1242 (N_1242,In_788,In_480);
and U1243 (N_1243,In_902,N_842);
xnor U1244 (N_1244,In_1493,N_924);
or U1245 (N_1245,N_353,In_432);
nor U1246 (N_1246,In_2207,In_1594);
xnor U1247 (N_1247,In_1287,N_569);
xor U1248 (N_1248,In_2353,In_1478);
or U1249 (N_1249,In_1836,N_19);
xnor U1250 (N_1250,In_2548,In_2982);
or U1251 (N_1251,N_659,In_408);
xnor U1252 (N_1252,N_557,In_844);
nand U1253 (N_1253,In_1665,In_1797);
or U1254 (N_1254,N_909,N_670);
and U1255 (N_1255,N_443,N_560);
nor U1256 (N_1256,In_1161,In_1246);
and U1257 (N_1257,In_150,In_1299);
or U1258 (N_1258,In_1039,In_935);
and U1259 (N_1259,N_607,In_974);
xor U1260 (N_1260,In_2077,N_901);
and U1261 (N_1261,N_174,In_1345);
xnor U1262 (N_1262,N_921,N_902);
nor U1263 (N_1263,N_298,In_214);
nand U1264 (N_1264,In_2280,N_774);
nor U1265 (N_1265,In_2656,N_874);
and U1266 (N_1266,N_634,N_816);
nor U1267 (N_1267,In_1589,In_2903);
and U1268 (N_1268,N_623,N_770);
nand U1269 (N_1269,N_686,In_592);
nor U1270 (N_1270,N_453,N_414);
nor U1271 (N_1271,In_753,In_1205);
xor U1272 (N_1272,In_431,In_2498);
and U1273 (N_1273,N_214,In_713);
xor U1274 (N_1274,In_91,N_985);
nand U1275 (N_1275,In_2793,In_1637);
and U1276 (N_1276,In_1645,N_692);
xnor U1277 (N_1277,N_173,In_1658);
xor U1278 (N_1278,In_855,In_1474);
nor U1279 (N_1279,N_395,N_638);
nor U1280 (N_1280,In_2846,N_349);
or U1281 (N_1281,In_870,In_2986);
xnor U1282 (N_1282,N_926,In_287);
and U1283 (N_1283,In_436,In_2282);
or U1284 (N_1284,N_96,In_1777);
or U1285 (N_1285,In_142,In_2758);
nor U1286 (N_1286,N_285,In_50);
or U1287 (N_1287,In_117,In_1892);
xnor U1288 (N_1288,In_817,In_1158);
nor U1289 (N_1289,N_763,N_809);
nor U1290 (N_1290,In_223,N_206);
and U1291 (N_1291,In_2789,N_601);
or U1292 (N_1292,In_2467,N_980);
nand U1293 (N_1293,In_2521,In_1122);
nor U1294 (N_1294,N_991,In_129);
and U1295 (N_1295,In_2026,In_1431);
and U1296 (N_1296,In_1867,N_611);
and U1297 (N_1297,In_2686,N_250);
xor U1298 (N_1298,N_104,N_823);
xor U1299 (N_1299,In_306,N_651);
and U1300 (N_1300,N_382,N_721);
nand U1301 (N_1301,N_654,In_1076);
and U1302 (N_1302,N_824,In_541);
nor U1303 (N_1303,N_532,N_570);
xor U1304 (N_1304,In_416,In_1407);
nor U1305 (N_1305,N_36,N_944);
and U1306 (N_1306,In_657,In_1646);
xor U1307 (N_1307,In_2468,In_2643);
and U1308 (N_1308,N_758,In_1606);
xnor U1309 (N_1309,N_476,In_2126);
nand U1310 (N_1310,N_188,In_660);
nand U1311 (N_1311,In_110,In_1571);
xor U1312 (N_1312,N_810,In_1414);
nand U1313 (N_1313,In_1079,In_1717);
and U1314 (N_1314,In_2613,N_331);
xnor U1315 (N_1315,In_1147,In_2890);
nand U1316 (N_1316,N_875,N_342);
nand U1317 (N_1317,N_239,N_201);
xor U1318 (N_1318,In_729,N_597);
and U1319 (N_1319,N_522,N_359);
xor U1320 (N_1320,In_700,In_1418);
xor U1321 (N_1321,N_442,In_538);
or U1322 (N_1322,N_811,In_9);
xnor U1323 (N_1323,In_2076,In_484);
nor U1324 (N_1324,N_593,In_1420);
or U1325 (N_1325,In_600,N_291);
nand U1326 (N_1326,In_2011,In_1901);
or U1327 (N_1327,N_249,N_499);
xor U1328 (N_1328,In_1395,In_790);
xnor U1329 (N_1329,In_2216,In_398);
xor U1330 (N_1330,N_513,In_1887);
nand U1331 (N_1331,N_101,In_2732);
or U1332 (N_1332,In_2742,N_880);
and U1333 (N_1333,N_583,N_545);
xor U1334 (N_1334,In_2180,N_895);
or U1335 (N_1335,In_371,N_441);
and U1336 (N_1336,In_2275,N_975);
nand U1337 (N_1337,In_2005,In_337);
or U1338 (N_1338,N_889,In_1919);
nand U1339 (N_1339,In_2432,N_94);
or U1340 (N_1340,In_461,N_643);
and U1341 (N_1341,N_986,N_205);
xor U1342 (N_1342,In_75,N_535);
and U1343 (N_1343,N_438,N_26);
nor U1344 (N_1344,In_1557,In_550);
nand U1345 (N_1345,In_2418,N_2);
nand U1346 (N_1346,In_1127,In_2694);
or U1347 (N_1347,N_676,In_1373);
nor U1348 (N_1348,N_619,In_473);
and U1349 (N_1349,In_1940,In_1604);
nand U1350 (N_1350,In_1762,In_451);
or U1351 (N_1351,In_750,N_937);
xor U1352 (N_1352,In_96,In_2137);
xnor U1353 (N_1353,In_2617,In_2118);
xnor U1354 (N_1354,In_494,In_574);
or U1355 (N_1355,In_849,N_367);
or U1356 (N_1356,N_802,N_642);
or U1357 (N_1357,In_1049,In_1148);
xor U1358 (N_1358,N_417,In_422);
nor U1359 (N_1359,N_171,N_667);
xor U1360 (N_1360,N_928,In_1747);
nor U1361 (N_1361,In_1950,In_426);
nor U1362 (N_1362,In_2039,In_507);
nand U1363 (N_1363,In_401,In_2724);
and U1364 (N_1364,N_995,In_2258);
nor U1365 (N_1365,In_46,N_674);
or U1366 (N_1366,N_949,In_2315);
nor U1367 (N_1367,N_286,N_129);
and U1368 (N_1368,In_354,In_1012);
nand U1369 (N_1369,In_518,In_1799);
or U1370 (N_1370,N_970,In_84);
nand U1371 (N_1371,In_918,In_33);
nand U1372 (N_1372,In_1311,N_516);
nor U1373 (N_1373,In_2809,N_31);
and U1374 (N_1374,In_2641,In_235);
and U1375 (N_1375,In_1070,In_2892);
or U1376 (N_1376,N_28,In_2907);
nor U1377 (N_1377,N_78,N_829);
and U1378 (N_1378,N_867,In_1558);
and U1379 (N_1379,In_886,In_1573);
and U1380 (N_1380,N_33,N_57);
and U1381 (N_1381,In_1553,N_428);
and U1382 (N_1382,In_1358,N_122);
nand U1383 (N_1383,N_796,N_248);
nand U1384 (N_1384,In_311,N_925);
and U1385 (N_1385,In_948,In_1471);
nand U1386 (N_1386,In_1229,N_324);
xnor U1387 (N_1387,In_895,In_1129);
and U1388 (N_1388,In_1915,In_811);
nand U1389 (N_1389,N_401,In_1017);
nand U1390 (N_1390,N_307,In_1219);
nand U1391 (N_1391,N_501,In_926);
nand U1392 (N_1392,In_295,In_1909);
xnor U1393 (N_1393,In_1236,In_2814);
xnor U1394 (N_1394,In_1351,In_993);
and U1395 (N_1395,In_2893,In_909);
and U1396 (N_1396,In_1314,In_1086);
or U1397 (N_1397,N_664,In_835);
xnor U1398 (N_1398,In_2852,N_750);
and U1399 (N_1399,In_2410,In_367);
or U1400 (N_1400,In_1053,N_389);
nor U1401 (N_1401,N_863,N_281);
and U1402 (N_1402,N_752,N_568);
or U1403 (N_1403,In_465,N_482);
xnor U1404 (N_1404,In_735,In_717);
and U1405 (N_1405,In_158,In_1615);
and U1406 (N_1406,In_2534,In_664);
xor U1407 (N_1407,N_550,N_615);
xnor U1408 (N_1408,N_494,In_2801);
nand U1409 (N_1409,N_747,In_321);
nor U1410 (N_1410,In_1509,In_189);
nand U1411 (N_1411,N_160,N_475);
xor U1412 (N_1412,In_97,N_699);
xor U1413 (N_1413,N_738,In_1789);
xnor U1414 (N_1414,N_539,N_994);
or U1415 (N_1415,N_323,In_2940);
xor U1416 (N_1416,In_1904,In_1274);
xnor U1417 (N_1417,In_1490,In_218);
or U1418 (N_1418,N_776,In_1180);
xor U1419 (N_1419,N_780,In_1850);
and U1420 (N_1420,N_600,N_961);
xor U1421 (N_1421,In_1009,In_1683);
xor U1422 (N_1422,In_530,In_1999);
and U1423 (N_1423,N_661,In_2700);
xnor U1424 (N_1424,In_961,N_139);
and U1425 (N_1425,In_942,In_2144);
nor U1426 (N_1426,In_2474,In_1422);
nor U1427 (N_1427,In_1399,In_614);
nor U1428 (N_1428,In_2197,In_665);
nand U1429 (N_1429,In_1933,In_893);
and U1430 (N_1430,N_740,In_869);
or U1431 (N_1431,N_149,N_585);
nand U1432 (N_1432,N_252,In_1978);
nand U1433 (N_1433,In_1501,In_1531);
or U1434 (N_1434,N_633,N_517);
and U1435 (N_1435,N_10,In_2316);
or U1436 (N_1436,In_2095,In_2147);
or U1437 (N_1437,In_1801,N_689);
nor U1438 (N_1438,N_213,In_1383);
nor U1439 (N_1439,N_423,In_2967);
xor U1440 (N_1440,In_409,In_683);
and U1441 (N_1441,N_119,In_1469);
xor U1442 (N_1442,In_1988,N_946);
nor U1443 (N_1443,N_549,In_2441);
nand U1444 (N_1444,N_301,In_2130);
and U1445 (N_1445,In_1359,In_2373);
xor U1446 (N_1446,N_284,In_2994);
nor U1447 (N_1447,In_1258,In_1638);
xor U1448 (N_1448,In_2704,In_2593);
or U1449 (N_1449,In_2376,In_2526);
nand U1450 (N_1450,N_574,In_2257);
nand U1451 (N_1451,In_1566,In_813);
nor U1452 (N_1452,In_915,N_591);
xor U1453 (N_1453,In_2056,N_972);
nor U1454 (N_1454,In_2356,In_758);
nor U1455 (N_1455,In_131,N_525);
nor U1456 (N_1456,In_2813,In_1106);
nor U1457 (N_1457,In_1917,In_1824);
nor U1458 (N_1458,In_705,N_705);
xnor U1459 (N_1459,In_1536,N_533);
nor U1460 (N_1460,In_1282,N_211);
nand U1461 (N_1461,In_1149,N_420);
nand U1462 (N_1462,In_1580,In_531);
xor U1463 (N_1463,N_30,N_318);
nand U1464 (N_1464,In_1032,In_1786);
nor U1465 (N_1465,N_596,In_618);
and U1466 (N_1466,In_11,N_854);
nand U1467 (N_1467,In_2333,In_2326);
or U1468 (N_1468,In_2650,In_2380);
or U1469 (N_1469,In_149,In_2998);
xnor U1470 (N_1470,In_201,N_717);
nor U1471 (N_1471,N_605,N_783);
xnor U1472 (N_1472,N_753,In_2206);
and U1473 (N_1473,In_2850,N_576);
nor U1474 (N_1474,N_785,In_658);
and U1475 (N_1475,In_1724,N_391);
nand U1476 (N_1476,In_2583,In_1652);
and U1477 (N_1477,N_375,In_2177);
and U1478 (N_1478,N_303,In_930);
nor U1479 (N_1479,In_1628,In_2276);
nor U1480 (N_1480,In_2375,In_1337);
nand U1481 (N_1481,N_27,In_613);
and U1482 (N_1482,N_77,In_74);
and U1483 (N_1483,N_960,N_162);
nand U1484 (N_1484,In_324,N_16);
and U1485 (N_1485,In_2358,In_1832);
or U1486 (N_1486,In_1998,N_939);
nand U1487 (N_1487,N_653,In_2673);
or U1488 (N_1488,N_210,In_1119);
nor U1489 (N_1489,N_806,In_2831);
nand U1490 (N_1490,N_480,In_1470);
nor U1491 (N_1491,In_475,In_982);
xnor U1492 (N_1492,In_2341,In_1178);
or U1493 (N_1493,N_862,In_814);
or U1494 (N_1494,N_894,N_760);
or U1495 (N_1495,In_1213,N_648);
xnor U1496 (N_1496,N_613,N_178);
xor U1497 (N_1497,In_393,N_716);
or U1498 (N_1498,In_1852,In_1625);
nor U1499 (N_1499,In_612,N_333);
nand U1500 (N_1500,N_929,N_652);
nand U1501 (N_1501,N_1203,N_172);
or U1502 (N_1502,N_588,N_524);
xor U1503 (N_1503,N_481,N_1340);
xor U1504 (N_1504,In_1827,N_512);
or U1505 (N_1505,N_1336,N_743);
xor U1506 (N_1506,N_974,In_2030);
nor U1507 (N_1507,N_1307,In_2488);
and U1508 (N_1508,N_1104,In_2446);
and U1509 (N_1509,N_1197,N_1069);
and U1510 (N_1510,N_97,N_744);
and U1511 (N_1511,In_1301,N_1244);
nand U1512 (N_1512,N_1414,N_1402);
xnor U1513 (N_1513,N_1446,N_1057);
nor U1514 (N_1514,In_365,N_541);
or U1515 (N_1515,N_685,In_2838);
nand U1516 (N_1516,N_851,In_526);
and U1517 (N_1517,N_53,N_1385);
nand U1518 (N_1518,N_1186,N_882);
nand U1519 (N_1519,In_2589,In_1268);
xnor U1520 (N_1520,In_2431,In_1111);
and U1521 (N_1521,In_148,N_1391);
or U1522 (N_1522,In_330,N_840);
xnor U1523 (N_1523,N_1062,In_2784);
or U1524 (N_1524,N_1048,N_784);
xor U1525 (N_1525,N_764,In_2001);
xnor U1526 (N_1526,N_1320,N_860);
xor U1527 (N_1527,N_1352,N_1079);
or U1528 (N_1528,In_2384,In_2988);
nand U1529 (N_1529,In_2861,N_1233);
nor U1530 (N_1530,N_883,N_1457);
or U1531 (N_1531,In_491,In_2270);
nand U1532 (N_1532,In_1980,N_1006);
nor U1533 (N_1533,N_1015,N_1158);
xor U1534 (N_1534,In_2948,N_1054);
or U1535 (N_1535,In_1081,N_1004);
nand U1536 (N_1536,In_2181,N_1433);
and U1537 (N_1537,In_2804,In_1389);
nand U1538 (N_1538,In_2501,N_977);
xor U1539 (N_1539,In_206,In_1393);
or U1540 (N_1540,N_564,In_1203);
nand U1541 (N_1541,In_2103,N_7);
nor U1542 (N_1542,N_1217,In_2604);
nand U1543 (N_1543,N_105,In_763);
or U1544 (N_1544,N_629,In_2097);
nand U1545 (N_1545,N_1293,In_1477);
and U1546 (N_1546,In_2674,In_2817);
nor U1547 (N_1547,In_2135,N_408);
nor U1548 (N_1548,In_602,N_1035);
or U1549 (N_1549,In_1811,N_771);
nor U1550 (N_1550,N_566,In_1649);
nand U1551 (N_1551,N_843,N_280);
xor U1552 (N_1552,In_1413,N_936);
nand U1553 (N_1553,In_178,In_2564);
or U1554 (N_1554,N_769,N_1332);
or U1555 (N_1555,In_1795,In_1907);
and U1556 (N_1556,N_255,In_2695);
xor U1557 (N_1557,N_1163,N_787);
xnor U1558 (N_1558,N_1132,In_1209);
and U1559 (N_1559,N_1437,In_2330);
and U1560 (N_1560,In_2926,N_1084);
xnor U1561 (N_1561,In_2644,In_1020);
nand U1562 (N_1562,N_581,N_754);
or U1563 (N_1563,N_267,In_1873);
or U1564 (N_1564,N_962,N_1359);
and U1565 (N_1565,In_421,N_1440);
and U1566 (N_1566,In_989,N_800);
xor U1567 (N_1567,In_1014,In_2507);
xnor U1568 (N_1568,In_1060,N_509);
and U1569 (N_1569,N_1283,N_133);
and U1570 (N_1570,N_736,N_1496);
nor U1571 (N_1571,In_1196,N_159);
xnor U1572 (N_1572,In_967,In_146);
and U1573 (N_1573,N_1129,In_1921);
xor U1574 (N_1574,N_1474,N_1326);
nand U1575 (N_1575,N_1370,N_114);
nor U1576 (N_1576,N_573,In_2363);
xnor U1577 (N_1577,In_1976,In_1764);
and U1578 (N_1578,In_1375,N_1232);
and U1579 (N_1579,N_1353,In_1331);
nor U1580 (N_1580,N_1063,In_2873);
or U1581 (N_1581,In_2173,In_1264);
nor U1582 (N_1582,N_1207,In_2828);
nor U1583 (N_1583,N_1341,N_1486);
nor U1584 (N_1584,N_625,N_1087);
xnor U1585 (N_1585,N_1322,In_2226);
nor U1586 (N_1586,In_2236,N_143);
or U1587 (N_1587,N_679,N_1361);
or U1588 (N_1588,N_1431,N_1014);
nand U1589 (N_1589,In_1733,N_1327);
and U1590 (N_1590,N_1255,In_2539);
and U1591 (N_1591,N_1031,In_154);
nor U1592 (N_1592,N_1149,N_616);
and U1593 (N_1593,In_582,N_1438);
or U1594 (N_1594,N_1463,N_1234);
or U1595 (N_1595,In_985,In_560);
nor U1596 (N_1596,N_1127,In_2713);
nand U1597 (N_1597,N_598,In_1438);
xnor U1598 (N_1598,N_79,N_1383);
nand U1599 (N_1599,N_429,N_1258);
xor U1600 (N_1600,N_614,N_567);
nor U1601 (N_1601,In_889,N_951);
and U1602 (N_1602,N_1102,In_1969);
nand U1603 (N_1603,N_14,In_903);
and U1604 (N_1604,In_128,N_1112);
or U1605 (N_1605,N_1076,N_1181);
nand U1606 (N_1606,In_2354,N_1144);
nor U1607 (N_1607,In_439,N_988);
nand U1608 (N_1608,N_1419,N_1267);
nand U1609 (N_1609,N_1298,In_2058);
and U1610 (N_1610,N_580,N_293);
or U1611 (N_1611,N_1130,N_1401);
xnor U1612 (N_1612,In_2263,N_1115);
or U1613 (N_1613,N_1490,N_1125);
nand U1614 (N_1614,N_1138,In_2016);
nand U1615 (N_1615,In_1071,N_772);
xnor U1616 (N_1616,In_285,N_1188);
nand U1617 (N_1617,In_1453,N_1107);
xnor U1618 (N_1618,In_2336,In_1931);
nor U1619 (N_1619,In_1618,N_1075);
nand U1620 (N_1620,N_845,N_1051);
or U1621 (N_1621,N_742,N_1036);
xor U1622 (N_1622,N_1049,N_1109);
or U1623 (N_1623,In_1991,N_1262);
nand U1624 (N_1624,N_1268,In_2222);
xor U1625 (N_1625,N_1093,In_1104);
or U1626 (N_1626,N_906,In_513);
nand U1627 (N_1627,N_1466,In_1349);
xnor U1628 (N_1628,N_1142,N_751);
xor U1629 (N_1629,N_24,N_1042);
or U1630 (N_1630,N_799,N_1065);
or U1631 (N_1631,N_1174,N_1055);
nor U1632 (N_1632,N_602,N_687);
nor U1633 (N_1633,In_765,N_885);
or U1634 (N_1634,N_1371,In_2992);
nand U1635 (N_1635,N_1047,N_1291);
nor U1636 (N_1636,In_888,In_1128);
nor U1637 (N_1637,N_1476,In_1457);
nor U1638 (N_1638,N_1228,N_344);
or U1639 (N_1639,N_1071,N_1400);
nand U1640 (N_1640,N_1318,In_2856);
and U1641 (N_1641,N_1434,In_1290);
and U1642 (N_1642,N_953,N_1261);
or U1643 (N_1643,N_1199,N_1397);
or U1644 (N_1644,N_1089,N_1281);
and U1645 (N_1645,N_22,N_123);
nand U1646 (N_1646,In_676,N_185);
nand U1647 (N_1647,In_1357,N_1090);
xnor U1648 (N_1648,N_1098,N_161);
and U1649 (N_1649,In_1130,N_50);
or U1650 (N_1650,In_1228,N_935);
nor U1651 (N_1651,In_192,In_949);
and U1652 (N_1652,N_1470,In_2779);
nand U1653 (N_1653,In_1785,N_433);
or U1654 (N_1654,In_1896,N_690);
xor U1655 (N_1655,In_2952,N_543);
xnor U1656 (N_1656,In_305,In_1754);
xnor U1657 (N_1657,In_781,N_1027);
nand U1658 (N_1658,In_2629,In_1871);
nor U1659 (N_1659,N_1083,N_603);
nand U1660 (N_1660,In_107,In_2425);
nor U1661 (N_1661,In_496,N_620);
or U1662 (N_1662,N_1243,In_1289);
and U1663 (N_1663,N_340,N_1034);
nand U1664 (N_1664,In_2797,In_1105);
xor U1665 (N_1665,In_824,N_268);
xnor U1666 (N_1666,N_1299,N_1404);
nor U1667 (N_1667,N_814,In_1737);
and U1668 (N_1668,N_112,In_1216);
nand U1669 (N_1669,N_1208,In_2603);
or U1670 (N_1670,In_1080,In_1093);
and U1671 (N_1671,N_1369,In_988);
xor U1672 (N_1672,N_1046,N_1000);
nor U1673 (N_1673,In_1179,N_1002);
nand U1674 (N_1674,N_264,N_1415);
xnor U1675 (N_1675,N_1282,N_1222);
nor U1676 (N_1676,N_1312,In_108);
or U1677 (N_1677,In_1975,In_772);
or U1678 (N_1678,In_2288,In_238);
and U1679 (N_1679,N_158,In_2146);
nor U1680 (N_1680,N_1377,In_1091);
nor U1681 (N_1681,N_1343,N_1113);
nor U1682 (N_1682,In_2990,N_1236);
and U1683 (N_1683,In_1011,N_1491);
xnor U1684 (N_1684,In_2402,N_68);
xnor U1685 (N_1685,N_1276,N_959);
nor U1686 (N_1686,In_2023,N_1339);
xor U1687 (N_1687,N_1161,In_553);
xor U1688 (N_1688,N_1350,In_2883);
or U1689 (N_1689,N_1141,In_2634);
xor U1690 (N_1690,In_2905,N_456);
xor U1691 (N_1691,N_244,N_519);
or U1692 (N_1692,In_693,N_956);
and U1693 (N_1693,N_852,N_766);
and U1694 (N_1694,In_2381,In_1496);
nor U1695 (N_1695,N_76,N_1373);
nor U1696 (N_1696,In_2832,In_1912);
xor U1697 (N_1697,N_390,In_2739);
nand U1698 (N_1698,In_57,N_1306);
nand U1699 (N_1699,N_1043,In_1159);
nor U1700 (N_1700,N_515,N_1499);
nand U1701 (N_1701,In_2958,N_807);
nor U1702 (N_1702,N_908,N_495);
xor U1703 (N_1703,In_2371,N_942);
nor U1704 (N_1704,N_1099,N_632);
nor U1705 (N_1705,In_1700,N_1347);
nor U1706 (N_1706,N_1478,In_1233);
nand U1707 (N_1707,N_1424,In_232);
nand U1708 (N_1708,N_931,N_203);
nand U1709 (N_1709,N_1365,N_1372);
and U1710 (N_1710,In_1113,N_1059);
and U1711 (N_1711,N_628,N_1477);
nor U1712 (N_1712,In_2606,N_226);
nor U1713 (N_1713,N_1338,N_1018);
and U1714 (N_1714,N_886,In_578);
xnor U1715 (N_1715,In_2193,N_815);
and U1716 (N_1716,N_1037,N_1259);
nor U1717 (N_1717,N_1252,N_730);
and U1718 (N_1718,N_1484,N_1164);
and U1719 (N_1719,In_2047,N_888);
and U1720 (N_1720,N_893,N_551);
and U1721 (N_1721,N_1003,N_242);
nor U1722 (N_1722,N_910,N_316);
or U1723 (N_1723,N_731,N_1133);
xor U1724 (N_1724,N_462,N_1272);
or U1725 (N_1725,In_1985,N_1356);
nand U1726 (N_1726,N_537,In_2179);
nor U1727 (N_1727,In_731,In_2586);
or U1728 (N_1728,N_1488,N_630);
nor U1729 (N_1729,N_1449,In_1023);
nor U1730 (N_1730,N_465,In_1953);
or U1731 (N_1731,In_448,N_881);
xnor U1732 (N_1732,In_118,N_813);
nor U1733 (N_1733,N_1456,In_1752);
xor U1734 (N_1734,N_1078,In_1972);
xor U1735 (N_1735,In_962,In_2176);
nor U1736 (N_1736,In_2949,N_979);
nor U1737 (N_1737,N_1230,N_1167);
or U1738 (N_1738,N_1331,N_1481);
or U1739 (N_1739,N_884,N_1165);
xnor U1740 (N_1740,N_1464,In_2985);
or U1741 (N_1741,In_707,In_1316);
or U1742 (N_1742,In_342,In_1879);
or U1743 (N_1743,N_1273,N_1333);
nor U1744 (N_1744,In_1692,N_641);
or U1745 (N_1745,N_1183,N_1498);
or U1746 (N_1746,N_335,In_1636);
nor U1747 (N_1747,In_2301,N_1194);
or U1748 (N_1748,N_1417,N_899);
nor U1749 (N_1749,N_671,In_18);
nor U1750 (N_1750,In_2253,N_1074);
xnor U1751 (N_1751,N_1452,N_1250);
and U1752 (N_1752,N_1200,N_1066);
or U1753 (N_1753,N_45,N_1060);
xor U1754 (N_1754,In_1947,In_2688);
nor U1755 (N_1755,N_1028,In_492);
nand U1756 (N_1756,N_1162,In_68);
and U1757 (N_1757,In_2516,In_927);
nand U1758 (N_1758,In_1284,In_2932);
nand U1759 (N_1759,N_1489,N_708);
or U1760 (N_1760,In_2329,In_1034);
nand U1761 (N_1761,N_184,N_69);
and U1762 (N_1762,N_822,N_198);
xor U1763 (N_1763,N_669,N_963);
nor U1764 (N_1764,N_790,N_713);
or U1765 (N_1765,In_2851,N_707);
or U1766 (N_1766,N_1119,In_2827);
or U1767 (N_1767,N_812,In_725);
or U1768 (N_1768,N_1393,In_347);
nor U1769 (N_1769,N_1411,N_1136);
or U1770 (N_1770,N_1346,N_658);
and U1771 (N_1771,N_553,N_982);
and U1772 (N_1772,In_234,N_672);
nor U1773 (N_1773,In_838,N_1439);
xnor U1774 (N_1774,In_1759,N_405);
and U1775 (N_1775,N_927,In_2537);
nor U1776 (N_1776,N_903,In_487);
nand U1777 (N_1777,N_1064,N_362);
and U1778 (N_1778,In_1798,In_1249);
or U1779 (N_1779,N_189,In_152);
nand U1780 (N_1780,N_1290,N_896);
xor U1781 (N_1781,N_1334,N_562);
nand U1782 (N_1782,N_1448,N_1460);
nor U1783 (N_1783,In_1110,In_740);
nand U1784 (N_1784,N_1175,N_644);
nor U1785 (N_1785,N_1313,N_1105);
and U1786 (N_1786,N_1295,In_2760);
nor U1787 (N_1787,N_759,N_1177);
nand U1788 (N_1788,N_622,In_586);
nand U1789 (N_1789,In_2800,In_637);
nor U1790 (N_1790,N_445,N_358);
nor U1791 (N_1791,In_1601,In_2737);
or U1792 (N_1792,In_505,N_1279);
xor U1793 (N_1793,N_1366,In_2924);
nand U1794 (N_1794,In_1097,N_873);
xnor U1795 (N_1795,N_1169,N_695);
nand U1796 (N_1796,N_1187,N_726);
nand U1797 (N_1797,N_0,N_471);
xor U1798 (N_1798,N_81,N_1381);
or U1799 (N_1799,N_1179,N_967);
nor U1800 (N_1800,In_563,N_1392);
nand U1801 (N_1801,N_838,In_2113);
nor U1802 (N_1802,N_1367,N_1170);
nor U1803 (N_1803,In_1404,N_1085);
xnor U1804 (N_1804,N_1245,In_1421);
nor U1805 (N_1805,N_725,In_1240);
and U1806 (N_1806,N_1248,N_1204);
nor U1807 (N_1807,N_1020,In_2221);
xnor U1808 (N_1808,N_1458,N_1189);
or U1809 (N_1809,N_1342,N_1455);
or U1810 (N_1810,In_1574,N_1495);
xor U1811 (N_1811,In_1563,N_1041);
xnor U1812 (N_1812,N_1153,N_1443);
xor U1813 (N_1813,N_287,In_932);
xnor U1814 (N_1814,In_1659,N_849);
or U1815 (N_1815,In_2495,N_1023);
or U1816 (N_1816,In_503,In_1579);
nand U1817 (N_1817,N_1052,N_1277);
or U1818 (N_1818,In_536,N_1390);
and U1819 (N_1819,In_1145,N_51);
nor U1820 (N_1820,N_681,N_256);
or U1821 (N_1821,N_868,In_2080);
xor U1822 (N_1822,N_1321,In_38);
nor U1823 (N_1823,N_1045,N_1469);
nor U1824 (N_1824,N_1374,In_1286);
nor U1825 (N_1825,N_329,N_943);
nand U1826 (N_1826,In_1551,N_678);
nor U1827 (N_1827,N_1468,N_647);
xnor U1828 (N_1828,In_1101,N_1030);
nor U1829 (N_1829,N_1150,N_177);
and U1830 (N_1830,In_1716,N_631);
and U1831 (N_1831,N_1427,N_1191);
and U1832 (N_1832,N_914,N_830);
nand U1833 (N_1833,In_458,N_1447);
and U1834 (N_1834,N_1219,In_2247);
xnor U1835 (N_1835,N_1429,N_1011);
and U1836 (N_1836,N_1025,In_2712);
nor U1837 (N_1837,In_1406,In_1283);
and U1838 (N_1838,N_898,In_876);
or U1839 (N_1839,N_1103,N_976);
and U1840 (N_1840,N_265,N_38);
or U1841 (N_1841,N_1348,In_2387);
nand U1842 (N_1842,In_999,N_314);
nor U1843 (N_1843,In_2914,N_955);
nor U1844 (N_1844,In_590,In_1296);
and U1845 (N_1845,In_2741,N_1121);
xor U1846 (N_1846,In_871,In_1542);
nor U1847 (N_1847,N_1305,N_624);
or U1848 (N_1848,In_2386,N_1344);
nor U1849 (N_1849,N_724,In_1963);
or U1850 (N_1850,N_450,In_1168);
or U1851 (N_1851,In_1788,N_680);
nand U1852 (N_1852,N_734,N_1155);
nor U1853 (N_1853,In_1889,In_2502);
nor U1854 (N_1854,N_1413,N_698);
nand U1855 (N_1855,N_1317,N_386);
nand U1856 (N_1856,N_1024,In_2675);
nor U1857 (N_1857,In_2066,N_1206);
xor U1858 (N_1858,N_997,N_332);
nand U1859 (N_1859,N_1311,N_1435);
and U1860 (N_1860,N_584,In_2414);
nor U1861 (N_1861,N_1038,N_1441);
and U1862 (N_1862,In_2217,N_548);
nor U1863 (N_1863,N_305,N_745);
and U1864 (N_1864,In_867,In_1271);
nor U1865 (N_1865,In_251,N_1122);
nand U1866 (N_1866,In_506,N_166);
or U1867 (N_1867,N_1309,In_1587);
and U1868 (N_1868,N_1190,In_2964);
nor U1869 (N_1869,N_604,N_304);
nand U1870 (N_1870,In_872,N_108);
and U1871 (N_1871,N_1152,In_1102);
xor U1872 (N_1872,N_1224,In_2672);
or U1873 (N_1873,In_821,N_684);
xor U1874 (N_1874,N_663,N_1396);
nand U1875 (N_1875,N_507,N_1405);
and U1876 (N_1876,N_645,In_1066);
nand U1877 (N_1877,N_1101,N_193);
nor U1878 (N_1878,In_1325,In_79);
or U1879 (N_1879,N_788,N_748);
or U1880 (N_1880,N_682,In_1545);
and U1881 (N_1881,In_2408,In_2762);
nand U1882 (N_1882,N_1260,In_540);
nor U1883 (N_1883,N_283,In_2169);
xor U1884 (N_1884,In_2600,In_954);
nor U1885 (N_1885,N_1275,N_514);
nor U1886 (N_1886,N_317,N_578);
or U1887 (N_1887,In_489,N_1479);
xor U1888 (N_1888,In_566,N_35);
nor U1889 (N_1889,N_1185,In_1497);
xnor U1890 (N_1890,In_2119,N_1368);
or U1891 (N_1891,N_415,N_948);
nand U1892 (N_1892,N_1056,N_590);
nor U1893 (N_1893,N_1454,N_919);
and U1894 (N_1894,N_1242,In_796);
nand U1895 (N_1895,In_1770,In_1171);
nand U1896 (N_1896,N_1238,N_1382);
or U1897 (N_1897,In_185,N_1287);
xnor U1898 (N_1898,N_422,In_1095);
nand U1899 (N_1899,N_1247,In_706);
and U1900 (N_1900,N_1471,N_741);
or U1901 (N_1901,N_339,In_1321);
or U1902 (N_1902,N_1212,N_655);
nor U1903 (N_1903,N_196,In_2956);
xor U1904 (N_1904,N_938,N_1091);
and U1905 (N_1905,N_485,N_1358);
xor U1906 (N_1906,N_1398,In_2310);
or U1907 (N_1907,In_1059,N_1140);
xor U1908 (N_1908,N_586,In_1330);
xor U1909 (N_1909,In_1443,N_352);
nor U1910 (N_1910,In_1667,N_1461);
nor U1911 (N_1911,In_1761,N_1289);
nor U1912 (N_1912,In_2714,N_627);
xnor U1913 (N_1913,N_503,N_930);
nand U1914 (N_1914,In_547,In_2551);
or U1915 (N_1915,In_996,N_803);
and U1916 (N_1916,N_1092,In_2648);
nor U1917 (N_1917,N_1135,N_547);
and U1918 (N_1918,In_318,N_640);
nor U1919 (N_1919,N_370,In_2073);
nand U1920 (N_1920,In_1866,In_2499);
nor U1921 (N_1921,N_223,N_397);
nand U1922 (N_1922,N_558,In_1995);
nand U1923 (N_1923,In_2048,N_1120);
xor U1924 (N_1924,N_552,N_1029);
nand U1925 (N_1925,N_923,N_1081);
xnor U1926 (N_1926,N_540,In_917);
nand U1927 (N_1927,N_1406,In_2727);
nor U1928 (N_1928,N_1172,In_392);
nand U1929 (N_1929,In_2090,N_1073);
and U1930 (N_1930,In_807,N_1349);
nor U1931 (N_1931,In_2847,In_495);
xnor U1932 (N_1932,N_258,N_561);
and U1933 (N_1933,In_303,In_1005);
nand U1934 (N_1934,In_1044,N_1256);
and U1935 (N_1935,N_981,N_782);
nand U1936 (N_1936,N_1146,N_1375);
nor U1937 (N_1937,N_1384,In_2453);
or U1938 (N_1938,In_2582,N_1017);
or U1939 (N_1939,In_171,N_922);
xnor U1940 (N_1940,N_1410,N_1249);
xnor U1941 (N_1941,N_835,N_900);
nand U1942 (N_1942,N_918,N_1159);
nand U1943 (N_1943,In_2759,N_834);
nand U1944 (N_1944,In_2960,N_592);
nand U1945 (N_1945,N_1218,In_1903);
nor U1946 (N_1946,N_646,N_728);
xnor U1947 (N_1947,N_718,In_2708);
xnor U1948 (N_1948,In_1702,N_1462);
nor U1949 (N_1949,N_1335,N_1148);
and U1950 (N_1950,N_385,In_99);
nor U1951 (N_1951,N_1195,N_270);
nor U1952 (N_1952,In_1454,N_1001);
nand U1953 (N_1953,N_954,In_2975);
and U1954 (N_1954,N_1088,N_368);
nor U1955 (N_1955,N_887,N_1323);
nand U1956 (N_1956,In_1067,N_870);
xor U1957 (N_1957,In_1380,In_1859);
xnor U1958 (N_1958,In_180,N_795);
or U1959 (N_1959,In_1369,N_957);
or U1960 (N_1960,N_1117,N_144);
nor U1961 (N_1961,In_1000,In_456);
xor U1962 (N_1962,N_1016,N_587);
or U1963 (N_1963,N_534,N_1214);
nand U1964 (N_1964,N_1176,In_236);
and U1965 (N_1965,N_1193,In_1547);
and U1966 (N_1966,N_932,In_2212);
or U1967 (N_1967,N_1239,In_2357);
xnor U1968 (N_1968,N_124,In_49);
and U1969 (N_1969,N_1157,In_2374);
nor U1970 (N_1970,In_714,N_1053);
and U1971 (N_1971,N_905,N_1451);
nor U1972 (N_1972,N_1171,In_1576);
nand U1973 (N_1973,N_186,In_852);
nor U1974 (N_1974,In_1778,In_2152);
xor U1975 (N_1975,In_1986,N_1237);
nand U1976 (N_1976,In_77,N_1240);
or U1977 (N_1977,N_1426,In_1370);
or U1978 (N_1978,N_1241,In_924);
and U1979 (N_1979,N_618,In_2157);
or U1980 (N_1980,N_498,In_319);
nor U1981 (N_1981,N_529,N_786);
xnor U1982 (N_1982,N_1096,N_1097);
nor U1983 (N_1983,N_1210,In_81);
xnor U1984 (N_1984,In_359,N_855);
nand U1985 (N_1985,N_132,N_330);
nand U1986 (N_1986,In_1958,N_1297);
nor U1987 (N_1987,In_2580,In_1480);
nor U1988 (N_1988,In_362,In_2504);
xor U1989 (N_1989,N_154,In_839);
and U1990 (N_1990,In_5,N_1111);
and U1991 (N_1991,N_338,In_481);
or U1992 (N_1992,In_2200,N_181);
and U1993 (N_1993,N_222,In_2059);
or U1994 (N_1994,N_1012,In_608);
xor U1995 (N_1995,In_2415,N_1108);
and U1996 (N_1996,In_1440,In_4);
xor U1997 (N_1997,N_4,In_2881);
nand U1998 (N_1998,N_1403,In_2803);
xnor U1999 (N_1999,N_818,N_1286);
nor U2000 (N_2000,In_751,N_1655);
and U2001 (N_2001,N_1690,N_1418);
nand U2002 (N_2002,N_1386,N_1032);
nor U2003 (N_2003,In_605,N_1779);
and U2004 (N_2004,N_1007,N_637);
xor U2005 (N_2005,N_1430,N_1839);
xor U2006 (N_2006,In_1136,N_1607);
nand U2007 (N_2007,In_1112,N_1205);
or U2008 (N_2008,In_1269,N_243);
or U2009 (N_2009,N_1972,N_1733);
xor U2010 (N_2010,N_1754,N_749);
nand U2011 (N_2011,N_1717,N_1493);
nor U2012 (N_2012,N_1630,N_1658);
nor U2013 (N_2013,N_1954,N_1269);
and U2014 (N_2014,N_572,In_699);
nand U2015 (N_2015,In_21,In_51);
nor U2016 (N_2016,N_1982,N_1100);
and U2017 (N_2017,In_511,N_1855);
or U2018 (N_2018,In_2428,N_1882);
nand U2019 (N_2019,In_425,N_1944);
nand U2020 (N_2020,N_1787,N_1571);
xnor U2021 (N_2021,In_972,N_1894);
and U2022 (N_2022,In_795,N_1723);
or U2023 (N_2023,N_1849,In_2046);
nand U2024 (N_2024,N_1663,N_1612);
nand U2025 (N_2025,N_1363,N_1966);
nand U2026 (N_2026,N_1211,N_1670);
nand U2027 (N_2027,N_1831,N_106);
and U2028 (N_2028,N_1220,N_1131);
nor U2029 (N_2029,N_1969,N_1801);
xor U2030 (N_2030,N_933,N_1525);
nor U2031 (N_2031,N_1985,In_603);
nor U2032 (N_2032,N_1620,N_1453);
nor U2033 (N_2033,In_1954,N_1933);
nand U2034 (N_2034,N_1784,N_1409);
and U2035 (N_2035,N_1616,N_1772);
nand U2036 (N_2036,N_1548,N_1702);
or U2037 (N_2037,N_1379,N_1927);
or U2038 (N_2038,N_1715,N_1851);
nand U2039 (N_2039,N_1749,N_1202);
nor U2040 (N_2040,N_1879,In_812);
xnor U2041 (N_2041,N_1337,In_1926);
or U2042 (N_2042,In_1983,N_1705);
or U2043 (N_2043,In_2815,N_1492);
nor U2044 (N_2044,N_1033,N_636);
nor U2045 (N_2045,N_460,N_1292);
xnor U2046 (N_2046,N_1910,In_1227);
nand U2047 (N_2047,N_1639,N_1818);
nor U2048 (N_2048,In_2601,In_2979);
nor U2049 (N_2049,In_2684,N_1529);
xnor U2050 (N_2050,In_532,N_1380);
xor U2051 (N_2051,N_864,In_2751);
nor U2052 (N_2052,N_1505,N_1533);
nor U2053 (N_2053,N_1826,In_703);
and U2054 (N_2054,N_1815,In_322);
and U2055 (N_2055,In_1107,N_1916);
nor U2056 (N_2056,N_1977,N_706);
nor U2057 (N_2057,N_1538,N_1951);
and U2058 (N_2058,In_2897,N_1513);
xnor U2059 (N_2059,N_1914,N_1251);
xnor U2060 (N_2060,N_831,In_2670);
xor U2061 (N_2061,N_1834,N_1619);
or U2062 (N_2062,N_1946,N_1934);
nor U2063 (N_2063,N_464,N_1050);
xnor U2064 (N_2064,In_922,In_925);
and U2065 (N_2065,N_1960,In_1398);
nor U2066 (N_2066,N_1802,N_1436);
nand U2067 (N_2067,N_83,N_1930);
nand U2068 (N_2068,N_1147,N_857);
or U2069 (N_2069,N_398,N_1294);
nand U2070 (N_2070,In_2676,N_1825);
or U2071 (N_2071,N_1911,N_232);
nor U2072 (N_2072,N_1939,N_1932);
or U2073 (N_2073,N_1701,N_1794);
and U2074 (N_2074,N_1757,In_1177);
nand U2075 (N_2075,N_1626,N_1537);
xnor U2076 (N_2076,N_1806,N_542);
or U2077 (N_2077,N_1123,N_1816);
nand U2078 (N_2078,N_1893,N_1770);
or U2079 (N_2079,N_1667,In_1857);
nor U2080 (N_2080,N_1067,N_1432);
or U2081 (N_2081,N_1734,In_1016);
or U2082 (N_2082,N_1072,N_1653);
nor U2083 (N_2083,N_1895,N_1576);
and U2084 (N_2084,N_1617,N_1459);
nand U2085 (N_2085,N_1948,N_1859);
nor U2086 (N_2086,N_1585,N_1615);
xor U2087 (N_2087,In_2917,N_1395);
and U2088 (N_2088,N_1955,N_1080);
xor U2089 (N_2089,N_1679,N_773);
or U2090 (N_2090,N_1225,N_1989);
nand U2091 (N_2091,N_1673,N_1565);
nand U2092 (N_2092,N_459,N_1590);
or U2093 (N_2093,N_449,N_892);
nand U2094 (N_2094,In_2519,N_992);
nand U2095 (N_2095,N_1082,In_1519);
nand U2096 (N_2096,N_1166,N_1578);
nand U2097 (N_2097,N_1664,In_947);
xor U2098 (N_2098,N_1022,N_1721);
nor U2099 (N_2099,N_1886,N_1755);
xnor U2100 (N_2100,N_1345,N_1675);
or U2101 (N_2101,N_1502,In_767);
nand U2102 (N_2102,N_1741,In_2728);
nand U2103 (N_2103,N_1857,N_1995);
and U2104 (N_2104,N_1531,N_1887);
nand U2105 (N_2105,In_567,In_1841);
xnor U2106 (N_2106,N_1254,N_1534);
or U2107 (N_2107,N_1569,In_2239);
nor U2108 (N_2108,N_1304,N_1512);
nand U2109 (N_2109,N_1913,N_1523);
xnor U2110 (N_2110,N_1591,N_1582);
or U2111 (N_2111,N_1388,N_1316);
and U2112 (N_2112,N_269,N_1645);
nor U2113 (N_2113,N_1556,In_26);
nand U2114 (N_2114,N_1983,N_1751);
or U2115 (N_2115,N_1450,In_164);
and U2116 (N_2116,In_2264,N_1919);
nor U2117 (N_2117,N_1678,N_1901);
nor U2118 (N_2118,N_1725,In_1704);
and U2119 (N_2119,In_1024,N_1209);
xnor U2120 (N_2120,N_1627,N_1536);
or U2121 (N_2121,In_955,N_1040);
or U2122 (N_2122,N_1891,N_1737);
and U2123 (N_2123,N_1931,In_1920);
xnor U2124 (N_2124,N_1600,N_1213);
and U2125 (N_2125,N_1889,In_1214);
nand U2126 (N_2126,N_999,N_1997);
nor U2127 (N_2127,N_1423,N_1661);
nor U2128 (N_2128,N_1549,N_1868);
or U2129 (N_2129,N_1603,N_1708);
nor U2130 (N_2130,In_2249,N_1876);
xnor U2131 (N_2131,In_1900,N_1828);
nor U2132 (N_2132,N_1707,N_469);
and U2133 (N_2133,N_1724,N_1465);
xnor U2134 (N_2134,N_1561,N_1573);
nand U2135 (N_2135,In_1883,N_1771);
nand U2136 (N_2136,N_1445,In_591);
and U2137 (N_2137,N_1551,N_1687);
nand U2138 (N_2138,N_1399,In_1270);
and U2139 (N_2139,In_2974,N_1557);
xor U2140 (N_2140,In_2578,N_1274);
nand U2141 (N_2141,N_520,N_1722);
nand U2142 (N_2142,N_1915,In_1742);
nand U2143 (N_2143,In_1230,N_1510);
nand U2144 (N_2144,N_373,N_1683);
xnor U2145 (N_2145,N_915,N_1785);
nand U2146 (N_2146,N_1278,N_1235);
nor U2147 (N_2147,N_998,In_2040);
or U2148 (N_2148,N_1881,N_1738);
and U2149 (N_2149,N_1360,N_1727);
and U2150 (N_2150,N_1480,N_1812);
nand U2151 (N_2151,N_472,N_1923);
and U2152 (N_2152,N_1813,N_1145);
xor U2153 (N_2153,N_1599,In_2433);
or U2154 (N_2154,In_1250,In_1291);
or U2155 (N_2155,N_1714,N_1928);
xor U2156 (N_2156,In_1769,N_1792);
xor U2157 (N_2157,In_2839,N_1648);
nor U2158 (N_2158,N_1953,N_609);
xnor U2159 (N_2159,N_1957,In_1503);
nor U2160 (N_2160,In_1342,N_1508);
or U2161 (N_2161,N_1408,N_1970);
or U2162 (N_2162,N_1711,In_2523);
xor U2163 (N_2163,In_2311,N_1005);
nor U2164 (N_2164,N_1647,In_802);
and U2165 (N_2165,N_1795,N_1503);
nor U2166 (N_2166,N_1128,N_1602);
nand U2167 (N_2167,In_1218,In_2017);
nand U2168 (N_2168,N_1842,In_2853);
nor U2169 (N_2169,In_1937,In_1760);
xnor U2170 (N_2170,In_478,N_1657);
nor U2171 (N_2171,N_1070,N_1581);
xnor U2172 (N_2172,N_1967,N_1998);
or U2173 (N_2173,N_1958,In_1960);
nor U2174 (N_2174,N_1671,N_1753);
or U2175 (N_2175,N_1285,N_1810);
xnor U2176 (N_2176,N_1594,N_1897);
nor U2177 (N_2177,N_1938,N_1629);
nand U2178 (N_2178,N_1584,N_1762);
and U2179 (N_2179,N_1837,In_931);
nand U2180 (N_2180,N_697,N_1692);
nand U2181 (N_2181,N_727,N_1610);
and U2182 (N_2182,N_1324,N_565);
nor U2183 (N_2183,N_1357,N_1284);
or U2184 (N_2184,In_161,N_1971);
nand U2185 (N_2185,N_40,N_1964);
nor U2186 (N_2186,N_1888,N_474);
xnor U2187 (N_2187,N_1819,N_1257);
nor U2188 (N_2188,N_1325,N_1118);
xnor U2189 (N_2189,N_1703,N_1900);
xnor U2190 (N_2190,In_1189,N_1829);
or U2191 (N_2191,N_1917,N_1173);
xor U2192 (N_2192,N_1959,N_732);
or U2193 (N_2193,N_1906,N_1226);
nor U2194 (N_2194,In_1807,N_1929);
nand U2195 (N_2195,N_1867,In_1541);
and U2196 (N_2196,N_1735,N_1740);
nand U2197 (N_2197,In_98,N_1376);
xor U2198 (N_2198,N_1180,In_865);
nor U2199 (N_2199,N_1871,N_1963);
and U2200 (N_2200,N_861,In_2585);
xnor U2201 (N_2201,N_1682,N_1800);
nor U2202 (N_2202,N_1821,N_461);
or U2203 (N_2203,In_89,N_1746);
nand U2204 (N_2204,N_1807,N_1649);
xnor U2205 (N_2205,In_1809,N_714);
xor U2206 (N_2206,N_1907,N_1700);
and U2207 (N_2207,N_1598,N_1674);
xnor U2208 (N_2208,In_1524,N_1416);
or U2209 (N_2209,N_1862,N_1330);
and U2210 (N_2210,N_1314,N_1988);
xor U2211 (N_2211,N_75,N_1778);
and U2212 (N_2212,In_294,N_1691);
nor U2213 (N_2213,In_1458,N_147);
nor U2214 (N_2214,N_1765,N_1562);
and U2215 (N_2215,N_1184,N_1838);
and U2216 (N_2216,N_762,N_1803);
or U2217 (N_2217,N_528,N_1822);
nand U2218 (N_2218,In_1552,N_1712);
nor U2219 (N_2219,N_1196,N_292);
and U2220 (N_2220,N_1774,N_1856);
and U2221 (N_2221,N_467,N_1912);
xnor U2222 (N_2222,In_575,In_2777);
xnor U2223 (N_2223,N_1543,N_1542);
or U2224 (N_2224,N_1216,N_1710);
xor U2225 (N_2225,N_1019,N_1168);
nand U2226 (N_2226,In_1927,N_668);
or U2227 (N_2227,N_220,N_1756);
or U2228 (N_2228,N_1182,In_279);
xor U2229 (N_2229,N_1793,N_1558);
or U2230 (N_2230,N_1010,N_1640);
nand U2231 (N_2231,N_1947,N_1902);
or U2232 (N_2232,N_1884,N_1497);
xor U2233 (N_2233,N_1805,N_1631);
nor U2234 (N_2234,In_52,N_793);
and U2235 (N_2235,N_1310,N_1328);
nand U2236 (N_2236,N_1634,N_1789);
or U2237 (N_2237,N_1973,N_1730);
and U2238 (N_2238,N_1126,N_1726);
or U2239 (N_2239,In_1208,N_1545);
nor U2240 (N_2240,N_1606,N_720);
xor U2241 (N_2241,N_1880,N_64);
or U2242 (N_2242,N_712,In_1498);
or U2243 (N_2243,N_1614,N_1935);
xor U2244 (N_2244,N_1528,N_546);
nand U2245 (N_2245,N_1768,N_610);
or U2246 (N_2246,N_1848,N_989);
nor U2247 (N_2247,N_37,N_297);
nand U2248 (N_2248,N_121,N_1719);
or U2249 (N_2249,N_56,N_1521);
or U2250 (N_2250,In_165,N_1875);
nor U2251 (N_2251,N_1364,N_1783);
nand U2252 (N_2252,N_1979,N_1597);
and U2253 (N_2253,N_1039,N_657);
xnor U2254 (N_2254,In_2863,N_1987);
nor U2255 (N_2255,N_1685,N_1716);
nor U2256 (N_2256,N_1552,N_1500);
nand U2257 (N_2257,N_850,N_1798);
nor U2258 (N_2258,N_1999,N_1699);
nand U2259 (N_2259,N_1583,N_1709);
and U2260 (N_2260,In_1965,In_880);
nor U2261 (N_2261,N_1519,N_1026);
and U2262 (N_2262,N_1588,N_1319);
nand U2263 (N_2263,N_1920,N_1693);
nor U2264 (N_2264,N_1593,In_2229);
and U2265 (N_2265,N_1547,N_1178);
xor U2266 (N_2266,N_1656,In_105);
nand U2267 (N_2267,N_1009,N_848);
and U2268 (N_2268,N_1713,N_1767);
xnor U2269 (N_2269,N_1743,In_2715);
and U2270 (N_2270,N_1574,N_1866);
or U2271 (N_2271,N_1835,N_1706);
xor U2272 (N_2272,N_1758,N_1790);
or U2273 (N_2273,N_719,N_993);
and U2274 (N_2274,N_1854,N_1263);
and U2275 (N_2275,N_934,N_1869);
xnor U2276 (N_2276,N_1936,N_1846);
nor U2277 (N_2277,N_1922,N_715);
and U2278 (N_2278,N_1520,N_1942);
nand U2279 (N_2279,N_1151,N_1086);
nand U2280 (N_2280,In_1021,N_1442);
nand U2281 (N_2281,N_1467,N_1472);
xnor U2282 (N_2282,N_1681,In_2454);
nor U2283 (N_2283,N_1483,N_492);
nor U2284 (N_2284,In_216,N_1227);
nand U2285 (N_2285,N_1444,N_1650);
and U2286 (N_2286,N_1501,N_1684);
and U2287 (N_2287,N_1861,N_1665);
nand U2288 (N_2288,N_1301,In_2753);
and U2289 (N_2289,N_1921,In_1666);
nor U2290 (N_2290,N_599,N_1137);
nor U2291 (N_2291,N_1781,N_1506);
nand U2292 (N_2292,N_1378,N_1986);
nand U2293 (N_2293,N_544,N_1058);
and U2294 (N_2294,In_606,N_1270);
nor U2295 (N_2295,N_1223,N_8);
nor U2296 (N_2296,N_1586,N_1300);
and U2297 (N_2297,N_1651,N_1515);
xor U2298 (N_2298,N_1694,N_1745);
nor U2299 (N_2299,N_1992,N_1596);
nor U2300 (N_2300,N_1752,N_733);
or U2301 (N_2301,N_1154,N_1874);
nor U2302 (N_2302,N_1546,N_209);
or U2303 (N_2303,In_1243,N_1124);
or U2304 (N_2304,In_666,N_1739);
nand U2305 (N_2305,N_1539,N_1788);
nand U2306 (N_2306,N_1580,N_1903);
or U2307 (N_2307,In_2128,N_1773);
nand U2308 (N_2308,N_191,N_1303);
or U2309 (N_2309,N_1736,N_666);
and U2310 (N_2310,N_1698,In_2308);
and U2311 (N_2311,N_447,N_1980);
and U2312 (N_2312,N_1680,N_1566);
nor U2313 (N_2313,In_2150,In_2227);
nand U2314 (N_2314,N_1761,N_1622);
and U2315 (N_2315,N_1271,In_2201);
or U2316 (N_2316,In_1964,N_1635);
and U2317 (N_2317,N_399,N_1797);
nor U2318 (N_2318,In_598,In_2443);
nor U2319 (N_2319,N_917,N_1808);
nor U2320 (N_2320,N_1864,N_1485);
and U2321 (N_2321,N_1564,N_282);
xnor U2322 (N_2322,N_907,N_828);
nand U2323 (N_2323,N_1747,In_1335);
xor U2324 (N_2324,N_673,N_1844);
or U2325 (N_2325,N_1116,N_489);
nand U2326 (N_2326,N_1198,N_1421);
nand U2327 (N_2327,N_1672,In_205);
nand U2328 (N_2328,N_1511,N_984);
and U2329 (N_2329,N_1021,N_1504);
nand U2330 (N_2330,N_1494,N_9);
or U2331 (N_2331,In_277,N_1530);
nor U2332 (N_2332,N_656,In_2278);
nor U2333 (N_2333,N_1796,N_1666);
nor U2334 (N_2334,N_1229,N_1908);
xnor U2335 (N_2335,In_568,In_565);
xnor U2336 (N_2336,N_1791,N_1139);
nand U2337 (N_2337,N_1994,In_450);
nor U2338 (N_2338,N_1830,N_1660);
and U2339 (N_2339,N_1845,N_1362);
xor U2340 (N_2340,N_91,In_2277);
or U2341 (N_2341,N_660,In_2469);
nand U2342 (N_2342,N_1759,N_110);
nor U2343 (N_2343,N_1008,N_1308);
or U2344 (N_2344,N_1925,N_1628);
nand U2345 (N_2345,In_2574,In_1441);
and U2346 (N_2346,N_1618,N_877);
nor U2347 (N_2347,N_1646,N_1720);
and U2348 (N_2348,N_1873,N_1697);
xor U2349 (N_2349,In_1994,In_2818);
and U2350 (N_2350,N_1993,N_1686);
or U2351 (N_2351,N_1990,N_233);
or U2352 (N_2352,In_2323,N_767);
and U2353 (N_2353,N_1221,In_483);
or U2354 (N_2354,In_265,N_1896);
nand U2355 (N_2355,N_1264,N_1652);
and U2356 (N_2356,N_1991,N_639);
nor U2357 (N_2357,In_1730,In_2299);
xor U2358 (N_2358,N_1892,N_479);
or U2359 (N_2359,N_1728,N_523);
nor U2360 (N_2360,In_2802,N_696);
nor U2361 (N_2361,N_950,N_141);
and U2362 (N_2362,N_1625,N_1296);
or U2363 (N_2363,N_1804,N_1689);
or U2364 (N_2364,N_1847,N_1563);
nand U2365 (N_2365,N_1560,N_1094);
and U2366 (N_2366,In_914,N_1507);
xnor U2367 (N_2367,N_1924,N_804);
nor U2368 (N_2368,In_2632,N_1114);
xor U2369 (N_2369,In_747,N_1143);
nand U2370 (N_2370,N_1817,N_675);
and U2371 (N_2371,N_844,N_1676);
or U2372 (N_2372,N_1823,N_1577);
xnor U2373 (N_2373,N_836,N_582);
xor U2374 (N_2374,In_2127,N_1518);
xor U2375 (N_2375,N_1532,In_162);
nand U2376 (N_2376,N_1763,N_1962);
nor U2377 (N_2377,N_1509,N_1412);
and U2378 (N_2378,N_1068,N_1592);
or U2379 (N_2379,N_1013,In_877);
nand U2380 (N_2380,In_845,N_29);
nand U2381 (N_2381,N_1280,N_1981);
nand U2382 (N_2382,In_283,N_1905);
nand U2383 (N_2383,N_1613,In_1599);
nand U2384 (N_2384,N_1748,N_1742);
xor U2385 (N_2385,N_1201,N_1731);
nor U2386 (N_2386,N_1595,N_1061);
xnor U2387 (N_2387,In_2693,N_1918);
nor U2388 (N_2388,N_1949,N_1633);
or U2389 (N_2389,N_1636,N_1688);
nor U2390 (N_2390,N_1836,N_235);
and U2391 (N_2391,N_1950,In_1688);
nor U2392 (N_2392,N_1799,N_1780);
nor U2393 (N_2393,N_1550,In_2256);
xnor U2394 (N_2394,N_1786,In_2202);
or U2395 (N_2395,N_1246,N_1482);
nor U2396 (N_2396,In_1560,N_1898);
or U2397 (N_2397,In_1622,N_1637);
and U2398 (N_2398,N_1394,N_1865);
or U2399 (N_2399,N_1570,N_1654);
xor U2400 (N_2400,N_1354,N_505);
xor U2401 (N_2401,N_1832,N_1863);
or U2402 (N_2402,N_1351,N_1750);
nand U2403 (N_2403,N_1077,N_457);
nand U2404 (N_2404,N_1764,In_2806);
or U2405 (N_2405,In_411,N_1775);
nor U2406 (N_2406,N_1288,N_216);
and U2407 (N_2407,N_1777,N_1425);
nand U2408 (N_2408,N_1695,N_971);
xnor U2409 (N_2409,N_1890,N_1744);
or U2410 (N_2410,N_1870,N_1624);
and U2411 (N_2411,In_2364,In_920);
nand U2412 (N_2412,N_1860,N_1522);
and U2413 (N_2413,In_2199,N_1555);
nor U2414 (N_2414,N_1608,N_1669);
nor U2415 (N_2415,N_1540,N_1315);
nand U2416 (N_2416,N_1638,In_1565);
or U2417 (N_2417,N_1134,N_1943);
or U2418 (N_2418,N_1514,N_1517);
nor U2419 (N_2419,N_1544,N_1541);
nand U2420 (N_2420,In_2204,In_1640);
and U2421 (N_2421,N_1611,N_1704);
and U2422 (N_2422,N_1776,N_300);
xnor U2423 (N_2423,In_1206,In_1619);
or U2424 (N_2424,N_1840,N_1878);
and U2425 (N_2425,N_328,N_775);
nor U2426 (N_2426,N_1231,In_308);
nand U2427 (N_2427,N_1843,N_1718);
and U2428 (N_2428,N_1852,N_1110);
nor U2429 (N_2429,N_1814,N_978);
nor U2430 (N_2430,In_502,N_1095);
or U2431 (N_2431,N_1766,N_1696);
and U2432 (N_2432,N_1975,N_1587);
nor U2433 (N_2433,N_1553,N_1853);
xor U2434 (N_2434,N_650,N_440);
and U2435 (N_2435,N_1659,N_1782);
xnor U2436 (N_2436,In_298,N_1389);
nor U2437 (N_2437,In_1657,N_826);
nor U2438 (N_2438,N_1899,N_1642);
or U2439 (N_2439,In_2100,N_1732);
and U2440 (N_2440,N_1926,N_1965);
xnor U2441 (N_2441,N_1524,N_1850);
nor U2442 (N_2442,N_381,N_1428);
nand U2443 (N_2443,In_2951,N_1885);
nor U2444 (N_2444,N_274,N_1609);
xnor U2445 (N_2445,In_2448,N_1572);
xor U2446 (N_2446,N_1605,N_1568);
or U2447 (N_2447,N_1858,N_1841);
xor U2448 (N_2448,N_1535,N_662);
and U2449 (N_2449,N_1769,In_1893);
xor U2450 (N_2450,N_1968,N_1641);
xor U2451 (N_2451,In_2503,N_530);
and U2452 (N_2452,N_1601,N_1407);
xnor U2453 (N_2453,N_1623,N_1554);
nand U2454 (N_2454,N_1820,N_940);
nand U2455 (N_2455,N_1941,N_1579);
nand U2456 (N_2456,In_2660,In_2623);
and U2457 (N_2457,N_1833,In_1899);
nor U2458 (N_2458,N_1473,N_1937);
or U2459 (N_2459,N_916,N_1355);
xnor U2460 (N_2460,N_1575,N_341);
and U2461 (N_2461,In_1676,N_1662);
and U2462 (N_2462,N_1475,N_410);
nand U2463 (N_2463,N_400,N_1559);
nand U2464 (N_2464,N_1996,N_1956);
xor U2465 (N_2465,N_1974,N_941);
xor U2466 (N_2466,N_1824,N_1156);
and U2467 (N_2467,In_1135,In_1749);
and U2468 (N_2468,N_1760,In_1939);
or U2469 (N_2469,N_1106,In_2331);
xor U2470 (N_2470,N_841,N_1677);
and U2471 (N_2471,N_1387,N_1266);
nor U2472 (N_2472,N_1160,In_1910);
and U2473 (N_2473,In_1038,N_1215);
nor U2474 (N_2474,N_310,N_1909);
nand U2475 (N_2475,In_2882,In_859);
and U2476 (N_2476,N_1621,In_2912);
nor U2477 (N_2477,N_1329,In_738);
or U2478 (N_2478,N_418,N_1877);
xnor U2479 (N_2479,N_1567,In_198);
or U2480 (N_2480,N_1729,N_1978);
and U2481 (N_2481,N_1984,N_1044);
nand U2482 (N_2482,N_1302,N_1253);
xnor U2483 (N_2483,N_1604,In_941);
and U2484 (N_2484,N_1952,In_296);
xnor U2485 (N_2485,N_1961,In_1740);
nand U2486 (N_2486,N_1904,N_1422);
nor U2487 (N_2487,N_1811,N_1827);
and U2488 (N_2488,N_1527,N_1632);
xor U2489 (N_2489,N_1872,N_1643);
and U2490 (N_2490,N_65,N_412);
nand U2491 (N_2491,N_228,N_1420);
nor U2492 (N_2492,N_1265,In_35);
xnor U2493 (N_2493,N_1516,N_1809);
or U2494 (N_2494,N_1883,N_1940);
xnor U2495 (N_2495,N_1526,N_1644);
nand U2496 (N_2496,N_1589,In_1109);
nor U2497 (N_2497,In_1052,N_1945);
xnor U2498 (N_2498,N_1487,N_1192);
xnor U2499 (N_2499,N_1976,N_1668);
and U2500 (N_2500,N_2033,N_2253);
and U2501 (N_2501,N_2173,N_2238);
xnor U2502 (N_2502,N_2326,N_2183);
or U2503 (N_2503,N_2341,N_2276);
or U2504 (N_2504,N_2155,N_2418);
and U2505 (N_2505,N_2289,N_2411);
nor U2506 (N_2506,N_2120,N_2438);
and U2507 (N_2507,N_2452,N_2271);
xnor U2508 (N_2508,N_2085,N_2390);
or U2509 (N_2509,N_2045,N_2479);
nor U2510 (N_2510,N_2021,N_2492);
nor U2511 (N_2511,N_2177,N_2208);
and U2512 (N_2512,N_2082,N_2362);
nor U2513 (N_2513,N_2137,N_2196);
and U2514 (N_2514,N_2039,N_2342);
xor U2515 (N_2515,N_2099,N_2240);
or U2516 (N_2516,N_2234,N_2169);
and U2517 (N_2517,N_2018,N_2496);
nor U2518 (N_2518,N_2201,N_2353);
nor U2519 (N_2519,N_2441,N_2279);
or U2520 (N_2520,N_2393,N_2142);
or U2521 (N_2521,N_2006,N_2288);
nand U2522 (N_2522,N_2159,N_2422);
and U2523 (N_2523,N_2112,N_2087);
or U2524 (N_2524,N_2197,N_2054);
nor U2525 (N_2525,N_2057,N_2325);
nand U2526 (N_2526,N_2221,N_2375);
and U2527 (N_2527,N_2449,N_2491);
nand U2528 (N_2528,N_2048,N_2065);
nor U2529 (N_2529,N_2285,N_2040);
xor U2530 (N_2530,N_2214,N_2030);
nor U2531 (N_2531,N_2320,N_2073);
or U2532 (N_2532,N_2464,N_2321);
or U2533 (N_2533,N_2114,N_2364);
or U2534 (N_2534,N_2058,N_2029);
nand U2535 (N_2535,N_2211,N_2127);
xor U2536 (N_2536,N_2022,N_2306);
nand U2537 (N_2537,N_2494,N_2052);
xor U2538 (N_2538,N_2247,N_2227);
and U2539 (N_2539,N_2350,N_2181);
nand U2540 (N_2540,N_2000,N_2059);
nor U2541 (N_2541,N_2463,N_2144);
xor U2542 (N_2542,N_2194,N_2304);
xor U2543 (N_2543,N_2232,N_2151);
and U2544 (N_2544,N_2445,N_2356);
nand U2545 (N_2545,N_2163,N_2213);
and U2546 (N_2546,N_2161,N_2396);
and U2547 (N_2547,N_2079,N_2458);
nand U2548 (N_2548,N_2074,N_2239);
xnor U2549 (N_2549,N_2269,N_2041);
or U2550 (N_2550,N_2373,N_2091);
nor U2551 (N_2551,N_2335,N_2126);
xor U2552 (N_2552,N_2190,N_2435);
or U2553 (N_2553,N_2005,N_2402);
nor U2554 (N_2554,N_2345,N_2188);
xor U2555 (N_2555,N_2186,N_2361);
nor U2556 (N_2556,N_2377,N_2410);
nor U2557 (N_2557,N_2358,N_2062);
nand U2558 (N_2558,N_2466,N_2078);
or U2559 (N_2559,N_2106,N_2277);
and U2560 (N_2560,N_2031,N_2296);
or U2561 (N_2561,N_2017,N_2193);
nor U2562 (N_2562,N_2158,N_2164);
and U2563 (N_2563,N_2272,N_2412);
nor U2564 (N_2564,N_2318,N_2268);
nand U2565 (N_2565,N_2104,N_2135);
or U2566 (N_2566,N_2439,N_2050);
and U2567 (N_2567,N_2488,N_2053);
xnor U2568 (N_2568,N_2243,N_2471);
nor U2569 (N_2569,N_2171,N_2357);
or U2570 (N_2570,N_2266,N_2365);
or U2571 (N_2571,N_2367,N_2076);
nand U2572 (N_2572,N_2185,N_2477);
xor U2573 (N_2573,N_2308,N_2472);
nor U2574 (N_2574,N_2119,N_2003);
and U2575 (N_2575,N_2111,N_2363);
xnor U2576 (N_2576,N_2340,N_2475);
and U2577 (N_2577,N_2148,N_2386);
and U2578 (N_2578,N_2343,N_2069);
nor U2579 (N_2579,N_2369,N_2245);
xnor U2580 (N_2580,N_2001,N_2476);
xor U2581 (N_2581,N_2176,N_2336);
nand U2582 (N_2582,N_2132,N_2225);
or U2583 (N_2583,N_2486,N_2125);
or U2584 (N_2584,N_2218,N_2376);
and U2585 (N_2585,N_2314,N_2408);
and U2586 (N_2586,N_2372,N_2292);
or U2587 (N_2587,N_2401,N_2224);
nand U2588 (N_2588,N_2027,N_2019);
nand U2589 (N_2589,N_2419,N_2397);
or U2590 (N_2590,N_2293,N_2013);
nor U2591 (N_2591,N_2089,N_2425);
and U2592 (N_2592,N_2102,N_2140);
or U2593 (N_2593,N_2175,N_2436);
or U2594 (N_2594,N_2283,N_2299);
nand U2595 (N_2595,N_2042,N_2080);
and U2596 (N_2596,N_2117,N_2428);
and U2597 (N_2597,N_2023,N_2311);
or U2598 (N_2598,N_2490,N_2007);
and U2599 (N_2599,N_2061,N_2448);
nand U2600 (N_2600,N_2028,N_2354);
nor U2601 (N_2601,N_2374,N_2118);
or U2602 (N_2602,N_2179,N_2067);
and U2603 (N_2603,N_2322,N_2382);
nor U2604 (N_2604,N_2160,N_2098);
nand U2605 (N_2605,N_2399,N_2414);
nand U2606 (N_2606,N_2295,N_2116);
nand U2607 (N_2607,N_2010,N_2313);
nand U2608 (N_2608,N_2205,N_2170);
or U2609 (N_2609,N_2047,N_2310);
or U2610 (N_2610,N_2286,N_2199);
nand U2611 (N_2611,N_2407,N_2433);
nand U2612 (N_2612,N_2038,N_2035);
nor U2613 (N_2613,N_2037,N_2260);
or U2614 (N_2614,N_2011,N_2474);
or U2615 (N_2615,N_2478,N_2424);
or U2616 (N_2616,N_2025,N_2481);
nor U2617 (N_2617,N_2191,N_2446);
or U2618 (N_2618,N_2133,N_2338);
or U2619 (N_2619,N_2219,N_2157);
xnor U2620 (N_2620,N_2290,N_2398);
nor U2621 (N_2621,N_2257,N_2090);
nand U2622 (N_2622,N_2060,N_2432);
and U2623 (N_2623,N_2131,N_2495);
or U2624 (N_2624,N_2317,N_2444);
nor U2625 (N_2625,N_2235,N_2404);
nand U2626 (N_2626,N_2145,N_2055);
and U2627 (N_2627,N_2077,N_2002);
nor U2628 (N_2628,N_2450,N_2141);
nand U2629 (N_2629,N_2459,N_2044);
nand U2630 (N_2630,N_2200,N_2451);
xnor U2631 (N_2631,N_2294,N_2093);
nand U2632 (N_2632,N_2154,N_2207);
nand U2633 (N_2633,N_2046,N_2440);
or U2634 (N_2634,N_2259,N_2330);
and U2635 (N_2635,N_2113,N_2282);
or U2636 (N_2636,N_2278,N_2136);
nand U2637 (N_2637,N_2122,N_2456);
nand U2638 (N_2638,N_2216,N_2437);
nor U2639 (N_2639,N_2334,N_2258);
nor U2640 (N_2640,N_2182,N_2034);
nor U2641 (N_2641,N_2291,N_2051);
nor U2642 (N_2642,N_2101,N_2187);
nor U2643 (N_2643,N_2248,N_2056);
and U2644 (N_2644,N_2236,N_2300);
nor U2645 (N_2645,N_2230,N_2360);
and U2646 (N_2646,N_2265,N_2231);
nor U2647 (N_2647,N_2139,N_2264);
or U2648 (N_2648,N_2071,N_2379);
nor U2649 (N_2649,N_2426,N_2442);
nand U2650 (N_2650,N_2315,N_2233);
xor U2651 (N_2651,N_2489,N_2094);
nand U2652 (N_2652,N_2096,N_2174);
nand U2653 (N_2653,N_2487,N_2166);
or U2654 (N_2654,N_2123,N_2406);
and U2655 (N_2655,N_2332,N_2128);
or U2656 (N_2656,N_2012,N_2206);
nand U2657 (N_2657,N_2391,N_2454);
nor U2658 (N_2658,N_2134,N_2388);
or U2659 (N_2659,N_2072,N_2327);
or U2660 (N_2660,N_2121,N_2172);
or U2661 (N_2661,N_2246,N_2380);
nand U2662 (N_2662,N_2331,N_2480);
xor U2663 (N_2663,N_2337,N_2431);
and U2664 (N_2664,N_2413,N_2270);
nor U2665 (N_2665,N_2430,N_2081);
nor U2666 (N_2666,N_2405,N_2415);
or U2667 (N_2667,N_2150,N_2009);
xnor U2668 (N_2668,N_2349,N_2149);
and U2669 (N_2669,N_2324,N_2064);
nor U2670 (N_2670,N_2036,N_2394);
and U2671 (N_2671,N_2355,N_2015);
nand U2672 (N_2672,N_2403,N_2274);
and U2673 (N_2673,N_2366,N_2319);
nor U2674 (N_2674,N_2075,N_2420);
or U2675 (N_2675,N_2129,N_2223);
xnor U2676 (N_2676,N_2146,N_2004);
nor U2677 (N_2677,N_2251,N_2421);
xnor U2678 (N_2678,N_2095,N_2086);
nand U2679 (N_2679,N_2016,N_2088);
and U2680 (N_2680,N_2287,N_2470);
xnor U2681 (N_2681,N_2305,N_2469);
and U2682 (N_2682,N_2254,N_2184);
or U2683 (N_2683,N_2180,N_2312);
nand U2684 (N_2684,N_2465,N_2153);
or U2685 (N_2685,N_2329,N_2392);
nand U2686 (N_2686,N_2237,N_2309);
or U2687 (N_2687,N_2302,N_2109);
and U2688 (N_2688,N_2417,N_2100);
nor U2689 (N_2689,N_2255,N_2195);
nand U2690 (N_2690,N_2473,N_2165);
nand U2691 (N_2691,N_2250,N_2348);
nand U2692 (N_2692,N_2307,N_2152);
nand U2693 (N_2693,N_2267,N_2462);
xor U2694 (N_2694,N_2162,N_2143);
and U2695 (N_2695,N_2378,N_2226);
or U2696 (N_2696,N_2359,N_2498);
nor U2697 (N_2697,N_2273,N_2383);
and U2698 (N_2698,N_2178,N_2263);
or U2699 (N_2699,N_2387,N_2108);
and U2700 (N_2700,N_2229,N_2499);
or U2701 (N_2701,N_2138,N_2423);
xnor U2702 (N_2702,N_2261,N_2284);
and U2703 (N_2703,N_2014,N_2147);
xor U2704 (N_2704,N_2351,N_2124);
or U2705 (N_2705,N_2217,N_2066);
nand U2706 (N_2706,N_2210,N_2241);
or U2707 (N_2707,N_2275,N_2222);
xnor U2708 (N_2708,N_2156,N_2097);
nor U2709 (N_2709,N_2434,N_2083);
nor U2710 (N_2710,N_2242,N_2228);
nor U2711 (N_2711,N_2385,N_2352);
xnor U2712 (N_2712,N_2384,N_2020);
nand U2713 (N_2713,N_2482,N_2468);
xnor U2714 (N_2714,N_2460,N_2297);
and U2715 (N_2715,N_2068,N_2280);
nand U2716 (N_2716,N_2070,N_2301);
nor U2717 (N_2717,N_2103,N_2008);
and U2718 (N_2718,N_2262,N_2107);
xnor U2719 (N_2719,N_2344,N_2092);
and U2720 (N_2720,N_2429,N_2453);
nor U2721 (N_2721,N_2281,N_2447);
and U2722 (N_2722,N_2400,N_2333);
and U2723 (N_2723,N_2368,N_2209);
or U2724 (N_2724,N_2130,N_2497);
xor U2725 (N_2725,N_2202,N_2167);
and U2726 (N_2726,N_2370,N_2416);
or U2727 (N_2727,N_2105,N_2484);
and U2728 (N_2728,N_2457,N_2256);
xor U2729 (N_2729,N_2461,N_2043);
or U2730 (N_2730,N_2168,N_2409);
nand U2731 (N_2731,N_2189,N_2249);
nor U2732 (N_2732,N_2347,N_2493);
nor U2733 (N_2733,N_2316,N_2427);
or U2734 (N_2734,N_2328,N_2049);
and U2735 (N_2735,N_2252,N_2024);
or U2736 (N_2736,N_2212,N_2220);
or U2737 (N_2737,N_2204,N_2395);
and U2738 (N_2738,N_2026,N_2485);
nand U2739 (N_2739,N_2443,N_2215);
xnor U2740 (N_2740,N_2371,N_2389);
or U2741 (N_2741,N_2192,N_2346);
or U2742 (N_2742,N_2110,N_2063);
or U2743 (N_2743,N_2244,N_2339);
xnor U2744 (N_2744,N_2323,N_2455);
nor U2745 (N_2745,N_2467,N_2032);
nand U2746 (N_2746,N_2298,N_2203);
xnor U2747 (N_2747,N_2483,N_2303);
xor U2748 (N_2748,N_2381,N_2198);
nor U2749 (N_2749,N_2115,N_2084);
nor U2750 (N_2750,N_2280,N_2221);
nand U2751 (N_2751,N_2004,N_2398);
and U2752 (N_2752,N_2169,N_2453);
and U2753 (N_2753,N_2238,N_2102);
and U2754 (N_2754,N_2324,N_2255);
xnor U2755 (N_2755,N_2143,N_2478);
xnor U2756 (N_2756,N_2270,N_2345);
xnor U2757 (N_2757,N_2182,N_2128);
xor U2758 (N_2758,N_2177,N_2084);
and U2759 (N_2759,N_2118,N_2325);
or U2760 (N_2760,N_2121,N_2076);
and U2761 (N_2761,N_2123,N_2137);
nor U2762 (N_2762,N_2224,N_2428);
or U2763 (N_2763,N_2469,N_2013);
xor U2764 (N_2764,N_2420,N_2273);
and U2765 (N_2765,N_2094,N_2223);
nand U2766 (N_2766,N_2108,N_2085);
nand U2767 (N_2767,N_2292,N_2279);
xnor U2768 (N_2768,N_2207,N_2151);
xor U2769 (N_2769,N_2330,N_2099);
or U2770 (N_2770,N_2211,N_2232);
nor U2771 (N_2771,N_2411,N_2053);
nor U2772 (N_2772,N_2410,N_2329);
and U2773 (N_2773,N_2095,N_2034);
xnor U2774 (N_2774,N_2117,N_2407);
or U2775 (N_2775,N_2001,N_2184);
nor U2776 (N_2776,N_2111,N_2373);
xnor U2777 (N_2777,N_2354,N_2335);
xor U2778 (N_2778,N_2452,N_2009);
and U2779 (N_2779,N_2165,N_2077);
nor U2780 (N_2780,N_2153,N_2081);
xnor U2781 (N_2781,N_2320,N_2463);
nand U2782 (N_2782,N_2461,N_2486);
xnor U2783 (N_2783,N_2005,N_2070);
nand U2784 (N_2784,N_2468,N_2313);
xor U2785 (N_2785,N_2357,N_2043);
or U2786 (N_2786,N_2394,N_2056);
and U2787 (N_2787,N_2488,N_2484);
or U2788 (N_2788,N_2498,N_2360);
xor U2789 (N_2789,N_2060,N_2409);
and U2790 (N_2790,N_2127,N_2482);
xnor U2791 (N_2791,N_2259,N_2208);
nand U2792 (N_2792,N_2033,N_2323);
xor U2793 (N_2793,N_2267,N_2469);
nand U2794 (N_2794,N_2352,N_2304);
nor U2795 (N_2795,N_2383,N_2098);
nand U2796 (N_2796,N_2036,N_2490);
nor U2797 (N_2797,N_2423,N_2046);
or U2798 (N_2798,N_2053,N_2434);
xnor U2799 (N_2799,N_2422,N_2210);
nand U2800 (N_2800,N_2408,N_2044);
nand U2801 (N_2801,N_2100,N_2288);
nand U2802 (N_2802,N_2449,N_2267);
nor U2803 (N_2803,N_2452,N_2034);
or U2804 (N_2804,N_2292,N_2177);
and U2805 (N_2805,N_2466,N_2329);
or U2806 (N_2806,N_2334,N_2091);
nor U2807 (N_2807,N_2267,N_2383);
nor U2808 (N_2808,N_2051,N_2466);
nand U2809 (N_2809,N_2150,N_2476);
nor U2810 (N_2810,N_2454,N_2076);
nand U2811 (N_2811,N_2077,N_2138);
xor U2812 (N_2812,N_2096,N_2378);
and U2813 (N_2813,N_2201,N_2160);
nor U2814 (N_2814,N_2139,N_2476);
or U2815 (N_2815,N_2326,N_2416);
nor U2816 (N_2816,N_2347,N_2155);
nand U2817 (N_2817,N_2294,N_2006);
nor U2818 (N_2818,N_2313,N_2269);
and U2819 (N_2819,N_2360,N_2307);
or U2820 (N_2820,N_2445,N_2233);
or U2821 (N_2821,N_2469,N_2404);
nand U2822 (N_2822,N_2413,N_2017);
and U2823 (N_2823,N_2268,N_2259);
or U2824 (N_2824,N_2401,N_2474);
or U2825 (N_2825,N_2000,N_2072);
nor U2826 (N_2826,N_2086,N_2352);
xnor U2827 (N_2827,N_2171,N_2400);
nor U2828 (N_2828,N_2120,N_2093);
and U2829 (N_2829,N_2176,N_2353);
and U2830 (N_2830,N_2318,N_2215);
nor U2831 (N_2831,N_2132,N_2196);
and U2832 (N_2832,N_2267,N_2095);
and U2833 (N_2833,N_2139,N_2111);
and U2834 (N_2834,N_2318,N_2213);
nand U2835 (N_2835,N_2397,N_2486);
nor U2836 (N_2836,N_2364,N_2107);
nor U2837 (N_2837,N_2028,N_2171);
nor U2838 (N_2838,N_2471,N_2277);
xnor U2839 (N_2839,N_2177,N_2385);
and U2840 (N_2840,N_2065,N_2070);
xnor U2841 (N_2841,N_2336,N_2414);
and U2842 (N_2842,N_2214,N_2419);
nor U2843 (N_2843,N_2433,N_2194);
and U2844 (N_2844,N_2339,N_2179);
or U2845 (N_2845,N_2134,N_2362);
and U2846 (N_2846,N_2314,N_2274);
nand U2847 (N_2847,N_2347,N_2075);
and U2848 (N_2848,N_2450,N_2127);
nand U2849 (N_2849,N_2488,N_2296);
nand U2850 (N_2850,N_2362,N_2079);
and U2851 (N_2851,N_2079,N_2212);
or U2852 (N_2852,N_2483,N_2376);
and U2853 (N_2853,N_2256,N_2274);
or U2854 (N_2854,N_2300,N_2355);
nor U2855 (N_2855,N_2401,N_2369);
xor U2856 (N_2856,N_2340,N_2421);
or U2857 (N_2857,N_2050,N_2056);
nor U2858 (N_2858,N_2135,N_2101);
nor U2859 (N_2859,N_2017,N_2195);
or U2860 (N_2860,N_2126,N_2026);
nand U2861 (N_2861,N_2455,N_2368);
nand U2862 (N_2862,N_2477,N_2325);
or U2863 (N_2863,N_2351,N_2326);
nand U2864 (N_2864,N_2273,N_2208);
and U2865 (N_2865,N_2293,N_2172);
nand U2866 (N_2866,N_2012,N_2104);
or U2867 (N_2867,N_2162,N_2235);
or U2868 (N_2868,N_2140,N_2125);
and U2869 (N_2869,N_2114,N_2068);
or U2870 (N_2870,N_2008,N_2115);
nor U2871 (N_2871,N_2273,N_2436);
and U2872 (N_2872,N_2047,N_2080);
or U2873 (N_2873,N_2197,N_2004);
nor U2874 (N_2874,N_2057,N_2099);
nand U2875 (N_2875,N_2469,N_2122);
and U2876 (N_2876,N_2421,N_2323);
xor U2877 (N_2877,N_2248,N_2060);
or U2878 (N_2878,N_2043,N_2229);
or U2879 (N_2879,N_2486,N_2450);
or U2880 (N_2880,N_2004,N_2037);
nand U2881 (N_2881,N_2198,N_2094);
or U2882 (N_2882,N_2293,N_2192);
xor U2883 (N_2883,N_2196,N_2487);
and U2884 (N_2884,N_2425,N_2286);
xnor U2885 (N_2885,N_2409,N_2038);
xor U2886 (N_2886,N_2066,N_2215);
nor U2887 (N_2887,N_2048,N_2495);
or U2888 (N_2888,N_2120,N_2207);
and U2889 (N_2889,N_2174,N_2030);
and U2890 (N_2890,N_2038,N_2326);
nand U2891 (N_2891,N_2048,N_2154);
xor U2892 (N_2892,N_2198,N_2010);
and U2893 (N_2893,N_2235,N_2290);
xor U2894 (N_2894,N_2048,N_2300);
nor U2895 (N_2895,N_2286,N_2344);
xnor U2896 (N_2896,N_2433,N_2402);
or U2897 (N_2897,N_2489,N_2085);
nand U2898 (N_2898,N_2341,N_2329);
nor U2899 (N_2899,N_2477,N_2063);
nand U2900 (N_2900,N_2319,N_2431);
nand U2901 (N_2901,N_2367,N_2433);
xnor U2902 (N_2902,N_2426,N_2254);
or U2903 (N_2903,N_2139,N_2391);
or U2904 (N_2904,N_2091,N_2390);
nor U2905 (N_2905,N_2180,N_2021);
nor U2906 (N_2906,N_2412,N_2341);
or U2907 (N_2907,N_2138,N_2333);
nand U2908 (N_2908,N_2032,N_2305);
nor U2909 (N_2909,N_2219,N_2326);
or U2910 (N_2910,N_2338,N_2200);
nand U2911 (N_2911,N_2329,N_2180);
or U2912 (N_2912,N_2040,N_2335);
xnor U2913 (N_2913,N_2444,N_2238);
xnor U2914 (N_2914,N_2463,N_2378);
xor U2915 (N_2915,N_2386,N_2375);
nor U2916 (N_2916,N_2465,N_2493);
and U2917 (N_2917,N_2313,N_2413);
xor U2918 (N_2918,N_2184,N_2035);
nor U2919 (N_2919,N_2294,N_2326);
xor U2920 (N_2920,N_2022,N_2359);
and U2921 (N_2921,N_2415,N_2377);
and U2922 (N_2922,N_2402,N_2368);
or U2923 (N_2923,N_2128,N_2031);
nor U2924 (N_2924,N_2479,N_2122);
and U2925 (N_2925,N_2129,N_2027);
nand U2926 (N_2926,N_2075,N_2226);
or U2927 (N_2927,N_2409,N_2344);
nor U2928 (N_2928,N_2311,N_2087);
xor U2929 (N_2929,N_2154,N_2063);
xnor U2930 (N_2930,N_2166,N_2258);
and U2931 (N_2931,N_2057,N_2380);
nor U2932 (N_2932,N_2382,N_2277);
nor U2933 (N_2933,N_2277,N_2332);
and U2934 (N_2934,N_2345,N_2090);
and U2935 (N_2935,N_2383,N_2459);
and U2936 (N_2936,N_2459,N_2289);
and U2937 (N_2937,N_2471,N_2206);
or U2938 (N_2938,N_2344,N_2400);
and U2939 (N_2939,N_2472,N_2197);
nor U2940 (N_2940,N_2337,N_2359);
xor U2941 (N_2941,N_2114,N_2216);
nand U2942 (N_2942,N_2073,N_2000);
or U2943 (N_2943,N_2223,N_2485);
nand U2944 (N_2944,N_2014,N_2475);
or U2945 (N_2945,N_2379,N_2200);
and U2946 (N_2946,N_2228,N_2213);
or U2947 (N_2947,N_2489,N_2360);
nand U2948 (N_2948,N_2031,N_2237);
xnor U2949 (N_2949,N_2144,N_2145);
xor U2950 (N_2950,N_2181,N_2414);
nor U2951 (N_2951,N_2419,N_2376);
and U2952 (N_2952,N_2136,N_2197);
nor U2953 (N_2953,N_2170,N_2452);
or U2954 (N_2954,N_2344,N_2422);
or U2955 (N_2955,N_2140,N_2261);
or U2956 (N_2956,N_2301,N_2213);
xnor U2957 (N_2957,N_2325,N_2066);
or U2958 (N_2958,N_2093,N_2086);
xor U2959 (N_2959,N_2379,N_2133);
nand U2960 (N_2960,N_2155,N_2343);
nor U2961 (N_2961,N_2192,N_2021);
nand U2962 (N_2962,N_2370,N_2354);
or U2963 (N_2963,N_2473,N_2299);
nor U2964 (N_2964,N_2370,N_2194);
nor U2965 (N_2965,N_2021,N_2319);
and U2966 (N_2966,N_2480,N_2239);
and U2967 (N_2967,N_2170,N_2300);
or U2968 (N_2968,N_2183,N_2467);
or U2969 (N_2969,N_2409,N_2040);
xnor U2970 (N_2970,N_2193,N_2091);
or U2971 (N_2971,N_2393,N_2050);
nor U2972 (N_2972,N_2305,N_2219);
and U2973 (N_2973,N_2332,N_2431);
and U2974 (N_2974,N_2212,N_2169);
or U2975 (N_2975,N_2197,N_2035);
nand U2976 (N_2976,N_2291,N_2375);
and U2977 (N_2977,N_2028,N_2018);
and U2978 (N_2978,N_2132,N_2029);
xnor U2979 (N_2979,N_2157,N_2436);
and U2980 (N_2980,N_2252,N_2145);
or U2981 (N_2981,N_2240,N_2429);
nand U2982 (N_2982,N_2455,N_2371);
nand U2983 (N_2983,N_2448,N_2170);
nor U2984 (N_2984,N_2059,N_2197);
nor U2985 (N_2985,N_2385,N_2018);
or U2986 (N_2986,N_2121,N_2174);
nor U2987 (N_2987,N_2387,N_2004);
nand U2988 (N_2988,N_2145,N_2126);
and U2989 (N_2989,N_2203,N_2127);
nor U2990 (N_2990,N_2249,N_2314);
or U2991 (N_2991,N_2219,N_2224);
nand U2992 (N_2992,N_2267,N_2114);
nand U2993 (N_2993,N_2221,N_2242);
nand U2994 (N_2994,N_2276,N_2205);
and U2995 (N_2995,N_2347,N_2092);
nand U2996 (N_2996,N_2333,N_2385);
and U2997 (N_2997,N_2022,N_2310);
and U2998 (N_2998,N_2478,N_2323);
and U2999 (N_2999,N_2426,N_2088);
and U3000 (N_3000,N_2680,N_2952);
nor U3001 (N_3001,N_2571,N_2934);
nor U3002 (N_3002,N_2697,N_2693);
nor U3003 (N_3003,N_2899,N_2734);
nor U3004 (N_3004,N_2913,N_2821);
nand U3005 (N_3005,N_2553,N_2735);
xnor U3006 (N_3006,N_2590,N_2521);
nand U3007 (N_3007,N_2600,N_2976);
nor U3008 (N_3008,N_2798,N_2831);
nor U3009 (N_3009,N_2878,N_2668);
nand U3010 (N_3010,N_2621,N_2835);
xor U3011 (N_3011,N_2613,N_2716);
or U3012 (N_3012,N_2961,N_2933);
or U3013 (N_3013,N_2591,N_2706);
xor U3014 (N_3014,N_2917,N_2622);
or U3015 (N_3015,N_2906,N_2566);
nor U3016 (N_3016,N_2596,N_2719);
nor U3017 (N_3017,N_2903,N_2788);
or U3018 (N_3018,N_2604,N_2919);
and U3019 (N_3019,N_2850,N_2580);
and U3020 (N_3020,N_2760,N_2931);
and U3021 (N_3021,N_2500,N_2864);
and U3022 (N_3022,N_2843,N_2807);
and U3023 (N_3023,N_2890,N_2990);
xnor U3024 (N_3024,N_2897,N_2721);
nor U3025 (N_3025,N_2692,N_2809);
nand U3026 (N_3026,N_2649,N_2808);
nand U3027 (N_3027,N_2993,N_2607);
nand U3028 (N_3028,N_2524,N_2756);
nand U3029 (N_3029,N_2516,N_2767);
nor U3030 (N_3030,N_2520,N_2626);
and U3031 (N_3031,N_2761,N_2551);
and U3032 (N_3032,N_2802,N_2603);
and U3033 (N_3033,N_2606,N_2656);
or U3034 (N_3034,N_2836,N_2558);
or U3035 (N_3035,N_2766,N_2886);
and U3036 (N_3036,N_2855,N_2661);
or U3037 (N_3037,N_2646,N_2686);
or U3038 (N_3038,N_2550,N_2689);
or U3039 (N_3039,N_2896,N_2823);
and U3040 (N_3040,N_2773,N_2667);
nand U3041 (N_3041,N_2912,N_2800);
nor U3042 (N_3042,N_2617,N_2932);
nand U3043 (N_3043,N_2926,N_2837);
or U3044 (N_3044,N_2778,N_2819);
nor U3045 (N_3045,N_2842,N_2510);
nor U3046 (N_3046,N_2943,N_2775);
nor U3047 (N_3047,N_2883,N_2794);
xor U3048 (N_3048,N_2841,N_2895);
and U3049 (N_3049,N_2724,N_2793);
xor U3050 (N_3050,N_2951,N_2738);
and U3051 (N_3051,N_2705,N_2691);
nor U3052 (N_3052,N_2753,N_2790);
xor U3053 (N_3053,N_2568,N_2810);
nand U3054 (N_3054,N_2945,N_2955);
nor U3055 (N_3055,N_2511,N_2923);
or U3056 (N_3056,N_2629,N_2700);
nor U3057 (N_3057,N_2844,N_2789);
nor U3058 (N_3058,N_2556,N_2829);
nand U3059 (N_3059,N_2666,N_2662);
nor U3060 (N_3060,N_2852,N_2665);
or U3061 (N_3061,N_2517,N_2805);
and U3062 (N_3062,N_2612,N_2598);
and U3063 (N_3063,N_2901,N_2542);
xnor U3064 (N_3064,N_2688,N_2927);
nor U3065 (N_3065,N_2948,N_2824);
nor U3066 (N_3066,N_2815,N_2935);
or U3067 (N_3067,N_2969,N_2696);
xor U3068 (N_3068,N_2588,N_2676);
xor U3069 (N_3069,N_2817,N_2527);
and U3070 (N_3070,N_2546,N_2732);
nor U3071 (N_3071,N_2519,N_2728);
nand U3072 (N_3072,N_2783,N_2543);
xor U3073 (N_3073,N_2674,N_2533);
nor U3074 (N_3074,N_2583,N_2547);
nand U3075 (N_3075,N_2988,N_2536);
nor U3076 (N_3076,N_2655,N_2509);
and U3077 (N_3077,N_2982,N_2981);
nand U3078 (N_3078,N_2914,N_2586);
and U3079 (N_3079,N_2576,N_2502);
xnor U3080 (N_3080,N_2960,N_2538);
or U3081 (N_3081,N_2838,N_2845);
xor U3082 (N_3082,N_2949,N_2544);
and U3083 (N_3083,N_2675,N_2745);
or U3084 (N_3084,N_2698,N_2594);
nand U3085 (N_3085,N_2880,N_2652);
and U3086 (N_3086,N_2518,N_2818);
nand U3087 (N_3087,N_2907,N_2900);
and U3088 (N_3088,N_2846,N_2638);
xor U3089 (N_3089,N_2685,N_2814);
and U3090 (N_3090,N_2643,N_2560);
nand U3091 (N_3091,N_2953,N_2534);
nand U3092 (N_3092,N_2859,N_2565);
nor U3093 (N_3093,N_2757,N_2763);
nand U3094 (N_3094,N_2820,N_2701);
and U3095 (N_3095,N_2862,N_2531);
nor U3096 (N_3096,N_2507,N_2740);
nand U3097 (N_3097,N_2867,N_2530);
nor U3098 (N_3098,N_2780,N_2523);
nand U3099 (N_3099,N_2879,N_2541);
or U3100 (N_3100,N_2968,N_2991);
or U3101 (N_3101,N_2540,N_2548);
or U3102 (N_3102,N_2937,N_2659);
nand U3103 (N_3103,N_2731,N_2830);
xor U3104 (N_3104,N_2825,N_2506);
nor U3105 (N_3105,N_2634,N_2645);
nand U3106 (N_3106,N_2816,N_2853);
or U3107 (N_3107,N_2671,N_2592);
and U3108 (N_3108,N_2654,N_2958);
and U3109 (N_3109,N_2641,N_2796);
or U3110 (N_3110,N_2909,N_2737);
xnor U3111 (N_3111,N_2888,N_2751);
nor U3112 (N_3112,N_2752,N_2625);
and U3113 (N_3113,N_2552,N_2749);
or U3114 (N_3114,N_2683,N_2774);
xor U3115 (N_3115,N_2669,N_2562);
nand U3116 (N_3116,N_2574,N_2729);
nand U3117 (N_3117,N_2681,N_2615);
or U3118 (N_3118,N_2918,N_2563);
nand U3119 (N_3119,N_2595,N_2840);
nand U3120 (N_3120,N_2972,N_2711);
or U3121 (N_3121,N_2985,N_2549);
or U3122 (N_3122,N_2658,N_2730);
and U3123 (N_3123,N_2539,N_2892);
nor U3124 (N_3124,N_2857,N_2827);
nand U3125 (N_3125,N_2522,N_2791);
and U3126 (N_3126,N_2833,N_2602);
nor U3127 (N_3127,N_2723,N_2532);
xor U3128 (N_3128,N_2851,N_2882);
xor U3129 (N_3129,N_2694,N_2860);
nand U3130 (N_3130,N_2922,N_2639);
xnor U3131 (N_3131,N_2806,N_2707);
xor U3132 (N_3132,N_2572,N_2877);
nand U3133 (N_3133,N_2936,N_2505);
nor U3134 (N_3134,N_2647,N_2942);
or U3135 (N_3135,N_2997,N_2679);
and U3136 (N_3136,N_2528,N_2980);
or U3137 (N_3137,N_2725,N_2946);
xnor U3138 (N_3138,N_2770,N_2925);
nor U3139 (N_3139,N_2894,N_2664);
and U3140 (N_3140,N_2584,N_2525);
or U3141 (N_3141,N_2636,N_2944);
or U3142 (N_3142,N_2635,N_2781);
or U3143 (N_3143,N_2742,N_2672);
nor U3144 (N_3144,N_2708,N_2581);
xor U3145 (N_3145,N_2768,N_2983);
xnor U3146 (N_3146,N_2986,N_2736);
nand U3147 (N_3147,N_2627,N_2984);
xor U3148 (N_3148,N_2797,N_2537);
or U3149 (N_3149,N_2573,N_2501);
or U3150 (N_3150,N_2784,N_2630);
xor U3151 (N_3151,N_2526,N_2748);
and U3152 (N_3152,N_2508,N_2966);
xor U3153 (N_3153,N_2994,N_2999);
or U3154 (N_3154,N_2856,N_2564);
and U3155 (N_3155,N_2776,N_2947);
and U3156 (N_3156,N_2908,N_2938);
nor U3157 (N_3157,N_2582,N_2765);
xnor U3158 (N_3158,N_2929,N_2861);
nand U3159 (N_3159,N_2624,N_2759);
nor U3160 (N_3160,N_2799,N_2832);
xor U3161 (N_3161,N_2754,N_2597);
xor U3162 (N_3162,N_2872,N_2561);
and U3163 (N_3163,N_2939,N_2535);
or U3164 (N_3164,N_2812,N_2995);
and U3165 (N_3165,N_2712,N_2803);
or U3166 (N_3166,N_2640,N_2764);
and U3167 (N_3167,N_2839,N_2967);
or U3168 (N_3168,N_2747,N_2924);
or U3169 (N_3169,N_2682,N_2777);
and U3170 (N_3170,N_2915,N_2695);
nand U3171 (N_3171,N_2996,N_2554);
or U3172 (N_3172,N_2620,N_2977);
nand U3173 (N_3173,N_2632,N_2930);
and U3174 (N_3174,N_2755,N_2718);
or U3175 (N_3175,N_2875,N_2762);
xnor U3176 (N_3176,N_2657,N_2964);
xor U3177 (N_3177,N_2889,N_2514);
and U3178 (N_3178,N_2870,N_2989);
xor U3179 (N_3179,N_2921,N_2744);
or U3180 (N_3180,N_2954,N_2717);
nor U3181 (N_3181,N_2578,N_2727);
and U3182 (N_3182,N_2504,N_2605);
or U3183 (N_3183,N_2739,N_2979);
xnor U3184 (N_3184,N_2569,N_2848);
nor U3185 (N_3185,N_2741,N_2710);
xor U3186 (N_3186,N_2699,N_2973);
nor U3187 (N_3187,N_2957,N_2893);
nand U3188 (N_3188,N_2795,N_2904);
or U3189 (N_3189,N_2673,N_2963);
nor U3190 (N_3190,N_2651,N_2813);
nand U3191 (N_3191,N_2720,N_2771);
and U3192 (N_3192,N_2557,N_2920);
nor U3193 (N_3193,N_2503,N_2992);
nand U3194 (N_3194,N_2865,N_2577);
xnor U3195 (N_3195,N_2608,N_2684);
xor U3196 (N_3196,N_2677,N_2847);
or U3197 (N_3197,N_2687,N_2916);
and U3198 (N_3198,N_2704,N_2702);
nand U3199 (N_3199,N_2962,N_2941);
nand U3200 (N_3200,N_2950,N_2690);
and U3201 (N_3201,N_2746,N_2905);
and U3202 (N_3202,N_2902,N_2910);
nand U3203 (N_3203,N_2772,N_2650);
xor U3204 (N_3204,N_2587,N_2792);
xor U3205 (N_3205,N_2599,N_2589);
nor U3206 (N_3206,N_2928,N_2633);
nand U3207 (N_3207,N_2616,N_2970);
nor U3208 (N_3208,N_2786,N_2898);
or U3209 (N_3209,N_2628,N_2849);
nor U3210 (N_3210,N_2758,N_2703);
nor U3211 (N_3211,N_2873,N_2884);
xnor U3212 (N_3212,N_2545,N_2866);
and U3213 (N_3213,N_2822,N_2610);
nand U3214 (N_3214,N_2513,N_2722);
nor U3215 (N_3215,N_2869,N_2974);
and U3216 (N_3216,N_2611,N_2956);
nand U3217 (N_3217,N_2785,N_2750);
or U3218 (N_3218,N_2601,N_2834);
nor U3219 (N_3219,N_2559,N_2678);
nand U3220 (N_3220,N_2868,N_2881);
xor U3221 (N_3221,N_2623,N_2648);
or U3222 (N_3222,N_2512,N_2940);
nand U3223 (N_3223,N_2959,N_2978);
or U3224 (N_3224,N_2911,N_2715);
or U3225 (N_3225,N_2726,N_2971);
nand U3226 (N_3226,N_2631,N_2987);
nand U3227 (N_3227,N_2782,N_2609);
or U3228 (N_3228,N_2828,N_2515);
nand U3229 (N_3229,N_2863,N_2663);
and U3230 (N_3230,N_2779,N_2614);
and U3231 (N_3231,N_2660,N_2804);
xnor U3232 (N_3232,N_2585,N_2801);
and U3233 (N_3233,N_2619,N_2618);
nand U3234 (N_3234,N_2998,N_2743);
or U3235 (N_3235,N_2887,N_2874);
nor U3236 (N_3236,N_2637,N_2670);
nand U3237 (N_3237,N_2891,N_2567);
and U3238 (N_3238,N_2858,N_2714);
or U3239 (N_3239,N_2653,N_2579);
nand U3240 (N_3240,N_2709,N_2644);
and U3241 (N_3241,N_2826,N_2733);
nand U3242 (N_3242,N_2769,N_2642);
xor U3243 (N_3243,N_2871,N_2555);
nor U3244 (N_3244,N_2575,N_2885);
and U3245 (N_3245,N_2965,N_2975);
nor U3246 (N_3246,N_2876,N_2811);
nand U3247 (N_3247,N_2593,N_2529);
xnor U3248 (N_3248,N_2787,N_2570);
nor U3249 (N_3249,N_2713,N_2854);
and U3250 (N_3250,N_2561,N_2865);
nand U3251 (N_3251,N_2660,N_2554);
and U3252 (N_3252,N_2755,N_2790);
nor U3253 (N_3253,N_2869,N_2718);
nor U3254 (N_3254,N_2629,N_2896);
nor U3255 (N_3255,N_2606,N_2593);
nor U3256 (N_3256,N_2807,N_2985);
or U3257 (N_3257,N_2537,N_2819);
xor U3258 (N_3258,N_2509,N_2677);
and U3259 (N_3259,N_2912,N_2688);
xor U3260 (N_3260,N_2938,N_2655);
and U3261 (N_3261,N_2945,N_2883);
xnor U3262 (N_3262,N_2955,N_2847);
and U3263 (N_3263,N_2975,N_2798);
and U3264 (N_3264,N_2779,N_2806);
nor U3265 (N_3265,N_2661,N_2571);
nor U3266 (N_3266,N_2755,N_2738);
and U3267 (N_3267,N_2736,N_2507);
xor U3268 (N_3268,N_2982,N_2621);
xnor U3269 (N_3269,N_2638,N_2841);
xor U3270 (N_3270,N_2676,N_2968);
nor U3271 (N_3271,N_2733,N_2580);
nor U3272 (N_3272,N_2985,N_2980);
and U3273 (N_3273,N_2802,N_2748);
xor U3274 (N_3274,N_2595,N_2811);
nor U3275 (N_3275,N_2856,N_2678);
and U3276 (N_3276,N_2915,N_2990);
or U3277 (N_3277,N_2757,N_2829);
nand U3278 (N_3278,N_2691,N_2695);
or U3279 (N_3279,N_2866,N_2658);
or U3280 (N_3280,N_2948,N_2622);
xor U3281 (N_3281,N_2874,N_2913);
or U3282 (N_3282,N_2567,N_2662);
nand U3283 (N_3283,N_2965,N_2776);
and U3284 (N_3284,N_2627,N_2736);
xnor U3285 (N_3285,N_2933,N_2852);
nand U3286 (N_3286,N_2831,N_2999);
and U3287 (N_3287,N_2532,N_2575);
or U3288 (N_3288,N_2570,N_2989);
nor U3289 (N_3289,N_2619,N_2701);
and U3290 (N_3290,N_2572,N_2923);
nor U3291 (N_3291,N_2567,N_2849);
nor U3292 (N_3292,N_2986,N_2826);
nor U3293 (N_3293,N_2867,N_2854);
nor U3294 (N_3294,N_2527,N_2924);
and U3295 (N_3295,N_2913,N_2681);
xor U3296 (N_3296,N_2685,N_2504);
and U3297 (N_3297,N_2791,N_2829);
or U3298 (N_3298,N_2960,N_2969);
nor U3299 (N_3299,N_2660,N_2869);
or U3300 (N_3300,N_2898,N_2530);
nor U3301 (N_3301,N_2535,N_2793);
nor U3302 (N_3302,N_2553,N_2588);
nor U3303 (N_3303,N_2700,N_2938);
nand U3304 (N_3304,N_2782,N_2500);
nor U3305 (N_3305,N_2679,N_2985);
nand U3306 (N_3306,N_2669,N_2640);
or U3307 (N_3307,N_2989,N_2963);
or U3308 (N_3308,N_2589,N_2943);
nor U3309 (N_3309,N_2526,N_2971);
xnor U3310 (N_3310,N_2658,N_2783);
or U3311 (N_3311,N_2899,N_2754);
nand U3312 (N_3312,N_2743,N_2991);
xor U3313 (N_3313,N_2786,N_2706);
nor U3314 (N_3314,N_2947,N_2795);
nand U3315 (N_3315,N_2686,N_2967);
nand U3316 (N_3316,N_2734,N_2677);
nor U3317 (N_3317,N_2727,N_2630);
and U3318 (N_3318,N_2970,N_2965);
and U3319 (N_3319,N_2625,N_2929);
and U3320 (N_3320,N_2554,N_2732);
xnor U3321 (N_3321,N_2770,N_2768);
nand U3322 (N_3322,N_2595,N_2553);
or U3323 (N_3323,N_2935,N_2523);
or U3324 (N_3324,N_2630,N_2773);
nand U3325 (N_3325,N_2796,N_2782);
nand U3326 (N_3326,N_2727,N_2700);
nor U3327 (N_3327,N_2906,N_2568);
xnor U3328 (N_3328,N_2720,N_2715);
xnor U3329 (N_3329,N_2921,N_2653);
xor U3330 (N_3330,N_2691,N_2572);
and U3331 (N_3331,N_2827,N_2972);
or U3332 (N_3332,N_2761,N_2547);
xor U3333 (N_3333,N_2686,N_2728);
xnor U3334 (N_3334,N_2564,N_2572);
xnor U3335 (N_3335,N_2581,N_2786);
xor U3336 (N_3336,N_2579,N_2809);
xor U3337 (N_3337,N_2905,N_2858);
or U3338 (N_3338,N_2768,N_2650);
nor U3339 (N_3339,N_2935,N_2789);
nand U3340 (N_3340,N_2982,N_2810);
xnor U3341 (N_3341,N_2546,N_2630);
or U3342 (N_3342,N_2768,N_2893);
nand U3343 (N_3343,N_2708,N_2826);
nor U3344 (N_3344,N_2695,N_2890);
or U3345 (N_3345,N_2513,N_2757);
nand U3346 (N_3346,N_2708,N_2984);
or U3347 (N_3347,N_2632,N_2782);
nand U3348 (N_3348,N_2799,N_2833);
nand U3349 (N_3349,N_2999,N_2715);
nor U3350 (N_3350,N_2729,N_2718);
nor U3351 (N_3351,N_2586,N_2833);
xnor U3352 (N_3352,N_2769,N_2951);
nand U3353 (N_3353,N_2921,N_2668);
and U3354 (N_3354,N_2758,N_2527);
and U3355 (N_3355,N_2568,N_2821);
xnor U3356 (N_3356,N_2819,N_2618);
and U3357 (N_3357,N_2670,N_2786);
and U3358 (N_3358,N_2680,N_2949);
and U3359 (N_3359,N_2650,N_2878);
xor U3360 (N_3360,N_2841,N_2597);
nor U3361 (N_3361,N_2609,N_2597);
and U3362 (N_3362,N_2839,N_2665);
nor U3363 (N_3363,N_2781,N_2502);
nor U3364 (N_3364,N_2894,N_2821);
nand U3365 (N_3365,N_2983,N_2852);
or U3366 (N_3366,N_2929,N_2791);
nand U3367 (N_3367,N_2717,N_2961);
nand U3368 (N_3368,N_2732,N_2520);
nor U3369 (N_3369,N_2842,N_2534);
and U3370 (N_3370,N_2866,N_2985);
xor U3371 (N_3371,N_2768,N_2531);
nor U3372 (N_3372,N_2687,N_2774);
nor U3373 (N_3373,N_2684,N_2704);
nor U3374 (N_3374,N_2759,N_2920);
or U3375 (N_3375,N_2514,N_2570);
and U3376 (N_3376,N_2661,N_2845);
and U3377 (N_3377,N_2705,N_2663);
nor U3378 (N_3378,N_2560,N_2738);
nand U3379 (N_3379,N_2745,N_2722);
or U3380 (N_3380,N_2649,N_2768);
or U3381 (N_3381,N_2505,N_2575);
nand U3382 (N_3382,N_2609,N_2592);
nand U3383 (N_3383,N_2972,N_2835);
or U3384 (N_3384,N_2949,N_2999);
nor U3385 (N_3385,N_2695,N_2832);
xnor U3386 (N_3386,N_2641,N_2996);
nand U3387 (N_3387,N_2609,N_2842);
and U3388 (N_3388,N_2654,N_2740);
nor U3389 (N_3389,N_2541,N_2753);
xnor U3390 (N_3390,N_2732,N_2872);
nand U3391 (N_3391,N_2876,N_2760);
or U3392 (N_3392,N_2676,N_2673);
or U3393 (N_3393,N_2704,N_2943);
nand U3394 (N_3394,N_2573,N_2596);
and U3395 (N_3395,N_2904,N_2615);
or U3396 (N_3396,N_2986,N_2934);
or U3397 (N_3397,N_2932,N_2863);
nor U3398 (N_3398,N_2592,N_2588);
and U3399 (N_3399,N_2992,N_2704);
or U3400 (N_3400,N_2880,N_2994);
xor U3401 (N_3401,N_2972,N_2725);
and U3402 (N_3402,N_2632,N_2939);
xor U3403 (N_3403,N_2999,N_2692);
xor U3404 (N_3404,N_2837,N_2680);
nor U3405 (N_3405,N_2908,N_2680);
and U3406 (N_3406,N_2898,N_2999);
nor U3407 (N_3407,N_2886,N_2930);
or U3408 (N_3408,N_2811,N_2852);
and U3409 (N_3409,N_2876,N_2971);
xnor U3410 (N_3410,N_2998,N_2913);
and U3411 (N_3411,N_2951,N_2524);
and U3412 (N_3412,N_2735,N_2566);
nand U3413 (N_3413,N_2754,N_2923);
xnor U3414 (N_3414,N_2846,N_2513);
xor U3415 (N_3415,N_2556,N_2690);
and U3416 (N_3416,N_2888,N_2645);
nand U3417 (N_3417,N_2908,N_2799);
nand U3418 (N_3418,N_2563,N_2873);
or U3419 (N_3419,N_2764,N_2570);
nand U3420 (N_3420,N_2631,N_2587);
nor U3421 (N_3421,N_2947,N_2542);
nor U3422 (N_3422,N_2819,N_2740);
xnor U3423 (N_3423,N_2915,N_2873);
or U3424 (N_3424,N_2723,N_2893);
xor U3425 (N_3425,N_2845,N_2737);
or U3426 (N_3426,N_2746,N_2886);
or U3427 (N_3427,N_2980,N_2764);
and U3428 (N_3428,N_2848,N_2737);
or U3429 (N_3429,N_2854,N_2864);
or U3430 (N_3430,N_2853,N_2686);
nor U3431 (N_3431,N_2624,N_2886);
nand U3432 (N_3432,N_2965,N_2806);
xnor U3433 (N_3433,N_2512,N_2786);
or U3434 (N_3434,N_2815,N_2712);
nor U3435 (N_3435,N_2862,N_2993);
or U3436 (N_3436,N_2642,N_2741);
or U3437 (N_3437,N_2593,N_2945);
and U3438 (N_3438,N_2848,N_2976);
and U3439 (N_3439,N_2917,N_2981);
or U3440 (N_3440,N_2935,N_2998);
nor U3441 (N_3441,N_2713,N_2507);
and U3442 (N_3442,N_2713,N_2926);
or U3443 (N_3443,N_2597,N_2669);
xor U3444 (N_3444,N_2720,N_2699);
and U3445 (N_3445,N_2832,N_2831);
nand U3446 (N_3446,N_2996,N_2635);
and U3447 (N_3447,N_2553,N_2875);
nand U3448 (N_3448,N_2663,N_2590);
nor U3449 (N_3449,N_2732,N_2798);
and U3450 (N_3450,N_2982,N_2583);
nor U3451 (N_3451,N_2534,N_2796);
xnor U3452 (N_3452,N_2798,N_2999);
xor U3453 (N_3453,N_2835,N_2935);
nor U3454 (N_3454,N_2943,N_2746);
or U3455 (N_3455,N_2523,N_2725);
or U3456 (N_3456,N_2669,N_2647);
and U3457 (N_3457,N_2886,N_2773);
nand U3458 (N_3458,N_2784,N_2774);
or U3459 (N_3459,N_2674,N_2811);
nand U3460 (N_3460,N_2631,N_2532);
nand U3461 (N_3461,N_2671,N_2559);
nand U3462 (N_3462,N_2950,N_2890);
nand U3463 (N_3463,N_2889,N_2814);
nand U3464 (N_3464,N_2739,N_2644);
nor U3465 (N_3465,N_2781,N_2842);
or U3466 (N_3466,N_2962,N_2966);
and U3467 (N_3467,N_2826,N_2983);
nand U3468 (N_3468,N_2917,N_2836);
nor U3469 (N_3469,N_2788,N_2982);
or U3470 (N_3470,N_2682,N_2737);
xor U3471 (N_3471,N_2699,N_2895);
and U3472 (N_3472,N_2751,N_2644);
nand U3473 (N_3473,N_2590,N_2769);
and U3474 (N_3474,N_2550,N_2642);
xnor U3475 (N_3475,N_2554,N_2951);
nand U3476 (N_3476,N_2659,N_2664);
nand U3477 (N_3477,N_2989,N_2884);
xnor U3478 (N_3478,N_2601,N_2577);
nor U3479 (N_3479,N_2856,N_2889);
and U3480 (N_3480,N_2649,N_2770);
and U3481 (N_3481,N_2889,N_2604);
or U3482 (N_3482,N_2556,N_2705);
xor U3483 (N_3483,N_2503,N_2815);
or U3484 (N_3484,N_2570,N_2609);
xor U3485 (N_3485,N_2779,N_2781);
and U3486 (N_3486,N_2730,N_2682);
nor U3487 (N_3487,N_2522,N_2984);
nand U3488 (N_3488,N_2951,N_2918);
nor U3489 (N_3489,N_2672,N_2902);
or U3490 (N_3490,N_2873,N_2731);
nor U3491 (N_3491,N_2742,N_2883);
or U3492 (N_3492,N_2826,N_2972);
nor U3493 (N_3493,N_2681,N_2753);
xor U3494 (N_3494,N_2894,N_2811);
or U3495 (N_3495,N_2940,N_2965);
or U3496 (N_3496,N_2505,N_2957);
nor U3497 (N_3497,N_2726,N_2513);
or U3498 (N_3498,N_2970,N_2710);
and U3499 (N_3499,N_2998,N_2595);
and U3500 (N_3500,N_3297,N_3094);
nor U3501 (N_3501,N_3149,N_3144);
xnor U3502 (N_3502,N_3290,N_3197);
xor U3503 (N_3503,N_3346,N_3456);
nor U3504 (N_3504,N_3276,N_3181);
or U3505 (N_3505,N_3172,N_3258);
nor U3506 (N_3506,N_3018,N_3118);
nand U3507 (N_3507,N_3283,N_3206);
nand U3508 (N_3508,N_3400,N_3281);
nand U3509 (N_3509,N_3405,N_3413);
nor U3510 (N_3510,N_3124,N_3292);
and U3511 (N_3511,N_3109,N_3257);
nor U3512 (N_3512,N_3389,N_3240);
nand U3513 (N_3513,N_3006,N_3313);
nand U3514 (N_3514,N_3351,N_3468);
or U3515 (N_3515,N_3287,N_3340);
nand U3516 (N_3516,N_3132,N_3021);
xnor U3517 (N_3517,N_3142,N_3384);
nand U3518 (N_3518,N_3294,N_3249);
nor U3519 (N_3519,N_3383,N_3376);
xnor U3520 (N_3520,N_3353,N_3199);
nand U3521 (N_3521,N_3422,N_3250);
xor U3522 (N_3522,N_3487,N_3026);
or U3523 (N_3523,N_3285,N_3083);
nand U3524 (N_3524,N_3230,N_3242);
nand U3525 (N_3525,N_3147,N_3348);
and U3526 (N_3526,N_3179,N_3238);
and U3527 (N_3527,N_3459,N_3282);
nor U3528 (N_3528,N_3491,N_3160);
or U3529 (N_3529,N_3274,N_3330);
nor U3530 (N_3530,N_3091,N_3084);
or U3531 (N_3531,N_3466,N_3039);
or U3532 (N_3532,N_3379,N_3477);
nor U3533 (N_3533,N_3038,N_3210);
or U3534 (N_3534,N_3056,N_3497);
xnor U3535 (N_3535,N_3471,N_3047);
nor U3536 (N_3536,N_3212,N_3417);
and U3537 (N_3537,N_3303,N_3222);
nor U3538 (N_3538,N_3234,N_3001);
nor U3539 (N_3539,N_3127,N_3409);
and U3540 (N_3540,N_3079,N_3218);
or U3541 (N_3541,N_3332,N_3223);
nor U3542 (N_3542,N_3399,N_3309);
nand U3543 (N_3543,N_3097,N_3366);
xnor U3544 (N_3544,N_3463,N_3163);
xor U3545 (N_3545,N_3397,N_3043);
and U3546 (N_3546,N_3485,N_3291);
xnor U3547 (N_3547,N_3102,N_3215);
or U3548 (N_3548,N_3357,N_3196);
nand U3549 (N_3549,N_3152,N_3385);
xor U3550 (N_3550,N_3436,N_3076);
nor U3551 (N_3551,N_3324,N_3099);
nand U3552 (N_3552,N_3065,N_3229);
nand U3553 (N_3553,N_3263,N_3003);
xor U3554 (N_3554,N_3123,N_3361);
xor U3555 (N_3555,N_3239,N_3489);
nand U3556 (N_3556,N_3386,N_3387);
nand U3557 (N_3557,N_3327,N_3075);
or U3558 (N_3558,N_3322,N_3002);
and U3559 (N_3559,N_3072,N_3219);
nand U3560 (N_3560,N_3209,N_3474);
nor U3561 (N_3561,N_3382,N_3183);
nor U3562 (N_3562,N_3341,N_3030);
nor U3563 (N_3563,N_3445,N_3236);
xnor U3564 (N_3564,N_3289,N_3381);
and U3565 (N_3565,N_3112,N_3494);
xnor U3566 (N_3566,N_3138,N_3165);
xor U3567 (N_3567,N_3055,N_3298);
and U3568 (N_3568,N_3469,N_3100);
or U3569 (N_3569,N_3279,N_3161);
nand U3570 (N_3570,N_3216,N_3339);
xor U3571 (N_3571,N_3137,N_3231);
nand U3572 (N_3572,N_3117,N_3246);
xnor U3573 (N_3573,N_3412,N_3203);
nor U3574 (N_3574,N_3490,N_3476);
xor U3575 (N_3575,N_3461,N_3156);
nor U3576 (N_3576,N_3153,N_3048);
or U3577 (N_3577,N_3051,N_3358);
and U3578 (N_3578,N_3221,N_3273);
nand U3579 (N_3579,N_3150,N_3325);
and U3580 (N_3580,N_3260,N_3368);
and U3581 (N_3581,N_3078,N_3244);
nand U3582 (N_3582,N_3068,N_3275);
nor U3583 (N_3583,N_3052,N_3040);
nor U3584 (N_3584,N_3464,N_3121);
or U3585 (N_3585,N_3071,N_3107);
xor U3586 (N_3586,N_3031,N_3146);
nor U3587 (N_3587,N_3269,N_3408);
xnor U3588 (N_3588,N_3119,N_3430);
and U3589 (N_3589,N_3355,N_3129);
nand U3590 (N_3590,N_3256,N_3151);
or U3591 (N_3591,N_3088,N_3085);
xor U3592 (N_3592,N_3278,N_3010);
nand U3593 (N_3593,N_3311,N_3407);
or U3594 (N_3594,N_3370,N_3074);
or U3595 (N_3595,N_3145,N_3095);
xnor U3596 (N_3596,N_3435,N_3182);
and U3597 (N_3597,N_3460,N_3217);
xnor U3598 (N_3598,N_3415,N_3000);
nand U3599 (N_3599,N_3470,N_3280);
nand U3600 (N_3600,N_3185,N_3125);
and U3601 (N_3601,N_3041,N_3053);
and U3602 (N_3602,N_3304,N_3406);
and U3603 (N_3603,N_3131,N_3180);
xnor U3604 (N_3604,N_3103,N_3493);
or U3605 (N_3605,N_3070,N_3403);
xnor U3606 (N_3606,N_3479,N_3308);
nor U3607 (N_3607,N_3194,N_3224);
nor U3608 (N_3608,N_3302,N_3089);
or U3609 (N_3609,N_3427,N_3005);
nand U3610 (N_3610,N_3315,N_3426);
nand U3611 (N_3611,N_3321,N_3081);
xor U3612 (N_3612,N_3451,N_3062);
nand U3613 (N_3613,N_3492,N_3367);
nand U3614 (N_3614,N_3438,N_3371);
nand U3615 (N_3615,N_3202,N_3017);
nand U3616 (N_3616,N_3188,N_3027);
and U3617 (N_3617,N_3044,N_3042);
nand U3618 (N_3618,N_3227,N_3440);
xor U3619 (N_3619,N_3004,N_3305);
xor U3620 (N_3620,N_3499,N_3296);
nor U3621 (N_3621,N_3465,N_3418);
or U3622 (N_3622,N_3190,N_3432);
xnor U3623 (N_3623,N_3186,N_3326);
or U3624 (N_3624,N_3488,N_3170);
nor U3625 (N_3625,N_3082,N_3114);
xor U3626 (N_3626,N_3356,N_3211);
xnor U3627 (N_3627,N_3111,N_3226);
nor U3628 (N_3628,N_3193,N_3155);
xor U3629 (N_3629,N_3016,N_3478);
nor U3630 (N_3630,N_3106,N_3028);
nand U3631 (N_3631,N_3232,N_3446);
xor U3632 (N_3632,N_3066,N_3423);
or U3633 (N_3633,N_3347,N_3344);
and U3634 (N_3634,N_3345,N_3058);
or U3635 (N_3635,N_3104,N_3191);
nand U3636 (N_3636,N_3034,N_3306);
nor U3637 (N_3637,N_3364,N_3388);
or U3638 (N_3638,N_3241,N_3266);
nand U3639 (N_3639,N_3243,N_3204);
and U3640 (N_3640,N_3277,N_3495);
xor U3641 (N_3641,N_3157,N_3380);
and U3642 (N_3642,N_3073,N_3301);
or U3643 (N_3643,N_3372,N_3428);
and U3644 (N_3644,N_3205,N_3447);
or U3645 (N_3645,N_3271,N_3267);
nand U3646 (N_3646,N_3067,N_3126);
nand U3647 (N_3647,N_3090,N_3248);
nand U3648 (N_3648,N_3333,N_3171);
or U3649 (N_3649,N_3268,N_3255);
xnor U3650 (N_3650,N_3293,N_3481);
nor U3651 (N_3651,N_3411,N_3086);
and U3652 (N_3652,N_3317,N_3424);
and U3653 (N_3653,N_3022,N_3024);
or U3654 (N_3654,N_3475,N_3013);
or U3655 (N_3655,N_3046,N_3375);
xor U3656 (N_3656,N_3128,N_3093);
and U3657 (N_3657,N_3176,N_3113);
nand U3658 (N_3658,N_3425,N_3329);
nand U3659 (N_3659,N_3164,N_3014);
nor U3660 (N_3660,N_3484,N_3323);
or U3661 (N_3661,N_3458,N_3262);
or U3662 (N_3662,N_3167,N_3015);
xnor U3663 (N_3663,N_3077,N_3120);
xnor U3664 (N_3664,N_3310,N_3336);
xnor U3665 (N_3665,N_3143,N_3110);
or U3666 (N_3666,N_3396,N_3228);
and U3667 (N_3667,N_3416,N_3162);
or U3668 (N_3668,N_3159,N_3420);
xor U3669 (N_3669,N_3300,N_3390);
or U3670 (N_3670,N_3166,N_3139);
and U3671 (N_3671,N_3272,N_3480);
xor U3672 (N_3672,N_3020,N_3254);
or U3673 (N_3673,N_3168,N_3235);
and U3674 (N_3674,N_3319,N_3178);
xor U3675 (N_3675,N_3135,N_3314);
or U3676 (N_3676,N_3369,N_3233);
and U3677 (N_3677,N_3195,N_3421);
nor U3678 (N_3678,N_3473,N_3395);
and U3679 (N_3679,N_3442,N_3472);
or U3680 (N_3680,N_3251,N_3105);
xnor U3681 (N_3681,N_3115,N_3116);
and U3682 (N_3682,N_3335,N_3069);
or U3683 (N_3683,N_3410,N_3350);
and U3684 (N_3684,N_3498,N_3286);
nor U3685 (N_3685,N_3063,N_3270);
and U3686 (N_3686,N_3404,N_3433);
nand U3687 (N_3687,N_3033,N_3101);
nand U3688 (N_3688,N_3441,N_3174);
and U3689 (N_3689,N_3439,N_3208);
or U3690 (N_3690,N_3331,N_3377);
xnor U3691 (N_3691,N_3252,N_3253);
nand U3692 (N_3692,N_3050,N_3337);
nand U3693 (N_3693,N_3402,N_3080);
xnor U3694 (N_3694,N_3496,N_3177);
nor U3695 (N_3695,N_3237,N_3312);
nor U3696 (N_3696,N_3141,N_3374);
xor U3697 (N_3697,N_3225,N_3295);
and U3698 (N_3698,N_3198,N_3365);
and U3699 (N_3699,N_3060,N_3247);
nor U3700 (N_3700,N_3354,N_3391);
and U3701 (N_3701,N_3437,N_3352);
xnor U3702 (N_3702,N_3061,N_3011);
or U3703 (N_3703,N_3134,N_3483);
xor U3704 (N_3704,N_3201,N_3299);
nor U3705 (N_3705,N_3029,N_3450);
nor U3706 (N_3706,N_3467,N_3455);
or U3707 (N_3707,N_3007,N_3059);
and U3708 (N_3708,N_3214,N_3360);
and U3709 (N_3709,N_3154,N_3245);
nor U3710 (N_3710,N_3023,N_3343);
and U3711 (N_3711,N_3362,N_3133);
or U3712 (N_3712,N_3032,N_3261);
and U3713 (N_3713,N_3429,N_3025);
nor U3714 (N_3714,N_3444,N_3359);
or U3715 (N_3715,N_3187,N_3035);
and U3716 (N_3716,N_3045,N_3414);
and U3717 (N_3717,N_3108,N_3307);
nor U3718 (N_3718,N_3009,N_3288);
xnor U3719 (N_3719,N_3200,N_3284);
nor U3720 (N_3720,N_3264,N_3169);
and U3721 (N_3721,N_3378,N_3318);
or U3722 (N_3722,N_3316,N_3452);
nand U3723 (N_3723,N_3008,N_3342);
nand U3724 (N_3724,N_3136,N_3462);
xor U3725 (N_3725,N_3393,N_3148);
and U3726 (N_3726,N_3012,N_3401);
and U3727 (N_3727,N_3448,N_3443);
nand U3728 (N_3728,N_3486,N_3173);
xnor U3729 (N_3729,N_3098,N_3431);
nand U3730 (N_3730,N_3158,N_3482);
xor U3731 (N_3731,N_3087,N_3140);
or U3732 (N_3732,N_3175,N_3363);
nand U3733 (N_3733,N_3394,N_3184);
nor U3734 (N_3734,N_3054,N_3434);
and U3735 (N_3735,N_3037,N_3064);
and U3736 (N_3736,N_3419,N_3122);
xnor U3737 (N_3737,N_3259,N_3265);
nand U3738 (N_3738,N_3192,N_3398);
nor U3739 (N_3739,N_3328,N_3213);
or U3740 (N_3740,N_3189,N_3454);
nor U3741 (N_3741,N_3220,N_3130);
and U3742 (N_3742,N_3349,N_3092);
xnor U3743 (N_3743,N_3334,N_3019);
nand U3744 (N_3744,N_3049,N_3457);
or U3745 (N_3745,N_3373,N_3320);
nor U3746 (N_3746,N_3096,N_3057);
nand U3747 (N_3747,N_3036,N_3207);
nand U3748 (N_3748,N_3449,N_3338);
xnor U3749 (N_3749,N_3392,N_3453);
nor U3750 (N_3750,N_3282,N_3093);
xnor U3751 (N_3751,N_3000,N_3417);
xor U3752 (N_3752,N_3119,N_3117);
nor U3753 (N_3753,N_3119,N_3299);
or U3754 (N_3754,N_3194,N_3474);
xnor U3755 (N_3755,N_3022,N_3103);
nand U3756 (N_3756,N_3415,N_3431);
xnor U3757 (N_3757,N_3493,N_3491);
nand U3758 (N_3758,N_3409,N_3195);
or U3759 (N_3759,N_3378,N_3026);
and U3760 (N_3760,N_3265,N_3099);
nand U3761 (N_3761,N_3151,N_3379);
xnor U3762 (N_3762,N_3002,N_3141);
nor U3763 (N_3763,N_3263,N_3050);
nor U3764 (N_3764,N_3187,N_3440);
nand U3765 (N_3765,N_3135,N_3172);
xor U3766 (N_3766,N_3120,N_3458);
and U3767 (N_3767,N_3088,N_3394);
xor U3768 (N_3768,N_3433,N_3168);
xor U3769 (N_3769,N_3330,N_3119);
nand U3770 (N_3770,N_3386,N_3372);
nand U3771 (N_3771,N_3399,N_3249);
nor U3772 (N_3772,N_3353,N_3383);
and U3773 (N_3773,N_3494,N_3080);
xnor U3774 (N_3774,N_3151,N_3259);
and U3775 (N_3775,N_3139,N_3205);
nand U3776 (N_3776,N_3443,N_3463);
and U3777 (N_3777,N_3294,N_3389);
nand U3778 (N_3778,N_3247,N_3221);
xnor U3779 (N_3779,N_3000,N_3172);
xnor U3780 (N_3780,N_3222,N_3338);
and U3781 (N_3781,N_3114,N_3199);
or U3782 (N_3782,N_3250,N_3203);
and U3783 (N_3783,N_3055,N_3284);
nor U3784 (N_3784,N_3379,N_3367);
nor U3785 (N_3785,N_3112,N_3096);
nor U3786 (N_3786,N_3016,N_3373);
xnor U3787 (N_3787,N_3469,N_3289);
nor U3788 (N_3788,N_3033,N_3434);
nor U3789 (N_3789,N_3492,N_3247);
and U3790 (N_3790,N_3448,N_3051);
nand U3791 (N_3791,N_3445,N_3046);
and U3792 (N_3792,N_3241,N_3142);
and U3793 (N_3793,N_3296,N_3253);
nand U3794 (N_3794,N_3118,N_3388);
xor U3795 (N_3795,N_3192,N_3476);
and U3796 (N_3796,N_3433,N_3386);
or U3797 (N_3797,N_3308,N_3493);
and U3798 (N_3798,N_3204,N_3432);
nand U3799 (N_3799,N_3345,N_3074);
xor U3800 (N_3800,N_3097,N_3029);
and U3801 (N_3801,N_3315,N_3073);
nor U3802 (N_3802,N_3102,N_3211);
or U3803 (N_3803,N_3021,N_3449);
and U3804 (N_3804,N_3329,N_3020);
xor U3805 (N_3805,N_3114,N_3360);
nor U3806 (N_3806,N_3375,N_3456);
or U3807 (N_3807,N_3408,N_3303);
and U3808 (N_3808,N_3134,N_3274);
and U3809 (N_3809,N_3127,N_3170);
and U3810 (N_3810,N_3133,N_3005);
or U3811 (N_3811,N_3201,N_3090);
xnor U3812 (N_3812,N_3280,N_3360);
and U3813 (N_3813,N_3121,N_3377);
xor U3814 (N_3814,N_3205,N_3437);
xnor U3815 (N_3815,N_3074,N_3478);
xor U3816 (N_3816,N_3097,N_3278);
nor U3817 (N_3817,N_3434,N_3364);
xnor U3818 (N_3818,N_3420,N_3148);
xor U3819 (N_3819,N_3388,N_3039);
or U3820 (N_3820,N_3367,N_3478);
xor U3821 (N_3821,N_3387,N_3411);
nand U3822 (N_3822,N_3465,N_3292);
or U3823 (N_3823,N_3234,N_3180);
or U3824 (N_3824,N_3463,N_3444);
nand U3825 (N_3825,N_3170,N_3159);
nor U3826 (N_3826,N_3224,N_3120);
and U3827 (N_3827,N_3080,N_3091);
nand U3828 (N_3828,N_3074,N_3242);
or U3829 (N_3829,N_3036,N_3473);
and U3830 (N_3830,N_3298,N_3144);
nand U3831 (N_3831,N_3304,N_3454);
xnor U3832 (N_3832,N_3077,N_3497);
nand U3833 (N_3833,N_3284,N_3480);
nor U3834 (N_3834,N_3138,N_3438);
xor U3835 (N_3835,N_3385,N_3394);
nor U3836 (N_3836,N_3008,N_3156);
nor U3837 (N_3837,N_3114,N_3331);
and U3838 (N_3838,N_3251,N_3481);
or U3839 (N_3839,N_3058,N_3243);
xnor U3840 (N_3840,N_3492,N_3263);
or U3841 (N_3841,N_3168,N_3228);
xnor U3842 (N_3842,N_3082,N_3426);
or U3843 (N_3843,N_3485,N_3304);
or U3844 (N_3844,N_3406,N_3385);
nand U3845 (N_3845,N_3168,N_3486);
nor U3846 (N_3846,N_3178,N_3218);
and U3847 (N_3847,N_3454,N_3050);
nand U3848 (N_3848,N_3293,N_3230);
nand U3849 (N_3849,N_3283,N_3064);
nand U3850 (N_3850,N_3047,N_3440);
and U3851 (N_3851,N_3178,N_3269);
or U3852 (N_3852,N_3301,N_3235);
xor U3853 (N_3853,N_3260,N_3353);
nand U3854 (N_3854,N_3001,N_3139);
and U3855 (N_3855,N_3137,N_3053);
xnor U3856 (N_3856,N_3282,N_3016);
nor U3857 (N_3857,N_3456,N_3093);
nor U3858 (N_3858,N_3095,N_3288);
nand U3859 (N_3859,N_3391,N_3385);
nand U3860 (N_3860,N_3435,N_3294);
nand U3861 (N_3861,N_3275,N_3433);
xor U3862 (N_3862,N_3297,N_3485);
and U3863 (N_3863,N_3192,N_3032);
and U3864 (N_3864,N_3376,N_3348);
and U3865 (N_3865,N_3000,N_3212);
nor U3866 (N_3866,N_3084,N_3305);
xnor U3867 (N_3867,N_3266,N_3038);
xnor U3868 (N_3868,N_3189,N_3420);
or U3869 (N_3869,N_3133,N_3248);
or U3870 (N_3870,N_3289,N_3052);
and U3871 (N_3871,N_3476,N_3215);
and U3872 (N_3872,N_3338,N_3121);
nand U3873 (N_3873,N_3385,N_3359);
and U3874 (N_3874,N_3203,N_3288);
xor U3875 (N_3875,N_3446,N_3488);
nor U3876 (N_3876,N_3225,N_3126);
or U3877 (N_3877,N_3475,N_3137);
nand U3878 (N_3878,N_3080,N_3104);
and U3879 (N_3879,N_3049,N_3153);
and U3880 (N_3880,N_3232,N_3489);
nor U3881 (N_3881,N_3075,N_3289);
and U3882 (N_3882,N_3245,N_3073);
and U3883 (N_3883,N_3389,N_3332);
and U3884 (N_3884,N_3063,N_3186);
nor U3885 (N_3885,N_3180,N_3418);
or U3886 (N_3886,N_3042,N_3176);
xor U3887 (N_3887,N_3364,N_3171);
nor U3888 (N_3888,N_3117,N_3302);
or U3889 (N_3889,N_3230,N_3430);
or U3890 (N_3890,N_3031,N_3279);
and U3891 (N_3891,N_3324,N_3290);
nor U3892 (N_3892,N_3309,N_3140);
or U3893 (N_3893,N_3022,N_3153);
nand U3894 (N_3894,N_3168,N_3033);
or U3895 (N_3895,N_3312,N_3382);
and U3896 (N_3896,N_3164,N_3336);
nor U3897 (N_3897,N_3335,N_3183);
or U3898 (N_3898,N_3463,N_3096);
and U3899 (N_3899,N_3209,N_3302);
and U3900 (N_3900,N_3017,N_3462);
or U3901 (N_3901,N_3400,N_3319);
xnor U3902 (N_3902,N_3005,N_3230);
or U3903 (N_3903,N_3331,N_3069);
nor U3904 (N_3904,N_3371,N_3383);
xor U3905 (N_3905,N_3029,N_3468);
or U3906 (N_3906,N_3476,N_3228);
nand U3907 (N_3907,N_3209,N_3058);
and U3908 (N_3908,N_3273,N_3452);
and U3909 (N_3909,N_3436,N_3169);
xor U3910 (N_3910,N_3013,N_3192);
nor U3911 (N_3911,N_3320,N_3131);
and U3912 (N_3912,N_3091,N_3436);
xor U3913 (N_3913,N_3003,N_3424);
nand U3914 (N_3914,N_3203,N_3106);
nand U3915 (N_3915,N_3052,N_3062);
or U3916 (N_3916,N_3148,N_3112);
or U3917 (N_3917,N_3390,N_3485);
and U3918 (N_3918,N_3178,N_3372);
nor U3919 (N_3919,N_3121,N_3409);
xnor U3920 (N_3920,N_3488,N_3216);
xnor U3921 (N_3921,N_3034,N_3291);
nand U3922 (N_3922,N_3082,N_3034);
xor U3923 (N_3923,N_3312,N_3219);
xor U3924 (N_3924,N_3077,N_3459);
or U3925 (N_3925,N_3385,N_3423);
nand U3926 (N_3926,N_3403,N_3158);
or U3927 (N_3927,N_3168,N_3443);
and U3928 (N_3928,N_3456,N_3453);
nor U3929 (N_3929,N_3324,N_3053);
nor U3930 (N_3930,N_3079,N_3413);
xor U3931 (N_3931,N_3222,N_3443);
nor U3932 (N_3932,N_3351,N_3187);
nor U3933 (N_3933,N_3292,N_3011);
xnor U3934 (N_3934,N_3401,N_3420);
and U3935 (N_3935,N_3120,N_3342);
nor U3936 (N_3936,N_3049,N_3354);
nor U3937 (N_3937,N_3058,N_3387);
nand U3938 (N_3938,N_3236,N_3390);
nor U3939 (N_3939,N_3192,N_3238);
xor U3940 (N_3940,N_3160,N_3248);
nand U3941 (N_3941,N_3419,N_3156);
nor U3942 (N_3942,N_3107,N_3230);
nor U3943 (N_3943,N_3153,N_3295);
xor U3944 (N_3944,N_3410,N_3397);
xnor U3945 (N_3945,N_3259,N_3264);
and U3946 (N_3946,N_3377,N_3242);
xnor U3947 (N_3947,N_3040,N_3180);
nor U3948 (N_3948,N_3459,N_3242);
xnor U3949 (N_3949,N_3374,N_3058);
or U3950 (N_3950,N_3452,N_3498);
and U3951 (N_3951,N_3074,N_3403);
nand U3952 (N_3952,N_3293,N_3266);
nor U3953 (N_3953,N_3234,N_3025);
xor U3954 (N_3954,N_3278,N_3290);
or U3955 (N_3955,N_3438,N_3338);
nand U3956 (N_3956,N_3487,N_3238);
nor U3957 (N_3957,N_3010,N_3456);
and U3958 (N_3958,N_3257,N_3004);
and U3959 (N_3959,N_3325,N_3388);
nand U3960 (N_3960,N_3458,N_3122);
or U3961 (N_3961,N_3089,N_3121);
xnor U3962 (N_3962,N_3323,N_3077);
xnor U3963 (N_3963,N_3249,N_3054);
xor U3964 (N_3964,N_3465,N_3486);
or U3965 (N_3965,N_3186,N_3497);
nand U3966 (N_3966,N_3121,N_3402);
nand U3967 (N_3967,N_3097,N_3310);
or U3968 (N_3968,N_3076,N_3284);
or U3969 (N_3969,N_3204,N_3172);
or U3970 (N_3970,N_3270,N_3264);
nand U3971 (N_3971,N_3176,N_3439);
and U3972 (N_3972,N_3244,N_3469);
nand U3973 (N_3973,N_3156,N_3307);
nand U3974 (N_3974,N_3167,N_3233);
or U3975 (N_3975,N_3470,N_3484);
xnor U3976 (N_3976,N_3242,N_3010);
or U3977 (N_3977,N_3415,N_3061);
nand U3978 (N_3978,N_3044,N_3271);
nor U3979 (N_3979,N_3163,N_3216);
nand U3980 (N_3980,N_3362,N_3092);
nand U3981 (N_3981,N_3472,N_3141);
and U3982 (N_3982,N_3246,N_3173);
xnor U3983 (N_3983,N_3165,N_3149);
nand U3984 (N_3984,N_3012,N_3245);
nor U3985 (N_3985,N_3288,N_3271);
xnor U3986 (N_3986,N_3098,N_3137);
and U3987 (N_3987,N_3440,N_3111);
or U3988 (N_3988,N_3336,N_3042);
xnor U3989 (N_3989,N_3331,N_3466);
xnor U3990 (N_3990,N_3331,N_3256);
and U3991 (N_3991,N_3430,N_3419);
nand U3992 (N_3992,N_3176,N_3237);
nand U3993 (N_3993,N_3375,N_3382);
and U3994 (N_3994,N_3105,N_3463);
nand U3995 (N_3995,N_3229,N_3116);
or U3996 (N_3996,N_3332,N_3221);
and U3997 (N_3997,N_3451,N_3493);
xor U3998 (N_3998,N_3391,N_3164);
xor U3999 (N_3999,N_3255,N_3460);
xor U4000 (N_4000,N_3990,N_3894);
or U4001 (N_4001,N_3573,N_3719);
or U4002 (N_4002,N_3622,N_3675);
or U4003 (N_4003,N_3604,N_3500);
nand U4004 (N_4004,N_3686,N_3738);
nor U4005 (N_4005,N_3948,N_3515);
nor U4006 (N_4006,N_3981,N_3683);
and U4007 (N_4007,N_3633,N_3890);
and U4008 (N_4008,N_3816,N_3749);
nor U4009 (N_4009,N_3586,N_3858);
or U4010 (N_4010,N_3626,N_3659);
and U4011 (N_4011,N_3510,N_3840);
nor U4012 (N_4012,N_3587,N_3759);
and U4013 (N_4013,N_3778,N_3875);
nor U4014 (N_4014,N_3791,N_3537);
or U4015 (N_4015,N_3852,N_3671);
or U4016 (N_4016,N_3975,N_3694);
nor U4017 (N_4017,N_3962,N_3946);
and U4018 (N_4018,N_3502,N_3649);
xor U4019 (N_4019,N_3889,N_3953);
or U4020 (N_4020,N_3985,N_3531);
nor U4021 (N_4021,N_3583,N_3901);
or U4022 (N_4022,N_3549,N_3927);
or U4023 (N_4023,N_3780,N_3730);
nor U4024 (N_4024,N_3781,N_3577);
nand U4025 (N_4025,N_3906,N_3922);
xor U4026 (N_4026,N_3844,N_3608);
and U4027 (N_4027,N_3525,N_3923);
xor U4028 (N_4028,N_3596,N_3945);
xnor U4029 (N_4029,N_3704,N_3881);
xnor U4030 (N_4030,N_3826,N_3580);
nor U4031 (N_4031,N_3550,N_3527);
nand U4032 (N_4032,N_3718,N_3555);
and U4033 (N_4033,N_3909,N_3862);
and U4034 (N_4034,N_3755,N_3884);
nand U4035 (N_4035,N_3857,N_3585);
nor U4036 (N_4036,N_3829,N_3554);
xor U4037 (N_4037,N_3993,N_3963);
xor U4038 (N_4038,N_3831,N_3853);
or U4039 (N_4039,N_3669,N_3711);
xnor U4040 (N_4040,N_3842,N_3956);
and U4041 (N_4041,N_3631,N_3815);
xnor U4042 (N_4042,N_3636,N_3790);
nand U4043 (N_4043,N_3805,N_3677);
and U4044 (N_4044,N_3760,N_3989);
nor U4045 (N_4045,N_3642,N_3972);
nand U4046 (N_4046,N_3827,N_3637);
and U4047 (N_4047,N_3582,N_3943);
nor U4048 (N_4048,N_3575,N_3775);
and U4049 (N_4049,N_3655,N_3559);
nand U4050 (N_4050,N_3746,N_3941);
xor U4051 (N_4051,N_3887,N_3632);
and U4052 (N_4052,N_3625,N_3744);
nand U4053 (N_4053,N_3662,N_3933);
nor U4054 (N_4054,N_3503,N_3732);
nor U4055 (N_4055,N_3828,N_3822);
nand U4056 (N_4056,N_3532,N_3770);
or U4057 (N_4057,N_3505,N_3609);
xnor U4058 (N_4058,N_3891,N_3942);
or U4059 (N_4059,N_3650,N_3562);
or U4060 (N_4060,N_3995,N_3673);
and U4061 (N_4061,N_3788,N_3839);
or U4062 (N_4062,N_3886,N_3638);
xor U4063 (N_4063,N_3877,N_3727);
nand U4064 (N_4064,N_3809,N_3773);
nor U4065 (N_4065,N_3740,N_3581);
nand U4066 (N_4066,N_3810,N_3610);
nor U4067 (N_4067,N_3911,N_3836);
and U4068 (N_4068,N_3986,N_3764);
nand U4069 (N_4069,N_3529,N_3691);
and U4070 (N_4070,N_3794,N_3926);
nand U4071 (N_4071,N_3651,N_3670);
or U4072 (N_4072,N_3695,N_3974);
nor U4073 (N_4073,N_3623,N_3590);
nand U4074 (N_4074,N_3854,N_3660);
and U4075 (N_4075,N_3874,N_3615);
nor U4076 (N_4076,N_3932,N_3705);
nand U4077 (N_4077,N_3793,N_3903);
nor U4078 (N_4078,N_3980,N_3769);
and U4079 (N_4079,N_3777,N_3726);
nand U4080 (N_4080,N_3750,N_3992);
nand U4081 (N_4081,N_3845,N_3850);
nand U4082 (N_4082,N_3849,N_3728);
nor U4083 (N_4083,N_3865,N_3762);
nand U4084 (N_4084,N_3818,N_3507);
nor U4085 (N_4085,N_3968,N_3912);
or U4086 (N_4086,N_3936,N_3612);
xnor U4087 (N_4087,N_3924,N_3944);
nor U4088 (N_4088,N_3663,N_3667);
and U4089 (N_4089,N_3544,N_3693);
or U4090 (N_4090,N_3518,N_3784);
and U4091 (N_4091,N_3878,N_3761);
xor U4092 (N_4092,N_3925,N_3699);
nor U4093 (N_4093,N_3592,N_3506);
or U4094 (N_4094,N_3534,N_3966);
and U4095 (N_4095,N_3617,N_3666);
or U4096 (N_4096,N_3949,N_3645);
nand U4097 (N_4097,N_3978,N_3568);
xnor U4098 (N_4098,N_3606,N_3861);
and U4099 (N_4099,N_3598,N_3792);
nor U4100 (N_4100,N_3516,N_3756);
or U4101 (N_4101,N_3997,N_3888);
nand U4102 (N_4102,N_3658,N_3751);
xor U4103 (N_4103,N_3823,N_3939);
nor U4104 (N_4104,N_3897,N_3834);
nor U4105 (N_4105,N_3648,N_3754);
or U4106 (N_4106,N_3843,N_3758);
nand U4107 (N_4107,N_3713,N_3514);
nand U4108 (N_4108,N_3921,N_3747);
nor U4109 (N_4109,N_3964,N_3847);
or U4110 (N_4110,N_3982,N_3766);
nor U4111 (N_4111,N_3902,N_3799);
nor U4112 (N_4112,N_3628,N_3552);
and U4113 (N_4113,N_3541,N_3951);
and U4114 (N_4114,N_3976,N_3715);
nand U4115 (N_4115,N_3971,N_3538);
or U4116 (N_4116,N_3918,N_3873);
nand U4117 (N_4117,N_3915,N_3787);
or U4118 (N_4118,N_3661,N_3629);
and U4119 (N_4119,N_3814,N_3914);
nor U4120 (N_4120,N_3748,N_3872);
or U4121 (N_4121,N_3556,N_3624);
xnor U4122 (N_4122,N_3947,N_3812);
and U4123 (N_4123,N_3690,N_3868);
or U4124 (N_4124,N_3863,N_3900);
xnor U4125 (N_4125,N_3571,N_3833);
and U4126 (N_4126,N_3572,N_3892);
xnor U4127 (N_4127,N_3907,N_3696);
xnor U4128 (N_4128,N_3689,N_3917);
xor U4129 (N_4129,N_3804,N_3593);
nor U4130 (N_4130,N_3916,N_3692);
nand U4131 (N_4131,N_3621,N_3929);
nor U4132 (N_4132,N_3513,N_3681);
nor U4133 (N_4133,N_3680,N_3603);
nand U4134 (N_4134,N_3664,N_3611);
nand U4135 (N_4135,N_3595,N_3722);
and U4136 (N_4136,N_3540,N_3825);
or U4137 (N_4137,N_3551,N_3896);
xor U4138 (N_4138,N_3731,N_3652);
and U4139 (N_4139,N_3521,N_3653);
or U4140 (N_4140,N_3709,N_3563);
or U4141 (N_4141,N_3801,N_3937);
or U4142 (N_4142,N_3984,N_3768);
xor U4143 (N_4143,N_3783,N_3883);
nor U4144 (N_4144,N_3739,N_3565);
or U4145 (N_4145,N_3765,N_3536);
or U4146 (N_4146,N_3898,N_3796);
nor U4147 (N_4147,N_3807,N_3987);
nand U4148 (N_4148,N_3772,N_3589);
nor U4149 (N_4149,N_3576,N_3588);
and U4150 (N_4150,N_3800,N_3880);
xor U4151 (N_4151,N_3720,N_3957);
or U4152 (N_4152,N_3910,N_3511);
and U4153 (N_4153,N_3996,N_3767);
nand U4154 (N_4154,N_3547,N_3570);
xor U4155 (N_4155,N_3859,N_3871);
xor U4156 (N_4156,N_3928,N_3950);
and U4157 (N_4157,N_3607,N_3931);
nand U4158 (N_4158,N_3753,N_3717);
nor U4159 (N_4159,N_3601,N_3647);
nand U4160 (N_4160,N_3991,N_3835);
or U4161 (N_4161,N_3630,N_3786);
nor U4162 (N_4162,N_3806,N_3895);
or U4163 (N_4163,N_3714,N_3602);
or U4164 (N_4164,N_3665,N_3882);
nand U4165 (N_4165,N_3560,N_3566);
xnor U4166 (N_4166,N_3960,N_3935);
or U4167 (N_4167,N_3741,N_3501);
or U4168 (N_4168,N_3522,N_3934);
xnor U4169 (N_4169,N_3742,N_3820);
nand U4170 (N_4170,N_3860,N_3548);
or U4171 (N_4171,N_3657,N_3724);
nor U4172 (N_4172,N_3605,N_3774);
and U4173 (N_4173,N_3701,N_3591);
and U4174 (N_4174,N_3994,N_3672);
xnor U4175 (N_4175,N_3830,N_3908);
nand U4176 (N_4176,N_3838,N_3509);
nand U4177 (N_4177,N_3557,N_3938);
and U4178 (N_4178,N_3876,N_3656);
xnor U4179 (N_4179,N_3599,N_3771);
or U4180 (N_4180,N_3619,N_3685);
nand U4181 (N_4181,N_3795,N_3940);
nor U4182 (N_4182,N_3885,N_3855);
or U4183 (N_4183,N_3779,N_3893);
nand U4184 (N_4184,N_3697,N_3654);
or U4185 (N_4185,N_3594,N_3763);
nor U4186 (N_4186,N_3620,N_3545);
xor U4187 (N_4187,N_3702,N_3600);
nand U4188 (N_4188,N_3999,N_3808);
or U4189 (N_4189,N_3710,N_3729);
and U4190 (N_4190,N_3578,N_3584);
or U4191 (N_4191,N_3523,N_3959);
or U4192 (N_4192,N_3954,N_3821);
xor U4193 (N_4193,N_3803,N_3819);
nor U4194 (N_4194,N_3967,N_3564);
nand U4195 (N_4195,N_3837,N_3782);
and U4196 (N_4196,N_3958,N_3614);
nor U4197 (N_4197,N_3635,N_3952);
nor U4198 (N_4198,N_3634,N_3866);
and U4199 (N_4199,N_3721,N_3678);
and U4200 (N_4200,N_3752,N_3688);
xor U4201 (N_4201,N_3668,N_3970);
xor U4202 (N_4202,N_3832,N_3641);
nand U4203 (N_4203,N_3703,N_3618);
or U4204 (N_4204,N_3524,N_3687);
or U4205 (N_4205,N_3539,N_3646);
or U4206 (N_4206,N_3579,N_3736);
nor U4207 (N_4207,N_3869,N_3899);
and U4208 (N_4208,N_3597,N_3789);
and U4209 (N_4209,N_3569,N_3969);
nand U4210 (N_4210,N_3674,N_3535);
and U4211 (N_4211,N_3616,N_3508);
nor U4212 (N_4212,N_3698,N_3627);
and U4213 (N_4213,N_3679,N_3920);
xor U4214 (N_4214,N_3824,N_3639);
nand U4215 (N_4215,N_3870,N_3977);
nor U4216 (N_4216,N_3706,N_3841);
nand U4217 (N_4217,N_3512,N_3640);
or U4218 (N_4218,N_3879,N_3817);
nand U4219 (N_4219,N_3567,N_3864);
nor U4220 (N_4220,N_3965,N_3743);
xor U4221 (N_4221,N_3961,N_3735);
nor U4222 (N_4222,N_3785,N_3676);
xnor U4223 (N_4223,N_3930,N_3848);
xnor U4224 (N_4224,N_3574,N_3988);
xor U4225 (N_4225,N_3561,N_3707);
nor U4226 (N_4226,N_3867,N_3643);
or U4227 (N_4227,N_3723,N_3983);
nand U4228 (N_4228,N_3973,N_3776);
or U4229 (N_4229,N_3558,N_3716);
xor U4230 (N_4230,N_3682,N_3734);
or U4231 (N_4231,N_3811,N_3613);
xnor U4232 (N_4232,N_3533,N_3644);
or U4233 (N_4233,N_3955,N_3851);
nand U4234 (N_4234,N_3998,N_3797);
and U4235 (N_4235,N_3737,N_3712);
nor U4236 (N_4236,N_3979,N_3543);
nand U4237 (N_4237,N_3745,N_3700);
or U4238 (N_4238,N_3684,N_3725);
nor U4239 (N_4239,N_3733,N_3846);
nor U4240 (N_4240,N_3905,N_3520);
and U4241 (N_4241,N_3526,N_3798);
nor U4242 (N_4242,N_3528,N_3519);
or U4243 (N_4243,N_3856,N_3504);
nor U4244 (N_4244,N_3757,N_3904);
and U4245 (N_4245,N_3708,N_3542);
and U4246 (N_4246,N_3546,N_3802);
nor U4247 (N_4247,N_3919,N_3913);
nand U4248 (N_4248,N_3813,N_3553);
or U4249 (N_4249,N_3530,N_3517);
and U4250 (N_4250,N_3636,N_3611);
nor U4251 (N_4251,N_3678,N_3758);
and U4252 (N_4252,N_3611,N_3717);
and U4253 (N_4253,N_3833,N_3570);
nand U4254 (N_4254,N_3893,N_3898);
nor U4255 (N_4255,N_3726,N_3677);
nand U4256 (N_4256,N_3809,N_3904);
xnor U4257 (N_4257,N_3916,N_3672);
nor U4258 (N_4258,N_3712,N_3864);
nor U4259 (N_4259,N_3744,N_3903);
nor U4260 (N_4260,N_3744,N_3885);
xor U4261 (N_4261,N_3903,N_3622);
nor U4262 (N_4262,N_3696,N_3753);
nand U4263 (N_4263,N_3652,N_3633);
nor U4264 (N_4264,N_3573,N_3967);
and U4265 (N_4265,N_3581,N_3803);
or U4266 (N_4266,N_3713,N_3742);
nor U4267 (N_4267,N_3759,N_3588);
and U4268 (N_4268,N_3970,N_3809);
nand U4269 (N_4269,N_3591,N_3940);
and U4270 (N_4270,N_3609,N_3755);
and U4271 (N_4271,N_3759,N_3650);
xor U4272 (N_4272,N_3731,N_3813);
xor U4273 (N_4273,N_3986,N_3973);
nor U4274 (N_4274,N_3802,N_3746);
nor U4275 (N_4275,N_3869,N_3828);
nor U4276 (N_4276,N_3814,N_3640);
and U4277 (N_4277,N_3609,N_3566);
nand U4278 (N_4278,N_3910,N_3601);
xor U4279 (N_4279,N_3983,N_3573);
or U4280 (N_4280,N_3925,N_3795);
and U4281 (N_4281,N_3805,N_3931);
nor U4282 (N_4282,N_3524,N_3848);
or U4283 (N_4283,N_3673,N_3682);
nand U4284 (N_4284,N_3667,N_3778);
nor U4285 (N_4285,N_3649,N_3889);
nand U4286 (N_4286,N_3575,N_3697);
or U4287 (N_4287,N_3976,N_3669);
xor U4288 (N_4288,N_3613,N_3633);
xor U4289 (N_4289,N_3516,N_3728);
nand U4290 (N_4290,N_3715,N_3564);
or U4291 (N_4291,N_3967,N_3808);
or U4292 (N_4292,N_3504,N_3576);
nand U4293 (N_4293,N_3692,N_3789);
and U4294 (N_4294,N_3957,N_3997);
xor U4295 (N_4295,N_3936,N_3984);
xnor U4296 (N_4296,N_3906,N_3988);
xnor U4297 (N_4297,N_3925,N_3643);
or U4298 (N_4298,N_3692,N_3732);
or U4299 (N_4299,N_3720,N_3940);
or U4300 (N_4300,N_3553,N_3723);
or U4301 (N_4301,N_3620,N_3610);
and U4302 (N_4302,N_3724,N_3988);
xnor U4303 (N_4303,N_3907,N_3882);
nand U4304 (N_4304,N_3571,N_3878);
or U4305 (N_4305,N_3661,N_3620);
nand U4306 (N_4306,N_3987,N_3803);
nor U4307 (N_4307,N_3744,N_3740);
nand U4308 (N_4308,N_3974,N_3617);
nor U4309 (N_4309,N_3610,N_3928);
xnor U4310 (N_4310,N_3596,N_3997);
nor U4311 (N_4311,N_3582,N_3923);
xnor U4312 (N_4312,N_3854,N_3513);
nor U4313 (N_4313,N_3611,N_3761);
xnor U4314 (N_4314,N_3827,N_3793);
nor U4315 (N_4315,N_3954,N_3581);
and U4316 (N_4316,N_3849,N_3566);
xor U4317 (N_4317,N_3586,N_3970);
and U4318 (N_4318,N_3783,N_3635);
nand U4319 (N_4319,N_3673,N_3866);
xor U4320 (N_4320,N_3767,N_3626);
or U4321 (N_4321,N_3527,N_3815);
nand U4322 (N_4322,N_3568,N_3546);
nand U4323 (N_4323,N_3884,N_3507);
or U4324 (N_4324,N_3751,N_3760);
nand U4325 (N_4325,N_3627,N_3702);
or U4326 (N_4326,N_3668,N_3941);
and U4327 (N_4327,N_3752,N_3922);
nand U4328 (N_4328,N_3580,N_3915);
or U4329 (N_4329,N_3946,N_3611);
or U4330 (N_4330,N_3648,N_3534);
xor U4331 (N_4331,N_3967,N_3503);
or U4332 (N_4332,N_3859,N_3548);
nand U4333 (N_4333,N_3877,N_3600);
nand U4334 (N_4334,N_3697,N_3849);
nand U4335 (N_4335,N_3771,N_3684);
nor U4336 (N_4336,N_3557,N_3893);
xor U4337 (N_4337,N_3925,N_3873);
or U4338 (N_4338,N_3814,N_3825);
and U4339 (N_4339,N_3967,N_3954);
nor U4340 (N_4340,N_3574,N_3999);
nand U4341 (N_4341,N_3725,N_3690);
xor U4342 (N_4342,N_3747,N_3929);
xor U4343 (N_4343,N_3848,N_3966);
or U4344 (N_4344,N_3987,N_3691);
xor U4345 (N_4345,N_3594,N_3670);
or U4346 (N_4346,N_3530,N_3846);
xor U4347 (N_4347,N_3619,N_3985);
xor U4348 (N_4348,N_3805,N_3820);
nand U4349 (N_4349,N_3621,N_3503);
xor U4350 (N_4350,N_3867,N_3735);
nand U4351 (N_4351,N_3631,N_3647);
nand U4352 (N_4352,N_3816,N_3536);
nor U4353 (N_4353,N_3874,N_3820);
or U4354 (N_4354,N_3761,N_3557);
and U4355 (N_4355,N_3832,N_3825);
xnor U4356 (N_4356,N_3885,N_3988);
nor U4357 (N_4357,N_3582,N_3734);
or U4358 (N_4358,N_3978,N_3838);
nor U4359 (N_4359,N_3643,N_3589);
and U4360 (N_4360,N_3521,N_3874);
xnor U4361 (N_4361,N_3677,N_3955);
nor U4362 (N_4362,N_3944,N_3718);
xor U4363 (N_4363,N_3542,N_3972);
nand U4364 (N_4364,N_3853,N_3511);
nand U4365 (N_4365,N_3585,N_3801);
nand U4366 (N_4366,N_3961,N_3865);
and U4367 (N_4367,N_3818,N_3635);
nand U4368 (N_4368,N_3815,N_3716);
xor U4369 (N_4369,N_3644,N_3604);
and U4370 (N_4370,N_3880,N_3694);
or U4371 (N_4371,N_3558,N_3838);
nand U4372 (N_4372,N_3899,N_3965);
and U4373 (N_4373,N_3666,N_3638);
xor U4374 (N_4374,N_3658,N_3827);
or U4375 (N_4375,N_3967,N_3508);
xnor U4376 (N_4376,N_3923,N_3626);
and U4377 (N_4377,N_3647,N_3590);
xor U4378 (N_4378,N_3839,N_3739);
nand U4379 (N_4379,N_3849,N_3704);
nor U4380 (N_4380,N_3730,N_3781);
and U4381 (N_4381,N_3536,N_3575);
xor U4382 (N_4382,N_3506,N_3837);
nand U4383 (N_4383,N_3783,N_3962);
and U4384 (N_4384,N_3885,N_3990);
nor U4385 (N_4385,N_3993,N_3945);
xor U4386 (N_4386,N_3998,N_3814);
nand U4387 (N_4387,N_3555,N_3732);
nor U4388 (N_4388,N_3717,N_3839);
xor U4389 (N_4389,N_3697,N_3587);
xnor U4390 (N_4390,N_3935,N_3899);
xnor U4391 (N_4391,N_3519,N_3542);
xnor U4392 (N_4392,N_3624,N_3960);
nor U4393 (N_4393,N_3579,N_3622);
nand U4394 (N_4394,N_3546,N_3538);
xnor U4395 (N_4395,N_3669,N_3527);
nand U4396 (N_4396,N_3908,N_3564);
nand U4397 (N_4397,N_3783,N_3678);
nor U4398 (N_4398,N_3523,N_3790);
nand U4399 (N_4399,N_3880,N_3638);
or U4400 (N_4400,N_3680,N_3859);
and U4401 (N_4401,N_3560,N_3837);
nand U4402 (N_4402,N_3871,N_3979);
nor U4403 (N_4403,N_3518,N_3502);
xor U4404 (N_4404,N_3516,N_3711);
nor U4405 (N_4405,N_3801,N_3853);
nand U4406 (N_4406,N_3616,N_3907);
and U4407 (N_4407,N_3929,N_3713);
nor U4408 (N_4408,N_3549,N_3807);
xor U4409 (N_4409,N_3880,N_3846);
xor U4410 (N_4410,N_3718,N_3716);
and U4411 (N_4411,N_3567,N_3675);
and U4412 (N_4412,N_3913,N_3835);
nor U4413 (N_4413,N_3540,N_3586);
nand U4414 (N_4414,N_3681,N_3872);
nand U4415 (N_4415,N_3638,N_3633);
nand U4416 (N_4416,N_3718,N_3922);
nand U4417 (N_4417,N_3597,N_3635);
nor U4418 (N_4418,N_3625,N_3910);
and U4419 (N_4419,N_3603,N_3612);
xor U4420 (N_4420,N_3714,N_3607);
or U4421 (N_4421,N_3850,N_3709);
xor U4422 (N_4422,N_3633,N_3658);
or U4423 (N_4423,N_3846,N_3715);
nand U4424 (N_4424,N_3637,N_3711);
and U4425 (N_4425,N_3739,N_3759);
xnor U4426 (N_4426,N_3535,N_3897);
or U4427 (N_4427,N_3686,N_3900);
or U4428 (N_4428,N_3916,N_3513);
or U4429 (N_4429,N_3642,N_3810);
and U4430 (N_4430,N_3598,N_3557);
and U4431 (N_4431,N_3985,N_3730);
xnor U4432 (N_4432,N_3886,N_3923);
xnor U4433 (N_4433,N_3975,N_3788);
xor U4434 (N_4434,N_3807,N_3655);
nor U4435 (N_4435,N_3500,N_3760);
nor U4436 (N_4436,N_3585,N_3710);
and U4437 (N_4437,N_3733,N_3665);
or U4438 (N_4438,N_3566,N_3684);
or U4439 (N_4439,N_3578,N_3761);
xnor U4440 (N_4440,N_3894,N_3898);
or U4441 (N_4441,N_3658,N_3690);
nand U4442 (N_4442,N_3690,N_3655);
nor U4443 (N_4443,N_3985,N_3818);
or U4444 (N_4444,N_3804,N_3947);
or U4445 (N_4445,N_3700,N_3564);
nor U4446 (N_4446,N_3579,N_3977);
nor U4447 (N_4447,N_3656,N_3873);
and U4448 (N_4448,N_3807,N_3522);
and U4449 (N_4449,N_3953,N_3720);
nor U4450 (N_4450,N_3571,N_3807);
nor U4451 (N_4451,N_3918,N_3980);
nand U4452 (N_4452,N_3677,N_3962);
and U4453 (N_4453,N_3899,N_3944);
nand U4454 (N_4454,N_3532,N_3975);
nor U4455 (N_4455,N_3958,N_3685);
or U4456 (N_4456,N_3747,N_3897);
nand U4457 (N_4457,N_3525,N_3920);
nand U4458 (N_4458,N_3977,N_3914);
or U4459 (N_4459,N_3788,N_3674);
or U4460 (N_4460,N_3736,N_3788);
or U4461 (N_4461,N_3784,N_3691);
xnor U4462 (N_4462,N_3607,N_3588);
or U4463 (N_4463,N_3783,N_3788);
nor U4464 (N_4464,N_3623,N_3529);
nand U4465 (N_4465,N_3774,N_3861);
nand U4466 (N_4466,N_3884,N_3623);
nor U4467 (N_4467,N_3613,N_3625);
and U4468 (N_4468,N_3903,N_3686);
and U4469 (N_4469,N_3694,N_3630);
or U4470 (N_4470,N_3870,N_3932);
xnor U4471 (N_4471,N_3870,N_3803);
xor U4472 (N_4472,N_3911,N_3818);
nand U4473 (N_4473,N_3674,N_3928);
and U4474 (N_4474,N_3897,N_3746);
or U4475 (N_4475,N_3890,N_3679);
xor U4476 (N_4476,N_3772,N_3643);
xnor U4477 (N_4477,N_3627,N_3545);
nand U4478 (N_4478,N_3635,N_3562);
xor U4479 (N_4479,N_3971,N_3707);
nor U4480 (N_4480,N_3903,N_3656);
nand U4481 (N_4481,N_3650,N_3518);
and U4482 (N_4482,N_3806,N_3833);
nor U4483 (N_4483,N_3938,N_3967);
and U4484 (N_4484,N_3723,N_3899);
nor U4485 (N_4485,N_3608,N_3834);
and U4486 (N_4486,N_3669,N_3672);
nor U4487 (N_4487,N_3743,N_3568);
and U4488 (N_4488,N_3862,N_3519);
nor U4489 (N_4489,N_3999,N_3751);
or U4490 (N_4490,N_3706,N_3818);
xnor U4491 (N_4491,N_3911,N_3882);
or U4492 (N_4492,N_3575,N_3968);
nor U4493 (N_4493,N_3987,N_3658);
xor U4494 (N_4494,N_3696,N_3688);
xnor U4495 (N_4495,N_3529,N_3556);
nor U4496 (N_4496,N_3597,N_3756);
nor U4497 (N_4497,N_3635,N_3731);
nor U4498 (N_4498,N_3929,N_3733);
xnor U4499 (N_4499,N_3659,N_3815);
nand U4500 (N_4500,N_4117,N_4242);
nor U4501 (N_4501,N_4044,N_4259);
and U4502 (N_4502,N_4414,N_4022);
xor U4503 (N_4503,N_4009,N_4263);
and U4504 (N_4504,N_4385,N_4171);
or U4505 (N_4505,N_4392,N_4389);
nand U4506 (N_4506,N_4461,N_4393);
and U4507 (N_4507,N_4473,N_4110);
and U4508 (N_4508,N_4452,N_4462);
or U4509 (N_4509,N_4293,N_4247);
and U4510 (N_4510,N_4339,N_4129);
nor U4511 (N_4511,N_4345,N_4152);
nor U4512 (N_4512,N_4341,N_4328);
nand U4513 (N_4513,N_4291,N_4451);
nor U4514 (N_4514,N_4337,N_4409);
nand U4515 (N_4515,N_4240,N_4364);
or U4516 (N_4516,N_4163,N_4442);
and U4517 (N_4517,N_4423,N_4243);
xnor U4518 (N_4518,N_4481,N_4324);
nand U4519 (N_4519,N_4230,N_4064);
nor U4520 (N_4520,N_4225,N_4281);
or U4521 (N_4521,N_4475,N_4241);
and U4522 (N_4522,N_4220,N_4161);
nor U4523 (N_4523,N_4459,N_4380);
nor U4524 (N_4524,N_4218,N_4173);
xor U4525 (N_4525,N_4100,N_4228);
and U4526 (N_4526,N_4415,N_4387);
nor U4527 (N_4527,N_4466,N_4209);
and U4528 (N_4528,N_4499,N_4321);
and U4529 (N_4529,N_4131,N_4288);
nand U4530 (N_4530,N_4125,N_4333);
xor U4531 (N_4531,N_4133,N_4268);
or U4532 (N_4532,N_4011,N_4322);
nor U4533 (N_4533,N_4377,N_4222);
or U4534 (N_4534,N_4060,N_4074);
nor U4535 (N_4535,N_4390,N_4493);
nand U4536 (N_4536,N_4115,N_4283);
nand U4537 (N_4537,N_4182,N_4176);
nand U4538 (N_4538,N_4353,N_4186);
nand U4539 (N_4539,N_4188,N_4034);
or U4540 (N_4540,N_4381,N_4257);
nand U4541 (N_4541,N_4486,N_4149);
or U4542 (N_4542,N_4492,N_4363);
nor U4543 (N_4543,N_4111,N_4172);
or U4544 (N_4544,N_4441,N_4114);
xor U4545 (N_4545,N_4443,N_4253);
nor U4546 (N_4546,N_4083,N_4248);
xor U4547 (N_4547,N_4208,N_4150);
or U4548 (N_4548,N_4046,N_4068);
xor U4549 (N_4549,N_4267,N_4061);
nor U4550 (N_4550,N_4103,N_4296);
xor U4551 (N_4551,N_4198,N_4168);
xnor U4552 (N_4552,N_4399,N_4453);
or U4553 (N_4553,N_4189,N_4421);
nand U4554 (N_4554,N_4223,N_4362);
and U4555 (N_4555,N_4106,N_4043);
or U4556 (N_4556,N_4093,N_4383);
nor U4557 (N_4557,N_4013,N_4231);
xnor U4558 (N_4558,N_4084,N_4407);
nand U4559 (N_4559,N_4138,N_4440);
nand U4560 (N_4560,N_4468,N_4330);
nor U4561 (N_4561,N_4266,N_4376);
and U4562 (N_4562,N_4478,N_4311);
nor U4563 (N_4563,N_4028,N_4431);
nand U4564 (N_4564,N_4275,N_4417);
nor U4565 (N_4565,N_4342,N_4327);
or U4566 (N_4566,N_4312,N_4388);
xor U4567 (N_4567,N_4020,N_4065);
nor U4568 (N_4568,N_4318,N_4360);
xnor U4569 (N_4569,N_4445,N_4206);
nor U4570 (N_4570,N_4356,N_4010);
and U4571 (N_4571,N_4447,N_4406);
and U4572 (N_4572,N_4494,N_4085);
nor U4573 (N_4573,N_4303,N_4167);
and U4574 (N_4574,N_4099,N_4137);
nand U4575 (N_4575,N_4118,N_4252);
nand U4576 (N_4576,N_4140,N_4373);
or U4577 (N_4577,N_4049,N_4207);
nor U4578 (N_4578,N_4216,N_4448);
and U4579 (N_4579,N_4410,N_4413);
nor U4580 (N_4580,N_4256,N_4199);
xor U4581 (N_4581,N_4480,N_4002);
and U4582 (N_4582,N_4098,N_4308);
xor U4583 (N_4583,N_4255,N_4159);
nand U4584 (N_4584,N_4430,N_4076);
or U4585 (N_4585,N_4039,N_4178);
or U4586 (N_4586,N_4316,N_4145);
nor U4587 (N_4587,N_4160,N_4460);
and U4588 (N_4588,N_4340,N_4096);
and U4589 (N_4589,N_4384,N_4403);
nor U4590 (N_4590,N_4136,N_4325);
and U4591 (N_4591,N_4192,N_4151);
xnor U4592 (N_4592,N_4346,N_4144);
xnor U4593 (N_4593,N_4365,N_4033);
nand U4594 (N_4594,N_4395,N_4491);
nor U4595 (N_4595,N_4404,N_4107);
and U4596 (N_4596,N_4334,N_4249);
xor U4597 (N_4597,N_4398,N_4250);
and U4598 (N_4598,N_4057,N_4239);
and U4599 (N_4599,N_4305,N_4052);
xor U4600 (N_4600,N_4338,N_4017);
and U4601 (N_4601,N_4471,N_4048);
xor U4602 (N_4602,N_4201,N_4411);
xor U4603 (N_4603,N_4170,N_4091);
nand U4604 (N_4604,N_4254,N_4235);
xor U4605 (N_4605,N_4246,N_4298);
nand U4606 (N_4606,N_4484,N_4059);
or U4607 (N_4607,N_4141,N_4264);
xor U4608 (N_4608,N_4361,N_4265);
and U4609 (N_4609,N_4439,N_4438);
xnor U4610 (N_4610,N_4301,N_4304);
or U4611 (N_4611,N_4236,N_4032);
nand U4612 (N_4612,N_4273,N_4184);
and U4613 (N_4613,N_4219,N_4154);
nor U4614 (N_4614,N_4300,N_4437);
nand U4615 (N_4615,N_4146,N_4350);
or U4616 (N_4616,N_4204,N_4436);
and U4617 (N_4617,N_4314,N_4457);
nand U4618 (N_4618,N_4205,N_4244);
and U4619 (N_4619,N_4294,N_4224);
nor U4620 (N_4620,N_4262,N_4130);
nand U4621 (N_4621,N_4344,N_4271);
or U4622 (N_4622,N_4086,N_4378);
nand U4623 (N_4623,N_4062,N_4112);
xor U4624 (N_4624,N_4348,N_4433);
and U4625 (N_4625,N_4435,N_4162);
and U4626 (N_4626,N_4232,N_4124);
nor U4627 (N_4627,N_4405,N_4464);
nor U4628 (N_4628,N_4297,N_4007);
and U4629 (N_4629,N_4102,N_4213);
xor U4630 (N_4630,N_4310,N_4026);
and U4631 (N_4631,N_4229,N_4191);
and U4632 (N_4632,N_4221,N_4488);
or U4633 (N_4633,N_4425,N_4142);
or U4634 (N_4634,N_4105,N_4181);
nand U4635 (N_4635,N_4025,N_4367);
xor U4636 (N_4636,N_4444,N_4290);
xor U4637 (N_4637,N_4490,N_4424);
or U4638 (N_4638,N_4183,N_4416);
and U4639 (N_4639,N_4418,N_4391);
nor U4640 (N_4640,N_4012,N_4309);
or U4641 (N_4641,N_4195,N_4200);
xnor U4642 (N_4642,N_4214,N_4428);
and U4643 (N_4643,N_4004,N_4332);
and U4644 (N_4644,N_4366,N_4371);
nor U4645 (N_4645,N_4122,N_4227);
and U4646 (N_4646,N_4212,N_4458);
and U4647 (N_4647,N_4030,N_4147);
xor U4648 (N_4648,N_4467,N_4479);
nor U4649 (N_4649,N_4126,N_4139);
or U4650 (N_4650,N_4067,N_4053);
xnor U4651 (N_4651,N_4238,N_4158);
xor U4652 (N_4652,N_4104,N_4092);
or U4653 (N_4653,N_4432,N_4292);
xor U4654 (N_4654,N_4394,N_4089);
and U4655 (N_4655,N_4317,N_4177);
xnor U4656 (N_4656,N_4455,N_4128);
nor U4657 (N_4657,N_4422,N_4497);
nor U4658 (N_4658,N_4258,N_4279);
and U4659 (N_4659,N_4454,N_4319);
nand U4660 (N_4660,N_4382,N_4295);
xor U4661 (N_4661,N_4023,N_4120);
or U4662 (N_4662,N_4323,N_4038);
and U4663 (N_4663,N_4166,N_4071);
and U4664 (N_4664,N_4108,N_4078);
or U4665 (N_4665,N_4101,N_4088);
nor U4666 (N_4666,N_4031,N_4251);
or U4667 (N_4667,N_4357,N_4097);
and U4668 (N_4668,N_4080,N_4193);
nor U4669 (N_4669,N_4489,N_4000);
nand U4670 (N_4670,N_4054,N_4370);
and U4671 (N_4671,N_4094,N_4197);
nor U4672 (N_4672,N_4226,N_4196);
nor U4673 (N_4673,N_4408,N_4179);
nand U4674 (N_4674,N_4487,N_4302);
nor U4675 (N_4675,N_4157,N_4018);
xnor U4676 (N_4676,N_4335,N_4359);
or U4677 (N_4677,N_4286,N_4374);
nor U4678 (N_4678,N_4355,N_4369);
nand U4679 (N_4679,N_4343,N_4400);
nand U4680 (N_4680,N_4045,N_4069);
nand U4681 (N_4681,N_4190,N_4450);
nor U4682 (N_4682,N_4202,N_4153);
xor U4683 (N_4683,N_4315,N_4278);
nand U4684 (N_4684,N_4477,N_4368);
nor U4685 (N_4685,N_4180,N_4483);
xor U4686 (N_4686,N_4001,N_4082);
nor U4687 (N_4687,N_4386,N_4014);
nand U4688 (N_4688,N_4029,N_4175);
nand U4689 (N_4689,N_4496,N_4051);
or U4690 (N_4690,N_4015,N_4066);
and U4691 (N_4691,N_4070,N_4155);
nand U4692 (N_4692,N_4073,N_4427);
or U4693 (N_4693,N_4289,N_4270);
nor U4694 (N_4694,N_4005,N_4063);
or U4695 (N_4695,N_4284,N_4470);
xnor U4696 (N_4696,N_4215,N_4463);
nor U4697 (N_4697,N_4174,N_4187);
or U4698 (N_4698,N_4260,N_4287);
xnor U4699 (N_4699,N_4021,N_4134);
xnor U4700 (N_4700,N_4465,N_4210);
nor U4701 (N_4701,N_4081,N_4148);
and U4702 (N_4702,N_4420,N_4320);
and U4703 (N_4703,N_4050,N_4397);
xnor U4704 (N_4704,N_4079,N_4003);
nand U4705 (N_4705,N_4027,N_4072);
or U4706 (N_4706,N_4402,N_4349);
or U4707 (N_4707,N_4041,N_4135);
and U4708 (N_4708,N_4412,N_4476);
and U4709 (N_4709,N_4285,N_4329);
xor U4710 (N_4710,N_4156,N_4047);
nor U4711 (N_4711,N_4211,N_4165);
nand U4712 (N_4712,N_4347,N_4234);
and U4713 (N_4713,N_4306,N_4396);
or U4714 (N_4714,N_4261,N_4495);
xnor U4715 (N_4715,N_4282,N_4113);
nand U4716 (N_4716,N_4237,N_4498);
nand U4717 (N_4717,N_4077,N_4016);
xor U4718 (N_4718,N_4307,N_4006);
and U4719 (N_4719,N_4426,N_4372);
and U4720 (N_4720,N_4109,N_4245);
xor U4721 (N_4721,N_4008,N_4035);
and U4722 (N_4722,N_4185,N_4469);
xnor U4723 (N_4723,N_4075,N_4269);
nand U4724 (N_4724,N_4331,N_4123);
nand U4725 (N_4725,N_4058,N_4419);
nor U4726 (N_4726,N_4090,N_4121);
or U4727 (N_4727,N_4401,N_4456);
nor U4728 (N_4728,N_4434,N_4169);
nand U4729 (N_4729,N_4233,N_4116);
xnor U4730 (N_4730,N_4379,N_4095);
nand U4731 (N_4731,N_4217,N_4272);
nor U4732 (N_4732,N_4040,N_4042);
xnor U4733 (N_4733,N_4351,N_4313);
and U4734 (N_4734,N_4299,N_4354);
nand U4735 (N_4735,N_4336,N_4352);
xnor U4736 (N_4736,N_4024,N_4056);
or U4737 (N_4737,N_4358,N_4485);
and U4738 (N_4738,N_4037,N_4429);
xnor U4739 (N_4739,N_4143,N_4132);
or U4740 (N_4740,N_4036,N_4277);
xnor U4741 (N_4741,N_4375,N_4127);
xnor U4742 (N_4742,N_4019,N_4087);
and U4743 (N_4743,N_4194,N_4055);
nor U4744 (N_4744,N_4326,N_4472);
or U4745 (N_4745,N_4274,N_4474);
xor U4746 (N_4746,N_4203,N_4164);
nand U4747 (N_4747,N_4280,N_4482);
or U4748 (N_4748,N_4446,N_4276);
nor U4749 (N_4749,N_4119,N_4449);
and U4750 (N_4750,N_4048,N_4194);
nor U4751 (N_4751,N_4100,N_4239);
nor U4752 (N_4752,N_4441,N_4489);
xor U4753 (N_4753,N_4442,N_4465);
nand U4754 (N_4754,N_4298,N_4046);
xor U4755 (N_4755,N_4167,N_4144);
nor U4756 (N_4756,N_4313,N_4398);
or U4757 (N_4757,N_4242,N_4161);
nand U4758 (N_4758,N_4444,N_4196);
or U4759 (N_4759,N_4076,N_4342);
and U4760 (N_4760,N_4377,N_4149);
and U4761 (N_4761,N_4007,N_4489);
and U4762 (N_4762,N_4407,N_4006);
nand U4763 (N_4763,N_4452,N_4345);
nor U4764 (N_4764,N_4206,N_4080);
nor U4765 (N_4765,N_4045,N_4144);
or U4766 (N_4766,N_4260,N_4381);
xor U4767 (N_4767,N_4194,N_4393);
or U4768 (N_4768,N_4012,N_4231);
xnor U4769 (N_4769,N_4374,N_4278);
nor U4770 (N_4770,N_4051,N_4188);
nand U4771 (N_4771,N_4342,N_4102);
xnor U4772 (N_4772,N_4328,N_4395);
nor U4773 (N_4773,N_4132,N_4179);
nand U4774 (N_4774,N_4412,N_4169);
and U4775 (N_4775,N_4277,N_4280);
and U4776 (N_4776,N_4442,N_4459);
or U4777 (N_4777,N_4008,N_4121);
and U4778 (N_4778,N_4411,N_4139);
nor U4779 (N_4779,N_4418,N_4202);
xor U4780 (N_4780,N_4149,N_4113);
xor U4781 (N_4781,N_4473,N_4412);
nand U4782 (N_4782,N_4316,N_4437);
xor U4783 (N_4783,N_4068,N_4448);
or U4784 (N_4784,N_4370,N_4232);
and U4785 (N_4785,N_4121,N_4224);
or U4786 (N_4786,N_4025,N_4389);
nand U4787 (N_4787,N_4213,N_4128);
and U4788 (N_4788,N_4176,N_4225);
and U4789 (N_4789,N_4004,N_4440);
and U4790 (N_4790,N_4090,N_4203);
and U4791 (N_4791,N_4142,N_4139);
xnor U4792 (N_4792,N_4107,N_4294);
nand U4793 (N_4793,N_4459,N_4422);
nand U4794 (N_4794,N_4045,N_4177);
nand U4795 (N_4795,N_4186,N_4154);
or U4796 (N_4796,N_4059,N_4391);
xor U4797 (N_4797,N_4218,N_4168);
or U4798 (N_4798,N_4379,N_4494);
and U4799 (N_4799,N_4237,N_4428);
nor U4800 (N_4800,N_4089,N_4041);
xor U4801 (N_4801,N_4043,N_4176);
xor U4802 (N_4802,N_4450,N_4320);
and U4803 (N_4803,N_4291,N_4186);
xnor U4804 (N_4804,N_4463,N_4056);
or U4805 (N_4805,N_4327,N_4086);
nor U4806 (N_4806,N_4011,N_4200);
and U4807 (N_4807,N_4130,N_4304);
and U4808 (N_4808,N_4479,N_4403);
xor U4809 (N_4809,N_4324,N_4193);
and U4810 (N_4810,N_4087,N_4360);
and U4811 (N_4811,N_4349,N_4026);
nor U4812 (N_4812,N_4449,N_4341);
and U4813 (N_4813,N_4188,N_4023);
xor U4814 (N_4814,N_4045,N_4075);
xor U4815 (N_4815,N_4076,N_4102);
and U4816 (N_4816,N_4017,N_4248);
or U4817 (N_4817,N_4472,N_4365);
and U4818 (N_4818,N_4326,N_4426);
and U4819 (N_4819,N_4480,N_4447);
and U4820 (N_4820,N_4394,N_4182);
xnor U4821 (N_4821,N_4157,N_4049);
nor U4822 (N_4822,N_4181,N_4329);
nor U4823 (N_4823,N_4445,N_4166);
nor U4824 (N_4824,N_4213,N_4494);
nor U4825 (N_4825,N_4072,N_4370);
nand U4826 (N_4826,N_4209,N_4278);
xor U4827 (N_4827,N_4093,N_4154);
and U4828 (N_4828,N_4415,N_4212);
or U4829 (N_4829,N_4156,N_4225);
nand U4830 (N_4830,N_4029,N_4496);
xor U4831 (N_4831,N_4358,N_4445);
and U4832 (N_4832,N_4007,N_4272);
nor U4833 (N_4833,N_4437,N_4318);
and U4834 (N_4834,N_4418,N_4246);
nor U4835 (N_4835,N_4025,N_4152);
or U4836 (N_4836,N_4263,N_4095);
and U4837 (N_4837,N_4349,N_4285);
nand U4838 (N_4838,N_4264,N_4397);
or U4839 (N_4839,N_4200,N_4305);
or U4840 (N_4840,N_4494,N_4316);
nand U4841 (N_4841,N_4123,N_4058);
or U4842 (N_4842,N_4074,N_4089);
and U4843 (N_4843,N_4495,N_4019);
xor U4844 (N_4844,N_4012,N_4458);
or U4845 (N_4845,N_4467,N_4272);
nor U4846 (N_4846,N_4060,N_4386);
nor U4847 (N_4847,N_4264,N_4275);
or U4848 (N_4848,N_4487,N_4054);
and U4849 (N_4849,N_4355,N_4392);
and U4850 (N_4850,N_4428,N_4462);
nor U4851 (N_4851,N_4449,N_4446);
nor U4852 (N_4852,N_4263,N_4224);
and U4853 (N_4853,N_4216,N_4073);
xnor U4854 (N_4854,N_4069,N_4065);
nand U4855 (N_4855,N_4090,N_4360);
xor U4856 (N_4856,N_4452,N_4394);
nand U4857 (N_4857,N_4314,N_4363);
and U4858 (N_4858,N_4199,N_4099);
nand U4859 (N_4859,N_4447,N_4382);
xnor U4860 (N_4860,N_4127,N_4067);
and U4861 (N_4861,N_4301,N_4220);
xnor U4862 (N_4862,N_4063,N_4125);
nor U4863 (N_4863,N_4465,N_4328);
or U4864 (N_4864,N_4323,N_4279);
and U4865 (N_4865,N_4437,N_4409);
nor U4866 (N_4866,N_4171,N_4353);
or U4867 (N_4867,N_4188,N_4423);
xnor U4868 (N_4868,N_4431,N_4495);
nor U4869 (N_4869,N_4036,N_4342);
and U4870 (N_4870,N_4347,N_4476);
xor U4871 (N_4871,N_4089,N_4266);
xor U4872 (N_4872,N_4423,N_4048);
nor U4873 (N_4873,N_4081,N_4169);
or U4874 (N_4874,N_4162,N_4110);
xor U4875 (N_4875,N_4279,N_4094);
nor U4876 (N_4876,N_4436,N_4383);
nand U4877 (N_4877,N_4481,N_4254);
nor U4878 (N_4878,N_4322,N_4007);
xor U4879 (N_4879,N_4241,N_4009);
and U4880 (N_4880,N_4415,N_4008);
xnor U4881 (N_4881,N_4348,N_4168);
and U4882 (N_4882,N_4489,N_4426);
nor U4883 (N_4883,N_4222,N_4415);
and U4884 (N_4884,N_4043,N_4268);
nor U4885 (N_4885,N_4095,N_4449);
and U4886 (N_4886,N_4246,N_4443);
nor U4887 (N_4887,N_4469,N_4068);
or U4888 (N_4888,N_4363,N_4203);
and U4889 (N_4889,N_4293,N_4312);
and U4890 (N_4890,N_4120,N_4098);
and U4891 (N_4891,N_4366,N_4026);
xnor U4892 (N_4892,N_4023,N_4499);
and U4893 (N_4893,N_4138,N_4391);
xor U4894 (N_4894,N_4174,N_4368);
nand U4895 (N_4895,N_4237,N_4010);
nor U4896 (N_4896,N_4281,N_4372);
or U4897 (N_4897,N_4319,N_4436);
nand U4898 (N_4898,N_4083,N_4389);
and U4899 (N_4899,N_4344,N_4135);
or U4900 (N_4900,N_4408,N_4287);
nor U4901 (N_4901,N_4263,N_4358);
or U4902 (N_4902,N_4213,N_4171);
and U4903 (N_4903,N_4059,N_4411);
nor U4904 (N_4904,N_4304,N_4442);
xnor U4905 (N_4905,N_4225,N_4311);
xnor U4906 (N_4906,N_4348,N_4250);
nor U4907 (N_4907,N_4144,N_4328);
and U4908 (N_4908,N_4125,N_4364);
and U4909 (N_4909,N_4007,N_4232);
nand U4910 (N_4910,N_4011,N_4483);
nand U4911 (N_4911,N_4356,N_4021);
nand U4912 (N_4912,N_4434,N_4177);
nand U4913 (N_4913,N_4006,N_4011);
xnor U4914 (N_4914,N_4158,N_4106);
and U4915 (N_4915,N_4440,N_4346);
or U4916 (N_4916,N_4180,N_4161);
and U4917 (N_4917,N_4235,N_4375);
or U4918 (N_4918,N_4402,N_4294);
xnor U4919 (N_4919,N_4426,N_4323);
or U4920 (N_4920,N_4474,N_4349);
xnor U4921 (N_4921,N_4363,N_4385);
nand U4922 (N_4922,N_4489,N_4309);
or U4923 (N_4923,N_4274,N_4243);
xnor U4924 (N_4924,N_4245,N_4195);
xnor U4925 (N_4925,N_4265,N_4046);
nand U4926 (N_4926,N_4264,N_4109);
nor U4927 (N_4927,N_4130,N_4038);
nand U4928 (N_4928,N_4170,N_4413);
nor U4929 (N_4929,N_4222,N_4338);
or U4930 (N_4930,N_4264,N_4170);
nand U4931 (N_4931,N_4418,N_4301);
nand U4932 (N_4932,N_4112,N_4123);
and U4933 (N_4933,N_4237,N_4158);
nor U4934 (N_4934,N_4452,N_4141);
or U4935 (N_4935,N_4334,N_4140);
nand U4936 (N_4936,N_4097,N_4497);
xnor U4937 (N_4937,N_4048,N_4033);
xnor U4938 (N_4938,N_4100,N_4332);
nor U4939 (N_4939,N_4320,N_4185);
nand U4940 (N_4940,N_4009,N_4448);
or U4941 (N_4941,N_4419,N_4013);
nor U4942 (N_4942,N_4058,N_4111);
or U4943 (N_4943,N_4185,N_4213);
and U4944 (N_4944,N_4273,N_4090);
nand U4945 (N_4945,N_4175,N_4366);
xnor U4946 (N_4946,N_4419,N_4410);
nand U4947 (N_4947,N_4113,N_4407);
or U4948 (N_4948,N_4108,N_4385);
nor U4949 (N_4949,N_4057,N_4455);
nand U4950 (N_4950,N_4140,N_4476);
xor U4951 (N_4951,N_4176,N_4232);
and U4952 (N_4952,N_4114,N_4263);
xnor U4953 (N_4953,N_4078,N_4127);
xnor U4954 (N_4954,N_4387,N_4209);
nor U4955 (N_4955,N_4342,N_4412);
nand U4956 (N_4956,N_4240,N_4370);
nand U4957 (N_4957,N_4042,N_4034);
or U4958 (N_4958,N_4477,N_4291);
xor U4959 (N_4959,N_4477,N_4353);
or U4960 (N_4960,N_4105,N_4407);
nor U4961 (N_4961,N_4301,N_4118);
nand U4962 (N_4962,N_4099,N_4425);
and U4963 (N_4963,N_4068,N_4285);
and U4964 (N_4964,N_4243,N_4493);
nand U4965 (N_4965,N_4462,N_4138);
xor U4966 (N_4966,N_4443,N_4231);
nor U4967 (N_4967,N_4383,N_4396);
and U4968 (N_4968,N_4174,N_4442);
nand U4969 (N_4969,N_4166,N_4444);
and U4970 (N_4970,N_4067,N_4169);
nand U4971 (N_4971,N_4439,N_4468);
xor U4972 (N_4972,N_4361,N_4004);
nand U4973 (N_4973,N_4272,N_4065);
nor U4974 (N_4974,N_4122,N_4379);
and U4975 (N_4975,N_4159,N_4443);
nor U4976 (N_4976,N_4062,N_4129);
nor U4977 (N_4977,N_4443,N_4143);
xor U4978 (N_4978,N_4319,N_4145);
nor U4979 (N_4979,N_4003,N_4389);
or U4980 (N_4980,N_4018,N_4290);
xnor U4981 (N_4981,N_4087,N_4188);
xor U4982 (N_4982,N_4259,N_4381);
nor U4983 (N_4983,N_4483,N_4447);
and U4984 (N_4984,N_4063,N_4483);
nand U4985 (N_4985,N_4188,N_4239);
nor U4986 (N_4986,N_4309,N_4367);
or U4987 (N_4987,N_4205,N_4285);
or U4988 (N_4988,N_4055,N_4057);
nor U4989 (N_4989,N_4449,N_4244);
nor U4990 (N_4990,N_4259,N_4187);
nand U4991 (N_4991,N_4177,N_4208);
nor U4992 (N_4992,N_4087,N_4176);
nand U4993 (N_4993,N_4251,N_4181);
and U4994 (N_4994,N_4446,N_4122);
or U4995 (N_4995,N_4193,N_4047);
nand U4996 (N_4996,N_4443,N_4008);
xor U4997 (N_4997,N_4463,N_4473);
nand U4998 (N_4998,N_4350,N_4241);
xor U4999 (N_4999,N_4392,N_4070);
or U5000 (N_5000,N_4591,N_4856);
xor U5001 (N_5001,N_4762,N_4649);
or U5002 (N_5002,N_4726,N_4703);
nor U5003 (N_5003,N_4826,N_4537);
nand U5004 (N_5004,N_4644,N_4954);
or U5005 (N_5005,N_4776,N_4522);
and U5006 (N_5006,N_4566,N_4584);
nand U5007 (N_5007,N_4756,N_4679);
and U5008 (N_5008,N_4560,N_4805);
and U5009 (N_5009,N_4643,N_4528);
nor U5010 (N_5010,N_4606,N_4747);
and U5011 (N_5011,N_4675,N_4695);
and U5012 (N_5012,N_4790,N_4562);
nand U5013 (N_5013,N_4975,N_4713);
nand U5014 (N_5014,N_4834,N_4853);
nor U5015 (N_5015,N_4585,N_4665);
xor U5016 (N_5016,N_4629,N_4851);
nor U5017 (N_5017,N_4594,N_4792);
nand U5018 (N_5018,N_4508,N_4933);
nand U5019 (N_5019,N_4773,N_4614);
and U5020 (N_5020,N_4619,N_4563);
nor U5021 (N_5021,N_4752,N_4577);
nand U5022 (N_5022,N_4727,N_4890);
or U5023 (N_5023,N_4961,N_4574);
xor U5024 (N_5024,N_4758,N_4955);
and U5025 (N_5025,N_4902,N_4876);
nand U5026 (N_5026,N_4745,N_4559);
nor U5027 (N_5027,N_4882,N_4832);
xor U5028 (N_5028,N_4770,N_4578);
or U5029 (N_5029,N_4716,N_4894);
and U5030 (N_5030,N_4945,N_4901);
nor U5031 (N_5031,N_4870,N_4929);
nor U5032 (N_5032,N_4605,N_4564);
xnor U5033 (N_5033,N_4788,N_4859);
nor U5034 (N_5034,N_4811,N_4728);
xnor U5035 (N_5035,N_4698,N_4922);
and U5036 (N_5036,N_4583,N_4668);
nor U5037 (N_5037,N_4991,N_4871);
xor U5038 (N_5038,N_4904,N_4608);
xnor U5039 (N_5039,N_4631,N_4927);
nor U5040 (N_5040,N_4514,N_4539);
or U5041 (N_5041,N_4828,N_4952);
or U5042 (N_5042,N_4587,N_4896);
or U5043 (N_5043,N_4694,N_4823);
and U5044 (N_5044,N_4979,N_4656);
xnor U5045 (N_5045,N_4915,N_4985);
xor U5046 (N_5046,N_4576,N_4877);
xor U5047 (N_5047,N_4573,N_4645);
or U5048 (N_5048,N_4857,N_4647);
nand U5049 (N_5049,N_4978,N_4742);
and U5050 (N_5050,N_4808,N_4994);
xor U5051 (N_5051,N_4569,N_4535);
nor U5052 (N_5052,N_4783,N_4542);
xnor U5053 (N_5053,N_4774,N_4516);
and U5054 (N_5054,N_4884,N_4504);
nand U5055 (N_5055,N_4527,N_4682);
nor U5056 (N_5056,N_4814,N_4612);
and U5057 (N_5057,N_4845,N_4532);
and U5058 (N_5058,N_4604,N_4976);
nand U5059 (N_5059,N_4864,N_4920);
nor U5060 (N_5060,N_4771,N_4586);
xnor U5061 (N_5061,N_4861,N_4930);
and U5062 (N_5062,N_4717,N_4813);
or U5063 (N_5063,N_4893,N_4900);
or U5064 (N_5064,N_4820,N_4767);
and U5065 (N_5065,N_4691,N_4670);
nand U5066 (N_5066,N_4720,N_4730);
nand U5067 (N_5067,N_4622,N_4638);
and U5068 (N_5068,N_4924,N_4648);
or U5069 (N_5069,N_4772,N_4939);
nor U5070 (N_5070,N_4719,N_4642);
nand U5071 (N_5071,N_4686,N_4872);
nor U5072 (N_5072,N_4570,N_4838);
or U5073 (N_5073,N_4709,N_4948);
xnor U5074 (N_5074,N_4541,N_4750);
xnor U5075 (N_5075,N_4699,N_4545);
xor U5076 (N_5076,N_4879,N_4715);
nor U5077 (N_5077,N_4690,N_4681);
xor U5078 (N_5078,N_4754,N_4751);
or U5079 (N_5079,N_4797,N_4941);
and U5080 (N_5080,N_4618,N_4530);
xnor U5081 (N_5081,N_4980,N_4867);
nand U5082 (N_5082,N_4819,N_4950);
nand U5083 (N_5083,N_4959,N_4844);
or U5084 (N_5084,N_4680,N_4780);
nor U5085 (N_5085,N_4520,N_4610);
nor U5086 (N_5086,N_4740,N_4887);
nand U5087 (N_5087,N_4692,N_4889);
nor U5088 (N_5088,N_4635,N_4982);
nand U5089 (N_5089,N_4916,N_4860);
and U5090 (N_5090,N_4589,N_4503);
xnor U5091 (N_5091,N_4966,N_4546);
xnor U5092 (N_5092,N_4628,N_4613);
nor U5093 (N_5093,N_4969,N_4880);
or U5094 (N_5094,N_4700,N_4934);
and U5095 (N_5095,N_4580,N_4689);
nor U5096 (N_5096,N_4718,N_4885);
nor U5097 (N_5097,N_4623,N_4654);
nand U5098 (N_5098,N_4662,N_4993);
xor U5099 (N_5099,N_4852,N_4624);
xor U5100 (N_5100,N_4911,N_4658);
xnor U5101 (N_5101,N_4509,N_4737);
xor U5102 (N_5102,N_4968,N_4626);
nor U5103 (N_5103,N_4803,N_4731);
nand U5104 (N_5104,N_4914,N_4734);
nand U5105 (N_5105,N_4725,N_4855);
nand U5106 (N_5106,N_4972,N_4723);
nand U5107 (N_5107,N_4651,N_4794);
or U5108 (N_5108,N_4778,N_4661);
and U5109 (N_5109,N_4843,N_4942);
nor U5110 (N_5110,N_4704,N_4502);
or U5111 (N_5111,N_4932,N_4536);
nor U5112 (N_5112,N_4678,N_4739);
nor U5113 (N_5113,N_4607,N_4997);
and U5114 (N_5114,N_4664,N_4946);
nor U5115 (N_5115,N_4990,N_4553);
xnor U5116 (N_5116,N_4749,N_4839);
xor U5117 (N_5117,N_4525,N_4974);
nand U5118 (N_5118,N_4673,N_4935);
xnor U5119 (N_5119,N_4873,N_4837);
and U5120 (N_5120,N_4706,N_4818);
or U5121 (N_5121,N_4995,N_4663);
or U5122 (N_5122,N_4903,N_4633);
or U5123 (N_5123,N_4555,N_4802);
or U5124 (N_5124,N_4722,N_4791);
xnor U5125 (N_5125,N_4676,N_4962);
or U5126 (N_5126,N_4599,N_4653);
nand U5127 (N_5127,N_4983,N_4785);
and U5128 (N_5128,N_4511,N_4895);
nor U5129 (N_5129,N_4641,N_4907);
nand U5130 (N_5130,N_4875,N_4593);
or U5131 (N_5131,N_4898,N_4846);
or U5132 (N_5132,N_4741,N_4830);
and U5133 (N_5133,N_4616,N_4765);
xnor U5134 (N_5134,N_4977,N_4971);
or U5135 (N_5135,N_4913,N_4646);
xnor U5136 (N_5136,N_4878,N_4696);
or U5137 (N_5137,N_4804,N_4840);
nand U5138 (N_5138,N_4825,N_4567);
nand U5139 (N_5139,N_4981,N_4669);
and U5140 (N_5140,N_4630,N_4777);
and U5141 (N_5141,N_4708,N_4923);
and U5142 (N_5142,N_4519,N_4921);
nand U5143 (N_5143,N_4824,N_4829);
nor U5144 (N_5144,N_4854,N_4781);
nor U5145 (N_5145,N_4822,N_4886);
nor U5146 (N_5146,N_4554,N_4620);
and U5147 (N_5147,N_4766,N_4501);
nand U5148 (N_5148,N_4906,N_4517);
or U5149 (N_5149,N_4757,N_4561);
or U5150 (N_5150,N_4634,N_4849);
and U5151 (N_5151,N_4659,N_4784);
or U5152 (N_5152,N_4833,N_4515);
nand U5153 (N_5153,N_4609,N_4547);
or U5154 (N_5154,N_4786,N_4986);
nand U5155 (N_5155,N_4523,N_4881);
nor U5156 (N_5156,N_4625,N_4711);
or U5157 (N_5157,N_4836,N_4685);
and U5158 (N_5158,N_4973,N_4568);
nor U5159 (N_5159,N_4600,N_4572);
nand U5160 (N_5160,N_4964,N_4735);
and U5161 (N_5161,N_4714,N_4697);
nand U5162 (N_5162,N_4759,N_4806);
xor U5163 (N_5163,N_4817,N_4831);
and U5164 (N_5164,N_4905,N_4672);
nand U5165 (N_5165,N_4755,N_4506);
nor U5166 (N_5166,N_4666,N_4926);
and U5167 (N_5167,N_4960,N_4603);
nor U5168 (N_5168,N_4507,N_4512);
nand U5169 (N_5169,N_4639,N_4958);
xnor U5170 (N_5170,N_4611,N_4534);
nand U5171 (N_5171,N_4588,N_4888);
and U5172 (N_5172,N_4571,N_4540);
nand U5173 (N_5173,N_4650,N_4866);
nand U5174 (N_5174,N_4892,N_4760);
xor U5175 (N_5175,N_4732,N_4556);
nand U5176 (N_5176,N_4660,N_4575);
nor U5177 (N_5177,N_4744,N_4524);
xor U5178 (N_5178,N_4816,N_4518);
or U5179 (N_5179,N_4917,N_4544);
or U5180 (N_5180,N_4531,N_4683);
or U5181 (N_5181,N_4827,N_4768);
and U5182 (N_5182,N_4919,N_4705);
xnor U5183 (N_5183,N_4500,N_4764);
or U5184 (N_5184,N_4931,N_4850);
xor U5185 (N_5185,N_4807,N_4565);
and U5186 (N_5186,N_4582,N_4733);
xor U5187 (N_5187,N_4912,N_4693);
nand U5188 (N_5188,N_4655,N_4842);
or U5189 (N_5189,N_4909,N_4949);
nor U5190 (N_5190,N_4763,N_4769);
nor U5191 (N_5191,N_4615,N_4543);
nor U5192 (N_5192,N_4748,N_4883);
nor U5193 (N_5193,N_4652,N_4590);
or U5194 (N_5194,N_4796,N_4897);
xor U5195 (N_5195,N_4684,N_4841);
and U5196 (N_5196,N_4538,N_4953);
and U5197 (N_5197,N_4989,N_4899);
nor U5198 (N_5198,N_4992,N_4812);
or U5199 (N_5199,N_4738,N_4984);
xor U5200 (N_5200,N_4549,N_4835);
nand U5201 (N_5201,N_4558,N_4918);
xor U5202 (N_5202,N_4598,N_4970);
and U5203 (N_5203,N_4956,N_4951);
xor U5204 (N_5204,N_4874,N_4782);
nor U5205 (N_5205,N_4967,N_4801);
xor U5206 (N_5206,N_4937,N_4550);
nand U5207 (N_5207,N_4637,N_4779);
and U5208 (N_5208,N_4848,N_4533);
xnor U5209 (N_5209,N_4677,N_4800);
nand U5210 (N_5210,N_4999,N_4761);
nand U5211 (N_5211,N_4721,N_4998);
nand U5212 (N_5212,N_4551,N_4938);
xnor U5213 (N_5213,N_4636,N_4557);
and U5214 (N_5214,N_4601,N_4908);
nor U5215 (N_5215,N_4710,N_4957);
xor U5216 (N_5216,N_4510,N_4799);
and U5217 (N_5217,N_4513,N_4940);
and U5218 (N_5218,N_4862,N_4775);
or U5219 (N_5219,N_4596,N_4526);
and U5220 (N_5220,N_4963,N_4858);
xnor U5221 (N_5221,N_4617,N_4701);
nand U5222 (N_5222,N_4793,N_4729);
xor U5223 (N_5223,N_4743,N_4687);
or U5224 (N_5224,N_4910,N_4815);
nand U5225 (N_5225,N_4809,N_4581);
nand U5226 (N_5226,N_4621,N_4505);
xor U5227 (N_5227,N_4521,N_4640);
nor U5228 (N_5228,N_4865,N_4746);
xnor U5229 (N_5229,N_4712,N_4552);
and U5230 (N_5230,N_4671,N_4579);
nor U5231 (N_5231,N_4529,N_4798);
xnor U5232 (N_5232,N_4702,N_4674);
nand U5233 (N_5233,N_4657,N_4928);
nand U5234 (N_5234,N_4548,N_4724);
and U5235 (N_5235,N_4996,N_4936);
or U5236 (N_5236,N_4868,N_4632);
xor U5237 (N_5237,N_4891,N_4592);
or U5238 (N_5238,N_4988,N_4863);
or U5239 (N_5239,N_4943,N_4627);
and U5240 (N_5240,N_4925,N_4821);
and U5241 (N_5241,N_4795,N_4789);
nand U5242 (N_5242,N_4602,N_4987);
or U5243 (N_5243,N_4667,N_4595);
nor U5244 (N_5244,N_4597,N_4965);
nor U5245 (N_5245,N_4688,N_4869);
xnor U5246 (N_5246,N_4944,N_4810);
xnor U5247 (N_5247,N_4736,N_4847);
xor U5248 (N_5248,N_4707,N_4947);
and U5249 (N_5249,N_4753,N_4787);
xor U5250 (N_5250,N_4868,N_4533);
and U5251 (N_5251,N_4818,N_4921);
xor U5252 (N_5252,N_4992,N_4691);
nand U5253 (N_5253,N_4544,N_4577);
nor U5254 (N_5254,N_4632,N_4919);
and U5255 (N_5255,N_4512,N_4683);
or U5256 (N_5256,N_4896,N_4906);
nand U5257 (N_5257,N_4831,N_4854);
and U5258 (N_5258,N_4651,N_4580);
xor U5259 (N_5259,N_4641,N_4539);
or U5260 (N_5260,N_4634,N_4970);
nor U5261 (N_5261,N_4893,N_4714);
nand U5262 (N_5262,N_4849,N_4547);
nand U5263 (N_5263,N_4584,N_4658);
nand U5264 (N_5264,N_4584,N_4512);
nand U5265 (N_5265,N_4693,N_4762);
xnor U5266 (N_5266,N_4947,N_4781);
nand U5267 (N_5267,N_4866,N_4738);
xnor U5268 (N_5268,N_4916,N_4681);
nor U5269 (N_5269,N_4901,N_4585);
and U5270 (N_5270,N_4501,N_4739);
nand U5271 (N_5271,N_4590,N_4879);
and U5272 (N_5272,N_4980,N_4509);
xnor U5273 (N_5273,N_4674,N_4736);
nand U5274 (N_5274,N_4852,N_4660);
and U5275 (N_5275,N_4988,N_4616);
or U5276 (N_5276,N_4823,N_4529);
nand U5277 (N_5277,N_4786,N_4880);
nand U5278 (N_5278,N_4697,N_4743);
and U5279 (N_5279,N_4853,N_4584);
nor U5280 (N_5280,N_4553,N_4837);
nor U5281 (N_5281,N_4675,N_4636);
nand U5282 (N_5282,N_4833,N_4809);
xor U5283 (N_5283,N_4757,N_4836);
and U5284 (N_5284,N_4604,N_4720);
nand U5285 (N_5285,N_4648,N_4610);
nand U5286 (N_5286,N_4872,N_4916);
xnor U5287 (N_5287,N_4836,N_4831);
nand U5288 (N_5288,N_4879,N_4611);
nand U5289 (N_5289,N_4915,N_4686);
nor U5290 (N_5290,N_4843,N_4875);
nor U5291 (N_5291,N_4985,N_4692);
or U5292 (N_5292,N_4979,N_4992);
and U5293 (N_5293,N_4539,N_4910);
or U5294 (N_5294,N_4645,N_4951);
and U5295 (N_5295,N_4774,N_4588);
or U5296 (N_5296,N_4677,N_4750);
nor U5297 (N_5297,N_4916,N_4888);
nand U5298 (N_5298,N_4875,N_4918);
nand U5299 (N_5299,N_4972,N_4727);
or U5300 (N_5300,N_4827,N_4881);
nor U5301 (N_5301,N_4631,N_4542);
nor U5302 (N_5302,N_4746,N_4695);
and U5303 (N_5303,N_4617,N_4918);
or U5304 (N_5304,N_4638,N_4619);
and U5305 (N_5305,N_4862,N_4746);
xor U5306 (N_5306,N_4683,N_4519);
and U5307 (N_5307,N_4609,N_4527);
nor U5308 (N_5308,N_4917,N_4683);
and U5309 (N_5309,N_4523,N_4508);
nor U5310 (N_5310,N_4539,N_4822);
or U5311 (N_5311,N_4949,N_4811);
and U5312 (N_5312,N_4946,N_4884);
nor U5313 (N_5313,N_4995,N_4771);
or U5314 (N_5314,N_4667,N_4811);
xor U5315 (N_5315,N_4573,N_4511);
nand U5316 (N_5316,N_4750,N_4593);
or U5317 (N_5317,N_4805,N_4571);
xnor U5318 (N_5318,N_4601,N_4507);
nand U5319 (N_5319,N_4807,N_4714);
nor U5320 (N_5320,N_4819,N_4644);
nand U5321 (N_5321,N_4641,N_4667);
or U5322 (N_5322,N_4956,N_4510);
or U5323 (N_5323,N_4961,N_4777);
and U5324 (N_5324,N_4514,N_4948);
xor U5325 (N_5325,N_4735,N_4884);
nand U5326 (N_5326,N_4730,N_4712);
xnor U5327 (N_5327,N_4772,N_4994);
xnor U5328 (N_5328,N_4543,N_4568);
or U5329 (N_5329,N_4606,N_4766);
nand U5330 (N_5330,N_4762,N_4522);
nor U5331 (N_5331,N_4772,N_4513);
nand U5332 (N_5332,N_4661,N_4779);
xor U5333 (N_5333,N_4771,N_4974);
or U5334 (N_5334,N_4914,N_4690);
xor U5335 (N_5335,N_4728,N_4887);
xor U5336 (N_5336,N_4742,N_4883);
xnor U5337 (N_5337,N_4749,N_4778);
nand U5338 (N_5338,N_4930,N_4909);
nand U5339 (N_5339,N_4837,N_4732);
or U5340 (N_5340,N_4998,N_4670);
or U5341 (N_5341,N_4592,N_4558);
nand U5342 (N_5342,N_4645,N_4653);
or U5343 (N_5343,N_4544,N_4903);
xor U5344 (N_5344,N_4831,N_4691);
nor U5345 (N_5345,N_4581,N_4664);
or U5346 (N_5346,N_4720,N_4685);
xor U5347 (N_5347,N_4985,N_4988);
xnor U5348 (N_5348,N_4971,N_4849);
and U5349 (N_5349,N_4587,N_4862);
nor U5350 (N_5350,N_4562,N_4569);
xor U5351 (N_5351,N_4888,N_4808);
nand U5352 (N_5352,N_4812,N_4525);
and U5353 (N_5353,N_4561,N_4980);
nand U5354 (N_5354,N_4655,N_4724);
nand U5355 (N_5355,N_4731,N_4771);
nand U5356 (N_5356,N_4509,N_4720);
xnor U5357 (N_5357,N_4719,N_4762);
nand U5358 (N_5358,N_4552,N_4566);
nor U5359 (N_5359,N_4659,N_4888);
nand U5360 (N_5360,N_4757,N_4870);
or U5361 (N_5361,N_4609,N_4928);
xor U5362 (N_5362,N_4798,N_4944);
and U5363 (N_5363,N_4638,N_4898);
and U5364 (N_5364,N_4911,N_4672);
nand U5365 (N_5365,N_4533,N_4806);
nand U5366 (N_5366,N_4821,N_4673);
or U5367 (N_5367,N_4602,N_4543);
or U5368 (N_5368,N_4963,N_4818);
nor U5369 (N_5369,N_4501,N_4528);
and U5370 (N_5370,N_4703,N_4587);
xnor U5371 (N_5371,N_4977,N_4634);
and U5372 (N_5372,N_4637,N_4652);
xnor U5373 (N_5373,N_4830,N_4751);
nand U5374 (N_5374,N_4518,N_4717);
nand U5375 (N_5375,N_4795,N_4635);
xor U5376 (N_5376,N_4918,N_4914);
nand U5377 (N_5377,N_4804,N_4667);
nor U5378 (N_5378,N_4739,N_4749);
xnor U5379 (N_5379,N_4925,N_4652);
nor U5380 (N_5380,N_4667,N_4750);
or U5381 (N_5381,N_4790,N_4781);
xnor U5382 (N_5382,N_4923,N_4574);
xor U5383 (N_5383,N_4866,N_4686);
xor U5384 (N_5384,N_4939,N_4538);
or U5385 (N_5385,N_4668,N_4572);
or U5386 (N_5386,N_4849,N_4765);
nor U5387 (N_5387,N_4518,N_4651);
xor U5388 (N_5388,N_4637,N_4769);
and U5389 (N_5389,N_4981,N_4947);
nand U5390 (N_5390,N_4654,N_4852);
and U5391 (N_5391,N_4770,N_4744);
or U5392 (N_5392,N_4775,N_4743);
nand U5393 (N_5393,N_4680,N_4884);
and U5394 (N_5394,N_4702,N_4523);
or U5395 (N_5395,N_4998,N_4926);
and U5396 (N_5396,N_4776,N_4907);
and U5397 (N_5397,N_4565,N_4715);
or U5398 (N_5398,N_4877,N_4672);
xnor U5399 (N_5399,N_4582,N_4835);
nor U5400 (N_5400,N_4594,N_4740);
nand U5401 (N_5401,N_4975,N_4870);
and U5402 (N_5402,N_4502,N_4791);
xor U5403 (N_5403,N_4991,N_4586);
and U5404 (N_5404,N_4674,N_4839);
or U5405 (N_5405,N_4882,N_4999);
and U5406 (N_5406,N_4931,N_4954);
xnor U5407 (N_5407,N_4964,N_4548);
or U5408 (N_5408,N_4625,N_4748);
xnor U5409 (N_5409,N_4917,N_4825);
xor U5410 (N_5410,N_4676,N_4588);
nand U5411 (N_5411,N_4814,N_4935);
or U5412 (N_5412,N_4511,N_4818);
or U5413 (N_5413,N_4869,N_4925);
xor U5414 (N_5414,N_4683,N_4518);
xnor U5415 (N_5415,N_4670,N_4568);
and U5416 (N_5416,N_4931,N_4839);
xnor U5417 (N_5417,N_4556,N_4833);
xor U5418 (N_5418,N_4715,N_4901);
or U5419 (N_5419,N_4759,N_4534);
or U5420 (N_5420,N_4618,N_4750);
or U5421 (N_5421,N_4931,N_4847);
or U5422 (N_5422,N_4531,N_4574);
xor U5423 (N_5423,N_4933,N_4688);
nor U5424 (N_5424,N_4959,N_4905);
and U5425 (N_5425,N_4524,N_4592);
or U5426 (N_5426,N_4613,N_4962);
xor U5427 (N_5427,N_4570,N_4921);
nand U5428 (N_5428,N_4871,N_4754);
and U5429 (N_5429,N_4584,N_4902);
or U5430 (N_5430,N_4833,N_4869);
nand U5431 (N_5431,N_4847,N_4828);
xor U5432 (N_5432,N_4806,N_4666);
xnor U5433 (N_5433,N_4715,N_4515);
nor U5434 (N_5434,N_4856,N_4740);
xnor U5435 (N_5435,N_4693,N_4875);
nor U5436 (N_5436,N_4793,N_4912);
nand U5437 (N_5437,N_4865,N_4738);
or U5438 (N_5438,N_4760,N_4527);
xor U5439 (N_5439,N_4778,N_4962);
and U5440 (N_5440,N_4573,N_4633);
or U5441 (N_5441,N_4630,N_4680);
nand U5442 (N_5442,N_4549,N_4842);
or U5443 (N_5443,N_4535,N_4741);
nand U5444 (N_5444,N_4778,N_4665);
xnor U5445 (N_5445,N_4650,N_4976);
nor U5446 (N_5446,N_4925,N_4803);
nor U5447 (N_5447,N_4502,N_4546);
and U5448 (N_5448,N_4950,N_4527);
and U5449 (N_5449,N_4825,N_4971);
or U5450 (N_5450,N_4933,N_4559);
or U5451 (N_5451,N_4977,N_4941);
and U5452 (N_5452,N_4836,N_4596);
xor U5453 (N_5453,N_4842,N_4913);
or U5454 (N_5454,N_4899,N_4609);
or U5455 (N_5455,N_4576,N_4580);
or U5456 (N_5456,N_4682,N_4735);
and U5457 (N_5457,N_4804,N_4501);
nand U5458 (N_5458,N_4998,N_4589);
and U5459 (N_5459,N_4706,N_4992);
nand U5460 (N_5460,N_4641,N_4673);
and U5461 (N_5461,N_4989,N_4716);
or U5462 (N_5462,N_4997,N_4924);
and U5463 (N_5463,N_4751,N_4935);
and U5464 (N_5464,N_4525,N_4857);
and U5465 (N_5465,N_4677,N_4514);
and U5466 (N_5466,N_4511,N_4703);
and U5467 (N_5467,N_4759,N_4645);
nor U5468 (N_5468,N_4968,N_4687);
or U5469 (N_5469,N_4967,N_4696);
and U5470 (N_5470,N_4553,N_4981);
and U5471 (N_5471,N_4687,N_4922);
and U5472 (N_5472,N_4652,N_4808);
nand U5473 (N_5473,N_4597,N_4744);
nand U5474 (N_5474,N_4851,N_4503);
nor U5475 (N_5475,N_4514,N_4581);
and U5476 (N_5476,N_4571,N_4867);
nand U5477 (N_5477,N_4867,N_4549);
nand U5478 (N_5478,N_4757,N_4754);
nand U5479 (N_5479,N_4915,N_4826);
or U5480 (N_5480,N_4712,N_4670);
nand U5481 (N_5481,N_4833,N_4684);
nor U5482 (N_5482,N_4643,N_4503);
nand U5483 (N_5483,N_4772,N_4912);
nor U5484 (N_5484,N_4940,N_4986);
xnor U5485 (N_5485,N_4820,N_4884);
nor U5486 (N_5486,N_4532,N_4747);
and U5487 (N_5487,N_4730,N_4547);
nor U5488 (N_5488,N_4562,N_4683);
nor U5489 (N_5489,N_4645,N_4836);
xor U5490 (N_5490,N_4730,N_4605);
nor U5491 (N_5491,N_4582,N_4555);
xnor U5492 (N_5492,N_4895,N_4992);
or U5493 (N_5493,N_4912,N_4684);
nor U5494 (N_5494,N_4877,N_4680);
xor U5495 (N_5495,N_4662,N_4792);
or U5496 (N_5496,N_4562,N_4667);
xnor U5497 (N_5497,N_4901,N_4505);
nor U5498 (N_5498,N_4643,N_4856);
xor U5499 (N_5499,N_4997,N_4646);
or U5500 (N_5500,N_5381,N_5037);
xor U5501 (N_5501,N_5483,N_5262);
xnor U5502 (N_5502,N_5428,N_5411);
or U5503 (N_5503,N_5215,N_5047);
or U5504 (N_5504,N_5020,N_5118);
or U5505 (N_5505,N_5424,N_5252);
or U5506 (N_5506,N_5277,N_5299);
nand U5507 (N_5507,N_5150,N_5358);
xor U5508 (N_5508,N_5220,N_5468);
or U5509 (N_5509,N_5155,N_5340);
nand U5510 (N_5510,N_5316,N_5264);
nor U5511 (N_5511,N_5269,N_5218);
xor U5512 (N_5512,N_5464,N_5423);
xor U5513 (N_5513,N_5078,N_5009);
nor U5514 (N_5514,N_5170,N_5221);
or U5515 (N_5515,N_5034,N_5489);
nor U5516 (N_5516,N_5117,N_5274);
xor U5517 (N_5517,N_5330,N_5430);
xnor U5518 (N_5518,N_5388,N_5088);
xnor U5519 (N_5519,N_5103,N_5421);
nand U5520 (N_5520,N_5311,N_5223);
or U5521 (N_5521,N_5392,N_5314);
or U5522 (N_5522,N_5279,N_5045);
and U5523 (N_5523,N_5325,N_5359);
nand U5524 (N_5524,N_5287,N_5005);
nor U5525 (N_5525,N_5444,N_5120);
nor U5526 (N_5526,N_5497,N_5235);
and U5527 (N_5527,N_5028,N_5452);
and U5528 (N_5528,N_5237,N_5227);
and U5529 (N_5529,N_5380,N_5039);
nor U5530 (N_5530,N_5082,N_5003);
or U5531 (N_5531,N_5178,N_5365);
and U5532 (N_5532,N_5337,N_5455);
nand U5533 (N_5533,N_5249,N_5168);
nor U5534 (N_5534,N_5152,N_5159);
nor U5535 (N_5535,N_5203,N_5070);
and U5536 (N_5536,N_5280,N_5375);
nor U5537 (N_5537,N_5270,N_5266);
nand U5538 (N_5538,N_5023,N_5393);
or U5539 (N_5539,N_5133,N_5377);
nand U5540 (N_5540,N_5156,N_5494);
or U5541 (N_5541,N_5238,N_5313);
nor U5542 (N_5542,N_5487,N_5473);
nand U5543 (N_5543,N_5233,N_5333);
nand U5544 (N_5544,N_5298,N_5477);
nor U5545 (N_5545,N_5355,N_5304);
nand U5546 (N_5546,N_5026,N_5171);
xor U5547 (N_5547,N_5437,N_5255);
and U5548 (N_5548,N_5211,N_5032);
and U5549 (N_5549,N_5465,N_5053);
nand U5550 (N_5550,N_5343,N_5177);
nor U5551 (N_5551,N_5008,N_5285);
xnor U5552 (N_5552,N_5107,N_5236);
nand U5553 (N_5553,N_5100,N_5334);
xor U5554 (N_5554,N_5471,N_5167);
nand U5555 (N_5555,N_5129,N_5414);
nor U5556 (N_5556,N_5385,N_5109);
and U5557 (N_5557,N_5401,N_5260);
nand U5558 (N_5558,N_5014,N_5391);
nand U5559 (N_5559,N_5172,N_5176);
xor U5560 (N_5560,N_5484,N_5022);
nor U5561 (N_5561,N_5289,N_5089);
xor U5562 (N_5562,N_5163,N_5371);
nor U5563 (N_5563,N_5482,N_5180);
and U5564 (N_5564,N_5449,N_5426);
or U5565 (N_5565,N_5186,N_5126);
nor U5566 (N_5566,N_5033,N_5329);
xnor U5567 (N_5567,N_5383,N_5087);
nor U5568 (N_5568,N_5438,N_5281);
or U5569 (N_5569,N_5164,N_5190);
nor U5570 (N_5570,N_5348,N_5035);
xor U5571 (N_5571,N_5001,N_5065);
or U5572 (N_5572,N_5386,N_5000);
xor U5573 (N_5573,N_5241,N_5323);
nand U5574 (N_5574,N_5369,N_5104);
or U5575 (N_5575,N_5301,N_5019);
or U5576 (N_5576,N_5072,N_5145);
xor U5577 (N_5577,N_5043,N_5328);
nand U5578 (N_5578,N_5091,N_5004);
or U5579 (N_5579,N_5011,N_5206);
nor U5580 (N_5580,N_5195,N_5353);
nand U5581 (N_5581,N_5283,N_5114);
and U5582 (N_5582,N_5061,N_5239);
or U5583 (N_5583,N_5336,N_5467);
nand U5584 (N_5584,N_5404,N_5111);
xnor U5585 (N_5585,N_5193,N_5453);
xor U5586 (N_5586,N_5422,N_5276);
xor U5587 (N_5587,N_5040,N_5138);
nand U5588 (N_5588,N_5419,N_5250);
nand U5589 (N_5589,N_5122,N_5116);
or U5590 (N_5590,N_5083,N_5013);
or U5591 (N_5591,N_5185,N_5029);
or U5592 (N_5592,N_5320,N_5051);
or U5593 (N_5593,N_5098,N_5036);
or U5594 (N_5594,N_5044,N_5134);
nand U5595 (N_5595,N_5272,N_5125);
nand U5596 (N_5596,N_5224,N_5364);
and U5597 (N_5597,N_5041,N_5303);
xor U5598 (N_5598,N_5253,N_5189);
xnor U5599 (N_5599,N_5286,N_5413);
nand U5600 (N_5600,N_5317,N_5427);
nor U5601 (N_5601,N_5173,N_5376);
and U5602 (N_5602,N_5174,N_5480);
nand U5603 (N_5603,N_5291,N_5209);
nor U5604 (N_5604,N_5310,N_5350);
or U5605 (N_5605,N_5228,N_5254);
and U5606 (N_5606,N_5148,N_5459);
and U5607 (N_5607,N_5093,N_5433);
or U5608 (N_5608,N_5259,N_5461);
or U5609 (N_5609,N_5256,N_5092);
and U5610 (N_5610,N_5055,N_5208);
nand U5611 (N_5611,N_5410,N_5481);
nand U5612 (N_5612,N_5207,N_5321);
nand U5613 (N_5613,N_5293,N_5384);
and U5614 (N_5614,N_5042,N_5360);
or U5615 (N_5615,N_5157,N_5394);
and U5616 (N_5616,N_5076,N_5132);
or U5617 (N_5617,N_5431,N_5031);
nand U5618 (N_5618,N_5346,N_5408);
and U5619 (N_5619,N_5101,N_5294);
or U5620 (N_5620,N_5382,N_5341);
and U5621 (N_5621,N_5389,N_5099);
nand U5622 (N_5622,N_5282,N_5425);
nor U5623 (N_5623,N_5131,N_5135);
and U5624 (N_5624,N_5257,N_5488);
and U5625 (N_5625,N_5158,N_5447);
nand U5626 (N_5626,N_5142,N_5307);
nand U5627 (N_5627,N_5012,N_5069);
or U5628 (N_5628,N_5338,N_5048);
or U5629 (N_5629,N_5054,N_5248);
nand U5630 (N_5630,N_5149,N_5309);
and U5631 (N_5631,N_5354,N_5418);
nor U5632 (N_5632,N_5015,N_5296);
xnor U5633 (N_5633,N_5137,N_5006);
nor U5634 (N_5634,N_5344,N_5457);
nand U5635 (N_5635,N_5327,N_5077);
nor U5636 (N_5636,N_5278,N_5197);
or U5637 (N_5637,N_5024,N_5067);
or U5638 (N_5638,N_5486,N_5368);
and U5639 (N_5639,N_5205,N_5139);
xnor U5640 (N_5640,N_5146,N_5182);
and U5641 (N_5641,N_5324,N_5361);
or U5642 (N_5642,N_5094,N_5016);
nand U5643 (N_5643,N_5308,N_5458);
and U5644 (N_5644,N_5038,N_5219);
nand U5645 (N_5645,N_5493,N_5181);
or U5646 (N_5646,N_5201,N_5108);
xor U5647 (N_5647,N_5415,N_5027);
nand U5648 (N_5648,N_5372,N_5002);
and U5649 (N_5649,N_5470,N_5096);
nor U5650 (N_5650,N_5443,N_5086);
nor U5651 (N_5651,N_5339,N_5058);
or U5652 (N_5652,N_5400,N_5492);
nand U5653 (N_5653,N_5121,N_5153);
or U5654 (N_5654,N_5062,N_5448);
xor U5655 (N_5655,N_5275,N_5243);
xnor U5656 (N_5656,N_5018,N_5284);
or U5657 (N_5657,N_5007,N_5200);
or U5658 (N_5658,N_5362,N_5246);
and U5659 (N_5659,N_5356,N_5349);
xor U5660 (N_5660,N_5297,N_5064);
xor U5661 (N_5661,N_5115,N_5268);
and U5662 (N_5662,N_5345,N_5475);
and U5663 (N_5663,N_5210,N_5409);
nand U5664 (N_5664,N_5143,N_5436);
nand U5665 (N_5665,N_5151,N_5073);
nor U5666 (N_5666,N_5021,N_5403);
and U5667 (N_5667,N_5119,N_5230);
nor U5668 (N_5668,N_5071,N_5102);
nand U5669 (N_5669,N_5095,N_5130);
nand U5670 (N_5670,N_5342,N_5194);
and U5671 (N_5671,N_5351,N_5198);
or U5672 (N_5672,N_5136,N_5397);
and U5673 (N_5673,N_5479,N_5335);
nor U5674 (N_5674,N_5216,N_5160);
and U5675 (N_5675,N_5416,N_5188);
xnor U5676 (N_5676,N_5440,N_5166);
or U5677 (N_5677,N_5030,N_5472);
nand U5678 (N_5678,N_5128,N_5331);
nand U5679 (N_5679,N_5288,N_5417);
or U5680 (N_5680,N_5312,N_5175);
nand U5681 (N_5681,N_5105,N_5196);
nand U5682 (N_5682,N_5315,N_5217);
xor U5683 (N_5683,N_5068,N_5097);
or U5684 (N_5684,N_5367,N_5106);
nor U5685 (N_5685,N_5242,N_5454);
or U5686 (N_5686,N_5295,N_5485);
nand U5687 (N_5687,N_5399,N_5231);
nor U5688 (N_5688,N_5451,N_5474);
xnor U5689 (N_5689,N_5169,N_5052);
nor U5690 (N_5690,N_5084,N_5056);
nand U5691 (N_5691,N_5491,N_5466);
xnor U5692 (N_5692,N_5214,N_5124);
nand U5693 (N_5693,N_5407,N_5441);
nand U5694 (N_5694,N_5445,N_5081);
nor U5695 (N_5695,N_5010,N_5460);
and U5696 (N_5696,N_5165,N_5113);
nor U5697 (N_5697,N_5267,N_5478);
nand U5698 (N_5698,N_5232,N_5378);
or U5699 (N_5699,N_5059,N_5302);
xor U5700 (N_5700,N_5370,N_5322);
nand U5701 (N_5701,N_5495,N_5379);
and U5702 (N_5702,N_5050,N_5412);
xnor U5703 (N_5703,N_5373,N_5347);
nand U5704 (N_5704,N_5429,N_5463);
xor U5705 (N_5705,N_5057,N_5390);
xor U5706 (N_5706,N_5366,N_5420);
xor U5707 (N_5707,N_5202,N_5079);
xnor U5708 (N_5708,N_5374,N_5306);
and U5709 (N_5709,N_5352,N_5187);
or U5710 (N_5710,N_5183,N_5046);
and U5711 (N_5711,N_5439,N_5405);
nor U5712 (N_5712,N_5462,N_5063);
nand U5713 (N_5713,N_5066,N_5363);
nand U5714 (N_5714,N_5127,N_5387);
nand U5715 (N_5715,N_5199,N_5442);
nor U5716 (N_5716,N_5212,N_5247);
xnor U5717 (N_5717,N_5222,N_5395);
and U5718 (N_5718,N_5225,N_5496);
or U5719 (N_5719,N_5112,N_5318);
nor U5720 (N_5720,N_5476,N_5326);
and U5721 (N_5721,N_5080,N_5123);
nand U5722 (N_5722,N_5271,N_5258);
nor U5723 (N_5723,N_5292,N_5406);
and U5724 (N_5724,N_5456,N_5147);
nand U5725 (N_5725,N_5110,N_5085);
xnor U5726 (N_5726,N_5162,N_5263);
nor U5727 (N_5727,N_5244,N_5499);
xnor U5728 (N_5728,N_5261,N_5245);
and U5729 (N_5729,N_5179,N_5319);
nand U5730 (N_5730,N_5191,N_5075);
nand U5731 (N_5731,N_5434,N_5300);
and U5732 (N_5732,N_5161,N_5490);
nor U5733 (N_5733,N_5396,N_5357);
nor U5734 (N_5734,N_5265,N_5435);
xor U5735 (N_5735,N_5273,N_5213);
nor U5736 (N_5736,N_5140,N_5498);
nand U5737 (N_5737,N_5049,N_5240);
and U5738 (N_5738,N_5251,N_5446);
and U5739 (N_5739,N_5305,N_5234);
xor U5740 (N_5740,N_5432,N_5204);
or U5741 (N_5741,N_5154,N_5469);
nor U5742 (N_5742,N_5450,N_5090);
and U5743 (N_5743,N_5192,N_5332);
nor U5744 (N_5744,N_5226,N_5141);
xor U5745 (N_5745,N_5184,N_5402);
nand U5746 (N_5746,N_5074,N_5144);
or U5747 (N_5747,N_5060,N_5398);
nor U5748 (N_5748,N_5025,N_5290);
or U5749 (N_5749,N_5229,N_5017);
nand U5750 (N_5750,N_5340,N_5388);
or U5751 (N_5751,N_5411,N_5062);
nor U5752 (N_5752,N_5188,N_5385);
nor U5753 (N_5753,N_5387,N_5252);
nand U5754 (N_5754,N_5258,N_5191);
and U5755 (N_5755,N_5233,N_5259);
nand U5756 (N_5756,N_5184,N_5354);
and U5757 (N_5757,N_5376,N_5433);
xor U5758 (N_5758,N_5485,N_5361);
nor U5759 (N_5759,N_5414,N_5080);
or U5760 (N_5760,N_5422,N_5310);
and U5761 (N_5761,N_5398,N_5039);
and U5762 (N_5762,N_5348,N_5253);
xnor U5763 (N_5763,N_5180,N_5434);
or U5764 (N_5764,N_5274,N_5053);
nor U5765 (N_5765,N_5340,N_5017);
xnor U5766 (N_5766,N_5117,N_5168);
and U5767 (N_5767,N_5268,N_5380);
nand U5768 (N_5768,N_5045,N_5427);
nor U5769 (N_5769,N_5003,N_5147);
xor U5770 (N_5770,N_5323,N_5350);
nand U5771 (N_5771,N_5336,N_5127);
xnor U5772 (N_5772,N_5146,N_5213);
and U5773 (N_5773,N_5404,N_5182);
and U5774 (N_5774,N_5058,N_5049);
or U5775 (N_5775,N_5122,N_5283);
nor U5776 (N_5776,N_5440,N_5165);
xnor U5777 (N_5777,N_5054,N_5245);
nand U5778 (N_5778,N_5057,N_5191);
or U5779 (N_5779,N_5029,N_5303);
or U5780 (N_5780,N_5132,N_5051);
or U5781 (N_5781,N_5482,N_5398);
and U5782 (N_5782,N_5393,N_5346);
xor U5783 (N_5783,N_5080,N_5109);
xor U5784 (N_5784,N_5273,N_5436);
and U5785 (N_5785,N_5459,N_5089);
nand U5786 (N_5786,N_5256,N_5099);
nand U5787 (N_5787,N_5480,N_5285);
and U5788 (N_5788,N_5055,N_5251);
or U5789 (N_5789,N_5386,N_5443);
or U5790 (N_5790,N_5006,N_5147);
xnor U5791 (N_5791,N_5004,N_5348);
and U5792 (N_5792,N_5471,N_5161);
or U5793 (N_5793,N_5200,N_5002);
and U5794 (N_5794,N_5031,N_5333);
or U5795 (N_5795,N_5217,N_5153);
nor U5796 (N_5796,N_5029,N_5320);
nor U5797 (N_5797,N_5357,N_5341);
nand U5798 (N_5798,N_5236,N_5128);
xnor U5799 (N_5799,N_5066,N_5406);
xor U5800 (N_5800,N_5199,N_5464);
nor U5801 (N_5801,N_5309,N_5460);
nand U5802 (N_5802,N_5198,N_5297);
nand U5803 (N_5803,N_5222,N_5475);
nand U5804 (N_5804,N_5382,N_5296);
nand U5805 (N_5805,N_5145,N_5006);
and U5806 (N_5806,N_5153,N_5262);
or U5807 (N_5807,N_5010,N_5166);
and U5808 (N_5808,N_5231,N_5274);
xor U5809 (N_5809,N_5420,N_5139);
nand U5810 (N_5810,N_5142,N_5156);
xor U5811 (N_5811,N_5371,N_5420);
nor U5812 (N_5812,N_5034,N_5411);
nor U5813 (N_5813,N_5067,N_5193);
and U5814 (N_5814,N_5375,N_5479);
xnor U5815 (N_5815,N_5453,N_5305);
nor U5816 (N_5816,N_5423,N_5188);
nand U5817 (N_5817,N_5267,N_5395);
and U5818 (N_5818,N_5308,N_5276);
or U5819 (N_5819,N_5183,N_5267);
or U5820 (N_5820,N_5354,N_5369);
xnor U5821 (N_5821,N_5345,N_5498);
and U5822 (N_5822,N_5207,N_5214);
nand U5823 (N_5823,N_5008,N_5026);
and U5824 (N_5824,N_5485,N_5062);
xnor U5825 (N_5825,N_5178,N_5064);
nor U5826 (N_5826,N_5352,N_5289);
xor U5827 (N_5827,N_5226,N_5308);
nor U5828 (N_5828,N_5233,N_5192);
and U5829 (N_5829,N_5036,N_5393);
nor U5830 (N_5830,N_5338,N_5042);
nor U5831 (N_5831,N_5413,N_5036);
nand U5832 (N_5832,N_5202,N_5150);
nor U5833 (N_5833,N_5025,N_5104);
and U5834 (N_5834,N_5355,N_5239);
xor U5835 (N_5835,N_5157,N_5196);
and U5836 (N_5836,N_5367,N_5060);
or U5837 (N_5837,N_5146,N_5492);
and U5838 (N_5838,N_5083,N_5407);
xnor U5839 (N_5839,N_5187,N_5190);
nor U5840 (N_5840,N_5259,N_5462);
or U5841 (N_5841,N_5013,N_5403);
or U5842 (N_5842,N_5180,N_5079);
xnor U5843 (N_5843,N_5262,N_5111);
and U5844 (N_5844,N_5363,N_5083);
nor U5845 (N_5845,N_5114,N_5358);
or U5846 (N_5846,N_5367,N_5370);
nor U5847 (N_5847,N_5301,N_5381);
xor U5848 (N_5848,N_5198,N_5257);
nor U5849 (N_5849,N_5343,N_5306);
or U5850 (N_5850,N_5055,N_5319);
or U5851 (N_5851,N_5351,N_5462);
nand U5852 (N_5852,N_5108,N_5072);
and U5853 (N_5853,N_5353,N_5286);
or U5854 (N_5854,N_5008,N_5103);
nor U5855 (N_5855,N_5256,N_5122);
nor U5856 (N_5856,N_5186,N_5063);
nor U5857 (N_5857,N_5224,N_5424);
nand U5858 (N_5858,N_5484,N_5386);
nor U5859 (N_5859,N_5377,N_5049);
or U5860 (N_5860,N_5411,N_5472);
nand U5861 (N_5861,N_5089,N_5469);
and U5862 (N_5862,N_5478,N_5292);
nor U5863 (N_5863,N_5002,N_5208);
or U5864 (N_5864,N_5010,N_5041);
or U5865 (N_5865,N_5157,N_5129);
or U5866 (N_5866,N_5215,N_5328);
nor U5867 (N_5867,N_5392,N_5093);
nor U5868 (N_5868,N_5167,N_5191);
nand U5869 (N_5869,N_5093,N_5414);
xor U5870 (N_5870,N_5215,N_5061);
nand U5871 (N_5871,N_5022,N_5219);
xor U5872 (N_5872,N_5233,N_5383);
or U5873 (N_5873,N_5197,N_5384);
or U5874 (N_5874,N_5485,N_5357);
xnor U5875 (N_5875,N_5403,N_5269);
nor U5876 (N_5876,N_5088,N_5402);
and U5877 (N_5877,N_5118,N_5126);
xnor U5878 (N_5878,N_5321,N_5162);
xnor U5879 (N_5879,N_5480,N_5191);
nor U5880 (N_5880,N_5472,N_5184);
nand U5881 (N_5881,N_5489,N_5107);
nor U5882 (N_5882,N_5469,N_5185);
or U5883 (N_5883,N_5236,N_5179);
and U5884 (N_5884,N_5099,N_5443);
nor U5885 (N_5885,N_5159,N_5156);
nand U5886 (N_5886,N_5082,N_5442);
and U5887 (N_5887,N_5232,N_5325);
nand U5888 (N_5888,N_5410,N_5344);
nor U5889 (N_5889,N_5185,N_5248);
xor U5890 (N_5890,N_5097,N_5378);
or U5891 (N_5891,N_5381,N_5126);
or U5892 (N_5892,N_5328,N_5394);
nand U5893 (N_5893,N_5453,N_5476);
nor U5894 (N_5894,N_5154,N_5189);
nor U5895 (N_5895,N_5216,N_5337);
nor U5896 (N_5896,N_5173,N_5478);
nor U5897 (N_5897,N_5269,N_5188);
and U5898 (N_5898,N_5153,N_5264);
nor U5899 (N_5899,N_5312,N_5282);
and U5900 (N_5900,N_5251,N_5440);
xnor U5901 (N_5901,N_5046,N_5467);
xnor U5902 (N_5902,N_5114,N_5461);
nand U5903 (N_5903,N_5211,N_5437);
nor U5904 (N_5904,N_5185,N_5425);
nor U5905 (N_5905,N_5377,N_5005);
nor U5906 (N_5906,N_5246,N_5447);
xnor U5907 (N_5907,N_5273,N_5298);
xnor U5908 (N_5908,N_5013,N_5350);
and U5909 (N_5909,N_5110,N_5159);
and U5910 (N_5910,N_5088,N_5134);
xor U5911 (N_5911,N_5334,N_5143);
or U5912 (N_5912,N_5461,N_5112);
nand U5913 (N_5913,N_5005,N_5353);
nor U5914 (N_5914,N_5117,N_5158);
nand U5915 (N_5915,N_5231,N_5372);
or U5916 (N_5916,N_5444,N_5159);
nor U5917 (N_5917,N_5134,N_5009);
nor U5918 (N_5918,N_5439,N_5085);
nand U5919 (N_5919,N_5239,N_5094);
nand U5920 (N_5920,N_5386,N_5411);
xnor U5921 (N_5921,N_5282,N_5172);
or U5922 (N_5922,N_5029,N_5327);
xnor U5923 (N_5923,N_5044,N_5080);
or U5924 (N_5924,N_5266,N_5228);
and U5925 (N_5925,N_5004,N_5324);
nor U5926 (N_5926,N_5010,N_5399);
xnor U5927 (N_5927,N_5230,N_5067);
nand U5928 (N_5928,N_5262,N_5043);
xor U5929 (N_5929,N_5204,N_5441);
nand U5930 (N_5930,N_5402,N_5375);
or U5931 (N_5931,N_5102,N_5203);
and U5932 (N_5932,N_5168,N_5392);
xor U5933 (N_5933,N_5226,N_5059);
nand U5934 (N_5934,N_5043,N_5332);
or U5935 (N_5935,N_5181,N_5283);
nand U5936 (N_5936,N_5112,N_5044);
or U5937 (N_5937,N_5351,N_5314);
nand U5938 (N_5938,N_5351,N_5105);
xnor U5939 (N_5939,N_5454,N_5275);
xnor U5940 (N_5940,N_5350,N_5330);
or U5941 (N_5941,N_5464,N_5269);
nand U5942 (N_5942,N_5030,N_5109);
nor U5943 (N_5943,N_5423,N_5119);
nand U5944 (N_5944,N_5102,N_5008);
nor U5945 (N_5945,N_5443,N_5080);
nand U5946 (N_5946,N_5255,N_5469);
xnor U5947 (N_5947,N_5234,N_5416);
nand U5948 (N_5948,N_5385,N_5133);
nor U5949 (N_5949,N_5120,N_5106);
and U5950 (N_5950,N_5494,N_5411);
or U5951 (N_5951,N_5027,N_5168);
nor U5952 (N_5952,N_5498,N_5252);
xnor U5953 (N_5953,N_5191,N_5312);
xor U5954 (N_5954,N_5454,N_5334);
xnor U5955 (N_5955,N_5134,N_5160);
and U5956 (N_5956,N_5163,N_5148);
and U5957 (N_5957,N_5275,N_5390);
xor U5958 (N_5958,N_5016,N_5118);
nand U5959 (N_5959,N_5238,N_5379);
nor U5960 (N_5960,N_5283,N_5091);
and U5961 (N_5961,N_5156,N_5215);
xnor U5962 (N_5962,N_5134,N_5414);
nand U5963 (N_5963,N_5312,N_5143);
nand U5964 (N_5964,N_5024,N_5213);
or U5965 (N_5965,N_5485,N_5134);
and U5966 (N_5966,N_5069,N_5497);
nand U5967 (N_5967,N_5152,N_5023);
and U5968 (N_5968,N_5188,N_5226);
or U5969 (N_5969,N_5447,N_5282);
or U5970 (N_5970,N_5285,N_5381);
xor U5971 (N_5971,N_5152,N_5456);
or U5972 (N_5972,N_5201,N_5024);
nand U5973 (N_5973,N_5414,N_5218);
nor U5974 (N_5974,N_5456,N_5448);
nand U5975 (N_5975,N_5007,N_5385);
or U5976 (N_5976,N_5456,N_5494);
nor U5977 (N_5977,N_5071,N_5197);
nand U5978 (N_5978,N_5329,N_5279);
xor U5979 (N_5979,N_5247,N_5289);
nor U5980 (N_5980,N_5442,N_5062);
xnor U5981 (N_5981,N_5304,N_5118);
xnor U5982 (N_5982,N_5011,N_5137);
nor U5983 (N_5983,N_5288,N_5448);
and U5984 (N_5984,N_5475,N_5160);
nor U5985 (N_5985,N_5334,N_5447);
nand U5986 (N_5986,N_5459,N_5242);
or U5987 (N_5987,N_5110,N_5223);
nand U5988 (N_5988,N_5238,N_5209);
and U5989 (N_5989,N_5149,N_5461);
xor U5990 (N_5990,N_5037,N_5142);
xnor U5991 (N_5991,N_5284,N_5274);
nor U5992 (N_5992,N_5433,N_5467);
nor U5993 (N_5993,N_5115,N_5086);
nand U5994 (N_5994,N_5282,N_5069);
and U5995 (N_5995,N_5198,N_5261);
xor U5996 (N_5996,N_5206,N_5102);
nand U5997 (N_5997,N_5060,N_5330);
nand U5998 (N_5998,N_5401,N_5495);
nor U5999 (N_5999,N_5102,N_5413);
nand U6000 (N_6000,N_5521,N_5957);
xor U6001 (N_6001,N_5599,N_5513);
or U6002 (N_6002,N_5978,N_5657);
xor U6003 (N_6003,N_5502,N_5701);
nand U6004 (N_6004,N_5645,N_5886);
nand U6005 (N_6005,N_5745,N_5563);
or U6006 (N_6006,N_5786,N_5698);
nor U6007 (N_6007,N_5555,N_5848);
and U6008 (N_6008,N_5649,N_5659);
nand U6009 (N_6009,N_5526,N_5836);
nand U6010 (N_6010,N_5717,N_5802);
xor U6011 (N_6011,N_5993,N_5816);
nor U6012 (N_6012,N_5708,N_5684);
nand U6013 (N_6013,N_5847,N_5895);
xnor U6014 (N_6014,N_5960,N_5784);
nor U6015 (N_6015,N_5742,N_5522);
nand U6016 (N_6016,N_5772,N_5743);
and U6017 (N_6017,N_5704,N_5729);
or U6018 (N_6018,N_5955,N_5686);
nor U6019 (N_6019,N_5589,N_5778);
or U6020 (N_6020,N_5905,N_5583);
or U6021 (N_6021,N_5682,N_5857);
nor U6022 (N_6022,N_5644,N_5953);
or U6023 (N_6023,N_5511,N_5741);
nor U6024 (N_6024,N_5576,N_5793);
and U6025 (N_6025,N_5790,N_5934);
nand U6026 (N_6026,N_5678,N_5537);
xnor U6027 (N_6027,N_5962,N_5918);
or U6028 (N_6028,N_5881,N_5766);
xor U6029 (N_6029,N_5952,N_5892);
nor U6030 (N_6030,N_5507,N_5618);
xor U6031 (N_6031,N_5610,N_5529);
nand U6032 (N_6032,N_5942,N_5725);
nor U6033 (N_6033,N_5959,N_5932);
nor U6034 (N_6034,N_5916,N_5887);
and U6035 (N_6035,N_5769,N_5607);
or U6036 (N_6036,N_5824,N_5780);
nand U6037 (N_6037,N_5876,N_5757);
or U6038 (N_6038,N_5530,N_5558);
nor U6039 (N_6039,N_5820,N_5969);
or U6040 (N_6040,N_5754,N_5667);
or U6041 (N_6041,N_5999,N_5949);
nand U6042 (N_6042,N_5984,N_5798);
nor U6043 (N_6043,N_5852,N_5861);
xnor U6044 (N_6044,N_5799,N_5570);
or U6045 (N_6045,N_5574,N_5773);
xnor U6046 (N_6046,N_5737,N_5501);
and U6047 (N_6047,N_5728,N_5992);
nor U6048 (N_6048,N_5747,N_5723);
or U6049 (N_6049,N_5720,N_5909);
nor U6050 (N_6050,N_5981,N_5781);
or U6051 (N_6051,N_5810,N_5750);
xor U6052 (N_6052,N_5765,N_5588);
nor U6053 (N_6053,N_5756,N_5967);
nor U6054 (N_6054,N_5715,N_5792);
nor U6055 (N_6055,N_5553,N_5691);
nor U6056 (N_6056,N_5807,N_5689);
and U6057 (N_6057,N_5907,N_5994);
nand U6058 (N_6058,N_5936,N_5722);
and U6059 (N_6059,N_5548,N_5998);
nor U6060 (N_6060,N_5544,N_5650);
nor U6061 (N_6061,N_5568,N_5956);
or U6062 (N_6062,N_5732,N_5523);
nor U6063 (N_6063,N_5894,N_5739);
nor U6064 (N_6064,N_5697,N_5731);
nand U6065 (N_6065,N_5559,N_5579);
or U6066 (N_6066,N_5573,N_5946);
and U6067 (N_6067,N_5621,N_5777);
and U6068 (N_6068,N_5623,N_5908);
or U6069 (N_6069,N_5768,N_5996);
or U6070 (N_6070,N_5629,N_5664);
and U6071 (N_6071,N_5995,N_5670);
and U6072 (N_6072,N_5878,N_5591);
nand U6073 (N_6073,N_5870,N_5867);
nand U6074 (N_6074,N_5580,N_5554);
and U6075 (N_6075,N_5520,N_5687);
xnor U6076 (N_6076,N_5590,N_5619);
nand U6077 (N_6077,N_5841,N_5843);
or U6078 (N_6078,N_5943,N_5904);
nor U6079 (N_6079,N_5945,N_5915);
nor U6080 (N_6080,N_5594,N_5617);
nor U6081 (N_6081,N_5801,N_5699);
and U6082 (N_6082,N_5740,N_5560);
and U6083 (N_6083,N_5791,N_5612);
and U6084 (N_6084,N_5823,N_5788);
or U6085 (N_6085,N_5517,N_5705);
nor U6086 (N_6086,N_5864,N_5817);
nor U6087 (N_6087,N_5724,N_5516);
or U6088 (N_6088,N_5855,N_5990);
nor U6089 (N_6089,N_5890,N_5826);
or U6090 (N_6090,N_5806,N_5979);
nand U6091 (N_6091,N_5928,N_5922);
nand U6092 (N_6092,N_5813,N_5811);
nand U6093 (N_6093,N_5730,N_5556);
nand U6094 (N_6094,N_5627,N_5504);
or U6095 (N_6095,N_5653,N_5693);
nor U6096 (N_6096,N_5666,N_5899);
and U6097 (N_6097,N_5850,N_5506);
nor U6098 (N_6098,N_5669,N_5938);
nor U6099 (N_6099,N_5885,N_5609);
nor U6100 (N_6100,N_5866,N_5608);
or U6101 (N_6101,N_5675,N_5789);
nor U6102 (N_6102,N_5726,N_5718);
or U6103 (N_6103,N_5571,N_5912);
or U6104 (N_6104,N_5825,N_5551);
or U6105 (N_6105,N_5891,N_5652);
and U6106 (N_6106,N_5510,N_5902);
nor U6107 (N_6107,N_5764,N_5628);
nand U6108 (N_6108,N_5771,N_5577);
and U6109 (N_6109,N_5803,N_5822);
xnor U6110 (N_6110,N_5707,N_5716);
or U6111 (N_6111,N_5661,N_5862);
or U6112 (N_6112,N_5988,N_5931);
nor U6113 (N_6113,N_5541,N_5989);
xnor U6114 (N_6114,N_5679,N_5869);
nor U6115 (N_6115,N_5635,N_5751);
xor U6116 (N_6116,N_5567,N_5838);
xor U6117 (N_6117,N_5547,N_5625);
xnor U6118 (N_6118,N_5896,N_5535);
nor U6119 (N_6119,N_5787,N_5688);
and U6120 (N_6120,N_5500,N_5566);
xnor U6121 (N_6121,N_5860,N_5971);
xor U6122 (N_6122,N_5968,N_5828);
nor U6123 (N_6123,N_5702,N_5776);
and U6124 (N_6124,N_5643,N_5681);
nor U6125 (N_6125,N_5703,N_5874);
nor U6126 (N_6126,N_5676,N_5927);
nand U6127 (N_6127,N_5897,N_5744);
xor U6128 (N_6128,N_5581,N_5797);
xor U6129 (N_6129,N_5545,N_5983);
nor U6130 (N_6130,N_5821,N_5602);
xnor U6131 (N_6131,N_5673,N_5569);
nor U6132 (N_6132,N_5964,N_5940);
xor U6133 (N_6133,N_5991,N_5846);
xor U6134 (N_6134,N_5626,N_5616);
or U6135 (N_6135,N_5795,N_5758);
nand U6136 (N_6136,N_5519,N_5719);
xnor U6137 (N_6137,N_5538,N_5770);
and U6138 (N_6138,N_5782,N_5671);
nor U6139 (N_6139,N_5598,N_5585);
and U6140 (N_6140,N_5593,N_5721);
or U6141 (N_6141,N_5898,N_5985);
or U6142 (N_6142,N_5525,N_5695);
nand U6143 (N_6143,N_5550,N_5534);
xnor U6144 (N_6144,N_5950,N_5763);
nand U6145 (N_6145,N_5575,N_5672);
and U6146 (N_6146,N_5884,N_5736);
and U6147 (N_6147,N_5840,N_5966);
or U6148 (N_6148,N_5651,N_5970);
xnor U6149 (N_6149,N_5913,N_5980);
or U6150 (N_6150,N_5900,N_5911);
or U6151 (N_6151,N_5982,N_5515);
or U6152 (N_6152,N_5965,N_5508);
and U6153 (N_6153,N_5595,N_5849);
and U6154 (N_6154,N_5925,N_5759);
xnor U6155 (N_6155,N_5646,N_5503);
or U6156 (N_6156,N_5963,N_5805);
nand U6157 (N_6157,N_5865,N_5856);
nand U6158 (N_6158,N_5549,N_5735);
or U6159 (N_6159,N_5562,N_5937);
nand U6160 (N_6160,N_5839,N_5713);
or U6161 (N_6161,N_5694,N_5976);
and U6162 (N_6162,N_5637,N_5712);
xnor U6163 (N_6163,N_5783,N_5604);
nand U6164 (N_6164,N_5578,N_5641);
nor U6165 (N_6165,N_5614,N_5597);
and U6166 (N_6166,N_5906,N_5640);
and U6167 (N_6167,N_5804,N_5620);
and U6168 (N_6168,N_5552,N_5714);
nand U6169 (N_6169,N_5833,N_5872);
nand U6170 (N_6170,N_5509,N_5648);
nor U6171 (N_6171,N_5622,N_5853);
xnor U6172 (N_6172,N_5903,N_5975);
and U6173 (N_6173,N_5746,N_5761);
xor U6174 (N_6174,N_5779,N_5829);
or U6175 (N_6175,N_5800,N_5926);
xnor U6176 (N_6176,N_5505,N_5873);
xnor U6177 (N_6177,N_5528,N_5524);
nor U6178 (N_6178,N_5532,N_5536);
nand U6179 (N_6179,N_5785,N_5518);
xnor U6180 (N_6180,N_5662,N_5924);
nor U6181 (N_6181,N_5920,N_5794);
nand U6182 (N_6182,N_5674,N_5706);
xnor U6183 (N_6183,N_5660,N_5951);
and U6184 (N_6184,N_5733,N_5947);
nor U6185 (N_6185,N_5748,N_5584);
nand U6186 (N_6186,N_5815,N_5592);
nor U6187 (N_6187,N_5539,N_5561);
nor U6188 (N_6188,N_5837,N_5775);
or U6189 (N_6189,N_5830,N_5889);
nand U6190 (N_6190,N_5546,N_5683);
or U6191 (N_6191,N_5812,N_5831);
and U6192 (N_6192,N_5647,N_5809);
nand U6193 (N_6193,N_5710,N_5600);
or U6194 (N_6194,N_5851,N_5677);
nand U6195 (N_6195,N_5808,N_5656);
and U6196 (N_6196,N_5727,N_5859);
and U6197 (N_6197,N_5533,N_5882);
nand U6198 (N_6198,N_5879,N_5929);
nor U6199 (N_6199,N_5734,N_5606);
nor U6200 (N_6200,N_5572,N_5910);
nor U6201 (N_6201,N_5961,N_5680);
or U6202 (N_6202,N_5753,N_5944);
and U6203 (N_6203,N_5512,N_5668);
xor U6204 (N_6204,N_5835,N_5973);
nor U6205 (N_6205,N_5917,N_5933);
and U6206 (N_6206,N_5954,N_5863);
xor U6207 (N_6207,N_5972,N_5930);
or U6208 (N_6208,N_5842,N_5540);
xnor U6209 (N_6209,N_5613,N_5711);
and U6210 (N_6210,N_5690,N_5948);
nor U6211 (N_6211,N_5615,N_5935);
nand U6212 (N_6212,N_5654,N_5919);
and U6213 (N_6213,N_5709,N_5639);
and U6214 (N_6214,N_5596,N_5767);
or U6215 (N_6215,N_5542,N_5752);
nand U6216 (N_6216,N_5760,N_5814);
nor U6217 (N_6217,N_5665,N_5663);
nand U6218 (N_6218,N_5543,N_5557);
or U6219 (N_6219,N_5755,N_5696);
nor U6220 (N_6220,N_5939,N_5692);
nor U6221 (N_6221,N_5997,N_5531);
and U6222 (N_6222,N_5834,N_5685);
xnor U6223 (N_6223,N_5700,N_5658);
and U6224 (N_6224,N_5774,N_5564);
xnor U6225 (N_6225,N_5601,N_5854);
or U6226 (N_6226,N_5636,N_5818);
nand U6227 (N_6227,N_5796,N_5941);
or U6228 (N_6228,N_5827,N_5868);
and U6229 (N_6229,N_5642,N_5749);
nor U6230 (N_6230,N_5611,N_5893);
xor U6231 (N_6231,N_5958,N_5587);
or U6232 (N_6232,N_5888,N_5514);
and U6233 (N_6233,N_5633,N_5858);
xor U6234 (N_6234,N_5527,N_5871);
nor U6235 (N_6235,N_5586,N_5914);
xnor U6236 (N_6236,N_5632,N_5921);
nor U6237 (N_6237,N_5565,N_5977);
nor U6238 (N_6238,N_5974,N_5762);
nand U6239 (N_6239,N_5638,N_5923);
nor U6240 (N_6240,N_5844,N_5832);
and U6241 (N_6241,N_5624,N_5631);
or U6242 (N_6242,N_5845,N_5634);
xnor U6243 (N_6243,N_5603,N_5875);
nor U6244 (N_6244,N_5883,N_5582);
xnor U6245 (N_6245,N_5630,N_5738);
and U6246 (N_6246,N_5880,N_5819);
and U6247 (N_6247,N_5655,N_5987);
or U6248 (N_6248,N_5901,N_5605);
nor U6249 (N_6249,N_5877,N_5986);
and U6250 (N_6250,N_5933,N_5867);
nor U6251 (N_6251,N_5983,N_5763);
and U6252 (N_6252,N_5892,N_5987);
xor U6253 (N_6253,N_5559,N_5850);
xnor U6254 (N_6254,N_5868,N_5629);
or U6255 (N_6255,N_5721,N_5538);
xor U6256 (N_6256,N_5910,N_5695);
or U6257 (N_6257,N_5997,N_5859);
nand U6258 (N_6258,N_5853,N_5621);
xnor U6259 (N_6259,N_5724,N_5785);
xnor U6260 (N_6260,N_5624,N_5676);
nor U6261 (N_6261,N_5835,N_5845);
or U6262 (N_6262,N_5924,N_5965);
nand U6263 (N_6263,N_5691,N_5922);
nor U6264 (N_6264,N_5959,N_5787);
nor U6265 (N_6265,N_5567,N_5585);
or U6266 (N_6266,N_5987,N_5821);
xor U6267 (N_6267,N_5657,N_5669);
nor U6268 (N_6268,N_5583,N_5666);
nor U6269 (N_6269,N_5885,N_5870);
or U6270 (N_6270,N_5870,N_5933);
and U6271 (N_6271,N_5729,N_5579);
nor U6272 (N_6272,N_5704,N_5998);
nand U6273 (N_6273,N_5763,N_5980);
and U6274 (N_6274,N_5729,N_5776);
nand U6275 (N_6275,N_5652,N_5768);
xor U6276 (N_6276,N_5674,N_5682);
xor U6277 (N_6277,N_5747,N_5665);
and U6278 (N_6278,N_5958,N_5832);
or U6279 (N_6279,N_5926,N_5921);
xnor U6280 (N_6280,N_5500,N_5585);
nand U6281 (N_6281,N_5736,N_5911);
nor U6282 (N_6282,N_5651,N_5584);
and U6283 (N_6283,N_5875,N_5796);
and U6284 (N_6284,N_5652,N_5539);
and U6285 (N_6285,N_5587,N_5976);
or U6286 (N_6286,N_5980,N_5762);
nand U6287 (N_6287,N_5983,N_5601);
xnor U6288 (N_6288,N_5541,N_5601);
or U6289 (N_6289,N_5612,N_5506);
nand U6290 (N_6290,N_5514,N_5781);
xor U6291 (N_6291,N_5695,N_5749);
nor U6292 (N_6292,N_5925,N_5635);
nor U6293 (N_6293,N_5695,N_5786);
xnor U6294 (N_6294,N_5821,N_5800);
nand U6295 (N_6295,N_5800,N_5773);
and U6296 (N_6296,N_5662,N_5586);
xor U6297 (N_6297,N_5799,N_5701);
or U6298 (N_6298,N_5567,N_5559);
or U6299 (N_6299,N_5761,N_5902);
or U6300 (N_6300,N_5645,N_5603);
xor U6301 (N_6301,N_5921,N_5552);
nand U6302 (N_6302,N_5805,N_5976);
and U6303 (N_6303,N_5657,N_5641);
nand U6304 (N_6304,N_5714,N_5697);
and U6305 (N_6305,N_5947,N_5868);
xor U6306 (N_6306,N_5719,N_5859);
nand U6307 (N_6307,N_5978,N_5831);
xor U6308 (N_6308,N_5624,N_5670);
nand U6309 (N_6309,N_5563,N_5773);
xor U6310 (N_6310,N_5543,N_5915);
or U6311 (N_6311,N_5571,N_5843);
or U6312 (N_6312,N_5594,N_5709);
and U6313 (N_6313,N_5740,N_5945);
and U6314 (N_6314,N_5500,N_5983);
and U6315 (N_6315,N_5526,N_5547);
nand U6316 (N_6316,N_5755,N_5975);
and U6317 (N_6317,N_5763,N_5907);
nor U6318 (N_6318,N_5518,N_5792);
or U6319 (N_6319,N_5580,N_5617);
or U6320 (N_6320,N_5843,N_5550);
or U6321 (N_6321,N_5785,N_5983);
or U6322 (N_6322,N_5615,N_5874);
and U6323 (N_6323,N_5510,N_5562);
nand U6324 (N_6324,N_5769,N_5636);
xor U6325 (N_6325,N_5968,N_5576);
or U6326 (N_6326,N_5796,N_5700);
nor U6327 (N_6327,N_5554,N_5822);
and U6328 (N_6328,N_5880,N_5754);
or U6329 (N_6329,N_5672,N_5728);
nand U6330 (N_6330,N_5511,N_5661);
nand U6331 (N_6331,N_5945,N_5602);
nor U6332 (N_6332,N_5925,N_5996);
and U6333 (N_6333,N_5819,N_5651);
and U6334 (N_6334,N_5737,N_5823);
and U6335 (N_6335,N_5879,N_5713);
or U6336 (N_6336,N_5682,N_5522);
and U6337 (N_6337,N_5575,N_5592);
nor U6338 (N_6338,N_5745,N_5910);
and U6339 (N_6339,N_5999,N_5763);
nor U6340 (N_6340,N_5635,N_5517);
nand U6341 (N_6341,N_5985,N_5831);
nor U6342 (N_6342,N_5817,N_5692);
nor U6343 (N_6343,N_5859,N_5823);
or U6344 (N_6344,N_5851,N_5639);
and U6345 (N_6345,N_5608,N_5695);
nor U6346 (N_6346,N_5737,N_5879);
nand U6347 (N_6347,N_5646,N_5987);
or U6348 (N_6348,N_5971,N_5930);
nor U6349 (N_6349,N_5629,N_5713);
xor U6350 (N_6350,N_5865,N_5965);
or U6351 (N_6351,N_5821,N_5581);
nand U6352 (N_6352,N_5900,N_5823);
or U6353 (N_6353,N_5614,N_5974);
nand U6354 (N_6354,N_5731,N_5859);
and U6355 (N_6355,N_5563,N_5823);
or U6356 (N_6356,N_5945,N_5906);
or U6357 (N_6357,N_5957,N_5925);
xnor U6358 (N_6358,N_5577,N_5966);
nor U6359 (N_6359,N_5670,N_5755);
nand U6360 (N_6360,N_5827,N_5972);
nor U6361 (N_6361,N_5510,N_5735);
or U6362 (N_6362,N_5849,N_5756);
and U6363 (N_6363,N_5929,N_5520);
nor U6364 (N_6364,N_5524,N_5616);
or U6365 (N_6365,N_5735,N_5636);
or U6366 (N_6366,N_5790,N_5565);
nand U6367 (N_6367,N_5956,N_5880);
nor U6368 (N_6368,N_5636,N_5974);
nand U6369 (N_6369,N_5624,N_5762);
nand U6370 (N_6370,N_5801,N_5696);
xor U6371 (N_6371,N_5567,N_5763);
or U6372 (N_6372,N_5652,N_5862);
and U6373 (N_6373,N_5833,N_5617);
and U6374 (N_6374,N_5671,N_5805);
and U6375 (N_6375,N_5522,N_5756);
nand U6376 (N_6376,N_5823,N_5664);
nand U6377 (N_6377,N_5526,N_5593);
nand U6378 (N_6378,N_5978,N_5957);
or U6379 (N_6379,N_5592,N_5627);
xor U6380 (N_6380,N_5943,N_5568);
and U6381 (N_6381,N_5508,N_5923);
or U6382 (N_6382,N_5722,N_5943);
xnor U6383 (N_6383,N_5806,N_5607);
nor U6384 (N_6384,N_5764,N_5955);
nand U6385 (N_6385,N_5764,N_5805);
nor U6386 (N_6386,N_5545,N_5719);
nor U6387 (N_6387,N_5745,N_5790);
or U6388 (N_6388,N_5892,N_5798);
nor U6389 (N_6389,N_5949,N_5991);
and U6390 (N_6390,N_5885,N_5977);
and U6391 (N_6391,N_5710,N_5695);
and U6392 (N_6392,N_5696,N_5908);
nor U6393 (N_6393,N_5826,N_5723);
or U6394 (N_6394,N_5846,N_5978);
or U6395 (N_6395,N_5758,N_5800);
and U6396 (N_6396,N_5947,N_5905);
nand U6397 (N_6397,N_5976,N_5972);
and U6398 (N_6398,N_5820,N_5779);
xor U6399 (N_6399,N_5944,N_5566);
and U6400 (N_6400,N_5838,N_5699);
and U6401 (N_6401,N_5817,N_5580);
and U6402 (N_6402,N_5717,N_5656);
and U6403 (N_6403,N_5574,N_5764);
xnor U6404 (N_6404,N_5572,N_5754);
xnor U6405 (N_6405,N_5698,N_5619);
nand U6406 (N_6406,N_5853,N_5663);
nand U6407 (N_6407,N_5905,N_5704);
or U6408 (N_6408,N_5943,N_5877);
xor U6409 (N_6409,N_5671,N_5601);
nand U6410 (N_6410,N_5533,N_5849);
nand U6411 (N_6411,N_5557,N_5704);
or U6412 (N_6412,N_5626,N_5941);
and U6413 (N_6413,N_5993,N_5745);
nor U6414 (N_6414,N_5562,N_5548);
or U6415 (N_6415,N_5697,N_5685);
xnor U6416 (N_6416,N_5671,N_5503);
xnor U6417 (N_6417,N_5553,N_5824);
and U6418 (N_6418,N_5580,N_5992);
nand U6419 (N_6419,N_5590,N_5681);
nor U6420 (N_6420,N_5802,N_5527);
nor U6421 (N_6421,N_5959,N_5539);
nand U6422 (N_6422,N_5610,N_5532);
or U6423 (N_6423,N_5829,N_5783);
xnor U6424 (N_6424,N_5705,N_5786);
nand U6425 (N_6425,N_5704,N_5709);
and U6426 (N_6426,N_5655,N_5703);
nor U6427 (N_6427,N_5952,N_5616);
nand U6428 (N_6428,N_5973,N_5593);
or U6429 (N_6429,N_5821,N_5950);
and U6430 (N_6430,N_5832,N_5634);
xnor U6431 (N_6431,N_5749,N_5675);
xnor U6432 (N_6432,N_5634,N_5510);
nor U6433 (N_6433,N_5663,N_5648);
nor U6434 (N_6434,N_5932,N_5986);
xnor U6435 (N_6435,N_5947,N_5862);
nand U6436 (N_6436,N_5861,N_5591);
nor U6437 (N_6437,N_5584,N_5980);
xor U6438 (N_6438,N_5505,N_5826);
or U6439 (N_6439,N_5557,N_5792);
nor U6440 (N_6440,N_5535,N_5704);
nor U6441 (N_6441,N_5735,N_5769);
xor U6442 (N_6442,N_5829,N_5541);
nor U6443 (N_6443,N_5945,N_5704);
nor U6444 (N_6444,N_5895,N_5707);
nand U6445 (N_6445,N_5703,N_5662);
and U6446 (N_6446,N_5684,N_5758);
or U6447 (N_6447,N_5604,N_5847);
nand U6448 (N_6448,N_5780,N_5684);
nor U6449 (N_6449,N_5740,N_5636);
nor U6450 (N_6450,N_5930,N_5987);
and U6451 (N_6451,N_5833,N_5822);
or U6452 (N_6452,N_5771,N_5760);
xor U6453 (N_6453,N_5792,N_5586);
nand U6454 (N_6454,N_5884,N_5947);
and U6455 (N_6455,N_5985,N_5649);
xor U6456 (N_6456,N_5868,N_5824);
or U6457 (N_6457,N_5601,N_5922);
nand U6458 (N_6458,N_5587,N_5642);
and U6459 (N_6459,N_5600,N_5933);
nor U6460 (N_6460,N_5732,N_5757);
nand U6461 (N_6461,N_5594,N_5710);
and U6462 (N_6462,N_5729,N_5746);
and U6463 (N_6463,N_5991,N_5772);
nor U6464 (N_6464,N_5777,N_5870);
or U6465 (N_6465,N_5764,N_5767);
xnor U6466 (N_6466,N_5960,N_5898);
nor U6467 (N_6467,N_5918,N_5532);
and U6468 (N_6468,N_5977,N_5748);
nor U6469 (N_6469,N_5870,N_5646);
and U6470 (N_6470,N_5523,N_5989);
nor U6471 (N_6471,N_5836,N_5625);
or U6472 (N_6472,N_5836,N_5849);
nand U6473 (N_6473,N_5674,N_5579);
nor U6474 (N_6474,N_5618,N_5604);
or U6475 (N_6475,N_5572,N_5825);
or U6476 (N_6476,N_5913,N_5725);
and U6477 (N_6477,N_5693,N_5798);
or U6478 (N_6478,N_5942,N_5825);
nand U6479 (N_6479,N_5854,N_5618);
nor U6480 (N_6480,N_5728,N_5739);
or U6481 (N_6481,N_5557,N_5955);
nand U6482 (N_6482,N_5993,N_5978);
nand U6483 (N_6483,N_5848,N_5831);
or U6484 (N_6484,N_5720,N_5953);
and U6485 (N_6485,N_5789,N_5659);
nor U6486 (N_6486,N_5942,N_5769);
nor U6487 (N_6487,N_5746,N_5850);
nand U6488 (N_6488,N_5868,N_5867);
nor U6489 (N_6489,N_5814,N_5798);
and U6490 (N_6490,N_5682,N_5971);
and U6491 (N_6491,N_5666,N_5682);
nand U6492 (N_6492,N_5743,N_5738);
xnor U6493 (N_6493,N_5637,N_5922);
xor U6494 (N_6494,N_5802,N_5701);
nand U6495 (N_6495,N_5538,N_5984);
and U6496 (N_6496,N_5677,N_5906);
nand U6497 (N_6497,N_5525,N_5865);
xnor U6498 (N_6498,N_5876,N_5660);
nor U6499 (N_6499,N_5750,N_5618);
xor U6500 (N_6500,N_6328,N_6359);
or U6501 (N_6501,N_6304,N_6310);
nor U6502 (N_6502,N_6248,N_6087);
nand U6503 (N_6503,N_6101,N_6277);
or U6504 (N_6504,N_6228,N_6287);
and U6505 (N_6505,N_6108,N_6435);
and U6506 (N_6506,N_6191,N_6021);
xnor U6507 (N_6507,N_6379,N_6195);
nand U6508 (N_6508,N_6452,N_6053);
or U6509 (N_6509,N_6352,N_6003);
or U6510 (N_6510,N_6010,N_6471);
nor U6511 (N_6511,N_6343,N_6148);
nor U6512 (N_6512,N_6281,N_6405);
nor U6513 (N_6513,N_6437,N_6472);
or U6514 (N_6514,N_6419,N_6460);
or U6515 (N_6515,N_6457,N_6229);
and U6516 (N_6516,N_6090,N_6263);
and U6517 (N_6517,N_6112,N_6387);
nand U6518 (N_6518,N_6200,N_6260);
or U6519 (N_6519,N_6430,N_6291);
nor U6520 (N_6520,N_6158,N_6015);
nand U6521 (N_6521,N_6062,N_6494);
nor U6522 (N_6522,N_6275,N_6209);
nor U6523 (N_6523,N_6089,N_6069);
xor U6524 (N_6524,N_6432,N_6177);
or U6525 (N_6525,N_6289,N_6383);
or U6526 (N_6526,N_6371,N_6088);
xnor U6527 (N_6527,N_6219,N_6412);
xor U6528 (N_6528,N_6315,N_6376);
and U6529 (N_6529,N_6034,N_6205);
and U6530 (N_6530,N_6011,N_6198);
nor U6531 (N_6531,N_6473,N_6042);
nand U6532 (N_6532,N_6001,N_6160);
and U6533 (N_6533,N_6331,N_6180);
nand U6534 (N_6534,N_6363,N_6243);
and U6535 (N_6535,N_6396,N_6490);
nand U6536 (N_6536,N_6082,N_6194);
xnor U6537 (N_6537,N_6240,N_6153);
xnor U6538 (N_6538,N_6215,N_6370);
or U6539 (N_6539,N_6360,N_6126);
or U6540 (N_6540,N_6325,N_6446);
or U6541 (N_6541,N_6161,N_6073);
and U6542 (N_6542,N_6369,N_6250);
or U6543 (N_6543,N_6211,N_6496);
xor U6544 (N_6544,N_6192,N_6280);
nand U6545 (N_6545,N_6463,N_6253);
xor U6546 (N_6546,N_6436,N_6057);
nand U6547 (N_6547,N_6348,N_6199);
or U6548 (N_6548,N_6407,N_6272);
xnor U6549 (N_6549,N_6155,N_6134);
and U6550 (N_6550,N_6074,N_6204);
and U6551 (N_6551,N_6400,N_6459);
nor U6552 (N_6552,N_6025,N_6080);
and U6553 (N_6553,N_6133,N_6347);
and U6554 (N_6554,N_6045,N_6314);
and U6555 (N_6555,N_6464,N_6488);
nor U6556 (N_6556,N_6138,N_6202);
nor U6557 (N_6557,N_6335,N_6079);
or U6558 (N_6558,N_6029,N_6351);
or U6559 (N_6559,N_6444,N_6023);
and U6560 (N_6560,N_6208,N_6367);
xor U6561 (N_6561,N_6416,N_6186);
xor U6562 (N_6562,N_6479,N_6125);
and U6563 (N_6563,N_6411,N_6004);
xor U6564 (N_6564,N_6068,N_6358);
and U6565 (N_6565,N_6095,N_6278);
nor U6566 (N_6566,N_6453,N_6041);
nor U6567 (N_6567,N_6420,N_6425);
and U6568 (N_6568,N_6308,N_6039);
nand U6569 (N_6569,N_6176,N_6413);
or U6570 (N_6570,N_6442,N_6454);
and U6571 (N_6571,N_6262,N_6267);
xnor U6572 (N_6572,N_6377,N_6316);
xor U6573 (N_6573,N_6391,N_6188);
or U6574 (N_6574,N_6334,N_6330);
xnor U6575 (N_6575,N_6285,N_6344);
xnor U6576 (N_6576,N_6338,N_6036);
or U6577 (N_6577,N_6382,N_6332);
and U6578 (N_6578,N_6486,N_6225);
nor U6579 (N_6579,N_6475,N_6336);
nor U6580 (N_6580,N_6051,N_6049);
xnor U6581 (N_6581,N_6439,N_6313);
and U6582 (N_6582,N_6178,N_6115);
xnor U6583 (N_6583,N_6426,N_6116);
nor U6584 (N_6584,N_6468,N_6164);
nor U6585 (N_6585,N_6124,N_6113);
or U6586 (N_6586,N_6165,N_6353);
xnor U6587 (N_6587,N_6384,N_6107);
xnor U6588 (N_6588,N_6491,N_6084);
nand U6589 (N_6589,N_6337,N_6206);
nand U6590 (N_6590,N_6072,N_6394);
nand U6591 (N_6591,N_6269,N_6233);
or U6592 (N_6592,N_6066,N_6499);
nand U6593 (N_6593,N_6480,N_6237);
or U6594 (N_6594,N_6128,N_6421);
nand U6595 (N_6595,N_6386,N_6127);
nand U6596 (N_6596,N_6103,N_6000);
xnor U6597 (N_6597,N_6060,N_6146);
and U6598 (N_6598,N_6427,N_6014);
nand U6599 (N_6599,N_6341,N_6255);
xnor U6600 (N_6600,N_6047,N_6329);
xnor U6601 (N_6601,N_6102,N_6147);
nor U6602 (N_6602,N_6461,N_6449);
xor U6603 (N_6603,N_6450,N_6410);
and U6604 (N_6604,N_6170,N_6027);
nor U6605 (N_6605,N_6122,N_6207);
nand U6606 (N_6606,N_6061,N_6302);
and U6607 (N_6607,N_6075,N_6136);
or U6608 (N_6608,N_6311,N_6462);
nand U6609 (N_6609,N_6284,N_6349);
xnor U6610 (N_6610,N_6213,N_6050);
or U6611 (N_6611,N_6117,N_6013);
and U6612 (N_6612,N_6143,N_6227);
and U6613 (N_6613,N_6409,N_6086);
xor U6614 (N_6614,N_6220,N_6100);
or U6615 (N_6615,N_6467,N_6094);
nand U6616 (N_6616,N_6171,N_6020);
nor U6617 (N_6617,N_6283,N_6048);
xor U6618 (N_6618,N_6231,N_6043);
xor U6619 (N_6619,N_6181,N_6381);
nand U6620 (N_6620,N_6234,N_6163);
or U6621 (N_6621,N_6466,N_6478);
xnor U6622 (N_6622,N_6266,N_6007);
nand U6623 (N_6623,N_6154,N_6241);
and U6624 (N_6624,N_6017,N_6168);
nor U6625 (N_6625,N_6299,N_6058);
nand U6626 (N_6626,N_6397,N_6390);
xnor U6627 (N_6627,N_6495,N_6238);
or U6628 (N_6628,N_6077,N_6368);
nand U6629 (N_6629,N_6149,N_6111);
nand U6630 (N_6630,N_6455,N_6012);
and U6631 (N_6631,N_6300,N_6135);
nand U6632 (N_6632,N_6270,N_6109);
nor U6633 (N_6633,N_6054,N_6433);
nand U6634 (N_6634,N_6070,N_6261);
xnor U6635 (N_6635,N_6055,N_6144);
xor U6636 (N_6636,N_6076,N_6242);
or U6637 (N_6637,N_6078,N_6414);
xnor U6638 (N_6638,N_6395,N_6422);
nand U6639 (N_6639,N_6301,N_6393);
nor U6640 (N_6640,N_6399,N_6424);
nand U6641 (N_6641,N_6320,N_6189);
xnor U6642 (N_6642,N_6440,N_6085);
or U6643 (N_6643,N_6037,N_6005);
xnor U6644 (N_6644,N_6448,N_6224);
xnor U6645 (N_6645,N_6326,N_6290);
nand U6646 (N_6646,N_6091,N_6221);
or U6647 (N_6647,N_6105,N_6477);
xor U6648 (N_6648,N_6481,N_6375);
nor U6649 (N_6649,N_6130,N_6465);
or U6650 (N_6650,N_6121,N_6245);
and U6651 (N_6651,N_6056,N_6096);
and U6652 (N_6652,N_6361,N_6032);
nand U6653 (N_6653,N_6374,N_6322);
nand U6654 (N_6654,N_6123,N_6190);
and U6655 (N_6655,N_6323,N_6031);
xor U6656 (N_6656,N_6276,N_6346);
or U6657 (N_6657,N_6418,N_6139);
or U6658 (N_6658,N_6286,N_6024);
nor U6659 (N_6659,N_6222,N_6497);
or U6660 (N_6660,N_6483,N_6309);
or U6661 (N_6661,N_6385,N_6474);
and U6662 (N_6662,N_6006,N_6244);
xnor U6663 (N_6663,N_6030,N_6182);
nand U6664 (N_6664,N_6265,N_6485);
nand U6665 (N_6665,N_6487,N_6451);
nor U6666 (N_6666,N_6114,N_6378);
nor U6667 (N_6667,N_6179,N_6493);
xor U6668 (N_6668,N_6099,N_6293);
nand U6669 (N_6669,N_6254,N_6119);
xor U6670 (N_6670,N_6110,N_6258);
and U6671 (N_6671,N_6438,N_6026);
xnor U6672 (N_6672,N_6141,N_6298);
nor U6673 (N_6673,N_6044,N_6246);
nor U6674 (N_6674,N_6256,N_6271);
and U6675 (N_6675,N_6307,N_6456);
xnor U6676 (N_6676,N_6132,N_6404);
or U6677 (N_6677,N_6447,N_6356);
nand U6678 (N_6678,N_6482,N_6216);
or U6679 (N_6679,N_6187,N_6193);
nor U6680 (N_6680,N_6357,N_6185);
or U6681 (N_6681,N_6097,N_6067);
xnor U6682 (N_6682,N_6212,N_6294);
or U6683 (N_6683,N_6431,N_6252);
and U6684 (N_6684,N_6040,N_6151);
nand U6685 (N_6685,N_6104,N_6305);
nand U6686 (N_6686,N_6098,N_6081);
or U6687 (N_6687,N_6035,N_6131);
and U6688 (N_6688,N_6365,N_6214);
nand U6689 (N_6689,N_6162,N_6340);
or U6690 (N_6690,N_6106,N_6366);
and U6691 (N_6691,N_6303,N_6273);
and U6692 (N_6692,N_6268,N_6288);
nand U6693 (N_6693,N_6470,N_6129);
and U6694 (N_6694,N_6247,N_6327);
or U6695 (N_6695,N_6434,N_6217);
xnor U6696 (N_6696,N_6052,N_6364);
nand U6697 (N_6697,N_6355,N_6150);
nor U6698 (N_6698,N_6443,N_6292);
nand U6699 (N_6699,N_6264,N_6373);
xnor U6700 (N_6700,N_6282,N_6321);
nor U6701 (N_6701,N_6428,N_6118);
nor U6702 (N_6702,N_6159,N_6235);
nand U6703 (N_6703,N_6295,N_6002);
xor U6704 (N_6704,N_6484,N_6092);
and U6705 (N_6705,N_6059,N_6372);
or U6706 (N_6706,N_6489,N_6259);
or U6707 (N_6707,N_6354,N_6333);
and U6708 (N_6708,N_6339,N_6389);
nor U6709 (N_6709,N_6423,N_6392);
or U6710 (N_6710,N_6184,N_6362);
and U6711 (N_6711,N_6140,N_6445);
and U6712 (N_6712,N_6174,N_6317);
xnor U6713 (N_6713,N_6152,N_6183);
nand U6714 (N_6714,N_6093,N_6019);
xor U6715 (N_6715,N_6458,N_6380);
or U6716 (N_6716,N_6306,N_6064);
or U6717 (N_6717,N_6145,N_6257);
xor U6718 (N_6718,N_6169,N_6028);
nand U6719 (N_6719,N_6166,N_6175);
nor U6720 (N_6720,N_6415,N_6249);
and U6721 (N_6721,N_6441,N_6312);
nand U6722 (N_6722,N_6398,N_6402);
and U6723 (N_6723,N_6230,N_6226);
and U6724 (N_6724,N_6251,N_6063);
and U6725 (N_6725,N_6236,N_6142);
xor U6726 (N_6726,N_6022,N_6469);
and U6727 (N_6727,N_6324,N_6196);
xnor U6728 (N_6728,N_6342,N_6046);
nor U6729 (N_6729,N_6388,N_6318);
xnor U6730 (N_6730,N_6476,N_6173);
and U6731 (N_6731,N_6232,N_6172);
and U6732 (N_6732,N_6018,N_6008);
nor U6733 (N_6733,N_6071,N_6345);
or U6734 (N_6734,N_6009,N_6137);
xnor U6735 (N_6735,N_6279,N_6296);
nor U6736 (N_6736,N_6429,N_6197);
nor U6737 (N_6737,N_6401,N_6417);
nor U6738 (N_6738,N_6218,N_6065);
xor U6739 (N_6739,N_6274,N_6408);
and U6740 (N_6740,N_6201,N_6016);
xnor U6741 (N_6741,N_6350,N_6223);
and U6742 (N_6742,N_6157,N_6297);
nand U6743 (N_6743,N_6033,N_6203);
nand U6744 (N_6744,N_6319,N_6120);
and U6745 (N_6745,N_6210,N_6239);
nor U6746 (N_6746,N_6156,N_6406);
and U6747 (N_6747,N_6498,N_6492);
xnor U6748 (N_6748,N_6083,N_6167);
xnor U6749 (N_6749,N_6038,N_6403);
nor U6750 (N_6750,N_6172,N_6372);
nand U6751 (N_6751,N_6286,N_6291);
nand U6752 (N_6752,N_6131,N_6386);
nor U6753 (N_6753,N_6066,N_6452);
xor U6754 (N_6754,N_6373,N_6191);
nand U6755 (N_6755,N_6426,N_6219);
nor U6756 (N_6756,N_6124,N_6233);
nor U6757 (N_6757,N_6400,N_6022);
or U6758 (N_6758,N_6443,N_6195);
nor U6759 (N_6759,N_6210,N_6394);
xor U6760 (N_6760,N_6198,N_6409);
nor U6761 (N_6761,N_6388,N_6349);
and U6762 (N_6762,N_6360,N_6450);
or U6763 (N_6763,N_6249,N_6014);
nand U6764 (N_6764,N_6406,N_6235);
or U6765 (N_6765,N_6320,N_6491);
and U6766 (N_6766,N_6221,N_6140);
or U6767 (N_6767,N_6119,N_6465);
and U6768 (N_6768,N_6425,N_6453);
xor U6769 (N_6769,N_6366,N_6212);
xor U6770 (N_6770,N_6010,N_6027);
and U6771 (N_6771,N_6494,N_6370);
or U6772 (N_6772,N_6115,N_6424);
and U6773 (N_6773,N_6389,N_6085);
nand U6774 (N_6774,N_6397,N_6307);
xor U6775 (N_6775,N_6441,N_6018);
xor U6776 (N_6776,N_6353,N_6326);
and U6777 (N_6777,N_6304,N_6484);
xnor U6778 (N_6778,N_6233,N_6034);
or U6779 (N_6779,N_6037,N_6186);
or U6780 (N_6780,N_6156,N_6355);
xor U6781 (N_6781,N_6001,N_6205);
and U6782 (N_6782,N_6273,N_6250);
nor U6783 (N_6783,N_6119,N_6134);
xor U6784 (N_6784,N_6460,N_6228);
and U6785 (N_6785,N_6023,N_6406);
or U6786 (N_6786,N_6368,N_6396);
xor U6787 (N_6787,N_6052,N_6155);
nand U6788 (N_6788,N_6295,N_6119);
or U6789 (N_6789,N_6105,N_6104);
xnor U6790 (N_6790,N_6483,N_6187);
and U6791 (N_6791,N_6302,N_6178);
nand U6792 (N_6792,N_6389,N_6466);
and U6793 (N_6793,N_6489,N_6215);
or U6794 (N_6794,N_6209,N_6036);
nand U6795 (N_6795,N_6378,N_6020);
nand U6796 (N_6796,N_6261,N_6212);
xnor U6797 (N_6797,N_6320,N_6362);
nor U6798 (N_6798,N_6066,N_6333);
and U6799 (N_6799,N_6460,N_6328);
nor U6800 (N_6800,N_6015,N_6296);
nor U6801 (N_6801,N_6274,N_6455);
or U6802 (N_6802,N_6193,N_6046);
or U6803 (N_6803,N_6173,N_6147);
nor U6804 (N_6804,N_6279,N_6320);
and U6805 (N_6805,N_6297,N_6351);
and U6806 (N_6806,N_6010,N_6456);
or U6807 (N_6807,N_6391,N_6221);
or U6808 (N_6808,N_6385,N_6215);
nand U6809 (N_6809,N_6025,N_6054);
and U6810 (N_6810,N_6293,N_6112);
or U6811 (N_6811,N_6392,N_6261);
nand U6812 (N_6812,N_6449,N_6423);
and U6813 (N_6813,N_6105,N_6180);
nand U6814 (N_6814,N_6333,N_6450);
nand U6815 (N_6815,N_6373,N_6443);
nand U6816 (N_6816,N_6135,N_6154);
and U6817 (N_6817,N_6140,N_6423);
and U6818 (N_6818,N_6398,N_6107);
nor U6819 (N_6819,N_6412,N_6095);
nor U6820 (N_6820,N_6265,N_6271);
nand U6821 (N_6821,N_6062,N_6124);
and U6822 (N_6822,N_6470,N_6188);
xor U6823 (N_6823,N_6438,N_6478);
nor U6824 (N_6824,N_6117,N_6459);
xnor U6825 (N_6825,N_6340,N_6193);
xor U6826 (N_6826,N_6482,N_6185);
xor U6827 (N_6827,N_6416,N_6443);
xor U6828 (N_6828,N_6418,N_6129);
and U6829 (N_6829,N_6038,N_6037);
or U6830 (N_6830,N_6391,N_6072);
nor U6831 (N_6831,N_6456,N_6385);
nand U6832 (N_6832,N_6296,N_6413);
and U6833 (N_6833,N_6298,N_6232);
nor U6834 (N_6834,N_6109,N_6423);
xor U6835 (N_6835,N_6247,N_6191);
xnor U6836 (N_6836,N_6018,N_6110);
nand U6837 (N_6837,N_6044,N_6005);
or U6838 (N_6838,N_6339,N_6255);
nand U6839 (N_6839,N_6167,N_6196);
xnor U6840 (N_6840,N_6281,N_6475);
or U6841 (N_6841,N_6046,N_6024);
or U6842 (N_6842,N_6418,N_6363);
nor U6843 (N_6843,N_6244,N_6039);
or U6844 (N_6844,N_6048,N_6378);
or U6845 (N_6845,N_6354,N_6428);
nor U6846 (N_6846,N_6288,N_6050);
or U6847 (N_6847,N_6424,N_6164);
xor U6848 (N_6848,N_6109,N_6302);
nand U6849 (N_6849,N_6400,N_6350);
or U6850 (N_6850,N_6099,N_6301);
and U6851 (N_6851,N_6060,N_6028);
nor U6852 (N_6852,N_6058,N_6136);
or U6853 (N_6853,N_6313,N_6355);
nor U6854 (N_6854,N_6083,N_6368);
and U6855 (N_6855,N_6245,N_6170);
and U6856 (N_6856,N_6427,N_6045);
xnor U6857 (N_6857,N_6329,N_6006);
nand U6858 (N_6858,N_6358,N_6059);
and U6859 (N_6859,N_6415,N_6059);
xnor U6860 (N_6860,N_6288,N_6488);
and U6861 (N_6861,N_6132,N_6074);
xnor U6862 (N_6862,N_6295,N_6418);
xor U6863 (N_6863,N_6452,N_6332);
xnor U6864 (N_6864,N_6427,N_6329);
xor U6865 (N_6865,N_6091,N_6343);
nand U6866 (N_6866,N_6419,N_6454);
nor U6867 (N_6867,N_6128,N_6378);
and U6868 (N_6868,N_6165,N_6125);
nor U6869 (N_6869,N_6299,N_6292);
nand U6870 (N_6870,N_6223,N_6095);
or U6871 (N_6871,N_6339,N_6351);
xnor U6872 (N_6872,N_6283,N_6288);
nand U6873 (N_6873,N_6051,N_6174);
nand U6874 (N_6874,N_6148,N_6484);
and U6875 (N_6875,N_6113,N_6460);
nand U6876 (N_6876,N_6471,N_6273);
nand U6877 (N_6877,N_6152,N_6277);
or U6878 (N_6878,N_6389,N_6268);
and U6879 (N_6879,N_6245,N_6414);
and U6880 (N_6880,N_6082,N_6045);
or U6881 (N_6881,N_6293,N_6488);
nor U6882 (N_6882,N_6125,N_6109);
or U6883 (N_6883,N_6490,N_6480);
xnor U6884 (N_6884,N_6239,N_6271);
and U6885 (N_6885,N_6131,N_6451);
xnor U6886 (N_6886,N_6019,N_6436);
or U6887 (N_6887,N_6077,N_6415);
and U6888 (N_6888,N_6194,N_6395);
xor U6889 (N_6889,N_6112,N_6287);
or U6890 (N_6890,N_6495,N_6110);
nand U6891 (N_6891,N_6420,N_6016);
or U6892 (N_6892,N_6088,N_6232);
or U6893 (N_6893,N_6120,N_6424);
and U6894 (N_6894,N_6026,N_6016);
nor U6895 (N_6895,N_6451,N_6192);
xor U6896 (N_6896,N_6476,N_6379);
or U6897 (N_6897,N_6389,N_6341);
nor U6898 (N_6898,N_6245,N_6494);
and U6899 (N_6899,N_6387,N_6010);
nor U6900 (N_6900,N_6271,N_6224);
and U6901 (N_6901,N_6434,N_6271);
and U6902 (N_6902,N_6145,N_6429);
xor U6903 (N_6903,N_6287,N_6210);
nor U6904 (N_6904,N_6110,N_6071);
or U6905 (N_6905,N_6425,N_6095);
nor U6906 (N_6906,N_6461,N_6357);
or U6907 (N_6907,N_6139,N_6326);
nand U6908 (N_6908,N_6144,N_6328);
xnor U6909 (N_6909,N_6102,N_6338);
or U6910 (N_6910,N_6073,N_6335);
or U6911 (N_6911,N_6223,N_6481);
and U6912 (N_6912,N_6410,N_6326);
and U6913 (N_6913,N_6053,N_6100);
or U6914 (N_6914,N_6027,N_6317);
nor U6915 (N_6915,N_6491,N_6032);
xor U6916 (N_6916,N_6207,N_6250);
nand U6917 (N_6917,N_6227,N_6332);
nor U6918 (N_6918,N_6150,N_6263);
nand U6919 (N_6919,N_6393,N_6007);
nor U6920 (N_6920,N_6325,N_6416);
xnor U6921 (N_6921,N_6412,N_6443);
nand U6922 (N_6922,N_6426,N_6026);
or U6923 (N_6923,N_6498,N_6340);
nor U6924 (N_6924,N_6311,N_6492);
nor U6925 (N_6925,N_6285,N_6260);
or U6926 (N_6926,N_6187,N_6218);
or U6927 (N_6927,N_6257,N_6342);
nor U6928 (N_6928,N_6479,N_6071);
nor U6929 (N_6929,N_6103,N_6131);
xor U6930 (N_6930,N_6184,N_6172);
xnor U6931 (N_6931,N_6044,N_6477);
xor U6932 (N_6932,N_6238,N_6068);
nor U6933 (N_6933,N_6259,N_6045);
and U6934 (N_6934,N_6377,N_6453);
and U6935 (N_6935,N_6168,N_6185);
nand U6936 (N_6936,N_6202,N_6208);
nand U6937 (N_6937,N_6035,N_6275);
nand U6938 (N_6938,N_6328,N_6423);
xor U6939 (N_6939,N_6137,N_6266);
xnor U6940 (N_6940,N_6426,N_6059);
xnor U6941 (N_6941,N_6251,N_6130);
or U6942 (N_6942,N_6310,N_6049);
and U6943 (N_6943,N_6016,N_6005);
nand U6944 (N_6944,N_6283,N_6396);
xor U6945 (N_6945,N_6190,N_6201);
and U6946 (N_6946,N_6089,N_6426);
xnor U6947 (N_6947,N_6434,N_6242);
nand U6948 (N_6948,N_6111,N_6134);
nand U6949 (N_6949,N_6078,N_6328);
xnor U6950 (N_6950,N_6098,N_6261);
or U6951 (N_6951,N_6236,N_6421);
xnor U6952 (N_6952,N_6396,N_6176);
nor U6953 (N_6953,N_6220,N_6435);
nor U6954 (N_6954,N_6287,N_6169);
or U6955 (N_6955,N_6087,N_6081);
or U6956 (N_6956,N_6008,N_6039);
nand U6957 (N_6957,N_6247,N_6455);
and U6958 (N_6958,N_6396,N_6164);
nor U6959 (N_6959,N_6099,N_6238);
or U6960 (N_6960,N_6244,N_6078);
nor U6961 (N_6961,N_6300,N_6222);
xor U6962 (N_6962,N_6463,N_6395);
and U6963 (N_6963,N_6297,N_6024);
nand U6964 (N_6964,N_6135,N_6385);
nor U6965 (N_6965,N_6302,N_6198);
nor U6966 (N_6966,N_6090,N_6162);
nand U6967 (N_6967,N_6366,N_6125);
nand U6968 (N_6968,N_6026,N_6216);
nand U6969 (N_6969,N_6144,N_6455);
xor U6970 (N_6970,N_6339,N_6062);
nor U6971 (N_6971,N_6107,N_6009);
or U6972 (N_6972,N_6117,N_6466);
xor U6973 (N_6973,N_6051,N_6433);
or U6974 (N_6974,N_6165,N_6352);
nand U6975 (N_6975,N_6198,N_6258);
nand U6976 (N_6976,N_6488,N_6379);
and U6977 (N_6977,N_6397,N_6296);
nand U6978 (N_6978,N_6265,N_6181);
and U6979 (N_6979,N_6338,N_6434);
or U6980 (N_6980,N_6087,N_6214);
or U6981 (N_6981,N_6213,N_6170);
nor U6982 (N_6982,N_6401,N_6480);
and U6983 (N_6983,N_6148,N_6366);
nor U6984 (N_6984,N_6314,N_6129);
xnor U6985 (N_6985,N_6061,N_6250);
xor U6986 (N_6986,N_6132,N_6356);
or U6987 (N_6987,N_6023,N_6073);
xnor U6988 (N_6988,N_6062,N_6380);
and U6989 (N_6989,N_6066,N_6268);
nand U6990 (N_6990,N_6475,N_6414);
nand U6991 (N_6991,N_6136,N_6315);
or U6992 (N_6992,N_6195,N_6484);
nor U6993 (N_6993,N_6417,N_6062);
xnor U6994 (N_6994,N_6309,N_6321);
xor U6995 (N_6995,N_6319,N_6315);
nand U6996 (N_6996,N_6494,N_6331);
and U6997 (N_6997,N_6031,N_6499);
nand U6998 (N_6998,N_6393,N_6165);
nand U6999 (N_6999,N_6393,N_6326);
or U7000 (N_7000,N_6898,N_6882);
nand U7001 (N_7001,N_6773,N_6657);
or U7002 (N_7002,N_6905,N_6530);
xor U7003 (N_7003,N_6635,N_6965);
xor U7004 (N_7004,N_6973,N_6795);
xnor U7005 (N_7005,N_6528,N_6870);
nand U7006 (N_7006,N_6514,N_6536);
or U7007 (N_7007,N_6871,N_6763);
and U7008 (N_7008,N_6515,N_6727);
or U7009 (N_7009,N_6619,N_6847);
or U7010 (N_7010,N_6687,N_6896);
nor U7011 (N_7011,N_6943,N_6910);
and U7012 (N_7012,N_6862,N_6928);
or U7013 (N_7013,N_6764,N_6921);
nor U7014 (N_7014,N_6704,N_6962);
xor U7015 (N_7015,N_6684,N_6550);
and U7016 (N_7016,N_6799,N_6927);
nor U7017 (N_7017,N_6913,N_6641);
and U7018 (N_7018,N_6892,N_6855);
xnor U7019 (N_7019,N_6613,N_6809);
nor U7020 (N_7020,N_6994,N_6523);
xor U7021 (N_7021,N_6946,N_6680);
and U7022 (N_7022,N_6573,N_6769);
xnor U7023 (N_7023,N_6903,N_6574);
or U7024 (N_7024,N_6673,N_6540);
and U7025 (N_7025,N_6741,N_6825);
nand U7026 (N_7026,N_6777,N_6885);
or U7027 (N_7027,N_6527,N_6650);
nand U7028 (N_7028,N_6959,N_6575);
or U7029 (N_7029,N_6979,N_6719);
nand U7030 (N_7030,N_6744,N_6817);
or U7031 (N_7031,N_6854,N_6788);
nand U7032 (N_7032,N_6751,N_6629);
nor U7033 (N_7033,N_6797,N_6700);
and U7034 (N_7034,N_6645,N_6577);
and U7035 (N_7035,N_6889,N_6596);
nor U7036 (N_7036,N_6620,N_6766);
nand U7037 (N_7037,N_6975,N_6688);
nor U7038 (N_7038,N_6553,N_6549);
nand U7039 (N_7039,N_6647,N_6614);
or U7040 (N_7040,N_6877,N_6634);
and U7041 (N_7041,N_6728,N_6661);
xnor U7042 (N_7042,N_6695,N_6958);
xor U7043 (N_7043,N_6589,N_6754);
nor U7044 (N_7044,N_6960,N_6895);
or U7045 (N_7045,N_6838,N_6762);
and U7046 (N_7046,N_6945,N_6559);
nand U7047 (N_7047,N_6894,N_6667);
xnor U7048 (N_7048,N_6588,N_6904);
nor U7049 (N_7049,N_6792,N_6692);
nor U7050 (N_7050,N_6972,N_6623);
or U7051 (N_7051,N_6839,N_6907);
and U7052 (N_7052,N_6991,N_6806);
or U7053 (N_7053,N_6986,N_6500);
and U7054 (N_7054,N_6569,N_6571);
nand U7055 (N_7055,N_6622,N_6947);
xnor U7056 (N_7056,N_6966,N_6646);
xnor U7057 (N_7057,N_6701,N_6875);
or U7058 (N_7058,N_6917,N_6970);
xor U7059 (N_7059,N_6659,N_6807);
and U7060 (N_7060,N_6976,N_6558);
or U7061 (N_7061,N_6978,N_6794);
nor U7062 (N_7062,N_6757,N_6507);
nor U7063 (N_7063,N_6509,N_6756);
and U7064 (N_7064,N_6802,N_6971);
nor U7065 (N_7065,N_6936,N_6785);
or U7066 (N_7066,N_6720,N_6824);
xor U7067 (N_7067,N_6955,N_6772);
xnor U7068 (N_7068,N_6732,N_6781);
xnor U7069 (N_7069,N_6826,N_6513);
nand U7070 (N_7070,N_6901,N_6520);
xnor U7071 (N_7071,N_6526,N_6676);
and U7072 (N_7072,N_6504,N_6615);
nand U7073 (N_7073,N_6546,N_6501);
xor U7074 (N_7074,N_6678,N_6830);
nor U7075 (N_7075,N_6572,N_6967);
xor U7076 (N_7076,N_6551,N_6938);
or U7077 (N_7077,N_6812,N_6793);
xor U7078 (N_7078,N_6831,N_6633);
xnor U7079 (N_7079,N_6656,N_6786);
and U7080 (N_7080,N_6524,N_6611);
and U7081 (N_7081,N_6833,N_6929);
or U7082 (N_7082,N_6547,N_6803);
or U7083 (N_7083,N_6580,N_6605);
xnor U7084 (N_7084,N_6583,N_6787);
and U7085 (N_7085,N_6995,N_6798);
nand U7086 (N_7086,N_6518,N_6937);
nand U7087 (N_7087,N_6874,N_6853);
and U7088 (N_7088,N_6506,N_6996);
nor U7089 (N_7089,N_6887,N_6821);
nand U7090 (N_7090,N_6753,N_6662);
nor U7091 (N_7091,N_6861,N_6800);
xnor U7092 (N_7092,N_6872,N_6693);
and U7093 (N_7093,N_6568,N_6674);
nor U7094 (N_7094,N_6671,N_6934);
or U7095 (N_7095,N_6522,N_6923);
nor U7096 (N_7096,N_6775,N_6685);
and U7097 (N_7097,N_6768,N_6598);
nor U7098 (N_7098,N_6990,N_6748);
xor U7099 (N_7099,N_6819,N_6922);
xor U7100 (N_7100,N_6867,N_6840);
xor U7101 (N_7101,N_6624,N_6618);
xnor U7102 (N_7102,N_6660,N_6737);
and U7103 (N_7103,N_6760,N_6724);
nor U7104 (N_7104,N_6810,N_6627);
or U7105 (N_7105,N_6954,N_6691);
nor U7106 (N_7106,N_6651,N_6632);
or U7107 (N_7107,N_6968,N_6811);
and U7108 (N_7108,N_6866,N_6638);
nor U7109 (N_7109,N_6716,N_6796);
or U7110 (N_7110,N_6570,N_6998);
nor U7111 (N_7111,N_6999,N_6805);
or U7112 (N_7112,N_6576,N_6582);
xor U7113 (N_7113,N_6816,N_6900);
or U7114 (N_7114,N_6738,N_6743);
nand U7115 (N_7115,N_6560,N_6782);
xor U7116 (N_7116,N_6599,N_6808);
and U7117 (N_7117,N_6940,N_6916);
xor U7118 (N_7118,N_6525,N_6658);
xnor U7119 (N_7119,N_6718,N_6567);
or U7120 (N_7120,N_6595,N_6630);
xnor U7121 (N_7121,N_6606,N_6565);
nand U7122 (N_7122,N_6883,N_6869);
or U7123 (N_7123,N_6736,N_6859);
nand U7124 (N_7124,N_6908,N_6696);
and U7125 (N_7125,N_6594,N_6578);
xnor U7126 (N_7126,N_6851,N_6542);
and U7127 (N_7127,N_6920,N_6552);
nor U7128 (N_7128,N_6535,N_6914);
or U7129 (N_7129,N_6909,N_6829);
nor U7130 (N_7130,N_6699,N_6663);
nor U7131 (N_7131,N_6915,N_6873);
nand U7132 (N_7132,N_6987,N_6664);
nor U7133 (N_7133,N_6884,N_6841);
and U7134 (N_7134,N_6850,N_6814);
and U7135 (N_7135,N_6944,N_6818);
and U7136 (N_7136,N_6963,N_6607);
xnor U7137 (N_7137,N_6698,N_6617);
and U7138 (N_7138,N_6876,N_6858);
or U7139 (N_7139,N_6655,N_6783);
xor U7140 (N_7140,N_6856,N_6951);
nor U7141 (N_7141,N_6670,N_6765);
nand U7142 (N_7142,N_6933,N_6935);
and U7143 (N_7143,N_6621,N_6521);
and U7144 (N_7144,N_6988,N_6926);
or U7145 (N_7145,N_6554,N_6612);
nor U7146 (N_7146,N_6984,N_6608);
nand U7147 (N_7147,N_6591,N_6712);
nor U7148 (N_7148,N_6654,N_6845);
xnor U7149 (N_7149,N_6843,N_6779);
xor U7150 (N_7150,N_6677,N_6532);
and U7151 (N_7151,N_6745,N_6886);
xor U7152 (N_7152,N_6879,N_6561);
nor U7153 (N_7153,N_6564,N_6868);
nand U7154 (N_7154,N_6834,N_6503);
and U7155 (N_7155,N_6842,N_6666);
nand U7156 (N_7156,N_6616,N_6848);
nor U7157 (N_7157,N_6759,N_6771);
or U7158 (N_7158,N_6537,N_6725);
nand U7159 (N_7159,N_6610,N_6815);
or U7160 (N_7160,N_6849,N_6707);
nand U7161 (N_7161,N_6502,N_6556);
and U7162 (N_7162,N_6878,N_6804);
nand U7163 (N_7163,N_6733,N_6604);
nor U7164 (N_7164,N_6893,N_6631);
and U7165 (N_7165,N_6906,N_6888);
nand U7166 (N_7166,N_6541,N_6653);
xnor U7167 (N_7167,N_6689,N_6585);
nor U7168 (N_7168,N_6918,N_6822);
or U7169 (N_7169,N_6890,N_6717);
xor U7170 (N_7170,N_6711,N_6600);
xnor U7171 (N_7171,N_6985,N_6681);
nor U7172 (N_7172,N_6703,N_6665);
nand U7173 (N_7173,N_6731,N_6579);
nand U7174 (N_7174,N_6636,N_6705);
nand U7175 (N_7175,N_6669,N_6562);
xnor U7176 (N_7176,N_6702,N_6950);
nand U7177 (N_7177,N_6778,N_6519);
or U7178 (N_7178,N_6683,N_6713);
nand U7179 (N_7179,N_6602,N_6891);
nand U7180 (N_7180,N_6593,N_6863);
nand U7181 (N_7181,N_6740,N_6969);
and U7182 (N_7182,N_6776,N_6813);
or U7183 (N_7183,N_6828,N_6827);
and U7184 (N_7184,N_6880,N_6601);
or U7185 (N_7185,N_6708,N_6790);
and U7186 (N_7186,N_6739,N_6581);
nand U7187 (N_7187,N_6742,N_6747);
xnor U7188 (N_7188,N_6902,N_6952);
xnor U7189 (N_7189,N_6857,N_6586);
nand U7190 (N_7190,N_6544,N_6648);
or U7191 (N_7191,N_6981,N_6837);
xor U7192 (N_7192,N_6690,N_6836);
nor U7193 (N_7193,N_6864,N_6820);
nand U7194 (N_7194,N_6628,N_6977);
nand U7195 (N_7195,N_6956,N_6603);
nor U7196 (N_7196,N_6925,N_6548);
xor U7197 (N_7197,N_6592,N_6942);
nand U7198 (N_7198,N_6860,N_6730);
nand U7199 (N_7199,N_6539,N_6563);
or U7200 (N_7200,N_6697,N_6715);
and U7201 (N_7201,N_6721,N_6557);
or U7202 (N_7202,N_6625,N_6590);
or U7203 (N_7203,N_6957,N_6714);
nor U7204 (N_7204,N_6538,N_6801);
xnor U7205 (N_7205,N_6533,N_6749);
and U7206 (N_7206,N_6789,N_6982);
xnor U7207 (N_7207,N_6939,N_6980);
nor U7208 (N_7208,N_6897,N_6675);
and U7209 (N_7209,N_6770,N_6709);
and U7210 (N_7210,N_6780,N_6516);
and U7211 (N_7211,N_6668,N_6609);
nor U7212 (N_7212,N_6729,N_6752);
or U7213 (N_7213,N_6642,N_6640);
nand U7214 (N_7214,N_6997,N_6948);
nand U7215 (N_7215,N_6597,N_6746);
xnor U7216 (N_7216,N_6531,N_6924);
nand U7217 (N_7217,N_6512,N_6511);
or U7218 (N_7218,N_6881,N_6706);
xor U7219 (N_7219,N_6832,N_6761);
xor U7220 (N_7220,N_6791,N_6543);
nand U7221 (N_7221,N_6755,N_6961);
xor U7222 (N_7222,N_6852,N_6643);
or U7223 (N_7223,N_6989,N_6774);
nand U7224 (N_7224,N_6510,N_6587);
nor U7225 (N_7225,N_6823,N_6931);
nand U7226 (N_7226,N_6734,N_6930);
nor U7227 (N_7227,N_6644,N_6844);
nor U7228 (N_7228,N_6584,N_6911);
nand U7229 (N_7229,N_6941,N_6992);
and U7230 (N_7230,N_6726,N_6964);
or U7231 (N_7231,N_6517,N_6767);
or U7232 (N_7232,N_6865,N_6639);
or U7233 (N_7233,N_6722,N_6899);
and U7234 (N_7234,N_6953,N_6652);
and U7235 (N_7235,N_6723,N_6649);
nor U7236 (N_7236,N_6626,N_6679);
nand U7237 (N_7237,N_6983,N_6637);
xor U7238 (N_7238,N_6682,N_6694);
nor U7239 (N_7239,N_6758,N_6932);
nor U7240 (N_7240,N_6534,N_6672);
nand U7241 (N_7241,N_6835,N_6735);
nand U7242 (N_7242,N_6508,N_6505);
nand U7243 (N_7243,N_6529,N_6566);
or U7244 (N_7244,N_6710,N_6555);
or U7245 (N_7245,N_6912,N_6949);
xor U7246 (N_7246,N_6993,N_6686);
nand U7247 (N_7247,N_6974,N_6846);
and U7248 (N_7248,N_6919,N_6545);
nand U7249 (N_7249,N_6750,N_6784);
or U7250 (N_7250,N_6982,N_6849);
and U7251 (N_7251,N_6758,N_6742);
and U7252 (N_7252,N_6763,N_6669);
xnor U7253 (N_7253,N_6561,N_6791);
nand U7254 (N_7254,N_6530,N_6833);
nor U7255 (N_7255,N_6891,N_6800);
or U7256 (N_7256,N_6623,N_6634);
xnor U7257 (N_7257,N_6718,N_6946);
nor U7258 (N_7258,N_6986,N_6747);
or U7259 (N_7259,N_6754,N_6547);
nand U7260 (N_7260,N_6821,N_6902);
nor U7261 (N_7261,N_6530,N_6557);
or U7262 (N_7262,N_6841,N_6524);
or U7263 (N_7263,N_6852,N_6536);
nor U7264 (N_7264,N_6767,N_6882);
nand U7265 (N_7265,N_6909,N_6696);
xnor U7266 (N_7266,N_6555,N_6922);
or U7267 (N_7267,N_6763,N_6726);
nor U7268 (N_7268,N_6880,N_6887);
or U7269 (N_7269,N_6683,N_6660);
nand U7270 (N_7270,N_6985,N_6942);
nor U7271 (N_7271,N_6648,N_6828);
and U7272 (N_7272,N_6587,N_6956);
nor U7273 (N_7273,N_6902,N_6501);
or U7274 (N_7274,N_6997,N_6598);
and U7275 (N_7275,N_6903,N_6961);
nor U7276 (N_7276,N_6978,N_6962);
or U7277 (N_7277,N_6527,N_6838);
nor U7278 (N_7278,N_6530,N_6970);
nor U7279 (N_7279,N_6855,N_6859);
nand U7280 (N_7280,N_6693,N_6923);
nor U7281 (N_7281,N_6551,N_6882);
or U7282 (N_7282,N_6925,N_6513);
xor U7283 (N_7283,N_6920,N_6716);
nor U7284 (N_7284,N_6979,N_6801);
nor U7285 (N_7285,N_6886,N_6631);
and U7286 (N_7286,N_6761,N_6534);
or U7287 (N_7287,N_6979,N_6821);
nor U7288 (N_7288,N_6510,N_6504);
or U7289 (N_7289,N_6717,N_6799);
xor U7290 (N_7290,N_6811,N_6762);
and U7291 (N_7291,N_6754,N_6893);
and U7292 (N_7292,N_6600,N_6792);
xor U7293 (N_7293,N_6888,N_6904);
nor U7294 (N_7294,N_6736,N_6660);
or U7295 (N_7295,N_6954,N_6715);
xnor U7296 (N_7296,N_6830,N_6917);
xnor U7297 (N_7297,N_6902,N_6596);
and U7298 (N_7298,N_6504,N_6884);
xor U7299 (N_7299,N_6571,N_6739);
nor U7300 (N_7300,N_6865,N_6883);
and U7301 (N_7301,N_6783,N_6780);
and U7302 (N_7302,N_6754,N_6540);
nand U7303 (N_7303,N_6740,N_6597);
and U7304 (N_7304,N_6741,N_6785);
and U7305 (N_7305,N_6507,N_6952);
nand U7306 (N_7306,N_6596,N_6973);
or U7307 (N_7307,N_6917,N_6945);
nand U7308 (N_7308,N_6985,N_6959);
nand U7309 (N_7309,N_6644,N_6608);
xnor U7310 (N_7310,N_6564,N_6629);
and U7311 (N_7311,N_6817,N_6616);
or U7312 (N_7312,N_6745,N_6998);
nand U7313 (N_7313,N_6891,N_6939);
or U7314 (N_7314,N_6625,N_6598);
and U7315 (N_7315,N_6693,N_6999);
xnor U7316 (N_7316,N_6847,N_6890);
and U7317 (N_7317,N_6797,N_6659);
and U7318 (N_7318,N_6607,N_6841);
nor U7319 (N_7319,N_6808,N_6771);
or U7320 (N_7320,N_6888,N_6870);
and U7321 (N_7321,N_6994,N_6602);
nand U7322 (N_7322,N_6867,N_6949);
nand U7323 (N_7323,N_6674,N_6936);
and U7324 (N_7324,N_6845,N_6759);
nor U7325 (N_7325,N_6652,N_6854);
nand U7326 (N_7326,N_6719,N_6860);
and U7327 (N_7327,N_6892,N_6820);
nor U7328 (N_7328,N_6517,N_6988);
xnor U7329 (N_7329,N_6690,N_6731);
or U7330 (N_7330,N_6628,N_6710);
nand U7331 (N_7331,N_6560,N_6689);
nand U7332 (N_7332,N_6662,N_6505);
nor U7333 (N_7333,N_6836,N_6969);
xor U7334 (N_7334,N_6787,N_6960);
or U7335 (N_7335,N_6649,N_6504);
and U7336 (N_7336,N_6952,N_6581);
xnor U7337 (N_7337,N_6990,N_6823);
or U7338 (N_7338,N_6908,N_6513);
or U7339 (N_7339,N_6885,N_6909);
nand U7340 (N_7340,N_6649,N_6827);
xor U7341 (N_7341,N_6983,N_6877);
nand U7342 (N_7342,N_6837,N_6961);
nand U7343 (N_7343,N_6662,N_6776);
nand U7344 (N_7344,N_6586,N_6546);
and U7345 (N_7345,N_6720,N_6647);
nor U7346 (N_7346,N_6847,N_6978);
nand U7347 (N_7347,N_6678,N_6656);
nor U7348 (N_7348,N_6804,N_6510);
nor U7349 (N_7349,N_6773,N_6531);
xnor U7350 (N_7350,N_6828,N_6708);
xnor U7351 (N_7351,N_6749,N_6979);
and U7352 (N_7352,N_6748,N_6870);
or U7353 (N_7353,N_6802,N_6763);
nand U7354 (N_7354,N_6971,N_6784);
or U7355 (N_7355,N_6796,N_6933);
and U7356 (N_7356,N_6794,N_6594);
and U7357 (N_7357,N_6681,N_6614);
nor U7358 (N_7358,N_6836,N_6522);
nor U7359 (N_7359,N_6989,N_6966);
nor U7360 (N_7360,N_6735,N_6677);
and U7361 (N_7361,N_6738,N_6764);
nand U7362 (N_7362,N_6681,N_6995);
xor U7363 (N_7363,N_6550,N_6858);
nor U7364 (N_7364,N_6890,N_6599);
xor U7365 (N_7365,N_6892,N_6624);
nor U7366 (N_7366,N_6515,N_6596);
or U7367 (N_7367,N_6894,N_6702);
or U7368 (N_7368,N_6829,N_6562);
nand U7369 (N_7369,N_6736,N_6942);
xnor U7370 (N_7370,N_6606,N_6633);
xor U7371 (N_7371,N_6957,N_6568);
or U7372 (N_7372,N_6809,N_6674);
nor U7373 (N_7373,N_6887,N_6818);
nor U7374 (N_7374,N_6901,N_6728);
and U7375 (N_7375,N_6881,N_6592);
nand U7376 (N_7376,N_6788,N_6502);
or U7377 (N_7377,N_6632,N_6800);
xor U7378 (N_7378,N_6711,N_6550);
or U7379 (N_7379,N_6625,N_6913);
nor U7380 (N_7380,N_6825,N_6824);
nor U7381 (N_7381,N_6714,N_6540);
or U7382 (N_7382,N_6853,N_6627);
xnor U7383 (N_7383,N_6991,N_6629);
nor U7384 (N_7384,N_6888,N_6983);
and U7385 (N_7385,N_6655,N_6779);
and U7386 (N_7386,N_6757,N_6847);
nand U7387 (N_7387,N_6897,N_6948);
nor U7388 (N_7388,N_6892,N_6754);
nand U7389 (N_7389,N_6931,N_6598);
and U7390 (N_7390,N_6949,N_6588);
and U7391 (N_7391,N_6854,N_6879);
xnor U7392 (N_7392,N_6983,N_6764);
nand U7393 (N_7393,N_6505,N_6844);
nor U7394 (N_7394,N_6910,N_6534);
xor U7395 (N_7395,N_6707,N_6542);
or U7396 (N_7396,N_6797,N_6845);
or U7397 (N_7397,N_6903,N_6692);
nor U7398 (N_7398,N_6944,N_6744);
and U7399 (N_7399,N_6595,N_6981);
xor U7400 (N_7400,N_6847,N_6985);
or U7401 (N_7401,N_6942,N_6608);
and U7402 (N_7402,N_6832,N_6603);
nand U7403 (N_7403,N_6825,N_6797);
nand U7404 (N_7404,N_6618,N_6819);
xor U7405 (N_7405,N_6793,N_6981);
or U7406 (N_7406,N_6562,N_6750);
or U7407 (N_7407,N_6856,N_6654);
xor U7408 (N_7408,N_6864,N_6537);
nor U7409 (N_7409,N_6928,N_6668);
nand U7410 (N_7410,N_6953,N_6657);
xor U7411 (N_7411,N_6628,N_6669);
nand U7412 (N_7412,N_6809,N_6879);
xor U7413 (N_7413,N_6553,N_6822);
nor U7414 (N_7414,N_6536,N_6825);
nor U7415 (N_7415,N_6756,N_6738);
nand U7416 (N_7416,N_6869,N_6560);
nand U7417 (N_7417,N_6961,N_6778);
nor U7418 (N_7418,N_6538,N_6670);
and U7419 (N_7419,N_6825,N_6855);
xnor U7420 (N_7420,N_6984,N_6620);
nand U7421 (N_7421,N_6831,N_6734);
xor U7422 (N_7422,N_6606,N_6526);
nand U7423 (N_7423,N_6926,N_6726);
nand U7424 (N_7424,N_6894,N_6810);
xnor U7425 (N_7425,N_6771,N_6650);
or U7426 (N_7426,N_6875,N_6984);
xnor U7427 (N_7427,N_6569,N_6647);
or U7428 (N_7428,N_6604,N_6615);
nand U7429 (N_7429,N_6782,N_6595);
or U7430 (N_7430,N_6678,N_6630);
or U7431 (N_7431,N_6782,N_6671);
xnor U7432 (N_7432,N_6816,N_6518);
nor U7433 (N_7433,N_6903,N_6595);
xnor U7434 (N_7434,N_6975,N_6727);
or U7435 (N_7435,N_6695,N_6755);
nor U7436 (N_7436,N_6761,N_6554);
nor U7437 (N_7437,N_6937,N_6887);
and U7438 (N_7438,N_6904,N_6815);
or U7439 (N_7439,N_6918,N_6798);
and U7440 (N_7440,N_6772,N_6872);
nand U7441 (N_7441,N_6832,N_6515);
or U7442 (N_7442,N_6612,N_6777);
and U7443 (N_7443,N_6724,N_6642);
nor U7444 (N_7444,N_6778,N_6516);
nand U7445 (N_7445,N_6864,N_6909);
nor U7446 (N_7446,N_6942,N_6752);
and U7447 (N_7447,N_6764,N_6561);
or U7448 (N_7448,N_6603,N_6621);
nor U7449 (N_7449,N_6833,N_6808);
or U7450 (N_7450,N_6837,N_6617);
and U7451 (N_7451,N_6868,N_6720);
xor U7452 (N_7452,N_6830,N_6837);
and U7453 (N_7453,N_6874,N_6731);
or U7454 (N_7454,N_6784,N_6716);
and U7455 (N_7455,N_6725,N_6953);
or U7456 (N_7456,N_6803,N_6900);
xnor U7457 (N_7457,N_6879,N_6788);
or U7458 (N_7458,N_6524,N_6667);
nor U7459 (N_7459,N_6884,N_6572);
or U7460 (N_7460,N_6655,N_6925);
nand U7461 (N_7461,N_6834,N_6789);
xnor U7462 (N_7462,N_6729,N_6592);
nor U7463 (N_7463,N_6768,N_6664);
and U7464 (N_7464,N_6906,N_6884);
and U7465 (N_7465,N_6731,N_6532);
and U7466 (N_7466,N_6843,N_6521);
nor U7467 (N_7467,N_6523,N_6879);
xor U7468 (N_7468,N_6989,N_6724);
or U7469 (N_7469,N_6780,N_6757);
xnor U7470 (N_7470,N_6683,N_6784);
nand U7471 (N_7471,N_6901,N_6663);
nand U7472 (N_7472,N_6700,N_6728);
nand U7473 (N_7473,N_6597,N_6724);
xor U7474 (N_7474,N_6896,N_6935);
or U7475 (N_7475,N_6824,N_6671);
nand U7476 (N_7476,N_6581,N_6974);
or U7477 (N_7477,N_6739,N_6710);
and U7478 (N_7478,N_6575,N_6518);
and U7479 (N_7479,N_6617,N_6611);
xnor U7480 (N_7480,N_6755,N_6517);
nand U7481 (N_7481,N_6502,N_6706);
nor U7482 (N_7482,N_6529,N_6558);
or U7483 (N_7483,N_6539,N_6763);
or U7484 (N_7484,N_6728,N_6501);
nor U7485 (N_7485,N_6797,N_6543);
or U7486 (N_7486,N_6814,N_6977);
nand U7487 (N_7487,N_6718,N_6741);
nand U7488 (N_7488,N_6871,N_6572);
nor U7489 (N_7489,N_6617,N_6824);
nor U7490 (N_7490,N_6979,N_6596);
or U7491 (N_7491,N_6554,N_6548);
and U7492 (N_7492,N_6848,N_6690);
or U7493 (N_7493,N_6673,N_6629);
xnor U7494 (N_7494,N_6553,N_6521);
and U7495 (N_7495,N_6577,N_6785);
nor U7496 (N_7496,N_6510,N_6954);
nand U7497 (N_7497,N_6602,N_6680);
or U7498 (N_7498,N_6961,N_6851);
or U7499 (N_7499,N_6948,N_6664);
xnor U7500 (N_7500,N_7287,N_7310);
nor U7501 (N_7501,N_7493,N_7169);
xor U7502 (N_7502,N_7379,N_7319);
or U7503 (N_7503,N_7035,N_7429);
or U7504 (N_7504,N_7057,N_7178);
or U7505 (N_7505,N_7220,N_7311);
xnor U7506 (N_7506,N_7361,N_7330);
nor U7507 (N_7507,N_7328,N_7273);
and U7508 (N_7508,N_7398,N_7478);
and U7509 (N_7509,N_7144,N_7142);
nor U7510 (N_7510,N_7143,N_7170);
nand U7511 (N_7511,N_7141,N_7078);
and U7512 (N_7512,N_7331,N_7329);
nor U7513 (N_7513,N_7115,N_7473);
xor U7514 (N_7514,N_7292,N_7200);
nand U7515 (N_7515,N_7425,N_7207);
nor U7516 (N_7516,N_7355,N_7348);
nand U7517 (N_7517,N_7135,N_7276);
or U7518 (N_7518,N_7041,N_7448);
and U7519 (N_7519,N_7288,N_7496);
and U7520 (N_7520,N_7214,N_7060);
xnor U7521 (N_7521,N_7353,N_7123);
xnor U7522 (N_7522,N_7300,N_7122);
or U7523 (N_7523,N_7295,N_7154);
nand U7524 (N_7524,N_7008,N_7106);
nand U7525 (N_7525,N_7388,N_7347);
nor U7526 (N_7526,N_7335,N_7212);
or U7527 (N_7527,N_7252,N_7087);
or U7528 (N_7528,N_7364,N_7127);
and U7529 (N_7529,N_7180,N_7437);
and U7530 (N_7530,N_7188,N_7133);
nand U7531 (N_7531,N_7334,N_7193);
nor U7532 (N_7532,N_7480,N_7371);
or U7533 (N_7533,N_7067,N_7419);
or U7534 (N_7534,N_7010,N_7080);
nor U7535 (N_7535,N_7337,N_7174);
or U7536 (N_7536,N_7377,N_7103);
or U7537 (N_7537,N_7420,N_7268);
xor U7538 (N_7538,N_7394,N_7303);
xnor U7539 (N_7539,N_7109,N_7269);
nand U7540 (N_7540,N_7224,N_7343);
nor U7541 (N_7541,N_7237,N_7153);
xor U7542 (N_7542,N_7484,N_7165);
nor U7543 (N_7543,N_7291,N_7223);
and U7544 (N_7544,N_7190,N_7294);
or U7545 (N_7545,N_7454,N_7168);
and U7546 (N_7546,N_7129,N_7023);
and U7547 (N_7547,N_7099,N_7069);
nand U7548 (N_7548,N_7261,N_7403);
nor U7549 (N_7549,N_7375,N_7382);
nand U7550 (N_7550,N_7018,N_7302);
nand U7551 (N_7551,N_7251,N_7322);
and U7552 (N_7552,N_7246,N_7274);
nand U7553 (N_7553,N_7068,N_7076);
or U7554 (N_7554,N_7009,N_7275);
and U7555 (N_7555,N_7461,N_7208);
or U7556 (N_7556,N_7264,N_7326);
nand U7557 (N_7557,N_7203,N_7259);
xnor U7558 (N_7558,N_7185,N_7105);
and U7559 (N_7559,N_7477,N_7043);
or U7560 (N_7560,N_7338,N_7148);
nor U7561 (N_7561,N_7137,N_7247);
or U7562 (N_7562,N_7464,N_7235);
or U7563 (N_7563,N_7262,N_7469);
and U7564 (N_7564,N_7071,N_7307);
nor U7565 (N_7565,N_7363,N_7152);
nor U7566 (N_7566,N_7086,N_7238);
nand U7567 (N_7567,N_7216,N_7255);
nand U7568 (N_7568,N_7050,N_7034);
nand U7569 (N_7569,N_7279,N_7245);
and U7570 (N_7570,N_7423,N_7108);
and U7571 (N_7571,N_7285,N_7431);
xnor U7572 (N_7572,N_7140,N_7472);
or U7573 (N_7573,N_7380,N_7352);
or U7574 (N_7574,N_7145,N_7362);
nand U7575 (N_7575,N_7440,N_7349);
and U7576 (N_7576,N_7485,N_7456);
nor U7577 (N_7577,N_7317,N_7387);
and U7578 (N_7578,N_7198,N_7128);
nor U7579 (N_7579,N_7400,N_7421);
xor U7580 (N_7580,N_7236,N_7230);
and U7581 (N_7581,N_7097,N_7098);
xnor U7582 (N_7582,N_7093,N_7408);
or U7583 (N_7583,N_7376,N_7160);
or U7584 (N_7584,N_7004,N_7030);
nand U7585 (N_7585,N_7181,N_7042);
xnor U7586 (N_7586,N_7370,N_7029);
nand U7587 (N_7587,N_7175,N_7323);
xnor U7588 (N_7588,N_7254,N_7470);
nor U7589 (N_7589,N_7197,N_7266);
or U7590 (N_7590,N_7290,N_7209);
and U7591 (N_7591,N_7217,N_7487);
nand U7592 (N_7592,N_7369,N_7150);
nand U7593 (N_7593,N_7455,N_7155);
nand U7594 (N_7594,N_7118,N_7418);
nand U7595 (N_7595,N_7022,N_7146);
or U7596 (N_7596,N_7013,N_7134);
or U7597 (N_7597,N_7281,N_7450);
nand U7598 (N_7598,N_7339,N_7182);
and U7599 (N_7599,N_7499,N_7164);
nor U7600 (N_7600,N_7066,N_7457);
or U7601 (N_7601,N_7244,N_7354);
nand U7602 (N_7602,N_7124,N_7063);
nor U7603 (N_7603,N_7490,N_7390);
or U7604 (N_7604,N_7094,N_7414);
nand U7605 (N_7605,N_7119,N_7359);
nor U7606 (N_7606,N_7081,N_7096);
and U7607 (N_7607,N_7441,N_7312);
and U7608 (N_7608,N_7072,N_7399);
nand U7609 (N_7609,N_7172,N_7020);
or U7610 (N_7610,N_7025,N_7346);
nor U7611 (N_7611,N_7271,N_7358);
nor U7612 (N_7612,N_7044,N_7495);
nand U7613 (N_7613,N_7491,N_7107);
xor U7614 (N_7614,N_7397,N_7006);
or U7615 (N_7615,N_7306,N_7250);
nand U7616 (N_7616,N_7201,N_7016);
nand U7617 (N_7617,N_7187,N_7471);
or U7618 (N_7618,N_7136,N_7131);
and U7619 (N_7619,N_7012,N_7070);
or U7620 (N_7620,N_7378,N_7406);
nor U7621 (N_7621,N_7301,N_7084);
or U7622 (N_7622,N_7412,N_7341);
and U7623 (N_7623,N_7219,N_7049);
nand U7624 (N_7624,N_7383,N_7202);
nand U7625 (N_7625,N_7272,N_7416);
and U7626 (N_7626,N_7167,N_7442);
nand U7627 (N_7627,N_7280,N_7054);
nor U7628 (N_7628,N_7260,N_7374);
nor U7629 (N_7629,N_7002,N_7407);
or U7630 (N_7630,N_7289,N_7233);
or U7631 (N_7631,N_7267,N_7433);
nand U7632 (N_7632,N_7462,N_7074);
nand U7633 (N_7633,N_7147,N_7100);
or U7634 (N_7634,N_7316,N_7062);
xnor U7635 (N_7635,N_7028,N_7075);
nor U7636 (N_7636,N_7277,N_7270);
or U7637 (N_7637,N_7263,N_7196);
or U7638 (N_7638,N_7253,N_7417);
xnor U7639 (N_7639,N_7007,N_7305);
and U7640 (N_7640,N_7422,N_7488);
nand U7641 (N_7641,N_7248,N_7432);
or U7642 (N_7642,N_7024,N_7117);
nor U7643 (N_7643,N_7090,N_7333);
nor U7644 (N_7644,N_7282,N_7411);
nand U7645 (N_7645,N_7315,N_7151);
nand U7646 (N_7646,N_7047,N_7226);
nor U7647 (N_7647,N_7475,N_7058);
xnor U7648 (N_7648,N_7194,N_7110);
or U7649 (N_7649,N_7061,N_7005);
nor U7650 (N_7650,N_7438,N_7113);
nand U7651 (N_7651,N_7498,N_7467);
and U7652 (N_7652,N_7381,N_7242);
nand U7653 (N_7653,N_7162,N_7221);
and U7654 (N_7654,N_7206,N_7130);
xor U7655 (N_7655,N_7336,N_7447);
nand U7656 (N_7656,N_7111,N_7227);
nand U7657 (N_7657,N_7458,N_7157);
nor U7658 (N_7658,N_7121,N_7396);
nand U7659 (N_7659,N_7304,N_7231);
xor U7660 (N_7660,N_7037,N_7017);
and U7661 (N_7661,N_7095,N_7345);
xnor U7662 (N_7662,N_7476,N_7278);
xor U7663 (N_7663,N_7021,N_7222);
and U7664 (N_7664,N_7159,N_7240);
or U7665 (N_7665,N_7173,N_7427);
or U7666 (N_7666,N_7318,N_7393);
and U7667 (N_7667,N_7356,N_7213);
and U7668 (N_7668,N_7309,N_7483);
nor U7669 (N_7669,N_7112,N_7052);
nand U7670 (N_7670,N_7365,N_7293);
and U7671 (N_7671,N_7019,N_7463);
and U7672 (N_7672,N_7039,N_7229);
and U7673 (N_7673,N_7126,N_7204);
nand U7674 (N_7674,N_7410,N_7497);
or U7675 (N_7675,N_7386,N_7139);
xnor U7676 (N_7676,N_7401,N_7104);
and U7677 (N_7677,N_7092,N_7055);
nand U7678 (N_7678,N_7205,N_7367);
nor U7679 (N_7679,N_7232,N_7031);
or U7680 (N_7680,N_7015,N_7073);
nand U7681 (N_7681,N_7439,N_7426);
nor U7682 (N_7682,N_7298,N_7184);
or U7683 (N_7683,N_7189,N_7166);
nor U7684 (N_7684,N_7389,N_7077);
xor U7685 (N_7685,N_7011,N_7195);
and U7686 (N_7686,N_7492,N_7296);
or U7687 (N_7687,N_7191,N_7065);
nand U7688 (N_7688,N_7038,N_7079);
and U7689 (N_7689,N_7340,N_7384);
nor U7690 (N_7690,N_7258,N_7284);
or U7691 (N_7691,N_7459,N_7372);
and U7692 (N_7692,N_7428,N_7199);
or U7693 (N_7693,N_7466,N_7132);
xnor U7694 (N_7694,N_7391,N_7064);
nor U7695 (N_7695,N_7368,N_7033);
nor U7696 (N_7696,N_7215,N_7460);
and U7697 (N_7697,N_7211,N_7045);
nand U7698 (N_7698,N_7056,N_7357);
and U7699 (N_7699,N_7489,N_7482);
xnor U7700 (N_7700,N_7149,N_7082);
or U7701 (N_7701,N_7360,N_7465);
nand U7702 (N_7702,N_7350,N_7083);
xnor U7703 (N_7703,N_7449,N_7225);
nor U7704 (N_7704,N_7046,N_7051);
and U7705 (N_7705,N_7210,N_7453);
xor U7706 (N_7706,N_7088,N_7243);
xnor U7707 (N_7707,N_7299,N_7228);
xnor U7708 (N_7708,N_7446,N_7395);
xnor U7709 (N_7709,N_7183,N_7451);
and U7710 (N_7710,N_7404,N_7313);
nor U7711 (N_7711,N_7102,N_7101);
nor U7712 (N_7712,N_7125,N_7314);
nand U7713 (N_7713,N_7032,N_7468);
nor U7714 (N_7714,N_7265,N_7014);
or U7715 (N_7715,N_7308,N_7001);
xor U7716 (N_7716,N_7089,N_7435);
or U7717 (N_7717,N_7256,N_7156);
nor U7718 (N_7718,N_7344,N_7324);
nor U7719 (N_7719,N_7486,N_7479);
nor U7720 (N_7720,N_7257,N_7320);
and U7721 (N_7721,N_7409,N_7239);
xor U7722 (N_7722,N_7163,N_7444);
or U7723 (N_7723,N_7436,N_7138);
and U7724 (N_7724,N_7218,N_7241);
nor U7725 (N_7725,N_7434,N_7116);
and U7726 (N_7726,N_7171,N_7120);
nand U7727 (N_7727,N_7003,N_7443);
nor U7728 (N_7728,N_7325,N_7161);
xor U7729 (N_7729,N_7297,N_7405);
nand U7730 (N_7730,N_7053,N_7192);
and U7731 (N_7731,N_7332,N_7283);
and U7732 (N_7732,N_7249,N_7481);
xor U7733 (N_7733,N_7402,N_7413);
or U7734 (N_7734,N_7114,N_7186);
nor U7735 (N_7735,N_7385,N_7430);
and U7736 (N_7736,N_7474,N_7286);
nand U7737 (N_7737,N_7366,N_7000);
and U7738 (N_7738,N_7321,N_7392);
nand U7739 (N_7739,N_7234,N_7452);
xnor U7740 (N_7740,N_7036,N_7026);
nand U7741 (N_7741,N_7424,N_7176);
xnor U7742 (N_7742,N_7027,N_7040);
or U7743 (N_7743,N_7091,N_7445);
xnor U7744 (N_7744,N_7179,N_7085);
and U7745 (N_7745,N_7327,N_7342);
or U7746 (N_7746,N_7373,N_7048);
or U7747 (N_7747,N_7177,N_7158);
nor U7748 (N_7748,N_7494,N_7351);
nand U7749 (N_7749,N_7415,N_7059);
nor U7750 (N_7750,N_7126,N_7220);
nor U7751 (N_7751,N_7025,N_7267);
nor U7752 (N_7752,N_7244,N_7376);
nand U7753 (N_7753,N_7290,N_7258);
xor U7754 (N_7754,N_7021,N_7285);
nor U7755 (N_7755,N_7089,N_7026);
or U7756 (N_7756,N_7395,N_7053);
or U7757 (N_7757,N_7080,N_7085);
nand U7758 (N_7758,N_7202,N_7425);
and U7759 (N_7759,N_7174,N_7113);
or U7760 (N_7760,N_7184,N_7359);
nand U7761 (N_7761,N_7084,N_7029);
nand U7762 (N_7762,N_7443,N_7252);
nor U7763 (N_7763,N_7026,N_7298);
xnor U7764 (N_7764,N_7266,N_7350);
nor U7765 (N_7765,N_7080,N_7017);
or U7766 (N_7766,N_7031,N_7465);
nor U7767 (N_7767,N_7249,N_7460);
xnor U7768 (N_7768,N_7264,N_7219);
nor U7769 (N_7769,N_7382,N_7091);
nor U7770 (N_7770,N_7495,N_7261);
nand U7771 (N_7771,N_7324,N_7390);
or U7772 (N_7772,N_7191,N_7003);
nand U7773 (N_7773,N_7183,N_7132);
and U7774 (N_7774,N_7364,N_7083);
nand U7775 (N_7775,N_7027,N_7029);
and U7776 (N_7776,N_7205,N_7046);
nand U7777 (N_7777,N_7474,N_7138);
or U7778 (N_7778,N_7187,N_7387);
nand U7779 (N_7779,N_7286,N_7423);
nand U7780 (N_7780,N_7173,N_7357);
and U7781 (N_7781,N_7105,N_7104);
nand U7782 (N_7782,N_7163,N_7132);
nor U7783 (N_7783,N_7467,N_7227);
and U7784 (N_7784,N_7288,N_7223);
nand U7785 (N_7785,N_7048,N_7491);
nand U7786 (N_7786,N_7334,N_7259);
or U7787 (N_7787,N_7276,N_7070);
xnor U7788 (N_7788,N_7404,N_7322);
nand U7789 (N_7789,N_7408,N_7422);
xor U7790 (N_7790,N_7382,N_7448);
nand U7791 (N_7791,N_7126,N_7473);
and U7792 (N_7792,N_7023,N_7094);
and U7793 (N_7793,N_7315,N_7147);
or U7794 (N_7794,N_7285,N_7151);
or U7795 (N_7795,N_7048,N_7285);
and U7796 (N_7796,N_7430,N_7493);
or U7797 (N_7797,N_7130,N_7067);
nand U7798 (N_7798,N_7018,N_7363);
nand U7799 (N_7799,N_7260,N_7019);
xor U7800 (N_7800,N_7478,N_7152);
and U7801 (N_7801,N_7208,N_7101);
xnor U7802 (N_7802,N_7399,N_7467);
xnor U7803 (N_7803,N_7027,N_7459);
xor U7804 (N_7804,N_7100,N_7129);
or U7805 (N_7805,N_7361,N_7469);
nand U7806 (N_7806,N_7171,N_7116);
or U7807 (N_7807,N_7240,N_7044);
and U7808 (N_7808,N_7312,N_7186);
xor U7809 (N_7809,N_7147,N_7179);
or U7810 (N_7810,N_7109,N_7208);
nor U7811 (N_7811,N_7207,N_7220);
nor U7812 (N_7812,N_7418,N_7236);
or U7813 (N_7813,N_7101,N_7142);
nor U7814 (N_7814,N_7354,N_7243);
or U7815 (N_7815,N_7011,N_7234);
nor U7816 (N_7816,N_7345,N_7059);
and U7817 (N_7817,N_7192,N_7099);
and U7818 (N_7818,N_7257,N_7126);
or U7819 (N_7819,N_7229,N_7099);
xnor U7820 (N_7820,N_7346,N_7100);
xnor U7821 (N_7821,N_7054,N_7072);
and U7822 (N_7822,N_7399,N_7209);
and U7823 (N_7823,N_7088,N_7083);
and U7824 (N_7824,N_7469,N_7242);
nand U7825 (N_7825,N_7262,N_7465);
nand U7826 (N_7826,N_7172,N_7214);
or U7827 (N_7827,N_7101,N_7448);
and U7828 (N_7828,N_7207,N_7394);
xnor U7829 (N_7829,N_7254,N_7092);
and U7830 (N_7830,N_7020,N_7131);
nand U7831 (N_7831,N_7147,N_7335);
xnor U7832 (N_7832,N_7071,N_7233);
nor U7833 (N_7833,N_7486,N_7455);
nand U7834 (N_7834,N_7156,N_7259);
and U7835 (N_7835,N_7057,N_7004);
or U7836 (N_7836,N_7226,N_7089);
nand U7837 (N_7837,N_7221,N_7235);
xor U7838 (N_7838,N_7190,N_7037);
nor U7839 (N_7839,N_7031,N_7352);
nor U7840 (N_7840,N_7323,N_7012);
xnor U7841 (N_7841,N_7399,N_7409);
nand U7842 (N_7842,N_7121,N_7093);
xor U7843 (N_7843,N_7051,N_7228);
xor U7844 (N_7844,N_7386,N_7025);
nor U7845 (N_7845,N_7043,N_7152);
nor U7846 (N_7846,N_7236,N_7348);
nor U7847 (N_7847,N_7083,N_7422);
and U7848 (N_7848,N_7136,N_7141);
and U7849 (N_7849,N_7423,N_7402);
nor U7850 (N_7850,N_7367,N_7402);
or U7851 (N_7851,N_7421,N_7127);
or U7852 (N_7852,N_7165,N_7172);
and U7853 (N_7853,N_7098,N_7354);
nor U7854 (N_7854,N_7039,N_7304);
nand U7855 (N_7855,N_7300,N_7139);
xor U7856 (N_7856,N_7360,N_7234);
xor U7857 (N_7857,N_7320,N_7150);
xnor U7858 (N_7858,N_7255,N_7166);
nand U7859 (N_7859,N_7400,N_7494);
nor U7860 (N_7860,N_7056,N_7484);
and U7861 (N_7861,N_7173,N_7326);
xnor U7862 (N_7862,N_7033,N_7121);
and U7863 (N_7863,N_7044,N_7434);
and U7864 (N_7864,N_7272,N_7028);
xnor U7865 (N_7865,N_7281,N_7411);
nor U7866 (N_7866,N_7351,N_7136);
nand U7867 (N_7867,N_7463,N_7467);
nor U7868 (N_7868,N_7471,N_7265);
and U7869 (N_7869,N_7323,N_7056);
or U7870 (N_7870,N_7256,N_7023);
nor U7871 (N_7871,N_7312,N_7391);
or U7872 (N_7872,N_7425,N_7238);
xnor U7873 (N_7873,N_7102,N_7071);
or U7874 (N_7874,N_7458,N_7062);
nor U7875 (N_7875,N_7328,N_7456);
or U7876 (N_7876,N_7490,N_7032);
xor U7877 (N_7877,N_7163,N_7293);
or U7878 (N_7878,N_7412,N_7225);
nand U7879 (N_7879,N_7194,N_7026);
nor U7880 (N_7880,N_7146,N_7393);
and U7881 (N_7881,N_7419,N_7372);
nor U7882 (N_7882,N_7202,N_7237);
or U7883 (N_7883,N_7190,N_7044);
nor U7884 (N_7884,N_7144,N_7130);
and U7885 (N_7885,N_7213,N_7086);
nor U7886 (N_7886,N_7181,N_7475);
or U7887 (N_7887,N_7129,N_7088);
nand U7888 (N_7888,N_7396,N_7087);
or U7889 (N_7889,N_7377,N_7478);
and U7890 (N_7890,N_7147,N_7234);
or U7891 (N_7891,N_7361,N_7349);
nor U7892 (N_7892,N_7037,N_7344);
nand U7893 (N_7893,N_7117,N_7006);
and U7894 (N_7894,N_7439,N_7014);
or U7895 (N_7895,N_7066,N_7336);
nand U7896 (N_7896,N_7265,N_7250);
nand U7897 (N_7897,N_7215,N_7216);
and U7898 (N_7898,N_7309,N_7399);
xor U7899 (N_7899,N_7388,N_7075);
nand U7900 (N_7900,N_7445,N_7149);
or U7901 (N_7901,N_7397,N_7384);
xor U7902 (N_7902,N_7308,N_7002);
and U7903 (N_7903,N_7111,N_7360);
nor U7904 (N_7904,N_7073,N_7336);
xnor U7905 (N_7905,N_7082,N_7220);
xnor U7906 (N_7906,N_7267,N_7084);
nor U7907 (N_7907,N_7312,N_7454);
xor U7908 (N_7908,N_7356,N_7150);
nor U7909 (N_7909,N_7397,N_7337);
xor U7910 (N_7910,N_7165,N_7157);
and U7911 (N_7911,N_7394,N_7152);
or U7912 (N_7912,N_7039,N_7182);
nand U7913 (N_7913,N_7489,N_7391);
nor U7914 (N_7914,N_7259,N_7284);
nand U7915 (N_7915,N_7013,N_7341);
nand U7916 (N_7916,N_7470,N_7443);
nand U7917 (N_7917,N_7393,N_7147);
nor U7918 (N_7918,N_7142,N_7233);
xnor U7919 (N_7919,N_7487,N_7122);
nand U7920 (N_7920,N_7367,N_7376);
nor U7921 (N_7921,N_7240,N_7060);
nand U7922 (N_7922,N_7154,N_7359);
and U7923 (N_7923,N_7359,N_7487);
or U7924 (N_7924,N_7050,N_7037);
nand U7925 (N_7925,N_7394,N_7331);
or U7926 (N_7926,N_7190,N_7223);
or U7927 (N_7927,N_7295,N_7303);
or U7928 (N_7928,N_7277,N_7114);
or U7929 (N_7929,N_7445,N_7268);
nand U7930 (N_7930,N_7360,N_7345);
nor U7931 (N_7931,N_7351,N_7147);
nor U7932 (N_7932,N_7125,N_7069);
nor U7933 (N_7933,N_7091,N_7085);
xor U7934 (N_7934,N_7191,N_7099);
or U7935 (N_7935,N_7194,N_7062);
and U7936 (N_7936,N_7373,N_7187);
xor U7937 (N_7937,N_7045,N_7161);
and U7938 (N_7938,N_7163,N_7326);
nand U7939 (N_7939,N_7154,N_7119);
xor U7940 (N_7940,N_7093,N_7289);
nand U7941 (N_7941,N_7429,N_7010);
and U7942 (N_7942,N_7120,N_7195);
xnor U7943 (N_7943,N_7462,N_7329);
nor U7944 (N_7944,N_7237,N_7067);
xnor U7945 (N_7945,N_7199,N_7488);
xnor U7946 (N_7946,N_7421,N_7482);
nand U7947 (N_7947,N_7223,N_7470);
nand U7948 (N_7948,N_7177,N_7142);
xnor U7949 (N_7949,N_7440,N_7467);
xor U7950 (N_7950,N_7439,N_7437);
nand U7951 (N_7951,N_7335,N_7129);
and U7952 (N_7952,N_7281,N_7142);
xnor U7953 (N_7953,N_7057,N_7249);
and U7954 (N_7954,N_7163,N_7233);
nand U7955 (N_7955,N_7337,N_7396);
and U7956 (N_7956,N_7150,N_7094);
and U7957 (N_7957,N_7375,N_7430);
and U7958 (N_7958,N_7288,N_7365);
nor U7959 (N_7959,N_7172,N_7438);
and U7960 (N_7960,N_7027,N_7440);
or U7961 (N_7961,N_7271,N_7299);
xor U7962 (N_7962,N_7379,N_7144);
nor U7963 (N_7963,N_7347,N_7093);
and U7964 (N_7964,N_7059,N_7324);
or U7965 (N_7965,N_7085,N_7307);
xor U7966 (N_7966,N_7411,N_7085);
nor U7967 (N_7967,N_7077,N_7349);
or U7968 (N_7968,N_7329,N_7191);
nor U7969 (N_7969,N_7441,N_7244);
nand U7970 (N_7970,N_7066,N_7339);
nand U7971 (N_7971,N_7034,N_7226);
nand U7972 (N_7972,N_7357,N_7413);
and U7973 (N_7973,N_7421,N_7163);
or U7974 (N_7974,N_7154,N_7011);
and U7975 (N_7975,N_7280,N_7293);
nor U7976 (N_7976,N_7438,N_7070);
nor U7977 (N_7977,N_7007,N_7444);
nor U7978 (N_7978,N_7061,N_7174);
nand U7979 (N_7979,N_7016,N_7358);
or U7980 (N_7980,N_7077,N_7087);
nand U7981 (N_7981,N_7492,N_7331);
nand U7982 (N_7982,N_7499,N_7385);
or U7983 (N_7983,N_7011,N_7389);
or U7984 (N_7984,N_7027,N_7106);
xor U7985 (N_7985,N_7271,N_7124);
and U7986 (N_7986,N_7282,N_7485);
and U7987 (N_7987,N_7450,N_7315);
nor U7988 (N_7988,N_7384,N_7206);
and U7989 (N_7989,N_7370,N_7057);
xor U7990 (N_7990,N_7450,N_7007);
nor U7991 (N_7991,N_7085,N_7108);
and U7992 (N_7992,N_7409,N_7489);
nor U7993 (N_7993,N_7431,N_7298);
xor U7994 (N_7994,N_7275,N_7336);
or U7995 (N_7995,N_7457,N_7406);
and U7996 (N_7996,N_7473,N_7222);
or U7997 (N_7997,N_7378,N_7273);
and U7998 (N_7998,N_7409,N_7235);
nor U7999 (N_7999,N_7421,N_7431);
or U8000 (N_8000,N_7657,N_7826);
or U8001 (N_8001,N_7516,N_7632);
xor U8002 (N_8002,N_7609,N_7899);
or U8003 (N_8003,N_7717,N_7754);
and U8004 (N_8004,N_7773,N_7944);
xnor U8005 (N_8005,N_7691,N_7786);
nand U8006 (N_8006,N_7770,N_7564);
and U8007 (N_8007,N_7812,N_7795);
xor U8008 (N_8008,N_7697,N_7558);
or U8009 (N_8009,N_7878,N_7517);
nand U8010 (N_8010,N_7612,N_7533);
nor U8011 (N_8011,N_7911,N_7521);
xnor U8012 (N_8012,N_7722,N_7654);
nand U8013 (N_8013,N_7872,N_7651);
and U8014 (N_8014,N_7844,N_7855);
and U8015 (N_8015,N_7822,N_7723);
or U8016 (N_8016,N_7730,N_7802);
nor U8017 (N_8017,N_7806,N_7928);
nand U8018 (N_8018,N_7737,N_7989);
nand U8019 (N_8019,N_7658,N_7853);
and U8020 (N_8020,N_7810,N_7715);
xnor U8021 (N_8021,N_7668,N_7549);
or U8022 (N_8022,N_7988,N_7663);
nand U8023 (N_8023,N_7809,N_7702);
nor U8024 (N_8024,N_7916,N_7856);
xnor U8025 (N_8025,N_7705,N_7774);
and U8026 (N_8026,N_7593,N_7743);
or U8027 (N_8027,N_7681,N_7985);
nand U8028 (N_8028,N_7947,N_7669);
and U8029 (N_8029,N_7778,N_7518);
xor U8030 (N_8030,N_7607,N_7502);
and U8031 (N_8031,N_7814,N_7863);
nor U8032 (N_8032,N_7596,N_7788);
or U8033 (N_8033,N_7652,N_7704);
and U8034 (N_8034,N_7628,N_7683);
nand U8035 (N_8035,N_7576,N_7676);
or U8036 (N_8036,N_7592,N_7962);
nand U8037 (N_8037,N_7557,N_7755);
and U8038 (N_8038,N_7957,N_7923);
or U8039 (N_8039,N_7567,N_7907);
or U8040 (N_8040,N_7610,N_7815);
nor U8041 (N_8041,N_7649,N_7700);
nor U8042 (N_8042,N_7752,N_7535);
nor U8043 (N_8043,N_7544,N_7677);
nor U8044 (N_8044,N_7827,N_7580);
nand U8045 (N_8045,N_7937,N_7572);
nand U8046 (N_8046,N_7581,N_7949);
nor U8047 (N_8047,N_7606,N_7884);
nand U8048 (N_8048,N_7945,N_7684);
or U8049 (N_8049,N_7685,N_7621);
nor U8050 (N_8050,N_7794,N_7779);
or U8051 (N_8051,N_7530,N_7742);
xnor U8052 (N_8052,N_7867,N_7999);
and U8053 (N_8053,N_7694,N_7699);
xnor U8054 (N_8054,N_7939,N_7843);
or U8055 (N_8055,N_7763,N_7909);
and U8056 (N_8056,N_7776,N_7725);
xnor U8057 (N_8057,N_7682,N_7539);
xnor U8058 (N_8058,N_7792,N_7751);
and U8059 (N_8059,N_7563,N_7602);
nand U8060 (N_8060,N_7793,N_7898);
xor U8061 (N_8061,N_7987,N_7970);
nor U8062 (N_8062,N_7869,N_7969);
nand U8063 (N_8063,N_7613,N_7588);
or U8064 (N_8064,N_7540,N_7750);
nor U8065 (N_8065,N_7775,N_7617);
or U8066 (N_8066,N_7847,N_7835);
or U8067 (N_8067,N_7706,N_7832);
nor U8068 (N_8068,N_7577,N_7645);
or U8069 (N_8069,N_7905,N_7870);
nand U8070 (N_8070,N_7789,N_7823);
or U8071 (N_8071,N_7862,N_7692);
nor U8072 (N_8072,N_7785,N_7841);
and U8073 (N_8073,N_7982,N_7967);
nor U8074 (N_8074,N_7858,N_7500);
nand U8075 (N_8075,N_7824,N_7696);
or U8076 (N_8076,N_7895,N_7943);
nor U8077 (N_8077,N_7514,N_7729);
nand U8078 (N_8078,N_7680,N_7532);
nand U8079 (N_8079,N_7719,N_7501);
or U8080 (N_8080,N_7850,N_7724);
xor U8081 (N_8081,N_7961,N_7587);
nand U8082 (N_8082,N_7687,N_7638);
nor U8083 (N_8083,N_7701,N_7805);
xnor U8084 (N_8084,N_7777,N_7511);
nand U8085 (N_8085,N_7546,N_7929);
and U8086 (N_8086,N_7974,N_7886);
nor U8087 (N_8087,N_7807,N_7594);
nand U8088 (N_8088,N_7551,N_7670);
or U8089 (N_8089,N_7880,N_7626);
and U8090 (N_8090,N_7507,N_7600);
and U8091 (N_8091,N_7978,N_7874);
or U8092 (N_8092,N_7550,N_7875);
or U8093 (N_8093,N_7510,N_7934);
nand U8094 (N_8094,N_7513,N_7848);
nand U8095 (N_8095,N_7762,N_7541);
and U8096 (N_8096,N_7548,N_7608);
xor U8097 (N_8097,N_7749,N_7710);
or U8098 (N_8098,N_7605,N_7857);
and U8099 (N_8099,N_7990,N_7842);
or U8100 (N_8100,N_7515,N_7634);
xor U8101 (N_8101,N_7619,N_7797);
nor U8102 (N_8102,N_7883,N_7915);
xnor U8103 (N_8103,N_7653,N_7554);
nor U8104 (N_8104,N_7868,N_7686);
nand U8105 (N_8105,N_7865,N_7964);
nand U8106 (N_8106,N_7845,N_7948);
or U8107 (N_8107,N_7721,N_7655);
and U8108 (N_8108,N_7647,N_7570);
nor U8109 (N_8109,N_7767,N_7735);
and U8110 (N_8110,N_7555,N_7892);
nand U8111 (N_8111,N_7582,N_7896);
nor U8112 (N_8112,N_7635,N_7958);
or U8113 (N_8113,N_7849,N_7831);
nand U8114 (N_8114,N_7666,N_7716);
nand U8115 (N_8115,N_7648,N_7575);
nand U8116 (N_8116,N_7796,N_7996);
nor U8117 (N_8117,N_7589,N_7938);
xor U8118 (N_8118,N_7525,N_7618);
or U8119 (N_8119,N_7667,N_7959);
nand U8120 (N_8120,N_7689,N_7556);
nor U8121 (N_8121,N_7597,N_7837);
or U8122 (N_8122,N_7818,N_7726);
nand U8123 (N_8123,N_7543,N_7674);
xnor U8124 (N_8124,N_7732,N_7560);
nor U8125 (N_8125,N_7906,N_7679);
xor U8126 (N_8126,N_7800,N_7568);
or U8127 (N_8127,N_7935,N_7641);
or U8128 (N_8128,N_7545,N_7889);
xnor U8129 (N_8129,N_7840,N_7665);
nor U8130 (N_8130,N_7698,N_7601);
nand U8131 (N_8131,N_7984,N_7995);
and U8132 (N_8132,N_7820,N_7506);
nand U8133 (N_8133,N_7912,N_7901);
and U8134 (N_8134,N_7552,N_7993);
xnor U8135 (N_8135,N_7897,N_7836);
or U8136 (N_8136,N_7972,N_7604);
nand U8137 (N_8137,N_7864,N_7917);
and U8138 (N_8138,N_7955,N_7900);
or U8139 (N_8139,N_7891,N_7718);
nor U8140 (N_8140,N_7761,N_7624);
nand U8141 (N_8141,N_7894,N_7930);
nand U8142 (N_8142,N_7965,N_7509);
and U8143 (N_8143,N_7565,N_7714);
nand U8144 (N_8144,N_7708,N_7925);
nor U8145 (N_8145,N_7813,N_7759);
nand U8146 (N_8146,N_7629,N_7747);
or U8147 (N_8147,N_7707,N_7586);
nand U8148 (N_8148,N_7914,N_7768);
nor U8149 (N_8149,N_7627,N_7711);
and U8150 (N_8150,N_7672,N_7839);
xor U8151 (N_8151,N_7838,N_7547);
or U8152 (N_8152,N_7656,N_7736);
nor U8153 (N_8153,N_7877,N_7744);
nand U8154 (N_8154,N_7566,N_7534);
and U8155 (N_8155,N_7713,N_7998);
and U8156 (N_8156,N_7904,N_7816);
nand U8157 (N_8157,N_7852,N_7756);
and U8158 (N_8158,N_7659,N_7598);
nor U8159 (N_8159,N_7631,N_7876);
nor U8160 (N_8160,N_7523,N_7526);
nor U8161 (N_8161,N_7646,N_7760);
and U8162 (N_8162,N_7956,N_7920);
xor U8163 (N_8163,N_7578,N_7520);
nor U8164 (N_8164,N_7553,N_7873);
xnor U8165 (N_8165,N_7908,N_7675);
xnor U8166 (N_8166,N_7579,N_7591);
and U8167 (N_8167,N_7660,N_7542);
or U8168 (N_8168,N_7829,N_7830);
and U8169 (N_8169,N_7936,N_7940);
xor U8170 (N_8170,N_7603,N_7615);
nand U8171 (N_8171,N_7924,N_7671);
and U8172 (N_8172,N_7893,N_7690);
nor U8173 (N_8173,N_7688,N_7882);
or U8174 (N_8174,N_7997,N_7951);
nand U8175 (N_8175,N_7712,N_7738);
xnor U8176 (N_8176,N_7790,N_7746);
nand U8177 (N_8177,N_7902,N_7804);
and U8178 (N_8178,N_7693,N_7650);
nor U8179 (N_8179,N_7950,N_7703);
and U8180 (N_8180,N_7503,N_7825);
or U8181 (N_8181,N_7860,N_7784);
nand U8182 (N_8182,N_7819,N_7765);
nand U8183 (N_8183,N_7888,N_7931);
xnor U8184 (N_8184,N_7573,N_7787);
or U8185 (N_8185,N_7524,N_7758);
and U8186 (N_8186,N_7817,N_7881);
or U8187 (N_8187,N_7887,N_7971);
xor U8188 (N_8188,N_7678,N_7623);
and U8189 (N_8189,N_7821,N_7527);
or U8190 (N_8190,N_7764,N_7782);
and U8191 (N_8191,N_7811,N_7953);
nor U8192 (N_8192,N_7536,N_7981);
nand U8193 (N_8193,N_7986,N_7834);
or U8194 (N_8194,N_7673,N_7584);
nor U8195 (N_8195,N_7640,N_7574);
nor U8196 (N_8196,N_7734,N_7808);
nand U8197 (N_8197,N_7846,N_7871);
xor U8198 (N_8198,N_7781,N_7505);
nand U8199 (N_8199,N_7637,N_7791);
xor U8200 (N_8200,N_7833,N_7583);
and U8201 (N_8201,N_7727,N_7932);
and U8202 (N_8202,N_7968,N_7620);
nand U8203 (N_8203,N_7769,N_7662);
or U8204 (N_8204,N_7960,N_7595);
and U8205 (N_8205,N_7661,N_7980);
nand U8206 (N_8206,N_7994,N_7508);
nor U8207 (N_8207,N_7740,N_7528);
nor U8208 (N_8208,N_7991,N_7798);
and U8209 (N_8209,N_7731,N_7910);
xnor U8210 (N_8210,N_7859,N_7919);
nand U8211 (N_8211,N_7538,N_7611);
xnor U8212 (N_8212,N_7977,N_7913);
nor U8213 (N_8213,N_7973,N_7630);
nand U8214 (N_8214,N_7512,N_7590);
or U8215 (N_8215,N_7625,N_7643);
nor U8216 (N_8216,N_7979,N_7622);
xnor U8217 (N_8217,N_7966,N_7745);
and U8218 (N_8218,N_7531,N_7633);
nand U8219 (N_8219,N_7780,N_7599);
nor U8220 (N_8220,N_7642,N_7571);
nor U8221 (N_8221,N_7954,N_7976);
nand U8222 (N_8222,N_7504,N_7921);
and U8223 (N_8223,N_7890,N_7561);
and U8224 (N_8224,N_7922,N_7733);
nand U8225 (N_8225,N_7772,N_7695);
nor U8226 (N_8226,N_7927,N_7861);
nor U8227 (N_8227,N_7992,N_7537);
or U8228 (N_8228,N_7941,N_7885);
nor U8229 (N_8229,N_7799,N_7720);
or U8230 (N_8230,N_7748,N_7879);
nor U8231 (N_8231,N_7562,N_7616);
nand U8232 (N_8232,N_7918,N_7709);
or U8233 (N_8233,N_7639,N_7801);
and U8234 (N_8234,N_7963,N_7903);
and U8235 (N_8235,N_7664,N_7728);
xnor U8236 (N_8236,N_7569,N_7766);
nand U8237 (N_8237,N_7952,N_7854);
nor U8238 (N_8238,N_7946,N_7741);
or U8239 (N_8239,N_7529,N_7783);
xnor U8240 (N_8240,N_7942,N_7975);
nand U8241 (N_8241,N_7614,N_7828);
nand U8242 (N_8242,N_7757,N_7983);
xnor U8243 (N_8243,N_7739,N_7926);
nand U8244 (N_8244,N_7851,N_7803);
nor U8245 (N_8245,N_7585,N_7753);
xor U8246 (N_8246,N_7636,N_7522);
nand U8247 (N_8247,N_7519,N_7866);
nand U8248 (N_8248,N_7559,N_7644);
or U8249 (N_8249,N_7771,N_7933);
and U8250 (N_8250,N_7554,N_7522);
nor U8251 (N_8251,N_7912,N_7515);
or U8252 (N_8252,N_7566,N_7726);
or U8253 (N_8253,N_7633,N_7893);
nand U8254 (N_8254,N_7840,N_7908);
and U8255 (N_8255,N_7656,N_7606);
nor U8256 (N_8256,N_7995,N_7952);
nor U8257 (N_8257,N_7527,N_7704);
or U8258 (N_8258,N_7871,N_7808);
or U8259 (N_8259,N_7642,N_7719);
or U8260 (N_8260,N_7584,N_7868);
nand U8261 (N_8261,N_7800,N_7504);
xor U8262 (N_8262,N_7836,N_7622);
nor U8263 (N_8263,N_7642,N_7754);
or U8264 (N_8264,N_7597,N_7630);
or U8265 (N_8265,N_7934,N_7910);
nand U8266 (N_8266,N_7732,N_7671);
and U8267 (N_8267,N_7837,N_7716);
nor U8268 (N_8268,N_7680,N_7827);
nor U8269 (N_8269,N_7667,N_7754);
nor U8270 (N_8270,N_7536,N_7977);
or U8271 (N_8271,N_7759,N_7744);
nand U8272 (N_8272,N_7783,N_7875);
nor U8273 (N_8273,N_7970,N_7547);
nor U8274 (N_8274,N_7735,N_7681);
nor U8275 (N_8275,N_7811,N_7864);
or U8276 (N_8276,N_7757,N_7614);
nor U8277 (N_8277,N_7534,N_7823);
and U8278 (N_8278,N_7545,N_7863);
nor U8279 (N_8279,N_7555,N_7500);
and U8280 (N_8280,N_7598,N_7940);
nor U8281 (N_8281,N_7558,N_7794);
or U8282 (N_8282,N_7544,N_7970);
nand U8283 (N_8283,N_7688,N_7894);
nor U8284 (N_8284,N_7967,N_7886);
and U8285 (N_8285,N_7868,N_7926);
or U8286 (N_8286,N_7547,N_7693);
nor U8287 (N_8287,N_7505,N_7562);
nor U8288 (N_8288,N_7965,N_7696);
xnor U8289 (N_8289,N_7681,N_7709);
xor U8290 (N_8290,N_7659,N_7925);
xor U8291 (N_8291,N_7724,N_7766);
or U8292 (N_8292,N_7618,N_7621);
xor U8293 (N_8293,N_7694,N_7510);
or U8294 (N_8294,N_7573,N_7550);
xor U8295 (N_8295,N_7886,N_7572);
nor U8296 (N_8296,N_7570,N_7686);
nand U8297 (N_8297,N_7576,N_7741);
nor U8298 (N_8298,N_7844,N_7766);
xor U8299 (N_8299,N_7572,N_7990);
and U8300 (N_8300,N_7524,N_7979);
nand U8301 (N_8301,N_7722,N_7695);
and U8302 (N_8302,N_7840,N_7992);
xor U8303 (N_8303,N_7936,N_7610);
and U8304 (N_8304,N_7868,N_7624);
nor U8305 (N_8305,N_7761,N_7800);
nand U8306 (N_8306,N_7513,N_7954);
xor U8307 (N_8307,N_7701,N_7616);
and U8308 (N_8308,N_7939,N_7542);
and U8309 (N_8309,N_7762,N_7623);
or U8310 (N_8310,N_7703,N_7534);
nand U8311 (N_8311,N_7844,N_7807);
nor U8312 (N_8312,N_7830,N_7892);
and U8313 (N_8313,N_7831,N_7813);
nor U8314 (N_8314,N_7739,N_7544);
nor U8315 (N_8315,N_7610,N_7825);
nand U8316 (N_8316,N_7543,N_7712);
and U8317 (N_8317,N_7776,N_7882);
xor U8318 (N_8318,N_7824,N_7676);
nor U8319 (N_8319,N_7831,N_7698);
nand U8320 (N_8320,N_7847,N_7808);
and U8321 (N_8321,N_7926,N_7769);
xor U8322 (N_8322,N_7837,N_7685);
xnor U8323 (N_8323,N_7957,N_7882);
nor U8324 (N_8324,N_7591,N_7972);
and U8325 (N_8325,N_7867,N_7832);
or U8326 (N_8326,N_7610,N_7970);
nand U8327 (N_8327,N_7778,N_7600);
nand U8328 (N_8328,N_7781,N_7938);
or U8329 (N_8329,N_7722,N_7667);
or U8330 (N_8330,N_7820,N_7813);
xor U8331 (N_8331,N_7656,N_7636);
and U8332 (N_8332,N_7549,N_7527);
xnor U8333 (N_8333,N_7803,N_7870);
nor U8334 (N_8334,N_7914,N_7922);
xor U8335 (N_8335,N_7914,N_7874);
nand U8336 (N_8336,N_7511,N_7642);
nand U8337 (N_8337,N_7905,N_7701);
nor U8338 (N_8338,N_7952,N_7745);
xnor U8339 (N_8339,N_7612,N_7773);
or U8340 (N_8340,N_7819,N_7643);
xnor U8341 (N_8341,N_7957,N_7603);
nand U8342 (N_8342,N_7683,N_7797);
xnor U8343 (N_8343,N_7623,N_7939);
and U8344 (N_8344,N_7648,N_7698);
nor U8345 (N_8345,N_7511,N_7889);
nand U8346 (N_8346,N_7777,N_7521);
nor U8347 (N_8347,N_7651,N_7694);
and U8348 (N_8348,N_7651,N_7754);
xnor U8349 (N_8349,N_7978,N_7733);
nor U8350 (N_8350,N_7813,N_7819);
and U8351 (N_8351,N_7706,N_7814);
and U8352 (N_8352,N_7911,N_7678);
xnor U8353 (N_8353,N_7762,N_7640);
nor U8354 (N_8354,N_7793,N_7526);
nand U8355 (N_8355,N_7838,N_7687);
xnor U8356 (N_8356,N_7973,N_7701);
xnor U8357 (N_8357,N_7542,N_7501);
xnor U8358 (N_8358,N_7714,N_7859);
nand U8359 (N_8359,N_7540,N_7552);
xor U8360 (N_8360,N_7748,N_7910);
xor U8361 (N_8361,N_7598,N_7987);
or U8362 (N_8362,N_7815,N_7687);
and U8363 (N_8363,N_7797,N_7933);
nor U8364 (N_8364,N_7753,N_7660);
nor U8365 (N_8365,N_7728,N_7869);
or U8366 (N_8366,N_7656,N_7810);
and U8367 (N_8367,N_7537,N_7866);
and U8368 (N_8368,N_7892,N_7931);
nand U8369 (N_8369,N_7959,N_7807);
nand U8370 (N_8370,N_7989,N_7986);
nand U8371 (N_8371,N_7895,N_7811);
nand U8372 (N_8372,N_7661,N_7863);
xnor U8373 (N_8373,N_7921,N_7810);
nand U8374 (N_8374,N_7846,N_7872);
xnor U8375 (N_8375,N_7826,N_7799);
xor U8376 (N_8376,N_7713,N_7682);
nand U8377 (N_8377,N_7861,N_7737);
or U8378 (N_8378,N_7762,N_7693);
nand U8379 (N_8379,N_7768,N_7763);
nand U8380 (N_8380,N_7526,N_7912);
nor U8381 (N_8381,N_7633,N_7935);
and U8382 (N_8382,N_7971,N_7857);
nor U8383 (N_8383,N_7926,N_7664);
nor U8384 (N_8384,N_7669,N_7578);
nand U8385 (N_8385,N_7611,N_7652);
nand U8386 (N_8386,N_7534,N_7973);
nand U8387 (N_8387,N_7579,N_7815);
nor U8388 (N_8388,N_7770,N_7771);
xnor U8389 (N_8389,N_7843,N_7744);
nor U8390 (N_8390,N_7590,N_7547);
or U8391 (N_8391,N_7873,N_7596);
or U8392 (N_8392,N_7533,N_7807);
nand U8393 (N_8393,N_7739,N_7676);
nand U8394 (N_8394,N_7979,N_7907);
nor U8395 (N_8395,N_7633,N_7922);
and U8396 (N_8396,N_7540,N_7787);
nor U8397 (N_8397,N_7837,N_7521);
or U8398 (N_8398,N_7789,N_7904);
xnor U8399 (N_8399,N_7880,N_7510);
and U8400 (N_8400,N_7774,N_7604);
nand U8401 (N_8401,N_7901,N_7508);
nor U8402 (N_8402,N_7509,N_7991);
nor U8403 (N_8403,N_7826,N_7703);
or U8404 (N_8404,N_7866,N_7653);
and U8405 (N_8405,N_7565,N_7507);
or U8406 (N_8406,N_7829,N_7843);
nand U8407 (N_8407,N_7958,N_7813);
nand U8408 (N_8408,N_7832,N_7740);
and U8409 (N_8409,N_7852,N_7609);
and U8410 (N_8410,N_7820,N_7950);
nand U8411 (N_8411,N_7815,N_7784);
nand U8412 (N_8412,N_7774,N_7790);
and U8413 (N_8413,N_7784,N_7851);
and U8414 (N_8414,N_7682,N_7525);
xnor U8415 (N_8415,N_7784,N_7752);
nand U8416 (N_8416,N_7976,N_7781);
and U8417 (N_8417,N_7854,N_7549);
xnor U8418 (N_8418,N_7838,N_7791);
or U8419 (N_8419,N_7916,N_7750);
xor U8420 (N_8420,N_7723,N_7580);
and U8421 (N_8421,N_7721,N_7886);
nor U8422 (N_8422,N_7601,N_7904);
nor U8423 (N_8423,N_7945,N_7743);
nand U8424 (N_8424,N_7997,N_7781);
xor U8425 (N_8425,N_7772,N_7657);
nand U8426 (N_8426,N_7773,N_7851);
or U8427 (N_8427,N_7600,N_7584);
and U8428 (N_8428,N_7658,N_7950);
nor U8429 (N_8429,N_7937,N_7612);
nor U8430 (N_8430,N_7542,N_7908);
or U8431 (N_8431,N_7721,N_7962);
xnor U8432 (N_8432,N_7662,N_7834);
and U8433 (N_8433,N_7643,N_7950);
and U8434 (N_8434,N_7705,N_7902);
xnor U8435 (N_8435,N_7860,N_7914);
nand U8436 (N_8436,N_7698,N_7650);
nand U8437 (N_8437,N_7849,N_7809);
xnor U8438 (N_8438,N_7566,N_7890);
or U8439 (N_8439,N_7723,N_7559);
or U8440 (N_8440,N_7739,N_7917);
xor U8441 (N_8441,N_7630,N_7960);
xor U8442 (N_8442,N_7517,N_7593);
nand U8443 (N_8443,N_7943,N_7933);
or U8444 (N_8444,N_7611,N_7891);
and U8445 (N_8445,N_7902,N_7589);
nor U8446 (N_8446,N_7643,N_7824);
nor U8447 (N_8447,N_7956,N_7625);
xnor U8448 (N_8448,N_7637,N_7952);
nor U8449 (N_8449,N_7584,N_7677);
nor U8450 (N_8450,N_7727,N_7970);
or U8451 (N_8451,N_7538,N_7669);
or U8452 (N_8452,N_7789,N_7962);
nand U8453 (N_8453,N_7725,N_7540);
nand U8454 (N_8454,N_7606,N_7702);
xnor U8455 (N_8455,N_7940,N_7862);
xnor U8456 (N_8456,N_7926,N_7841);
and U8457 (N_8457,N_7627,N_7572);
xnor U8458 (N_8458,N_7785,N_7695);
or U8459 (N_8459,N_7616,N_7631);
nand U8460 (N_8460,N_7970,N_7689);
xnor U8461 (N_8461,N_7674,N_7937);
nand U8462 (N_8462,N_7584,N_7505);
or U8463 (N_8463,N_7676,N_7714);
or U8464 (N_8464,N_7832,N_7968);
nand U8465 (N_8465,N_7890,N_7827);
nor U8466 (N_8466,N_7646,N_7717);
or U8467 (N_8467,N_7599,N_7578);
or U8468 (N_8468,N_7652,N_7578);
nor U8469 (N_8469,N_7713,N_7579);
and U8470 (N_8470,N_7627,N_7793);
nand U8471 (N_8471,N_7612,N_7753);
or U8472 (N_8472,N_7667,N_7671);
or U8473 (N_8473,N_7701,N_7718);
xor U8474 (N_8474,N_7519,N_7562);
nor U8475 (N_8475,N_7675,N_7516);
or U8476 (N_8476,N_7540,N_7796);
or U8477 (N_8477,N_7644,N_7758);
xor U8478 (N_8478,N_7986,N_7931);
xor U8479 (N_8479,N_7763,N_7852);
or U8480 (N_8480,N_7827,N_7552);
and U8481 (N_8481,N_7719,N_7981);
xnor U8482 (N_8482,N_7563,N_7567);
or U8483 (N_8483,N_7761,N_7584);
xnor U8484 (N_8484,N_7869,N_7920);
nor U8485 (N_8485,N_7505,N_7860);
nor U8486 (N_8486,N_7819,N_7522);
xnor U8487 (N_8487,N_7814,N_7541);
nand U8488 (N_8488,N_7897,N_7676);
nand U8489 (N_8489,N_7645,N_7586);
nor U8490 (N_8490,N_7860,N_7547);
and U8491 (N_8491,N_7552,N_7931);
xor U8492 (N_8492,N_7827,N_7836);
xnor U8493 (N_8493,N_7687,N_7869);
and U8494 (N_8494,N_7669,N_7587);
xor U8495 (N_8495,N_7518,N_7848);
and U8496 (N_8496,N_7522,N_7718);
or U8497 (N_8497,N_7769,N_7863);
or U8498 (N_8498,N_7698,N_7563);
xnor U8499 (N_8499,N_7640,N_7720);
or U8500 (N_8500,N_8297,N_8436);
nor U8501 (N_8501,N_8053,N_8285);
nor U8502 (N_8502,N_8481,N_8204);
nand U8503 (N_8503,N_8446,N_8465);
or U8504 (N_8504,N_8393,N_8493);
xnor U8505 (N_8505,N_8205,N_8447);
nor U8506 (N_8506,N_8093,N_8098);
xnor U8507 (N_8507,N_8176,N_8486);
and U8508 (N_8508,N_8475,N_8480);
or U8509 (N_8509,N_8333,N_8150);
xor U8510 (N_8510,N_8012,N_8131);
nor U8511 (N_8511,N_8173,N_8077);
nor U8512 (N_8512,N_8491,N_8284);
xor U8513 (N_8513,N_8373,N_8271);
nor U8514 (N_8514,N_8017,N_8055);
nand U8515 (N_8515,N_8001,N_8312);
or U8516 (N_8516,N_8223,N_8437);
nor U8517 (N_8517,N_8387,N_8018);
xnor U8518 (N_8518,N_8392,N_8498);
and U8519 (N_8519,N_8172,N_8209);
nand U8520 (N_8520,N_8303,N_8453);
or U8521 (N_8521,N_8352,N_8423);
xnor U8522 (N_8522,N_8109,N_8169);
xnor U8523 (N_8523,N_8319,N_8372);
nand U8524 (N_8524,N_8234,N_8263);
xor U8525 (N_8525,N_8376,N_8039);
nand U8526 (N_8526,N_8015,N_8395);
nand U8527 (N_8527,N_8167,N_8132);
nor U8528 (N_8528,N_8351,N_8243);
and U8529 (N_8529,N_8092,N_8033);
nor U8530 (N_8530,N_8404,N_8435);
and U8531 (N_8531,N_8200,N_8381);
xnor U8532 (N_8532,N_8145,N_8127);
and U8533 (N_8533,N_8218,N_8334);
and U8534 (N_8534,N_8143,N_8415);
and U8535 (N_8535,N_8264,N_8308);
nor U8536 (N_8536,N_8118,N_8377);
nor U8537 (N_8537,N_8097,N_8121);
nor U8538 (N_8538,N_8464,N_8443);
nor U8539 (N_8539,N_8311,N_8224);
or U8540 (N_8540,N_8065,N_8043);
xor U8541 (N_8541,N_8175,N_8003);
and U8542 (N_8542,N_8256,N_8170);
xnor U8543 (N_8543,N_8215,N_8379);
xnor U8544 (N_8544,N_8119,N_8096);
or U8545 (N_8545,N_8448,N_8081);
xnor U8546 (N_8546,N_8487,N_8482);
nand U8547 (N_8547,N_8116,N_8108);
and U8548 (N_8548,N_8348,N_8146);
nand U8549 (N_8549,N_8191,N_8196);
and U8550 (N_8550,N_8391,N_8009);
and U8551 (N_8551,N_8469,N_8231);
and U8552 (N_8552,N_8032,N_8104);
nand U8553 (N_8553,N_8149,N_8038);
nor U8554 (N_8554,N_8408,N_8247);
and U8555 (N_8555,N_8484,N_8051);
nor U8556 (N_8556,N_8367,N_8432);
xor U8557 (N_8557,N_8346,N_8087);
and U8558 (N_8558,N_8076,N_8088);
nor U8559 (N_8559,N_8291,N_8183);
nor U8560 (N_8560,N_8229,N_8279);
nor U8561 (N_8561,N_8318,N_8383);
or U8562 (N_8562,N_8139,N_8058);
xnor U8563 (N_8563,N_8124,N_8439);
nand U8564 (N_8564,N_8363,N_8474);
nand U8565 (N_8565,N_8241,N_8298);
nor U8566 (N_8566,N_8057,N_8222);
nor U8567 (N_8567,N_8296,N_8197);
xor U8568 (N_8568,N_8248,N_8180);
nand U8569 (N_8569,N_8240,N_8134);
nor U8570 (N_8570,N_8011,N_8130);
or U8571 (N_8571,N_8337,N_8460);
xor U8572 (N_8572,N_8328,N_8343);
nor U8573 (N_8573,N_8302,N_8013);
or U8574 (N_8574,N_8091,N_8049);
nor U8575 (N_8575,N_8041,N_8478);
nor U8576 (N_8576,N_8473,N_8008);
or U8577 (N_8577,N_8147,N_8181);
nor U8578 (N_8578,N_8035,N_8410);
nor U8579 (N_8579,N_8067,N_8470);
xnor U8580 (N_8580,N_8140,N_8288);
or U8581 (N_8581,N_8115,N_8389);
nand U8582 (N_8582,N_8066,N_8450);
nand U8583 (N_8583,N_8358,N_8061);
nor U8584 (N_8584,N_8133,N_8398);
xnor U8585 (N_8585,N_8195,N_8340);
nand U8586 (N_8586,N_8177,N_8314);
xnor U8587 (N_8587,N_8239,N_8322);
or U8588 (N_8588,N_8135,N_8186);
nand U8589 (N_8589,N_8022,N_8158);
or U8590 (N_8590,N_8471,N_8216);
xor U8591 (N_8591,N_8370,N_8299);
nand U8592 (N_8592,N_8499,N_8293);
and U8593 (N_8593,N_8152,N_8380);
or U8594 (N_8594,N_8037,N_8427);
and U8595 (N_8595,N_8048,N_8111);
or U8596 (N_8596,N_8384,N_8028);
xor U8597 (N_8597,N_8403,N_8361);
and U8598 (N_8598,N_8212,N_8286);
and U8599 (N_8599,N_8168,N_8341);
nor U8600 (N_8600,N_8120,N_8014);
and U8601 (N_8601,N_8227,N_8294);
xnor U8602 (N_8602,N_8153,N_8230);
xnor U8603 (N_8603,N_8488,N_8267);
nand U8604 (N_8604,N_8163,N_8306);
and U8605 (N_8605,N_8242,N_8084);
nand U8606 (N_8606,N_8203,N_8046);
and U8607 (N_8607,N_8074,N_8005);
nand U8608 (N_8608,N_8188,N_8010);
xor U8609 (N_8609,N_8266,N_8290);
xor U8610 (N_8610,N_8193,N_8187);
xor U8611 (N_8611,N_8324,N_8102);
nand U8612 (N_8612,N_8253,N_8273);
xnor U8613 (N_8613,N_8416,N_8394);
and U8614 (N_8614,N_8232,N_8354);
xor U8615 (N_8615,N_8162,N_8295);
and U8616 (N_8616,N_8344,N_8262);
nor U8617 (N_8617,N_8356,N_8040);
and U8618 (N_8618,N_8458,N_8495);
nand U8619 (N_8619,N_8249,N_8357);
xnor U8620 (N_8620,N_8114,N_8326);
nand U8621 (N_8621,N_8030,N_8476);
or U8622 (N_8622,N_8171,N_8086);
nor U8623 (N_8623,N_8424,N_8494);
and U8624 (N_8624,N_8252,N_8325);
or U8625 (N_8625,N_8259,N_8029);
and U8626 (N_8626,N_8479,N_8113);
xor U8627 (N_8627,N_8430,N_8422);
and U8628 (N_8628,N_8406,N_8129);
xor U8629 (N_8629,N_8100,N_8433);
xnor U8630 (N_8630,N_8221,N_8059);
nand U8631 (N_8631,N_8156,N_8411);
or U8632 (N_8632,N_8160,N_8440);
or U8633 (N_8633,N_8004,N_8069);
nand U8634 (N_8634,N_8428,N_8060);
or U8635 (N_8635,N_8278,N_8345);
nand U8636 (N_8636,N_8441,N_8456);
nor U8637 (N_8637,N_8207,N_8413);
nand U8638 (N_8638,N_8332,N_8414);
nand U8639 (N_8639,N_8025,N_8457);
nand U8640 (N_8640,N_8185,N_8396);
nand U8641 (N_8641,N_8485,N_8402);
nand U8642 (N_8642,N_8202,N_8117);
nor U8643 (N_8643,N_8154,N_8375);
and U8644 (N_8644,N_8075,N_8155);
nand U8645 (N_8645,N_8101,N_8031);
and U8646 (N_8646,N_8492,N_8412);
nor U8647 (N_8647,N_8426,N_8429);
nor U8648 (N_8648,N_8136,N_8161);
or U8649 (N_8649,N_8251,N_8257);
and U8650 (N_8650,N_8421,N_8021);
xor U8651 (N_8651,N_8378,N_8246);
xnor U8652 (N_8652,N_8417,N_8420);
nor U8653 (N_8653,N_8148,N_8225);
nand U8654 (N_8654,N_8276,N_8006);
xnor U8655 (N_8655,N_8250,N_8366);
and U8656 (N_8656,N_8407,N_8489);
xor U8657 (N_8657,N_8362,N_8477);
xnor U8658 (N_8658,N_8142,N_8144);
nand U8659 (N_8659,N_8268,N_8459);
or U8660 (N_8660,N_8419,N_8050);
or U8661 (N_8661,N_8463,N_8444);
nand U8662 (N_8662,N_8269,N_8374);
or U8663 (N_8663,N_8027,N_8189);
xnor U8664 (N_8664,N_8305,N_8355);
nand U8665 (N_8665,N_8137,N_8401);
nand U8666 (N_8666,N_8054,N_8369);
nor U8667 (N_8667,N_8452,N_8063);
nand U8668 (N_8668,N_8388,N_8281);
and U8669 (N_8669,N_8068,N_8199);
and U8670 (N_8670,N_8339,N_8327);
or U8671 (N_8671,N_8182,N_8034);
and U8672 (N_8672,N_8036,N_8198);
or U8673 (N_8673,N_8386,N_8128);
nand U8674 (N_8674,N_8347,N_8206);
and U8675 (N_8675,N_8090,N_8238);
nor U8676 (N_8676,N_8409,N_8258);
xor U8677 (N_8677,N_8461,N_8072);
or U8678 (N_8678,N_8174,N_8434);
and U8679 (N_8679,N_8110,N_8235);
and U8680 (N_8680,N_8157,N_8184);
nand U8681 (N_8681,N_8016,N_8236);
and U8682 (N_8682,N_8254,N_8304);
nand U8683 (N_8683,N_8213,N_8201);
or U8684 (N_8684,N_8282,N_8315);
xor U8685 (N_8685,N_8399,N_8083);
nor U8686 (N_8686,N_8042,N_8192);
or U8687 (N_8687,N_8277,N_8126);
or U8688 (N_8688,N_8064,N_8385);
nor U8689 (N_8689,N_8287,N_8071);
nor U8690 (N_8690,N_8107,N_8244);
nand U8691 (N_8691,N_8451,N_8310);
nor U8692 (N_8692,N_8497,N_8316);
xnor U8693 (N_8693,N_8194,N_8047);
nand U8694 (N_8694,N_8329,N_8467);
or U8695 (N_8695,N_8211,N_8044);
nand U8696 (N_8696,N_8080,N_8125);
or U8697 (N_8697,N_8237,N_8317);
nand U8698 (N_8698,N_8122,N_8445);
nor U8699 (N_8699,N_8289,N_8070);
and U8700 (N_8700,N_8472,N_8165);
or U8701 (N_8701,N_8026,N_8313);
xnor U8702 (N_8702,N_8007,N_8056);
and U8703 (N_8703,N_8292,N_8082);
and U8704 (N_8704,N_8438,N_8261);
xor U8705 (N_8705,N_8353,N_8260);
and U8706 (N_8706,N_8190,N_8159);
or U8707 (N_8707,N_8307,N_8309);
nor U8708 (N_8708,N_8272,N_8335);
nand U8709 (N_8709,N_8219,N_8265);
nor U8710 (N_8710,N_8364,N_8217);
nand U8711 (N_8711,N_8208,N_8331);
nor U8712 (N_8712,N_8442,N_8228);
or U8713 (N_8713,N_8255,N_8466);
and U8714 (N_8714,N_8179,N_8079);
or U8715 (N_8715,N_8359,N_8123);
and U8716 (N_8716,N_8073,N_8085);
nand U8717 (N_8717,N_8320,N_8233);
and U8718 (N_8718,N_8368,N_8095);
xnor U8719 (N_8719,N_8178,N_8210);
and U8720 (N_8720,N_8323,N_8338);
nand U8721 (N_8721,N_8089,N_8141);
or U8722 (N_8722,N_8301,N_8321);
nand U8723 (N_8723,N_8300,N_8226);
nor U8724 (N_8724,N_8000,N_8283);
nor U8725 (N_8725,N_8024,N_8496);
nor U8726 (N_8726,N_8002,N_8468);
or U8727 (N_8727,N_8103,N_8405);
xor U8728 (N_8728,N_8349,N_8045);
nand U8729 (N_8729,N_8099,N_8275);
nor U8730 (N_8730,N_8330,N_8455);
and U8731 (N_8731,N_8214,N_8138);
nand U8732 (N_8732,N_8164,N_8270);
xor U8733 (N_8733,N_8454,N_8020);
and U8734 (N_8734,N_8350,N_8462);
nor U8735 (N_8735,N_8105,N_8425);
nor U8736 (N_8736,N_8418,N_8336);
or U8737 (N_8737,N_8365,N_8371);
xor U8738 (N_8738,N_8245,N_8397);
nand U8739 (N_8739,N_8019,N_8106);
nor U8740 (N_8740,N_8023,N_8078);
and U8741 (N_8741,N_8390,N_8431);
or U8742 (N_8742,N_8052,N_8280);
and U8743 (N_8743,N_8490,N_8360);
or U8744 (N_8744,N_8112,N_8382);
nand U8745 (N_8745,N_8274,N_8342);
or U8746 (N_8746,N_8166,N_8483);
nand U8747 (N_8747,N_8151,N_8400);
nand U8748 (N_8748,N_8449,N_8062);
or U8749 (N_8749,N_8094,N_8220);
or U8750 (N_8750,N_8166,N_8449);
nand U8751 (N_8751,N_8305,N_8101);
or U8752 (N_8752,N_8014,N_8253);
nor U8753 (N_8753,N_8070,N_8032);
nand U8754 (N_8754,N_8072,N_8124);
and U8755 (N_8755,N_8439,N_8011);
nand U8756 (N_8756,N_8318,N_8305);
xnor U8757 (N_8757,N_8207,N_8040);
or U8758 (N_8758,N_8170,N_8270);
nand U8759 (N_8759,N_8193,N_8218);
xor U8760 (N_8760,N_8465,N_8469);
or U8761 (N_8761,N_8133,N_8126);
nand U8762 (N_8762,N_8371,N_8437);
nor U8763 (N_8763,N_8173,N_8273);
nor U8764 (N_8764,N_8354,N_8188);
xnor U8765 (N_8765,N_8004,N_8310);
or U8766 (N_8766,N_8288,N_8173);
and U8767 (N_8767,N_8394,N_8400);
or U8768 (N_8768,N_8030,N_8135);
and U8769 (N_8769,N_8229,N_8061);
xnor U8770 (N_8770,N_8123,N_8179);
and U8771 (N_8771,N_8458,N_8194);
nor U8772 (N_8772,N_8064,N_8259);
nand U8773 (N_8773,N_8460,N_8069);
nand U8774 (N_8774,N_8352,N_8406);
xor U8775 (N_8775,N_8126,N_8074);
xnor U8776 (N_8776,N_8096,N_8197);
xor U8777 (N_8777,N_8445,N_8463);
nand U8778 (N_8778,N_8126,N_8060);
or U8779 (N_8779,N_8290,N_8080);
nand U8780 (N_8780,N_8231,N_8120);
and U8781 (N_8781,N_8356,N_8041);
nor U8782 (N_8782,N_8283,N_8410);
and U8783 (N_8783,N_8188,N_8493);
nor U8784 (N_8784,N_8271,N_8126);
and U8785 (N_8785,N_8383,N_8258);
nor U8786 (N_8786,N_8042,N_8108);
and U8787 (N_8787,N_8115,N_8369);
or U8788 (N_8788,N_8278,N_8256);
nor U8789 (N_8789,N_8211,N_8315);
xnor U8790 (N_8790,N_8259,N_8088);
and U8791 (N_8791,N_8497,N_8056);
nor U8792 (N_8792,N_8448,N_8497);
or U8793 (N_8793,N_8478,N_8260);
xor U8794 (N_8794,N_8153,N_8253);
and U8795 (N_8795,N_8407,N_8060);
nor U8796 (N_8796,N_8021,N_8239);
and U8797 (N_8797,N_8160,N_8435);
nand U8798 (N_8798,N_8220,N_8299);
nor U8799 (N_8799,N_8227,N_8266);
and U8800 (N_8800,N_8308,N_8004);
nor U8801 (N_8801,N_8369,N_8093);
nor U8802 (N_8802,N_8400,N_8425);
or U8803 (N_8803,N_8152,N_8317);
nor U8804 (N_8804,N_8367,N_8364);
and U8805 (N_8805,N_8234,N_8061);
and U8806 (N_8806,N_8102,N_8008);
or U8807 (N_8807,N_8383,N_8075);
and U8808 (N_8808,N_8380,N_8162);
nand U8809 (N_8809,N_8321,N_8247);
xor U8810 (N_8810,N_8160,N_8100);
and U8811 (N_8811,N_8072,N_8168);
or U8812 (N_8812,N_8416,N_8193);
xor U8813 (N_8813,N_8300,N_8490);
nand U8814 (N_8814,N_8086,N_8121);
nand U8815 (N_8815,N_8250,N_8018);
nor U8816 (N_8816,N_8164,N_8058);
nor U8817 (N_8817,N_8489,N_8401);
nand U8818 (N_8818,N_8302,N_8454);
xnor U8819 (N_8819,N_8228,N_8213);
nor U8820 (N_8820,N_8023,N_8293);
or U8821 (N_8821,N_8382,N_8134);
nor U8822 (N_8822,N_8361,N_8379);
nor U8823 (N_8823,N_8477,N_8328);
nand U8824 (N_8824,N_8156,N_8478);
nand U8825 (N_8825,N_8157,N_8153);
and U8826 (N_8826,N_8293,N_8446);
and U8827 (N_8827,N_8118,N_8081);
and U8828 (N_8828,N_8318,N_8450);
and U8829 (N_8829,N_8104,N_8108);
xor U8830 (N_8830,N_8364,N_8416);
nor U8831 (N_8831,N_8113,N_8330);
and U8832 (N_8832,N_8242,N_8272);
nor U8833 (N_8833,N_8145,N_8208);
nor U8834 (N_8834,N_8383,N_8411);
and U8835 (N_8835,N_8471,N_8441);
nor U8836 (N_8836,N_8035,N_8264);
or U8837 (N_8837,N_8108,N_8409);
nand U8838 (N_8838,N_8427,N_8371);
or U8839 (N_8839,N_8487,N_8415);
or U8840 (N_8840,N_8338,N_8388);
nand U8841 (N_8841,N_8448,N_8174);
nand U8842 (N_8842,N_8194,N_8395);
or U8843 (N_8843,N_8455,N_8122);
xor U8844 (N_8844,N_8099,N_8186);
nand U8845 (N_8845,N_8186,N_8347);
nand U8846 (N_8846,N_8354,N_8071);
nor U8847 (N_8847,N_8012,N_8116);
or U8848 (N_8848,N_8093,N_8023);
or U8849 (N_8849,N_8048,N_8287);
and U8850 (N_8850,N_8040,N_8002);
nand U8851 (N_8851,N_8345,N_8095);
nor U8852 (N_8852,N_8006,N_8248);
nand U8853 (N_8853,N_8295,N_8056);
xor U8854 (N_8854,N_8321,N_8329);
or U8855 (N_8855,N_8000,N_8232);
nor U8856 (N_8856,N_8283,N_8015);
xnor U8857 (N_8857,N_8083,N_8328);
nor U8858 (N_8858,N_8464,N_8025);
or U8859 (N_8859,N_8434,N_8226);
and U8860 (N_8860,N_8376,N_8497);
and U8861 (N_8861,N_8076,N_8450);
xor U8862 (N_8862,N_8246,N_8273);
nor U8863 (N_8863,N_8348,N_8451);
nand U8864 (N_8864,N_8385,N_8438);
xnor U8865 (N_8865,N_8252,N_8300);
xor U8866 (N_8866,N_8127,N_8074);
or U8867 (N_8867,N_8340,N_8368);
nor U8868 (N_8868,N_8193,N_8054);
and U8869 (N_8869,N_8210,N_8352);
nand U8870 (N_8870,N_8347,N_8239);
nor U8871 (N_8871,N_8100,N_8180);
nand U8872 (N_8872,N_8454,N_8292);
nor U8873 (N_8873,N_8428,N_8347);
or U8874 (N_8874,N_8204,N_8193);
or U8875 (N_8875,N_8061,N_8086);
nand U8876 (N_8876,N_8266,N_8342);
nor U8877 (N_8877,N_8059,N_8341);
xnor U8878 (N_8878,N_8302,N_8052);
and U8879 (N_8879,N_8332,N_8216);
xor U8880 (N_8880,N_8127,N_8014);
and U8881 (N_8881,N_8337,N_8392);
or U8882 (N_8882,N_8094,N_8323);
and U8883 (N_8883,N_8362,N_8092);
xnor U8884 (N_8884,N_8317,N_8262);
and U8885 (N_8885,N_8203,N_8257);
nand U8886 (N_8886,N_8412,N_8259);
xor U8887 (N_8887,N_8240,N_8425);
nand U8888 (N_8888,N_8200,N_8305);
or U8889 (N_8889,N_8193,N_8156);
or U8890 (N_8890,N_8394,N_8238);
or U8891 (N_8891,N_8220,N_8038);
nor U8892 (N_8892,N_8453,N_8073);
and U8893 (N_8893,N_8409,N_8394);
nand U8894 (N_8894,N_8309,N_8329);
or U8895 (N_8895,N_8200,N_8285);
and U8896 (N_8896,N_8247,N_8340);
nor U8897 (N_8897,N_8388,N_8409);
xor U8898 (N_8898,N_8153,N_8181);
nand U8899 (N_8899,N_8299,N_8287);
and U8900 (N_8900,N_8002,N_8406);
or U8901 (N_8901,N_8131,N_8378);
nand U8902 (N_8902,N_8323,N_8034);
or U8903 (N_8903,N_8214,N_8428);
and U8904 (N_8904,N_8165,N_8440);
nand U8905 (N_8905,N_8453,N_8208);
nor U8906 (N_8906,N_8091,N_8433);
or U8907 (N_8907,N_8278,N_8159);
and U8908 (N_8908,N_8012,N_8362);
nand U8909 (N_8909,N_8489,N_8251);
nand U8910 (N_8910,N_8125,N_8124);
nand U8911 (N_8911,N_8348,N_8478);
nand U8912 (N_8912,N_8285,N_8165);
nand U8913 (N_8913,N_8244,N_8037);
or U8914 (N_8914,N_8166,N_8046);
nor U8915 (N_8915,N_8090,N_8358);
xor U8916 (N_8916,N_8056,N_8252);
or U8917 (N_8917,N_8135,N_8078);
and U8918 (N_8918,N_8250,N_8021);
xor U8919 (N_8919,N_8190,N_8316);
nor U8920 (N_8920,N_8056,N_8480);
nor U8921 (N_8921,N_8135,N_8233);
nand U8922 (N_8922,N_8337,N_8161);
and U8923 (N_8923,N_8103,N_8302);
xor U8924 (N_8924,N_8180,N_8283);
and U8925 (N_8925,N_8292,N_8270);
nor U8926 (N_8926,N_8344,N_8072);
and U8927 (N_8927,N_8000,N_8015);
xor U8928 (N_8928,N_8035,N_8110);
and U8929 (N_8929,N_8164,N_8168);
nand U8930 (N_8930,N_8352,N_8493);
nor U8931 (N_8931,N_8106,N_8434);
or U8932 (N_8932,N_8056,N_8149);
and U8933 (N_8933,N_8143,N_8063);
nand U8934 (N_8934,N_8119,N_8069);
xnor U8935 (N_8935,N_8324,N_8409);
or U8936 (N_8936,N_8345,N_8287);
and U8937 (N_8937,N_8158,N_8403);
or U8938 (N_8938,N_8021,N_8006);
nor U8939 (N_8939,N_8367,N_8282);
or U8940 (N_8940,N_8209,N_8141);
nand U8941 (N_8941,N_8271,N_8224);
nand U8942 (N_8942,N_8118,N_8170);
nor U8943 (N_8943,N_8009,N_8184);
and U8944 (N_8944,N_8152,N_8475);
and U8945 (N_8945,N_8297,N_8488);
nand U8946 (N_8946,N_8395,N_8242);
and U8947 (N_8947,N_8148,N_8081);
nor U8948 (N_8948,N_8373,N_8348);
nor U8949 (N_8949,N_8341,N_8027);
nand U8950 (N_8950,N_8332,N_8272);
xor U8951 (N_8951,N_8068,N_8123);
xnor U8952 (N_8952,N_8338,N_8136);
xnor U8953 (N_8953,N_8208,N_8063);
nor U8954 (N_8954,N_8319,N_8198);
or U8955 (N_8955,N_8395,N_8139);
nor U8956 (N_8956,N_8031,N_8361);
and U8957 (N_8957,N_8146,N_8212);
nor U8958 (N_8958,N_8128,N_8122);
or U8959 (N_8959,N_8377,N_8150);
or U8960 (N_8960,N_8090,N_8131);
xnor U8961 (N_8961,N_8212,N_8321);
nor U8962 (N_8962,N_8316,N_8287);
and U8963 (N_8963,N_8103,N_8489);
nand U8964 (N_8964,N_8080,N_8041);
xor U8965 (N_8965,N_8446,N_8046);
nor U8966 (N_8966,N_8066,N_8054);
nor U8967 (N_8967,N_8282,N_8143);
xor U8968 (N_8968,N_8306,N_8313);
nor U8969 (N_8969,N_8043,N_8267);
nand U8970 (N_8970,N_8332,N_8124);
xnor U8971 (N_8971,N_8198,N_8021);
and U8972 (N_8972,N_8091,N_8224);
nor U8973 (N_8973,N_8009,N_8471);
and U8974 (N_8974,N_8119,N_8166);
and U8975 (N_8975,N_8254,N_8073);
xnor U8976 (N_8976,N_8119,N_8085);
xnor U8977 (N_8977,N_8387,N_8239);
nor U8978 (N_8978,N_8426,N_8220);
nand U8979 (N_8979,N_8306,N_8177);
and U8980 (N_8980,N_8442,N_8123);
xnor U8981 (N_8981,N_8422,N_8390);
nand U8982 (N_8982,N_8395,N_8178);
nor U8983 (N_8983,N_8038,N_8147);
or U8984 (N_8984,N_8051,N_8205);
or U8985 (N_8985,N_8246,N_8355);
or U8986 (N_8986,N_8170,N_8438);
xor U8987 (N_8987,N_8409,N_8389);
nor U8988 (N_8988,N_8284,N_8091);
and U8989 (N_8989,N_8034,N_8419);
nand U8990 (N_8990,N_8478,N_8233);
nor U8991 (N_8991,N_8307,N_8484);
or U8992 (N_8992,N_8449,N_8167);
and U8993 (N_8993,N_8422,N_8388);
and U8994 (N_8994,N_8002,N_8095);
or U8995 (N_8995,N_8154,N_8422);
or U8996 (N_8996,N_8328,N_8204);
nor U8997 (N_8997,N_8091,N_8321);
and U8998 (N_8998,N_8212,N_8039);
and U8999 (N_8999,N_8205,N_8409);
nor U9000 (N_9000,N_8548,N_8779);
nand U9001 (N_9001,N_8620,N_8586);
and U9002 (N_9002,N_8964,N_8960);
xor U9003 (N_9003,N_8750,N_8785);
nor U9004 (N_9004,N_8688,N_8886);
nand U9005 (N_9005,N_8690,N_8885);
xnor U9006 (N_9006,N_8868,N_8918);
or U9007 (N_9007,N_8519,N_8741);
nor U9008 (N_9008,N_8603,N_8978);
and U9009 (N_9009,N_8717,N_8854);
nand U9010 (N_9010,N_8710,N_8762);
or U9011 (N_9011,N_8853,N_8666);
nand U9012 (N_9012,N_8569,N_8576);
nor U9013 (N_9013,N_8962,N_8510);
xor U9014 (N_9014,N_8580,N_8830);
nand U9015 (N_9015,N_8752,N_8618);
and U9016 (N_9016,N_8994,N_8869);
nor U9017 (N_9017,N_8973,N_8561);
or U9018 (N_9018,N_8661,N_8524);
nand U9019 (N_9019,N_8835,N_8759);
nand U9020 (N_9020,N_8686,N_8591);
and U9021 (N_9021,N_8725,N_8969);
nor U9022 (N_9022,N_8694,N_8995);
nand U9023 (N_9023,N_8513,N_8906);
and U9024 (N_9024,N_8795,N_8540);
xor U9025 (N_9025,N_8634,N_8874);
or U9026 (N_9026,N_8793,N_8997);
nand U9027 (N_9027,N_8756,N_8588);
nor U9028 (N_9028,N_8640,N_8977);
and U9029 (N_9029,N_8782,N_8593);
xnor U9030 (N_9030,N_8935,N_8972);
nand U9031 (N_9031,N_8776,N_8800);
or U9032 (N_9032,N_8975,N_8991);
or U9033 (N_9033,N_8898,N_8766);
xor U9034 (N_9034,N_8713,N_8679);
and U9035 (N_9035,N_8954,N_8594);
xor U9036 (N_9036,N_8656,N_8635);
and U9037 (N_9037,N_8908,N_8516);
or U9038 (N_9038,N_8814,N_8671);
xor U9039 (N_9039,N_8685,N_8573);
xor U9040 (N_9040,N_8667,N_8860);
nor U9041 (N_9041,N_8959,N_8742);
and U9042 (N_9042,N_8968,N_8809);
and U9043 (N_9043,N_8879,N_8735);
or U9044 (N_9044,N_8535,N_8834);
or U9045 (N_9045,N_8627,N_8642);
xnor U9046 (N_9046,N_8733,N_8663);
and U9047 (N_9047,N_8509,N_8796);
xnor U9048 (N_9048,N_8616,N_8677);
or U9049 (N_9049,N_8763,N_8613);
nor U9050 (N_9050,N_8765,N_8803);
nor U9051 (N_9051,N_8871,N_8948);
and U9052 (N_9052,N_8660,N_8696);
nor U9053 (N_9053,N_8719,N_8571);
or U9054 (N_9054,N_8738,N_8789);
xnor U9055 (N_9055,N_8630,N_8527);
and U9056 (N_9056,N_8970,N_8985);
nor U9057 (N_9057,N_8723,N_8683);
xnor U9058 (N_9058,N_8929,N_8979);
and U9059 (N_9059,N_8728,N_8749);
nand U9060 (N_9060,N_8881,N_8863);
nor U9061 (N_9061,N_8720,N_8739);
nand U9062 (N_9062,N_8986,N_8578);
nand U9063 (N_9063,N_8632,N_8743);
nor U9064 (N_9064,N_8624,N_8851);
xnor U9065 (N_9065,N_8857,N_8981);
xnor U9066 (N_9066,N_8887,N_8953);
or U9067 (N_9067,N_8774,N_8550);
and U9068 (N_9068,N_8617,N_8607);
and U9069 (N_9069,N_8729,N_8502);
nor U9070 (N_9070,N_8974,N_8826);
nand U9071 (N_9071,N_8700,N_8697);
and U9072 (N_9072,N_8744,N_8933);
nor U9073 (N_9073,N_8745,N_8651);
and U9074 (N_9074,N_8563,N_8517);
and U9075 (N_9075,N_8681,N_8768);
nor U9076 (N_9076,N_8736,N_8615);
and U9077 (N_9077,N_8769,N_8746);
and U9078 (N_9078,N_8945,N_8920);
nor U9079 (N_9079,N_8602,N_8990);
nand U9080 (N_9080,N_8731,N_8557);
and U9081 (N_9081,N_8568,N_8611);
or U9082 (N_9082,N_8849,N_8546);
or U9083 (N_9083,N_8629,N_8649);
xor U9084 (N_9084,N_8987,N_8506);
or U9085 (N_9085,N_8572,N_8841);
xnor U9086 (N_9086,N_8958,N_8805);
xnor U9087 (N_9087,N_8798,N_8547);
nand U9088 (N_9088,N_8598,N_8819);
xor U9089 (N_9089,N_8589,N_8790);
nand U9090 (N_9090,N_8664,N_8873);
or U9091 (N_9091,N_8810,N_8939);
nor U9092 (N_9092,N_8919,N_8967);
nand U9093 (N_9093,N_8715,N_8646);
and U9094 (N_9094,N_8996,N_8839);
or U9095 (N_9095,N_8876,N_8934);
and U9096 (N_9096,N_8812,N_8673);
nand U9097 (N_9097,N_8626,N_8522);
nand U9098 (N_9098,N_8647,N_8525);
xnor U9099 (N_9099,N_8855,N_8682);
or U9100 (N_9100,N_8889,N_8866);
xnor U9101 (N_9101,N_8605,N_8590);
or U9102 (N_9102,N_8890,N_8791);
nand U9103 (N_9103,N_8534,N_8816);
xnor U9104 (N_9104,N_8930,N_8570);
and U9105 (N_9105,N_8882,N_8832);
and U9106 (N_9106,N_8751,N_8505);
or U9107 (N_9107,N_8693,N_8755);
nand U9108 (N_9108,N_8772,N_8807);
and U9109 (N_9109,N_8587,N_8653);
or U9110 (N_9110,N_8904,N_8843);
xor U9111 (N_9111,N_8982,N_8998);
nor U9112 (N_9112,N_8583,N_8753);
nor U9113 (N_9113,N_8619,N_8722);
or U9114 (N_9114,N_8818,N_8614);
or U9115 (N_9115,N_8836,N_8709);
xor U9116 (N_9116,N_8950,N_8581);
nor U9117 (N_9117,N_8555,N_8699);
xor U9118 (N_9118,N_8907,N_8551);
nand U9119 (N_9119,N_8564,N_8781);
xnor U9120 (N_9120,N_8899,N_8971);
nor U9121 (N_9121,N_8560,N_8775);
and U9122 (N_9122,N_8846,N_8892);
xnor U9123 (N_9123,N_8533,N_8542);
nor U9124 (N_9124,N_8888,N_8965);
or U9125 (N_9125,N_8639,N_8747);
and U9126 (N_9126,N_8916,N_8956);
nor U9127 (N_9127,N_8706,N_8530);
and U9128 (N_9128,N_8622,N_8980);
xnor U9129 (N_9129,N_8575,N_8531);
xnor U9130 (N_9130,N_8915,N_8553);
nor U9131 (N_9131,N_8698,N_8737);
nand U9132 (N_9132,N_8532,N_8518);
xor U9133 (N_9133,N_8507,N_8712);
and U9134 (N_9134,N_8877,N_8925);
nand U9135 (N_9135,N_8872,N_8730);
or U9136 (N_9136,N_8884,N_8504);
or U9137 (N_9137,N_8652,N_8794);
nand U9138 (N_9138,N_8966,N_8902);
nor U9139 (N_9139,N_8610,N_8678);
and U9140 (N_9140,N_8927,N_8777);
nand U9141 (N_9141,N_8515,N_8914);
nor U9142 (N_9142,N_8597,N_8895);
xor U9143 (N_9143,N_8520,N_8512);
xor U9144 (N_9144,N_8764,N_8600);
nor U9145 (N_9145,N_8726,N_8878);
nand U9146 (N_9146,N_8549,N_8514);
and U9147 (N_9147,N_8668,N_8821);
or U9148 (N_9148,N_8599,N_8558);
nand U9149 (N_9149,N_8543,N_8859);
nor U9150 (N_9150,N_8711,N_8654);
xnor U9151 (N_9151,N_8701,N_8567);
and U9152 (N_9152,N_8951,N_8574);
or U9153 (N_9153,N_8705,N_8801);
xnor U9154 (N_9154,N_8724,N_8833);
or U9155 (N_9155,N_8633,N_8989);
or U9156 (N_9156,N_8670,N_8988);
nand U9157 (N_9157,N_8999,N_8928);
nand U9158 (N_9158,N_8662,N_8585);
or U9159 (N_9159,N_8862,N_8831);
nor U9160 (N_9160,N_8992,N_8896);
or U9161 (N_9161,N_8936,N_8707);
nand U9162 (N_9162,N_8984,N_8500);
nor U9163 (N_9163,N_8947,N_8941);
nand U9164 (N_9164,N_8802,N_8850);
or U9165 (N_9165,N_8923,N_8911);
nand U9166 (N_9166,N_8692,N_8838);
nand U9167 (N_9167,N_8659,N_8596);
nor U9168 (N_9168,N_8676,N_8526);
xnor U9169 (N_9169,N_8544,N_8924);
or U9170 (N_9170,N_8848,N_8921);
xnor U9171 (N_9171,N_8541,N_8903);
and U9172 (N_9172,N_8606,N_8845);
nor U9173 (N_9173,N_8638,N_8734);
nor U9174 (N_9174,N_8827,N_8894);
nand U9175 (N_9175,N_8680,N_8932);
and U9176 (N_9176,N_8856,N_8612);
or U9177 (N_9177,N_8865,N_8837);
xnor U9178 (N_9178,N_8815,N_8788);
xor U9179 (N_9179,N_8554,N_8565);
nor U9180 (N_9180,N_8909,N_8508);
xnor U9181 (N_9181,N_8949,N_8511);
nor U9182 (N_9182,N_8847,N_8529);
nor U9183 (N_9183,N_8536,N_8748);
or U9184 (N_9184,N_8625,N_8783);
nand U9185 (N_9185,N_8811,N_8708);
or U9186 (N_9186,N_8880,N_8786);
nand U9187 (N_9187,N_8584,N_8691);
and U9188 (N_9188,N_8806,N_8993);
xor U9189 (N_9189,N_8852,N_8944);
nand U9190 (N_9190,N_8840,N_8727);
nor U9191 (N_9191,N_8926,N_8637);
nand U9192 (N_9192,N_8784,N_8716);
nand U9193 (N_9193,N_8641,N_8608);
and U9194 (N_9194,N_8799,N_8897);
nor U9195 (N_9195,N_8797,N_8955);
and U9196 (N_9196,N_8937,N_8813);
and U9197 (N_9197,N_8644,N_8658);
nor U9198 (N_9198,N_8952,N_8957);
or U9199 (N_9199,N_8577,N_8537);
nor U9200 (N_9200,N_8760,N_8758);
and U9201 (N_9201,N_8754,N_8721);
xor U9202 (N_9202,N_8695,N_8931);
and U9203 (N_9203,N_8655,N_8961);
nand U9204 (N_9204,N_8870,N_8922);
and U9205 (N_9205,N_8672,N_8864);
nor U9206 (N_9206,N_8913,N_8761);
or U9207 (N_9207,N_8778,N_8645);
nand U9208 (N_9208,N_8891,N_8628);
or U9209 (N_9209,N_8650,N_8910);
and U9210 (N_9210,N_8674,N_8702);
and U9211 (N_9211,N_8905,N_8556);
and U9212 (N_9212,N_8545,N_8665);
or U9213 (N_9213,N_8643,N_8808);
nor U9214 (N_9214,N_8946,N_8901);
nand U9215 (N_9215,N_8780,N_8559);
nand U9216 (N_9216,N_8976,N_8767);
nor U9217 (N_9217,N_8552,N_8844);
nor U9218 (N_9218,N_8867,N_8773);
nand U9219 (N_9219,N_8770,N_8539);
and U9220 (N_9220,N_8669,N_8623);
nand U9221 (N_9221,N_8912,N_8503);
nor U9222 (N_9222,N_8963,N_8636);
nand U9223 (N_9223,N_8804,N_8704);
or U9224 (N_9224,N_8579,N_8883);
nand U9225 (N_9225,N_8538,N_8824);
or U9226 (N_9226,N_8621,N_8732);
and U9227 (N_9227,N_8757,N_8523);
nand U9228 (N_9228,N_8820,N_8829);
nor U9229 (N_9229,N_8595,N_8687);
nand U9230 (N_9230,N_8657,N_8823);
nand U9231 (N_9231,N_8900,N_8917);
or U9232 (N_9232,N_8825,N_8787);
nor U9233 (N_9233,N_8861,N_8501);
xnor U9234 (N_9234,N_8703,N_8648);
or U9235 (N_9235,N_8521,N_8893);
xor U9236 (N_9236,N_8875,N_8592);
and U9237 (N_9237,N_8792,N_8943);
nor U9238 (N_9238,N_8822,N_8940);
nand U9239 (N_9239,N_8828,N_8689);
nor U9240 (N_9240,N_8562,N_8604);
or U9241 (N_9241,N_8942,N_8609);
and U9242 (N_9242,N_8631,N_8684);
and U9243 (N_9243,N_8817,N_8858);
nand U9244 (N_9244,N_8740,N_8675);
and U9245 (N_9245,N_8938,N_8714);
xor U9246 (N_9246,N_8983,N_8771);
nor U9247 (N_9247,N_8718,N_8528);
xnor U9248 (N_9248,N_8601,N_8566);
and U9249 (N_9249,N_8842,N_8582);
nand U9250 (N_9250,N_8662,N_8538);
nor U9251 (N_9251,N_8835,N_8941);
and U9252 (N_9252,N_8586,N_8673);
nor U9253 (N_9253,N_8509,N_8924);
nand U9254 (N_9254,N_8562,N_8971);
or U9255 (N_9255,N_8796,N_8639);
xnor U9256 (N_9256,N_8550,N_8970);
or U9257 (N_9257,N_8754,N_8543);
xnor U9258 (N_9258,N_8806,N_8715);
and U9259 (N_9259,N_8662,N_8844);
and U9260 (N_9260,N_8617,N_8815);
and U9261 (N_9261,N_8861,N_8892);
or U9262 (N_9262,N_8683,N_8797);
xor U9263 (N_9263,N_8846,N_8682);
xor U9264 (N_9264,N_8976,N_8549);
or U9265 (N_9265,N_8942,N_8755);
and U9266 (N_9266,N_8582,N_8861);
nand U9267 (N_9267,N_8648,N_8627);
xnor U9268 (N_9268,N_8572,N_8743);
or U9269 (N_9269,N_8934,N_8712);
nor U9270 (N_9270,N_8633,N_8530);
xor U9271 (N_9271,N_8885,N_8928);
xnor U9272 (N_9272,N_8939,N_8903);
nand U9273 (N_9273,N_8719,N_8947);
xor U9274 (N_9274,N_8684,N_8757);
xor U9275 (N_9275,N_8536,N_8588);
or U9276 (N_9276,N_8926,N_8707);
and U9277 (N_9277,N_8581,N_8793);
nor U9278 (N_9278,N_8976,N_8751);
nor U9279 (N_9279,N_8764,N_8569);
or U9280 (N_9280,N_8759,N_8727);
and U9281 (N_9281,N_8531,N_8735);
xnor U9282 (N_9282,N_8829,N_8911);
nand U9283 (N_9283,N_8908,N_8581);
or U9284 (N_9284,N_8529,N_8766);
nor U9285 (N_9285,N_8682,N_8876);
nor U9286 (N_9286,N_8660,N_8700);
xnor U9287 (N_9287,N_8956,N_8500);
nand U9288 (N_9288,N_8546,N_8632);
nor U9289 (N_9289,N_8935,N_8817);
nor U9290 (N_9290,N_8804,N_8800);
nand U9291 (N_9291,N_8781,N_8596);
or U9292 (N_9292,N_8931,N_8817);
and U9293 (N_9293,N_8922,N_8743);
or U9294 (N_9294,N_8696,N_8989);
nand U9295 (N_9295,N_8579,N_8662);
nand U9296 (N_9296,N_8741,N_8886);
xnor U9297 (N_9297,N_8598,N_8763);
xnor U9298 (N_9298,N_8512,N_8758);
or U9299 (N_9299,N_8827,N_8851);
xor U9300 (N_9300,N_8574,N_8869);
or U9301 (N_9301,N_8878,N_8635);
nor U9302 (N_9302,N_8901,N_8504);
nor U9303 (N_9303,N_8871,N_8932);
or U9304 (N_9304,N_8601,N_8665);
or U9305 (N_9305,N_8728,N_8784);
or U9306 (N_9306,N_8791,N_8592);
nand U9307 (N_9307,N_8718,N_8844);
nand U9308 (N_9308,N_8928,N_8686);
nor U9309 (N_9309,N_8793,N_8583);
xor U9310 (N_9310,N_8618,N_8993);
nor U9311 (N_9311,N_8889,N_8686);
and U9312 (N_9312,N_8716,N_8813);
nand U9313 (N_9313,N_8961,N_8894);
nor U9314 (N_9314,N_8781,N_8762);
or U9315 (N_9315,N_8617,N_8520);
and U9316 (N_9316,N_8662,N_8970);
xnor U9317 (N_9317,N_8615,N_8692);
xnor U9318 (N_9318,N_8852,N_8593);
or U9319 (N_9319,N_8588,N_8737);
xnor U9320 (N_9320,N_8681,N_8551);
and U9321 (N_9321,N_8742,N_8624);
nor U9322 (N_9322,N_8920,N_8638);
and U9323 (N_9323,N_8776,N_8922);
or U9324 (N_9324,N_8869,N_8529);
or U9325 (N_9325,N_8715,N_8592);
or U9326 (N_9326,N_8709,N_8954);
xnor U9327 (N_9327,N_8609,N_8749);
nand U9328 (N_9328,N_8938,N_8552);
xor U9329 (N_9329,N_8659,N_8838);
nor U9330 (N_9330,N_8814,N_8575);
and U9331 (N_9331,N_8901,N_8909);
nand U9332 (N_9332,N_8877,N_8892);
xor U9333 (N_9333,N_8906,N_8695);
nand U9334 (N_9334,N_8553,N_8928);
and U9335 (N_9335,N_8775,N_8585);
nor U9336 (N_9336,N_8935,N_8977);
and U9337 (N_9337,N_8629,N_8871);
xnor U9338 (N_9338,N_8954,N_8850);
nor U9339 (N_9339,N_8618,N_8524);
nor U9340 (N_9340,N_8829,N_8822);
xnor U9341 (N_9341,N_8830,N_8929);
nor U9342 (N_9342,N_8798,N_8976);
nand U9343 (N_9343,N_8745,N_8835);
or U9344 (N_9344,N_8753,N_8880);
xor U9345 (N_9345,N_8661,N_8511);
nor U9346 (N_9346,N_8928,N_8530);
nor U9347 (N_9347,N_8913,N_8655);
or U9348 (N_9348,N_8740,N_8533);
nand U9349 (N_9349,N_8903,N_8651);
nand U9350 (N_9350,N_8789,N_8784);
nand U9351 (N_9351,N_8988,N_8588);
or U9352 (N_9352,N_8767,N_8974);
nor U9353 (N_9353,N_8962,N_8873);
or U9354 (N_9354,N_8605,N_8642);
or U9355 (N_9355,N_8972,N_8815);
or U9356 (N_9356,N_8792,N_8596);
xnor U9357 (N_9357,N_8934,N_8759);
or U9358 (N_9358,N_8841,N_8776);
nand U9359 (N_9359,N_8508,N_8829);
and U9360 (N_9360,N_8509,N_8794);
xnor U9361 (N_9361,N_8980,N_8666);
nor U9362 (N_9362,N_8788,N_8925);
xnor U9363 (N_9363,N_8982,N_8778);
nand U9364 (N_9364,N_8746,N_8992);
nor U9365 (N_9365,N_8769,N_8506);
and U9366 (N_9366,N_8758,N_8757);
xnor U9367 (N_9367,N_8627,N_8656);
xnor U9368 (N_9368,N_8835,N_8586);
or U9369 (N_9369,N_8838,N_8668);
or U9370 (N_9370,N_8956,N_8865);
xor U9371 (N_9371,N_8937,N_8914);
and U9372 (N_9372,N_8916,N_8819);
or U9373 (N_9373,N_8837,N_8954);
and U9374 (N_9374,N_8721,N_8711);
xor U9375 (N_9375,N_8888,N_8669);
nor U9376 (N_9376,N_8781,N_8740);
nand U9377 (N_9377,N_8852,N_8613);
or U9378 (N_9378,N_8505,N_8523);
or U9379 (N_9379,N_8771,N_8702);
and U9380 (N_9380,N_8741,N_8529);
xor U9381 (N_9381,N_8837,N_8565);
nor U9382 (N_9382,N_8886,N_8986);
or U9383 (N_9383,N_8529,N_8664);
nand U9384 (N_9384,N_8511,N_8662);
nor U9385 (N_9385,N_8930,N_8592);
or U9386 (N_9386,N_8968,N_8625);
nor U9387 (N_9387,N_8734,N_8925);
xnor U9388 (N_9388,N_8925,N_8825);
or U9389 (N_9389,N_8972,N_8720);
and U9390 (N_9390,N_8633,N_8872);
xor U9391 (N_9391,N_8750,N_8722);
and U9392 (N_9392,N_8905,N_8532);
and U9393 (N_9393,N_8693,N_8590);
xor U9394 (N_9394,N_8709,N_8852);
or U9395 (N_9395,N_8914,N_8683);
nor U9396 (N_9396,N_8924,N_8605);
nand U9397 (N_9397,N_8540,N_8815);
nor U9398 (N_9398,N_8536,N_8990);
and U9399 (N_9399,N_8778,N_8959);
and U9400 (N_9400,N_8880,N_8500);
and U9401 (N_9401,N_8847,N_8945);
xor U9402 (N_9402,N_8501,N_8671);
xor U9403 (N_9403,N_8622,N_8617);
nand U9404 (N_9404,N_8755,N_8745);
or U9405 (N_9405,N_8759,N_8589);
or U9406 (N_9406,N_8691,N_8602);
or U9407 (N_9407,N_8944,N_8850);
xor U9408 (N_9408,N_8918,N_8544);
nor U9409 (N_9409,N_8807,N_8820);
and U9410 (N_9410,N_8595,N_8514);
nor U9411 (N_9411,N_8708,N_8685);
nor U9412 (N_9412,N_8821,N_8600);
and U9413 (N_9413,N_8636,N_8864);
nand U9414 (N_9414,N_8584,N_8895);
and U9415 (N_9415,N_8878,N_8703);
and U9416 (N_9416,N_8869,N_8601);
nor U9417 (N_9417,N_8944,N_8743);
or U9418 (N_9418,N_8740,N_8609);
and U9419 (N_9419,N_8665,N_8878);
nor U9420 (N_9420,N_8864,N_8556);
and U9421 (N_9421,N_8696,N_8561);
or U9422 (N_9422,N_8568,N_8950);
xnor U9423 (N_9423,N_8819,N_8633);
and U9424 (N_9424,N_8637,N_8509);
nand U9425 (N_9425,N_8871,N_8819);
nor U9426 (N_9426,N_8975,N_8509);
or U9427 (N_9427,N_8618,N_8677);
xor U9428 (N_9428,N_8785,N_8677);
or U9429 (N_9429,N_8541,N_8584);
or U9430 (N_9430,N_8776,N_8739);
xor U9431 (N_9431,N_8522,N_8523);
and U9432 (N_9432,N_8782,N_8551);
and U9433 (N_9433,N_8957,N_8723);
xor U9434 (N_9434,N_8594,N_8513);
xor U9435 (N_9435,N_8952,N_8706);
and U9436 (N_9436,N_8769,N_8798);
nor U9437 (N_9437,N_8543,N_8548);
nor U9438 (N_9438,N_8592,N_8650);
or U9439 (N_9439,N_8585,N_8607);
nor U9440 (N_9440,N_8792,N_8876);
xor U9441 (N_9441,N_8596,N_8804);
nor U9442 (N_9442,N_8604,N_8693);
and U9443 (N_9443,N_8770,N_8772);
xor U9444 (N_9444,N_8956,N_8569);
or U9445 (N_9445,N_8561,N_8513);
xnor U9446 (N_9446,N_8567,N_8699);
or U9447 (N_9447,N_8962,N_8723);
and U9448 (N_9448,N_8892,N_8810);
or U9449 (N_9449,N_8872,N_8798);
xnor U9450 (N_9450,N_8527,N_8634);
xnor U9451 (N_9451,N_8528,N_8676);
nor U9452 (N_9452,N_8704,N_8839);
and U9453 (N_9453,N_8888,N_8515);
and U9454 (N_9454,N_8509,N_8904);
nand U9455 (N_9455,N_8987,N_8715);
nand U9456 (N_9456,N_8783,N_8643);
xor U9457 (N_9457,N_8644,N_8843);
nor U9458 (N_9458,N_8737,N_8541);
nor U9459 (N_9459,N_8764,N_8895);
nor U9460 (N_9460,N_8510,N_8839);
nor U9461 (N_9461,N_8887,N_8810);
or U9462 (N_9462,N_8591,N_8860);
nor U9463 (N_9463,N_8972,N_8500);
nor U9464 (N_9464,N_8636,N_8999);
nor U9465 (N_9465,N_8546,N_8687);
nor U9466 (N_9466,N_8876,N_8642);
nand U9467 (N_9467,N_8807,N_8984);
nor U9468 (N_9468,N_8911,N_8889);
xnor U9469 (N_9469,N_8976,N_8654);
nand U9470 (N_9470,N_8935,N_8739);
nor U9471 (N_9471,N_8884,N_8900);
or U9472 (N_9472,N_8854,N_8589);
nand U9473 (N_9473,N_8511,N_8938);
and U9474 (N_9474,N_8951,N_8549);
nor U9475 (N_9475,N_8571,N_8784);
nand U9476 (N_9476,N_8735,N_8607);
and U9477 (N_9477,N_8973,N_8612);
xor U9478 (N_9478,N_8531,N_8786);
xor U9479 (N_9479,N_8607,N_8996);
nand U9480 (N_9480,N_8621,N_8729);
or U9481 (N_9481,N_8736,N_8975);
and U9482 (N_9482,N_8550,N_8505);
nor U9483 (N_9483,N_8910,N_8676);
xor U9484 (N_9484,N_8876,N_8848);
xnor U9485 (N_9485,N_8545,N_8750);
and U9486 (N_9486,N_8894,N_8517);
nand U9487 (N_9487,N_8938,N_8581);
or U9488 (N_9488,N_8689,N_8643);
or U9489 (N_9489,N_8761,N_8973);
nand U9490 (N_9490,N_8601,N_8615);
and U9491 (N_9491,N_8949,N_8839);
or U9492 (N_9492,N_8531,N_8961);
nand U9493 (N_9493,N_8939,N_8860);
or U9494 (N_9494,N_8938,N_8879);
and U9495 (N_9495,N_8844,N_8752);
and U9496 (N_9496,N_8515,N_8607);
xor U9497 (N_9497,N_8756,N_8747);
or U9498 (N_9498,N_8819,N_8642);
nand U9499 (N_9499,N_8873,N_8898);
and U9500 (N_9500,N_9173,N_9255);
nand U9501 (N_9501,N_9087,N_9248);
nand U9502 (N_9502,N_9240,N_9368);
nor U9503 (N_9503,N_9011,N_9249);
xor U9504 (N_9504,N_9477,N_9130);
nor U9505 (N_9505,N_9127,N_9456);
xnor U9506 (N_9506,N_9306,N_9180);
xor U9507 (N_9507,N_9126,N_9488);
xor U9508 (N_9508,N_9146,N_9069);
and U9509 (N_9509,N_9238,N_9001);
or U9510 (N_9510,N_9359,N_9431);
or U9511 (N_9511,N_9288,N_9223);
or U9512 (N_9512,N_9334,N_9405);
xor U9513 (N_9513,N_9053,N_9467);
xnor U9514 (N_9514,N_9028,N_9203);
and U9515 (N_9515,N_9260,N_9473);
nor U9516 (N_9516,N_9090,N_9161);
or U9517 (N_9517,N_9188,N_9455);
nand U9518 (N_9518,N_9309,N_9262);
nor U9519 (N_9519,N_9354,N_9474);
and U9520 (N_9520,N_9142,N_9231);
xnor U9521 (N_9521,N_9493,N_9373);
nand U9522 (N_9522,N_9475,N_9264);
and U9523 (N_9523,N_9189,N_9035);
nand U9524 (N_9524,N_9453,N_9417);
nor U9525 (N_9525,N_9367,N_9463);
or U9526 (N_9526,N_9479,N_9027);
or U9527 (N_9527,N_9466,N_9224);
nor U9528 (N_9528,N_9084,N_9128);
nand U9529 (N_9529,N_9049,N_9254);
nand U9530 (N_9530,N_9406,N_9147);
or U9531 (N_9531,N_9149,N_9391);
and U9532 (N_9532,N_9386,N_9287);
and U9533 (N_9533,N_9423,N_9424);
and U9534 (N_9534,N_9039,N_9218);
and U9535 (N_9535,N_9194,N_9086);
nor U9536 (N_9536,N_9274,N_9232);
or U9537 (N_9537,N_9119,N_9332);
and U9538 (N_9538,N_9157,N_9046);
nor U9539 (N_9539,N_9132,N_9165);
and U9540 (N_9540,N_9044,N_9153);
nand U9541 (N_9541,N_9398,N_9206);
nand U9542 (N_9542,N_9158,N_9104);
and U9543 (N_9543,N_9250,N_9190);
nand U9544 (N_9544,N_9122,N_9056);
and U9545 (N_9545,N_9442,N_9022);
nand U9546 (N_9546,N_9394,N_9176);
xor U9547 (N_9547,N_9459,N_9333);
xnor U9548 (N_9548,N_9498,N_9380);
xnor U9549 (N_9549,N_9031,N_9003);
or U9550 (N_9550,N_9198,N_9246);
xnor U9551 (N_9551,N_9362,N_9308);
nand U9552 (N_9552,N_9045,N_9484);
nand U9553 (N_9553,N_9156,N_9166);
and U9554 (N_9554,N_9018,N_9050);
nand U9555 (N_9555,N_9286,N_9026);
or U9556 (N_9556,N_9441,N_9037);
and U9557 (N_9557,N_9416,N_9004);
xnor U9558 (N_9558,N_9000,N_9444);
nor U9559 (N_9559,N_9404,N_9296);
nand U9560 (N_9560,N_9034,N_9192);
nand U9561 (N_9561,N_9272,N_9413);
and U9562 (N_9562,N_9412,N_9201);
xnor U9563 (N_9563,N_9209,N_9105);
or U9564 (N_9564,N_9317,N_9136);
nor U9565 (N_9565,N_9275,N_9181);
nor U9566 (N_9566,N_9042,N_9364);
nor U9567 (N_9567,N_9108,N_9059);
and U9568 (N_9568,N_9419,N_9361);
nor U9569 (N_9569,N_9277,N_9338);
xor U9570 (N_9570,N_9174,N_9072);
nor U9571 (N_9571,N_9107,N_9326);
and U9572 (N_9572,N_9103,N_9392);
and U9573 (N_9573,N_9055,N_9278);
or U9574 (N_9574,N_9239,N_9213);
or U9575 (N_9575,N_9487,N_9483);
xnor U9576 (N_9576,N_9495,N_9196);
and U9577 (N_9577,N_9141,N_9124);
nor U9578 (N_9578,N_9490,N_9030);
nor U9579 (N_9579,N_9060,N_9081);
nor U9580 (N_9580,N_9307,N_9193);
nor U9581 (N_9581,N_9096,N_9305);
nand U9582 (N_9582,N_9251,N_9002);
xor U9583 (N_9583,N_9470,N_9175);
nor U9584 (N_9584,N_9397,N_9208);
and U9585 (N_9585,N_9065,N_9300);
xor U9586 (N_9586,N_9312,N_9331);
and U9587 (N_9587,N_9497,N_9010);
xor U9588 (N_9588,N_9471,N_9320);
and U9589 (N_9589,N_9123,N_9187);
nand U9590 (N_9590,N_9099,N_9408);
nor U9591 (N_9591,N_9183,N_9088);
xnor U9592 (N_9592,N_9178,N_9452);
nor U9593 (N_9593,N_9399,N_9427);
or U9594 (N_9594,N_9291,N_9294);
xnor U9595 (N_9595,N_9205,N_9265);
nor U9596 (N_9596,N_9169,N_9491);
nor U9597 (N_9597,N_9051,N_9472);
xnor U9598 (N_9598,N_9071,N_9390);
and U9599 (N_9599,N_9216,N_9219);
nand U9600 (N_9600,N_9339,N_9019);
and U9601 (N_9601,N_9095,N_9024);
nor U9602 (N_9602,N_9343,N_9379);
xnor U9603 (N_9603,N_9237,N_9435);
nor U9604 (N_9604,N_9225,N_9365);
nand U9605 (N_9605,N_9247,N_9014);
or U9606 (N_9606,N_9481,N_9243);
and U9607 (N_9607,N_9064,N_9043);
and U9608 (N_9608,N_9350,N_9324);
xor U9609 (N_9609,N_9450,N_9073);
xnor U9610 (N_9610,N_9315,N_9113);
or U9611 (N_9611,N_9370,N_9328);
nor U9612 (N_9612,N_9280,N_9252);
xor U9613 (N_9613,N_9438,N_9415);
xnor U9614 (N_9614,N_9335,N_9214);
xor U9615 (N_9615,N_9314,N_9047);
nor U9616 (N_9616,N_9369,N_9494);
xnor U9617 (N_9617,N_9330,N_9321);
and U9618 (N_9618,N_9139,N_9032);
or U9619 (N_9619,N_9179,N_9302);
xnor U9620 (N_9620,N_9215,N_9449);
or U9621 (N_9621,N_9461,N_9485);
xnor U9622 (N_9622,N_9110,N_9098);
and U9623 (N_9623,N_9229,N_9318);
and U9624 (N_9624,N_9411,N_9311);
xor U9625 (N_9625,N_9325,N_9385);
xnor U9626 (N_9626,N_9293,N_9348);
and U9627 (N_9627,N_9184,N_9100);
or U9628 (N_9628,N_9058,N_9245);
nor U9629 (N_9629,N_9410,N_9242);
or U9630 (N_9630,N_9268,N_9144);
nor U9631 (N_9631,N_9101,N_9109);
nor U9632 (N_9632,N_9094,N_9186);
nand U9633 (N_9633,N_9077,N_9222);
and U9634 (N_9634,N_9057,N_9261);
and U9635 (N_9635,N_9115,N_9038);
xor U9636 (N_9636,N_9227,N_9154);
nand U9637 (N_9637,N_9304,N_9396);
nor U9638 (N_9638,N_9148,N_9270);
nand U9639 (N_9639,N_9061,N_9244);
or U9640 (N_9640,N_9393,N_9257);
or U9641 (N_9641,N_9155,N_9355);
nand U9642 (N_9642,N_9151,N_9012);
xnor U9643 (N_9643,N_9292,N_9258);
or U9644 (N_9644,N_9421,N_9478);
nand U9645 (N_9645,N_9135,N_9269);
nor U9646 (N_9646,N_9353,N_9372);
xnor U9647 (N_9647,N_9211,N_9093);
and U9648 (N_9648,N_9160,N_9395);
nor U9649 (N_9649,N_9210,N_9138);
and U9650 (N_9650,N_9460,N_9167);
and U9651 (N_9651,N_9076,N_9233);
and U9652 (N_9652,N_9329,N_9499);
and U9653 (N_9653,N_9143,N_9054);
or U9654 (N_9654,N_9137,N_9120);
or U9655 (N_9655,N_9079,N_9383);
and U9656 (N_9656,N_9357,N_9066);
xor U9657 (N_9657,N_9008,N_9344);
nor U9658 (N_9658,N_9259,N_9133);
nor U9659 (N_9659,N_9041,N_9029);
or U9660 (N_9660,N_9033,N_9017);
and U9661 (N_9661,N_9145,N_9177);
and U9662 (N_9662,N_9407,N_9414);
or U9663 (N_9663,N_9439,N_9428);
and U9664 (N_9664,N_9204,N_9013);
nand U9665 (N_9665,N_9048,N_9068);
or U9666 (N_9666,N_9443,N_9235);
xor U9667 (N_9667,N_9284,N_9371);
or U9668 (N_9668,N_9476,N_9273);
xnor U9669 (N_9669,N_9400,N_9097);
and U9670 (N_9670,N_9106,N_9403);
and U9671 (N_9671,N_9020,N_9276);
and U9672 (N_9672,N_9164,N_9469);
xor U9673 (N_9673,N_9451,N_9360);
nor U9674 (N_9674,N_9062,N_9426);
nor U9675 (N_9675,N_9377,N_9376);
nand U9676 (N_9676,N_9346,N_9327);
or U9677 (N_9677,N_9425,N_9226);
nor U9678 (N_9678,N_9114,N_9290);
xor U9679 (N_9679,N_9436,N_9085);
xnor U9680 (N_9680,N_9468,N_9131);
or U9681 (N_9681,N_9492,N_9295);
nor U9682 (N_9682,N_9234,N_9375);
or U9683 (N_9683,N_9366,N_9125);
nand U9684 (N_9684,N_9263,N_9358);
or U9685 (N_9685,N_9285,N_9191);
xnor U9686 (N_9686,N_9299,N_9241);
and U9687 (N_9687,N_9462,N_9430);
or U9688 (N_9688,N_9134,N_9363);
and U9689 (N_9689,N_9384,N_9454);
nor U9690 (N_9690,N_9089,N_9091);
xor U9691 (N_9691,N_9313,N_9446);
nand U9692 (N_9692,N_9117,N_9422);
xor U9693 (N_9693,N_9070,N_9322);
or U9694 (N_9694,N_9195,N_9447);
and U9695 (N_9695,N_9199,N_9006);
nand U9696 (N_9696,N_9282,N_9389);
or U9697 (N_9697,N_9217,N_9075);
nor U9698 (N_9698,N_9168,N_9323);
nor U9699 (N_9699,N_9401,N_9440);
xor U9700 (N_9700,N_9342,N_9009);
nand U9701 (N_9701,N_9266,N_9007);
and U9702 (N_9702,N_9116,N_9170);
xnor U9703 (N_9703,N_9349,N_9200);
and U9704 (N_9704,N_9310,N_9387);
or U9705 (N_9705,N_9074,N_9297);
xor U9706 (N_9706,N_9303,N_9202);
nand U9707 (N_9707,N_9212,N_9301);
or U9708 (N_9708,N_9256,N_9092);
nor U9709 (N_9709,N_9437,N_9388);
or U9710 (N_9710,N_9221,N_9378);
nand U9711 (N_9711,N_9480,N_9253);
or U9712 (N_9712,N_9382,N_9159);
nor U9713 (N_9713,N_9345,N_9418);
or U9714 (N_9714,N_9220,N_9236);
nor U9715 (N_9715,N_9429,N_9036);
nor U9716 (N_9716,N_9351,N_9207);
and U9717 (N_9717,N_9316,N_9015);
nor U9718 (N_9718,N_9197,N_9352);
nor U9719 (N_9719,N_9172,N_9067);
nor U9720 (N_9720,N_9271,N_9083);
nand U9721 (N_9721,N_9347,N_9021);
xnor U9722 (N_9722,N_9063,N_9140);
or U9723 (N_9723,N_9129,N_9267);
nor U9724 (N_9724,N_9496,N_9080);
nor U9725 (N_9725,N_9171,N_9289);
xor U9726 (N_9726,N_9434,N_9111);
xor U9727 (N_9727,N_9005,N_9341);
nor U9728 (N_9728,N_9445,N_9102);
nand U9729 (N_9729,N_9230,N_9112);
or U9730 (N_9730,N_9409,N_9016);
and U9731 (N_9731,N_9228,N_9448);
and U9732 (N_9732,N_9185,N_9152);
xor U9733 (N_9733,N_9182,N_9118);
nor U9734 (N_9734,N_9340,N_9432);
nand U9735 (N_9735,N_9374,N_9281);
xnor U9736 (N_9736,N_9283,N_9457);
or U9737 (N_9737,N_9025,N_9464);
or U9738 (N_9738,N_9465,N_9433);
xor U9739 (N_9739,N_9458,N_9489);
and U9740 (N_9740,N_9402,N_9336);
nor U9741 (N_9741,N_9319,N_9337);
nand U9742 (N_9742,N_9052,N_9163);
nand U9743 (N_9743,N_9121,N_9040);
and U9744 (N_9744,N_9356,N_9023);
xor U9745 (N_9745,N_9162,N_9381);
or U9746 (N_9746,N_9150,N_9482);
or U9747 (N_9747,N_9420,N_9486);
nor U9748 (N_9748,N_9082,N_9279);
xor U9749 (N_9749,N_9078,N_9298);
nand U9750 (N_9750,N_9380,N_9279);
nand U9751 (N_9751,N_9088,N_9070);
nand U9752 (N_9752,N_9261,N_9324);
nor U9753 (N_9753,N_9008,N_9463);
or U9754 (N_9754,N_9447,N_9186);
nor U9755 (N_9755,N_9349,N_9088);
or U9756 (N_9756,N_9213,N_9106);
xnor U9757 (N_9757,N_9074,N_9368);
xor U9758 (N_9758,N_9041,N_9498);
nor U9759 (N_9759,N_9110,N_9140);
nor U9760 (N_9760,N_9486,N_9032);
or U9761 (N_9761,N_9486,N_9135);
and U9762 (N_9762,N_9042,N_9310);
nand U9763 (N_9763,N_9098,N_9194);
or U9764 (N_9764,N_9068,N_9044);
and U9765 (N_9765,N_9289,N_9368);
and U9766 (N_9766,N_9466,N_9299);
xor U9767 (N_9767,N_9245,N_9381);
xor U9768 (N_9768,N_9427,N_9052);
or U9769 (N_9769,N_9275,N_9089);
xor U9770 (N_9770,N_9465,N_9212);
or U9771 (N_9771,N_9192,N_9444);
or U9772 (N_9772,N_9263,N_9403);
and U9773 (N_9773,N_9000,N_9493);
nor U9774 (N_9774,N_9416,N_9180);
xnor U9775 (N_9775,N_9448,N_9188);
or U9776 (N_9776,N_9311,N_9346);
or U9777 (N_9777,N_9491,N_9320);
nand U9778 (N_9778,N_9435,N_9094);
or U9779 (N_9779,N_9430,N_9232);
nor U9780 (N_9780,N_9105,N_9217);
nor U9781 (N_9781,N_9371,N_9317);
nor U9782 (N_9782,N_9190,N_9125);
nor U9783 (N_9783,N_9183,N_9163);
nor U9784 (N_9784,N_9437,N_9131);
or U9785 (N_9785,N_9167,N_9127);
and U9786 (N_9786,N_9424,N_9358);
and U9787 (N_9787,N_9446,N_9181);
nand U9788 (N_9788,N_9406,N_9389);
xor U9789 (N_9789,N_9250,N_9369);
nand U9790 (N_9790,N_9246,N_9484);
or U9791 (N_9791,N_9067,N_9286);
and U9792 (N_9792,N_9373,N_9269);
xnor U9793 (N_9793,N_9028,N_9366);
nor U9794 (N_9794,N_9355,N_9123);
xnor U9795 (N_9795,N_9283,N_9364);
and U9796 (N_9796,N_9463,N_9024);
xor U9797 (N_9797,N_9105,N_9375);
nand U9798 (N_9798,N_9049,N_9239);
xnor U9799 (N_9799,N_9283,N_9101);
or U9800 (N_9800,N_9404,N_9043);
or U9801 (N_9801,N_9430,N_9258);
nor U9802 (N_9802,N_9325,N_9438);
nor U9803 (N_9803,N_9065,N_9106);
or U9804 (N_9804,N_9435,N_9318);
nand U9805 (N_9805,N_9297,N_9280);
or U9806 (N_9806,N_9475,N_9211);
or U9807 (N_9807,N_9359,N_9265);
or U9808 (N_9808,N_9071,N_9292);
or U9809 (N_9809,N_9155,N_9203);
xor U9810 (N_9810,N_9058,N_9164);
nor U9811 (N_9811,N_9278,N_9166);
or U9812 (N_9812,N_9320,N_9131);
and U9813 (N_9813,N_9494,N_9346);
xnor U9814 (N_9814,N_9323,N_9033);
nand U9815 (N_9815,N_9083,N_9241);
xor U9816 (N_9816,N_9347,N_9389);
nand U9817 (N_9817,N_9487,N_9243);
or U9818 (N_9818,N_9085,N_9180);
nor U9819 (N_9819,N_9235,N_9117);
or U9820 (N_9820,N_9325,N_9424);
and U9821 (N_9821,N_9404,N_9161);
or U9822 (N_9822,N_9365,N_9419);
and U9823 (N_9823,N_9326,N_9388);
or U9824 (N_9824,N_9009,N_9371);
nor U9825 (N_9825,N_9393,N_9326);
nand U9826 (N_9826,N_9435,N_9252);
nand U9827 (N_9827,N_9465,N_9469);
and U9828 (N_9828,N_9473,N_9485);
nand U9829 (N_9829,N_9213,N_9224);
and U9830 (N_9830,N_9151,N_9061);
and U9831 (N_9831,N_9024,N_9223);
nor U9832 (N_9832,N_9136,N_9013);
nor U9833 (N_9833,N_9070,N_9126);
nand U9834 (N_9834,N_9072,N_9207);
or U9835 (N_9835,N_9327,N_9093);
nor U9836 (N_9836,N_9368,N_9193);
xnor U9837 (N_9837,N_9037,N_9231);
nand U9838 (N_9838,N_9418,N_9237);
xor U9839 (N_9839,N_9161,N_9066);
and U9840 (N_9840,N_9015,N_9051);
and U9841 (N_9841,N_9293,N_9443);
xor U9842 (N_9842,N_9350,N_9475);
and U9843 (N_9843,N_9099,N_9180);
nand U9844 (N_9844,N_9431,N_9314);
nor U9845 (N_9845,N_9064,N_9406);
xor U9846 (N_9846,N_9445,N_9205);
or U9847 (N_9847,N_9407,N_9299);
xnor U9848 (N_9848,N_9405,N_9303);
nor U9849 (N_9849,N_9181,N_9067);
and U9850 (N_9850,N_9426,N_9034);
nor U9851 (N_9851,N_9322,N_9489);
xor U9852 (N_9852,N_9435,N_9086);
or U9853 (N_9853,N_9058,N_9289);
xnor U9854 (N_9854,N_9003,N_9226);
xor U9855 (N_9855,N_9324,N_9325);
nor U9856 (N_9856,N_9476,N_9057);
and U9857 (N_9857,N_9397,N_9049);
nand U9858 (N_9858,N_9355,N_9235);
and U9859 (N_9859,N_9210,N_9330);
xor U9860 (N_9860,N_9040,N_9182);
nor U9861 (N_9861,N_9329,N_9347);
or U9862 (N_9862,N_9068,N_9047);
nand U9863 (N_9863,N_9478,N_9126);
or U9864 (N_9864,N_9358,N_9088);
xnor U9865 (N_9865,N_9141,N_9148);
xor U9866 (N_9866,N_9374,N_9027);
and U9867 (N_9867,N_9112,N_9117);
xor U9868 (N_9868,N_9040,N_9097);
or U9869 (N_9869,N_9480,N_9008);
and U9870 (N_9870,N_9294,N_9338);
xor U9871 (N_9871,N_9258,N_9324);
xor U9872 (N_9872,N_9402,N_9487);
nand U9873 (N_9873,N_9088,N_9324);
nor U9874 (N_9874,N_9025,N_9290);
nor U9875 (N_9875,N_9478,N_9330);
and U9876 (N_9876,N_9487,N_9339);
nor U9877 (N_9877,N_9029,N_9406);
xnor U9878 (N_9878,N_9277,N_9296);
and U9879 (N_9879,N_9072,N_9471);
or U9880 (N_9880,N_9313,N_9411);
or U9881 (N_9881,N_9452,N_9104);
nor U9882 (N_9882,N_9431,N_9102);
and U9883 (N_9883,N_9001,N_9412);
nor U9884 (N_9884,N_9064,N_9051);
xor U9885 (N_9885,N_9218,N_9352);
xnor U9886 (N_9886,N_9445,N_9451);
and U9887 (N_9887,N_9030,N_9225);
xor U9888 (N_9888,N_9403,N_9230);
and U9889 (N_9889,N_9342,N_9424);
and U9890 (N_9890,N_9164,N_9088);
xnor U9891 (N_9891,N_9426,N_9228);
nand U9892 (N_9892,N_9190,N_9412);
nand U9893 (N_9893,N_9383,N_9128);
xor U9894 (N_9894,N_9233,N_9449);
nand U9895 (N_9895,N_9356,N_9141);
nor U9896 (N_9896,N_9244,N_9141);
nor U9897 (N_9897,N_9232,N_9499);
nand U9898 (N_9898,N_9416,N_9318);
and U9899 (N_9899,N_9076,N_9199);
and U9900 (N_9900,N_9376,N_9000);
nor U9901 (N_9901,N_9371,N_9421);
xnor U9902 (N_9902,N_9180,N_9458);
nand U9903 (N_9903,N_9198,N_9387);
nor U9904 (N_9904,N_9185,N_9274);
xnor U9905 (N_9905,N_9086,N_9215);
nand U9906 (N_9906,N_9208,N_9374);
or U9907 (N_9907,N_9272,N_9274);
or U9908 (N_9908,N_9061,N_9463);
nand U9909 (N_9909,N_9351,N_9236);
nor U9910 (N_9910,N_9098,N_9048);
nand U9911 (N_9911,N_9102,N_9108);
xor U9912 (N_9912,N_9231,N_9005);
nor U9913 (N_9913,N_9024,N_9292);
nand U9914 (N_9914,N_9220,N_9020);
xnor U9915 (N_9915,N_9433,N_9487);
nand U9916 (N_9916,N_9042,N_9456);
nand U9917 (N_9917,N_9283,N_9001);
xor U9918 (N_9918,N_9297,N_9285);
or U9919 (N_9919,N_9242,N_9160);
and U9920 (N_9920,N_9086,N_9436);
xor U9921 (N_9921,N_9116,N_9478);
and U9922 (N_9922,N_9033,N_9345);
and U9923 (N_9923,N_9437,N_9147);
xnor U9924 (N_9924,N_9001,N_9305);
and U9925 (N_9925,N_9442,N_9151);
and U9926 (N_9926,N_9268,N_9267);
xor U9927 (N_9927,N_9144,N_9215);
and U9928 (N_9928,N_9440,N_9132);
nand U9929 (N_9929,N_9090,N_9208);
xor U9930 (N_9930,N_9182,N_9094);
nor U9931 (N_9931,N_9296,N_9386);
and U9932 (N_9932,N_9159,N_9025);
xor U9933 (N_9933,N_9027,N_9272);
nand U9934 (N_9934,N_9265,N_9104);
nor U9935 (N_9935,N_9204,N_9100);
nand U9936 (N_9936,N_9012,N_9258);
nor U9937 (N_9937,N_9205,N_9199);
nor U9938 (N_9938,N_9315,N_9091);
xor U9939 (N_9939,N_9011,N_9376);
nand U9940 (N_9940,N_9417,N_9390);
and U9941 (N_9941,N_9090,N_9086);
or U9942 (N_9942,N_9175,N_9400);
and U9943 (N_9943,N_9122,N_9274);
xnor U9944 (N_9944,N_9241,N_9422);
and U9945 (N_9945,N_9297,N_9365);
nor U9946 (N_9946,N_9324,N_9275);
nor U9947 (N_9947,N_9123,N_9362);
xor U9948 (N_9948,N_9223,N_9405);
and U9949 (N_9949,N_9369,N_9216);
xnor U9950 (N_9950,N_9421,N_9292);
xnor U9951 (N_9951,N_9320,N_9202);
or U9952 (N_9952,N_9129,N_9309);
nor U9953 (N_9953,N_9401,N_9381);
nand U9954 (N_9954,N_9370,N_9402);
or U9955 (N_9955,N_9224,N_9226);
and U9956 (N_9956,N_9359,N_9262);
nand U9957 (N_9957,N_9437,N_9356);
or U9958 (N_9958,N_9146,N_9262);
nand U9959 (N_9959,N_9495,N_9380);
or U9960 (N_9960,N_9031,N_9016);
and U9961 (N_9961,N_9178,N_9416);
and U9962 (N_9962,N_9212,N_9252);
or U9963 (N_9963,N_9359,N_9170);
nor U9964 (N_9964,N_9245,N_9423);
nor U9965 (N_9965,N_9485,N_9130);
or U9966 (N_9966,N_9464,N_9265);
nand U9967 (N_9967,N_9465,N_9172);
xor U9968 (N_9968,N_9066,N_9148);
nand U9969 (N_9969,N_9492,N_9440);
and U9970 (N_9970,N_9224,N_9059);
and U9971 (N_9971,N_9106,N_9366);
nand U9972 (N_9972,N_9201,N_9004);
or U9973 (N_9973,N_9257,N_9146);
nand U9974 (N_9974,N_9487,N_9313);
nor U9975 (N_9975,N_9197,N_9319);
and U9976 (N_9976,N_9153,N_9158);
and U9977 (N_9977,N_9085,N_9162);
and U9978 (N_9978,N_9068,N_9160);
nand U9979 (N_9979,N_9481,N_9283);
or U9980 (N_9980,N_9011,N_9243);
and U9981 (N_9981,N_9248,N_9416);
or U9982 (N_9982,N_9046,N_9441);
nor U9983 (N_9983,N_9316,N_9309);
nand U9984 (N_9984,N_9384,N_9109);
nor U9985 (N_9985,N_9309,N_9290);
nand U9986 (N_9986,N_9461,N_9264);
and U9987 (N_9987,N_9248,N_9094);
and U9988 (N_9988,N_9285,N_9273);
nor U9989 (N_9989,N_9371,N_9017);
or U9990 (N_9990,N_9426,N_9359);
nor U9991 (N_9991,N_9270,N_9473);
nand U9992 (N_9992,N_9299,N_9221);
nor U9993 (N_9993,N_9269,N_9054);
nand U9994 (N_9994,N_9153,N_9213);
and U9995 (N_9995,N_9462,N_9412);
or U9996 (N_9996,N_9131,N_9008);
nand U9997 (N_9997,N_9137,N_9179);
or U9998 (N_9998,N_9441,N_9394);
nor U9999 (N_9999,N_9227,N_9043);
nand U10000 (N_10000,N_9711,N_9738);
xor U10001 (N_10001,N_9895,N_9724);
nand U10002 (N_10002,N_9777,N_9651);
nand U10003 (N_10003,N_9971,N_9575);
or U10004 (N_10004,N_9812,N_9698);
and U10005 (N_10005,N_9511,N_9980);
and U10006 (N_10006,N_9784,N_9705);
or U10007 (N_10007,N_9521,N_9569);
nand U10008 (N_10008,N_9645,N_9693);
or U10009 (N_10009,N_9778,N_9633);
nor U10010 (N_10010,N_9675,N_9737);
nand U10011 (N_10011,N_9930,N_9624);
nand U10012 (N_10012,N_9549,N_9665);
nand U10013 (N_10013,N_9764,N_9507);
or U10014 (N_10014,N_9600,N_9831);
xnor U10015 (N_10015,N_9866,N_9736);
or U10016 (N_10016,N_9938,N_9809);
or U10017 (N_10017,N_9918,N_9654);
or U10018 (N_10018,N_9849,N_9677);
nor U10019 (N_10019,N_9584,N_9560);
xnor U10020 (N_10020,N_9854,N_9772);
and U10021 (N_10021,N_9515,N_9689);
xor U10022 (N_10022,N_9529,N_9676);
nand U10023 (N_10023,N_9770,N_9609);
nor U10024 (N_10024,N_9695,N_9702);
nor U10025 (N_10025,N_9935,N_9659);
nand U10026 (N_10026,N_9712,N_9597);
or U10027 (N_10027,N_9986,N_9691);
or U10028 (N_10028,N_9740,N_9969);
xnor U10029 (N_10029,N_9857,N_9890);
nor U10030 (N_10030,N_9541,N_9502);
and U10031 (N_10031,N_9884,N_9836);
xnor U10032 (N_10032,N_9891,N_9623);
and U10033 (N_10033,N_9576,N_9927);
nor U10034 (N_10034,N_9943,N_9808);
and U10035 (N_10035,N_9604,N_9946);
nand U10036 (N_10036,N_9798,N_9819);
nor U10037 (N_10037,N_9843,N_9664);
nand U10038 (N_10038,N_9928,N_9699);
or U10039 (N_10039,N_9629,N_9828);
nand U10040 (N_10040,N_9883,N_9984);
and U10041 (N_10041,N_9720,N_9760);
or U10042 (N_10042,N_9769,N_9936);
nand U10043 (N_10043,N_9917,N_9746);
xor U10044 (N_10044,N_9981,N_9972);
or U10045 (N_10045,N_9611,N_9732);
nand U10046 (N_10046,N_9814,N_9783);
or U10047 (N_10047,N_9678,N_9723);
and U10048 (N_10048,N_9868,N_9513);
nor U10049 (N_10049,N_9733,N_9922);
nand U10050 (N_10050,N_9573,N_9617);
xor U10051 (N_10051,N_9768,N_9944);
and U10052 (N_10052,N_9717,N_9673);
or U10053 (N_10053,N_9873,N_9579);
xor U10054 (N_10054,N_9683,N_9729);
or U10055 (N_10055,N_9806,N_9697);
nor U10056 (N_10056,N_9979,N_9547);
nand U10057 (N_10057,N_9722,N_9779);
nor U10058 (N_10058,N_9878,N_9970);
nor U10059 (N_10059,N_9796,N_9949);
or U10060 (N_10060,N_9512,N_9679);
and U10061 (N_10061,N_9751,N_9688);
nand U10062 (N_10062,N_9838,N_9725);
nand U10063 (N_10063,N_9993,N_9948);
nand U10064 (N_10064,N_9505,N_9911);
xor U10065 (N_10065,N_9718,N_9593);
nand U10066 (N_10066,N_9940,N_9977);
xor U10067 (N_10067,N_9745,N_9627);
nand U10068 (N_10068,N_9754,N_9882);
xnor U10069 (N_10069,N_9839,N_9856);
and U10070 (N_10070,N_9792,N_9719);
nor U10071 (N_10071,N_9650,N_9947);
xnor U10072 (N_10072,N_9646,N_9802);
and U10073 (N_10073,N_9821,N_9861);
nor U10074 (N_10074,N_9880,N_9558);
xnor U10075 (N_10075,N_9537,N_9991);
nand U10076 (N_10076,N_9603,N_9731);
and U10077 (N_10077,N_9909,N_9807);
or U10078 (N_10078,N_9684,N_9516);
and U10079 (N_10079,N_9585,N_9789);
and U10080 (N_10080,N_9741,N_9658);
nor U10081 (N_10081,N_9615,N_9847);
and U10082 (N_10082,N_9990,N_9620);
nor U10083 (N_10083,N_9628,N_9811);
nand U10084 (N_10084,N_9956,N_9566);
xor U10085 (N_10085,N_9714,N_9780);
xor U10086 (N_10086,N_9610,N_9879);
xnor U10087 (N_10087,N_9613,N_9776);
nor U10088 (N_10088,N_9567,N_9716);
nand U10089 (N_10089,N_9832,N_9586);
nor U10090 (N_10090,N_9942,N_9692);
or U10091 (N_10091,N_9510,N_9619);
or U10092 (N_10092,N_9893,N_9605);
nand U10093 (N_10093,N_9929,N_9790);
nand U10094 (N_10094,N_9708,N_9581);
and U10095 (N_10095,N_9904,N_9632);
nand U10096 (N_10096,N_9548,N_9841);
xnor U10097 (N_10097,N_9687,N_9791);
xnor U10098 (N_10098,N_9815,N_9752);
nor U10099 (N_10099,N_9960,N_9899);
xnor U10100 (N_10100,N_9803,N_9703);
nor U10101 (N_10101,N_9570,N_9663);
and U10102 (N_10102,N_9713,N_9910);
and U10103 (N_10103,N_9855,N_9742);
and U10104 (N_10104,N_9998,N_9587);
nand U10105 (N_10105,N_9774,N_9588);
xor U10106 (N_10106,N_9864,N_9589);
or U10107 (N_10107,N_9959,N_9571);
and U10108 (N_10108,N_9996,N_9735);
nor U10109 (N_10109,N_9862,N_9859);
nand U10110 (N_10110,N_9788,N_9592);
or U10111 (N_10111,N_9534,N_9535);
nand U10112 (N_10112,N_9700,N_9544);
and U10113 (N_10113,N_9906,N_9925);
nor U10114 (N_10114,N_9647,N_9978);
nor U10115 (N_10115,N_9590,N_9823);
xnor U10116 (N_10116,N_9564,N_9975);
or U10117 (N_10117,N_9795,N_9835);
nand U10118 (N_10118,N_9853,N_9932);
and U10119 (N_10119,N_9924,N_9867);
nor U10120 (N_10120,N_9536,N_9897);
nand U10121 (N_10121,N_9989,N_9995);
nor U10122 (N_10122,N_9905,N_9870);
xnor U10123 (N_10123,N_9860,N_9591);
nand U10124 (N_10124,N_9945,N_9518);
nand U10125 (N_10125,N_9892,N_9520);
xnor U10126 (N_10126,N_9546,N_9608);
xor U10127 (N_10127,N_9953,N_9829);
and U10128 (N_10128,N_9539,N_9793);
nand U10129 (N_10129,N_9912,N_9509);
nand U10130 (N_10130,N_9639,N_9863);
xnor U10131 (N_10131,N_9921,N_9888);
and U10132 (N_10132,N_9726,N_9545);
nor U10133 (N_10133,N_9973,N_9640);
nand U10134 (N_10134,N_9550,N_9824);
or U10135 (N_10135,N_9680,N_9661);
or U10136 (N_10136,N_9626,N_9577);
xor U10137 (N_10137,N_9985,N_9682);
nand U10138 (N_10138,N_9822,N_9508);
nand U10139 (N_10139,N_9937,N_9637);
and U10140 (N_10140,N_9707,N_9710);
nand U10141 (N_10141,N_9997,N_9757);
or U10142 (N_10142,N_9950,N_9999);
xnor U10143 (N_10143,N_9988,N_9915);
or U10144 (N_10144,N_9887,N_9668);
and U10145 (N_10145,N_9920,N_9551);
nor U10146 (N_10146,N_9580,N_9900);
nor U10147 (N_10147,N_9903,N_9523);
or U10148 (N_10148,N_9876,N_9543);
xor U10149 (N_10149,N_9744,N_9885);
nand U10150 (N_10150,N_9503,N_9635);
nand U10151 (N_10151,N_9607,N_9506);
xnor U10152 (N_10152,N_9952,N_9643);
nor U10153 (N_10153,N_9706,N_9813);
and U10154 (N_10154,N_9553,N_9625);
nor U10155 (N_10155,N_9933,N_9612);
nor U10156 (N_10156,N_9907,N_9554);
nand U10157 (N_10157,N_9845,N_9636);
nand U10158 (N_10158,N_9763,N_9765);
nor U10159 (N_10159,N_9671,N_9622);
xnor U10160 (N_10160,N_9538,N_9753);
or U10161 (N_10161,N_9804,N_9800);
or U10162 (N_10162,N_9517,N_9834);
and U10163 (N_10163,N_9851,N_9652);
nor U10164 (N_10164,N_9786,N_9797);
nand U10165 (N_10165,N_9559,N_9552);
and U10166 (N_10166,N_9734,N_9721);
xor U10167 (N_10167,N_9583,N_9818);
and U10168 (N_10168,N_9974,N_9820);
nand U10169 (N_10169,N_9739,N_9670);
nor U10170 (N_10170,N_9524,N_9846);
or U10171 (N_10171,N_9923,N_9525);
xor U10172 (N_10172,N_9532,N_9842);
and U10173 (N_10173,N_9644,N_9825);
nor U10174 (N_10174,N_9799,N_9965);
xnor U10175 (N_10175,N_9748,N_9982);
and U10176 (N_10176,N_9653,N_9572);
nand U10177 (N_10177,N_9848,N_9992);
nor U10178 (N_10178,N_9962,N_9660);
and U10179 (N_10179,N_9672,N_9730);
xnor U10180 (N_10180,N_9694,N_9830);
xnor U10181 (N_10181,N_9727,N_9898);
xor U10182 (N_10182,N_9630,N_9913);
or U10183 (N_10183,N_9598,N_9785);
and U10184 (N_10184,N_9522,N_9666);
xor U10185 (N_10185,N_9568,N_9787);
nand U10186 (N_10186,N_9667,N_9877);
xnor U10187 (N_10187,N_9649,N_9773);
nor U10188 (N_10188,N_9526,N_9941);
nor U10189 (N_10189,N_9542,N_9685);
nand U10190 (N_10190,N_9728,N_9759);
xor U10191 (N_10191,N_9750,N_9563);
and U10192 (N_10192,N_9871,N_9634);
nor U10193 (N_10193,N_9919,N_9901);
nand U10194 (N_10194,N_9908,N_9963);
xor U10195 (N_10195,N_9987,N_9614);
or U10196 (N_10196,N_9852,N_9826);
and U10197 (N_10197,N_9638,N_9968);
nor U10198 (N_10198,N_9827,N_9964);
xnor U10199 (N_10199,N_9669,N_9967);
or U10200 (N_10200,N_9709,N_9858);
nand U10201 (N_10201,N_9565,N_9954);
nand U10202 (N_10202,N_9994,N_9865);
or U10203 (N_10203,N_9531,N_9926);
and U10204 (N_10204,N_9674,N_9844);
xnor U10205 (N_10205,N_9875,N_9556);
or U10206 (N_10206,N_9662,N_9951);
or U10207 (N_10207,N_9958,N_9771);
nor U10208 (N_10208,N_9775,N_9961);
nand U10209 (N_10209,N_9618,N_9805);
nor U10210 (N_10210,N_9602,N_9504);
or U10211 (N_10211,N_9648,N_9794);
and U10212 (N_10212,N_9533,N_9761);
and U10213 (N_10213,N_9896,N_9561);
and U10214 (N_10214,N_9519,N_9756);
or U10215 (N_10215,N_9766,N_9833);
nor U10216 (N_10216,N_9616,N_9976);
nor U10217 (N_10217,N_9701,N_9931);
and U10218 (N_10218,N_9743,N_9957);
and U10219 (N_10219,N_9655,N_9595);
or U10220 (N_10220,N_9801,N_9501);
xnor U10221 (N_10221,N_9850,N_9934);
and U10222 (N_10222,N_9816,N_9886);
and U10223 (N_10223,N_9690,N_9983);
xor U10224 (N_10224,N_9555,N_9500);
xnor U10225 (N_10225,N_9747,N_9657);
nor U10226 (N_10226,N_9704,N_9869);
or U10227 (N_10227,N_9762,N_9902);
nor U10228 (N_10228,N_9749,N_9540);
nor U10229 (N_10229,N_9557,N_9817);
xnor U10230 (N_10230,N_9642,N_9955);
xnor U10231 (N_10231,N_9767,N_9596);
nor U10232 (N_10232,N_9574,N_9599);
or U10233 (N_10233,N_9594,N_9889);
xor U10234 (N_10234,N_9916,N_9562);
xor U10235 (N_10235,N_9914,N_9696);
xnor U10236 (N_10236,N_9601,N_9641);
and U10237 (N_10237,N_9656,N_9755);
and U10238 (N_10238,N_9606,N_9514);
xor U10239 (N_10239,N_9681,N_9527);
xor U10240 (N_10240,N_9840,N_9578);
nor U10241 (N_10241,N_9621,N_9530);
nand U10242 (N_10242,N_9758,N_9810);
nor U10243 (N_10243,N_9686,N_9837);
xor U10244 (N_10244,N_9631,N_9528);
nand U10245 (N_10245,N_9939,N_9874);
nand U10246 (N_10246,N_9582,N_9782);
and U10247 (N_10247,N_9715,N_9966);
nor U10248 (N_10248,N_9872,N_9781);
nand U10249 (N_10249,N_9894,N_9881);
or U10250 (N_10250,N_9591,N_9545);
nand U10251 (N_10251,N_9641,N_9649);
nand U10252 (N_10252,N_9911,N_9634);
xnor U10253 (N_10253,N_9543,N_9943);
xor U10254 (N_10254,N_9608,N_9533);
or U10255 (N_10255,N_9569,N_9514);
and U10256 (N_10256,N_9649,N_9875);
or U10257 (N_10257,N_9737,N_9702);
nor U10258 (N_10258,N_9690,N_9731);
and U10259 (N_10259,N_9838,N_9504);
or U10260 (N_10260,N_9502,N_9832);
and U10261 (N_10261,N_9621,N_9550);
or U10262 (N_10262,N_9865,N_9898);
and U10263 (N_10263,N_9520,N_9628);
or U10264 (N_10264,N_9947,N_9866);
or U10265 (N_10265,N_9828,N_9766);
or U10266 (N_10266,N_9971,N_9672);
xor U10267 (N_10267,N_9610,N_9529);
xor U10268 (N_10268,N_9701,N_9852);
nand U10269 (N_10269,N_9612,N_9869);
nor U10270 (N_10270,N_9644,N_9831);
nor U10271 (N_10271,N_9783,N_9995);
xnor U10272 (N_10272,N_9699,N_9594);
nand U10273 (N_10273,N_9655,N_9667);
nor U10274 (N_10274,N_9513,N_9957);
nor U10275 (N_10275,N_9787,N_9871);
nand U10276 (N_10276,N_9619,N_9690);
xnor U10277 (N_10277,N_9695,N_9512);
nor U10278 (N_10278,N_9922,N_9841);
nor U10279 (N_10279,N_9807,N_9983);
nand U10280 (N_10280,N_9952,N_9603);
xnor U10281 (N_10281,N_9855,N_9656);
nand U10282 (N_10282,N_9575,N_9675);
xor U10283 (N_10283,N_9567,N_9977);
xnor U10284 (N_10284,N_9942,N_9671);
xor U10285 (N_10285,N_9776,N_9535);
nand U10286 (N_10286,N_9718,N_9754);
xor U10287 (N_10287,N_9872,N_9768);
xor U10288 (N_10288,N_9715,N_9924);
and U10289 (N_10289,N_9817,N_9561);
nand U10290 (N_10290,N_9683,N_9530);
and U10291 (N_10291,N_9908,N_9924);
xor U10292 (N_10292,N_9508,N_9781);
or U10293 (N_10293,N_9634,N_9961);
or U10294 (N_10294,N_9609,N_9679);
nor U10295 (N_10295,N_9547,N_9504);
and U10296 (N_10296,N_9563,N_9624);
xnor U10297 (N_10297,N_9655,N_9837);
nor U10298 (N_10298,N_9983,N_9905);
and U10299 (N_10299,N_9861,N_9915);
and U10300 (N_10300,N_9640,N_9586);
nand U10301 (N_10301,N_9622,N_9896);
xnor U10302 (N_10302,N_9790,N_9607);
nand U10303 (N_10303,N_9535,N_9661);
and U10304 (N_10304,N_9793,N_9581);
and U10305 (N_10305,N_9501,N_9530);
nand U10306 (N_10306,N_9688,N_9951);
nand U10307 (N_10307,N_9827,N_9992);
nand U10308 (N_10308,N_9533,N_9963);
and U10309 (N_10309,N_9607,N_9852);
nand U10310 (N_10310,N_9854,N_9876);
and U10311 (N_10311,N_9933,N_9884);
or U10312 (N_10312,N_9802,N_9851);
and U10313 (N_10313,N_9837,N_9563);
and U10314 (N_10314,N_9893,N_9714);
or U10315 (N_10315,N_9868,N_9596);
or U10316 (N_10316,N_9655,N_9600);
and U10317 (N_10317,N_9905,N_9590);
nor U10318 (N_10318,N_9670,N_9881);
xor U10319 (N_10319,N_9840,N_9630);
nor U10320 (N_10320,N_9850,N_9826);
or U10321 (N_10321,N_9777,N_9614);
xnor U10322 (N_10322,N_9922,N_9636);
and U10323 (N_10323,N_9561,N_9946);
nor U10324 (N_10324,N_9635,N_9705);
and U10325 (N_10325,N_9973,N_9751);
nand U10326 (N_10326,N_9665,N_9674);
xnor U10327 (N_10327,N_9607,N_9689);
and U10328 (N_10328,N_9716,N_9846);
or U10329 (N_10329,N_9743,N_9730);
nor U10330 (N_10330,N_9509,N_9659);
nand U10331 (N_10331,N_9755,N_9575);
and U10332 (N_10332,N_9842,N_9567);
nand U10333 (N_10333,N_9618,N_9919);
xnor U10334 (N_10334,N_9538,N_9936);
xor U10335 (N_10335,N_9598,N_9553);
or U10336 (N_10336,N_9985,N_9922);
and U10337 (N_10337,N_9639,N_9927);
nand U10338 (N_10338,N_9977,N_9621);
xor U10339 (N_10339,N_9901,N_9872);
nor U10340 (N_10340,N_9828,N_9543);
nor U10341 (N_10341,N_9908,N_9812);
nand U10342 (N_10342,N_9621,N_9672);
nor U10343 (N_10343,N_9640,N_9608);
xor U10344 (N_10344,N_9933,N_9892);
nand U10345 (N_10345,N_9581,N_9814);
nor U10346 (N_10346,N_9624,N_9691);
or U10347 (N_10347,N_9517,N_9842);
or U10348 (N_10348,N_9569,N_9860);
nor U10349 (N_10349,N_9503,N_9962);
and U10350 (N_10350,N_9799,N_9608);
nand U10351 (N_10351,N_9875,N_9779);
nor U10352 (N_10352,N_9800,N_9823);
xnor U10353 (N_10353,N_9894,N_9689);
nor U10354 (N_10354,N_9581,N_9537);
xnor U10355 (N_10355,N_9860,N_9791);
and U10356 (N_10356,N_9677,N_9814);
nor U10357 (N_10357,N_9523,N_9645);
nand U10358 (N_10358,N_9961,N_9750);
nand U10359 (N_10359,N_9532,N_9907);
nand U10360 (N_10360,N_9994,N_9583);
xor U10361 (N_10361,N_9573,N_9748);
and U10362 (N_10362,N_9589,N_9655);
and U10363 (N_10363,N_9992,N_9808);
and U10364 (N_10364,N_9942,N_9614);
or U10365 (N_10365,N_9555,N_9668);
nor U10366 (N_10366,N_9816,N_9716);
nor U10367 (N_10367,N_9990,N_9814);
xor U10368 (N_10368,N_9623,N_9860);
xnor U10369 (N_10369,N_9788,N_9521);
or U10370 (N_10370,N_9842,N_9773);
xnor U10371 (N_10371,N_9970,N_9872);
and U10372 (N_10372,N_9877,N_9767);
nor U10373 (N_10373,N_9711,N_9553);
and U10374 (N_10374,N_9861,N_9590);
or U10375 (N_10375,N_9675,N_9994);
xor U10376 (N_10376,N_9926,N_9672);
or U10377 (N_10377,N_9695,N_9699);
or U10378 (N_10378,N_9593,N_9709);
or U10379 (N_10379,N_9946,N_9755);
or U10380 (N_10380,N_9897,N_9954);
or U10381 (N_10381,N_9798,N_9835);
nand U10382 (N_10382,N_9822,N_9519);
and U10383 (N_10383,N_9734,N_9547);
nor U10384 (N_10384,N_9527,N_9671);
nor U10385 (N_10385,N_9572,N_9669);
or U10386 (N_10386,N_9652,N_9750);
nand U10387 (N_10387,N_9974,N_9781);
xor U10388 (N_10388,N_9798,N_9528);
and U10389 (N_10389,N_9964,N_9891);
nor U10390 (N_10390,N_9629,N_9963);
nand U10391 (N_10391,N_9643,N_9565);
nand U10392 (N_10392,N_9957,N_9673);
nor U10393 (N_10393,N_9699,N_9994);
xnor U10394 (N_10394,N_9860,N_9919);
and U10395 (N_10395,N_9931,N_9551);
nand U10396 (N_10396,N_9822,N_9668);
nand U10397 (N_10397,N_9977,N_9561);
nand U10398 (N_10398,N_9777,N_9853);
xor U10399 (N_10399,N_9667,N_9848);
or U10400 (N_10400,N_9928,N_9870);
nor U10401 (N_10401,N_9861,N_9785);
or U10402 (N_10402,N_9983,N_9748);
and U10403 (N_10403,N_9629,N_9925);
nor U10404 (N_10404,N_9588,N_9612);
and U10405 (N_10405,N_9954,N_9725);
or U10406 (N_10406,N_9608,N_9512);
or U10407 (N_10407,N_9652,N_9888);
nor U10408 (N_10408,N_9662,N_9585);
xor U10409 (N_10409,N_9693,N_9772);
or U10410 (N_10410,N_9672,N_9530);
nand U10411 (N_10411,N_9517,N_9933);
nor U10412 (N_10412,N_9534,N_9520);
nand U10413 (N_10413,N_9527,N_9856);
nor U10414 (N_10414,N_9913,N_9932);
and U10415 (N_10415,N_9915,N_9609);
and U10416 (N_10416,N_9615,N_9917);
xor U10417 (N_10417,N_9570,N_9535);
nor U10418 (N_10418,N_9881,N_9744);
nand U10419 (N_10419,N_9893,N_9797);
or U10420 (N_10420,N_9905,N_9676);
nor U10421 (N_10421,N_9841,N_9799);
and U10422 (N_10422,N_9916,N_9973);
and U10423 (N_10423,N_9685,N_9553);
or U10424 (N_10424,N_9510,N_9732);
nor U10425 (N_10425,N_9725,N_9698);
or U10426 (N_10426,N_9954,N_9889);
nand U10427 (N_10427,N_9817,N_9720);
and U10428 (N_10428,N_9763,N_9972);
and U10429 (N_10429,N_9959,N_9822);
or U10430 (N_10430,N_9834,N_9679);
nand U10431 (N_10431,N_9766,N_9687);
and U10432 (N_10432,N_9909,N_9986);
or U10433 (N_10433,N_9793,N_9697);
or U10434 (N_10434,N_9727,N_9630);
or U10435 (N_10435,N_9890,N_9989);
and U10436 (N_10436,N_9510,N_9904);
nor U10437 (N_10437,N_9893,N_9598);
and U10438 (N_10438,N_9711,N_9774);
xnor U10439 (N_10439,N_9822,N_9644);
nand U10440 (N_10440,N_9801,N_9585);
xnor U10441 (N_10441,N_9579,N_9690);
nand U10442 (N_10442,N_9756,N_9510);
and U10443 (N_10443,N_9619,N_9776);
and U10444 (N_10444,N_9573,N_9638);
and U10445 (N_10445,N_9718,N_9900);
nor U10446 (N_10446,N_9797,N_9784);
nor U10447 (N_10447,N_9622,N_9961);
or U10448 (N_10448,N_9907,N_9591);
nand U10449 (N_10449,N_9516,N_9916);
nor U10450 (N_10450,N_9987,N_9701);
nor U10451 (N_10451,N_9966,N_9785);
nor U10452 (N_10452,N_9596,N_9952);
nand U10453 (N_10453,N_9910,N_9968);
xnor U10454 (N_10454,N_9723,N_9646);
xor U10455 (N_10455,N_9880,N_9501);
nor U10456 (N_10456,N_9817,N_9968);
or U10457 (N_10457,N_9962,N_9813);
and U10458 (N_10458,N_9751,N_9839);
or U10459 (N_10459,N_9539,N_9559);
xor U10460 (N_10460,N_9879,N_9807);
xor U10461 (N_10461,N_9563,N_9961);
nor U10462 (N_10462,N_9749,N_9722);
nor U10463 (N_10463,N_9531,N_9816);
xor U10464 (N_10464,N_9793,N_9544);
nand U10465 (N_10465,N_9820,N_9504);
xnor U10466 (N_10466,N_9582,N_9982);
and U10467 (N_10467,N_9527,N_9604);
nor U10468 (N_10468,N_9719,N_9920);
nand U10469 (N_10469,N_9556,N_9613);
or U10470 (N_10470,N_9524,N_9605);
and U10471 (N_10471,N_9835,N_9968);
nor U10472 (N_10472,N_9696,N_9936);
nand U10473 (N_10473,N_9791,N_9899);
or U10474 (N_10474,N_9603,N_9744);
nor U10475 (N_10475,N_9681,N_9760);
nor U10476 (N_10476,N_9527,N_9968);
nand U10477 (N_10477,N_9978,N_9849);
and U10478 (N_10478,N_9684,N_9872);
and U10479 (N_10479,N_9707,N_9750);
xnor U10480 (N_10480,N_9720,N_9591);
and U10481 (N_10481,N_9822,N_9587);
nor U10482 (N_10482,N_9755,N_9569);
and U10483 (N_10483,N_9670,N_9511);
nor U10484 (N_10484,N_9946,N_9775);
nor U10485 (N_10485,N_9894,N_9811);
nand U10486 (N_10486,N_9710,N_9513);
or U10487 (N_10487,N_9767,N_9516);
nand U10488 (N_10488,N_9515,N_9729);
nor U10489 (N_10489,N_9851,N_9600);
nor U10490 (N_10490,N_9968,N_9735);
nand U10491 (N_10491,N_9643,N_9929);
xor U10492 (N_10492,N_9582,N_9878);
or U10493 (N_10493,N_9655,N_9804);
or U10494 (N_10494,N_9754,N_9592);
and U10495 (N_10495,N_9759,N_9865);
nand U10496 (N_10496,N_9904,N_9694);
xor U10497 (N_10497,N_9753,N_9666);
or U10498 (N_10498,N_9825,N_9754);
nand U10499 (N_10499,N_9989,N_9716);
nand U10500 (N_10500,N_10090,N_10214);
or U10501 (N_10501,N_10388,N_10289);
nor U10502 (N_10502,N_10022,N_10242);
xor U10503 (N_10503,N_10279,N_10073);
or U10504 (N_10504,N_10141,N_10127);
xor U10505 (N_10505,N_10470,N_10384);
and U10506 (N_10506,N_10474,N_10266);
xor U10507 (N_10507,N_10259,N_10060);
xor U10508 (N_10508,N_10081,N_10399);
and U10509 (N_10509,N_10114,N_10423);
nor U10510 (N_10510,N_10247,N_10257);
or U10511 (N_10511,N_10430,N_10130);
xor U10512 (N_10512,N_10305,N_10014);
and U10513 (N_10513,N_10164,N_10340);
nor U10514 (N_10514,N_10248,N_10366);
nand U10515 (N_10515,N_10131,N_10333);
xnor U10516 (N_10516,N_10410,N_10211);
or U10517 (N_10517,N_10074,N_10077);
xnor U10518 (N_10518,N_10465,N_10479);
or U10519 (N_10519,N_10491,N_10427);
and U10520 (N_10520,N_10433,N_10346);
nor U10521 (N_10521,N_10380,N_10219);
xor U10522 (N_10522,N_10455,N_10158);
nand U10523 (N_10523,N_10484,N_10237);
nor U10524 (N_10524,N_10405,N_10363);
nor U10525 (N_10525,N_10009,N_10026);
or U10526 (N_10526,N_10300,N_10374);
nor U10527 (N_10527,N_10353,N_10042);
nor U10528 (N_10528,N_10359,N_10162);
and U10529 (N_10529,N_10451,N_10458);
nor U10530 (N_10530,N_10281,N_10370);
nand U10531 (N_10531,N_10093,N_10489);
xor U10532 (N_10532,N_10097,N_10311);
nor U10533 (N_10533,N_10201,N_10082);
or U10534 (N_10534,N_10499,N_10364);
and U10535 (N_10535,N_10239,N_10179);
nor U10536 (N_10536,N_10395,N_10284);
or U10537 (N_10537,N_10061,N_10249);
xnor U10538 (N_10538,N_10347,N_10415);
and U10539 (N_10539,N_10062,N_10016);
and U10540 (N_10540,N_10051,N_10182);
xor U10541 (N_10541,N_10367,N_10029);
or U10542 (N_10542,N_10393,N_10390);
and U10543 (N_10543,N_10025,N_10421);
nor U10544 (N_10544,N_10122,N_10135);
nand U10545 (N_10545,N_10139,N_10002);
nand U10546 (N_10546,N_10027,N_10498);
xnor U10547 (N_10547,N_10050,N_10231);
and U10548 (N_10548,N_10113,N_10208);
nor U10549 (N_10549,N_10270,N_10110);
nor U10550 (N_10550,N_10048,N_10161);
nand U10551 (N_10551,N_10487,N_10024);
xnor U10552 (N_10552,N_10083,N_10315);
nand U10553 (N_10553,N_10040,N_10102);
or U10554 (N_10554,N_10117,N_10381);
or U10555 (N_10555,N_10397,N_10106);
nand U10556 (N_10556,N_10039,N_10291);
or U10557 (N_10557,N_10124,N_10096);
nor U10558 (N_10558,N_10207,N_10243);
or U10559 (N_10559,N_10089,N_10056);
and U10560 (N_10560,N_10168,N_10403);
nor U10561 (N_10561,N_10256,N_10385);
and U10562 (N_10562,N_10358,N_10301);
nand U10563 (N_10563,N_10041,N_10112);
nor U10564 (N_10564,N_10298,N_10453);
nand U10565 (N_10565,N_10345,N_10422);
xnor U10566 (N_10566,N_10375,N_10057);
xor U10567 (N_10567,N_10013,N_10290);
or U10568 (N_10568,N_10398,N_10206);
or U10569 (N_10569,N_10052,N_10120);
and U10570 (N_10570,N_10307,N_10003);
or U10571 (N_10571,N_10235,N_10389);
and U10572 (N_10572,N_10407,N_10138);
nor U10573 (N_10573,N_10007,N_10287);
nor U10574 (N_10574,N_10319,N_10230);
nand U10575 (N_10575,N_10197,N_10037);
nor U10576 (N_10576,N_10222,N_10000);
nor U10577 (N_10577,N_10176,N_10280);
and U10578 (N_10578,N_10303,N_10169);
nand U10579 (N_10579,N_10355,N_10494);
nand U10580 (N_10580,N_10149,N_10323);
nand U10581 (N_10581,N_10084,N_10314);
nand U10582 (N_10582,N_10332,N_10001);
or U10583 (N_10583,N_10456,N_10265);
nor U10584 (N_10584,N_10209,N_10111);
or U10585 (N_10585,N_10163,N_10481);
nand U10586 (N_10586,N_10383,N_10460);
and U10587 (N_10587,N_10473,N_10476);
nand U10588 (N_10588,N_10190,N_10441);
xnor U10589 (N_10589,N_10282,N_10108);
nor U10590 (N_10590,N_10272,N_10070);
and U10591 (N_10591,N_10485,N_10442);
nand U10592 (N_10592,N_10199,N_10251);
or U10593 (N_10593,N_10192,N_10099);
xnor U10594 (N_10594,N_10440,N_10072);
nand U10595 (N_10595,N_10414,N_10254);
nand U10596 (N_10596,N_10264,N_10371);
nor U10597 (N_10597,N_10185,N_10101);
or U10598 (N_10598,N_10086,N_10234);
nor U10599 (N_10599,N_10244,N_10392);
and U10600 (N_10600,N_10053,N_10351);
xor U10601 (N_10601,N_10288,N_10200);
xnor U10602 (N_10602,N_10373,N_10409);
nand U10603 (N_10603,N_10121,N_10140);
and U10604 (N_10604,N_10186,N_10170);
or U10605 (N_10605,N_10262,N_10069);
xnor U10606 (N_10606,N_10233,N_10151);
or U10607 (N_10607,N_10166,N_10401);
or U10608 (N_10608,N_10193,N_10005);
or U10609 (N_10609,N_10335,N_10350);
or U10610 (N_10610,N_10210,N_10324);
nand U10611 (N_10611,N_10361,N_10238);
or U10612 (N_10612,N_10047,N_10480);
or U10613 (N_10613,N_10283,N_10105);
and U10614 (N_10614,N_10461,N_10236);
or U10615 (N_10615,N_10155,N_10225);
nor U10616 (N_10616,N_10495,N_10354);
xor U10617 (N_10617,N_10134,N_10116);
nand U10618 (N_10618,N_10369,N_10276);
or U10619 (N_10619,N_10146,N_10478);
and U10620 (N_10620,N_10420,N_10220);
or U10621 (N_10621,N_10488,N_10376);
or U10622 (N_10622,N_10462,N_10482);
nor U10623 (N_10623,N_10228,N_10100);
nand U10624 (N_10624,N_10203,N_10339);
and U10625 (N_10625,N_10080,N_10469);
or U10626 (N_10626,N_10172,N_10154);
and U10627 (N_10627,N_10277,N_10309);
and U10628 (N_10628,N_10152,N_10028);
nor U10629 (N_10629,N_10360,N_10076);
xnor U10630 (N_10630,N_10142,N_10320);
or U10631 (N_10631,N_10299,N_10258);
nand U10632 (N_10632,N_10180,N_10091);
or U10633 (N_10633,N_10297,N_10269);
nor U10634 (N_10634,N_10221,N_10344);
xnor U10635 (N_10635,N_10377,N_10464);
and U10636 (N_10636,N_10107,N_10044);
nor U10637 (N_10637,N_10012,N_10095);
and U10638 (N_10638,N_10133,N_10349);
and U10639 (N_10639,N_10457,N_10015);
or U10640 (N_10640,N_10011,N_10227);
xnor U10641 (N_10641,N_10125,N_10429);
xor U10642 (N_10642,N_10490,N_10425);
nand U10643 (N_10643,N_10017,N_10246);
nand U10644 (N_10644,N_10098,N_10156);
xor U10645 (N_10645,N_10295,N_10065);
or U10646 (N_10646,N_10318,N_10067);
xor U10647 (N_10647,N_10132,N_10063);
and U10648 (N_10648,N_10436,N_10036);
nor U10649 (N_10649,N_10205,N_10338);
nand U10650 (N_10650,N_10181,N_10471);
nand U10651 (N_10651,N_10342,N_10365);
or U10652 (N_10652,N_10147,N_10159);
nor U10653 (N_10653,N_10202,N_10391);
nor U10654 (N_10654,N_10034,N_10263);
and U10655 (N_10655,N_10337,N_10394);
and U10656 (N_10656,N_10419,N_10454);
or U10657 (N_10657,N_10018,N_10313);
nand U10658 (N_10658,N_10088,N_10126);
or U10659 (N_10659,N_10261,N_10408);
or U10660 (N_10660,N_10217,N_10452);
or U10661 (N_10661,N_10055,N_10432);
nand U10662 (N_10662,N_10123,N_10446);
xnor U10663 (N_10663,N_10068,N_10428);
and U10664 (N_10664,N_10443,N_10326);
nor U10665 (N_10665,N_10020,N_10439);
nor U10666 (N_10666,N_10023,N_10431);
nor U10667 (N_10667,N_10448,N_10218);
and U10668 (N_10668,N_10255,N_10145);
nor U10669 (N_10669,N_10157,N_10341);
and U10670 (N_10670,N_10304,N_10348);
or U10671 (N_10671,N_10136,N_10045);
xor U10672 (N_10672,N_10187,N_10308);
and U10673 (N_10673,N_10165,N_10273);
nor U10674 (N_10674,N_10293,N_10006);
or U10675 (N_10675,N_10387,N_10204);
xnor U10676 (N_10676,N_10396,N_10174);
nor U10677 (N_10677,N_10294,N_10194);
xor U10678 (N_10678,N_10372,N_10330);
and U10679 (N_10679,N_10173,N_10064);
or U10680 (N_10680,N_10467,N_10325);
or U10681 (N_10681,N_10416,N_10412);
nor U10682 (N_10682,N_10215,N_10316);
xnor U10683 (N_10683,N_10066,N_10071);
nor U10684 (N_10684,N_10411,N_10444);
xor U10685 (N_10685,N_10357,N_10144);
or U10686 (N_10686,N_10362,N_10400);
or U10687 (N_10687,N_10224,N_10030);
or U10688 (N_10688,N_10035,N_10085);
xor U10689 (N_10689,N_10477,N_10449);
or U10690 (N_10690,N_10004,N_10038);
xnor U10691 (N_10691,N_10128,N_10223);
nor U10692 (N_10692,N_10368,N_10483);
xor U10693 (N_10693,N_10286,N_10328);
and U10694 (N_10694,N_10497,N_10292);
xor U10695 (N_10695,N_10336,N_10195);
or U10696 (N_10696,N_10115,N_10271);
or U10697 (N_10697,N_10310,N_10404);
nand U10698 (N_10698,N_10008,N_10183);
or U10699 (N_10699,N_10229,N_10213);
nor U10700 (N_10700,N_10232,N_10253);
or U10701 (N_10701,N_10212,N_10317);
nor U10702 (N_10702,N_10417,N_10260);
xor U10703 (N_10703,N_10418,N_10379);
nand U10704 (N_10704,N_10177,N_10196);
nand U10705 (N_10705,N_10267,N_10033);
and U10706 (N_10706,N_10343,N_10463);
nor U10707 (N_10707,N_10321,N_10153);
nand U10708 (N_10708,N_10119,N_10109);
nor U10709 (N_10709,N_10167,N_10486);
nor U10710 (N_10710,N_10043,N_10075);
nor U10711 (N_10711,N_10306,N_10496);
xnor U10712 (N_10712,N_10331,N_10129);
nand U10713 (N_10713,N_10492,N_10059);
nand U10714 (N_10714,N_10058,N_10475);
and U10715 (N_10715,N_10278,N_10493);
and U10716 (N_10716,N_10078,N_10216);
nand U10717 (N_10717,N_10143,N_10092);
or U10718 (N_10718,N_10175,N_10178);
nand U10719 (N_10719,N_10472,N_10447);
xnor U10720 (N_10720,N_10437,N_10296);
nand U10721 (N_10721,N_10302,N_10160);
xnor U10722 (N_10722,N_10184,N_10334);
and U10723 (N_10723,N_10445,N_10468);
xnor U10724 (N_10724,N_10046,N_10049);
xor U10725 (N_10725,N_10275,N_10032);
and U10726 (N_10726,N_10241,N_10434);
or U10727 (N_10727,N_10021,N_10188);
or U10728 (N_10728,N_10189,N_10226);
nor U10729 (N_10729,N_10329,N_10356);
and U10730 (N_10730,N_10378,N_10438);
and U10731 (N_10731,N_10150,N_10386);
nand U10732 (N_10732,N_10352,N_10103);
nor U10733 (N_10733,N_10322,N_10010);
or U10734 (N_10734,N_10054,N_10094);
nand U10735 (N_10735,N_10148,N_10466);
nor U10736 (N_10736,N_10450,N_10191);
and U10737 (N_10737,N_10079,N_10382);
nor U10738 (N_10738,N_10031,N_10087);
nand U10739 (N_10739,N_10459,N_10274);
and U10740 (N_10740,N_10435,N_10171);
and U10741 (N_10741,N_10426,N_10312);
or U10742 (N_10742,N_10413,N_10327);
nor U10743 (N_10743,N_10019,N_10245);
and U10744 (N_10744,N_10137,N_10252);
nor U10745 (N_10745,N_10118,N_10250);
and U10746 (N_10746,N_10104,N_10240);
xor U10747 (N_10747,N_10406,N_10268);
nand U10748 (N_10748,N_10424,N_10402);
or U10749 (N_10749,N_10198,N_10285);
nor U10750 (N_10750,N_10056,N_10181);
nor U10751 (N_10751,N_10312,N_10123);
xor U10752 (N_10752,N_10028,N_10381);
and U10753 (N_10753,N_10495,N_10070);
xor U10754 (N_10754,N_10396,N_10089);
xor U10755 (N_10755,N_10164,N_10248);
or U10756 (N_10756,N_10446,N_10121);
or U10757 (N_10757,N_10324,N_10107);
nand U10758 (N_10758,N_10358,N_10270);
nor U10759 (N_10759,N_10117,N_10270);
or U10760 (N_10760,N_10477,N_10298);
nor U10761 (N_10761,N_10324,N_10337);
nand U10762 (N_10762,N_10014,N_10114);
nand U10763 (N_10763,N_10250,N_10247);
or U10764 (N_10764,N_10206,N_10103);
and U10765 (N_10765,N_10370,N_10005);
or U10766 (N_10766,N_10096,N_10092);
xnor U10767 (N_10767,N_10483,N_10332);
xor U10768 (N_10768,N_10052,N_10031);
and U10769 (N_10769,N_10272,N_10477);
xnor U10770 (N_10770,N_10471,N_10029);
nor U10771 (N_10771,N_10327,N_10168);
nor U10772 (N_10772,N_10066,N_10070);
xor U10773 (N_10773,N_10367,N_10306);
xor U10774 (N_10774,N_10408,N_10003);
or U10775 (N_10775,N_10282,N_10226);
xor U10776 (N_10776,N_10036,N_10393);
or U10777 (N_10777,N_10193,N_10441);
and U10778 (N_10778,N_10320,N_10074);
nor U10779 (N_10779,N_10061,N_10174);
nor U10780 (N_10780,N_10362,N_10471);
or U10781 (N_10781,N_10097,N_10217);
xor U10782 (N_10782,N_10340,N_10024);
nand U10783 (N_10783,N_10091,N_10112);
and U10784 (N_10784,N_10193,N_10307);
and U10785 (N_10785,N_10077,N_10191);
or U10786 (N_10786,N_10028,N_10247);
xor U10787 (N_10787,N_10123,N_10038);
xnor U10788 (N_10788,N_10233,N_10001);
or U10789 (N_10789,N_10069,N_10088);
or U10790 (N_10790,N_10033,N_10118);
nor U10791 (N_10791,N_10035,N_10075);
or U10792 (N_10792,N_10427,N_10200);
or U10793 (N_10793,N_10494,N_10302);
or U10794 (N_10794,N_10263,N_10028);
nand U10795 (N_10795,N_10044,N_10368);
nand U10796 (N_10796,N_10426,N_10214);
nor U10797 (N_10797,N_10236,N_10222);
nand U10798 (N_10798,N_10356,N_10304);
or U10799 (N_10799,N_10069,N_10203);
nor U10800 (N_10800,N_10202,N_10309);
xor U10801 (N_10801,N_10485,N_10473);
and U10802 (N_10802,N_10254,N_10160);
nor U10803 (N_10803,N_10473,N_10364);
nor U10804 (N_10804,N_10168,N_10420);
nand U10805 (N_10805,N_10276,N_10096);
xnor U10806 (N_10806,N_10217,N_10236);
or U10807 (N_10807,N_10056,N_10386);
nor U10808 (N_10808,N_10170,N_10048);
nand U10809 (N_10809,N_10201,N_10014);
xnor U10810 (N_10810,N_10362,N_10001);
xor U10811 (N_10811,N_10214,N_10096);
or U10812 (N_10812,N_10020,N_10172);
xnor U10813 (N_10813,N_10262,N_10473);
xnor U10814 (N_10814,N_10468,N_10356);
nor U10815 (N_10815,N_10285,N_10130);
xor U10816 (N_10816,N_10066,N_10249);
xnor U10817 (N_10817,N_10363,N_10307);
and U10818 (N_10818,N_10446,N_10368);
nand U10819 (N_10819,N_10355,N_10458);
nor U10820 (N_10820,N_10392,N_10296);
nand U10821 (N_10821,N_10461,N_10420);
xor U10822 (N_10822,N_10309,N_10438);
xor U10823 (N_10823,N_10440,N_10124);
or U10824 (N_10824,N_10340,N_10439);
xor U10825 (N_10825,N_10230,N_10119);
or U10826 (N_10826,N_10323,N_10366);
nand U10827 (N_10827,N_10023,N_10435);
xnor U10828 (N_10828,N_10011,N_10188);
nor U10829 (N_10829,N_10382,N_10162);
or U10830 (N_10830,N_10136,N_10360);
and U10831 (N_10831,N_10290,N_10440);
or U10832 (N_10832,N_10289,N_10420);
and U10833 (N_10833,N_10296,N_10245);
xor U10834 (N_10834,N_10082,N_10256);
or U10835 (N_10835,N_10380,N_10462);
nand U10836 (N_10836,N_10211,N_10184);
and U10837 (N_10837,N_10347,N_10266);
xor U10838 (N_10838,N_10341,N_10186);
nand U10839 (N_10839,N_10237,N_10037);
nand U10840 (N_10840,N_10201,N_10249);
or U10841 (N_10841,N_10107,N_10204);
nand U10842 (N_10842,N_10066,N_10043);
nor U10843 (N_10843,N_10421,N_10397);
nor U10844 (N_10844,N_10038,N_10364);
nor U10845 (N_10845,N_10375,N_10234);
xnor U10846 (N_10846,N_10010,N_10294);
nor U10847 (N_10847,N_10465,N_10023);
or U10848 (N_10848,N_10290,N_10399);
and U10849 (N_10849,N_10350,N_10084);
nand U10850 (N_10850,N_10444,N_10490);
and U10851 (N_10851,N_10180,N_10414);
xor U10852 (N_10852,N_10443,N_10344);
nand U10853 (N_10853,N_10382,N_10255);
and U10854 (N_10854,N_10330,N_10473);
or U10855 (N_10855,N_10351,N_10025);
and U10856 (N_10856,N_10288,N_10356);
nand U10857 (N_10857,N_10398,N_10229);
and U10858 (N_10858,N_10010,N_10318);
nand U10859 (N_10859,N_10020,N_10288);
nand U10860 (N_10860,N_10174,N_10122);
or U10861 (N_10861,N_10161,N_10293);
xor U10862 (N_10862,N_10080,N_10356);
xor U10863 (N_10863,N_10447,N_10457);
nor U10864 (N_10864,N_10104,N_10126);
nor U10865 (N_10865,N_10118,N_10108);
and U10866 (N_10866,N_10020,N_10239);
nand U10867 (N_10867,N_10024,N_10372);
and U10868 (N_10868,N_10328,N_10050);
or U10869 (N_10869,N_10060,N_10307);
or U10870 (N_10870,N_10393,N_10193);
or U10871 (N_10871,N_10007,N_10474);
nor U10872 (N_10872,N_10179,N_10022);
xnor U10873 (N_10873,N_10491,N_10303);
and U10874 (N_10874,N_10402,N_10084);
or U10875 (N_10875,N_10377,N_10346);
nor U10876 (N_10876,N_10471,N_10027);
nor U10877 (N_10877,N_10477,N_10169);
and U10878 (N_10878,N_10417,N_10202);
xor U10879 (N_10879,N_10297,N_10119);
nor U10880 (N_10880,N_10276,N_10274);
xor U10881 (N_10881,N_10215,N_10469);
nor U10882 (N_10882,N_10221,N_10118);
or U10883 (N_10883,N_10350,N_10231);
nand U10884 (N_10884,N_10188,N_10148);
nand U10885 (N_10885,N_10109,N_10248);
nand U10886 (N_10886,N_10184,N_10182);
or U10887 (N_10887,N_10167,N_10248);
or U10888 (N_10888,N_10062,N_10434);
or U10889 (N_10889,N_10268,N_10336);
nor U10890 (N_10890,N_10154,N_10096);
xnor U10891 (N_10891,N_10144,N_10115);
nand U10892 (N_10892,N_10066,N_10240);
and U10893 (N_10893,N_10417,N_10489);
nand U10894 (N_10894,N_10478,N_10397);
or U10895 (N_10895,N_10465,N_10403);
or U10896 (N_10896,N_10209,N_10305);
nor U10897 (N_10897,N_10485,N_10180);
and U10898 (N_10898,N_10365,N_10384);
xor U10899 (N_10899,N_10027,N_10253);
nand U10900 (N_10900,N_10270,N_10149);
and U10901 (N_10901,N_10238,N_10320);
nor U10902 (N_10902,N_10047,N_10167);
xnor U10903 (N_10903,N_10195,N_10325);
and U10904 (N_10904,N_10086,N_10228);
and U10905 (N_10905,N_10120,N_10140);
nand U10906 (N_10906,N_10327,N_10316);
xor U10907 (N_10907,N_10266,N_10205);
or U10908 (N_10908,N_10007,N_10481);
nand U10909 (N_10909,N_10426,N_10489);
nor U10910 (N_10910,N_10248,N_10316);
xnor U10911 (N_10911,N_10060,N_10267);
or U10912 (N_10912,N_10337,N_10334);
or U10913 (N_10913,N_10236,N_10026);
or U10914 (N_10914,N_10241,N_10487);
and U10915 (N_10915,N_10480,N_10052);
nor U10916 (N_10916,N_10259,N_10473);
or U10917 (N_10917,N_10239,N_10305);
nand U10918 (N_10918,N_10137,N_10359);
nand U10919 (N_10919,N_10252,N_10169);
nor U10920 (N_10920,N_10360,N_10056);
and U10921 (N_10921,N_10032,N_10166);
nor U10922 (N_10922,N_10086,N_10341);
nor U10923 (N_10923,N_10097,N_10269);
nor U10924 (N_10924,N_10378,N_10144);
or U10925 (N_10925,N_10416,N_10417);
or U10926 (N_10926,N_10214,N_10390);
or U10927 (N_10927,N_10175,N_10406);
xnor U10928 (N_10928,N_10000,N_10416);
and U10929 (N_10929,N_10315,N_10367);
nor U10930 (N_10930,N_10074,N_10310);
or U10931 (N_10931,N_10353,N_10314);
xor U10932 (N_10932,N_10353,N_10313);
and U10933 (N_10933,N_10498,N_10479);
xnor U10934 (N_10934,N_10281,N_10298);
xor U10935 (N_10935,N_10029,N_10290);
nor U10936 (N_10936,N_10246,N_10125);
or U10937 (N_10937,N_10443,N_10368);
nand U10938 (N_10938,N_10272,N_10068);
xor U10939 (N_10939,N_10478,N_10451);
nor U10940 (N_10940,N_10338,N_10223);
nand U10941 (N_10941,N_10177,N_10087);
nor U10942 (N_10942,N_10428,N_10226);
or U10943 (N_10943,N_10400,N_10421);
or U10944 (N_10944,N_10204,N_10478);
or U10945 (N_10945,N_10258,N_10456);
and U10946 (N_10946,N_10440,N_10403);
nor U10947 (N_10947,N_10329,N_10497);
and U10948 (N_10948,N_10473,N_10413);
or U10949 (N_10949,N_10469,N_10301);
xor U10950 (N_10950,N_10321,N_10207);
and U10951 (N_10951,N_10101,N_10457);
and U10952 (N_10952,N_10278,N_10481);
xor U10953 (N_10953,N_10355,N_10031);
or U10954 (N_10954,N_10339,N_10062);
xnor U10955 (N_10955,N_10261,N_10433);
nor U10956 (N_10956,N_10192,N_10301);
nor U10957 (N_10957,N_10459,N_10484);
and U10958 (N_10958,N_10099,N_10283);
or U10959 (N_10959,N_10286,N_10184);
and U10960 (N_10960,N_10148,N_10275);
nand U10961 (N_10961,N_10076,N_10163);
or U10962 (N_10962,N_10192,N_10321);
nand U10963 (N_10963,N_10323,N_10492);
nor U10964 (N_10964,N_10221,N_10171);
nand U10965 (N_10965,N_10000,N_10410);
and U10966 (N_10966,N_10024,N_10132);
and U10967 (N_10967,N_10236,N_10404);
nor U10968 (N_10968,N_10101,N_10455);
xnor U10969 (N_10969,N_10116,N_10363);
and U10970 (N_10970,N_10230,N_10206);
or U10971 (N_10971,N_10122,N_10330);
nor U10972 (N_10972,N_10173,N_10199);
nor U10973 (N_10973,N_10406,N_10251);
xor U10974 (N_10974,N_10494,N_10260);
nand U10975 (N_10975,N_10211,N_10472);
nor U10976 (N_10976,N_10010,N_10383);
nand U10977 (N_10977,N_10303,N_10290);
or U10978 (N_10978,N_10134,N_10449);
nand U10979 (N_10979,N_10408,N_10467);
and U10980 (N_10980,N_10299,N_10286);
nor U10981 (N_10981,N_10215,N_10104);
nor U10982 (N_10982,N_10270,N_10163);
or U10983 (N_10983,N_10466,N_10145);
or U10984 (N_10984,N_10494,N_10293);
and U10985 (N_10985,N_10286,N_10195);
nor U10986 (N_10986,N_10347,N_10346);
nor U10987 (N_10987,N_10319,N_10398);
nor U10988 (N_10988,N_10183,N_10232);
nor U10989 (N_10989,N_10372,N_10025);
nor U10990 (N_10990,N_10111,N_10208);
nor U10991 (N_10991,N_10296,N_10043);
xnor U10992 (N_10992,N_10449,N_10401);
nand U10993 (N_10993,N_10058,N_10335);
xnor U10994 (N_10994,N_10135,N_10159);
nor U10995 (N_10995,N_10287,N_10277);
nor U10996 (N_10996,N_10492,N_10462);
nand U10997 (N_10997,N_10370,N_10270);
nand U10998 (N_10998,N_10088,N_10269);
and U10999 (N_10999,N_10436,N_10350);
nand U11000 (N_11000,N_10991,N_10740);
and U11001 (N_11001,N_10751,N_10502);
nand U11002 (N_11002,N_10772,N_10704);
xnor U11003 (N_11003,N_10800,N_10706);
xnor U11004 (N_11004,N_10965,N_10955);
nor U11005 (N_11005,N_10849,N_10983);
and U11006 (N_11006,N_10789,N_10691);
nor U11007 (N_11007,N_10805,N_10945);
nor U11008 (N_11008,N_10899,N_10645);
nand U11009 (N_11009,N_10911,N_10625);
nor U11010 (N_11010,N_10641,N_10501);
and U11011 (N_11011,N_10560,N_10700);
and U11012 (N_11012,N_10540,N_10715);
xor U11013 (N_11013,N_10635,N_10898);
nor U11014 (N_11014,N_10707,N_10595);
nor U11015 (N_11015,N_10782,N_10949);
xor U11016 (N_11016,N_10537,N_10923);
xnor U11017 (N_11017,N_10827,N_10950);
nor U11018 (N_11018,N_10576,N_10790);
nor U11019 (N_11019,N_10640,N_10663);
or U11020 (N_11020,N_10791,N_10553);
and U11021 (N_11021,N_10703,N_10749);
xor U11022 (N_11022,N_10906,N_10729);
or U11023 (N_11023,N_10676,N_10655);
or U11024 (N_11024,N_10508,N_10738);
xnor U11025 (N_11025,N_10781,N_10986);
nor U11026 (N_11026,N_10727,N_10889);
nor U11027 (N_11027,N_10821,N_10522);
or U11028 (N_11028,N_10633,N_10823);
and U11029 (N_11029,N_10555,N_10910);
nor U11030 (N_11030,N_10828,N_10961);
nand U11031 (N_11031,N_10932,N_10505);
nor U11032 (N_11032,N_10632,N_10539);
nand U11033 (N_11033,N_10708,N_10993);
xor U11034 (N_11034,N_10658,N_10756);
nand U11035 (N_11035,N_10669,N_10973);
and U11036 (N_11036,N_10531,N_10812);
nor U11037 (N_11037,N_10615,N_10690);
and U11038 (N_11038,N_10673,N_10594);
xor U11039 (N_11039,N_10864,N_10754);
xnor U11040 (N_11040,N_10928,N_10847);
or U11041 (N_11041,N_10734,N_10867);
nand U11042 (N_11042,N_10830,N_10564);
xor U11043 (N_11043,N_10880,N_10649);
nor U11044 (N_11044,N_10612,N_10848);
nand U11045 (N_11045,N_10688,N_10523);
xnor U11046 (N_11046,N_10692,N_10783);
xor U11047 (N_11047,N_10992,N_10631);
nand U11048 (N_11048,N_10872,N_10826);
and U11049 (N_11049,N_10512,N_10750);
nor U11050 (N_11050,N_10574,N_10988);
nand U11051 (N_11051,N_10536,N_10568);
or U11052 (N_11052,N_10682,N_10657);
and U11053 (N_11053,N_10905,N_10630);
xor U11054 (N_11054,N_10580,N_10908);
nor U11055 (N_11055,N_10759,N_10882);
xor U11056 (N_11056,N_10689,N_10694);
or U11057 (N_11057,N_10546,N_10760);
xnor U11058 (N_11058,N_10958,N_10987);
or U11059 (N_11059,N_10600,N_10963);
nand U11060 (N_11060,N_10968,N_10693);
and U11061 (N_11061,N_10709,N_10593);
nand U11062 (N_11062,N_10775,N_10578);
and U11063 (N_11063,N_10535,N_10811);
nor U11064 (N_11064,N_10995,N_10582);
xor U11065 (N_11065,N_10935,N_10562);
or U11066 (N_11066,N_10721,N_10770);
nand U11067 (N_11067,N_10556,N_10807);
nand U11068 (N_11068,N_10589,N_10852);
xor U11069 (N_11069,N_10953,N_10617);
xor U11070 (N_11070,N_10662,N_10808);
and U11071 (N_11071,N_10552,N_10607);
or U11072 (N_11072,N_10611,N_10804);
or U11073 (N_11073,N_10944,N_10571);
nor U11074 (N_11074,N_10897,N_10936);
nand U11075 (N_11075,N_10695,N_10894);
nor U11076 (N_11076,N_10855,N_10887);
xor U11077 (N_11077,N_10860,N_10835);
and U11078 (N_11078,N_10724,N_10976);
or U11079 (N_11079,N_10646,N_10573);
nand U11080 (N_11080,N_10836,N_10744);
nor U11081 (N_11081,N_10597,N_10957);
and U11082 (N_11082,N_10529,N_10981);
and U11083 (N_11083,N_10996,N_10519);
or U11084 (N_11084,N_10650,N_10506);
or U11085 (N_11085,N_10865,N_10551);
xnor U11086 (N_11086,N_10956,N_10664);
nor U11087 (N_11087,N_10975,N_10858);
and U11088 (N_11088,N_10873,N_10614);
xor U11089 (N_11089,N_10565,N_10814);
or U11090 (N_11090,N_10798,N_10851);
xnor U11091 (N_11091,N_10675,N_10659);
xor U11092 (N_11092,N_10525,N_10773);
and U11093 (N_11093,N_10974,N_10888);
nand U11094 (N_11094,N_10603,N_10609);
or U11095 (N_11095,N_10970,N_10857);
and U11096 (N_11096,N_10696,N_10710);
and U11097 (N_11097,N_10871,N_10656);
or U11098 (N_11098,N_10969,N_10748);
and U11099 (N_11099,N_10538,N_10904);
nand U11100 (N_11100,N_10838,N_10892);
nor U11101 (N_11101,N_10731,N_10862);
xnor U11102 (N_11102,N_10639,N_10672);
nor U11103 (N_11103,N_10515,N_10739);
nand U11104 (N_11104,N_10528,N_10843);
nor U11105 (N_11105,N_10629,N_10642);
nor U11106 (N_11106,N_10792,N_10559);
xnor U11107 (N_11107,N_10776,N_10705);
and U11108 (N_11108,N_10893,N_10841);
or U11109 (N_11109,N_10507,N_10520);
xor U11110 (N_11110,N_10686,N_10541);
nand U11111 (N_11111,N_10926,N_10765);
xor U11112 (N_11112,N_10952,N_10997);
nor U11113 (N_11113,N_10984,N_10511);
nand U11114 (N_11114,N_10517,N_10876);
nand U11115 (N_11115,N_10769,N_10521);
and U11116 (N_11116,N_10624,N_10934);
nand U11117 (N_11117,N_10803,N_10883);
or U11118 (N_11118,N_10766,N_10549);
xnor U11119 (N_11119,N_10667,N_10654);
nor U11120 (N_11120,N_10683,N_10621);
nor U11121 (N_11121,N_10854,N_10687);
nor U11122 (N_11122,N_10819,N_10543);
nor U11123 (N_11123,N_10728,N_10570);
xor U11124 (N_11124,N_10563,N_10581);
and U11125 (N_11125,N_10868,N_10637);
and U11126 (N_11126,N_10985,N_10885);
nand U11127 (N_11127,N_10891,N_10752);
nor U11128 (N_11128,N_10813,N_10757);
nor U11129 (N_11129,N_10636,N_10758);
nor U11130 (N_11130,N_10532,N_10712);
nor U11131 (N_11131,N_10810,N_10665);
or U11132 (N_11132,N_10567,N_10701);
nand U11133 (N_11133,N_10774,N_10939);
nor U11134 (N_11134,N_10685,N_10504);
nor U11135 (N_11135,N_10833,N_10741);
or U11136 (N_11136,N_10959,N_10998);
or U11137 (N_11137,N_10550,N_10954);
and U11138 (N_11138,N_10920,N_10542);
or U11139 (N_11139,N_10747,N_10626);
or U11140 (N_11140,N_10585,N_10534);
and U11141 (N_11141,N_10746,N_10711);
or U11142 (N_11142,N_10972,N_10861);
nand U11143 (N_11143,N_10586,N_10768);
or U11144 (N_11144,N_10616,N_10764);
xor U11145 (N_11145,N_10743,N_10591);
nor U11146 (N_11146,N_10797,N_10733);
nor U11147 (N_11147,N_10584,N_10620);
and U11148 (N_11148,N_10674,N_10762);
or U11149 (N_11149,N_10719,N_10948);
nand U11150 (N_11150,N_10583,N_10726);
nor U11151 (N_11151,N_10648,N_10527);
nor U11152 (N_11152,N_10503,N_10869);
or U11153 (N_11153,N_10702,N_10666);
xor U11154 (N_11154,N_10572,N_10671);
and U11155 (N_11155,N_10599,N_10767);
and U11156 (N_11156,N_10856,N_10921);
nand U11157 (N_11157,N_10784,N_10575);
xor U11158 (N_11158,N_10561,N_10647);
or U11159 (N_11159,N_10548,N_10837);
nand U11160 (N_11160,N_10755,N_10994);
xor U11161 (N_11161,N_10802,N_10951);
or U11162 (N_11162,N_10788,N_10643);
xor U11163 (N_11163,N_10979,N_10787);
or U11164 (N_11164,N_10853,N_10866);
and U11165 (N_11165,N_10518,N_10623);
or U11166 (N_11166,N_10627,N_10877);
or U11167 (N_11167,N_10638,N_10907);
xnor U11168 (N_11168,N_10793,N_10634);
or U11169 (N_11169,N_10879,N_10681);
and U11170 (N_11170,N_10592,N_10924);
nand U11171 (N_11171,N_10832,N_10874);
xnor U11172 (N_11172,N_10844,N_10806);
xnor U11173 (N_11173,N_10780,N_10510);
nand U11174 (N_11174,N_10699,N_10713);
nand U11175 (N_11175,N_10735,N_10863);
nor U11176 (N_11176,N_10610,N_10809);
xor U11177 (N_11177,N_10799,N_10516);
nand U11178 (N_11178,N_10778,N_10794);
and U11179 (N_11179,N_10929,N_10698);
or U11180 (N_11180,N_10547,N_10668);
xor U11181 (N_11181,N_10901,N_10557);
nor U11182 (N_11182,N_10825,N_10895);
and U11183 (N_11183,N_10596,N_10509);
or U11184 (N_11184,N_10818,N_10622);
and U11185 (N_11185,N_10918,N_10941);
xor U11186 (N_11186,N_10903,N_10661);
or U11187 (N_11187,N_10608,N_10777);
nor U11188 (N_11188,N_10902,N_10822);
and U11189 (N_11189,N_10930,N_10878);
or U11190 (N_11190,N_10737,N_10978);
nand U11191 (N_11191,N_10846,N_10618);
xor U11192 (N_11192,N_10881,N_10915);
nand U11193 (N_11193,N_10619,N_10913);
xor U11194 (N_11194,N_10900,N_10697);
or U11195 (N_11195,N_10566,N_10628);
nand U11196 (N_11196,N_10919,N_10514);
xnor U11197 (N_11197,N_10989,N_10653);
nand U11198 (N_11198,N_10717,N_10533);
nand U11199 (N_11199,N_10530,N_10545);
or U11200 (N_11200,N_10587,N_10500);
or U11201 (N_11201,N_10786,N_10684);
or U11202 (N_11202,N_10933,N_10670);
and U11203 (N_11203,N_10980,N_10912);
nand U11204 (N_11204,N_10723,N_10820);
xor U11205 (N_11205,N_10815,N_10937);
and U11206 (N_11206,N_10613,N_10962);
nand U11207 (N_11207,N_10725,N_10999);
and U11208 (N_11208,N_10753,N_10524);
xnor U11209 (N_11209,N_10842,N_10736);
xnor U11210 (N_11210,N_10716,N_10795);
and U11211 (N_11211,N_10817,N_10971);
nor U11212 (N_11212,N_10890,N_10884);
xnor U11213 (N_11213,N_10678,N_10982);
xor U11214 (N_11214,N_10644,N_10834);
xnor U11215 (N_11215,N_10839,N_10745);
or U11216 (N_11216,N_10742,N_10680);
nand U11217 (N_11217,N_10569,N_10870);
or U11218 (N_11218,N_10829,N_10677);
and U11219 (N_11219,N_10925,N_10602);
nor U11220 (N_11220,N_10558,N_10605);
or U11221 (N_11221,N_10922,N_10914);
or U11222 (N_11222,N_10845,N_10960);
and U11223 (N_11223,N_10601,N_10886);
nand U11224 (N_11224,N_10917,N_10947);
and U11225 (N_11225,N_10824,N_10577);
and U11226 (N_11226,N_10720,N_10718);
nor U11227 (N_11227,N_10943,N_10785);
and U11228 (N_11228,N_10554,N_10801);
and U11229 (N_11229,N_10938,N_10590);
nand U11230 (N_11230,N_10544,N_10840);
or U11231 (N_11231,N_10763,N_10732);
and U11232 (N_11232,N_10604,N_10940);
and U11233 (N_11233,N_10660,N_10896);
or U11234 (N_11234,N_10977,N_10771);
nand U11235 (N_11235,N_10850,N_10598);
xnor U11236 (N_11236,N_10579,N_10916);
xnor U11237 (N_11237,N_10714,N_10816);
or U11238 (N_11238,N_10796,N_10651);
nor U11239 (N_11239,N_10513,N_10722);
and U11240 (N_11240,N_10946,N_10859);
nand U11241 (N_11241,N_10779,N_10931);
nor U11242 (N_11242,N_10606,N_10966);
and U11243 (N_11243,N_10875,N_10679);
and U11244 (N_11244,N_10927,N_10909);
nor U11245 (N_11245,N_10761,N_10964);
nor U11246 (N_11246,N_10730,N_10942);
nor U11247 (N_11247,N_10990,N_10526);
nor U11248 (N_11248,N_10588,N_10967);
and U11249 (N_11249,N_10831,N_10652);
nand U11250 (N_11250,N_10914,N_10873);
and U11251 (N_11251,N_10928,N_10526);
xor U11252 (N_11252,N_10736,N_10685);
or U11253 (N_11253,N_10607,N_10711);
nand U11254 (N_11254,N_10793,N_10857);
nand U11255 (N_11255,N_10644,N_10717);
or U11256 (N_11256,N_10611,N_10989);
and U11257 (N_11257,N_10592,N_10744);
xor U11258 (N_11258,N_10775,N_10831);
or U11259 (N_11259,N_10583,N_10920);
or U11260 (N_11260,N_10708,N_10992);
and U11261 (N_11261,N_10778,N_10758);
or U11262 (N_11262,N_10791,N_10812);
and U11263 (N_11263,N_10823,N_10868);
nor U11264 (N_11264,N_10792,N_10720);
nand U11265 (N_11265,N_10863,N_10542);
or U11266 (N_11266,N_10573,N_10529);
or U11267 (N_11267,N_10628,N_10993);
nand U11268 (N_11268,N_10787,N_10905);
nand U11269 (N_11269,N_10693,N_10591);
xnor U11270 (N_11270,N_10651,N_10702);
or U11271 (N_11271,N_10931,N_10936);
or U11272 (N_11272,N_10774,N_10771);
xnor U11273 (N_11273,N_10976,N_10504);
or U11274 (N_11274,N_10867,N_10791);
or U11275 (N_11275,N_10757,N_10954);
nor U11276 (N_11276,N_10623,N_10890);
or U11277 (N_11277,N_10969,N_10822);
xnor U11278 (N_11278,N_10816,N_10705);
xor U11279 (N_11279,N_10990,N_10695);
nor U11280 (N_11280,N_10914,N_10935);
xnor U11281 (N_11281,N_10773,N_10942);
or U11282 (N_11282,N_10693,N_10658);
xnor U11283 (N_11283,N_10518,N_10516);
or U11284 (N_11284,N_10995,N_10736);
or U11285 (N_11285,N_10549,N_10765);
xnor U11286 (N_11286,N_10674,N_10879);
and U11287 (N_11287,N_10964,N_10515);
nor U11288 (N_11288,N_10515,N_10996);
or U11289 (N_11289,N_10663,N_10709);
xnor U11290 (N_11290,N_10825,N_10961);
nor U11291 (N_11291,N_10636,N_10594);
and U11292 (N_11292,N_10529,N_10757);
or U11293 (N_11293,N_10542,N_10654);
or U11294 (N_11294,N_10987,N_10685);
or U11295 (N_11295,N_10595,N_10824);
xnor U11296 (N_11296,N_10788,N_10586);
xnor U11297 (N_11297,N_10873,N_10797);
nor U11298 (N_11298,N_10813,N_10796);
nor U11299 (N_11299,N_10757,N_10775);
nor U11300 (N_11300,N_10716,N_10946);
nand U11301 (N_11301,N_10965,N_10689);
or U11302 (N_11302,N_10564,N_10789);
nand U11303 (N_11303,N_10973,N_10821);
nor U11304 (N_11304,N_10509,N_10830);
nor U11305 (N_11305,N_10900,N_10680);
and U11306 (N_11306,N_10549,N_10762);
xor U11307 (N_11307,N_10780,N_10756);
and U11308 (N_11308,N_10751,N_10813);
and U11309 (N_11309,N_10655,N_10713);
nor U11310 (N_11310,N_10547,N_10736);
or U11311 (N_11311,N_10936,N_10985);
xor U11312 (N_11312,N_10792,N_10747);
or U11313 (N_11313,N_10692,N_10926);
xor U11314 (N_11314,N_10862,N_10885);
or U11315 (N_11315,N_10710,N_10865);
nor U11316 (N_11316,N_10514,N_10746);
xnor U11317 (N_11317,N_10977,N_10556);
nor U11318 (N_11318,N_10794,N_10982);
nor U11319 (N_11319,N_10794,N_10926);
xor U11320 (N_11320,N_10758,N_10923);
nand U11321 (N_11321,N_10922,N_10830);
or U11322 (N_11322,N_10594,N_10815);
or U11323 (N_11323,N_10685,N_10879);
and U11324 (N_11324,N_10556,N_10728);
or U11325 (N_11325,N_10796,N_10512);
and U11326 (N_11326,N_10669,N_10975);
or U11327 (N_11327,N_10889,N_10956);
nor U11328 (N_11328,N_10988,N_10964);
nand U11329 (N_11329,N_10635,N_10568);
nand U11330 (N_11330,N_10768,N_10640);
nand U11331 (N_11331,N_10970,N_10568);
nor U11332 (N_11332,N_10859,N_10616);
nor U11333 (N_11333,N_10687,N_10703);
nor U11334 (N_11334,N_10751,N_10922);
xor U11335 (N_11335,N_10889,N_10700);
or U11336 (N_11336,N_10928,N_10797);
nor U11337 (N_11337,N_10561,N_10977);
nand U11338 (N_11338,N_10546,N_10543);
nor U11339 (N_11339,N_10840,N_10775);
or U11340 (N_11340,N_10750,N_10834);
and U11341 (N_11341,N_10630,N_10650);
and U11342 (N_11342,N_10585,N_10524);
nand U11343 (N_11343,N_10752,N_10884);
nand U11344 (N_11344,N_10676,N_10543);
xor U11345 (N_11345,N_10502,N_10741);
and U11346 (N_11346,N_10940,N_10531);
nand U11347 (N_11347,N_10610,N_10512);
xor U11348 (N_11348,N_10952,N_10798);
nor U11349 (N_11349,N_10704,N_10553);
nor U11350 (N_11350,N_10687,N_10869);
or U11351 (N_11351,N_10996,N_10743);
xnor U11352 (N_11352,N_10834,N_10537);
xor U11353 (N_11353,N_10557,N_10735);
nor U11354 (N_11354,N_10832,N_10664);
nor U11355 (N_11355,N_10509,N_10965);
xor U11356 (N_11356,N_10782,N_10514);
and U11357 (N_11357,N_10577,N_10503);
nand U11358 (N_11358,N_10794,N_10780);
nand U11359 (N_11359,N_10515,N_10609);
or U11360 (N_11360,N_10903,N_10746);
and U11361 (N_11361,N_10677,N_10750);
nor U11362 (N_11362,N_10983,N_10824);
nand U11363 (N_11363,N_10661,N_10654);
xor U11364 (N_11364,N_10830,N_10763);
nor U11365 (N_11365,N_10969,N_10943);
xor U11366 (N_11366,N_10948,N_10953);
or U11367 (N_11367,N_10952,N_10530);
and U11368 (N_11368,N_10580,N_10634);
nor U11369 (N_11369,N_10971,N_10895);
nor U11370 (N_11370,N_10685,N_10639);
or U11371 (N_11371,N_10501,N_10992);
nand U11372 (N_11372,N_10587,N_10531);
and U11373 (N_11373,N_10947,N_10908);
nand U11374 (N_11374,N_10790,N_10694);
nor U11375 (N_11375,N_10986,N_10541);
and U11376 (N_11376,N_10960,N_10899);
xor U11377 (N_11377,N_10822,N_10901);
and U11378 (N_11378,N_10721,N_10976);
or U11379 (N_11379,N_10859,N_10541);
nor U11380 (N_11380,N_10979,N_10820);
nand U11381 (N_11381,N_10526,N_10794);
or U11382 (N_11382,N_10936,N_10829);
and U11383 (N_11383,N_10895,N_10507);
or U11384 (N_11384,N_10958,N_10959);
and U11385 (N_11385,N_10568,N_10978);
or U11386 (N_11386,N_10714,N_10673);
or U11387 (N_11387,N_10894,N_10829);
xnor U11388 (N_11388,N_10834,N_10717);
xnor U11389 (N_11389,N_10876,N_10916);
nor U11390 (N_11390,N_10825,N_10980);
and U11391 (N_11391,N_10568,N_10504);
nor U11392 (N_11392,N_10890,N_10923);
and U11393 (N_11393,N_10948,N_10945);
nor U11394 (N_11394,N_10595,N_10999);
xnor U11395 (N_11395,N_10737,N_10991);
xnor U11396 (N_11396,N_10949,N_10950);
nor U11397 (N_11397,N_10739,N_10631);
nand U11398 (N_11398,N_10636,N_10554);
nand U11399 (N_11399,N_10975,N_10883);
nand U11400 (N_11400,N_10954,N_10747);
or U11401 (N_11401,N_10850,N_10605);
or U11402 (N_11402,N_10786,N_10852);
xor U11403 (N_11403,N_10662,N_10611);
nor U11404 (N_11404,N_10883,N_10931);
xor U11405 (N_11405,N_10777,N_10888);
xor U11406 (N_11406,N_10698,N_10856);
nand U11407 (N_11407,N_10841,N_10677);
xor U11408 (N_11408,N_10944,N_10631);
and U11409 (N_11409,N_10999,N_10767);
xor U11410 (N_11410,N_10710,N_10533);
or U11411 (N_11411,N_10621,N_10722);
nor U11412 (N_11412,N_10722,N_10754);
nor U11413 (N_11413,N_10637,N_10610);
and U11414 (N_11414,N_10969,N_10992);
or U11415 (N_11415,N_10928,N_10551);
and U11416 (N_11416,N_10965,N_10720);
or U11417 (N_11417,N_10837,N_10666);
and U11418 (N_11418,N_10999,N_10947);
nand U11419 (N_11419,N_10691,N_10869);
xor U11420 (N_11420,N_10875,N_10590);
nand U11421 (N_11421,N_10735,N_10762);
xor U11422 (N_11422,N_10906,N_10563);
xnor U11423 (N_11423,N_10722,N_10598);
xnor U11424 (N_11424,N_10685,N_10615);
and U11425 (N_11425,N_10906,N_10749);
xor U11426 (N_11426,N_10887,N_10946);
nor U11427 (N_11427,N_10599,N_10801);
xor U11428 (N_11428,N_10780,N_10867);
and U11429 (N_11429,N_10920,N_10785);
nand U11430 (N_11430,N_10749,N_10800);
or U11431 (N_11431,N_10900,N_10505);
nand U11432 (N_11432,N_10550,N_10810);
nand U11433 (N_11433,N_10814,N_10512);
or U11434 (N_11434,N_10752,N_10836);
nand U11435 (N_11435,N_10575,N_10870);
xnor U11436 (N_11436,N_10805,N_10542);
xnor U11437 (N_11437,N_10929,N_10991);
and U11438 (N_11438,N_10511,N_10624);
and U11439 (N_11439,N_10681,N_10973);
nand U11440 (N_11440,N_10544,N_10702);
xor U11441 (N_11441,N_10903,N_10727);
or U11442 (N_11442,N_10989,N_10767);
and U11443 (N_11443,N_10846,N_10862);
nor U11444 (N_11444,N_10645,N_10596);
or U11445 (N_11445,N_10900,N_10935);
and U11446 (N_11446,N_10865,N_10514);
nor U11447 (N_11447,N_10967,N_10926);
nand U11448 (N_11448,N_10850,N_10622);
or U11449 (N_11449,N_10937,N_10649);
nor U11450 (N_11450,N_10809,N_10515);
nand U11451 (N_11451,N_10686,N_10679);
nor U11452 (N_11452,N_10627,N_10784);
nor U11453 (N_11453,N_10842,N_10881);
nor U11454 (N_11454,N_10714,N_10708);
nor U11455 (N_11455,N_10887,N_10812);
xnor U11456 (N_11456,N_10709,N_10646);
xor U11457 (N_11457,N_10969,N_10710);
or U11458 (N_11458,N_10716,N_10894);
or U11459 (N_11459,N_10701,N_10811);
nand U11460 (N_11460,N_10998,N_10745);
and U11461 (N_11461,N_10555,N_10805);
nor U11462 (N_11462,N_10697,N_10706);
xor U11463 (N_11463,N_10699,N_10574);
and U11464 (N_11464,N_10513,N_10989);
xor U11465 (N_11465,N_10622,N_10857);
or U11466 (N_11466,N_10938,N_10594);
or U11467 (N_11467,N_10637,N_10586);
or U11468 (N_11468,N_10936,N_10786);
or U11469 (N_11469,N_10993,N_10543);
or U11470 (N_11470,N_10745,N_10608);
or U11471 (N_11471,N_10893,N_10945);
nand U11472 (N_11472,N_10722,N_10556);
and U11473 (N_11473,N_10723,N_10802);
xor U11474 (N_11474,N_10797,N_10771);
nand U11475 (N_11475,N_10517,N_10754);
and U11476 (N_11476,N_10586,N_10600);
and U11477 (N_11477,N_10555,N_10556);
and U11478 (N_11478,N_10603,N_10944);
and U11479 (N_11479,N_10926,N_10521);
and U11480 (N_11480,N_10863,N_10910);
nor U11481 (N_11481,N_10942,N_10908);
nand U11482 (N_11482,N_10849,N_10827);
nand U11483 (N_11483,N_10544,N_10737);
or U11484 (N_11484,N_10772,N_10592);
or U11485 (N_11485,N_10991,N_10916);
nand U11486 (N_11486,N_10889,N_10959);
and U11487 (N_11487,N_10819,N_10800);
nand U11488 (N_11488,N_10923,N_10754);
or U11489 (N_11489,N_10652,N_10525);
or U11490 (N_11490,N_10597,N_10580);
and U11491 (N_11491,N_10993,N_10989);
or U11492 (N_11492,N_10650,N_10862);
xor U11493 (N_11493,N_10562,N_10861);
and U11494 (N_11494,N_10949,N_10691);
or U11495 (N_11495,N_10501,N_10960);
nand U11496 (N_11496,N_10521,N_10826);
or U11497 (N_11497,N_10665,N_10970);
and U11498 (N_11498,N_10721,N_10518);
or U11499 (N_11499,N_10900,N_10724);
xor U11500 (N_11500,N_11008,N_11011);
or U11501 (N_11501,N_11143,N_11004);
or U11502 (N_11502,N_11262,N_11351);
and U11503 (N_11503,N_11325,N_11141);
xnor U11504 (N_11504,N_11232,N_11222);
xnor U11505 (N_11505,N_11120,N_11314);
nand U11506 (N_11506,N_11181,N_11253);
or U11507 (N_11507,N_11461,N_11256);
or U11508 (N_11508,N_11052,N_11311);
or U11509 (N_11509,N_11341,N_11303);
nor U11510 (N_11510,N_11286,N_11006);
xnor U11511 (N_11511,N_11049,N_11000);
nor U11512 (N_11512,N_11276,N_11496);
and U11513 (N_11513,N_11147,N_11072);
nand U11514 (N_11514,N_11384,N_11194);
xnor U11515 (N_11515,N_11137,N_11283);
nand U11516 (N_11516,N_11162,N_11487);
nor U11517 (N_11517,N_11345,N_11423);
nor U11518 (N_11518,N_11178,N_11398);
nand U11519 (N_11519,N_11173,N_11393);
nand U11520 (N_11520,N_11266,N_11333);
xnor U11521 (N_11521,N_11105,N_11148);
nor U11522 (N_11522,N_11484,N_11458);
nor U11523 (N_11523,N_11473,N_11093);
or U11524 (N_11524,N_11056,N_11323);
and U11525 (N_11525,N_11350,N_11275);
and U11526 (N_11526,N_11490,N_11434);
nor U11527 (N_11527,N_11277,N_11353);
xnor U11528 (N_11528,N_11339,N_11357);
nor U11529 (N_11529,N_11269,N_11344);
and U11530 (N_11530,N_11376,N_11374);
nand U11531 (N_11531,N_11085,N_11227);
nor U11532 (N_11532,N_11214,N_11456);
xor U11533 (N_11533,N_11245,N_11302);
or U11534 (N_11534,N_11444,N_11083);
nand U11535 (N_11535,N_11103,N_11386);
nor U11536 (N_11536,N_11097,N_11062);
and U11537 (N_11537,N_11205,N_11310);
or U11538 (N_11538,N_11439,N_11076);
and U11539 (N_11539,N_11322,N_11098);
nor U11540 (N_11540,N_11370,N_11243);
and U11541 (N_11541,N_11217,N_11047);
and U11542 (N_11542,N_11027,N_11328);
nand U11543 (N_11543,N_11356,N_11365);
and U11544 (N_11544,N_11415,N_11051);
and U11545 (N_11545,N_11016,N_11079);
and U11546 (N_11546,N_11193,N_11208);
nand U11547 (N_11547,N_11175,N_11142);
or U11548 (N_11548,N_11034,N_11369);
nor U11549 (N_11549,N_11089,N_11424);
xnor U11550 (N_11550,N_11371,N_11126);
nand U11551 (N_11551,N_11234,N_11019);
xnor U11552 (N_11552,N_11184,N_11071);
nand U11553 (N_11553,N_11191,N_11028);
or U11554 (N_11554,N_11426,N_11244);
xnor U11555 (N_11555,N_11497,N_11338);
xnor U11556 (N_11556,N_11037,N_11468);
and U11557 (N_11557,N_11239,N_11372);
nor U11558 (N_11558,N_11088,N_11274);
or U11559 (N_11559,N_11154,N_11287);
xor U11560 (N_11560,N_11235,N_11094);
xnor U11561 (N_11561,N_11130,N_11259);
or U11562 (N_11562,N_11348,N_11242);
and U11563 (N_11563,N_11430,N_11488);
or U11564 (N_11564,N_11293,N_11395);
or U11565 (N_11565,N_11321,N_11122);
and U11566 (N_11566,N_11409,N_11313);
xor U11567 (N_11567,N_11144,N_11421);
nor U11568 (N_11568,N_11331,N_11174);
nand U11569 (N_11569,N_11260,N_11419);
or U11570 (N_11570,N_11161,N_11200);
or U11571 (N_11571,N_11138,N_11009);
nor U11572 (N_11572,N_11149,N_11020);
and U11573 (N_11573,N_11319,N_11084);
or U11574 (N_11574,N_11204,N_11474);
or U11575 (N_11575,N_11078,N_11170);
and U11576 (N_11576,N_11166,N_11045);
xnor U11577 (N_11577,N_11192,N_11146);
nor U11578 (N_11578,N_11157,N_11383);
nor U11579 (N_11579,N_11493,N_11249);
and U11580 (N_11580,N_11414,N_11437);
and U11581 (N_11581,N_11063,N_11317);
nand U11582 (N_11582,N_11460,N_11332);
nand U11583 (N_11583,N_11377,N_11452);
or U11584 (N_11584,N_11258,N_11254);
and U11585 (N_11585,N_11381,N_11436);
nand U11586 (N_11586,N_11033,N_11199);
nor U11587 (N_11587,N_11448,N_11038);
nand U11588 (N_11588,N_11366,N_11400);
nand U11589 (N_11589,N_11086,N_11113);
nand U11590 (N_11590,N_11077,N_11355);
nand U11591 (N_11591,N_11268,N_11050);
and U11592 (N_11592,N_11305,N_11104);
nand U11593 (N_11593,N_11307,N_11003);
xor U11594 (N_11594,N_11058,N_11330);
xor U11595 (N_11595,N_11294,N_11462);
or U11596 (N_11596,N_11443,N_11112);
or U11597 (N_11597,N_11335,N_11030);
nand U11598 (N_11598,N_11136,N_11291);
nor U11599 (N_11599,N_11359,N_11225);
and U11600 (N_11600,N_11091,N_11196);
and U11601 (N_11601,N_11096,N_11403);
nand U11602 (N_11602,N_11435,N_11485);
and U11603 (N_11603,N_11354,N_11111);
xor U11604 (N_11604,N_11282,N_11476);
and U11605 (N_11605,N_11236,N_11080);
nand U11606 (N_11606,N_11228,N_11151);
and U11607 (N_11607,N_11429,N_11233);
nor U11608 (N_11608,N_11231,N_11406);
xor U11609 (N_11609,N_11186,N_11095);
xor U11610 (N_11610,N_11055,N_11402);
or U11611 (N_11611,N_11257,N_11117);
xnor U11612 (N_11612,N_11362,N_11238);
nor U11613 (N_11613,N_11125,N_11230);
xor U11614 (N_11614,N_11410,N_11489);
nand U11615 (N_11615,N_11032,N_11379);
or U11616 (N_11616,N_11300,N_11201);
nor U11617 (N_11617,N_11241,N_11378);
or U11618 (N_11618,N_11285,N_11198);
nor U11619 (N_11619,N_11005,N_11367);
or U11620 (N_11620,N_11445,N_11023);
and U11621 (N_11621,N_11250,N_11425);
xnor U11622 (N_11622,N_11248,N_11385);
nand U11623 (N_11623,N_11334,N_11464);
xor U11624 (N_11624,N_11290,N_11106);
and U11625 (N_11625,N_11479,N_11431);
nor U11626 (N_11626,N_11320,N_11336);
and U11627 (N_11627,N_11002,N_11392);
nor U11628 (N_11628,N_11451,N_11364);
and U11629 (N_11629,N_11075,N_11035);
and U11630 (N_11630,N_11029,N_11115);
nand U11631 (N_11631,N_11447,N_11301);
or U11632 (N_11632,N_11446,N_11212);
xor U11633 (N_11633,N_11221,N_11494);
nand U11634 (N_11634,N_11169,N_11480);
nand U11635 (N_11635,N_11396,N_11329);
or U11636 (N_11636,N_11213,N_11206);
or U11637 (N_11637,N_11007,N_11407);
nor U11638 (N_11638,N_11306,N_11340);
xnor U11639 (N_11639,N_11012,N_11134);
nand U11640 (N_11640,N_11498,N_11255);
nand U11641 (N_11641,N_11048,N_11054);
and U11642 (N_11642,N_11152,N_11132);
or U11643 (N_11643,N_11203,N_11455);
nand U11644 (N_11644,N_11172,N_11017);
and U11645 (N_11645,N_11352,N_11160);
nand U11646 (N_11646,N_11159,N_11229);
nand U11647 (N_11647,N_11195,N_11189);
xor U11648 (N_11648,N_11440,N_11124);
xnor U11649 (N_11649,N_11165,N_11467);
nor U11650 (N_11650,N_11237,N_11408);
or U11651 (N_11651,N_11486,N_11216);
xor U11652 (N_11652,N_11343,N_11135);
nand U11653 (N_11653,N_11449,N_11495);
and U11654 (N_11654,N_11273,N_11289);
or U11655 (N_11655,N_11388,N_11001);
nand U11656 (N_11656,N_11316,N_11271);
xor U11657 (N_11657,N_11399,N_11108);
nor U11658 (N_11658,N_11481,N_11265);
nand U11659 (N_11659,N_11390,N_11482);
and U11660 (N_11660,N_11463,N_11240);
or U11661 (N_11661,N_11133,N_11279);
and U11662 (N_11662,N_11197,N_11140);
and U11663 (N_11663,N_11375,N_11309);
nor U11664 (N_11664,N_11121,N_11069);
nand U11665 (N_11665,N_11131,N_11110);
or U11666 (N_11666,N_11139,N_11156);
nand U11667 (N_11667,N_11471,N_11036);
nor U11668 (N_11668,N_11267,N_11066);
xor U11669 (N_11669,N_11278,N_11065);
and U11670 (N_11670,N_11288,N_11185);
and U11671 (N_11671,N_11044,N_11246);
and U11672 (N_11672,N_11281,N_11059);
or U11673 (N_11673,N_11041,N_11039);
xor U11674 (N_11674,N_11380,N_11010);
and U11675 (N_11675,N_11129,N_11296);
nand U11676 (N_11676,N_11031,N_11101);
nand U11677 (N_11677,N_11465,N_11413);
nand U11678 (N_11678,N_11297,N_11167);
and U11679 (N_11679,N_11470,N_11459);
or U11680 (N_11680,N_11412,N_11128);
nor U11681 (N_11681,N_11304,N_11109);
nor U11682 (N_11682,N_11179,N_11469);
or U11683 (N_11683,N_11068,N_11155);
nor U11684 (N_11684,N_11411,N_11090);
nor U11685 (N_11685,N_11438,N_11272);
xor U11686 (N_11686,N_11158,N_11107);
or U11687 (N_11687,N_11123,N_11046);
or U11688 (N_11688,N_11102,N_11363);
nor U11689 (N_11689,N_11114,N_11491);
or U11690 (N_11690,N_11092,N_11067);
nand U11691 (N_11691,N_11346,N_11164);
nor U11692 (N_11692,N_11119,N_11427);
or U11693 (N_11693,N_11295,N_11209);
nor U11694 (N_11694,N_11026,N_11418);
or U11695 (N_11695,N_11433,N_11315);
nor U11696 (N_11696,N_11177,N_11064);
or U11697 (N_11697,N_11116,N_11299);
xnor U11698 (N_11698,N_11171,N_11040);
xnor U11699 (N_11699,N_11450,N_11391);
or U11700 (N_11700,N_11024,N_11368);
nor U11701 (N_11701,N_11180,N_11337);
nor U11702 (N_11702,N_11223,N_11422);
xnor U11703 (N_11703,N_11483,N_11404);
or U11704 (N_11704,N_11478,N_11298);
xor U11705 (N_11705,N_11210,N_11499);
xnor U11706 (N_11706,N_11373,N_11387);
or U11707 (N_11707,N_11349,N_11327);
nand U11708 (N_11708,N_11013,N_11432);
nor U11709 (N_11709,N_11347,N_11401);
and U11710 (N_11710,N_11428,N_11168);
and U11711 (N_11711,N_11018,N_11252);
and U11712 (N_11712,N_11153,N_11057);
and U11713 (N_11713,N_11382,N_11043);
xor U11714 (N_11714,N_11454,N_11264);
nand U11715 (N_11715,N_11318,N_11308);
nor U11716 (N_11716,N_11270,N_11263);
or U11717 (N_11717,N_11219,N_11207);
nand U11718 (N_11718,N_11015,N_11188);
and U11719 (N_11719,N_11021,N_11280);
xnor U11720 (N_11720,N_11224,N_11326);
nand U11721 (N_11721,N_11358,N_11457);
or U11722 (N_11722,N_11202,N_11442);
or U11723 (N_11723,N_11215,N_11211);
xor U11724 (N_11724,N_11389,N_11226);
or U11725 (N_11725,N_11453,N_11190);
xor U11726 (N_11726,N_11261,N_11441);
xor U11727 (N_11727,N_11042,N_11312);
nand U11728 (N_11728,N_11247,N_11284);
or U11729 (N_11729,N_11475,N_11472);
nand U11730 (N_11730,N_11150,N_11163);
nand U11731 (N_11731,N_11118,N_11176);
nand U11732 (N_11732,N_11360,N_11324);
xnor U11733 (N_11733,N_11022,N_11361);
xor U11734 (N_11734,N_11342,N_11220);
nand U11735 (N_11735,N_11087,N_11182);
nand U11736 (N_11736,N_11187,N_11420);
xnor U11737 (N_11737,N_11127,N_11183);
xnor U11738 (N_11738,N_11405,N_11466);
xnor U11739 (N_11739,N_11417,N_11025);
and U11740 (N_11740,N_11073,N_11014);
or U11741 (N_11741,N_11061,N_11060);
or U11742 (N_11742,N_11218,N_11099);
nand U11743 (N_11743,N_11416,N_11053);
xor U11744 (N_11744,N_11292,N_11251);
and U11745 (N_11745,N_11477,N_11100);
xnor U11746 (N_11746,N_11492,N_11394);
nor U11747 (N_11747,N_11397,N_11070);
or U11748 (N_11748,N_11145,N_11081);
or U11749 (N_11749,N_11082,N_11074);
and U11750 (N_11750,N_11384,N_11071);
nand U11751 (N_11751,N_11124,N_11096);
xnor U11752 (N_11752,N_11356,N_11052);
nor U11753 (N_11753,N_11177,N_11324);
xor U11754 (N_11754,N_11382,N_11141);
nor U11755 (N_11755,N_11317,N_11460);
nor U11756 (N_11756,N_11295,N_11387);
nand U11757 (N_11757,N_11260,N_11286);
or U11758 (N_11758,N_11238,N_11432);
nor U11759 (N_11759,N_11099,N_11184);
or U11760 (N_11760,N_11015,N_11496);
nand U11761 (N_11761,N_11481,N_11057);
and U11762 (N_11762,N_11216,N_11002);
nand U11763 (N_11763,N_11004,N_11365);
nand U11764 (N_11764,N_11454,N_11154);
or U11765 (N_11765,N_11479,N_11271);
xnor U11766 (N_11766,N_11415,N_11477);
nand U11767 (N_11767,N_11375,N_11212);
xnor U11768 (N_11768,N_11130,N_11065);
xnor U11769 (N_11769,N_11052,N_11148);
or U11770 (N_11770,N_11195,N_11199);
and U11771 (N_11771,N_11320,N_11441);
xnor U11772 (N_11772,N_11121,N_11198);
xor U11773 (N_11773,N_11156,N_11476);
and U11774 (N_11774,N_11165,N_11186);
nor U11775 (N_11775,N_11180,N_11062);
xnor U11776 (N_11776,N_11023,N_11345);
xor U11777 (N_11777,N_11367,N_11378);
xor U11778 (N_11778,N_11248,N_11170);
nand U11779 (N_11779,N_11388,N_11062);
xor U11780 (N_11780,N_11485,N_11273);
xor U11781 (N_11781,N_11238,N_11195);
xnor U11782 (N_11782,N_11170,N_11395);
nand U11783 (N_11783,N_11004,N_11001);
nand U11784 (N_11784,N_11095,N_11052);
xnor U11785 (N_11785,N_11254,N_11203);
xnor U11786 (N_11786,N_11358,N_11388);
nor U11787 (N_11787,N_11297,N_11023);
nor U11788 (N_11788,N_11444,N_11152);
xor U11789 (N_11789,N_11383,N_11277);
xnor U11790 (N_11790,N_11201,N_11165);
nor U11791 (N_11791,N_11109,N_11250);
and U11792 (N_11792,N_11013,N_11382);
nor U11793 (N_11793,N_11096,N_11070);
nor U11794 (N_11794,N_11053,N_11078);
nor U11795 (N_11795,N_11189,N_11006);
and U11796 (N_11796,N_11076,N_11062);
xor U11797 (N_11797,N_11474,N_11277);
nor U11798 (N_11798,N_11427,N_11294);
nor U11799 (N_11799,N_11259,N_11178);
or U11800 (N_11800,N_11050,N_11222);
xnor U11801 (N_11801,N_11032,N_11123);
nor U11802 (N_11802,N_11167,N_11108);
nor U11803 (N_11803,N_11148,N_11096);
and U11804 (N_11804,N_11410,N_11289);
xnor U11805 (N_11805,N_11270,N_11058);
xnor U11806 (N_11806,N_11180,N_11055);
xnor U11807 (N_11807,N_11213,N_11184);
or U11808 (N_11808,N_11217,N_11462);
nor U11809 (N_11809,N_11220,N_11063);
or U11810 (N_11810,N_11178,N_11377);
nand U11811 (N_11811,N_11306,N_11369);
nor U11812 (N_11812,N_11405,N_11430);
xnor U11813 (N_11813,N_11041,N_11030);
xor U11814 (N_11814,N_11063,N_11382);
and U11815 (N_11815,N_11239,N_11182);
and U11816 (N_11816,N_11072,N_11149);
nor U11817 (N_11817,N_11242,N_11006);
nor U11818 (N_11818,N_11065,N_11066);
or U11819 (N_11819,N_11484,N_11121);
xor U11820 (N_11820,N_11461,N_11077);
or U11821 (N_11821,N_11408,N_11045);
nor U11822 (N_11822,N_11372,N_11053);
or U11823 (N_11823,N_11104,N_11477);
and U11824 (N_11824,N_11037,N_11445);
xnor U11825 (N_11825,N_11187,N_11110);
and U11826 (N_11826,N_11340,N_11279);
and U11827 (N_11827,N_11201,N_11215);
xnor U11828 (N_11828,N_11407,N_11390);
nor U11829 (N_11829,N_11133,N_11499);
xnor U11830 (N_11830,N_11176,N_11013);
or U11831 (N_11831,N_11199,N_11249);
and U11832 (N_11832,N_11338,N_11432);
xnor U11833 (N_11833,N_11062,N_11256);
or U11834 (N_11834,N_11425,N_11237);
xor U11835 (N_11835,N_11395,N_11129);
or U11836 (N_11836,N_11323,N_11061);
and U11837 (N_11837,N_11465,N_11018);
xor U11838 (N_11838,N_11001,N_11035);
xor U11839 (N_11839,N_11148,N_11330);
nor U11840 (N_11840,N_11096,N_11291);
nor U11841 (N_11841,N_11112,N_11264);
xor U11842 (N_11842,N_11319,N_11062);
xor U11843 (N_11843,N_11462,N_11417);
nor U11844 (N_11844,N_11149,N_11322);
nor U11845 (N_11845,N_11051,N_11042);
nand U11846 (N_11846,N_11155,N_11231);
or U11847 (N_11847,N_11113,N_11325);
or U11848 (N_11848,N_11329,N_11467);
and U11849 (N_11849,N_11454,N_11435);
nor U11850 (N_11850,N_11274,N_11473);
or U11851 (N_11851,N_11379,N_11399);
and U11852 (N_11852,N_11280,N_11108);
or U11853 (N_11853,N_11131,N_11064);
nor U11854 (N_11854,N_11106,N_11034);
nor U11855 (N_11855,N_11303,N_11036);
and U11856 (N_11856,N_11344,N_11100);
nand U11857 (N_11857,N_11416,N_11303);
xor U11858 (N_11858,N_11480,N_11300);
and U11859 (N_11859,N_11370,N_11015);
and U11860 (N_11860,N_11016,N_11136);
nor U11861 (N_11861,N_11477,N_11494);
or U11862 (N_11862,N_11470,N_11332);
nand U11863 (N_11863,N_11436,N_11416);
nand U11864 (N_11864,N_11454,N_11378);
and U11865 (N_11865,N_11323,N_11438);
or U11866 (N_11866,N_11037,N_11219);
nor U11867 (N_11867,N_11376,N_11193);
or U11868 (N_11868,N_11106,N_11043);
or U11869 (N_11869,N_11350,N_11034);
and U11870 (N_11870,N_11039,N_11171);
or U11871 (N_11871,N_11369,N_11102);
and U11872 (N_11872,N_11364,N_11479);
nor U11873 (N_11873,N_11088,N_11390);
and U11874 (N_11874,N_11217,N_11271);
xnor U11875 (N_11875,N_11206,N_11268);
nand U11876 (N_11876,N_11194,N_11035);
or U11877 (N_11877,N_11208,N_11106);
nand U11878 (N_11878,N_11016,N_11265);
nand U11879 (N_11879,N_11452,N_11047);
nor U11880 (N_11880,N_11066,N_11190);
or U11881 (N_11881,N_11428,N_11205);
or U11882 (N_11882,N_11437,N_11204);
nor U11883 (N_11883,N_11379,N_11075);
nand U11884 (N_11884,N_11370,N_11087);
nand U11885 (N_11885,N_11399,N_11294);
or U11886 (N_11886,N_11191,N_11206);
xnor U11887 (N_11887,N_11377,N_11061);
or U11888 (N_11888,N_11290,N_11181);
nand U11889 (N_11889,N_11191,N_11212);
xor U11890 (N_11890,N_11425,N_11012);
nand U11891 (N_11891,N_11046,N_11425);
nand U11892 (N_11892,N_11338,N_11347);
or U11893 (N_11893,N_11388,N_11137);
and U11894 (N_11894,N_11300,N_11347);
nand U11895 (N_11895,N_11454,N_11415);
xor U11896 (N_11896,N_11058,N_11489);
and U11897 (N_11897,N_11067,N_11158);
or U11898 (N_11898,N_11174,N_11197);
or U11899 (N_11899,N_11134,N_11023);
xor U11900 (N_11900,N_11424,N_11418);
nand U11901 (N_11901,N_11224,N_11199);
nand U11902 (N_11902,N_11277,N_11319);
nand U11903 (N_11903,N_11412,N_11318);
nand U11904 (N_11904,N_11478,N_11214);
nand U11905 (N_11905,N_11248,N_11132);
nand U11906 (N_11906,N_11098,N_11463);
and U11907 (N_11907,N_11448,N_11274);
nand U11908 (N_11908,N_11185,N_11126);
nor U11909 (N_11909,N_11327,N_11023);
and U11910 (N_11910,N_11416,N_11317);
nor U11911 (N_11911,N_11300,N_11365);
xnor U11912 (N_11912,N_11423,N_11124);
or U11913 (N_11913,N_11256,N_11309);
nand U11914 (N_11914,N_11292,N_11326);
or U11915 (N_11915,N_11250,N_11031);
nor U11916 (N_11916,N_11269,N_11471);
xor U11917 (N_11917,N_11269,N_11403);
nand U11918 (N_11918,N_11415,N_11115);
nand U11919 (N_11919,N_11122,N_11412);
xor U11920 (N_11920,N_11188,N_11085);
or U11921 (N_11921,N_11146,N_11410);
and U11922 (N_11922,N_11172,N_11101);
and U11923 (N_11923,N_11337,N_11338);
or U11924 (N_11924,N_11344,N_11369);
and U11925 (N_11925,N_11113,N_11085);
nand U11926 (N_11926,N_11461,N_11216);
or U11927 (N_11927,N_11188,N_11481);
or U11928 (N_11928,N_11332,N_11258);
and U11929 (N_11929,N_11313,N_11076);
nor U11930 (N_11930,N_11443,N_11314);
nand U11931 (N_11931,N_11407,N_11362);
nor U11932 (N_11932,N_11044,N_11168);
nand U11933 (N_11933,N_11287,N_11218);
and U11934 (N_11934,N_11002,N_11107);
or U11935 (N_11935,N_11044,N_11438);
nand U11936 (N_11936,N_11390,N_11098);
xnor U11937 (N_11937,N_11205,N_11149);
nor U11938 (N_11938,N_11143,N_11476);
or U11939 (N_11939,N_11014,N_11445);
nor U11940 (N_11940,N_11425,N_11117);
or U11941 (N_11941,N_11027,N_11292);
xor U11942 (N_11942,N_11374,N_11238);
and U11943 (N_11943,N_11348,N_11375);
nor U11944 (N_11944,N_11454,N_11078);
and U11945 (N_11945,N_11468,N_11198);
nor U11946 (N_11946,N_11265,N_11449);
xor U11947 (N_11947,N_11422,N_11257);
nand U11948 (N_11948,N_11267,N_11373);
xor U11949 (N_11949,N_11375,N_11111);
nand U11950 (N_11950,N_11101,N_11486);
nor U11951 (N_11951,N_11303,N_11329);
xnor U11952 (N_11952,N_11382,N_11131);
nand U11953 (N_11953,N_11375,N_11264);
or U11954 (N_11954,N_11013,N_11001);
nor U11955 (N_11955,N_11282,N_11434);
and U11956 (N_11956,N_11026,N_11376);
and U11957 (N_11957,N_11165,N_11360);
and U11958 (N_11958,N_11053,N_11499);
or U11959 (N_11959,N_11338,N_11433);
or U11960 (N_11960,N_11480,N_11389);
or U11961 (N_11961,N_11130,N_11323);
nand U11962 (N_11962,N_11317,N_11313);
nand U11963 (N_11963,N_11277,N_11184);
and U11964 (N_11964,N_11197,N_11004);
xor U11965 (N_11965,N_11162,N_11326);
xnor U11966 (N_11966,N_11054,N_11293);
nand U11967 (N_11967,N_11169,N_11103);
or U11968 (N_11968,N_11013,N_11261);
xor U11969 (N_11969,N_11390,N_11130);
nand U11970 (N_11970,N_11199,N_11013);
nand U11971 (N_11971,N_11181,N_11058);
nor U11972 (N_11972,N_11286,N_11084);
or U11973 (N_11973,N_11429,N_11040);
xnor U11974 (N_11974,N_11289,N_11165);
nor U11975 (N_11975,N_11474,N_11479);
xnor U11976 (N_11976,N_11407,N_11013);
xor U11977 (N_11977,N_11483,N_11395);
or U11978 (N_11978,N_11109,N_11286);
xnor U11979 (N_11979,N_11267,N_11172);
or U11980 (N_11980,N_11406,N_11117);
and U11981 (N_11981,N_11358,N_11027);
xor U11982 (N_11982,N_11498,N_11311);
nor U11983 (N_11983,N_11348,N_11493);
and U11984 (N_11984,N_11335,N_11194);
nor U11985 (N_11985,N_11451,N_11499);
xnor U11986 (N_11986,N_11104,N_11098);
or U11987 (N_11987,N_11246,N_11465);
xor U11988 (N_11988,N_11100,N_11197);
nand U11989 (N_11989,N_11066,N_11313);
nor U11990 (N_11990,N_11374,N_11472);
xor U11991 (N_11991,N_11048,N_11265);
and U11992 (N_11992,N_11236,N_11229);
nor U11993 (N_11993,N_11492,N_11146);
and U11994 (N_11994,N_11215,N_11179);
or U11995 (N_11995,N_11005,N_11112);
or U11996 (N_11996,N_11300,N_11293);
nand U11997 (N_11997,N_11129,N_11278);
or U11998 (N_11998,N_11497,N_11193);
or U11999 (N_11999,N_11463,N_11310);
or U12000 (N_12000,N_11891,N_11691);
xor U12001 (N_12001,N_11780,N_11841);
or U12002 (N_12002,N_11956,N_11705);
nor U12003 (N_12003,N_11865,N_11829);
nand U12004 (N_12004,N_11781,N_11807);
nor U12005 (N_12005,N_11557,N_11798);
xor U12006 (N_12006,N_11912,N_11657);
xnor U12007 (N_12007,N_11839,N_11972);
xor U12008 (N_12008,N_11523,N_11538);
nor U12009 (N_12009,N_11675,N_11717);
nor U12010 (N_12010,N_11643,N_11968);
or U12011 (N_12011,N_11812,N_11710);
and U12012 (N_12012,N_11613,N_11656);
and U12013 (N_12013,N_11728,N_11535);
or U12014 (N_12014,N_11754,N_11867);
nor U12015 (N_12015,N_11712,N_11616);
or U12016 (N_12016,N_11633,N_11795);
and U12017 (N_12017,N_11810,N_11857);
and U12018 (N_12018,N_11703,N_11879);
xor U12019 (N_12019,N_11859,N_11826);
nand U12020 (N_12020,N_11825,N_11687);
and U12021 (N_12021,N_11597,N_11636);
or U12022 (N_12022,N_11836,N_11734);
or U12023 (N_12023,N_11869,N_11991);
nor U12024 (N_12024,N_11609,N_11843);
or U12025 (N_12025,N_11581,N_11670);
xnor U12026 (N_12026,N_11804,N_11603);
or U12027 (N_12027,N_11593,N_11901);
xor U12028 (N_12028,N_11700,N_11676);
or U12029 (N_12029,N_11686,N_11773);
or U12030 (N_12030,N_11929,N_11583);
and U12031 (N_12031,N_11787,N_11904);
nand U12032 (N_12032,N_11548,N_11562);
xnor U12033 (N_12033,N_11560,N_11961);
or U12034 (N_12034,N_11527,N_11702);
or U12035 (N_12035,N_11601,N_11666);
or U12036 (N_12036,N_11847,N_11600);
nor U12037 (N_12037,N_11720,N_11753);
and U12038 (N_12038,N_11989,N_11940);
or U12039 (N_12039,N_11598,N_11910);
nand U12040 (N_12040,N_11987,N_11574);
and U12041 (N_12041,N_11817,N_11532);
or U12042 (N_12042,N_11797,N_11762);
and U12043 (N_12043,N_11694,N_11564);
nor U12044 (N_12044,N_11567,N_11701);
and U12045 (N_12045,N_11944,N_11775);
nor U12046 (N_12046,N_11552,N_11800);
nand U12047 (N_12047,N_11665,N_11755);
or U12048 (N_12048,N_11861,N_11791);
nand U12049 (N_12049,N_11974,N_11536);
nand U12050 (N_12050,N_11856,N_11945);
and U12051 (N_12051,N_11632,N_11623);
nor U12052 (N_12052,N_11683,N_11556);
and U12053 (N_12053,N_11794,N_11913);
nand U12054 (N_12054,N_11577,N_11559);
nor U12055 (N_12055,N_11948,N_11640);
and U12056 (N_12056,N_11652,N_11501);
nand U12057 (N_12057,N_11772,N_11846);
nand U12058 (N_12058,N_11522,N_11838);
nor U12059 (N_12059,N_11752,N_11881);
nor U12060 (N_12060,N_11938,N_11892);
nor U12061 (N_12061,N_11530,N_11515);
nand U12062 (N_12062,N_11539,N_11934);
or U12063 (N_12063,N_11953,N_11635);
xnor U12064 (N_12064,N_11801,N_11506);
or U12065 (N_12065,N_11872,N_11950);
and U12066 (N_12066,N_11648,N_11627);
or U12067 (N_12067,N_11820,N_11840);
or U12068 (N_12068,N_11588,N_11570);
nor U12069 (N_12069,N_11928,N_11844);
and U12070 (N_12070,N_11771,N_11650);
or U12071 (N_12071,N_11965,N_11511);
or U12072 (N_12072,N_11898,N_11606);
nor U12073 (N_12073,N_11995,N_11799);
nor U12074 (N_12074,N_11905,N_11960);
nor U12075 (N_12075,N_11866,N_11526);
xor U12076 (N_12076,N_11713,N_11599);
xor U12077 (N_12077,N_11774,N_11823);
or U12078 (N_12078,N_11568,N_11977);
and U12079 (N_12079,N_11628,N_11980);
xor U12080 (N_12080,N_11500,N_11963);
or U12081 (N_12081,N_11925,N_11604);
nor U12082 (N_12082,N_11900,N_11602);
or U12083 (N_12083,N_11765,N_11620);
and U12084 (N_12084,N_11646,N_11607);
nor U12085 (N_12085,N_11890,N_11739);
xnor U12086 (N_12086,N_11626,N_11575);
and U12087 (N_12087,N_11951,N_11757);
nand U12088 (N_12088,N_11582,N_11924);
nor U12089 (N_12089,N_11727,N_11885);
nor U12090 (N_12090,N_11550,N_11692);
and U12091 (N_12091,N_11964,N_11661);
xnor U12092 (N_12092,N_11664,N_11874);
nor U12093 (N_12093,N_11814,N_11729);
nand U12094 (N_12094,N_11918,N_11811);
and U12095 (N_12095,N_11561,N_11507);
or U12096 (N_12096,N_11743,N_11681);
nor U12097 (N_12097,N_11596,N_11707);
or U12098 (N_12098,N_11615,N_11962);
nand U12099 (N_12099,N_11726,N_11576);
nand U12100 (N_12100,N_11992,N_11519);
or U12101 (N_12101,N_11883,N_11782);
and U12102 (N_12102,N_11572,N_11592);
nor U12103 (N_12103,N_11863,N_11818);
or U12104 (N_12104,N_11653,N_11723);
or U12105 (N_12105,N_11858,N_11809);
or U12106 (N_12106,N_11966,N_11554);
nand U12107 (N_12107,N_11513,N_11789);
nor U12108 (N_12108,N_11860,N_11880);
xor U12109 (N_12109,N_11978,N_11751);
nand U12110 (N_12110,N_11837,N_11591);
and U12111 (N_12111,N_11544,N_11645);
and U12112 (N_12112,N_11864,N_11677);
xnor U12113 (N_12113,N_11954,N_11595);
or U12114 (N_12114,N_11721,N_11736);
or U12115 (N_12115,N_11622,N_11630);
or U12116 (N_12116,N_11541,N_11853);
nand U12117 (N_12117,N_11673,N_11612);
nor U12118 (N_12118,N_11589,N_11709);
nand U12119 (N_12119,N_11540,N_11788);
and U12120 (N_12120,N_11927,N_11660);
or U12121 (N_12121,N_11768,N_11767);
nand U12122 (N_12122,N_11505,N_11842);
nand U12123 (N_12123,N_11999,N_11618);
or U12124 (N_12124,N_11899,N_11914);
and U12125 (N_12125,N_11770,N_11947);
xnor U12126 (N_12126,N_11931,N_11619);
and U12127 (N_12127,N_11587,N_11525);
nor U12128 (N_12128,N_11868,N_11921);
xnor U12129 (N_12129,N_11850,N_11672);
nand U12130 (N_12130,N_11573,N_11735);
nand U12131 (N_12131,N_11737,N_11512);
xnor U12132 (N_12132,N_11920,N_11827);
nand U12133 (N_12133,N_11537,N_11534);
nand U12134 (N_12134,N_11509,N_11808);
nor U12135 (N_12135,N_11908,N_11689);
and U12136 (N_12136,N_11680,N_11786);
and U12137 (N_12137,N_11877,N_11549);
xnor U12138 (N_12138,N_11870,N_11916);
nor U12139 (N_12139,N_11822,N_11806);
xnor U12140 (N_12140,N_11888,N_11696);
or U12141 (N_12141,N_11551,N_11990);
nand U12142 (N_12142,N_11835,N_11919);
xnor U12143 (N_12143,N_11516,N_11684);
nor U12144 (N_12144,N_11738,N_11655);
nand U12145 (N_12145,N_11979,N_11503);
xor U12146 (N_12146,N_11886,N_11502);
or U12147 (N_12147,N_11876,N_11805);
and U12148 (N_12148,N_11518,N_11543);
nor U12149 (N_12149,N_11862,N_11558);
or U12150 (N_12150,N_11796,N_11637);
nor U12151 (N_12151,N_11894,N_11639);
nor U12152 (N_12152,N_11975,N_11504);
nor U12153 (N_12153,N_11642,N_11741);
or U12154 (N_12154,N_11941,N_11629);
nand U12155 (N_12155,N_11832,N_11802);
nor U12156 (N_12156,N_11679,N_11730);
or U12157 (N_12157,N_11624,N_11658);
or U12158 (N_12158,N_11764,N_11893);
nand U12159 (N_12159,N_11942,N_11760);
and U12160 (N_12160,N_11834,N_11959);
xor U12161 (N_12161,N_11663,N_11711);
nand U12162 (N_12162,N_11614,N_11563);
xor U12163 (N_12163,N_11889,N_11824);
nand U12164 (N_12164,N_11569,N_11545);
xor U12165 (N_12165,N_11958,N_11813);
nand U12166 (N_12166,N_11937,N_11976);
or U12167 (N_12167,N_11785,N_11546);
nand U12168 (N_12168,N_11533,N_11725);
nand U12169 (N_12169,N_11933,N_11678);
nor U12170 (N_12170,N_11625,N_11565);
nand U12171 (N_12171,N_11731,N_11580);
and U12172 (N_12172,N_11510,N_11952);
nor U12173 (N_12173,N_11708,N_11685);
or U12174 (N_12174,N_11668,N_11514);
xor U12175 (N_12175,N_11578,N_11936);
and U12176 (N_12176,N_11698,N_11855);
xnor U12177 (N_12177,N_11585,N_11766);
nand U12178 (N_12178,N_11555,N_11831);
nor U12179 (N_12179,N_11553,N_11981);
or U12180 (N_12180,N_11902,N_11695);
or U12181 (N_12181,N_11520,N_11949);
nand U12182 (N_12182,N_11884,N_11641);
or U12183 (N_12183,N_11793,N_11719);
and U12184 (N_12184,N_11943,N_11667);
or U12185 (N_12185,N_11631,N_11848);
or U12186 (N_12186,N_11756,N_11605);
and U12187 (N_12187,N_11815,N_11531);
nand U12188 (N_12188,N_11651,N_11547);
or U12189 (N_12189,N_11654,N_11878);
nand U12190 (N_12190,N_11758,N_11983);
nand U12191 (N_12191,N_11988,N_11955);
nand U12192 (N_12192,N_11833,N_11996);
nor U12193 (N_12193,N_11821,N_11871);
or U12194 (N_12194,N_11907,N_11986);
nand U12195 (N_12195,N_11887,N_11749);
and U12196 (N_12196,N_11994,N_11524);
nand U12197 (N_12197,N_11790,N_11896);
and U12198 (N_12198,N_11644,N_11993);
xnor U12199 (N_12199,N_11732,N_11769);
nand U12200 (N_12200,N_11517,N_11688);
or U12201 (N_12201,N_11682,N_11971);
nand U12202 (N_12202,N_11716,N_11845);
nor U12203 (N_12203,N_11747,N_11939);
nand U12204 (N_12204,N_11828,N_11935);
and U12205 (N_12205,N_11528,N_11669);
xor U12206 (N_12206,N_11699,N_11763);
nand U12207 (N_12207,N_11610,N_11917);
nor U12208 (N_12208,N_11715,N_11903);
nor U12209 (N_12209,N_11674,N_11508);
or U12210 (N_12210,N_11816,N_11590);
and U12211 (N_12211,N_11617,N_11759);
xor U12212 (N_12212,N_11932,N_11671);
or U12213 (N_12213,N_11748,N_11895);
or U12214 (N_12214,N_11690,N_11579);
and U12215 (N_12215,N_11985,N_11875);
or U12216 (N_12216,N_11529,N_11973);
and U12217 (N_12217,N_11566,N_11697);
or U12218 (N_12218,N_11778,N_11718);
nor U12219 (N_12219,N_11706,N_11922);
and U12220 (N_12220,N_11571,N_11744);
nand U12221 (N_12221,N_11957,N_11647);
and U12222 (N_12222,N_11634,N_11882);
or U12223 (N_12223,N_11909,N_11819);
nand U12224 (N_12224,N_11792,N_11930);
nor U12225 (N_12225,N_11873,N_11946);
xnor U12226 (N_12226,N_11594,N_11969);
nand U12227 (N_12227,N_11722,N_11733);
or U12228 (N_12228,N_11746,N_11659);
or U12229 (N_12229,N_11621,N_11750);
nor U12230 (N_12230,N_11982,N_11608);
xor U12231 (N_12231,N_11693,N_11662);
and U12232 (N_12232,N_11830,N_11586);
or U12233 (N_12233,N_11854,N_11997);
xor U12234 (N_12234,N_11915,N_11776);
xnor U12235 (N_12235,N_11638,N_11852);
nand U12236 (N_12236,N_11911,N_11851);
nand U12237 (N_12237,N_11906,N_11745);
and U12238 (N_12238,N_11724,N_11779);
or U12239 (N_12239,N_11611,N_11542);
nor U12240 (N_12240,N_11923,N_11783);
or U12241 (N_12241,N_11967,N_11521);
nand U12242 (N_12242,N_11784,N_11649);
nand U12243 (N_12243,N_11998,N_11803);
nand U12244 (N_12244,N_11984,N_11926);
and U12245 (N_12245,N_11761,N_11849);
or U12246 (N_12246,N_11970,N_11777);
nor U12247 (N_12247,N_11704,N_11584);
nand U12248 (N_12248,N_11714,N_11897);
or U12249 (N_12249,N_11740,N_11742);
and U12250 (N_12250,N_11618,N_11505);
or U12251 (N_12251,N_11888,N_11803);
nand U12252 (N_12252,N_11976,N_11785);
xor U12253 (N_12253,N_11666,N_11787);
or U12254 (N_12254,N_11828,N_11677);
xor U12255 (N_12255,N_11722,N_11954);
nor U12256 (N_12256,N_11768,N_11819);
xor U12257 (N_12257,N_11903,N_11723);
nor U12258 (N_12258,N_11899,N_11910);
xor U12259 (N_12259,N_11864,N_11621);
nor U12260 (N_12260,N_11752,N_11674);
xor U12261 (N_12261,N_11930,N_11559);
and U12262 (N_12262,N_11808,N_11799);
and U12263 (N_12263,N_11662,N_11990);
nand U12264 (N_12264,N_11916,N_11766);
and U12265 (N_12265,N_11914,N_11924);
or U12266 (N_12266,N_11756,N_11617);
nand U12267 (N_12267,N_11522,N_11853);
nor U12268 (N_12268,N_11508,N_11592);
or U12269 (N_12269,N_11506,N_11511);
nor U12270 (N_12270,N_11736,N_11550);
or U12271 (N_12271,N_11662,N_11863);
or U12272 (N_12272,N_11540,N_11918);
nand U12273 (N_12273,N_11945,N_11659);
or U12274 (N_12274,N_11588,N_11876);
nor U12275 (N_12275,N_11974,N_11956);
nor U12276 (N_12276,N_11762,N_11546);
nor U12277 (N_12277,N_11993,N_11879);
nor U12278 (N_12278,N_11829,N_11981);
nand U12279 (N_12279,N_11788,N_11585);
and U12280 (N_12280,N_11920,N_11669);
or U12281 (N_12281,N_11702,N_11863);
or U12282 (N_12282,N_11780,N_11741);
xor U12283 (N_12283,N_11630,N_11852);
nand U12284 (N_12284,N_11590,N_11689);
nor U12285 (N_12285,N_11885,N_11711);
or U12286 (N_12286,N_11978,N_11825);
nand U12287 (N_12287,N_11575,N_11910);
nand U12288 (N_12288,N_11745,N_11964);
and U12289 (N_12289,N_11709,N_11613);
xor U12290 (N_12290,N_11969,N_11995);
nand U12291 (N_12291,N_11747,N_11706);
nand U12292 (N_12292,N_11895,N_11838);
or U12293 (N_12293,N_11628,N_11881);
nor U12294 (N_12294,N_11644,N_11788);
nand U12295 (N_12295,N_11813,N_11718);
nand U12296 (N_12296,N_11615,N_11537);
nand U12297 (N_12297,N_11886,N_11724);
nand U12298 (N_12298,N_11767,N_11709);
and U12299 (N_12299,N_11656,N_11524);
nand U12300 (N_12300,N_11618,N_11566);
xor U12301 (N_12301,N_11589,N_11547);
nand U12302 (N_12302,N_11697,N_11935);
nor U12303 (N_12303,N_11717,N_11514);
nor U12304 (N_12304,N_11620,N_11885);
nand U12305 (N_12305,N_11569,N_11998);
nand U12306 (N_12306,N_11975,N_11564);
xnor U12307 (N_12307,N_11859,N_11593);
xor U12308 (N_12308,N_11720,N_11654);
or U12309 (N_12309,N_11595,N_11836);
or U12310 (N_12310,N_11777,N_11742);
xor U12311 (N_12311,N_11924,N_11741);
nand U12312 (N_12312,N_11896,N_11568);
and U12313 (N_12313,N_11691,N_11930);
xnor U12314 (N_12314,N_11962,N_11584);
nor U12315 (N_12315,N_11999,N_11976);
or U12316 (N_12316,N_11669,N_11981);
and U12317 (N_12317,N_11873,N_11867);
or U12318 (N_12318,N_11985,N_11610);
nand U12319 (N_12319,N_11988,N_11942);
nand U12320 (N_12320,N_11894,N_11775);
nand U12321 (N_12321,N_11626,N_11589);
xor U12322 (N_12322,N_11765,N_11979);
nand U12323 (N_12323,N_11770,N_11821);
nand U12324 (N_12324,N_11808,N_11652);
or U12325 (N_12325,N_11798,N_11962);
nor U12326 (N_12326,N_11590,N_11942);
or U12327 (N_12327,N_11794,N_11781);
nand U12328 (N_12328,N_11519,N_11617);
nand U12329 (N_12329,N_11971,N_11901);
and U12330 (N_12330,N_11589,N_11787);
and U12331 (N_12331,N_11615,N_11743);
or U12332 (N_12332,N_11812,N_11589);
or U12333 (N_12333,N_11581,N_11920);
or U12334 (N_12334,N_11627,N_11707);
nand U12335 (N_12335,N_11894,N_11898);
nor U12336 (N_12336,N_11542,N_11895);
nor U12337 (N_12337,N_11600,N_11698);
nor U12338 (N_12338,N_11736,N_11916);
xor U12339 (N_12339,N_11855,N_11646);
xor U12340 (N_12340,N_11731,N_11704);
xnor U12341 (N_12341,N_11623,N_11861);
or U12342 (N_12342,N_11940,N_11792);
nand U12343 (N_12343,N_11775,N_11626);
nor U12344 (N_12344,N_11944,N_11870);
or U12345 (N_12345,N_11611,N_11882);
nand U12346 (N_12346,N_11565,N_11997);
and U12347 (N_12347,N_11673,N_11736);
or U12348 (N_12348,N_11586,N_11613);
or U12349 (N_12349,N_11595,N_11901);
nor U12350 (N_12350,N_11661,N_11617);
nand U12351 (N_12351,N_11957,N_11609);
and U12352 (N_12352,N_11656,N_11733);
xnor U12353 (N_12353,N_11714,N_11689);
and U12354 (N_12354,N_11518,N_11822);
and U12355 (N_12355,N_11628,N_11803);
nand U12356 (N_12356,N_11835,N_11649);
nand U12357 (N_12357,N_11642,N_11714);
or U12358 (N_12358,N_11769,N_11615);
nor U12359 (N_12359,N_11941,N_11739);
or U12360 (N_12360,N_11522,N_11592);
xor U12361 (N_12361,N_11666,N_11798);
or U12362 (N_12362,N_11849,N_11786);
nor U12363 (N_12363,N_11502,N_11909);
xnor U12364 (N_12364,N_11666,N_11931);
and U12365 (N_12365,N_11600,N_11976);
xor U12366 (N_12366,N_11781,N_11598);
xnor U12367 (N_12367,N_11873,N_11648);
nor U12368 (N_12368,N_11647,N_11520);
or U12369 (N_12369,N_11770,N_11578);
nor U12370 (N_12370,N_11830,N_11880);
and U12371 (N_12371,N_11529,N_11952);
or U12372 (N_12372,N_11805,N_11645);
nand U12373 (N_12373,N_11870,N_11769);
xor U12374 (N_12374,N_11708,N_11912);
nand U12375 (N_12375,N_11959,N_11815);
or U12376 (N_12376,N_11909,N_11733);
or U12377 (N_12377,N_11929,N_11925);
or U12378 (N_12378,N_11568,N_11658);
and U12379 (N_12379,N_11838,N_11951);
nor U12380 (N_12380,N_11596,N_11900);
xor U12381 (N_12381,N_11661,N_11677);
and U12382 (N_12382,N_11699,N_11754);
nor U12383 (N_12383,N_11996,N_11927);
and U12384 (N_12384,N_11823,N_11717);
or U12385 (N_12385,N_11786,N_11742);
or U12386 (N_12386,N_11983,N_11666);
xnor U12387 (N_12387,N_11908,N_11948);
xor U12388 (N_12388,N_11896,N_11970);
nand U12389 (N_12389,N_11835,N_11719);
nor U12390 (N_12390,N_11624,N_11541);
or U12391 (N_12391,N_11743,N_11586);
and U12392 (N_12392,N_11991,N_11645);
xnor U12393 (N_12393,N_11738,N_11683);
nand U12394 (N_12394,N_11991,N_11992);
and U12395 (N_12395,N_11692,N_11534);
or U12396 (N_12396,N_11659,N_11767);
nand U12397 (N_12397,N_11787,N_11768);
nand U12398 (N_12398,N_11888,N_11750);
nor U12399 (N_12399,N_11680,N_11957);
and U12400 (N_12400,N_11837,N_11865);
nand U12401 (N_12401,N_11744,N_11659);
xor U12402 (N_12402,N_11897,N_11855);
or U12403 (N_12403,N_11657,N_11731);
nand U12404 (N_12404,N_11732,N_11688);
or U12405 (N_12405,N_11779,N_11623);
and U12406 (N_12406,N_11737,N_11647);
xnor U12407 (N_12407,N_11896,N_11621);
and U12408 (N_12408,N_11919,N_11718);
and U12409 (N_12409,N_11835,N_11822);
or U12410 (N_12410,N_11732,N_11500);
xnor U12411 (N_12411,N_11575,N_11759);
nor U12412 (N_12412,N_11618,N_11883);
and U12413 (N_12413,N_11912,N_11856);
xnor U12414 (N_12414,N_11689,N_11632);
and U12415 (N_12415,N_11600,N_11536);
and U12416 (N_12416,N_11760,N_11627);
or U12417 (N_12417,N_11979,N_11974);
nand U12418 (N_12418,N_11517,N_11589);
xnor U12419 (N_12419,N_11875,N_11958);
or U12420 (N_12420,N_11539,N_11612);
nor U12421 (N_12421,N_11591,N_11924);
and U12422 (N_12422,N_11683,N_11583);
nand U12423 (N_12423,N_11853,N_11839);
or U12424 (N_12424,N_11721,N_11541);
or U12425 (N_12425,N_11534,N_11744);
and U12426 (N_12426,N_11761,N_11607);
nand U12427 (N_12427,N_11763,N_11754);
nand U12428 (N_12428,N_11633,N_11784);
xnor U12429 (N_12429,N_11909,N_11732);
xnor U12430 (N_12430,N_11692,N_11779);
nor U12431 (N_12431,N_11688,N_11604);
nor U12432 (N_12432,N_11573,N_11682);
nand U12433 (N_12433,N_11677,N_11573);
and U12434 (N_12434,N_11523,N_11666);
xor U12435 (N_12435,N_11850,N_11717);
nand U12436 (N_12436,N_11571,N_11636);
xnor U12437 (N_12437,N_11873,N_11552);
nor U12438 (N_12438,N_11508,N_11996);
nand U12439 (N_12439,N_11786,N_11785);
nor U12440 (N_12440,N_11670,N_11659);
xnor U12441 (N_12441,N_11960,N_11583);
xor U12442 (N_12442,N_11919,N_11951);
and U12443 (N_12443,N_11994,N_11992);
nor U12444 (N_12444,N_11948,N_11568);
or U12445 (N_12445,N_11958,N_11973);
nand U12446 (N_12446,N_11788,N_11694);
or U12447 (N_12447,N_11641,N_11818);
nand U12448 (N_12448,N_11955,N_11985);
and U12449 (N_12449,N_11562,N_11944);
xnor U12450 (N_12450,N_11796,N_11636);
xor U12451 (N_12451,N_11530,N_11926);
nand U12452 (N_12452,N_11547,N_11683);
and U12453 (N_12453,N_11524,N_11893);
nor U12454 (N_12454,N_11829,N_11951);
nand U12455 (N_12455,N_11540,N_11849);
nand U12456 (N_12456,N_11661,N_11957);
or U12457 (N_12457,N_11588,N_11796);
or U12458 (N_12458,N_11627,N_11973);
nor U12459 (N_12459,N_11686,N_11559);
or U12460 (N_12460,N_11982,N_11947);
nor U12461 (N_12461,N_11676,N_11947);
nor U12462 (N_12462,N_11947,N_11813);
or U12463 (N_12463,N_11876,N_11810);
nand U12464 (N_12464,N_11564,N_11611);
xnor U12465 (N_12465,N_11742,N_11764);
xor U12466 (N_12466,N_11629,N_11806);
or U12467 (N_12467,N_11567,N_11627);
or U12468 (N_12468,N_11534,N_11943);
or U12469 (N_12469,N_11814,N_11785);
nand U12470 (N_12470,N_11747,N_11885);
xnor U12471 (N_12471,N_11885,N_11702);
nand U12472 (N_12472,N_11691,N_11562);
xnor U12473 (N_12473,N_11770,N_11645);
or U12474 (N_12474,N_11902,N_11986);
or U12475 (N_12475,N_11989,N_11744);
nor U12476 (N_12476,N_11571,N_11666);
and U12477 (N_12477,N_11725,N_11723);
and U12478 (N_12478,N_11859,N_11845);
nor U12479 (N_12479,N_11622,N_11713);
or U12480 (N_12480,N_11914,N_11665);
nor U12481 (N_12481,N_11500,N_11865);
xnor U12482 (N_12482,N_11953,N_11847);
nand U12483 (N_12483,N_11559,N_11875);
nand U12484 (N_12484,N_11598,N_11966);
nor U12485 (N_12485,N_11987,N_11542);
nand U12486 (N_12486,N_11976,N_11569);
xor U12487 (N_12487,N_11776,N_11860);
nor U12488 (N_12488,N_11829,N_11719);
nand U12489 (N_12489,N_11991,N_11915);
xor U12490 (N_12490,N_11628,N_11712);
and U12491 (N_12491,N_11951,N_11586);
nand U12492 (N_12492,N_11695,N_11590);
or U12493 (N_12493,N_11631,N_11892);
or U12494 (N_12494,N_11921,N_11738);
and U12495 (N_12495,N_11964,N_11680);
xnor U12496 (N_12496,N_11936,N_11616);
nor U12497 (N_12497,N_11504,N_11816);
and U12498 (N_12498,N_11705,N_11666);
nor U12499 (N_12499,N_11583,N_11581);
nand U12500 (N_12500,N_12358,N_12123);
nand U12501 (N_12501,N_12429,N_12459);
nand U12502 (N_12502,N_12023,N_12419);
nand U12503 (N_12503,N_12461,N_12261);
nor U12504 (N_12504,N_12345,N_12487);
and U12505 (N_12505,N_12154,N_12399);
and U12506 (N_12506,N_12485,N_12428);
nand U12507 (N_12507,N_12439,N_12478);
and U12508 (N_12508,N_12258,N_12144);
nand U12509 (N_12509,N_12114,N_12296);
nor U12510 (N_12510,N_12218,N_12375);
nand U12511 (N_12511,N_12432,N_12416);
nor U12512 (N_12512,N_12221,N_12318);
or U12513 (N_12513,N_12119,N_12196);
or U12514 (N_12514,N_12105,N_12452);
and U12515 (N_12515,N_12092,N_12472);
and U12516 (N_12516,N_12165,N_12143);
and U12517 (N_12517,N_12276,N_12403);
xor U12518 (N_12518,N_12083,N_12237);
xor U12519 (N_12519,N_12268,N_12273);
and U12520 (N_12520,N_12166,N_12342);
nor U12521 (N_12521,N_12423,N_12017);
or U12522 (N_12522,N_12495,N_12010);
nand U12523 (N_12523,N_12393,N_12175);
and U12524 (N_12524,N_12027,N_12022);
nand U12525 (N_12525,N_12104,N_12325);
or U12526 (N_12526,N_12142,N_12064);
nand U12527 (N_12527,N_12321,N_12238);
xnor U12528 (N_12528,N_12414,N_12217);
xor U12529 (N_12529,N_12449,N_12193);
xnor U12530 (N_12530,N_12251,N_12016);
or U12531 (N_12531,N_12332,N_12267);
or U12532 (N_12532,N_12149,N_12320);
xor U12533 (N_12533,N_12112,N_12444);
nor U12534 (N_12534,N_12089,N_12365);
or U12535 (N_12535,N_12397,N_12011);
nor U12536 (N_12536,N_12229,N_12265);
nand U12537 (N_12537,N_12285,N_12479);
xnor U12538 (N_12538,N_12354,N_12041);
xor U12539 (N_12539,N_12454,N_12313);
nor U12540 (N_12540,N_12445,N_12434);
nor U12541 (N_12541,N_12197,N_12029);
nand U12542 (N_12542,N_12299,N_12422);
or U12543 (N_12543,N_12006,N_12385);
xnor U12544 (N_12544,N_12033,N_12326);
xor U12545 (N_12545,N_12132,N_12026);
and U12546 (N_12546,N_12443,N_12486);
and U12547 (N_12547,N_12097,N_12341);
xnor U12548 (N_12548,N_12427,N_12236);
xor U12549 (N_12549,N_12338,N_12304);
xor U12550 (N_12550,N_12492,N_12073);
and U12551 (N_12551,N_12187,N_12199);
nand U12552 (N_12552,N_12362,N_12188);
xor U12553 (N_12553,N_12205,N_12139);
nand U12554 (N_12554,N_12038,N_12030);
nor U12555 (N_12555,N_12171,N_12085);
and U12556 (N_12556,N_12093,N_12348);
nor U12557 (N_12557,N_12135,N_12212);
nand U12558 (N_12558,N_12448,N_12283);
xnor U12559 (N_12559,N_12252,N_12044);
nand U12560 (N_12560,N_12262,N_12308);
or U12561 (N_12561,N_12344,N_12213);
nand U12562 (N_12562,N_12015,N_12303);
nand U12563 (N_12563,N_12413,N_12256);
and U12564 (N_12564,N_12289,N_12189);
and U12565 (N_12565,N_12441,N_12369);
or U12566 (N_12566,N_12014,N_12065);
nor U12567 (N_12567,N_12491,N_12079);
xnor U12568 (N_12568,N_12248,N_12253);
or U12569 (N_12569,N_12179,N_12355);
nand U12570 (N_12570,N_12181,N_12328);
nand U12571 (N_12571,N_12271,N_12186);
and U12572 (N_12572,N_12447,N_12130);
or U12573 (N_12573,N_12474,N_12060);
nand U12574 (N_12574,N_12408,N_12168);
or U12575 (N_12575,N_12316,N_12162);
and U12576 (N_12576,N_12002,N_12282);
xnor U12577 (N_12577,N_12336,N_12363);
xnor U12578 (N_12578,N_12476,N_12263);
xor U12579 (N_12579,N_12215,N_12400);
or U12580 (N_12580,N_12438,N_12203);
xor U12581 (N_12581,N_12047,N_12176);
xnor U12582 (N_12582,N_12124,N_12008);
and U12583 (N_12583,N_12173,N_12298);
or U12584 (N_12584,N_12395,N_12402);
xnor U12585 (N_12585,N_12063,N_12466);
xnor U12586 (N_12586,N_12169,N_12202);
or U12587 (N_12587,N_12453,N_12074);
and U12588 (N_12588,N_12421,N_12319);
or U12589 (N_12589,N_12086,N_12446);
and U12590 (N_12590,N_12099,N_12228);
nand U12591 (N_12591,N_12482,N_12350);
and U12592 (N_12592,N_12425,N_12394);
nand U12593 (N_12593,N_12100,N_12404);
nor U12594 (N_12594,N_12084,N_12061);
and U12595 (N_12595,N_12147,N_12463);
xor U12596 (N_12596,N_12172,N_12386);
or U12597 (N_12597,N_12158,N_12223);
and U12598 (N_12598,N_12225,N_12066);
nand U12599 (N_12599,N_12483,N_12475);
nor U12600 (N_12600,N_12286,N_12052);
and U12601 (N_12601,N_12347,N_12120);
xnor U12602 (N_12602,N_12156,N_12163);
nand U12603 (N_12603,N_12108,N_12287);
and U12604 (N_12604,N_12309,N_12246);
or U12605 (N_12605,N_12259,N_12284);
and U12606 (N_12606,N_12349,N_12426);
nor U12607 (N_12607,N_12109,N_12324);
nor U12608 (N_12608,N_12477,N_12496);
nand U12609 (N_12609,N_12056,N_12059);
and U12610 (N_12610,N_12398,N_12323);
nor U12611 (N_12611,N_12220,N_12437);
or U12612 (N_12612,N_12161,N_12288);
or U12613 (N_12613,N_12281,N_12095);
or U12614 (N_12614,N_12494,N_12498);
and U12615 (N_12615,N_12372,N_12230);
nor U12616 (N_12616,N_12357,N_12035);
and U12617 (N_12617,N_12159,N_12242);
xor U12618 (N_12618,N_12300,N_12272);
or U12619 (N_12619,N_12037,N_12315);
and U12620 (N_12620,N_12388,N_12292);
nor U12621 (N_12621,N_12160,N_12270);
nand U12622 (N_12622,N_12103,N_12182);
and U12623 (N_12623,N_12127,N_12266);
and U12624 (N_12624,N_12293,N_12210);
nand U12625 (N_12625,N_12361,N_12028);
xor U12626 (N_12626,N_12232,N_12126);
or U12627 (N_12627,N_12254,N_12250);
nor U12628 (N_12628,N_12106,N_12180);
or U12629 (N_12629,N_12279,N_12122);
or U12630 (N_12630,N_12275,N_12264);
and U12631 (N_12631,N_12136,N_12278);
nand U12632 (N_12632,N_12244,N_12077);
nor U12633 (N_12633,N_12457,N_12098);
nand U12634 (N_12634,N_12311,N_12484);
xnor U12635 (N_12635,N_12116,N_12024);
or U12636 (N_12636,N_12164,N_12465);
xor U12637 (N_12637,N_12378,N_12310);
and U12638 (N_12638,N_12231,N_12013);
xnor U12639 (N_12639,N_12034,N_12260);
nand U12640 (N_12640,N_12201,N_12155);
and U12641 (N_12641,N_12359,N_12392);
nor U12642 (N_12642,N_12499,N_12115);
and U12643 (N_12643,N_12456,N_12227);
or U12644 (N_12644,N_12054,N_12473);
nand U12645 (N_12645,N_12157,N_12036);
and U12646 (N_12646,N_12051,N_12458);
and U12647 (N_12647,N_12269,N_12333);
or U12648 (N_12648,N_12235,N_12364);
or U12649 (N_12649,N_12469,N_12101);
xnor U12650 (N_12650,N_12433,N_12405);
xnor U12651 (N_12651,N_12080,N_12178);
nand U12652 (N_12652,N_12489,N_12368);
and U12653 (N_12653,N_12078,N_12317);
xnor U12654 (N_12654,N_12409,N_12045);
nand U12655 (N_12655,N_12490,N_12305);
nor U12656 (N_12656,N_12071,N_12468);
or U12657 (N_12657,N_12396,N_12090);
or U12658 (N_12658,N_12440,N_12493);
or U12659 (N_12659,N_12420,N_12330);
nor U12660 (N_12660,N_12206,N_12129);
xor U12661 (N_12661,N_12376,N_12185);
xor U12662 (N_12662,N_12379,N_12401);
nor U12663 (N_12663,N_12407,N_12069);
nor U12664 (N_12664,N_12214,N_12410);
and U12665 (N_12665,N_12110,N_12340);
nand U12666 (N_12666,N_12343,N_12140);
and U12667 (N_12667,N_12255,N_12111);
nor U12668 (N_12668,N_12004,N_12001);
xor U12669 (N_12669,N_12249,N_12216);
or U12670 (N_12670,N_12137,N_12222);
xnor U12671 (N_12671,N_12418,N_12415);
and U12672 (N_12672,N_12057,N_12053);
or U12673 (N_12673,N_12153,N_12209);
xnor U12674 (N_12674,N_12234,N_12373);
or U12675 (N_12675,N_12370,N_12005);
nor U12676 (N_12676,N_12346,N_12204);
nand U12677 (N_12677,N_12380,N_12208);
xnor U12678 (N_12678,N_12068,N_12226);
xor U12679 (N_12679,N_12207,N_12290);
or U12680 (N_12680,N_12128,N_12058);
nor U12681 (N_12681,N_12134,N_12314);
nor U12682 (N_12682,N_12480,N_12460);
nor U12683 (N_12683,N_12118,N_12088);
nand U12684 (N_12684,N_12383,N_12121);
nor U12685 (N_12685,N_12335,N_12436);
xnor U12686 (N_12686,N_12481,N_12020);
or U12687 (N_12687,N_12012,N_12067);
nand U12688 (N_12688,N_12257,N_12497);
xor U12689 (N_12689,N_12007,N_12455);
xnor U12690 (N_12690,N_12025,N_12247);
nand U12691 (N_12691,N_12450,N_12471);
xor U12692 (N_12692,N_12046,N_12451);
nor U12693 (N_12693,N_12224,N_12243);
or U12694 (N_12694,N_12072,N_12151);
nor U12695 (N_12695,N_12177,N_12117);
nor U12696 (N_12696,N_12003,N_12170);
nand U12697 (N_12697,N_12371,N_12145);
nand U12698 (N_12698,N_12240,N_12295);
and U12699 (N_12699,N_12055,N_12239);
and U12700 (N_12700,N_12138,N_12424);
and U12701 (N_12701,N_12417,N_12076);
or U12702 (N_12702,N_12096,N_12062);
nor U12703 (N_12703,N_12102,N_12150);
nor U12704 (N_12704,N_12297,N_12019);
or U12705 (N_12705,N_12294,N_12352);
and U12706 (N_12706,N_12133,N_12322);
nor U12707 (N_12707,N_12339,N_12241);
and U12708 (N_12708,N_12442,N_12167);
xnor U12709 (N_12709,N_12467,N_12391);
xor U12710 (N_12710,N_12430,N_12356);
and U12711 (N_12711,N_12087,N_12192);
nand U12712 (N_12712,N_12367,N_12000);
and U12713 (N_12713,N_12245,N_12462);
nand U12714 (N_12714,N_12184,N_12406);
nand U12715 (N_12715,N_12374,N_12306);
nand U12716 (N_12716,N_12190,N_12148);
xnor U12717 (N_12717,N_12048,N_12360);
xnor U12718 (N_12718,N_12377,N_12031);
and U12719 (N_12719,N_12280,N_12146);
nor U12720 (N_12720,N_12301,N_12277);
xor U12721 (N_12721,N_12195,N_12329);
nor U12722 (N_12722,N_12113,N_12435);
and U12723 (N_12723,N_12381,N_12039);
nor U12724 (N_12724,N_12040,N_12200);
xor U12725 (N_12725,N_12464,N_12312);
and U12726 (N_12726,N_12152,N_12291);
nor U12727 (N_12727,N_12387,N_12141);
and U12728 (N_12728,N_12183,N_12351);
and U12729 (N_12729,N_12081,N_12198);
and U12730 (N_12730,N_12082,N_12233);
and U12731 (N_12731,N_12337,N_12032);
nand U12732 (N_12732,N_12353,N_12470);
nand U12733 (N_12733,N_12049,N_12043);
or U12734 (N_12734,N_12411,N_12125);
nor U12735 (N_12735,N_12382,N_12050);
and U12736 (N_12736,N_12307,N_12091);
and U12737 (N_12737,N_12219,N_12131);
nor U12738 (N_12738,N_12274,N_12021);
or U12739 (N_12739,N_12327,N_12174);
nor U12740 (N_12740,N_12390,N_12384);
nor U12741 (N_12741,N_12191,N_12302);
or U12742 (N_12742,N_12488,N_12018);
and U12743 (N_12743,N_12334,N_12331);
nor U12744 (N_12744,N_12070,N_12094);
nor U12745 (N_12745,N_12042,N_12075);
xnor U12746 (N_12746,N_12366,N_12211);
or U12747 (N_12747,N_12107,N_12389);
or U12748 (N_12748,N_12194,N_12009);
nand U12749 (N_12749,N_12412,N_12431);
and U12750 (N_12750,N_12042,N_12218);
and U12751 (N_12751,N_12063,N_12393);
or U12752 (N_12752,N_12254,N_12454);
or U12753 (N_12753,N_12282,N_12371);
and U12754 (N_12754,N_12404,N_12381);
and U12755 (N_12755,N_12301,N_12186);
nand U12756 (N_12756,N_12317,N_12185);
or U12757 (N_12757,N_12479,N_12027);
nor U12758 (N_12758,N_12402,N_12238);
nand U12759 (N_12759,N_12411,N_12224);
xor U12760 (N_12760,N_12435,N_12180);
nand U12761 (N_12761,N_12220,N_12462);
xor U12762 (N_12762,N_12461,N_12447);
nor U12763 (N_12763,N_12286,N_12032);
nand U12764 (N_12764,N_12426,N_12086);
or U12765 (N_12765,N_12370,N_12380);
nor U12766 (N_12766,N_12080,N_12316);
and U12767 (N_12767,N_12021,N_12192);
or U12768 (N_12768,N_12438,N_12386);
xnor U12769 (N_12769,N_12446,N_12063);
and U12770 (N_12770,N_12224,N_12041);
nand U12771 (N_12771,N_12368,N_12315);
and U12772 (N_12772,N_12389,N_12370);
nor U12773 (N_12773,N_12416,N_12176);
nor U12774 (N_12774,N_12221,N_12026);
xnor U12775 (N_12775,N_12153,N_12369);
or U12776 (N_12776,N_12341,N_12139);
nand U12777 (N_12777,N_12350,N_12156);
and U12778 (N_12778,N_12493,N_12264);
nor U12779 (N_12779,N_12343,N_12224);
nor U12780 (N_12780,N_12295,N_12289);
and U12781 (N_12781,N_12376,N_12239);
and U12782 (N_12782,N_12221,N_12200);
nor U12783 (N_12783,N_12219,N_12096);
and U12784 (N_12784,N_12405,N_12331);
or U12785 (N_12785,N_12107,N_12461);
xnor U12786 (N_12786,N_12143,N_12365);
nor U12787 (N_12787,N_12055,N_12312);
xor U12788 (N_12788,N_12421,N_12185);
xor U12789 (N_12789,N_12401,N_12196);
and U12790 (N_12790,N_12124,N_12445);
xor U12791 (N_12791,N_12084,N_12206);
or U12792 (N_12792,N_12335,N_12297);
nand U12793 (N_12793,N_12459,N_12298);
nand U12794 (N_12794,N_12256,N_12283);
nor U12795 (N_12795,N_12406,N_12426);
nor U12796 (N_12796,N_12331,N_12481);
nand U12797 (N_12797,N_12077,N_12087);
nand U12798 (N_12798,N_12448,N_12467);
or U12799 (N_12799,N_12390,N_12488);
and U12800 (N_12800,N_12193,N_12155);
and U12801 (N_12801,N_12430,N_12224);
or U12802 (N_12802,N_12032,N_12120);
or U12803 (N_12803,N_12222,N_12276);
and U12804 (N_12804,N_12204,N_12077);
and U12805 (N_12805,N_12435,N_12426);
nand U12806 (N_12806,N_12464,N_12336);
or U12807 (N_12807,N_12003,N_12140);
nor U12808 (N_12808,N_12074,N_12393);
xnor U12809 (N_12809,N_12011,N_12396);
and U12810 (N_12810,N_12196,N_12457);
and U12811 (N_12811,N_12147,N_12066);
or U12812 (N_12812,N_12166,N_12128);
xor U12813 (N_12813,N_12045,N_12496);
nor U12814 (N_12814,N_12409,N_12275);
nor U12815 (N_12815,N_12006,N_12043);
nand U12816 (N_12816,N_12382,N_12238);
xnor U12817 (N_12817,N_12130,N_12149);
nand U12818 (N_12818,N_12382,N_12240);
or U12819 (N_12819,N_12361,N_12069);
and U12820 (N_12820,N_12311,N_12485);
xnor U12821 (N_12821,N_12066,N_12345);
xor U12822 (N_12822,N_12045,N_12073);
xor U12823 (N_12823,N_12450,N_12205);
and U12824 (N_12824,N_12245,N_12391);
nor U12825 (N_12825,N_12235,N_12489);
xnor U12826 (N_12826,N_12468,N_12331);
and U12827 (N_12827,N_12257,N_12256);
nor U12828 (N_12828,N_12379,N_12158);
or U12829 (N_12829,N_12178,N_12236);
xnor U12830 (N_12830,N_12481,N_12146);
xor U12831 (N_12831,N_12126,N_12038);
or U12832 (N_12832,N_12392,N_12272);
nor U12833 (N_12833,N_12386,N_12144);
xnor U12834 (N_12834,N_12264,N_12199);
nand U12835 (N_12835,N_12479,N_12421);
xor U12836 (N_12836,N_12347,N_12107);
nor U12837 (N_12837,N_12262,N_12130);
or U12838 (N_12838,N_12162,N_12491);
xor U12839 (N_12839,N_12223,N_12119);
and U12840 (N_12840,N_12248,N_12027);
and U12841 (N_12841,N_12036,N_12127);
and U12842 (N_12842,N_12384,N_12241);
or U12843 (N_12843,N_12467,N_12067);
or U12844 (N_12844,N_12188,N_12218);
nand U12845 (N_12845,N_12474,N_12212);
or U12846 (N_12846,N_12115,N_12109);
nor U12847 (N_12847,N_12351,N_12045);
and U12848 (N_12848,N_12247,N_12027);
xnor U12849 (N_12849,N_12189,N_12474);
or U12850 (N_12850,N_12475,N_12341);
xor U12851 (N_12851,N_12151,N_12088);
or U12852 (N_12852,N_12229,N_12361);
or U12853 (N_12853,N_12037,N_12380);
nand U12854 (N_12854,N_12108,N_12121);
nand U12855 (N_12855,N_12303,N_12121);
nor U12856 (N_12856,N_12213,N_12150);
xor U12857 (N_12857,N_12161,N_12025);
nand U12858 (N_12858,N_12198,N_12259);
nor U12859 (N_12859,N_12313,N_12124);
xnor U12860 (N_12860,N_12193,N_12122);
xnor U12861 (N_12861,N_12139,N_12317);
and U12862 (N_12862,N_12412,N_12287);
xnor U12863 (N_12863,N_12355,N_12465);
nand U12864 (N_12864,N_12359,N_12095);
and U12865 (N_12865,N_12357,N_12011);
and U12866 (N_12866,N_12462,N_12104);
nor U12867 (N_12867,N_12361,N_12239);
or U12868 (N_12868,N_12117,N_12248);
nand U12869 (N_12869,N_12009,N_12178);
nor U12870 (N_12870,N_12158,N_12277);
nor U12871 (N_12871,N_12401,N_12482);
or U12872 (N_12872,N_12224,N_12165);
or U12873 (N_12873,N_12430,N_12223);
or U12874 (N_12874,N_12026,N_12029);
nor U12875 (N_12875,N_12456,N_12441);
nor U12876 (N_12876,N_12081,N_12276);
and U12877 (N_12877,N_12207,N_12163);
nor U12878 (N_12878,N_12390,N_12346);
nor U12879 (N_12879,N_12136,N_12284);
or U12880 (N_12880,N_12331,N_12417);
nor U12881 (N_12881,N_12054,N_12411);
nand U12882 (N_12882,N_12348,N_12267);
nand U12883 (N_12883,N_12354,N_12022);
nand U12884 (N_12884,N_12412,N_12271);
xnor U12885 (N_12885,N_12039,N_12397);
or U12886 (N_12886,N_12033,N_12131);
nor U12887 (N_12887,N_12485,N_12010);
nor U12888 (N_12888,N_12444,N_12207);
nor U12889 (N_12889,N_12299,N_12451);
nor U12890 (N_12890,N_12029,N_12172);
xnor U12891 (N_12891,N_12006,N_12351);
and U12892 (N_12892,N_12272,N_12296);
and U12893 (N_12893,N_12422,N_12374);
and U12894 (N_12894,N_12474,N_12419);
nand U12895 (N_12895,N_12265,N_12288);
nand U12896 (N_12896,N_12355,N_12391);
and U12897 (N_12897,N_12446,N_12088);
and U12898 (N_12898,N_12372,N_12448);
xor U12899 (N_12899,N_12290,N_12040);
or U12900 (N_12900,N_12035,N_12298);
nor U12901 (N_12901,N_12038,N_12231);
nor U12902 (N_12902,N_12129,N_12119);
nand U12903 (N_12903,N_12184,N_12490);
and U12904 (N_12904,N_12168,N_12176);
and U12905 (N_12905,N_12161,N_12314);
or U12906 (N_12906,N_12000,N_12327);
nor U12907 (N_12907,N_12423,N_12417);
nand U12908 (N_12908,N_12477,N_12083);
nor U12909 (N_12909,N_12381,N_12493);
nand U12910 (N_12910,N_12302,N_12452);
or U12911 (N_12911,N_12166,N_12326);
or U12912 (N_12912,N_12303,N_12481);
or U12913 (N_12913,N_12361,N_12149);
xnor U12914 (N_12914,N_12016,N_12150);
or U12915 (N_12915,N_12240,N_12192);
and U12916 (N_12916,N_12391,N_12222);
xnor U12917 (N_12917,N_12126,N_12304);
xor U12918 (N_12918,N_12454,N_12388);
nor U12919 (N_12919,N_12374,N_12423);
nand U12920 (N_12920,N_12233,N_12077);
xor U12921 (N_12921,N_12008,N_12459);
nand U12922 (N_12922,N_12370,N_12001);
and U12923 (N_12923,N_12189,N_12343);
nor U12924 (N_12924,N_12021,N_12070);
and U12925 (N_12925,N_12278,N_12233);
nor U12926 (N_12926,N_12419,N_12000);
nor U12927 (N_12927,N_12458,N_12404);
nand U12928 (N_12928,N_12048,N_12215);
or U12929 (N_12929,N_12153,N_12307);
nor U12930 (N_12930,N_12455,N_12344);
or U12931 (N_12931,N_12188,N_12290);
nor U12932 (N_12932,N_12126,N_12005);
xnor U12933 (N_12933,N_12230,N_12276);
or U12934 (N_12934,N_12393,N_12448);
or U12935 (N_12935,N_12072,N_12248);
nor U12936 (N_12936,N_12088,N_12325);
nor U12937 (N_12937,N_12105,N_12003);
xor U12938 (N_12938,N_12299,N_12472);
nor U12939 (N_12939,N_12429,N_12244);
xnor U12940 (N_12940,N_12447,N_12279);
nor U12941 (N_12941,N_12151,N_12458);
nor U12942 (N_12942,N_12492,N_12055);
nor U12943 (N_12943,N_12487,N_12046);
nor U12944 (N_12944,N_12225,N_12267);
and U12945 (N_12945,N_12425,N_12286);
and U12946 (N_12946,N_12231,N_12164);
nor U12947 (N_12947,N_12194,N_12372);
or U12948 (N_12948,N_12321,N_12259);
or U12949 (N_12949,N_12263,N_12472);
or U12950 (N_12950,N_12279,N_12285);
and U12951 (N_12951,N_12496,N_12302);
and U12952 (N_12952,N_12446,N_12409);
and U12953 (N_12953,N_12418,N_12056);
xor U12954 (N_12954,N_12134,N_12130);
nor U12955 (N_12955,N_12343,N_12193);
or U12956 (N_12956,N_12352,N_12072);
and U12957 (N_12957,N_12188,N_12462);
nand U12958 (N_12958,N_12193,N_12194);
nor U12959 (N_12959,N_12366,N_12338);
nand U12960 (N_12960,N_12280,N_12476);
and U12961 (N_12961,N_12194,N_12138);
or U12962 (N_12962,N_12258,N_12132);
or U12963 (N_12963,N_12411,N_12484);
or U12964 (N_12964,N_12264,N_12386);
nand U12965 (N_12965,N_12193,N_12008);
nor U12966 (N_12966,N_12235,N_12111);
and U12967 (N_12967,N_12216,N_12053);
and U12968 (N_12968,N_12120,N_12270);
nand U12969 (N_12969,N_12007,N_12299);
nand U12970 (N_12970,N_12166,N_12363);
xnor U12971 (N_12971,N_12236,N_12185);
or U12972 (N_12972,N_12294,N_12040);
nand U12973 (N_12973,N_12071,N_12480);
xor U12974 (N_12974,N_12424,N_12000);
or U12975 (N_12975,N_12253,N_12074);
xnor U12976 (N_12976,N_12356,N_12463);
or U12977 (N_12977,N_12002,N_12000);
and U12978 (N_12978,N_12246,N_12433);
nand U12979 (N_12979,N_12352,N_12276);
nor U12980 (N_12980,N_12143,N_12422);
and U12981 (N_12981,N_12167,N_12471);
nor U12982 (N_12982,N_12220,N_12203);
xor U12983 (N_12983,N_12210,N_12277);
nand U12984 (N_12984,N_12395,N_12308);
or U12985 (N_12985,N_12340,N_12009);
and U12986 (N_12986,N_12409,N_12278);
nand U12987 (N_12987,N_12468,N_12201);
xor U12988 (N_12988,N_12496,N_12283);
nand U12989 (N_12989,N_12084,N_12382);
and U12990 (N_12990,N_12088,N_12369);
and U12991 (N_12991,N_12198,N_12476);
xor U12992 (N_12992,N_12442,N_12185);
nor U12993 (N_12993,N_12425,N_12056);
nand U12994 (N_12994,N_12380,N_12221);
nand U12995 (N_12995,N_12369,N_12351);
and U12996 (N_12996,N_12192,N_12293);
or U12997 (N_12997,N_12226,N_12431);
nand U12998 (N_12998,N_12205,N_12327);
nor U12999 (N_12999,N_12471,N_12402);
nor U13000 (N_13000,N_12899,N_12952);
nor U13001 (N_13001,N_12789,N_12800);
nor U13002 (N_13002,N_12583,N_12860);
and U13003 (N_13003,N_12825,N_12528);
or U13004 (N_13004,N_12763,N_12891);
or U13005 (N_13005,N_12549,N_12653);
nand U13006 (N_13006,N_12513,N_12775);
nand U13007 (N_13007,N_12957,N_12872);
nor U13008 (N_13008,N_12881,N_12719);
or U13009 (N_13009,N_12792,N_12539);
nor U13010 (N_13010,N_12691,N_12954);
and U13011 (N_13011,N_12540,N_12922);
nand U13012 (N_13012,N_12764,N_12534);
nand U13013 (N_13013,N_12698,N_12831);
nor U13014 (N_13014,N_12619,N_12914);
or U13015 (N_13015,N_12934,N_12562);
and U13016 (N_13016,N_12620,N_12658);
xnor U13017 (N_13017,N_12911,N_12876);
or U13018 (N_13018,N_12675,N_12989);
and U13019 (N_13019,N_12793,N_12900);
nand U13020 (N_13020,N_12638,N_12595);
nand U13021 (N_13021,N_12566,N_12561);
xor U13022 (N_13022,N_12557,N_12897);
nand U13023 (N_13023,N_12754,N_12915);
or U13024 (N_13024,N_12762,N_12918);
nand U13025 (N_13025,N_12559,N_12929);
nand U13026 (N_13026,N_12538,N_12959);
and U13027 (N_13027,N_12953,N_12965);
nand U13028 (N_13028,N_12688,N_12515);
nor U13029 (N_13029,N_12741,N_12544);
and U13030 (N_13030,N_12610,N_12862);
nor U13031 (N_13031,N_12814,N_12655);
nand U13032 (N_13032,N_12973,N_12893);
xnor U13033 (N_13033,N_12986,N_12652);
xnor U13034 (N_13034,N_12988,N_12773);
xor U13035 (N_13035,N_12596,N_12783);
nand U13036 (N_13036,N_12729,N_12924);
xnor U13037 (N_13037,N_12590,N_12752);
nand U13038 (N_13038,N_12506,N_12903);
or U13039 (N_13039,N_12739,N_12581);
or U13040 (N_13040,N_12657,N_12574);
and U13041 (N_13041,N_12509,N_12999);
or U13042 (N_13042,N_12709,N_12807);
nand U13043 (N_13043,N_12605,N_12951);
and U13044 (N_13044,N_12659,N_12548);
xor U13045 (N_13045,N_12908,N_12874);
nand U13046 (N_13046,N_12694,N_12601);
and U13047 (N_13047,N_12907,N_12730);
xor U13048 (N_13048,N_12527,N_12828);
and U13049 (N_13049,N_12611,N_12718);
or U13050 (N_13050,N_12749,N_12871);
nand U13051 (N_13051,N_12904,N_12910);
nor U13052 (N_13052,N_12816,N_12555);
or U13053 (N_13053,N_12661,N_12568);
and U13054 (N_13054,N_12837,N_12936);
xor U13055 (N_13055,N_12608,N_12594);
nor U13056 (N_13056,N_12768,N_12507);
nand U13057 (N_13057,N_12683,N_12640);
nor U13058 (N_13058,N_12624,N_12844);
nor U13059 (N_13059,N_12933,N_12612);
xnor U13060 (N_13060,N_12804,N_12708);
nand U13061 (N_13061,N_12879,N_12846);
and U13062 (N_13062,N_12761,N_12817);
or U13063 (N_13063,N_12628,N_12545);
and U13064 (N_13064,N_12656,N_12788);
nor U13065 (N_13065,N_12790,N_12756);
nand U13066 (N_13066,N_12554,N_12815);
nand U13067 (N_13067,N_12669,N_12553);
and U13068 (N_13068,N_12636,N_12923);
and U13069 (N_13069,N_12695,N_12533);
xnor U13070 (N_13070,N_12976,N_12531);
nor U13071 (N_13071,N_12940,N_12913);
xor U13072 (N_13072,N_12681,N_12905);
xor U13073 (N_13073,N_12699,N_12550);
nor U13074 (N_13074,N_12985,N_12526);
xnor U13075 (N_13075,N_12827,N_12702);
or U13076 (N_13076,N_12774,N_12974);
and U13077 (N_13077,N_12753,N_12705);
or U13078 (N_13078,N_12637,N_12882);
or U13079 (N_13079,N_12570,N_12946);
nand U13080 (N_13080,N_12822,N_12607);
xor U13081 (N_13081,N_12832,N_12942);
or U13082 (N_13082,N_12689,N_12693);
nand U13083 (N_13083,N_12671,N_12824);
xnor U13084 (N_13084,N_12678,N_12686);
xnor U13085 (N_13085,N_12869,N_12706);
xor U13086 (N_13086,N_12674,N_12898);
xor U13087 (N_13087,N_12745,N_12618);
xor U13088 (N_13088,N_12925,N_12944);
nand U13089 (N_13089,N_12941,N_12982);
or U13090 (N_13090,N_12609,N_12731);
xnor U13091 (N_13091,N_12838,N_12896);
nor U13092 (N_13092,N_12803,N_12567);
xor U13093 (N_13093,N_12598,N_12703);
or U13094 (N_13094,N_12630,N_12808);
xnor U13095 (N_13095,N_12734,N_12950);
xnor U13096 (N_13096,N_12632,N_12737);
xnor U13097 (N_13097,N_12795,N_12516);
or U13098 (N_13098,N_12569,N_12573);
xor U13099 (N_13099,N_12771,N_12784);
and U13100 (N_13100,N_12810,N_12625);
nor U13101 (N_13101,N_12841,N_12717);
nand U13102 (N_13102,N_12585,N_12912);
xor U13103 (N_13103,N_12839,N_12766);
nor U13104 (N_13104,N_12701,N_12818);
and U13105 (N_13105,N_12530,N_12552);
nand U13106 (N_13106,N_12798,N_12830);
nor U13107 (N_13107,N_12856,N_12857);
nor U13108 (N_13108,N_12981,N_12760);
xor U13109 (N_13109,N_12820,N_12735);
xnor U13110 (N_13110,N_12592,N_12850);
or U13111 (N_13111,N_12885,N_12654);
nor U13112 (N_13112,N_12560,N_12931);
nand U13113 (N_13113,N_12575,N_12726);
nand U13114 (N_13114,N_12963,N_12863);
xnor U13115 (N_13115,N_12571,N_12895);
nor U13116 (N_13116,N_12748,N_12819);
or U13117 (N_13117,N_12889,N_12725);
nor U13118 (N_13118,N_12578,N_12835);
nand U13119 (N_13119,N_12712,N_12504);
nor U13120 (N_13120,N_12853,N_12958);
or U13121 (N_13121,N_12584,N_12955);
and U13122 (N_13122,N_12642,N_12978);
nand U13123 (N_13123,N_12859,N_12649);
or U13124 (N_13124,N_12597,N_12870);
nor U13125 (N_13125,N_12517,N_12909);
nand U13126 (N_13126,N_12970,N_12956);
nand U13127 (N_13127,N_12687,N_12582);
xor U13128 (N_13128,N_12697,N_12794);
nand U13129 (N_13129,N_12556,N_12679);
and U13130 (N_13130,N_12997,N_12892);
or U13131 (N_13131,N_12563,N_12724);
nor U13132 (N_13132,N_12537,N_12888);
nand U13133 (N_13133,N_12932,N_12576);
nand U13134 (N_13134,N_12919,N_12779);
or U13135 (N_13135,N_12736,N_12617);
xnor U13136 (N_13136,N_12716,N_12969);
and U13137 (N_13137,N_12738,N_12759);
nor U13138 (N_13138,N_12616,N_12505);
or U13139 (N_13139,N_12778,N_12720);
nand U13140 (N_13140,N_12510,N_12785);
and U13141 (N_13141,N_12602,N_12710);
and U13142 (N_13142,N_12757,N_12996);
nand U13143 (N_13143,N_12666,N_12979);
and U13144 (N_13144,N_12964,N_12938);
or U13145 (N_13145,N_12672,N_12707);
or U13146 (N_13146,N_12777,N_12690);
and U13147 (N_13147,N_12858,N_12758);
xor U13148 (N_13148,N_12629,N_12968);
nand U13149 (N_13149,N_12975,N_12711);
xor U13150 (N_13150,N_12668,N_12829);
and U13151 (N_13151,N_12811,N_12751);
xnor U13152 (N_13152,N_12535,N_12984);
nor U13153 (N_13153,N_12769,N_12713);
and U13154 (N_13154,N_12645,N_12805);
xnor U13155 (N_13155,N_12917,N_12728);
nor U13156 (N_13156,N_12781,N_12930);
xor U13157 (N_13157,N_12864,N_12770);
nor U13158 (N_13158,N_12623,N_12962);
nor U13159 (N_13159,N_12500,N_12626);
and U13160 (N_13160,N_12782,N_12866);
or U13161 (N_13161,N_12662,N_12684);
or U13162 (N_13162,N_12727,N_12511);
xor U13163 (N_13163,N_12847,N_12627);
nand U13164 (N_13164,N_12600,N_12884);
nor U13165 (N_13165,N_12966,N_12586);
and U13166 (N_13166,N_12634,N_12842);
and U13167 (N_13167,N_12843,N_12521);
or U13168 (N_13168,N_12833,N_12519);
xnor U13169 (N_13169,N_12767,N_12880);
nand U13170 (N_13170,N_12865,N_12928);
xnor U13171 (N_13171,N_12685,N_12834);
nor U13172 (N_13172,N_12755,N_12797);
xor U13173 (N_13173,N_12921,N_12851);
and U13174 (N_13174,N_12868,N_12643);
nor U13175 (N_13175,N_12796,N_12971);
nor U13176 (N_13176,N_12740,N_12939);
or U13177 (N_13177,N_12927,N_12572);
and U13178 (N_13178,N_12890,N_12812);
xor U13179 (N_13179,N_12967,N_12823);
xor U13180 (N_13180,N_12902,N_12943);
nand U13181 (N_13181,N_12765,N_12524);
and U13182 (N_13182,N_12503,N_12518);
nor U13183 (N_13183,N_12883,N_12821);
and U13184 (N_13184,N_12786,N_12682);
or U13185 (N_13185,N_12743,N_12648);
xor U13186 (N_13186,N_12848,N_12604);
and U13187 (N_13187,N_12529,N_12660);
xnor U13188 (N_13188,N_12680,N_12836);
or U13189 (N_13189,N_12663,N_12665);
and U13190 (N_13190,N_12901,N_12840);
nand U13191 (N_13191,N_12977,N_12809);
or U13192 (N_13192,N_12613,N_12746);
nand U13193 (N_13193,N_12541,N_12606);
xnor U13194 (N_13194,N_12960,N_12644);
and U13195 (N_13195,N_12692,N_12508);
or U13196 (N_13196,N_12599,N_12514);
xor U13197 (N_13197,N_12747,N_12700);
nand U13198 (N_13198,N_12993,N_12945);
nand U13199 (N_13199,N_12543,N_12854);
or U13200 (N_13200,N_12587,N_12542);
nor U13201 (N_13201,N_12802,N_12502);
nor U13202 (N_13202,N_12961,N_12995);
xor U13203 (N_13203,N_12520,N_12744);
nor U13204 (N_13204,N_12916,N_12647);
or U13205 (N_13205,N_12875,N_12546);
and U13206 (N_13206,N_12565,N_12992);
nand U13207 (N_13207,N_12532,N_12667);
xor U13208 (N_13208,N_12906,N_12806);
and U13209 (N_13209,N_12987,N_12877);
and U13210 (N_13210,N_12670,N_12501);
nand U13211 (N_13211,N_12742,N_12926);
and U13212 (N_13212,N_12633,N_12732);
xor U13213 (N_13213,N_12935,N_12715);
xnor U13214 (N_13214,N_12733,N_12826);
nor U13215 (N_13215,N_12522,N_12886);
or U13216 (N_13216,N_12991,N_12887);
xor U13217 (N_13217,N_12878,N_12676);
nor U13218 (N_13218,N_12787,N_12750);
nand U13219 (N_13219,N_12791,N_12949);
or U13220 (N_13220,N_12948,N_12635);
xor U13221 (N_13221,N_12813,N_12650);
xor U13222 (N_13222,N_12947,N_12799);
nor U13223 (N_13223,N_12696,N_12998);
nor U13224 (N_13224,N_12867,N_12801);
nand U13225 (N_13225,N_12536,N_12920);
nand U13226 (N_13226,N_12994,N_12722);
xnor U13227 (N_13227,N_12937,N_12631);
nand U13228 (N_13228,N_12646,N_12547);
nor U13229 (N_13229,N_12855,N_12614);
or U13230 (N_13230,N_12714,N_12641);
or U13231 (N_13231,N_12593,N_12983);
nor U13232 (N_13232,N_12564,N_12639);
nand U13233 (N_13233,N_12551,N_12673);
and U13234 (N_13234,N_12622,N_12591);
or U13235 (N_13235,N_12776,N_12664);
nor U13236 (N_13236,N_12990,N_12603);
and U13237 (N_13237,N_12723,N_12651);
and U13238 (N_13238,N_12980,N_12525);
nand U13239 (N_13239,N_12615,N_12577);
or U13240 (N_13240,N_12512,N_12523);
nor U13241 (N_13241,N_12721,N_12780);
nand U13242 (N_13242,N_12621,N_12852);
nand U13243 (N_13243,N_12589,N_12558);
xor U13244 (N_13244,N_12845,N_12580);
and U13245 (N_13245,N_12849,N_12861);
or U13246 (N_13246,N_12894,N_12704);
nand U13247 (N_13247,N_12677,N_12972);
xnor U13248 (N_13248,N_12579,N_12873);
nand U13249 (N_13249,N_12588,N_12772);
nor U13250 (N_13250,N_12869,N_12516);
nor U13251 (N_13251,N_12757,N_12849);
nor U13252 (N_13252,N_12532,N_12907);
xnor U13253 (N_13253,N_12764,N_12993);
nand U13254 (N_13254,N_12668,N_12666);
nor U13255 (N_13255,N_12807,N_12594);
nand U13256 (N_13256,N_12713,N_12506);
nor U13257 (N_13257,N_12985,N_12730);
nor U13258 (N_13258,N_12877,N_12504);
nand U13259 (N_13259,N_12823,N_12565);
nand U13260 (N_13260,N_12539,N_12921);
or U13261 (N_13261,N_12818,N_12893);
nor U13262 (N_13262,N_12741,N_12724);
and U13263 (N_13263,N_12765,N_12971);
nor U13264 (N_13264,N_12712,N_12567);
and U13265 (N_13265,N_12719,N_12870);
and U13266 (N_13266,N_12849,N_12585);
nor U13267 (N_13267,N_12684,N_12916);
xnor U13268 (N_13268,N_12661,N_12988);
nor U13269 (N_13269,N_12890,N_12622);
nor U13270 (N_13270,N_12621,N_12529);
or U13271 (N_13271,N_12558,N_12836);
xor U13272 (N_13272,N_12652,N_12928);
or U13273 (N_13273,N_12891,N_12864);
and U13274 (N_13274,N_12893,N_12947);
nor U13275 (N_13275,N_12728,N_12863);
nor U13276 (N_13276,N_12705,N_12859);
nor U13277 (N_13277,N_12890,N_12835);
nand U13278 (N_13278,N_12960,N_12828);
xor U13279 (N_13279,N_12686,N_12999);
xnor U13280 (N_13280,N_12782,N_12600);
or U13281 (N_13281,N_12881,N_12604);
or U13282 (N_13282,N_12795,N_12697);
nand U13283 (N_13283,N_12785,N_12638);
or U13284 (N_13284,N_12865,N_12671);
xor U13285 (N_13285,N_12984,N_12739);
xnor U13286 (N_13286,N_12726,N_12981);
nor U13287 (N_13287,N_12922,N_12576);
or U13288 (N_13288,N_12620,N_12661);
nand U13289 (N_13289,N_12645,N_12927);
nand U13290 (N_13290,N_12796,N_12699);
xnor U13291 (N_13291,N_12928,N_12513);
nor U13292 (N_13292,N_12902,N_12670);
nor U13293 (N_13293,N_12816,N_12864);
xnor U13294 (N_13294,N_12941,N_12593);
xnor U13295 (N_13295,N_12575,N_12549);
nor U13296 (N_13296,N_12950,N_12536);
and U13297 (N_13297,N_12896,N_12964);
nand U13298 (N_13298,N_12670,N_12926);
or U13299 (N_13299,N_12740,N_12810);
nand U13300 (N_13300,N_12911,N_12555);
nand U13301 (N_13301,N_12732,N_12523);
nor U13302 (N_13302,N_12694,N_12503);
nor U13303 (N_13303,N_12857,N_12879);
xnor U13304 (N_13304,N_12512,N_12698);
or U13305 (N_13305,N_12719,N_12981);
xor U13306 (N_13306,N_12689,N_12536);
nor U13307 (N_13307,N_12673,N_12776);
nor U13308 (N_13308,N_12766,N_12820);
xnor U13309 (N_13309,N_12983,N_12818);
or U13310 (N_13310,N_12586,N_12529);
or U13311 (N_13311,N_12889,N_12500);
and U13312 (N_13312,N_12587,N_12823);
nand U13313 (N_13313,N_12589,N_12672);
nand U13314 (N_13314,N_12959,N_12662);
nand U13315 (N_13315,N_12713,N_12545);
nand U13316 (N_13316,N_12726,N_12771);
and U13317 (N_13317,N_12895,N_12630);
and U13318 (N_13318,N_12841,N_12750);
nand U13319 (N_13319,N_12793,N_12591);
and U13320 (N_13320,N_12822,N_12818);
xnor U13321 (N_13321,N_12880,N_12939);
xor U13322 (N_13322,N_12788,N_12833);
or U13323 (N_13323,N_12888,N_12973);
nor U13324 (N_13324,N_12607,N_12553);
nand U13325 (N_13325,N_12645,N_12647);
and U13326 (N_13326,N_12539,N_12793);
nor U13327 (N_13327,N_12746,N_12865);
or U13328 (N_13328,N_12990,N_12997);
nor U13329 (N_13329,N_12548,N_12692);
or U13330 (N_13330,N_12564,N_12539);
and U13331 (N_13331,N_12905,N_12978);
or U13332 (N_13332,N_12986,N_12959);
xor U13333 (N_13333,N_12711,N_12990);
or U13334 (N_13334,N_12639,N_12962);
nand U13335 (N_13335,N_12738,N_12977);
or U13336 (N_13336,N_12670,N_12619);
or U13337 (N_13337,N_12989,N_12533);
xor U13338 (N_13338,N_12916,N_12691);
and U13339 (N_13339,N_12802,N_12571);
and U13340 (N_13340,N_12763,N_12761);
and U13341 (N_13341,N_12965,N_12780);
nor U13342 (N_13342,N_12700,N_12701);
nand U13343 (N_13343,N_12744,N_12614);
and U13344 (N_13344,N_12623,N_12894);
nor U13345 (N_13345,N_12818,N_12674);
nor U13346 (N_13346,N_12838,N_12783);
nand U13347 (N_13347,N_12545,N_12647);
nor U13348 (N_13348,N_12956,N_12858);
nor U13349 (N_13349,N_12996,N_12686);
nor U13350 (N_13350,N_12552,N_12882);
nor U13351 (N_13351,N_12554,N_12518);
nand U13352 (N_13352,N_12795,N_12870);
or U13353 (N_13353,N_12955,N_12970);
nand U13354 (N_13354,N_12595,N_12931);
and U13355 (N_13355,N_12679,N_12939);
and U13356 (N_13356,N_12654,N_12795);
or U13357 (N_13357,N_12803,N_12549);
xor U13358 (N_13358,N_12583,N_12890);
xor U13359 (N_13359,N_12812,N_12650);
or U13360 (N_13360,N_12956,N_12738);
and U13361 (N_13361,N_12503,N_12569);
or U13362 (N_13362,N_12983,N_12909);
nand U13363 (N_13363,N_12548,N_12641);
or U13364 (N_13364,N_12544,N_12960);
xor U13365 (N_13365,N_12640,N_12904);
or U13366 (N_13366,N_12772,N_12813);
or U13367 (N_13367,N_12877,N_12639);
nor U13368 (N_13368,N_12582,N_12514);
and U13369 (N_13369,N_12681,N_12657);
nand U13370 (N_13370,N_12728,N_12567);
xnor U13371 (N_13371,N_12583,N_12832);
xor U13372 (N_13372,N_12695,N_12923);
xnor U13373 (N_13373,N_12527,N_12873);
and U13374 (N_13374,N_12612,N_12611);
and U13375 (N_13375,N_12741,N_12958);
nand U13376 (N_13376,N_12929,N_12538);
nor U13377 (N_13377,N_12559,N_12983);
and U13378 (N_13378,N_12617,N_12650);
nor U13379 (N_13379,N_12766,N_12852);
nand U13380 (N_13380,N_12610,N_12674);
nor U13381 (N_13381,N_12618,N_12754);
nand U13382 (N_13382,N_12700,N_12835);
nand U13383 (N_13383,N_12608,N_12658);
or U13384 (N_13384,N_12672,N_12568);
or U13385 (N_13385,N_12988,N_12733);
nand U13386 (N_13386,N_12632,N_12761);
or U13387 (N_13387,N_12646,N_12504);
nor U13388 (N_13388,N_12543,N_12521);
xnor U13389 (N_13389,N_12618,N_12639);
and U13390 (N_13390,N_12951,N_12777);
xor U13391 (N_13391,N_12879,N_12885);
nand U13392 (N_13392,N_12832,N_12815);
or U13393 (N_13393,N_12513,N_12895);
and U13394 (N_13394,N_12603,N_12963);
xor U13395 (N_13395,N_12679,N_12909);
nand U13396 (N_13396,N_12882,N_12517);
xnor U13397 (N_13397,N_12632,N_12666);
and U13398 (N_13398,N_12564,N_12718);
and U13399 (N_13399,N_12790,N_12822);
and U13400 (N_13400,N_12901,N_12722);
xnor U13401 (N_13401,N_12785,N_12726);
or U13402 (N_13402,N_12953,N_12690);
or U13403 (N_13403,N_12864,N_12729);
nand U13404 (N_13404,N_12717,N_12978);
and U13405 (N_13405,N_12511,N_12876);
nor U13406 (N_13406,N_12542,N_12576);
or U13407 (N_13407,N_12961,N_12595);
nor U13408 (N_13408,N_12923,N_12564);
and U13409 (N_13409,N_12679,N_12595);
nor U13410 (N_13410,N_12870,N_12987);
nor U13411 (N_13411,N_12800,N_12804);
nor U13412 (N_13412,N_12896,N_12798);
nand U13413 (N_13413,N_12683,N_12917);
nor U13414 (N_13414,N_12628,N_12563);
nand U13415 (N_13415,N_12686,N_12568);
xnor U13416 (N_13416,N_12921,N_12689);
and U13417 (N_13417,N_12599,N_12976);
xor U13418 (N_13418,N_12987,N_12993);
nand U13419 (N_13419,N_12728,N_12797);
nand U13420 (N_13420,N_12996,N_12578);
nand U13421 (N_13421,N_12925,N_12719);
nand U13422 (N_13422,N_12907,N_12784);
xor U13423 (N_13423,N_12704,N_12711);
nand U13424 (N_13424,N_12576,N_12606);
nor U13425 (N_13425,N_12624,N_12725);
xnor U13426 (N_13426,N_12790,N_12583);
nand U13427 (N_13427,N_12924,N_12987);
and U13428 (N_13428,N_12576,N_12724);
nand U13429 (N_13429,N_12636,N_12889);
or U13430 (N_13430,N_12800,N_12664);
and U13431 (N_13431,N_12778,N_12925);
or U13432 (N_13432,N_12962,N_12668);
nor U13433 (N_13433,N_12779,N_12966);
nor U13434 (N_13434,N_12645,N_12971);
and U13435 (N_13435,N_12728,N_12875);
nor U13436 (N_13436,N_12783,N_12575);
and U13437 (N_13437,N_12715,N_12627);
or U13438 (N_13438,N_12916,N_12589);
and U13439 (N_13439,N_12870,N_12563);
nand U13440 (N_13440,N_12957,N_12572);
nand U13441 (N_13441,N_12857,N_12845);
and U13442 (N_13442,N_12750,N_12946);
or U13443 (N_13443,N_12959,N_12943);
nand U13444 (N_13444,N_12646,N_12989);
xor U13445 (N_13445,N_12716,N_12749);
nand U13446 (N_13446,N_12921,N_12823);
nor U13447 (N_13447,N_12858,N_12993);
nor U13448 (N_13448,N_12697,N_12844);
or U13449 (N_13449,N_12793,N_12828);
and U13450 (N_13450,N_12844,N_12957);
xor U13451 (N_13451,N_12716,N_12661);
xor U13452 (N_13452,N_12709,N_12583);
or U13453 (N_13453,N_12509,N_12511);
and U13454 (N_13454,N_12998,N_12759);
xor U13455 (N_13455,N_12701,N_12638);
or U13456 (N_13456,N_12785,N_12704);
nor U13457 (N_13457,N_12679,N_12932);
and U13458 (N_13458,N_12526,N_12850);
or U13459 (N_13459,N_12590,N_12724);
nor U13460 (N_13460,N_12853,N_12907);
and U13461 (N_13461,N_12541,N_12669);
xor U13462 (N_13462,N_12937,N_12813);
nor U13463 (N_13463,N_12726,N_12927);
or U13464 (N_13464,N_12702,N_12640);
or U13465 (N_13465,N_12583,N_12593);
nor U13466 (N_13466,N_12980,N_12783);
xnor U13467 (N_13467,N_12581,N_12863);
xnor U13468 (N_13468,N_12950,N_12712);
or U13469 (N_13469,N_12697,N_12754);
xnor U13470 (N_13470,N_12922,N_12776);
and U13471 (N_13471,N_12733,N_12631);
xnor U13472 (N_13472,N_12974,N_12662);
or U13473 (N_13473,N_12595,N_12501);
nand U13474 (N_13474,N_12831,N_12994);
nand U13475 (N_13475,N_12704,N_12600);
nor U13476 (N_13476,N_12983,N_12585);
or U13477 (N_13477,N_12753,N_12807);
nand U13478 (N_13478,N_12659,N_12808);
and U13479 (N_13479,N_12733,N_12806);
and U13480 (N_13480,N_12956,N_12905);
and U13481 (N_13481,N_12754,N_12792);
nor U13482 (N_13482,N_12728,N_12685);
and U13483 (N_13483,N_12969,N_12672);
nand U13484 (N_13484,N_12501,N_12644);
and U13485 (N_13485,N_12881,N_12688);
nand U13486 (N_13486,N_12652,N_12511);
nor U13487 (N_13487,N_12953,N_12659);
nand U13488 (N_13488,N_12972,N_12779);
or U13489 (N_13489,N_12847,N_12897);
nand U13490 (N_13490,N_12891,N_12707);
nand U13491 (N_13491,N_12665,N_12781);
nand U13492 (N_13492,N_12590,N_12937);
xor U13493 (N_13493,N_12660,N_12746);
xnor U13494 (N_13494,N_12736,N_12987);
and U13495 (N_13495,N_12518,N_12739);
nand U13496 (N_13496,N_12576,N_12693);
nor U13497 (N_13497,N_12703,N_12787);
nor U13498 (N_13498,N_12597,N_12552);
nor U13499 (N_13499,N_12851,N_12685);
and U13500 (N_13500,N_13106,N_13147);
nand U13501 (N_13501,N_13341,N_13288);
xnor U13502 (N_13502,N_13200,N_13324);
or U13503 (N_13503,N_13107,N_13226);
and U13504 (N_13504,N_13054,N_13008);
or U13505 (N_13505,N_13334,N_13067);
and U13506 (N_13506,N_13385,N_13303);
nor U13507 (N_13507,N_13449,N_13378);
or U13508 (N_13508,N_13379,N_13150);
nand U13509 (N_13509,N_13279,N_13464);
nand U13510 (N_13510,N_13138,N_13495);
nor U13511 (N_13511,N_13352,N_13422);
nand U13512 (N_13512,N_13483,N_13048);
nand U13513 (N_13513,N_13477,N_13498);
nand U13514 (N_13514,N_13451,N_13316);
or U13515 (N_13515,N_13083,N_13411);
nand U13516 (N_13516,N_13125,N_13033);
xor U13517 (N_13517,N_13466,N_13036);
and U13518 (N_13518,N_13425,N_13227);
nand U13519 (N_13519,N_13358,N_13052);
nand U13520 (N_13520,N_13260,N_13369);
and U13521 (N_13521,N_13374,N_13395);
and U13522 (N_13522,N_13120,N_13259);
nor U13523 (N_13523,N_13264,N_13305);
nand U13524 (N_13524,N_13326,N_13224);
nand U13525 (N_13525,N_13338,N_13016);
xor U13526 (N_13526,N_13251,N_13021);
xor U13527 (N_13527,N_13127,N_13100);
nand U13528 (N_13528,N_13415,N_13160);
nor U13529 (N_13529,N_13213,N_13429);
and U13530 (N_13530,N_13295,N_13207);
and U13531 (N_13531,N_13486,N_13382);
xnor U13532 (N_13532,N_13297,N_13433);
nand U13533 (N_13533,N_13491,N_13062);
xnor U13534 (N_13534,N_13030,N_13301);
or U13535 (N_13535,N_13056,N_13381);
nor U13536 (N_13536,N_13257,N_13255);
and U13537 (N_13537,N_13427,N_13093);
and U13538 (N_13538,N_13191,N_13313);
nand U13539 (N_13539,N_13091,N_13244);
or U13540 (N_13540,N_13402,N_13468);
or U13541 (N_13541,N_13201,N_13342);
nor U13542 (N_13542,N_13212,N_13102);
nor U13543 (N_13543,N_13024,N_13470);
or U13544 (N_13544,N_13068,N_13077);
and U13545 (N_13545,N_13168,N_13026);
xor U13546 (N_13546,N_13157,N_13265);
and U13547 (N_13547,N_13070,N_13423);
nor U13548 (N_13548,N_13443,N_13139);
nand U13549 (N_13549,N_13489,N_13481);
or U13550 (N_13550,N_13073,N_13171);
and U13551 (N_13551,N_13214,N_13431);
xor U13552 (N_13552,N_13234,N_13285);
nor U13553 (N_13553,N_13004,N_13323);
and U13554 (N_13554,N_13393,N_13453);
or U13555 (N_13555,N_13084,N_13447);
and U13556 (N_13556,N_13497,N_13045);
xor U13557 (N_13557,N_13430,N_13105);
nand U13558 (N_13558,N_13266,N_13432);
or U13559 (N_13559,N_13267,N_13383);
and U13560 (N_13560,N_13315,N_13019);
or U13561 (N_13561,N_13010,N_13001);
xnor U13562 (N_13562,N_13081,N_13158);
or U13563 (N_13563,N_13050,N_13069);
or U13564 (N_13564,N_13245,N_13319);
and U13565 (N_13565,N_13335,N_13231);
xnor U13566 (N_13566,N_13198,N_13141);
nor U13567 (N_13567,N_13273,N_13480);
nand U13568 (N_13568,N_13118,N_13347);
and U13569 (N_13569,N_13462,N_13331);
nor U13570 (N_13570,N_13282,N_13325);
nand U13571 (N_13571,N_13327,N_13344);
and U13572 (N_13572,N_13185,N_13205);
and U13573 (N_13573,N_13005,N_13365);
and U13574 (N_13574,N_13405,N_13277);
xor U13575 (N_13575,N_13299,N_13209);
xor U13576 (N_13576,N_13322,N_13275);
nor U13577 (N_13577,N_13418,N_13044);
xnor U13578 (N_13578,N_13167,N_13129);
and U13579 (N_13579,N_13281,N_13444);
nand U13580 (N_13580,N_13496,N_13330);
xnor U13581 (N_13581,N_13041,N_13009);
nor U13582 (N_13582,N_13333,N_13146);
nor U13583 (N_13583,N_13293,N_13302);
nor U13584 (N_13584,N_13484,N_13228);
and U13585 (N_13585,N_13237,N_13471);
nor U13586 (N_13586,N_13190,N_13003);
nand U13587 (N_13587,N_13194,N_13308);
and U13588 (N_13588,N_13442,N_13271);
and U13589 (N_13589,N_13022,N_13294);
and U13590 (N_13590,N_13252,N_13397);
nor U13591 (N_13591,N_13448,N_13454);
and U13592 (N_13592,N_13391,N_13363);
and U13593 (N_13593,N_13356,N_13473);
xor U13594 (N_13594,N_13494,N_13222);
or U13595 (N_13595,N_13398,N_13066);
xor U13596 (N_13596,N_13388,N_13350);
and U13597 (N_13597,N_13246,N_13371);
and U13598 (N_13598,N_13206,N_13403);
and U13599 (N_13599,N_13248,N_13040);
xor U13600 (N_13600,N_13186,N_13258);
xnor U13601 (N_13601,N_13204,N_13140);
xor U13602 (N_13602,N_13332,N_13085);
or U13603 (N_13603,N_13469,N_13002);
nand U13604 (N_13604,N_13110,N_13283);
or U13605 (N_13605,N_13208,N_13057);
xor U13606 (N_13606,N_13154,N_13460);
and U13607 (N_13607,N_13309,N_13181);
or U13608 (N_13608,N_13372,N_13413);
or U13609 (N_13609,N_13328,N_13351);
nor U13610 (N_13610,N_13475,N_13098);
xor U13611 (N_13611,N_13452,N_13268);
and U13612 (N_13612,N_13360,N_13317);
and U13613 (N_13613,N_13321,N_13135);
nand U13614 (N_13614,N_13131,N_13375);
nand U13615 (N_13615,N_13238,N_13235);
or U13616 (N_13616,N_13012,N_13396);
xor U13617 (N_13617,N_13132,N_13488);
xnor U13618 (N_13618,N_13148,N_13380);
xnor U13619 (N_13619,N_13446,N_13339);
and U13620 (N_13620,N_13249,N_13095);
and U13621 (N_13621,N_13126,N_13182);
nor U13622 (N_13622,N_13063,N_13337);
and U13623 (N_13623,N_13242,N_13278);
nand U13624 (N_13624,N_13035,N_13343);
or U13625 (N_13625,N_13287,N_13203);
nor U13626 (N_13626,N_13192,N_13291);
xnor U13627 (N_13627,N_13384,N_13220);
nand U13628 (N_13628,N_13134,N_13362);
and U13629 (N_13629,N_13434,N_13074);
or U13630 (N_13630,N_13230,N_13058);
or U13631 (N_13631,N_13346,N_13053);
or U13632 (N_13632,N_13112,N_13218);
or U13633 (N_13633,N_13221,N_13031);
nand U13634 (N_13634,N_13136,N_13162);
or U13635 (N_13635,N_13113,N_13478);
nand U13636 (N_13636,N_13086,N_13312);
xor U13637 (N_13637,N_13304,N_13320);
xor U13638 (N_13638,N_13013,N_13104);
nand U13639 (N_13639,N_13065,N_13366);
and U13640 (N_13640,N_13006,N_13314);
nor U13641 (N_13641,N_13361,N_13092);
or U13642 (N_13642,N_13000,N_13094);
nand U13643 (N_13643,N_13306,N_13175);
nor U13644 (N_13644,N_13261,N_13336);
or U13645 (N_13645,N_13472,N_13143);
nor U13646 (N_13646,N_13087,N_13329);
xnor U13647 (N_13647,N_13456,N_13310);
and U13648 (N_13648,N_13210,N_13133);
nand U13649 (N_13649,N_13490,N_13420);
and U13650 (N_13650,N_13159,N_13286);
nor U13651 (N_13651,N_13438,N_13239);
nand U13652 (N_13652,N_13049,N_13280);
or U13653 (N_13653,N_13137,N_13399);
nand U13654 (N_13654,N_13025,N_13276);
xnor U13655 (N_13655,N_13169,N_13130);
or U13656 (N_13656,N_13170,N_13368);
and U13657 (N_13657,N_13233,N_13038);
nand U13658 (N_13658,N_13055,N_13428);
and U13659 (N_13659,N_13082,N_13116);
nor U13660 (N_13660,N_13284,N_13034);
or U13661 (N_13661,N_13436,N_13492);
nor U13662 (N_13662,N_13177,N_13060);
xor U13663 (N_13663,N_13075,N_13482);
xnor U13664 (N_13664,N_13243,N_13188);
nand U13665 (N_13665,N_13318,N_13270);
or U13666 (N_13666,N_13476,N_13401);
nor U13667 (N_13667,N_13046,N_13172);
nor U13668 (N_13668,N_13029,N_13364);
and U13669 (N_13669,N_13232,N_13079);
and U13670 (N_13670,N_13345,N_13421);
or U13671 (N_13671,N_13197,N_13439);
or U13672 (N_13672,N_13011,N_13023);
nand U13673 (N_13673,N_13144,N_13414);
nor U13674 (N_13674,N_13290,N_13459);
nor U13675 (N_13675,N_13410,N_13254);
nor U13676 (N_13676,N_13196,N_13155);
nor U13677 (N_13677,N_13020,N_13153);
nor U13678 (N_13678,N_13457,N_13419);
nand U13679 (N_13679,N_13152,N_13078);
nor U13680 (N_13680,N_13216,N_13461);
xor U13681 (N_13681,N_13219,N_13376);
xor U13682 (N_13682,N_13353,N_13247);
nand U13683 (N_13683,N_13357,N_13406);
or U13684 (N_13684,N_13463,N_13064);
nor U13685 (N_13685,N_13349,N_13250);
xnor U13686 (N_13686,N_13193,N_13354);
nor U13687 (N_13687,N_13416,N_13103);
nor U13688 (N_13688,N_13474,N_13014);
and U13689 (N_13689,N_13435,N_13455);
and U13690 (N_13690,N_13088,N_13184);
nand U13691 (N_13691,N_13311,N_13047);
and U13692 (N_13692,N_13007,N_13142);
or U13693 (N_13693,N_13386,N_13032);
and U13694 (N_13694,N_13289,N_13018);
xor U13695 (N_13695,N_13412,N_13487);
nand U13696 (N_13696,N_13307,N_13465);
xnor U13697 (N_13697,N_13042,N_13109);
nand U13698 (N_13698,N_13298,N_13467);
xor U13699 (N_13699,N_13479,N_13404);
nand U13700 (N_13700,N_13180,N_13370);
and U13701 (N_13701,N_13389,N_13485);
nor U13702 (N_13702,N_13176,N_13187);
nand U13703 (N_13703,N_13199,N_13156);
nand U13704 (N_13704,N_13348,N_13458);
xor U13705 (N_13705,N_13076,N_13121);
xnor U13706 (N_13706,N_13061,N_13355);
or U13707 (N_13707,N_13367,N_13256);
or U13708 (N_13708,N_13359,N_13164);
nor U13709 (N_13709,N_13114,N_13437);
and U13710 (N_13710,N_13373,N_13450);
or U13711 (N_13711,N_13417,N_13394);
xor U13712 (N_13712,N_13409,N_13499);
xor U13713 (N_13713,N_13128,N_13089);
xor U13714 (N_13714,N_13202,N_13173);
xor U13715 (N_13715,N_13183,N_13390);
nor U13716 (N_13716,N_13392,N_13225);
xor U13717 (N_13717,N_13090,N_13178);
xor U13718 (N_13718,N_13099,N_13240);
nor U13719 (N_13719,N_13215,N_13493);
or U13720 (N_13720,N_13424,N_13229);
xnor U13721 (N_13721,N_13151,N_13124);
and U13722 (N_13722,N_13039,N_13195);
nor U13723 (N_13723,N_13017,N_13387);
or U13724 (N_13724,N_13377,N_13441);
xnor U13725 (N_13725,N_13051,N_13269);
nand U13726 (N_13726,N_13445,N_13189);
nor U13727 (N_13727,N_13272,N_13340);
nand U13728 (N_13728,N_13096,N_13408);
nand U13729 (N_13729,N_13211,N_13292);
nor U13730 (N_13730,N_13262,N_13300);
nand U13731 (N_13731,N_13122,N_13080);
and U13732 (N_13732,N_13145,N_13071);
and U13733 (N_13733,N_13440,N_13400);
nor U13734 (N_13734,N_13015,N_13111);
or U13735 (N_13735,N_13296,N_13097);
nor U13736 (N_13736,N_13123,N_13149);
or U13737 (N_13737,N_13174,N_13179);
nand U13738 (N_13738,N_13101,N_13253);
nand U13739 (N_13739,N_13274,N_13119);
or U13740 (N_13740,N_13072,N_13028);
or U13741 (N_13741,N_13163,N_13043);
nand U13742 (N_13742,N_13165,N_13059);
or U13743 (N_13743,N_13027,N_13037);
nor U13744 (N_13744,N_13108,N_13223);
nand U13745 (N_13745,N_13115,N_13161);
or U13746 (N_13746,N_13166,N_13117);
and U13747 (N_13747,N_13407,N_13236);
or U13748 (N_13748,N_13241,N_13217);
xnor U13749 (N_13749,N_13426,N_13263);
and U13750 (N_13750,N_13100,N_13013);
xnor U13751 (N_13751,N_13389,N_13176);
nand U13752 (N_13752,N_13342,N_13332);
xnor U13753 (N_13753,N_13442,N_13053);
nor U13754 (N_13754,N_13216,N_13350);
and U13755 (N_13755,N_13418,N_13426);
and U13756 (N_13756,N_13107,N_13049);
nor U13757 (N_13757,N_13163,N_13494);
or U13758 (N_13758,N_13211,N_13411);
and U13759 (N_13759,N_13209,N_13257);
and U13760 (N_13760,N_13072,N_13415);
nor U13761 (N_13761,N_13389,N_13310);
nor U13762 (N_13762,N_13291,N_13135);
nand U13763 (N_13763,N_13291,N_13229);
and U13764 (N_13764,N_13226,N_13251);
nand U13765 (N_13765,N_13314,N_13347);
nor U13766 (N_13766,N_13143,N_13222);
nor U13767 (N_13767,N_13207,N_13098);
xor U13768 (N_13768,N_13087,N_13347);
or U13769 (N_13769,N_13403,N_13109);
xnor U13770 (N_13770,N_13274,N_13423);
or U13771 (N_13771,N_13412,N_13140);
xor U13772 (N_13772,N_13437,N_13166);
xor U13773 (N_13773,N_13318,N_13298);
xnor U13774 (N_13774,N_13183,N_13179);
nor U13775 (N_13775,N_13191,N_13267);
nand U13776 (N_13776,N_13064,N_13172);
nor U13777 (N_13777,N_13443,N_13168);
or U13778 (N_13778,N_13155,N_13124);
or U13779 (N_13779,N_13398,N_13101);
or U13780 (N_13780,N_13237,N_13437);
or U13781 (N_13781,N_13406,N_13211);
nor U13782 (N_13782,N_13367,N_13313);
nand U13783 (N_13783,N_13152,N_13410);
nand U13784 (N_13784,N_13027,N_13314);
and U13785 (N_13785,N_13201,N_13034);
nor U13786 (N_13786,N_13116,N_13303);
or U13787 (N_13787,N_13138,N_13122);
or U13788 (N_13788,N_13379,N_13064);
nand U13789 (N_13789,N_13198,N_13258);
nand U13790 (N_13790,N_13366,N_13268);
and U13791 (N_13791,N_13129,N_13346);
nand U13792 (N_13792,N_13470,N_13372);
nand U13793 (N_13793,N_13054,N_13478);
nor U13794 (N_13794,N_13485,N_13463);
nor U13795 (N_13795,N_13251,N_13266);
nor U13796 (N_13796,N_13320,N_13393);
nand U13797 (N_13797,N_13023,N_13300);
nor U13798 (N_13798,N_13245,N_13198);
xor U13799 (N_13799,N_13008,N_13156);
nand U13800 (N_13800,N_13151,N_13234);
and U13801 (N_13801,N_13073,N_13018);
nand U13802 (N_13802,N_13205,N_13154);
nor U13803 (N_13803,N_13409,N_13046);
or U13804 (N_13804,N_13303,N_13117);
xnor U13805 (N_13805,N_13467,N_13171);
nor U13806 (N_13806,N_13393,N_13395);
nor U13807 (N_13807,N_13185,N_13224);
xor U13808 (N_13808,N_13209,N_13369);
nand U13809 (N_13809,N_13338,N_13305);
nor U13810 (N_13810,N_13481,N_13412);
xor U13811 (N_13811,N_13338,N_13105);
nand U13812 (N_13812,N_13479,N_13079);
xnor U13813 (N_13813,N_13077,N_13421);
and U13814 (N_13814,N_13045,N_13442);
nor U13815 (N_13815,N_13147,N_13330);
xor U13816 (N_13816,N_13024,N_13390);
nand U13817 (N_13817,N_13206,N_13202);
nor U13818 (N_13818,N_13476,N_13029);
and U13819 (N_13819,N_13193,N_13163);
or U13820 (N_13820,N_13184,N_13180);
or U13821 (N_13821,N_13215,N_13216);
xor U13822 (N_13822,N_13218,N_13332);
or U13823 (N_13823,N_13353,N_13462);
or U13824 (N_13824,N_13137,N_13111);
and U13825 (N_13825,N_13020,N_13474);
xnor U13826 (N_13826,N_13215,N_13280);
or U13827 (N_13827,N_13417,N_13085);
xor U13828 (N_13828,N_13341,N_13316);
and U13829 (N_13829,N_13339,N_13146);
nor U13830 (N_13830,N_13265,N_13200);
nor U13831 (N_13831,N_13422,N_13364);
nor U13832 (N_13832,N_13147,N_13021);
and U13833 (N_13833,N_13241,N_13353);
nor U13834 (N_13834,N_13198,N_13347);
xnor U13835 (N_13835,N_13110,N_13123);
nor U13836 (N_13836,N_13400,N_13192);
nor U13837 (N_13837,N_13233,N_13351);
nor U13838 (N_13838,N_13384,N_13276);
and U13839 (N_13839,N_13458,N_13387);
and U13840 (N_13840,N_13098,N_13392);
or U13841 (N_13841,N_13188,N_13321);
nor U13842 (N_13842,N_13242,N_13411);
or U13843 (N_13843,N_13029,N_13452);
nand U13844 (N_13844,N_13094,N_13355);
and U13845 (N_13845,N_13439,N_13269);
nand U13846 (N_13846,N_13077,N_13494);
nand U13847 (N_13847,N_13114,N_13228);
xor U13848 (N_13848,N_13264,N_13335);
and U13849 (N_13849,N_13238,N_13472);
and U13850 (N_13850,N_13337,N_13194);
xor U13851 (N_13851,N_13273,N_13274);
or U13852 (N_13852,N_13477,N_13027);
nor U13853 (N_13853,N_13040,N_13411);
nand U13854 (N_13854,N_13125,N_13408);
or U13855 (N_13855,N_13496,N_13281);
or U13856 (N_13856,N_13301,N_13124);
and U13857 (N_13857,N_13203,N_13011);
nor U13858 (N_13858,N_13371,N_13382);
xor U13859 (N_13859,N_13492,N_13265);
nand U13860 (N_13860,N_13437,N_13496);
nor U13861 (N_13861,N_13009,N_13183);
nor U13862 (N_13862,N_13100,N_13252);
or U13863 (N_13863,N_13099,N_13268);
nand U13864 (N_13864,N_13195,N_13232);
nand U13865 (N_13865,N_13379,N_13109);
nor U13866 (N_13866,N_13447,N_13366);
or U13867 (N_13867,N_13090,N_13140);
or U13868 (N_13868,N_13395,N_13256);
or U13869 (N_13869,N_13051,N_13401);
nand U13870 (N_13870,N_13266,N_13278);
nand U13871 (N_13871,N_13083,N_13460);
nand U13872 (N_13872,N_13369,N_13323);
nand U13873 (N_13873,N_13441,N_13145);
nor U13874 (N_13874,N_13460,N_13358);
nand U13875 (N_13875,N_13397,N_13462);
nor U13876 (N_13876,N_13320,N_13300);
and U13877 (N_13877,N_13171,N_13334);
nand U13878 (N_13878,N_13411,N_13200);
nor U13879 (N_13879,N_13330,N_13131);
nor U13880 (N_13880,N_13413,N_13010);
or U13881 (N_13881,N_13187,N_13461);
and U13882 (N_13882,N_13276,N_13182);
or U13883 (N_13883,N_13453,N_13233);
and U13884 (N_13884,N_13478,N_13190);
nand U13885 (N_13885,N_13349,N_13432);
xnor U13886 (N_13886,N_13399,N_13391);
and U13887 (N_13887,N_13139,N_13425);
nor U13888 (N_13888,N_13310,N_13464);
or U13889 (N_13889,N_13236,N_13334);
nand U13890 (N_13890,N_13429,N_13326);
nor U13891 (N_13891,N_13108,N_13061);
or U13892 (N_13892,N_13217,N_13356);
nor U13893 (N_13893,N_13125,N_13166);
and U13894 (N_13894,N_13490,N_13200);
nor U13895 (N_13895,N_13149,N_13270);
nand U13896 (N_13896,N_13171,N_13354);
and U13897 (N_13897,N_13132,N_13495);
and U13898 (N_13898,N_13043,N_13010);
nor U13899 (N_13899,N_13092,N_13320);
or U13900 (N_13900,N_13304,N_13331);
and U13901 (N_13901,N_13089,N_13044);
nor U13902 (N_13902,N_13465,N_13207);
xor U13903 (N_13903,N_13173,N_13428);
or U13904 (N_13904,N_13262,N_13165);
or U13905 (N_13905,N_13411,N_13491);
nor U13906 (N_13906,N_13156,N_13288);
xnor U13907 (N_13907,N_13444,N_13453);
or U13908 (N_13908,N_13276,N_13415);
xnor U13909 (N_13909,N_13394,N_13123);
xor U13910 (N_13910,N_13174,N_13135);
or U13911 (N_13911,N_13003,N_13474);
or U13912 (N_13912,N_13425,N_13039);
and U13913 (N_13913,N_13291,N_13236);
or U13914 (N_13914,N_13284,N_13222);
nor U13915 (N_13915,N_13469,N_13202);
or U13916 (N_13916,N_13148,N_13124);
and U13917 (N_13917,N_13283,N_13159);
nand U13918 (N_13918,N_13314,N_13001);
and U13919 (N_13919,N_13365,N_13043);
or U13920 (N_13920,N_13149,N_13020);
nor U13921 (N_13921,N_13295,N_13241);
xor U13922 (N_13922,N_13118,N_13404);
or U13923 (N_13923,N_13150,N_13405);
and U13924 (N_13924,N_13258,N_13450);
or U13925 (N_13925,N_13151,N_13227);
or U13926 (N_13926,N_13157,N_13173);
nor U13927 (N_13927,N_13467,N_13154);
nor U13928 (N_13928,N_13189,N_13475);
or U13929 (N_13929,N_13482,N_13473);
and U13930 (N_13930,N_13191,N_13118);
and U13931 (N_13931,N_13287,N_13212);
nor U13932 (N_13932,N_13408,N_13376);
nor U13933 (N_13933,N_13211,N_13403);
nand U13934 (N_13934,N_13092,N_13201);
and U13935 (N_13935,N_13313,N_13251);
nor U13936 (N_13936,N_13434,N_13389);
nor U13937 (N_13937,N_13326,N_13267);
nand U13938 (N_13938,N_13280,N_13411);
and U13939 (N_13939,N_13425,N_13281);
or U13940 (N_13940,N_13444,N_13098);
xor U13941 (N_13941,N_13196,N_13191);
or U13942 (N_13942,N_13273,N_13105);
or U13943 (N_13943,N_13382,N_13073);
or U13944 (N_13944,N_13187,N_13172);
and U13945 (N_13945,N_13123,N_13091);
nor U13946 (N_13946,N_13325,N_13249);
xnor U13947 (N_13947,N_13096,N_13090);
xnor U13948 (N_13948,N_13468,N_13033);
or U13949 (N_13949,N_13457,N_13194);
and U13950 (N_13950,N_13485,N_13209);
nor U13951 (N_13951,N_13246,N_13283);
nand U13952 (N_13952,N_13356,N_13197);
nand U13953 (N_13953,N_13172,N_13388);
nand U13954 (N_13954,N_13125,N_13152);
nand U13955 (N_13955,N_13318,N_13437);
nand U13956 (N_13956,N_13158,N_13101);
xnor U13957 (N_13957,N_13388,N_13026);
and U13958 (N_13958,N_13262,N_13221);
nor U13959 (N_13959,N_13057,N_13059);
and U13960 (N_13960,N_13312,N_13157);
nor U13961 (N_13961,N_13112,N_13288);
or U13962 (N_13962,N_13015,N_13190);
xor U13963 (N_13963,N_13065,N_13454);
or U13964 (N_13964,N_13348,N_13159);
or U13965 (N_13965,N_13456,N_13357);
and U13966 (N_13966,N_13491,N_13222);
nand U13967 (N_13967,N_13160,N_13090);
nor U13968 (N_13968,N_13284,N_13463);
or U13969 (N_13969,N_13283,N_13187);
xnor U13970 (N_13970,N_13022,N_13363);
xor U13971 (N_13971,N_13120,N_13049);
and U13972 (N_13972,N_13413,N_13470);
nor U13973 (N_13973,N_13201,N_13402);
xor U13974 (N_13974,N_13451,N_13109);
or U13975 (N_13975,N_13082,N_13150);
nor U13976 (N_13976,N_13453,N_13495);
nand U13977 (N_13977,N_13103,N_13330);
nor U13978 (N_13978,N_13076,N_13296);
nor U13979 (N_13979,N_13200,N_13388);
or U13980 (N_13980,N_13138,N_13221);
nor U13981 (N_13981,N_13412,N_13032);
or U13982 (N_13982,N_13137,N_13208);
nand U13983 (N_13983,N_13398,N_13205);
or U13984 (N_13984,N_13031,N_13125);
or U13985 (N_13985,N_13170,N_13456);
xor U13986 (N_13986,N_13368,N_13226);
nor U13987 (N_13987,N_13274,N_13308);
and U13988 (N_13988,N_13257,N_13320);
xor U13989 (N_13989,N_13083,N_13453);
xnor U13990 (N_13990,N_13098,N_13295);
nand U13991 (N_13991,N_13071,N_13257);
nand U13992 (N_13992,N_13005,N_13086);
or U13993 (N_13993,N_13124,N_13020);
nand U13994 (N_13994,N_13096,N_13273);
nor U13995 (N_13995,N_13394,N_13035);
or U13996 (N_13996,N_13195,N_13134);
nand U13997 (N_13997,N_13065,N_13188);
xor U13998 (N_13998,N_13287,N_13130);
xnor U13999 (N_13999,N_13452,N_13461);
xor U14000 (N_14000,N_13944,N_13616);
and U14001 (N_14001,N_13754,N_13620);
or U14002 (N_14002,N_13538,N_13781);
nand U14003 (N_14003,N_13871,N_13810);
or U14004 (N_14004,N_13572,N_13615);
nand U14005 (N_14005,N_13654,N_13518);
nor U14006 (N_14006,N_13599,N_13551);
nor U14007 (N_14007,N_13909,N_13792);
xnor U14008 (N_14008,N_13914,N_13831);
or U14009 (N_14009,N_13829,N_13541);
xor U14010 (N_14010,N_13861,N_13507);
or U14011 (N_14011,N_13711,N_13648);
nand U14012 (N_14012,N_13812,N_13593);
and U14013 (N_14013,N_13546,N_13913);
nor U14014 (N_14014,N_13783,N_13664);
nor U14015 (N_14015,N_13626,N_13922);
xnor U14016 (N_14016,N_13882,N_13935);
and U14017 (N_14017,N_13787,N_13624);
xor U14018 (N_14018,N_13556,N_13553);
xnor U14019 (N_14019,N_13960,N_13953);
and U14020 (N_14020,N_13930,N_13618);
and U14021 (N_14021,N_13919,N_13672);
and U14022 (N_14022,N_13799,N_13999);
nor U14023 (N_14023,N_13660,N_13657);
xnor U14024 (N_14024,N_13977,N_13817);
and U14025 (N_14025,N_13682,N_13506);
xnor U14026 (N_14026,N_13993,N_13929);
or U14027 (N_14027,N_13696,N_13517);
xnor U14028 (N_14028,N_13559,N_13653);
or U14029 (N_14029,N_13955,N_13803);
nand U14030 (N_14030,N_13918,N_13877);
xnor U14031 (N_14031,N_13681,N_13834);
nand U14032 (N_14032,N_13590,N_13673);
and U14033 (N_14033,N_13786,N_13661);
nor U14034 (N_14034,N_13649,N_13500);
nand U14035 (N_14035,N_13899,N_13561);
xor U14036 (N_14036,N_13560,N_13602);
and U14037 (N_14037,N_13818,N_13571);
nand U14038 (N_14038,N_13569,N_13804);
nand U14039 (N_14039,N_13723,N_13897);
or U14040 (N_14040,N_13652,N_13731);
nand U14041 (N_14041,N_13874,N_13585);
nor U14042 (N_14042,N_13703,N_13575);
and U14043 (N_14043,N_13509,N_13766);
nor U14044 (N_14044,N_13634,N_13980);
and U14045 (N_14045,N_13837,N_13565);
or U14046 (N_14046,N_13570,N_13784);
and U14047 (N_14047,N_13827,N_13925);
and U14048 (N_14048,N_13677,N_13869);
or U14049 (N_14049,N_13687,N_13636);
xor U14050 (N_14050,N_13957,N_13535);
nor U14051 (N_14051,N_13520,N_13676);
nor U14052 (N_14052,N_13939,N_13764);
and U14053 (N_14053,N_13592,N_13641);
and U14054 (N_14054,N_13646,N_13921);
xor U14055 (N_14055,N_13911,N_13916);
nor U14056 (N_14056,N_13519,N_13666);
nor U14057 (N_14057,N_13611,N_13849);
or U14058 (N_14058,N_13850,N_13749);
nand U14059 (N_14059,N_13512,N_13979);
xnor U14060 (N_14060,N_13567,N_13639);
nor U14061 (N_14061,N_13968,N_13958);
and U14062 (N_14062,N_13508,N_13580);
nor U14063 (N_14063,N_13531,N_13997);
xor U14064 (N_14064,N_13986,N_13795);
nor U14065 (N_14065,N_13751,N_13765);
nor U14066 (N_14066,N_13767,N_13617);
nor U14067 (N_14067,N_13876,N_13791);
or U14068 (N_14068,N_13932,N_13926);
nand U14069 (N_14069,N_13898,N_13655);
nor U14070 (N_14070,N_13591,N_13527);
and U14071 (N_14071,N_13726,N_13858);
nor U14072 (N_14072,N_13706,N_13972);
and U14073 (N_14073,N_13836,N_13776);
nand U14074 (N_14074,N_13699,N_13890);
or U14075 (N_14075,N_13642,N_13978);
nor U14076 (N_14076,N_13524,N_13934);
or U14077 (N_14077,N_13772,N_13540);
nor U14078 (N_14078,N_13697,N_13713);
nor U14079 (N_14079,N_13905,N_13698);
xnor U14080 (N_14080,N_13564,N_13838);
nor U14081 (N_14081,N_13847,N_13940);
nand U14082 (N_14082,N_13788,N_13854);
or U14083 (N_14083,N_13712,N_13920);
nand U14084 (N_14084,N_13862,N_13917);
xnor U14085 (N_14085,N_13832,N_13963);
and U14086 (N_14086,N_13878,N_13965);
nor U14087 (N_14087,N_13895,N_13529);
and U14088 (N_14088,N_13948,N_13604);
xor U14089 (N_14089,N_13746,N_13758);
and U14090 (N_14090,N_13692,N_13610);
xor U14091 (N_14091,N_13742,N_13557);
or U14092 (N_14092,N_13846,N_13716);
and U14093 (N_14093,N_13865,N_13802);
nand U14094 (N_14094,N_13720,N_13824);
and U14095 (N_14095,N_13684,N_13663);
or U14096 (N_14096,N_13555,N_13554);
nand U14097 (N_14097,N_13770,N_13533);
nand U14098 (N_14098,N_13737,N_13577);
nand U14099 (N_14099,N_13609,N_13650);
or U14100 (N_14100,N_13596,N_13937);
xnor U14101 (N_14101,N_13852,N_13727);
and U14102 (N_14102,N_13900,N_13562);
or U14103 (N_14103,N_13981,N_13782);
and U14104 (N_14104,N_13842,N_13798);
and U14105 (N_14105,N_13830,N_13548);
nor U14106 (N_14106,N_13969,N_13902);
and U14107 (N_14107,N_13760,N_13821);
nand U14108 (N_14108,N_13694,N_13801);
xnor U14109 (N_14109,N_13975,N_13608);
xnor U14110 (N_14110,N_13959,N_13651);
nand U14111 (N_14111,N_13819,N_13743);
xnor U14112 (N_14112,N_13915,N_13674);
or U14113 (N_14113,N_13885,N_13759);
or U14114 (N_14114,N_13883,N_13991);
nor U14115 (N_14115,N_13528,N_13733);
xor U14116 (N_14116,N_13923,N_13532);
nor U14117 (N_14117,N_13927,N_13583);
or U14118 (N_14118,N_13825,N_13621);
or U14119 (N_14119,N_13568,N_13870);
nand U14120 (N_14120,N_13947,N_13628);
nor U14121 (N_14121,N_13873,N_13748);
nand U14122 (N_14122,N_13543,N_13683);
nor U14123 (N_14123,N_13815,N_13576);
or U14124 (N_14124,N_13526,N_13891);
nand U14125 (N_14125,N_13721,N_13597);
or U14126 (N_14126,N_13725,N_13893);
nor U14127 (N_14127,N_13779,N_13867);
nand U14128 (N_14128,N_13558,N_13632);
or U14129 (N_14129,N_13522,N_13924);
or U14130 (N_14130,N_13625,N_13658);
nand U14131 (N_14131,N_13987,N_13627);
nor U14132 (N_14132,N_13603,N_13613);
nand U14133 (N_14133,N_13662,N_13724);
or U14134 (N_14134,N_13643,N_13954);
nand U14135 (N_14135,N_13521,N_13586);
nand U14136 (N_14136,N_13722,N_13800);
xor U14137 (N_14137,N_13894,N_13933);
and U14138 (N_14138,N_13702,N_13606);
xor U14139 (N_14139,N_13769,N_13690);
nor U14140 (N_14140,N_13806,N_13729);
nand U14141 (N_14141,N_13984,N_13605);
nand U14142 (N_14142,N_13600,N_13689);
or U14143 (N_14143,N_13719,N_13728);
and U14144 (N_14144,N_13503,N_13739);
and U14145 (N_14145,N_13872,N_13730);
and U14146 (N_14146,N_13892,N_13949);
and U14147 (N_14147,N_13516,N_13594);
and U14148 (N_14148,N_13705,N_13581);
nand U14149 (N_14149,N_13989,N_13707);
xor U14150 (N_14150,N_13717,N_13966);
nor U14151 (N_14151,N_13691,N_13752);
nand U14152 (N_14152,N_13549,N_13973);
nor U14153 (N_14153,N_13504,N_13709);
and U14154 (N_14154,N_13951,N_13584);
or U14155 (N_14155,N_13908,N_13995);
and U14156 (N_14156,N_13835,N_13701);
nand U14157 (N_14157,N_13845,N_13794);
nand U14158 (N_14158,N_13678,N_13734);
and U14159 (N_14159,N_13823,N_13887);
xnor U14160 (N_14160,N_13715,N_13839);
nor U14161 (N_14161,N_13856,N_13644);
or U14162 (N_14162,N_13886,N_13542);
nor U14163 (N_14163,N_13811,N_13988);
nor U14164 (N_14164,N_13735,N_13985);
or U14165 (N_14165,N_13544,N_13945);
nor U14166 (N_14166,N_13879,N_13808);
xor U14167 (N_14167,N_13840,N_13612);
and U14168 (N_14168,N_13539,N_13679);
xor U14169 (N_14169,N_13595,N_13668);
nand U14170 (N_14170,N_13515,N_13967);
and U14171 (N_14171,N_13863,N_13964);
or U14172 (N_14172,N_13797,N_13901);
or U14173 (N_14173,N_13623,N_13907);
nand U14174 (N_14174,N_13910,N_13640);
nand U14175 (N_14175,N_13855,N_13753);
nor U14176 (N_14176,N_13755,N_13950);
nand U14177 (N_14177,N_13669,N_13601);
xor U14178 (N_14178,N_13813,N_13671);
and U14179 (N_14179,N_13700,N_13670);
and U14180 (N_14180,N_13884,N_13693);
nor U14181 (N_14181,N_13807,N_13744);
and U14182 (N_14182,N_13763,N_13866);
nor U14183 (N_14183,N_13631,N_13550);
or U14184 (N_14184,N_13629,N_13675);
nor U14185 (N_14185,N_13983,N_13545);
and U14186 (N_14186,N_13857,N_13974);
nand U14187 (N_14187,N_13566,N_13931);
and U14188 (N_14188,N_13790,N_13768);
xor U14189 (N_14189,N_13547,N_13563);
nand U14190 (N_14190,N_13708,N_13614);
nand U14191 (N_14191,N_13868,N_13552);
or U14192 (N_14192,N_13537,N_13578);
or U14193 (N_14193,N_13853,N_13525);
nor U14194 (N_14194,N_13637,N_13573);
nor U14195 (N_14195,N_13502,N_13982);
and U14196 (N_14196,N_13633,N_13645);
nand U14197 (N_14197,N_13912,N_13942);
nand U14198 (N_14198,N_13741,N_13761);
xnor U14199 (N_14199,N_13688,N_13771);
or U14200 (N_14200,N_13619,N_13738);
nand U14201 (N_14201,N_13848,N_13864);
or U14202 (N_14202,N_13750,N_13789);
nor U14203 (N_14203,N_13956,N_13828);
and U14204 (N_14204,N_13534,N_13622);
xor U14205 (N_14205,N_13667,N_13875);
and U14206 (N_14206,N_13816,N_13574);
nand U14207 (N_14207,N_13896,N_13809);
and U14208 (N_14208,N_13774,N_13511);
nand U14209 (N_14209,N_13505,N_13785);
nand U14210 (N_14210,N_13820,N_13928);
or U14211 (N_14211,N_13793,N_13607);
nor U14212 (N_14212,N_13747,N_13513);
xnor U14213 (N_14213,N_13822,N_13745);
xor U14214 (N_14214,N_13962,N_13756);
nand U14215 (N_14215,N_13946,N_13579);
and U14216 (N_14216,N_13714,N_13904);
and U14217 (N_14217,N_13656,N_13970);
or U14218 (N_14218,N_13589,N_13971);
or U14219 (N_14219,N_13536,N_13844);
or U14220 (N_14220,N_13665,N_13903);
xor U14221 (N_14221,N_13941,N_13704);
or U14222 (N_14222,N_13998,N_13647);
xor U14223 (N_14223,N_13736,N_13588);
or U14224 (N_14224,N_13659,N_13952);
nand U14225 (N_14225,N_13685,N_13686);
xnor U14226 (N_14226,N_13757,N_13777);
or U14227 (N_14227,N_13740,N_13530);
or U14228 (N_14228,N_13976,N_13889);
nand U14229 (N_14229,N_13638,N_13992);
xnor U14230 (N_14230,N_13936,N_13833);
xor U14231 (N_14231,N_13906,N_13851);
xnor U14232 (N_14232,N_13961,N_13990);
and U14233 (N_14233,N_13710,N_13805);
xor U14234 (N_14234,N_13880,N_13514);
or U14235 (N_14235,N_13938,N_13881);
or U14236 (N_14236,N_13630,N_13510);
or U14237 (N_14237,N_13587,N_13732);
nor U14238 (N_14238,N_13796,N_13695);
or U14239 (N_14239,N_13859,N_13826);
nand U14240 (N_14240,N_13582,N_13843);
and U14241 (N_14241,N_13718,N_13841);
or U14242 (N_14242,N_13598,N_13501);
and U14243 (N_14243,N_13996,N_13780);
xnor U14244 (N_14244,N_13860,N_13943);
nand U14245 (N_14245,N_13775,N_13773);
or U14246 (N_14246,N_13523,N_13778);
and U14247 (N_14247,N_13888,N_13635);
or U14248 (N_14248,N_13680,N_13762);
nand U14249 (N_14249,N_13994,N_13814);
nor U14250 (N_14250,N_13695,N_13978);
or U14251 (N_14251,N_13906,N_13611);
or U14252 (N_14252,N_13529,N_13558);
or U14253 (N_14253,N_13928,N_13848);
or U14254 (N_14254,N_13913,N_13692);
xor U14255 (N_14255,N_13882,N_13728);
and U14256 (N_14256,N_13836,N_13589);
or U14257 (N_14257,N_13555,N_13855);
xor U14258 (N_14258,N_13971,N_13784);
or U14259 (N_14259,N_13936,N_13543);
xor U14260 (N_14260,N_13698,N_13599);
nand U14261 (N_14261,N_13821,N_13807);
nand U14262 (N_14262,N_13895,N_13796);
nand U14263 (N_14263,N_13809,N_13546);
xor U14264 (N_14264,N_13744,N_13588);
or U14265 (N_14265,N_13769,N_13670);
or U14266 (N_14266,N_13585,N_13530);
nor U14267 (N_14267,N_13940,N_13843);
and U14268 (N_14268,N_13925,N_13513);
nand U14269 (N_14269,N_13995,N_13666);
nor U14270 (N_14270,N_13690,N_13925);
and U14271 (N_14271,N_13651,N_13759);
and U14272 (N_14272,N_13849,N_13647);
or U14273 (N_14273,N_13999,N_13564);
xor U14274 (N_14274,N_13809,N_13531);
nor U14275 (N_14275,N_13622,N_13815);
or U14276 (N_14276,N_13662,N_13735);
and U14277 (N_14277,N_13649,N_13824);
xnor U14278 (N_14278,N_13704,N_13730);
or U14279 (N_14279,N_13894,N_13531);
xnor U14280 (N_14280,N_13896,N_13598);
nor U14281 (N_14281,N_13598,N_13618);
nor U14282 (N_14282,N_13814,N_13725);
and U14283 (N_14283,N_13641,N_13636);
nand U14284 (N_14284,N_13906,N_13993);
or U14285 (N_14285,N_13892,N_13956);
or U14286 (N_14286,N_13943,N_13765);
and U14287 (N_14287,N_13569,N_13825);
and U14288 (N_14288,N_13919,N_13547);
nand U14289 (N_14289,N_13801,N_13777);
nand U14290 (N_14290,N_13682,N_13607);
nand U14291 (N_14291,N_13943,N_13848);
and U14292 (N_14292,N_13520,N_13573);
nor U14293 (N_14293,N_13921,N_13930);
or U14294 (N_14294,N_13522,N_13694);
and U14295 (N_14295,N_13877,N_13614);
and U14296 (N_14296,N_13669,N_13780);
nor U14297 (N_14297,N_13929,N_13982);
and U14298 (N_14298,N_13619,N_13973);
nor U14299 (N_14299,N_13778,N_13681);
xnor U14300 (N_14300,N_13789,N_13656);
or U14301 (N_14301,N_13563,N_13953);
or U14302 (N_14302,N_13682,N_13850);
xor U14303 (N_14303,N_13746,N_13948);
or U14304 (N_14304,N_13865,N_13609);
xnor U14305 (N_14305,N_13775,N_13544);
nand U14306 (N_14306,N_13707,N_13804);
xor U14307 (N_14307,N_13595,N_13805);
or U14308 (N_14308,N_13759,N_13932);
xor U14309 (N_14309,N_13635,N_13807);
and U14310 (N_14310,N_13600,N_13884);
xor U14311 (N_14311,N_13578,N_13779);
xnor U14312 (N_14312,N_13689,N_13991);
and U14313 (N_14313,N_13793,N_13959);
nor U14314 (N_14314,N_13903,N_13860);
xor U14315 (N_14315,N_13792,N_13703);
nor U14316 (N_14316,N_13931,N_13811);
or U14317 (N_14317,N_13611,N_13795);
nor U14318 (N_14318,N_13506,N_13728);
and U14319 (N_14319,N_13593,N_13975);
or U14320 (N_14320,N_13965,N_13830);
and U14321 (N_14321,N_13524,N_13602);
and U14322 (N_14322,N_13977,N_13593);
and U14323 (N_14323,N_13821,N_13617);
nor U14324 (N_14324,N_13817,N_13645);
and U14325 (N_14325,N_13901,N_13781);
xor U14326 (N_14326,N_13884,N_13621);
or U14327 (N_14327,N_13586,N_13951);
or U14328 (N_14328,N_13808,N_13683);
and U14329 (N_14329,N_13867,N_13679);
nand U14330 (N_14330,N_13974,N_13867);
xnor U14331 (N_14331,N_13522,N_13801);
nor U14332 (N_14332,N_13807,N_13783);
nand U14333 (N_14333,N_13641,N_13720);
xnor U14334 (N_14334,N_13999,N_13893);
nor U14335 (N_14335,N_13743,N_13674);
nor U14336 (N_14336,N_13528,N_13915);
or U14337 (N_14337,N_13844,N_13836);
xor U14338 (N_14338,N_13770,N_13972);
nand U14339 (N_14339,N_13740,N_13731);
or U14340 (N_14340,N_13575,N_13891);
xnor U14341 (N_14341,N_13806,N_13918);
nand U14342 (N_14342,N_13665,N_13817);
nand U14343 (N_14343,N_13789,N_13545);
xor U14344 (N_14344,N_13612,N_13802);
nor U14345 (N_14345,N_13621,N_13728);
and U14346 (N_14346,N_13952,N_13829);
nand U14347 (N_14347,N_13693,N_13969);
and U14348 (N_14348,N_13883,N_13972);
nor U14349 (N_14349,N_13565,N_13642);
and U14350 (N_14350,N_13719,N_13872);
and U14351 (N_14351,N_13519,N_13985);
or U14352 (N_14352,N_13520,N_13991);
nor U14353 (N_14353,N_13536,N_13764);
nand U14354 (N_14354,N_13698,N_13988);
xnor U14355 (N_14355,N_13711,N_13553);
and U14356 (N_14356,N_13604,N_13680);
and U14357 (N_14357,N_13645,N_13720);
xnor U14358 (N_14358,N_13969,N_13916);
nand U14359 (N_14359,N_13798,N_13989);
and U14360 (N_14360,N_13673,N_13852);
nor U14361 (N_14361,N_13767,N_13630);
xnor U14362 (N_14362,N_13677,N_13542);
and U14363 (N_14363,N_13999,N_13618);
and U14364 (N_14364,N_13973,N_13673);
nand U14365 (N_14365,N_13618,N_13845);
nand U14366 (N_14366,N_13661,N_13850);
or U14367 (N_14367,N_13995,N_13964);
or U14368 (N_14368,N_13585,N_13968);
and U14369 (N_14369,N_13572,N_13952);
xnor U14370 (N_14370,N_13605,N_13845);
xor U14371 (N_14371,N_13638,N_13720);
and U14372 (N_14372,N_13988,N_13710);
nand U14373 (N_14373,N_13764,N_13502);
nor U14374 (N_14374,N_13834,N_13571);
nor U14375 (N_14375,N_13856,N_13534);
nand U14376 (N_14376,N_13774,N_13813);
nand U14377 (N_14377,N_13508,N_13799);
xnor U14378 (N_14378,N_13679,N_13986);
or U14379 (N_14379,N_13889,N_13833);
or U14380 (N_14380,N_13872,N_13620);
and U14381 (N_14381,N_13757,N_13508);
xnor U14382 (N_14382,N_13736,N_13790);
nand U14383 (N_14383,N_13962,N_13599);
nand U14384 (N_14384,N_13956,N_13706);
nor U14385 (N_14385,N_13584,N_13578);
xnor U14386 (N_14386,N_13804,N_13791);
xnor U14387 (N_14387,N_13604,N_13724);
xnor U14388 (N_14388,N_13709,N_13875);
or U14389 (N_14389,N_13874,N_13534);
and U14390 (N_14390,N_13812,N_13565);
nor U14391 (N_14391,N_13617,N_13895);
or U14392 (N_14392,N_13964,N_13840);
or U14393 (N_14393,N_13902,N_13954);
and U14394 (N_14394,N_13586,N_13804);
and U14395 (N_14395,N_13726,N_13940);
or U14396 (N_14396,N_13558,N_13750);
or U14397 (N_14397,N_13826,N_13502);
xor U14398 (N_14398,N_13768,N_13950);
and U14399 (N_14399,N_13623,N_13500);
xnor U14400 (N_14400,N_13862,N_13534);
xor U14401 (N_14401,N_13520,N_13954);
xnor U14402 (N_14402,N_13731,N_13643);
or U14403 (N_14403,N_13788,N_13771);
nand U14404 (N_14404,N_13557,N_13506);
nand U14405 (N_14405,N_13919,N_13950);
or U14406 (N_14406,N_13585,N_13555);
nor U14407 (N_14407,N_13754,N_13717);
xor U14408 (N_14408,N_13706,N_13585);
nand U14409 (N_14409,N_13860,N_13988);
nand U14410 (N_14410,N_13987,N_13728);
and U14411 (N_14411,N_13586,N_13700);
xor U14412 (N_14412,N_13678,N_13570);
nand U14413 (N_14413,N_13934,N_13660);
nor U14414 (N_14414,N_13844,N_13975);
xnor U14415 (N_14415,N_13871,N_13914);
or U14416 (N_14416,N_13647,N_13960);
nand U14417 (N_14417,N_13504,N_13913);
xor U14418 (N_14418,N_13878,N_13815);
or U14419 (N_14419,N_13948,N_13736);
xnor U14420 (N_14420,N_13528,N_13506);
xor U14421 (N_14421,N_13744,N_13954);
or U14422 (N_14422,N_13931,N_13558);
nand U14423 (N_14423,N_13730,N_13719);
nand U14424 (N_14424,N_13766,N_13983);
nor U14425 (N_14425,N_13604,N_13669);
nor U14426 (N_14426,N_13580,N_13825);
nor U14427 (N_14427,N_13578,N_13675);
or U14428 (N_14428,N_13930,N_13958);
or U14429 (N_14429,N_13519,N_13552);
nand U14430 (N_14430,N_13693,N_13561);
or U14431 (N_14431,N_13731,N_13952);
and U14432 (N_14432,N_13933,N_13620);
or U14433 (N_14433,N_13970,N_13637);
nor U14434 (N_14434,N_13928,N_13557);
and U14435 (N_14435,N_13884,N_13652);
xnor U14436 (N_14436,N_13713,N_13601);
and U14437 (N_14437,N_13655,N_13934);
nand U14438 (N_14438,N_13851,N_13566);
nor U14439 (N_14439,N_13517,N_13633);
nand U14440 (N_14440,N_13819,N_13578);
and U14441 (N_14441,N_13655,N_13731);
nand U14442 (N_14442,N_13646,N_13774);
xor U14443 (N_14443,N_13975,N_13917);
nand U14444 (N_14444,N_13875,N_13958);
nor U14445 (N_14445,N_13882,N_13550);
and U14446 (N_14446,N_13665,N_13697);
nand U14447 (N_14447,N_13878,N_13762);
or U14448 (N_14448,N_13921,N_13659);
and U14449 (N_14449,N_13742,N_13977);
nand U14450 (N_14450,N_13706,N_13809);
and U14451 (N_14451,N_13942,N_13505);
nand U14452 (N_14452,N_13644,N_13549);
or U14453 (N_14453,N_13638,N_13783);
nand U14454 (N_14454,N_13518,N_13551);
or U14455 (N_14455,N_13543,N_13802);
xnor U14456 (N_14456,N_13568,N_13729);
or U14457 (N_14457,N_13851,N_13587);
nor U14458 (N_14458,N_13619,N_13576);
or U14459 (N_14459,N_13652,N_13605);
xnor U14460 (N_14460,N_13694,N_13662);
nand U14461 (N_14461,N_13691,N_13787);
nor U14462 (N_14462,N_13971,N_13558);
xor U14463 (N_14463,N_13954,N_13932);
nor U14464 (N_14464,N_13957,N_13577);
nand U14465 (N_14465,N_13874,N_13851);
nor U14466 (N_14466,N_13540,N_13680);
xor U14467 (N_14467,N_13695,N_13610);
nor U14468 (N_14468,N_13541,N_13532);
or U14469 (N_14469,N_13503,N_13759);
nor U14470 (N_14470,N_13936,N_13894);
xor U14471 (N_14471,N_13948,N_13507);
or U14472 (N_14472,N_13938,N_13673);
nand U14473 (N_14473,N_13838,N_13697);
or U14474 (N_14474,N_13583,N_13681);
nand U14475 (N_14475,N_13618,N_13701);
or U14476 (N_14476,N_13614,N_13569);
nand U14477 (N_14477,N_13998,N_13696);
nand U14478 (N_14478,N_13982,N_13983);
nand U14479 (N_14479,N_13860,N_13675);
and U14480 (N_14480,N_13655,N_13849);
or U14481 (N_14481,N_13590,N_13503);
and U14482 (N_14482,N_13982,N_13873);
nor U14483 (N_14483,N_13985,N_13969);
and U14484 (N_14484,N_13870,N_13821);
and U14485 (N_14485,N_13559,N_13513);
and U14486 (N_14486,N_13739,N_13718);
xnor U14487 (N_14487,N_13529,N_13523);
nand U14488 (N_14488,N_13970,N_13844);
nor U14489 (N_14489,N_13772,N_13599);
or U14490 (N_14490,N_13734,N_13574);
or U14491 (N_14491,N_13621,N_13965);
or U14492 (N_14492,N_13598,N_13732);
nor U14493 (N_14493,N_13808,N_13967);
and U14494 (N_14494,N_13679,N_13747);
nand U14495 (N_14495,N_13797,N_13530);
nand U14496 (N_14496,N_13513,N_13712);
xnor U14497 (N_14497,N_13511,N_13925);
and U14498 (N_14498,N_13625,N_13849);
nand U14499 (N_14499,N_13622,N_13904);
nand U14500 (N_14500,N_14234,N_14224);
and U14501 (N_14501,N_14100,N_14111);
and U14502 (N_14502,N_14069,N_14495);
or U14503 (N_14503,N_14028,N_14050);
xor U14504 (N_14504,N_14214,N_14181);
nand U14505 (N_14505,N_14494,N_14479);
and U14506 (N_14506,N_14299,N_14078);
nand U14507 (N_14507,N_14052,N_14219);
nand U14508 (N_14508,N_14484,N_14316);
xor U14509 (N_14509,N_14195,N_14089);
nand U14510 (N_14510,N_14136,N_14368);
nand U14511 (N_14511,N_14308,N_14105);
nor U14512 (N_14512,N_14126,N_14481);
nor U14513 (N_14513,N_14034,N_14048);
nor U14514 (N_14514,N_14325,N_14376);
or U14515 (N_14515,N_14120,N_14182);
or U14516 (N_14516,N_14393,N_14141);
nand U14517 (N_14517,N_14337,N_14019);
and U14518 (N_14518,N_14146,N_14360);
nor U14519 (N_14519,N_14400,N_14338);
or U14520 (N_14520,N_14040,N_14462);
or U14521 (N_14521,N_14386,N_14109);
and U14522 (N_14522,N_14327,N_14118);
or U14523 (N_14523,N_14364,N_14446);
or U14524 (N_14524,N_14199,N_14018);
nand U14525 (N_14525,N_14450,N_14275);
nand U14526 (N_14526,N_14084,N_14254);
or U14527 (N_14527,N_14047,N_14403);
nand U14528 (N_14528,N_14440,N_14432);
nor U14529 (N_14529,N_14188,N_14090);
and U14530 (N_14530,N_14178,N_14119);
xnor U14531 (N_14531,N_14391,N_14080);
nor U14532 (N_14532,N_14343,N_14443);
nor U14533 (N_14533,N_14057,N_14056);
and U14534 (N_14534,N_14483,N_14285);
nor U14535 (N_14535,N_14428,N_14197);
nor U14536 (N_14536,N_14005,N_14332);
nor U14537 (N_14537,N_14088,N_14253);
xor U14538 (N_14538,N_14326,N_14274);
or U14539 (N_14539,N_14405,N_14128);
and U14540 (N_14540,N_14221,N_14485);
or U14541 (N_14541,N_14074,N_14108);
or U14542 (N_14542,N_14045,N_14349);
or U14543 (N_14543,N_14346,N_14211);
nor U14544 (N_14544,N_14022,N_14054);
and U14545 (N_14545,N_14116,N_14377);
nand U14546 (N_14546,N_14044,N_14137);
nand U14547 (N_14547,N_14430,N_14016);
nor U14548 (N_14548,N_14342,N_14294);
nor U14549 (N_14549,N_14063,N_14099);
or U14550 (N_14550,N_14310,N_14236);
nor U14551 (N_14551,N_14464,N_14408);
xor U14552 (N_14552,N_14114,N_14431);
nor U14553 (N_14553,N_14046,N_14129);
nand U14554 (N_14554,N_14399,N_14055);
xnor U14555 (N_14555,N_14010,N_14470);
and U14556 (N_14556,N_14421,N_14363);
or U14557 (N_14557,N_14015,N_14142);
or U14558 (N_14558,N_14249,N_14272);
nand U14559 (N_14559,N_14499,N_14395);
and U14560 (N_14560,N_14060,N_14365);
or U14561 (N_14561,N_14148,N_14175);
xnor U14562 (N_14562,N_14351,N_14061);
nor U14563 (N_14563,N_14264,N_14230);
and U14564 (N_14564,N_14110,N_14257);
nor U14565 (N_14565,N_14345,N_14389);
xnor U14566 (N_14566,N_14314,N_14058);
nor U14567 (N_14567,N_14165,N_14134);
nand U14568 (N_14568,N_14107,N_14466);
and U14569 (N_14569,N_14328,N_14177);
and U14570 (N_14570,N_14172,N_14087);
or U14571 (N_14571,N_14176,N_14472);
nand U14572 (N_14572,N_14256,N_14280);
nor U14573 (N_14573,N_14038,N_14497);
or U14574 (N_14574,N_14453,N_14324);
nand U14575 (N_14575,N_14179,N_14416);
nor U14576 (N_14576,N_14384,N_14482);
nor U14577 (N_14577,N_14398,N_14448);
or U14578 (N_14578,N_14232,N_14245);
nand U14579 (N_14579,N_14438,N_14309);
or U14580 (N_14580,N_14281,N_14139);
xnor U14581 (N_14581,N_14207,N_14027);
and U14582 (N_14582,N_14258,N_14273);
or U14583 (N_14583,N_14457,N_14315);
nor U14584 (N_14584,N_14298,N_14373);
or U14585 (N_14585,N_14321,N_14460);
and U14586 (N_14586,N_14348,N_14155);
and U14587 (N_14587,N_14132,N_14076);
and U14588 (N_14588,N_14041,N_14077);
or U14589 (N_14589,N_14218,N_14255);
xor U14590 (N_14590,N_14478,N_14117);
and U14591 (N_14591,N_14357,N_14292);
and U14592 (N_14592,N_14250,N_14290);
nor U14593 (N_14593,N_14169,N_14289);
xor U14594 (N_14594,N_14190,N_14334);
nand U14595 (N_14595,N_14268,N_14192);
or U14596 (N_14596,N_14106,N_14020);
nor U14597 (N_14597,N_14419,N_14387);
or U14598 (N_14598,N_14458,N_14480);
or U14599 (N_14599,N_14378,N_14157);
xnor U14600 (N_14600,N_14124,N_14282);
nand U14601 (N_14601,N_14145,N_14210);
xnor U14602 (N_14602,N_14051,N_14156);
nand U14603 (N_14603,N_14201,N_14433);
nand U14604 (N_14604,N_14390,N_14449);
or U14605 (N_14605,N_14239,N_14371);
xor U14606 (N_14606,N_14380,N_14067);
xor U14607 (N_14607,N_14247,N_14293);
nor U14608 (N_14608,N_14000,N_14070);
or U14609 (N_14609,N_14208,N_14341);
and U14610 (N_14610,N_14414,N_14131);
nand U14611 (N_14611,N_14217,N_14185);
nand U14612 (N_14612,N_14152,N_14191);
and U14613 (N_14613,N_14382,N_14103);
xnor U14614 (N_14614,N_14062,N_14427);
and U14615 (N_14615,N_14461,N_14468);
or U14616 (N_14616,N_14270,N_14033);
nand U14617 (N_14617,N_14323,N_14251);
and U14618 (N_14618,N_14037,N_14228);
and U14619 (N_14619,N_14196,N_14276);
and U14620 (N_14620,N_14227,N_14222);
or U14621 (N_14621,N_14333,N_14154);
xor U14622 (N_14622,N_14417,N_14489);
nand U14623 (N_14623,N_14161,N_14407);
nand U14624 (N_14624,N_14490,N_14159);
or U14625 (N_14625,N_14434,N_14306);
xor U14626 (N_14626,N_14189,N_14486);
nand U14627 (N_14627,N_14260,N_14241);
xnor U14628 (N_14628,N_14335,N_14204);
and U14629 (N_14629,N_14355,N_14474);
nand U14630 (N_14630,N_14029,N_14082);
nand U14631 (N_14631,N_14259,N_14238);
and U14632 (N_14632,N_14226,N_14149);
nor U14633 (N_14633,N_14001,N_14085);
nor U14634 (N_14634,N_14475,N_14375);
nor U14635 (N_14635,N_14206,N_14144);
nor U14636 (N_14636,N_14053,N_14354);
nand U14637 (N_14637,N_14340,N_14115);
or U14638 (N_14638,N_14445,N_14477);
and U14639 (N_14639,N_14243,N_14094);
and U14640 (N_14640,N_14198,N_14496);
xnor U14641 (N_14641,N_14168,N_14415);
nand U14642 (N_14642,N_14125,N_14064);
nor U14643 (N_14643,N_14488,N_14014);
or U14644 (N_14644,N_14013,N_14130);
and U14645 (N_14645,N_14491,N_14498);
and U14646 (N_14646,N_14411,N_14353);
and U14647 (N_14647,N_14248,N_14300);
and U14648 (N_14648,N_14233,N_14113);
nand U14649 (N_14649,N_14223,N_14404);
nand U14650 (N_14650,N_14262,N_14469);
xnor U14651 (N_14651,N_14383,N_14009);
nor U14652 (N_14652,N_14283,N_14442);
or U14653 (N_14653,N_14213,N_14406);
nand U14654 (N_14654,N_14359,N_14303);
nor U14655 (N_14655,N_14127,N_14288);
nand U14656 (N_14656,N_14456,N_14329);
xnor U14657 (N_14657,N_14073,N_14180);
nor U14658 (N_14658,N_14344,N_14410);
or U14659 (N_14659,N_14279,N_14418);
xnor U14660 (N_14660,N_14002,N_14122);
nor U14661 (N_14661,N_14467,N_14297);
xnor U14662 (N_14662,N_14271,N_14339);
nor U14663 (N_14663,N_14413,N_14242);
xnor U14664 (N_14664,N_14350,N_14347);
or U14665 (N_14665,N_14066,N_14187);
xnor U14666 (N_14666,N_14059,N_14231);
or U14667 (N_14667,N_14437,N_14296);
nor U14668 (N_14668,N_14140,N_14287);
or U14669 (N_14669,N_14035,N_14476);
or U14670 (N_14670,N_14183,N_14162);
xor U14671 (N_14671,N_14394,N_14269);
or U14672 (N_14672,N_14240,N_14021);
nor U14673 (N_14673,N_14039,N_14401);
nand U14674 (N_14674,N_14225,N_14277);
xor U14675 (N_14675,N_14186,N_14244);
nand U14676 (N_14676,N_14302,N_14291);
xnor U14677 (N_14677,N_14312,N_14263);
nor U14678 (N_14678,N_14409,N_14043);
and U14679 (N_14679,N_14374,N_14311);
xor U14680 (N_14680,N_14220,N_14435);
nand U14681 (N_14681,N_14330,N_14003);
nor U14682 (N_14682,N_14305,N_14093);
and U14683 (N_14683,N_14164,N_14397);
xnor U14684 (N_14684,N_14200,N_14265);
xor U14685 (N_14685,N_14203,N_14202);
nand U14686 (N_14686,N_14174,N_14096);
nor U14687 (N_14687,N_14487,N_14492);
nand U14688 (N_14688,N_14173,N_14024);
xnor U14689 (N_14689,N_14246,N_14006);
and U14690 (N_14690,N_14454,N_14423);
xor U14691 (N_14691,N_14036,N_14007);
nor U14692 (N_14692,N_14158,N_14095);
and U14693 (N_14693,N_14163,N_14138);
or U14694 (N_14694,N_14356,N_14235);
and U14695 (N_14695,N_14193,N_14170);
nand U14696 (N_14696,N_14104,N_14429);
or U14697 (N_14697,N_14216,N_14361);
nor U14698 (N_14698,N_14295,N_14215);
or U14699 (N_14699,N_14011,N_14367);
nor U14700 (N_14700,N_14284,N_14008);
nor U14701 (N_14701,N_14097,N_14150);
nand U14702 (N_14702,N_14121,N_14012);
nor U14703 (N_14703,N_14352,N_14369);
xor U14704 (N_14704,N_14102,N_14091);
nor U14705 (N_14705,N_14471,N_14366);
or U14706 (N_14706,N_14455,N_14465);
xor U14707 (N_14707,N_14304,N_14023);
nor U14708 (N_14708,N_14322,N_14370);
nor U14709 (N_14709,N_14336,N_14436);
or U14710 (N_14710,N_14439,N_14166);
and U14711 (N_14711,N_14313,N_14318);
and U14712 (N_14712,N_14194,N_14143);
xnor U14713 (N_14713,N_14301,N_14004);
and U14714 (N_14714,N_14133,N_14017);
nand U14715 (N_14715,N_14042,N_14065);
or U14716 (N_14716,N_14151,N_14071);
nor U14717 (N_14717,N_14463,N_14135);
and U14718 (N_14718,N_14030,N_14026);
nand U14719 (N_14719,N_14459,N_14426);
and U14720 (N_14720,N_14101,N_14153);
and U14721 (N_14721,N_14286,N_14331);
or U14722 (N_14722,N_14424,N_14031);
and U14723 (N_14723,N_14025,N_14184);
nor U14724 (N_14724,N_14320,N_14392);
nand U14725 (N_14725,N_14441,N_14420);
nor U14726 (N_14726,N_14229,N_14092);
and U14727 (N_14727,N_14388,N_14160);
nand U14728 (N_14728,N_14317,N_14307);
xor U14729 (N_14729,N_14086,N_14147);
nand U14730 (N_14730,N_14081,N_14451);
nor U14731 (N_14731,N_14425,N_14205);
and U14732 (N_14732,N_14412,N_14123);
nand U14733 (N_14733,N_14252,N_14452);
nand U14734 (N_14734,N_14098,N_14171);
nor U14735 (N_14735,N_14396,N_14237);
nand U14736 (N_14736,N_14266,N_14493);
and U14737 (N_14737,N_14267,N_14385);
nand U14738 (N_14738,N_14362,N_14422);
nand U14739 (N_14739,N_14049,N_14072);
nand U14740 (N_14740,N_14261,N_14075);
nand U14741 (N_14741,N_14372,N_14083);
and U14742 (N_14742,N_14319,N_14032);
xnor U14743 (N_14743,N_14209,N_14278);
and U14744 (N_14744,N_14212,N_14402);
nand U14745 (N_14745,N_14167,N_14068);
nand U14746 (N_14746,N_14444,N_14358);
or U14747 (N_14747,N_14447,N_14079);
xor U14748 (N_14748,N_14379,N_14381);
nand U14749 (N_14749,N_14473,N_14112);
or U14750 (N_14750,N_14276,N_14361);
nand U14751 (N_14751,N_14491,N_14221);
and U14752 (N_14752,N_14112,N_14409);
xnor U14753 (N_14753,N_14226,N_14432);
xnor U14754 (N_14754,N_14362,N_14163);
nand U14755 (N_14755,N_14184,N_14485);
xor U14756 (N_14756,N_14271,N_14003);
xnor U14757 (N_14757,N_14183,N_14352);
nor U14758 (N_14758,N_14427,N_14092);
nand U14759 (N_14759,N_14067,N_14187);
xnor U14760 (N_14760,N_14148,N_14216);
nor U14761 (N_14761,N_14490,N_14497);
or U14762 (N_14762,N_14035,N_14493);
nand U14763 (N_14763,N_14304,N_14303);
or U14764 (N_14764,N_14110,N_14430);
and U14765 (N_14765,N_14323,N_14267);
xnor U14766 (N_14766,N_14099,N_14389);
nor U14767 (N_14767,N_14158,N_14186);
nor U14768 (N_14768,N_14070,N_14071);
and U14769 (N_14769,N_14156,N_14319);
or U14770 (N_14770,N_14433,N_14081);
nand U14771 (N_14771,N_14483,N_14036);
and U14772 (N_14772,N_14265,N_14068);
nor U14773 (N_14773,N_14290,N_14496);
xnor U14774 (N_14774,N_14297,N_14441);
xnor U14775 (N_14775,N_14494,N_14403);
or U14776 (N_14776,N_14111,N_14118);
nor U14777 (N_14777,N_14092,N_14217);
nand U14778 (N_14778,N_14073,N_14050);
nor U14779 (N_14779,N_14071,N_14390);
and U14780 (N_14780,N_14039,N_14273);
xor U14781 (N_14781,N_14280,N_14342);
nand U14782 (N_14782,N_14025,N_14307);
nand U14783 (N_14783,N_14074,N_14029);
nand U14784 (N_14784,N_14051,N_14471);
or U14785 (N_14785,N_14273,N_14074);
xnor U14786 (N_14786,N_14232,N_14247);
nor U14787 (N_14787,N_14035,N_14202);
and U14788 (N_14788,N_14361,N_14306);
or U14789 (N_14789,N_14172,N_14439);
or U14790 (N_14790,N_14319,N_14294);
nor U14791 (N_14791,N_14479,N_14287);
xnor U14792 (N_14792,N_14074,N_14466);
and U14793 (N_14793,N_14137,N_14018);
or U14794 (N_14794,N_14379,N_14119);
nand U14795 (N_14795,N_14411,N_14321);
nand U14796 (N_14796,N_14481,N_14007);
and U14797 (N_14797,N_14385,N_14043);
and U14798 (N_14798,N_14173,N_14134);
or U14799 (N_14799,N_14153,N_14484);
or U14800 (N_14800,N_14286,N_14158);
and U14801 (N_14801,N_14112,N_14467);
xnor U14802 (N_14802,N_14151,N_14483);
or U14803 (N_14803,N_14305,N_14231);
and U14804 (N_14804,N_14115,N_14428);
and U14805 (N_14805,N_14441,N_14172);
or U14806 (N_14806,N_14318,N_14353);
nor U14807 (N_14807,N_14268,N_14001);
or U14808 (N_14808,N_14220,N_14099);
nor U14809 (N_14809,N_14100,N_14477);
or U14810 (N_14810,N_14356,N_14472);
or U14811 (N_14811,N_14106,N_14261);
and U14812 (N_14812,N_14328,N_14184);
xor U14813 (N_14813,N_14168,N_14013);
xor U14814 (N_14814,N_14399,N_14379);
and U14815 (N_14815,N_14002,N_14436);
or U14816 (N_14816,N_14344,N_14420);
and U14817 (N_14817,N_14141,N_14279);
nor U14818 (N_14818,N_14144,N_14003);
nand U14819 (N_14819,N_14218,N_14018);
and U14820 (N_14820,N_14177,N_14131);
and U14821 (N_14821,N_14442,N_14416);
xor U14822 (N_14822,N_14268,N_14422);
nand U14823 (N_14823,N_14164,N_14227);
and U14824 (N_14824,N_14233,N_14367);
nand U14825 (N_14825,N_14366,N_14354);
and U14826 (N_14826,N_14486,N_14289);
or U14827 (N_14827,N_14295,N_14199);
nor U14828 (N_14828,N_14031,N_14462);
xor U14829 (N_14829,N_14194,N_14438);
nand U14830 (N_14830,N_14133,N_14413);
and U14831 (N_14831,N_14288,N_14276);
or U14832 (N_14832,N_14175,N_14295);
or U14833 (N_14833,N_14230,N_14378);
or U14834 (N_14834,N_14071,N_14394);
xnor U14835 (N_14835,N_14446,N_14181);
nand U14836 (N_14836,N_14146,N_14085);
nand U14837 (N_14837,N_14425,N_14152);
nor U14838 (N_14838,N_14129,N_14187);
xnor U14839 (N_14839,N_14244,N_14421);
nand U14840 (N_14840,N_14245,N_14202);
or U14841 (N_14841,N_14043,N_14047);
nor U14842 (N_14842,N_14159,N_14430);
and U14843 (N_14843,N_14221,N_14278);
and U14844 (N_14844,N_14106,N_14005);
xnor U14845 (N_14845,N_14421,N_14189);
nor U14846 (N_14846,N_14101,N_14176);
xor U14847 (N_14847,N_14179,N_14101);
xor U14848 (N_14848,N_14406,N_14156);
or U14849 (N_14849,N_14462,N_14213);
nand U14850 (N_14850,N_14081,N_14149);
or U14851 (N_14851,N_14192,N_14372);
and U14852 (N_14852,N_14444,N_14220);
or U14853 (N_14853,N_14272,N_14268);
nand U14854 (N_14854,N_14087,N_14005);
and U14855 (N_14855,N_14273,N_14249);
nand U14856 (N_14856,N_14293,N_14110);
and U14857 (N_14857,N_14446,N_14198);
xnor U14858 (N_14858,N_14319,N_14285);
nand U14859 (N_14859,N_14114,N_14423);
or U14860 (N_14860,N_14357,N_14356);
nand U14861 (N_14861,N_14313,N_14496);
nor U14862 (N_14862,N_14159,N_14116);
nor U14863 (N_14863,N_14238,N_14229);
and U14864 (N_14864,N_14039,N_14329);
and U14865 (N_14865,N_14138,N_14103);
and U14866 (N_14866,N_14036,N_14324);
nor U14867 (N_14867,N_14304,N_14013);
nand U14868 (N_14868,N_14347,N_14085);
xor U14869 (N_14869,N_14318,N_14472);
or U14870 (N_14870,N_14375,N_14109);
xor U14871 (N_14871,N_14385,N_14158);
nand U14872 (N_14872,N_14139,N_14126);
xor U14873 (N_14873,N_14350,N_14331);
or U14874 (N_14874,N_14165,N_14179);
or U14875 (N_14875,N_14385,N_14474);
nand U14876 (N_14876,N_14423,N_14245);
or U14877 (N_14877,N_14212,N_14351);
and U14878 (N_14878,N_14170,N_14430);
and U14879 (N_14879,N_14455,N_14250);
and U14880 (N_14880,N_14029,N_14451);
xor U14881 (N_14881,N_14282,N_14426);
or U14882 (N_14882,N_14190,N_14269);
nand U14883 (N_14883,N_14060,N_14449);
nor U14884 (N_14884,N_14050,N_14280);
nor U14885 (N_14885,N_14327,N_14344);
and U14886 (N_14886,N_14309,N_14384);
xnor U14887 (N_14887,N_14220,N_14256);
nand U14888 (N_14888,N_14019,N_14232);
and U14889 (N_14889,N_14294,N_14129);
nor U14890 (N_14890,N_14320,N_14445);
or U14891 (N_14891,N_14403,N_14298);
xnor U14892 (N_14892,N_14347,N_14297);
xor U14893 (N_14893,N_14339,N_14362);
and U14894 (N_14894,N_14079,N_14011);
and U14895 (N_14895,N_14376,N_14331);
or U14896 (N_14896,N_14132,N_14170);
xor U14897 (N_14897,N_14251,N_14241);
and U14898 (N_14898,N_14143,N_14030);
nand U14899 (N_14899,N_14029,N_14410);
or U14900 (N_14900,N_14040,N_14171);
and U14901 (N_14901,N_14318,N_14052);
nand U14902 (N_14902,N_14247,N_14168);
and U14903 (N_14903,N_14072,N_14262);
nand U14904 (N_14904,N_14381,N_14349);
nor U14905 (N_14905,N_14339,N_14402);
xor U14906 (N_14906,N_14358,N_14497);
nand U14907 (N_14907,N_14447,N_14444);
and U14908 (N_14908,N_14264,N_14244);
or U14909 (N_14909,N_14483,N_14100);
xor U14910 (N_14910,N_14326,N_14120);
nand U14911 (N_14911,N_14338,N_14183);
and U14912 (N_14912,N_14349,N_14135);
and U14913 (N_14913,N_14365,N_14147);
nor U14914 (N_14914,N_14042,N_14455);
nor U14915 (N_14915,N_14490,N_14421);
xor U14916 (N_14916,N_14368,N_14302);
nand U14917 (N_14917,N_14455,N_14367);
nand U14918 (N_14918,N_14130,N_14250);
nand U14919 (N_14919,N_14348,N_14150);
xor U14920 (N_14920,N_14224,N_14009);
and U14921 (N_14921,N_14292,N_14399);
and U14922 (N_14922,N_14355,N_14060);
nand U14923 (N_14923,N_14313,N_14474);
and U14924 (N_14924,N_14319,N_14138);
or U14925 (N_14925,N_14490,N_14018);
nor U14926 (N_14926,N_14025,N_14353);
nand U14927 (N_14927,N_14340,N_14059);
and U14928 (N_14928,N_14465,N_14240);
xnor U14929 (N_14929,N_14275,N_14486);
or U14930 (N_14930,N_14221,N_14025);
nor U14931 (N_14931,N_14127,N_14391);
nand U14932 (N_14932,N_14074,N_14173);
nor U14933 (N_14933,N_14473,N_14217);
and U14934 (N_14934,N_14254,N_14484);
nand U14935 (N_14935,N_14365,N_14394);
and U14936 (N_14936,N_14418,N_14423);
nor U14937 (N_14937,N_14161,N_14340);
or U14938 (N_14938,N_14414,N_14015);
xor U14939 (N_14939,N_14269,N_14294);
nor U14940 (N_14940,N_14162,N_14030);
xor U14941 (N_14941,N_14427,N_14423);
nor U14942 (N_14942,N_14214,N_14082);
nand U14943 (N_14943,N_14124,N_14008);
nor U14944 (N_14944,N_14159,N_14015);
and U14945 (N_14945,N_14035,N_14297);
nor U14946 (N_14946,N_14107,N_14028);
nor U14947 (N_14947,N_14368,N_14249);
xor U14948 (N_14948,N_14447,N_14460);
xor U14949 (N_14949,N_14180,N_14206);
and U14950 (N_14950,N_14439,N_14239);
and U14951 (N_14951,N_14480,N_14454);
nand U14952 (N_14952,N_14245,N_14124);
xor U14953 (N_14953,N_14168,N_14149);
nor U14954 (N_14954,N_14486,N_14365);
or U14955 (N_14955,N_14325,N_14101);
xnor U14956 (N_14956,N_14473,N_14265);
xor U14957 (N_14957,N_14231,N_14129);
nand U14958 (N_14958,N_14032,N_14166);
nor U14959 (N_14959,N_14248,N_14115);
nand U14960 (N_14960,N_14128,N_14414);
or U14961 (N_14961,N_14001,N_14018);
nor U14962 (N_14962,N_14032,N_14053);
and U14963 (N_14963,N_14497,N_14074);
xnor U14964 (N_14964,N_14430,N_14149);
or U14965 (N_14965,N_14134,N_14279);
nand U14966 (N_14966,N_14215,N_14290);
xnor U14967 (N_14967,N_14053,N_14266);
xor U14968 (N_14968,N_14323,N_14361);
nand U14969 (N_14969,N_14302,N_14102);
nor U14970 (N_14970,N_14373,N_14097);
nand U14971 (N_14971,N_14314,N_14317);
and U14972 (N_14972,N_14235,N_14056);
and U14973 (N_14973,N_14419,N_14066);
nor U14974 (N_14974,N_14416,N_14162);
nor U14975 (N_14975,N_14332,N_14279);
or U14976 (N_14976,N_14206,N_14197);
and U14977 (N_14977,N_14093,N_14046);
nor U14978 (N_14978,N_14248,N_14460);
and U14979 (N_14979,N_14301,N_14349);
nand U14980 (N_14980,N_14189,N_14078);
nand U14981 (N_14981,N_14259,N_14320);
and U14982 (N_14982,N_14305,N_14215);
and U14983 (N_14983,N_14488,N_14097);
or U14984 (N_14984,N_14110,N_14114);
xor U14985 (N_14985,N_14450,N_14499);
xor U14986 (N_14986,N_14499,N_14385);
or U14987 (N_14987,N_14206,N_14097);
xnor U14988 (N_14988,N_14396,N_14197);
or U14989 (N_14989,N_14410,N_14231);
nand U14990 (N_14990,N_14254,N_14416);
or U14991 (N_14991,N_14349,N_14221);
nand U14992 (N_14992,N_14368,N_14268);
nor U14993 (N_14993,N_14477,N_14227);
or U14994 (N_14994,N_14061,N_14077);
nand U14995 (N_14995,N_14209,N_14034);
and U14996 (N_14996,N_14227,N_14292);
nand U14997 (N_14997,N_14247,N_14000);
nand U14998 (N_14998,N_14226,N_14232);
or U14999 (N_14999,N_14496,N_14038);
nor U15000 (N_15000,N_14762,N_14542);
nor U15001 (N_15001,N_14525,N_14776);
xor U15002 (N_15002,N_14872,N_14867);
xnor U15003 (N_15003,N_14725,N_14620);
nor U15004 (N_15004,N_14902,N_14691);
nor U15005 (N_15005,N_14837,N_14755);
and U15006 (N_15006,N_14571,N_14971);
and U15007 (N_15007,N_14685,N_14675);
nand U15008 (N_15008,N_14860,N_14652);
nand U15009 (N_15009,N_14640,N_14711);
nor U15010 (N_15010,N_14738,N_14764);
nand U15011 (N_15011,N_14884,N_14927);
and U15012 (N_15012,N_14680,N_14946);
and U15013 (N_15013,N_14744,N_14706);
or U15014 (N_15014,N_14752,N_14812);
or U15015 (N_15015,N_14952,N_14826);
and U15016 (N_15016,N_14741,N_14750);
xnor U15017 (N_15017,N_14507,N_14650);
and U15018 (N_15018,N_14881,N_14642);
or U15019 (N_15019,N_14958,N_14560);
nor U15020 (N_15020,N_14536,N_14736);
nand U15021 (N_15021,N_14777,N_14585);
and U15022 (N_15022,N_14552,N_14689);
nor U15023 (N_15023,N_14861,N_14687);
nand U15024 (N_15024,N_14989,N_14982);
nor U15025 (N_15025,N_14981,N_14896);
nand U15026 (N_15026,N_14576,N_14524);
or U15027 (N_15027,N_14765,N_14830);
or U15028 (N_15028,N_14817,N_14683);
and U15029 (N_15029,N_14802,N_14705);
or U15030 (N_15030,N_14639,N_14596);
nor U15031 (N_15031,N_14723,N_14920);
nand U15032 (N_15032,N_14806,N_14894);
nor U15033 (N_15033,N_14726,N_14681);
nor U15034 (N_15034,N_14959,N_14868);
nand U15035 (N_15035,N_14746,N_14663);
nand U15036 (N_15036,N_14579,N_14692);
and U15037 (N_15037,N_14513,N_14586);
nor U15038 (N_15038,N_14730,N_14630);
nor U15039 (N_15039,N_14561,N_14819);
nand U15040 (N_15040,N_14587,N_14781);
nor U15041 (N_15041,N_14924,N_14610);
nor U15042 (N_15042,N_14594,N_14724);
xnor U15043 (N_15043,N_14885,N_14835);
nand U15044 (N_15044,N_14537,N_14528);
or U15045 (N_15045,N_14916,N_14983);
nor U15046 (N_15046,N_14641,N_14954);
xnor U15047 (N_15047,N_14843,N_14574);
xnor U15048 (N_15048,N_14856,N_14974);
nor U15049 (N_15049,N_14996,N_14906);
xor U15050 (N_15050,N_14609,N_14719);
or U15051 (N_15051,N_14809,N_14508);
nor U15052 (N_15052,N_14666,N_14527);
and U15053 (N_15053,N_14753,N_14945);
nand U15054 (N_15054,N_14504,N_14673);
or U15055 (N_15055,N_14859,N_14688);
nand U15056 (N_15056,N_14814,N_14970);
nand U15057 (N_15057,N_14785,N_14852);
or U15058 (N_15058,N_14873,N_14702);
nor U15059 (N_15059,N_14577,N_14986);
nor U15060 (N_15060,N_14922,N_14784);
nand U15061 (N_15061,N_14758,N_14909);
xnor U15062 (N_15062,N_14729,N_14882);
nor U15063 (N_15063,N_14509,N_14997);
nor U15064 (N_15064,N_14540,N_14770);
or U15065 (N_15065,N_14716,N_14792);
or U15066 (N_15066,N_14998,N_14622);
and U15067 (N_15067,N_14883,N_14766);
or U15068 (N_15068,N_14644,N_14779);
and U15069 (N_15069,N_14858,N_14933);
and U15070 (N_15070,N_14538,N_14635);
nand U15071 (N_15071,N_14928,N_14891);
or U15072 (N_15072,N_14942,N_14512);
and U15073 (N_15073,N_14960,N_14510);
nand U15074 (N_15074,N_14601,N_14818);
and U15075 (N_15075,N_14619,N_14994);
nor U15076 (N_15076,N_14964,N_14816);
xor U15077 (N_15077,N_14667,N_14892);
nand U15078 (N_15078,N_14707,N_14783);
or U15079 (N_15079,N_14502,N_14682);
xor U15080 (N_15080,N_14651,N_14904);
or U15081 (N_15081,N_14780,N_14771);
xnor U15082 (N_15082,N_14742,N_14862);
nand U15083 (N_15083,N_14949,N_14799);
nand U15084 (N_15084,N_14602,N_14815);
xnor U15085 (N_15085,N_14853,N_14804);
nor U15086 (N_15086,N_14846,N_14511);
or U15087 (N_15087,N_14595,N_14539);
or U15088 (N_15088,N_14940,N_14962);
or U15089 (N_15089,N_14645,N_14794);
and U15090 (N_15090,N_14612,N_14751);
nand U15091 (N_15091,N_14695,N_14950);
or U15092 (N_15092,N_14624,N_14598);
or U15093 (N_15093,N_14931,N_14734);
and U15094 (N_15094,N_14939,N_14563);
nor U15095 (N_15095,N_14914,N_14877);
nand U15096 (N_15096,N_14921,N_14968);
and U15097 (N_15097,N_14824,N_14703);
xnor U15098 (N_15098,N_14544,N_14721);
nand U15099 (N_15099,N_14731,N_14580);
and U15100 (N_15100,N_14938,N_14732);
nand U15101 (N_15101,N_14828,N_14661);
xor U15102 (N_15102,N_14932,N_14791);
xnor U15103 (N_15103,N_14555,N_14674);
nor U15104 (N_15104,N_14615,N_14786);
or U15105 (N_15105,N_14572,N_14985);
or U15106 (N_15106,N_14978,N_14649);
nand U15107 (N_15107,N_14693,N_14850);
or U15108 (N_15108,N_14569,N_14517);
xor U15109 (N_15109,N_14531,N_14564);
nor U15110 (N_15110,N_14628,N_14889);
xnor U15111 (N_15111,N_14669,N_14941);
nor U15112 (N_15112,N_14590,N_14518);
nand U15113 (N_15113,N_14728,N_14761);
or U15114 (N_15114,N_14911,N_14803);
xor U15115 (N_15115,N_14603,N_14926);
or U15116 (N_15116,N_14915,N_14529);
nand U15117 (N_15117,N_14829,N_14821);
xor U15118 (N_15118,N_14581,N_14638);
nor U15119 (N_15119,N_14516,N_14717);
and U15120 (N_15120,N_14697,N_14797);
or U15121 (N_15121,N_14643,N_14584);
and U15122 (N_15122,N_14627,N_14832);
nor U15123 (N_15123,N_14648,N_14844);
or U15124 (N_15124,N_14760,N_14617);
nor U15125 (N_15125,N_14745,N_14676);
xor U15126 (N_15126,N_14589,N_14554);
or U15127 (N_15127,N_14629,N_14870);
and U15128 (N_15128,N_14514,N_14957);
nand U15129 (N_15129,N_14879,N_14696);
and U15130 (N_15130,N_14593,N_14948);
nand U15131 (N_15131,N_14965,N_14910);
or U15132 (N_15132,N_14551,N_14848);
nand U15133 (N_15133,N_14637,N_14671);
and U15134 (N_15134,N_14709,N_14523);
xor U15135 (N_15135,N_14833,N_14621);
or U15136 (N_15136,N_14588,N_14546);
xnor U15137 (N_15137,N_14878,N_14698);
nand U15138 (N_15138,N_14570,N_14710);
and U15139 (N_15139,N_14825,N_14715);
nand U15140 (N_15140,N_14718,N_14790);
nand U15141 (N_15141,N_14634,N_14831);
nor U15142 (N_15142,N_14684,N_14827);
nor U15143 (N_15143,N_14953,N_14653);
nand U15144 (N_15144,N_14714,N_14756);
nor U15145 (N_15145,N_14701,N_14887);
or U15146 (N_15146,N_14712,N_14966);
nand U15147 (N_15147,N_14987,N_14795);
or U15148 (N_15148,N_14558,N_14519);
xnor U15149 (N_15149,N_14805,N_14727);
and U15150 (N_15150,N_14599,N_14566);
and U15151 (N_15151,N_14614,N_14611);
or U15152 (N_15152,N_14636,N_14659);
and U15153 (N_15153,N_14631,N_14632);
nor U15154 (N_15154,N_14567,N_14845);
and U15155 (N_15155,N_14789,N_14658);
nor U15156 (N_15156,N_14735,N_14704);
xor U15157 (N_15157,N_14912,N_14907);
or U15158 (N_15158,N_14763,N_14925);
or U15159 (N_15159,N_14670,N_14600);
and U15160 (N_15160,N_14506,N_14759);
xor U15161 (N_15161,N_14810,N_14607);
and U15162 (N_15162,N_14591,N_14672);
xor U15163 (N_15163,N_14993,N_14657);
nand U15164 (N_15164,N_14582,N_14967);
xor U15165 (N_15165,N_14854,N_14740);
nor U15166 (N_15166,N_14545,N_14562);
nor U15167 (N_15167,N_14866,N_14984);
nand U15168 (N_15168,N_14871,N_14908);
and U15169 (N_15169,N_14975,N_14913);
xor U15170 (N_15170,N_14768,N_14800);
and U15171 (N_15171,N_14535,N_14820);
nor U15172 (N_15172,N_14923,N_14990);
nand U15173 (N_15173,N_14654,N_14847);
or U15174 (N_15174,N_14530,N_14855);
nand U15175 (N_15175,N_14647,N_14841);
nor U15176 (N_15176,N_14834,N_14583);
or U15177 (N_15177,N_14869,N_14995);
nand U15178 (N_15178,N_14888,N_14793);
xor U15179 (N_15179,N_14597,N_14655);
nor U15180 (N_15180,N_14905,N_14747);
nand U15181 (N_15181,N_14743,N_14739);
nor U15182 (N_15182,N_14733,N_14899);
xnor U15183 (N_15183,N_14898,N_14501);
nor U15184 (N_15184,N_14573,N_14972);
and U15185 (N_15185,N_14565,N_14807);
nor U15186 (N_15186,N_14690,N_14893);
xnor U15187 (N_15187,N_14973,N_14662);
or U15188 (N_15188,N_14618,N_14991);
nor U15189 (N_15189,N_14961,N_14875);
nor U15190 (N_15190,N_14956,N_14936);
nand U15191 (N_15191,N_14808,N_14935);
nor U15192 (N_15192,N_14969,N_14778);
xnor U15193 (N_15193,N_14823,N_14616);
nand U15194 (N_15194,N_14575,N_14988);
nor U15195 (N_15195,N_14947,N_14608);
xor U15196 (N_15196,N_14559,N_14606);
or U15197 (N_15197,N_14665,N_14592);
or U15198 (N_15198,N_14677,N_14532);
nor U15199 (N_15199,N_14801,N_14526);
and U15200 (N_15200,N_14919,N_14775);
xor U15201 (N_15201,N_14543,N_14534);
nor U15202 (N_15202,N_14839,N_14623);
or U15203 (N_15203,N_14686,N_14521);
and U15204 (N_15204,N_14664,N_14749);
or U15205 (N_15205,N_14976,N_14787);
nand U15206 (N_15206,N_14633,N_14656);
and U15207 (N_15207,N_14550,N_14500);
xor U15208 (N_15208,N_14865,N_14668);
or U15209 (N_15209,N_14798,N_14992);
nand U15210 (N_15210,N_14930,N_14694);
and U15211 (N_15211,N_14604,N_14757);
or U15212 (N_15212,N_14886,N_14660);
nand U15213 (N_15213,N_14900,N_14748);
or U15214 (N_15214,N_14520,N_14549);
nand U15215 (N_15215,N_14568,N_14917);
xor U15216 (N_15216,N_14864,N_14813);
nor U15217 (N_15217,N_14977,N_14713);
and U15218 (N_15218,N_14773,N_14944);
and U15219 (N_15219,N_14943,N_14822);
or U15220 (N_15220,N_14774,N_14720);
nor U15221 (N_15221,N_14842,N_14838);
xnor U15222 (N_15222,N_14836,N_14840);
or U15223 (N_15223,N_14699,N_14541);
or U15224 (N_15224,N_14708,N_14737);
nor U15225 (N_15225,N_14548,N_14999);
nand U15226 (N_15226,N_14918,N_14951);
and U15227 (N_15227,N_14782,N_14980);
or U15228 (N_15228,N_14897,N_14955);
nand U15229 (N_15229,N_14722,N_14890);
or U15230 (N_15230,N_14811,N_14613);
xnor U15231 (N_15231,N_14788,N_14929);
and U15232 (N_15232,N_14937,N_14515);
nor U15233 (N_15233,N_14796,N_14678);
nand U15234 (N_15234,N_14863,N_14849);
or U15235 (N_15235,N_14533,N_14503);
nor U15236 (N_15236,N_14646,N_14625);
nand U15237 (N_15237,N_14963,N_14874);
and U15238 (N_15238,N_14522,N_14679);
nand U15239 (N_15239,N_14578,N_14605);
and U15240 (N_15240,N_14767,N_14880);
and U15241 (N_15241,N_14876,N_14772);
and U15242 (N_15242,N_14556,N_14547);
and U15243 (N_15243,N_14505,N_14557);
and U15244 (N_15244,N_14979,N_14934);
xor U15245 (N_15245,N_14903,N_14851);
xnor U15246 (N_15246,N_14626,N_14769);
and U15247 (N_15247,N_14895,N_14754);
or U15248 (N_15248,N_14857,N_14700);
or U15249 (N_15249,N_14553,N_14901);
xor U15250 (N_15250,N_14511,N_14975);
or U15251 (N_15251,N_14895,N_14786);
nor U15252 (N_15252,N_14937,N_14999);
nor U15253 (N_15253,N_14854,N_14961);
or U15254 (N_15254,N_14783,N_14621);
xor U15255 (N_15255,N_14818,N_14729);
and U15256 (N_15256,N_14654,N_14943);
and U15257 (N_15257,N_14647,N_14794);
nor U15258 (N_15258,N_14906,N_14948);
and U15259 (N_15259,N_14819,N_14822);
nor U15260 (N_15260,N_14701,N_14746);
and U15261 (N_15261,N_14503,N_14612);
nand U15262 (N_15262,N_14549,N_14702);
or U15263 (N_15263,N_14958,N_14525);
and U15264 (N_15264,N_14510,N_14664);
nand U15265 (N_15265,N_14962,N_14935);
nor U15266 (N_15266,N_14708,N_14951);
xor U15267 (N_15267,N_14595,N_14599);
nor U15268 (N_15268,N_14913,N_14667);
xor U15269 (N_15269,N_14720,N_14873);
xnor U15270 (N_15270,N_14512,N_14920);
xnor U15271 (N_15271,N_14600,N_14506);
nand U15272 (N_15272,N_14733,N_14938);
nor U15273 (N_15273,N_14513,N_14761);
nor U15274 (N_15274,N_14980,N_14961);
xor U15275 (N_15275,N_14797,N_14635);
or U15276 (N_15276,N_14948,N_14857);
nor U15277 (N_15277,N_14790,N_14511);
xor U15278 (N_15278,N_14617,N_14813);
and U15279 (N_15279,N_14971,N_14661);
nand U15280 (N_15280,N_14772,N_14959);
and U15281 (N_15281,N_14700,N_14640);
xor U15282 (N_15282,N_14973,N_14891);
or U15283 (N_15283,N_14892,N_14893);
xnor U15284 (N_15284,N_14809,N_14797);
and U15285 (N_15285,N_14751,N_14735);
and U15286 (N_15286,N_14628,N_14817);
or U15287 (N_15287,N_14890,N_14648);
xnor U15288 (N_15288,N_14549,N_14611);
nand U15289 (N_15289,N_14819,N_14565);
and U15290 (N_15290,N_14741,N_14749);
nor U15291 (N_15291,N_14581,N_14644);
and U15292 (N_15292,N_14892,N_14645);
and U15293 (N_15293,N_14646,N_14573);
nand U15294 (N_15294,N_14696,N_14766);
or U15295 (N_15295,N_14556,N_14630);
and U15296 (N_15296,N_14769,N_14752);
nand U15297 (N_15297,N_14584,N_14718);
nor U15298 (N_15298,N_14773,N_14612);
nor U15299 (N_15299,N_14934,N_14847);
and U15300 (N_15300,N_14657,N_14550);
nand U15301 (N_15301,N_14777,N_14602);
nor U15302 (N_15302,N_14919,N_14585);
or U15303 (N_15303,N_14732,N_14714);
xor U15304 (N_15304,N_14553,N_14882);
and U15305 (N_15305,N_14651,N_14853);
xnor U15306 (N_15306,N_14515,N_14820);
and U15307 (N_15307,N_14557,N_14863);
nand U15308 (N_15308,N_14611,N_14624);
and U15309 (N_15309,N_14522,N_14845);
nor U15310 (N_15310,N_14875,N_14987);
nand U15311 (N_15311,N_14671,N_14990);
xor U15312 (N_15312,N_14999,N_14507);
or U15313 (N_15313,N_14801,N_14657);
or U15314 (N_15314,N_14809,N_14746);
or U15315 (N_15315,N_14935,N_14777);
nor U15316 (N_15316,N_14724,N_14722);
and U15317 (N_15317,N_14886,N_14793);
nor U15318 (N_15318,N_14767,N_14588);
and U15319 (N_15319,N_14676,N_14663);
and U15320 (N_15320,N_14879,N_14640);
or U15321 (N_15321,N_14893,N_14821);
xor U15322 (N_15322,N_14865,N_14532);
xor U15323 (N_15323,N_14869,N_14617);
or U15324 (N_15324,N_14807,N_14988);
and U15325 (N_15325,N_14912,N_14653);
or U15326 (N_15326,N_14596,N_14662);
and U15327 (N_15327,N_14976,N_14845);
nand U15328 (N_15328,N_14757,N_14664);
xnor U15329 (N_15329,N_14541,N_14580);
and U15330 (N_15330,N_14818,N_14949);
nor U15331 (N_15331,N_14735,N_14870);
nor U15332 (N_15332,N_14907,N_14995);
nand U15333 (N_15333,N_14619,N_14832);
nor U15334 (N_15334,N_14943,N_14940);
xnor U15335 (N_15335,N_14546,N_14601);
xnor U15336 (N_15336,N_14651,N_14576);
and U15337 (N_15337,N_14808,N_14707);
xnor U15338 (N_15338,N_14552,N_14995);
xnor U15339 (N_15339,N_14802,N_14666);
and U15340 (N_15340,N_14579,N_14866);
nor U15341 (N_15341,N_14522,N_14869);
nand U15342 (N_15342,N_14784,N_14551);
nor U15343 (N_15343,N_14838,N_14864);
and U15344 (N_15344,N_14997,N_14689);
nor U15345 (N_15345,N_14580,N_14906);
and U15346 (N_15346,N_14988,N_14784);
xor U15347 (N_15347,N_14754,N_14584);
or U15348 (N_15348,N_14994,N_14675);
xnor U15349 (N_15349,N_14603,N_14758);
and U15350 (N_15350,N_14612,N_14519);
nand U15351 (N_15351,N_14613,N_14719);
nand U15352 (N_15352,N_14867,N_14991);
nor U15353 (N_15353,N_14760,N_14887);
xor U15354 (N_15354,N_14608,N_14747);
nand U15355 (N_15355,N_14683,N_14855);
xnor U15356 (N_15356,N_14571,N_14722);
or U15357 (N_15357,N_14959,N_14754);
nor U15358 (N_15358,N_14536,N_14936);
or U15359 (N_15359,N_14981,N_14620);
nand U15360 (N_15360,N_14998,N_14706);
and U15361 (N_15361,N_14803,N_14930);
nor U15362 (N_15362,N_14774,N_14558);
and U15363 (N_15363,N_14917,N_14935);
xor U15364 (N_15364,N_14935,N_14654);
xnor U15365 (N_15365,N_14507,N_14967);
xnor U15366 (N_15366,N_14982,N_14809);
xnor U15367 (N_15367,N_14656,N_14706);
or U15368 (N_15368,N_14745,N_14876);
nor U15369 (N_15369,N_14873,N_14681);
nand U15370 (N_15370,N_14623,N_14693);
nand U15371 (N_15371,N_14774,N_14750);
and U15372 (N_15372,N_14773,N_14744);
and U15373 (N_15373,N_14875,N_14976);
nand U15374 (N_15374,N_14693,N_14805);
nand U15375 (N_15375,N_14806,N_14776);
nor U15376 (N_15376,N_14843,N_14928);
and U15377 (N_15377,N_14608,N_14830);
and U15378 (N_15378,N_14609,N_14913);
and U15379 (N_15379,N_14975,N_14508);
nor U15380 (N_15380,N_14875,N_14537);
nor U15381 (N_15381,N_14847,N_14671);
and U15382 (N_15382,N_14888,N_14887);
nor U15383 (N_15383,N_14962,N_14540);
and U15384 (N_15384,N_14976,N_14857);
xor U15385 (N_15385,N_14828,N_14912);
nand U15386 (N_15386,N_14918,N_14611);
nand U15387 (N_15387,N_14581,N_14768);
nor U15388 (N_15388,N_14743,N_14709);
nor U15389 (N_15389,N_14709,N_14611);
xnor U15390 (N_15390,N_14920,N_14914);
xnor U15391 (N_15391,N_14866,N_14673);
xor U15392 (N_15392,N_14504,N_14852);
nand U15393 (N_15393,N_14649,N_14913);
and U15394 (N_15394,N_14734,N_14908);
nand U15395 (N_15395,N_14542,N_14735);
nand U15396 (N_15396,N_14740,N_14917);
nand U15397 (N_15397,N_14560,N_14502);
xnor U15398 (N_15398,N_14958,N_14539);
and U15399 (N_15399,N_14737,N_14562);
nor U15400 (N_15400,N_14695,N_14566);
nand U15401 (N_15401,N_14569,N_14920);
xor U15402 (N_15402,N_14719,N_14957);
nand U15403 (N_15403,N_14718,N_14645);
xnor U15404 (N_15404,N_14954,N_14598);
or U15405 (N_15405,N_14516,N_14608);
nor U15406 (N_15406,N_14822,N_14901);
or U15407 (N_15407,N_14597,N_14782);
and U15408 (N_15408,N_14995,N_14671);
nand U15409 (N_15409,N_14929,N_14562);
nand U15410 (N_15410,N_14942,N_14818);
nor U15411 (N_15411,N_14878,N_14595);
nand U15412 (N_15412,N_14527,N_14525);
nand U15413 (N_15413,N_14616,N_14604);
nand U15414 (N_15414,N_14717,N_14931);
and U15415 (N_15415,N_14890,N_14573);
nor U15416 (N_15416,N_14537,N_14878);
xor U15417 (N_15417,N_14675,N_14971);
nor U15418 (N_15418,N_14970,N_14629);
nand U15419 (N_15419,N_14515,N_14999);
nand U15420 (N_15420,N_14907,N_14746);
xnor U15421 (N_15421,N_14832,N_14875);
or U15422 (N_15422,N_14702,N_14756);
xor U15423 (N_15423,N_14524,N_14673);
nand U15424 (N_15424,N_14900,N_14599);
nor U15425 (N_15425,N_14876,N_14626);
nor U15426 (N_15426,N_14634,N_14797);
and U15427 (N_15427,N_14580,N_14707);
nand U15428 (N_15428,N_14609,N_14648);
xor U15429 (N_15429,N_14527,N_14636);
or U15430 (N_15430,N_14622,N_14530);
xor U15431 (N_15431,N_14546,N_14945);
or U15432 (N_15432,N_14911,N_14776);
nand U15433 (N_15433,N_14794,N_14567);
or U15434 (N_15434,N_14600,N_14882);
nand U15435 (N_15435,N_14563,N_14907);
and U15436 (N_15436,N_14603,N_14883);
xnor U15437 (N_15437,N_14907,N_14899);
nor U15438 (N_15438,N_14686,N_14537);
and U15439 (N_15439,N_14793,N_14505);
nor U15440 (N_15440,N_14609,N_14667);
nor U15441 (N_15441,N_14622,N_14670);
nand U15442 (N_15442,N_14858,N_14859);
nor U15443 (N_15443,N_14548,N_14926);
xor U15444 (N_15444,N_14540,N_14550);
xnor U15445 (N_15445,N_14886,N_14760);
xnor U15446 (N_15446,N_14503,N_14941);
or U15447 (N_15447,N_14845,N_14769);
nor U15448 (N_15448,N_14964,N_14819);
nand U15449 (N_15449,N_14625,N_14895);
nand U15450 (N_15450,N_14988,N_14857);
nor U15451 (N_15451,N_14841,N_14748);
and U15452 (N_15452,N_14970,N_14813);
or U15453 (N_15453,N_14899,N_14970);
xor U15454 (N_15454,N_14878,N_14590);
and U15455 (N_15455,N_14531,N_14991);
nor U15456 (N_15456,N_14582,N_14522);
and U15457 (N_15457,N_14758,N_14689);
nand U15458 (N_15458,N_14798,N_14926);
and U15459 (N_15459,N_14917,N_14560);
nand U15460 (N_15460,N_14516,N_14685);
and U15461 (N_15461,N_14788,N_14933);
or U15462 (N_15462,N_14702,N_14736);
nor U15463 (N_15463,N_14814,N_14870);
nor U15464 (N_15464,N_14908,N_14897);
and U15465 (N_15465,N_14910,N_14676);
and U15466 (N_15466,N_14671,N_14933);
and U15467 (N_15467,N_14699,N_14660);
xnor U15468 (N_15468,N_14822,N_14790);
nand U15469 (N_15469,N_14742,N_14880);
xor U15470 (N_15470,N_14621,N_14547);
or U15471 (N_15471,N_14607,N_14513);
and U15472 (N_15472,N_14644,N_14831);
nand U15473 (N_15473,N_14641,N_14974);
nand U15474 (N_15474,N_14932,N_14794);
or U15475 (N_15475,N_14795,N_14957);
nor U15476 (N_15476,N_14742,N_14592);
and U15477 (N_15477,N_14649,N_14561);
xnor U15478 (N_15478,N_14966,N_14579);
xnor U15479 (N_15479,N_14797,N_14922);
or U15480 (N_15480,N_14582,N_14998);
xnor U15481 (N_15481,N_14990,N_14968);
or U15482 (N_15482,N_14986,N_14838);
nor U15483 (N_15483,N_14790,N_14731);
or U15484 (N_15484,N_14979,N_14727);
and U15485 (N_15485,N_14818,N_14739);
nand U15486 (N_15486,N_14976,N_14913);
xor U15487 (N_15487,N_14871,N_14688);
and U15488 (N_15488,N_14767,N_14929);
nor U15489 (N_15489,N_14805,N_14751);
and U15490 (N_15490,N_14531,N_14627);
or U15491 (N_15491,N_14528,N_14692);
nor U15492 (N_15492,N_14620,N_14829);
or U15493 (N_15493,N_14939,N_14555);
nor U15494 (N_15494,N_14537,N_14899);
or U15495 (N_15495,N_14662,N_14583);
and U15496 (N_15496,N_14723,N_14769);
or U15497 (N_15497,N_14602,N_14909);
or U15498 (N_15498,N_14906,N_14923);
nor U15499 (N_15499,N_14599,N_14731);
nand U15500 (N_15500,N_15057,N_15327);
nor U15501 (N_15501,N_15390,N_15141);
nor U15502 (N_15502,N_15249,N_15181);
nor U15503 (N_15503,N_15040,N_15140);
or U15504 (N_15504,N_15029,N_15497);
nor U15505 (N_15505,N_15469,N_15100);
or U15506 (N_15506,N_15190,N_15160);
nand U15507 (N_15507,N_15232,N_15371);
and U15508 (N_15508,N_15191,N_15300);
nand U15509 (N_15509,N_15401,N_15094);
nor U15510 (N_15510,N_15086,N_15240);
or U15511 (N_15511,N_15087,N_15070);
and U15512 (N_15512,N_15247,N_15259);
nand U15513 (N_15513,N_15097,N_15061);
or U15514 (N_15514,N_15293,N_15216);
and U15515 (N_15515,N_15143,N_15137);
xnor U15516 (N_15516,N_15149,N_15256);
and U15517 (N_15517,N_15051,N_15235);
xnor U15518 (N_15518,N_15242,N_15276);
xnor U15519 (N_15519,N_15020,N_15344);
and U15520 (N_15520,N_15136,N_15330);
nor U15521 (N_15521,N_15313,N_15208);
xnor U15522 (N_15522,N_15386,N_15387);
nor U15523 (N_15523,N_15161,N_15021);
xor U15524 (N_15524,N_15362,N_15227);
nor U15525 (N_15525,N_15119,N_15305);
or U15526 (N_15526,N_15066,N_15373);
xnor U15527 (N_15527,N_15289,N_15267);
and U15528 (N_15528,N_15319,N_15287);
nor U15529 (N_15529,N_15328,N_15432);
xnor U15530 (N_15530,N_15003,N_15367);
or U15531 (N_15531,N_15494,N_15151);
nand U15532 (N_15532,N_15467,N_15063);
xnor U15533 (N_15533,N_15203,N_15303);
xnor U15534 (N_15534,N_15439,N_15171);
nor U15535 (N_15535,N_15333,N_15117);
nor U15536 (N_15536,N_15134,N_15340);
nand U15537 (N_15537,N_15363,N_15298);
nor U15538 (N_15538,N_15355,N_15446);
and U15539 (N_15539,N_15343,N_15156);
nand U15540 (N_15540,N_15316,N_15164);
nand U15541 (N_15541,N_15039,N_15102);
nand U15542 (N_15542,N_15459,N_15427);
xnor U15543 (N_15543,N_15351,N_15440);
and U15544 (N_15544,N_15348,N_15412);
and U15545 (N_15545,N_15280,N_15286);
and U15546 (N_15546,N_15475,N_15153);
xor U15547 (N_15547,N_15205,N_15483);
xnor U15548 (N_15548,N_15217,N_15488);
or U15549 (N_15549,N_15194,N_15179);
xnor U15550 (N_15550,N_15168,N_15248);
or U15551 (N_15551,N_15172,N_15499);
nand U15552 (N_15552,N_15402,N_15449);
xor U15553 (N_15553,N_15368,N_15487);
nor U15554 (N_15554,N_15109,N_15255);
or U15555 (N_15555,N_15283,N_15321);
or U15556 (N_15556,N_15346,N_15403);
xnor U15557 (N_15557,N_15049,N_15491);
xor U15558 (N_15558,N_15000,N_15007);
or U15559 (N_15559,N_15126,N_15473);
and U15560 (N_15560,N_15031,N_15133);
nand U15561 (N_15561,N_15043,N_15393);
nor U15562 (N_15562,N_15498,N_15442);
nand U15563 (N_15563,N_15139,N_15106);
nand U15564 (N_15564,N_15050,N_15092);
nand U15565 (N_15565,N_15324,N_15381);
and U15566 (N_15566,N_15204,N_15400);
nor U15567 (N_15567,N_15329,N_15273);
nor U15568 (N_15568,N_15493,N_15023);
and U15569 (N_15569,N_15269,N_15476);
nand U15570 (N_15570,N_15365,N_15350);
or U15571 (N_15571,N_15192,N_15444);
nor U15572 (N_15572,N_15067,N_15101);
nand U15573 (N_15573,N_15048,N_15285);
nor U15574 (N_15574,N_15076,N_15001);
xor U15575 (N_15575,N_15122,N_15214);
or U15576 (N_15576,N_15434,N_15155);
or U15577 (N_15577,N_15486,N_15452);
xnor U15578 (N_15578,N_15152,N_15489);
nor U15579 (N_15579,N_15364,N_15099);
nand U15580 (N_15580,N_15047,N_15291);
xnor U15581 (N_15581,N_15084,N_15166);
or U15582 (N_15582,N_15068,N_15071);
nand U15583 (N_15583,N_15098,N_15175);
or U15584 (N_15584,N_15404,N_15073);
nor U15585 (N_15585,N_15124,N_15022);
or U15586 (N_15586,N_15264,N_15394);
and U15587 (N_15587,N_15339,N_15210);
xor U15588 (N_15588,N_15301,N_15399);
nor U15589 (N_15589,N_15145,N_15197);
xor U15590 (N_15590,N_15461,N_15443);
and U15591 (N_15591,N_15081,N_15104);
nor U15592 (N_15592,N_15279,N_15238);
nand U15593 (N_15593,N_15123,N_15079);
xnor U15594 (N_15594,N_15195,N_15025);
and U15595 (N_15595,N_15306,N_15323);
nor U15596 (N_15596,N_15069,N_15481);
xor U15597 (N_15597,N_15221,N_15460);
and U15598 (N_15598,N_15018,N_15308);
or U15599 (N_15599,N_15093,N_15392);
nand U15600 (N_15600,N_15370,N_15389);
and U15601 (N_15601,N_15448,N_15230);
xor U15602 (N_15602,N_15014,N_15163);
and U15603 (N_15603,N_15055,N_15085);
and U15604 (N_15604,N_15431,N_15418);
xor U15605 (N_15605,N_15275,N_15028);
or U15606 (N_15606,N_15215,N_15095);
nor U15607 (N_15607,N_15184,N_15125);
or U15608 (N_15608,N_15035,N_15015);
and U15609 (N_15609,N_15356,N_15245);
xnor U15610 (N_15610,N_15118,N_15397);
nand U15611 (N_15611,N_15395,N_15360);
or U15612 (N_15612,N_15244,N_15024);
nor U15613 (N_15613,N_15490,N_15121);
and U15614 (N_15614,N_15077,N_15262);
xnor U15615 (N_15615,N_15435,N_15458);
nor U15616 (N_15616,N_15228,N_15385);
nor U15617 (N_15617,N_15246,N_15016);
and U15618 (N_15618,N_15429,N_15380);
nand U15619 (N_15619,N_15496,N_15229);
xor U15620 (N_15620,N_15417,N_15284);
and U15621 (N_15621,N_15189,N_15292);
and U15622 (N_15622,N_15222,N_15359);
or U15623 (N_15623,N_15254,N_15008);
nand U15624 (N_15624,N_15445,N_15456);
and U15625 (N_15625,N_15416,N_15302);
nand U15626 (N_15626,N_15271,N_15377);
xnor U15627 (N_15627,N_15422,N_15480);
xnor U15628 (N_15628,N_15470,N_15052);
xnor U15629 (N_15629,N_15388,N_15193);
nand U15630 (N_15630,N_15142,N_15318);
nand U15631 (N_15631,N_15423,N_15369);
and U15632 (N_15632,N_15110,N_15220);
or U15633 (N_15633,N_15144,N_15114);
xor U15634 (N_15634,N_15492,N_15041);
xnor U15635 (N_15635,N_15354,N_15266);
or U15636 (N_15636,N_15309,N_15006);
nor U15637 (N_15637,N_15116,N_15111);
nor U15638 (N_15638,N_15234,N_15132);
xnor U15639 (N_15639,N_15382,N_15338);
xnor U15640 (N_15640,N_15297,N_15415);
xnor U15641 (N_15641,N_15185,N_15211);
and U15642 (N_15642,N_15105,N_15304);
or U15643 (N_15643,N_15011,N_15180);
and U15644 (N_15644,N_15378,N_15294);
or U15645 (N_15645,N_15436,N_15188);
xor U15646 (N_15646,N_15201,N_15322);
nand U15647 (N_15647,N_15361,N_15233);
nor U15648 (N_15648,N_15146,N_15037);
nand U15649 (N_15649,N_15374,N_15103);
or U15650 (N_15650,N_15078,N_15209);
xor U15651 (N_15651,N_15251,N_15463);
nand U15652 (N_15652,N_15157,N_15383);
nand U15653 (N_15653,N_15075,N_15257);
and U15654 (N_15654,N_15224,N_15046);
nor U15655 (N_15655,N_15112,N_15465);
or U15656 (N_15656,N_15150,N_15128);
nand U15657 (N_15657,N_15162,N_15182);
and U15658 (N_15658,N_15282,N_15464);
and U15659 (N_15659,N_15058,N_15384);
nor U15660 (N_15660,N_15457,N_15196);
xor U15661 (N_15661,N_15263,N_15186);
xnor U15662 (N_15662,N_15372,N_15495);
or U15663 (N_15663,N_15411,N_15425);
and U15664 (N_15664,N_15223,N_15455);
and U15665 (N_15665,N_15310,N_15409);
nand U15666 (N_15666,N_15226,N_15213);
nor U15667 (N_15667,N_15341,N_15472);
nor U15668 (N_15668,N_15038,N_15207);
xnor U15669 (N_15669,N_15349,N_15199);
nand U15670 (N_15670,N_15054,N_15082);
nor U15671 (N_15671,N_15258,N_15295);
nor U15672 (N_15672,N_15345,N_15420);
nor U15673 (N_15673,N_15010,N_15060);
and U15674 (N_15674,N_15120,N_15113);
nand U15675 (N_15675,N_15200,N_15438);
and U15676 (N_15676,N_15278,N_15004);
nand U15677 (N_15677,N_15272,N_15296);
and U15678 (N_15678,N_15342,N_15253);
and U15679 (N_15679,N_15288,N_15270);
nand U15680 (N_15680,N_15260,N_15331);
and U15681 (N_15681,N_15375,N_15053);
or U15682 (N_15682,N_15312,N_15017);
nor U15683 (N_15683,N_15379,N_15290);
or U15684 (N_15684,N_15468,N_15454);
nand U15685 (N_15685,N_15090,N_15072);
nand U15686 (N_15686,N_15419,N_15236);
or U15687 (N_15687,N_15413,N_15414);
or U15688 (N_15688,N_15332,N_15453);
or U15689 (N_15689,N_15410,N_15398);
xor U15690 (N_15690,N_15437,N_15315);
nand U15691 (N_15691,N_15281,N_15243);
or U15692 (N_15692,N_15042,N_15034);
and U15693 (N_15693,N_15219,N_15135);
or U15694 (N_15694,N_15074,N_15013);
or U15695 (N_15695,N_15430,N_15408);
and U15696 (N_15696,N_15441,N_15177);
and U15697 (N_15697,N_15165,N_15424);
or U15698 (N_15698,N_15334,N_15130);
and U15699 (N_15699,N_15426,N_15127);
or U15700 (N_15700,N_15148,N_15129);
or U15701 (N_15701,N_15406,N_15059);
or U15702 (N_15702,N_15108,N_15352);
and U15703 (N_15703,N_15484,N_15080);
and U15704 (N_15704,N_15336,N_15187);
or U15705 (N_15705,N_15450,N_15032);
and U15706 (N_15706,N_15250,N_15482);
xor U15707 (N_15707,N_15169,N_15391);
and U15708 (N_15708,N_15471,N_15252);
nand U15709 (N_15709,N_15451,N_15198);
xnor U15710 (N_15710,N_15178,N_15159);
and U15711 (N_15711,N_15147,N_15237);
and U15712 (N_15712,N_15033,N_15056);
or U15713 (N_15713,N_15268,N_15009);
nand U15714 (N_15714,N_15005,N_15261);
or U15715 (N_15715,N_15096,N_15447);
and U15716 (N_15716,N_15421,N_15407);
or U15717 (N_15717,N_15299,N_15167);
nor U15718 (N_15718,N_15091,N_15019);
or U15719 (N_15719,N_15320,N_15478);
nand U15720 (N_15720,N_15307,N_15030);
and U15721 (N_15721,N_15376,N_15138);
or U15722 (N_15722,N_15474,N_15335);
nor U15723 (N_15723,N_15089,N_15206);
nor U15724 (N_15724,N_15154,N_15107);
xnor U15725 (N_15725,N_15347,N_15174);
xnor U15726 (N_15726,N_15045,N_15325);
nor U15727 (N_15727,N_15183,N_15466);
nor U15728 (N_15728,N_15012,N_15170);
nand U15729 (N_15729,N_15231,N_15002);
or U15730 (N_15730,N_15088,N_15366);
and U15731 (N_15731,N_15317,N_15311);
xor U15732 (N_15732,N_15158,N_15212);
xnor U15733 (N_15733,N_15173,N_15044);
or U15734 (N_15734,N_15358,N_15062);
nor U15735 (N_15735,N_15277,N_15083);
nor U15736 (N_15736,N_15353,N_15462);
or U15737 (N_15737,N_15218,N_15176);
xnor U15738 (N_15738,N_15274,N_15241);
or U15739 (N_15739,N_15027,N_15428);
or U15740 (N_15740,N_15479,N_15485);
nand U15741 (N_15741,N_15326,N_15225);
nand U15742 (N_15742,N_15314,N_15131);
and U15743 (N_15743,N_15433,N_15026);
and U15744 (N_15744,N_15477,N_15115);
xor U15745 (N_15745,N_15357,N_15065);
and U15746 (N_15746,N_15265,N_15064);
nor U15747 (N_15747,N_15396,N_15337);
and U15748 (N_15748,N_15405,N_15239);
nor U15749 (N_15749,N_15036,N_15202);
and U15750 (N_15750,N_15474,N_15247);
xor U15751 (N_15751,N_15106,N_15346);
and U15752 (N_15752,N_15103,N_15090);
or U15753 (N_15753,N_15196,N_15062);
nand U15754 (N_15754,N_15444,N_15038);
nand U15755 (N_15755,N_15154,N_15209);
or U15756 (N_15756,N_15468,N_15071);
xnor U15757 (N_15757,N_15486,N_15398);
xor U15758 (N_15758,N_15101,N_15383);
xnor U15759 (N_15759,N_15306,N_15403);
nor U15760 (N_15760,N_15305,N_15299);
xor U15761 (N_15761,N_15167,N_15343);
or U15762 (N_15762,N_15468,N_15065);
or U15763 (N_15763,N_15051,N_15307);
nand U15764 (N_15764,N_15190,N_15067);
nor U15765 (N_15765,N_15026,N_15387);
xnor U15766 (N_15766,N_15073,N_15488);
or U15767 (N_15767,N_15124,N_15391);
xor U15768 (N_15768,N_15177,N_15373);
nand U15769 (N_15769,N_15453,N_15033);
or U15770 (N_15770,N_15134,N_15220);
nand U15771 (N_15771,N_15445,N_15307);
nor U15772 (N_15772,N_15208,N_15445);
and U15773 (N_15773,N_15088,N_15377);
nor U15774 (N_15774,N_15393,N_15026);
nand U15775 (N_15775,N_15236,N_15073);
nand U15776 (N_15776,N_15006,N_15431);
and U15777 (N_15777,N_15143,N_15224);
xnor U15778 (N_15778,N_15202,N_15288);
or U15779 (N_15779,N_15198,N_15083);
nor U15780 (N_15780,N_15429,N_15435);
nor U15781 (N_15781,N_15036,N_15482);
and U15782 (N_15782,N_15377,N_15105);
nor U15783 (N_15783,N_15191,N_15125);
nor U15784 (N_15784,N_15174,N_15304);
and U15785 (N_15785,N_15211,N_15261);
nor U15786 (N_15786,N_15268,N_15298);
or U15787 (N_15787,N_15313,N_15135);
nand U15788 (N_15788,N_15222,N_15290);
and U15789 (N_15789,N_15390,N_15422);
or U15790 (N_15790,N_15359,N_15068);
or U15791 (N_15791,N_15414,N_15167);
nor U15792 (N_15792,N_15309,N_15001);
nand U15793 (N_15793,N_15412,N_15318);
xor U15794 (N_15794,N_15130,N_15441);
xnor U15795 (N_15795,N_15309,N_15131);
nand U15796 (N_15796,N_15294,N_15158);
and U15797 (N_15797,N_15337,N_15044);
nand U15798 (N_15798,N_15053,N_15281);
or U15799 (N_15799,N_15398,N_15214);
nor U15800 (N_15800,N_15049,N_15302);
xnor U15801 (N_15801,N_15016,N_15259);
xor U15802 (N_15802,N_15246,N_15471);
and U15803 (N_15803,N_15034,N_15145);
or U15804 (N_15804,N_15050,N_15341);
or U15805 (N_15805,N_15128,N_15209);
nand U15806 (N_15806,N_15309,N_15276);
and U15807 (N_15807,N_15306,N_15071);
or U15808 (N_15808,N_15161,N_15389);
nand U15809 (N_15809,N_15210,N_15252);
or U15810 (N_15810,N_15327,N_15203);
or U15811 (N_15811,N_15492,N_15060);
nand U15812 (N_15812,N_15324,N_15417);
and U15813 (N_15813,N_15379,N_15293);
and U15814 (N_15814,N_15234,N_15256);
nand U15815 (N_15815,N_15379,N_15088);
nand U15816 (N_15816,N_15423,N_15375);
nor U15817 (N_15817,N_15268,N_15063);
nor U15818 (N_15818,N_15465,N_15082);
and U15819 (N_15819,N_15029,N_15231);
nor U15820 (N_15820,N_15024,N_15007);
xor U15821 (N_15821,N_15052,N_15391);
or U15822 (N_15822,N_15319,N_15164);
nand U15823 (N_15823,N_15142,N_15174);
nand U15824 (N_15824,N_15235,N_15118);
xor U15825 (N_15825,N_15248,N_15402);
nand U15826 (N_15826,N_15451,N_15086);
or U15827 (N_15827,N_15379,N_15030);
or U15828 (N_15828,N_15011,N_15089);
and U15829 (N_15829,N_15203,N_15000);
nand U15830 (N_15830,N_15141,N_15345);
and U15831 (N_15831,N_15254,N_15192);
and U15832 (N_15832,N_15249,N_15358);
nor U15833 (N_15833,N_15485,N_15021);
and U15834 (N_15834,N_15245,N_15270);
nor U15835 (N_15835,N_15273,N_15181);
nand U15836 (N_15836,N_15352,N_15075);
nor U15837 (N_15837,N_15434,N_15074);
or U15838 (N_15838,N_15202,N_15274);
or U15839 (N_15839,N_15475,N_15432);
or U15840 (N_15840,N_15194,N_15299);
or U15841 (N_15841,N_15382,N_15381);
xor U15842 (N_15842,N_15216,N_15124);
xor U15843 (N_15843,N_15491,N_15328);
nor U15844 (N_15844,N_15431,N_15306);
nor U15845 (N_15845,N_15408,N_15462);
nor U15846 (N_15846,N_15048,N_15090);
nand U15847 (N_15847,N_15210,N_15290);
xnor U15848 (N_15848,N_15366,N_15296);
nor U15849 (N_15849,N_15369,N_15037);
nor U15850 (N_15850,N_15260,N_15229);
nand U15851 (N_15851,N_15242,N_15458);
or U15852 (N_15852,N_15437,N_15413);
nor U15853 (N_15853,N_15244,N_15228);
or U15854 (N_15854,N_15135,N_15029);
and U15855 (N_15855,N_15131,N_15339);
and U15856 (N_15856,N_15250,N_15214);
xor U15857 (N_15857,N_15207,N_15298);
and U15858 (N_15858,N_15137,N_15151);
xnor U15859 (N_15859,N_15036,N_15059);
xor U15860 (N_15860,N_15057,N_15307);
xor U15861 (N_15861,N_15494,N_15115);
and U15862 (N_15862,N_15338,N_15286);
nor U15863 (N_15863,N_15148,N_15330);
nor U15864 (N_15864,N_15058,N_15304);
and U15865 (N_15865,N_15170,N_15471);
or U15866 (N_15866,N_15038,N_15012);
xnor U15867 (N_15867,N_15237,N_15016);
or U15868 (N_15868,N_15112,N_15184);
and U15869 (N_15869,N_15445,N_15463);
nor U15870 (N_15870,N_15331,N_15355);
and U15871 (N_15871,N_15453,N_15394);
or U15872 (N_15872,N_15006,N_15015);
and U15873 (N_15873,N_15388,N_15238);
and U15874 (N_15874,N_15264,N_15231);
nor U15875 (N_15875,N_15015,N_15004);
nor U15876 (N_15876,N_15202,N_15491);
xor U15877 (N_15877,N_15256,N_15033);
or U15878 (N_15878,N_15354,N_15450);
nor U15879 (N_15879,N_15471,N_15457);
nand U15880 (N_15880,N_15295,N_15155);
and U15881 (N_15881,N_15453,N_15343);
xor U15882 (N_15882,N_15439,N_15196);
nand U15883 (N_15883,N_15497,N_15445);
and U15884 (N_15884,N_15244,N_15121);
nand U15885 (N_15885,N_15415,N_15429);
xor U15886 (N_15886,N_15451,N_15306);
nand U15887 (N_15887,N_15219,N_15080);
nor U15888 (N_15888,N_15396,N_15002);
nor U15889 (N_15889,N_15210,N_15461);
or U15890 (N_15890,N_15094,N_15291);
nand U15891 (N_15891,N_15028,N_15411);
xnor U15892 (N_15892,N_15300,N_15246);
and U15893 (N_15893,N_15099,N_15084);
or U15894 (N_15894,N_15395,N_15069);
and U15895 (N_15895,N_15103,N_15182);
or U15896 (N_15896,N_15350,N_15212);
or U15897 (N_15897,N_15036,N_15219);
nand U15898 (N_15898,N_15058,N_15146);
nand U15899 (N_15899,N_15169,N_15197);
nand U15900 (N_15900,N_15172,N_15480);
nor U15901 (N_15901,N_15318,N_15399);
nand U15902 (N_15902,N_15107,N_15015);
or U15903 (N_15903,N_15123,N_15467);
and U15904 (N_15904,N_15039,N_15192);
or U15905 (N_15905,N_15371,N_15115);
nor U15906 (N_15906,N_15007,N_15233);
xnor U15907 (N_15907,N_15473,N_15193);
nor U15908 (N_15908,N_15166,N_15013);
or U15909 (N_15909,N_15191,N_15244);
or U15910 (N_15910,N_15204,N_15263);
or U15911 (N_15911,N_15230,N_15330);
nor U15912 (N_15912,N_15390,N_15163);
xnor U15913 (N_15913,N_15382,N_15035);
nand U15914 (N_15914,N_15043,N_15211);
nor U15915 (N_15915,N_15399,N_15205);
xnor U15916 (N_15916,N_15244,N_15252);
and U15917 (N_15917,N_15449,N_15018);
nor U15918 (N_15918,N_15393,N_15150);
and U15919 (N_15919,N_15335,N_15480);
nor U15920 (N_15920,N_15442,N_15348);
xnor U15921 (N_15921,N_15253,N_15289);
and U15922 (N_15922,N_15153,N_15371);
and U15923 (N_15923,N_15127,N_15300);
or U15924 (N_15924,N_15365,N_15278);
and U15925 (N_15925,N_15284,N_15321);
and U15926 (N_15926,N_15171,N_15151);
nand U15927 (N_15927,N_15239,N_15134);
nor U15928 (N_15928,N_15481,N_15065);
xnor U15929 (N_15929,N_15049,N_15055);
and U15930 (N_15930,N_15433,N_15194);
or U15931 (N_15931,N_15202,N_15418);
or U15932 (N_15932,N_15416,N_15447);
nand U15933 (N_15933,N_15447,N_15458);
or U15934 (N_15934,N_15112,N_15376);
xor U15935 (N_15935,N_15061,N_15003);
or U15936 (N_15936,N_15274,N_15352);
or U15937 (N_15937,N_15238,N_15040);
nand U15938 (N_15938,N_15131,N_15262);
xnor U15939 (N_15939,N_15165,N_15022);
xnor U15940 (N_15940,N_15080,N_15474);
xnor U15941 (N_15941,N_15034,N_15499);
or U15942 (N_15942,N_15279,N_15150);
nand U15943 (N_15943,N_15353,N_15425);
nand U15944 (N_15944,N_15444,N_15384);
and U15945 (N_15945,N_15013,N_15113);
or U15946 (N_15946,N_15264,N_15049);
or U15947 (N_15947,N_15212,N_15376);
nand U15948 (N_15948,N_15466,N_15192);
nand U15949 (N_15949,N_15196,N_15253);
xor U15950 (N_15950,N_15482,N_15498);
xor U15951 (N_15951,N_15200,N_15144);
and U15952 (N_15952,N_15006,N_15146);
or U15953 (N_15953,N_15174,N_15104);
xnor U15954 (N_15954,N_15323,N_15038);
and U15955 (N_15955,N_15195,N_15342);
and U15956 (N_15956,N_15184,N_15068);
nor U15957 (N_15957,N_15267,N_15174);
and U15958 (N_15958,N_15462,N_15405);
and U15959 (N_15959,N_15037,N_15127);
and U15960 (N_15960,N_15296,N_15146);
xor U15961 (N_15961,N_15295,N_15107);
and U15962 (N_15962,N_15476,N_15139);
or U15963 (N_15963,N_15368,N_15022);
xor U15964 (N_15964,N_15233,N_15294);
nor U15965 (N_15965,N_15385,N_15066);
or U15966 (N_15966,N_15224,N_15319);
or U15967 (N_15967,N_15418,N_15287);
or U15968 (N_15968,N_15336,N_15165);
or U15969 (N_15969,N_15478,N_15246);
and U15970 (N_15970,N_15356,N_15147);
nand U15971 (N_15971,N_15347,N_15282);
nand U15972 (N_15972,N_15467,N_15310);
and U15973 (N_15973,N_15425,N_15090);
xor U15974 (N_15974,N_15256,N_15491);
nand U15975 (N_15975,N_15400,N_15174);
or U15976 (N_15976,N_15431,N_15463);
xor U15977 (N_15977,N_15319,N_15043);
and U15978 (N_15978,N_15448,N_15342);
nand U15979 (N_15979,N_15435,N_15467);
nand U15980 (N_15980,N_15192,N_15201);
or U15981 (N_15981,N_15201,N_15311);
and U15982 (N_15982,N_15406,N_15107);
nand U15983 (N_15983,N_15188,N_15050);
xor U15984 (N_15984,N_15418,N_15496);
and U15985 (N_15985,N_15168,N_15188);
xnor U15986 (N_15986,N_15024,N_15288);
nand U15987 (N_15987,N_15249,N_15025);
or U15988 (N_15988,N_15070,N_15054);
xor U15989 (N_15989,N_15298,N_15418);
or U15990 (N_15990,N_15233,N_15048);
or U15991 (N_15991,N_15243,N_15391);
nor U15992 (N_15992,N_15323,N_15449);
and U15993 (N_15993,N_15254,N_15329);
or U15994 (N_15994,N_15344,N_15207);
and U15995 (N_15995,N_15227,N_15139);
xor U15996 (N_15996,N_15225,N_15282);
and U15997 (N_15997,N_15126,N_15425);
nand U15998 (N_15998,N_15205,N_15444);
nand U15999 (N_15999,N_15103,N_15168);
nand U16000 (N_16000,N_15751,N_15793);
nand U16001 (N_16001,N_15593,N_15948);
xnor U16002 (N_16002,N_15997,N_15781);
and U16003 (N_16003,N_15723,N_15848);
nand U16004 (N_16004,N_15621,N_15553);
or U16005 (N_16005,N_15810,N_15919);
nor U16006 (N_16006,N_15992,N_15841);
nand U16007 (N_16007,N_15551,N_15645);
and U16008 (N_16008,N_15705,N_15995);
and U16009 (N_16009,N_15935,N_15986);
or U16010 (N_16010,N_15687,N_15649);
xor U16011 (N_16011,N_15929,N_15719);
and U16012 (N_16012,N_15637,N_15753);
and U16013 (N_16013,N_15557,N_15655);
nor U16014 (N_16014,N_15767,N_15511);
or U16015 (N_16015,N_15825,N_15913);
xor U16016 (N_16016,N_15534,N_15897);
nor U16017 (N_16017,N_15692,N_15900);
xnor U16018 (N_16018,N_15567,N_15581);
xor U16019 (N_16019,N_15710,N_15860);
nor U16020 (N_16020,N_15609,N_15506);
xor U16021 (N_16021,N_15693,N_15709);
or U16022 (N_16022,N_15875,N_15790);
and U16023 (N_16023,N_15616,N_15777);
nor U16024 (N_16024,N_15749,N_15894);
nand U16025 (N_16025,N_15839,N_15982);
xnor U16026 (N_16026,N_15940,N_15836);
nor U16027 (N_16027,N_15826,N_15611);
and U16028 (N_16028,N_15872,N_15961);
xor U16029 (N_16029,N_15548,N_15617);
nor U16030 (N_16030,N_15726,N_15656);
or U16031 (N_16031,N_15519,N_15559);
xnor U16032 (N_16032,N_15994,N_15625);
nand U16033 (N_16033,N_15996,N_15973);
xnor U16034 (N_16034,N_15689,N_15500);
nand U16035 (N_16035,N_15993,N_15846);
nor U16036 (N_16036,N_15729,N_15772);
nor U16037 (N_16037,N_15960,N_15647);
xor U16038 (N_16038,N_15515,N_15967);
and U16039 (N_16039,N_15759,N_15804);
nor U16040 (N_16040,N_15914,N_15654);
or U16041 (N_16041,N_15785,N_15657);
xnor U16042 (N_16042,N_15981,N_15761);
nand U16043 (N_16043,N_15901,N_15861);
and U16044 (N_16044,N_15776,N_15596);
or U16045 (N_16045,N_15849,N_15983);
xnor U16046 (N_16046,N_15651,N_15924);
or U16047 (N_16047,N_15818,N_15667);
nand U16048 (N_16048,N_15912,N_15533);
xnor U16049 (N_16049,N_15583,N_15957);
xor U16050 (N_16050,N_15895,N_15661);
xnor U16051 (N_16051,N_15678,N_15739);
and U16052 (N_16052,N_15873,N_15813);
xor U16053 (N_16053,N_15535,N_15779);
and U16054 (N_16054,N_15505,N_15757);
or U16055 (N_16055,N_15544,N_15816);
nor U16056 (N_16056,N_15707,N_15613);
nor U16057 (N_16057,N_15720,N_15918);
xnor U16058 (N_16058,N_15903,N_15815);
and U16059 (N_16059,N_15740,N_15629);
and U16060 (N_16060,N_15568,N_15564);
nand U16061 (N_16061,N_15928,N_15831);
nand U16062 (N_16062,N_15532,N_15788);
xnor U16063 (N_16063,N_15669,N_15812);
and U16064 (N_16064,N_15646,N_15868);
xnor U16065 (N_16065,N_15938,N_15561);
and U16066 (N_16066,N_15999,N_15843);
nand U16067 (N_16067,N_15712,N_15699);
nor U16068 (N_16068,N_15905,N_15955);
and U16069 (N_16069,N_15612,N_15560);
nand U16070 (N_16070,N_15630,N_15518);
xor U16071 (N_16071,N_15576,N_15507);
nor U16072 (N_16072,N_15852,N_15586);
xor U16073 (N_16073,N_15664,N_15605);
xor U16074 (N_16074,N_15536,N_15700);
or U16075 (N_16075,N_15768,N_15943);
nand U16076 (N_16076,N_15744,N_15618);
xor U16077 (N_16077,N_15563,N_15789);
nand U16078 (N_16078,N_15603,N_15668);
nor U16079 (N_16079,N_15892,N_15545);
or U16080 (N_16080,N_15811,N_15610);
nand U16081 (N_16081,N_15771,N_15604);
and U16082 (N_16082,N_15711,N_15975);
nand U16083 (N_16083,N_15676,N_15514);
xnor U16084 (N_16084,N_15595,N_15909);
nand U16085 (N_16085,N_15716,N_15525);
nor U16086 (N_16086,N_15939,N_15896);
xor U16087 (N_16087,N_15856,N_15837);
and U16088 (N_16088,N_15835,N_15864);
and U16089 (N_16089,N_15934,N_15965);
or U16090 (N_16090,N_15732,N_15631);
xnor U16091 (N_16091,N_15990,N_15888);
and U16092 (N_16092,N_15585,N_15643);
and U16093 (N_16093,N_15708,N_15638);
or U16094 (N_16094,N_15869,N_15589);
nor U16095 (N_16095,N_15718,N_15800);
nor U16096 (N_16096,N_15794,N_15898);
xnor U16097 (N_16097,N_15956,N_15877);
xnor U16098 (N_16098,N_15714,N_15778);
xor U16099 (N_16099,N_15865,N_15642);
xor U16100 (N_16100,N_15902,N_15842);
or U16101 (N_16101,N_15874,N_15802);
and U16102 (N_16102,N_15683,N_15921);
nand U16103 (N_16103,N_15787,N_15893);
and U16104 (N_16104,N_15733,N_15819);
nor U16105 (N_16105,N_15857,N_15552);
nand U16106 (N_16106,N_15773,N_15660);
xor U16107 (N_16107,N_15575,N_15666);
nor U16108 (N_16108,N_15926,N_15858);
nor U16109 (N_16109,N_15847,N_15809);
or U16110 (N_16110,N_15704,N_15952);
nor U16111 (N_16111,N_15522,N_15915);
nand U16112 (N_16112,N_15731,N_15976);
nand U16113 (N_16113,N_15597,N_15962);
or U16114 (N_16114,N_15795,N_15725);
nor U16115 (N_16115,N_15702,N_15820);
and U16116 (N_16116,N_15531,N_15520);
nor U16117 (N_16117,N_15538,N_15906);
and U16118 (N_16118,N_15598,N_15946);
xnor U16119 (N_16119,N_15556,N_15754);
or U16120 (N_16120,N_15743,N_15608);
nand U16121 (N_16121,N_15622,N_15969);
or U16122 (N_16122,N_15572,N_15959);
xor U16123 (N_16123,N_15587,N_15673);
and U16124 (N_16124,N_15659,N_15882);
nand U16125 (N_16125,N_15584,N_15991);
and U16126 (N_16126,N_15644,N_15695);
or U16127 (N_16127,N_15713,N_15549);
nand U16128 (N_16128,N_15775,N_15565);
nor U16129 (N_16129,N_15876,N_15987);
nand U16130 (N_16130,N_15878,N_15635);
nand U16131 (N_16131,N_15574,N_15680);
nor U16132 (N_16132,N_15750,N_15879);
and U16133 (N_16133,N_15758,N_15528);
xor U16134 (N_16134,N_15728,N_15850);
and U16135 (N_16135,N_15838,N_15675);
nand U16136 (N_16136,N_15814,N_15966);
and U16137 (N_16137,N_15917,N_15805);
and U16138 (N_16138,N_15828,N_15807);
nor U16139 (N_16139,N_15591,N_15592);
or U16140 (N_16140,N_15867,N_15951);
and U16141 (N_16141,N_15715,N_15931);
nand U16142 (N_16142,N_15797,N_15899);
nor U16143 (N_16143,N_15769,N_15851);
nor U16144 (N_16144,N_15974,N_15658);
or U16145 (N_16145,N_15989,N_15889);
or U16146 (N_16146,N_15569,N_15833);
and U16147 (N_16147,N_15817,N_15911);
nand U16148 (N_16148,N_15840,N_15977);
nor U16149 (N_16149,N_15958,N_15717);
nand U16150 (N_16150,N_15942,N_15640);
or U16151 (N_16151,N_15891,N_15886);
nand U16152 (N_16152,N_15542,N_15663);
nand U16153 (N_16153,N_15694,N_15541);
and U16154 (N_16154,N_15827,N_15685);
xor U16155 (N_16155,N_15682,N_15524);
or U16156 (N_16156,N_15530,N_15681);
nand U16157 (N_16157,N_15984,N_15735);
and U16158 (N_16158,N_15970,N_15870);
xor U16159 (N_16159,N_15502,N_15748);
or U16160 (N_16160,N_15786,N_15526);
xnor U16161 (N_16161,N_15601,N_15504);
and U16162 (N_16162,N_15766,N_15980);
nor U16163 (N_16163,N_15745,N_15762);
xor U16164 (N_16164,N_15634,N_15600);
nor U16165 (N_16165,N_15696,N_15988);
and U16166 (N_16166,N_15932,N_15998);
xor U16167 (N_16167,N_15619,N_15606);
nand U16168 (N_16168,N_15550,N_15916);
and U16169 (N_16169,N_15510,N_15527);
nand U16170 (N_16170,N_15562,N_15883);
nor U16171 (N_16171,N_15904,N_15599);
and U16172 (N_16172,N_15501,N_15624);
or U16173 (N_16173,N_15736,N_15653);
xor U16174 (N_16174,N_15626,N_15920);
xnor U16175 (N_16175,N_15871,N_15925);
nand U16176 (N_16176,N_15615,N_15845);
nand U16177 (N_16177,N_15949,N_15954);
nor U16178 (N_16178,N_15944,N_15854);
or U16179 (N_16179,N_15799,N_15798);
or U16180 (N_16180,N_15590,N_15674);
and U16181 (N_16181,N_15947,N_15979);
nor U16182 (N_16182,N_15679,N_15730);
xnor U16183 (N_16183,N_15641,N_15796);
nand U16184 (N_16184,N_15742,N_15950);
nand U16185 (N_16185,N_15547,N_15594);
xor U16186 (N_16186,N_15523,N_15513);
or U16187 (N_16187,N_15537,N_15806);
and U16188 (N_16188,N_15887,N_15570);
xor U16189 (N_16189,N_15862,N_15941);
nand U16190 (N_16190,N_15910,N_15824);
nand U16191 (N_16191,N_15890,N_15512);
or U16192 (N_16192,N_15652,N_15801);
or U16193 (N_16193,N_15830,N_15834);
and U16194 (N_16194,N_15691,N_15884);
or U16195 (N_16195,N_15539,N_15546);
nand U16196 (N_16196,N_15540,N_15945);
nor U16197 (N_16197,N_15578,N_15756);
and U16198 (N_16198,N_15620,N_15573);
and U16199 (N_16199,N_15509,N_15724);
nor U16200 (N_16200,N_15521,N_15737);
xor U16201 (N_16201,N_15671,N_15953);
and U16202 (N_16202,N_15670,N_15698);
xnor U16203 (N_16203,N_15855,N_15686);
or U16204 (N_16204,N_15752,N_15844);
nand U16205 (N_16205,N_15722,N_15684);
or U16206 (N_16206,N_15580,N_15690);
or U16207 (N_16207,N_15627,N_15746);
nand U16208 (N_16208,N_15971,N_15577);
or U16209 (N_16209,N_15662,N_15963);
or U16210 (N_16210,N_15738,N_15881);
xor U16211 (N_16211,N_15936,N_15829);
nand U16212 (N_16212,N_15880,N_15791);
or U16213 (N_16213,N_15672,N_15516);
nand U16214 (N_16214,N_15529,N_15803);
nor U16215 (N_16215,N_15543,N_15822);
or U16216 (N_16216,N_15677,N_15648);
nor U16217 (N_16217,N_15933,N_15555);
nor U16218 (N_16218,N_15747,N_15607);
and U16219 (N_16219,N_15602,N_15863);
nand U16220 (N_16220,N_15508,N_15639);
nand U16221 (N_16221,N_15571,N_15628);
or U16222 (N_16222,N_15760,N_15808);
xor U16223 (N_16223,N_15579,N_15517);
and U16224 (N_16224,N_15633,N_15582);
nor U16225 (N_16225,N_15985,N_15688);
and U16226 (N_16226,N_15937,N_15972);
or U16227 (N_16227,N_15701,N_15554);
xnor U16228 (N_16228,N_15832,N_15930);
nor U16229 (N_16229,N_15632,N_15764);
or U16230 (N_16230,N_15907,N_15770);
nand U16231 (N_16231,N_15978,N_15623);
and U16232 (N_16232,N_15866,N_15650);
and U16233 (N_16233,N_15636,N_15558);
nand U16234 (N_16234,N_15703,N_15927);
nand U16235 (N_16235,N_15964,N_15774);
nand U16236 (N_16236,N_15784,N_15783);
nor U16237 (N_16237,N_15614,N_15697);
nor U16238 (N_16238,N_15665,N_15706);
nand U16239 (N_16239,N_15885,N_15859);
nor U16240 (N_16240,N_15908,N_15922);
nand U16241 (N_16241,N_15853,N_15588);
or U16242 (N_16242,N_15755,N_15765);
or U16243 (N_16243,N_15792,N_15823);
xor U16244 (N_16244,N_15821,N_15741);
nor U16245 (N_16245,N_15763,N_15734);
xor U16246 (N_16246,N_15923,N_15727);
and U16247 (N_16247,N_15566,N_15780);
or U16248 (N_16248,N_15782,N_15968);
xnor U16249 (N_16249,N_15721,N_15503);
and U16250 (N_16250,N_15872,N_15726);
nand U16251 (N_16251,N_15546,N_15516);
and U16252 (N_16252,N_15912,N_15991);
or U16253 (N_16253,N_15701,N_15857);
nor U16254 (N_16254,N_15867,N_15738);
xor U16255 (N_16255,N_15667,N_15952);
nor U16256 (N_16256,N_15919,N_15936);
nand U16257 (N_16257,N_15950,N_15506);
nor U16258 (N_16258,N_15607,N_15778);
xor U16259 (N_16259,N_15697,N_15772);
and U16260 (N_16260,N_15876,N_15804);
xnor U16261 (N_16261,N_15924,N_15858);
or U16262 (N_16262,N_15917,N_15539);
and U16263 (N_16263,N_15598,N_15765);
and U16264 (N_16264,N_15967,N_15628);
or U16265 (N_16265,N_15835,N_15736);
nor U16266 (N_16266,N_15786,N_15714);
or U16267 (N_16267,N_15546,N_15558);
and U16268 (N_16268,N_15668,N_15969);
xnor U16269 (N_16269,N_15935,N_15690);
xnor U16270 (N_16270,N_15859,N_15972);
and U16271 (N_16271,N_15677,N_15894);
or U16272 (N_16272,N_15926,N_15806);
nand U16273 (N_16273,N_15629,N_15712);
or U16274 (N_16274,N_15868,N_15849);
nand U16275 (N_16275,N_15903,N_15809);
or U16276 (N_16276,N_15858,N_15543);
nor U16277 (N_16277,N_15633,N_15878);
and U16278 (N_16278,N_15936,N_15818);
xnor U16279 (N_16279,N_15801,N_15924);
and U16280 (N_16280,N_15636,N_15732);
xnor U16281 (N_16281,N_15676,N_15746);
nor U16282 (N_16282,N_15865,N_15724);
nor U16283 (N_16283,N_15854,N_15644);
nand U16284 (N_16284,N_15967,N_15851);
nor U16285 (N_16285,N_15696,N_15730);
nand U16286 (N_16286,N_15878,N_15801);
and U16287 (N_16287,N_15811,N_15691);
or U16288 (N_16288,N_15824,N_15631);
or U16289 (N_16289,N_15799,N_15891);
nor U16290 (N_16290,N_15988,N_15876);
nand U16291 (N_16291,N_15796,N_15880);
nand U16292 (N_16292,N_15954,N_15874);
nand U16293 (N_16293,N_15805,N_15716);
or U16294 (N_16294,N_15992,N_15790);
xnor U16295 (N_16295,N_15935,N_15972);
xnor U16296 (N_16296,N_15919,N_15712);
nor U16297 (N_16297,N_15897,N_15509);
or U16298 (N_16298,N_15773,N_15512);
and U16299 (N_16299,N_15737,N_15507);
xor U16300 (N_16300,N_15544,N_15642);
nand U16301 (N_16301,N_15953,N_15574);
and U16302 (N_16302,N_15563,N_15887);
or U16303 (N_16303,N_15860,N_15503);
and U16304 (N_16304,N_15712,N_15770);
xor U16305 (N_16305,N_15690,N_15913);
nand U16306 (N_16306,N_15937,N_15753);
nand U16307 (N_16307,N_15750,N_15818);
nor U16308 (N_16308,N_15541,N_15799);
and U16309 (N_16309,N_15566,N_15749);
and U16310 (N_16310,N_15990,N_15615);
and U16311 (N_16311,N_15863,N_15519);
nor U16312 (N_16312,N_15553,N_15737);
and U16313 (N_16313,N_15875,N_15697);
nand U16314 (N_16314,N_15838,N_15680);
nor U16315 (N_16315,N_15520,N_15503);
xnor U16316 (N_16316,N_15553,N_15826);
and U16317 (N_16317,N_15609,N_15873);
and U16318 (N_16318,N_15949,N_15970);
or U16319 (N_16319,N_15527,N_15730);
or U16320 (N_16320,N_15541,N_15884);
or U16321 (N_16321,N_15573,N_15786);
and U16322 (N_16322,N_15838,N_15866);
and U16323 (N_16323,N_15840,N_15857);
and U16324 (N_16324,N_15621,N_15682);
nand U16325 (N_16325,N_15964,N_15952);
or U16326 (N_16326,N_15716,N_15963);
and U16327 (N_16327,N_15577,N_15582);
and U16328 (N_16328,N_15769,N_15579);
and U16329 (N_16329,N_15669,N_15659);
or U16330 (N_16330,N_15540,N_15542);
nand U16331 (N_16331,N_15650,N_15781);
and U16332 (N_16332,N_15962,N_15979);
or U16333 (N_16333,N_15651,N_15731);
nand U16334 (N_16334,N_15875,N_15746);
and U16335 (N_16335,N_15912,N_15609);
nor U16336 (N_16336,N_15832,N_15874);
and U16337 (N_16337,N_15835,N_15613);
and U16338 (N_16338,N_15596,N_15721);
and U16339 (N_16339,N_15762,N_15885);
nand U16340 (N_16340,N_15617,N_15967);
nor U16341 (N_16341,N_15971,N_15767);
and U16342 (N_16342,N_15823,N_15577);
or U16343 (N_16343,N_15959,N_15518);
and U16344 (N_16344,N_15737,N_15527);
and U16345 (N_16345,N_15548,N_15850);
xor U16346 (N_16346,N_15773,N_15532);
or U16347 (N_16347,N_15838,N_15676);
nand U16348 (N_16348,N_15864,N_15685);
nor U16349 (N_16349,N_15530,N_15512);
nor U16350 (N_16350,N_15814,N_15871);
nor U16351 (N_16351,N_15917,N_15987);
xor U16352 (N_16352,N_15942,N_15784);
nor U16353 (N_16353,N_15993,N_15584);
xor U16354 (N_16354,N_15597,N_15753);
and U16355 (N_16355,N_15647,N_15987);
or U16356 (N_16356,N_15954,N_15985);
nor U16357 (N_16357,N_15763,N_15652);
xnor U16358 (N_16358,N_15833,N_15876);
and U16359 (N_16359,N_15824,N_15604);
nand U16360 (N_16360,N_15732,N_15737);
and U16361 (N_16361,N_15893,N_15659);
nor U16362 (N_16362,N_15997,N_15884);
and U16363 (N_16363,N_15935,N_15713);
nand U16364 (N_16364,N_15849,N_15507);
and U16365 (N_16365,N_15516,N_15507);
nor U16366 (N_16366,N_15684,N_15948);
nand U16367 (N_16367,N_15591,N_15856);
nand U16368 (N_16368,N_15619,N_15640);
xnor U16369 (N_16369,N_15646,N_15562);
xnor U16370 (N_16370,N_15771,N_15840);
nand U16371 (N_16371,N_15913,N_15673);
nor U16372 (N_16372,N_15852,N_15665);
or U16373 (N_16373,N_15685,N_15627);
or U16374 (N_16374,N_15639,N_15804);
or U16375 (N_16375,N_15818,N_15920);
and U16376 (N_16376,N_15522,N_15684);
nor U16377 (N_16377,N_15746,N_15712);
xnor U16378 (N_16378,N_15789,N_15718);
or U16379 (N_16379,N_15675,N_15857);
nand U16380 (N_16380,N_15748,N_15968);
nand U16381 (N_16381,N_15950,N_15517);
xnor U16382 (N_16382,N_15788,N_15809);
nand U16383 (N_16383,N_15504,N_15833);
and U16384 (N_16384,N_15849,N_15805);
or U16385 (N_16385,N_15766,N_15837);
nand U16386 (N_16386,N_15535,N_15787);
or U16387 (N_16387,N_15528,N_15965);
xor U16388 (N_16388,N_15593,N_15758);
nor U16389 (N_16389,N_15647,N_15658);
xnor U16390 (N_16390,N_15854,N_15578);
xor U16391 (N_16391,N_15847,N_15996);
xnor U16392 (N_16392,N_15560,N_15762);
nor U16393 (N_16393,N_15913,N_15541);
nor U16394 (N_16394,N_15821,N_15600);
nand U16395 (N_16395,N_15894,N_15671);
or U16396 (N_16396,N_15998,N_15721);
or U16397 (N_16397,N_15988,N_15920);
nor U16398 (N_16398,N_15636,N_15610);
xor U16399 (N_16399,N_15803,N_15858);
or U16400 (N_16400,N_15948,N_15549);
and U16401 (N_16401,N_15900,N_15572);
xor U16402 (N_16402,N_15583,N_15781);
nand U16403 (N_16403,N_15972,N_15842);
and U16404 (N_16404,N_15839,N_15975);
xnor U16405 (N_16405,N_15534,N_15700);
and U16406 (N_16406,N_15948,N_15997);
xnor U16407 (N_16407,N_15649,N_15559);
and U16408 (N_16408,N_15781,N_15895);
nor U16409 (N_16409,N_15518,N_15918);
xnor U16410 (N_16410,N_15901,N_15972);
and U16411 (N_16411,N_15655,N_15605);
xor U16412 (N_16412,N_15603,N_15791);
xor U16413 (N_16413,N_15639,N_15553);
nor U16414 (N_16414,N_15591,N_15643);
and U16415 (N_16415,N_15706,N_15523);
and U16416 (N_16416,N_15991,N_15901);
nand U16417 (N_16417,N_15772,N_15960);
or U16418 (N_16418,N_15624,N_15891);
nand U16419 (N_16419,N_15645,N_15994);
xor U16420 (N_16420,N_15517,N_15643);
nand U16421 (N_16421,N_15587,N_15646);
nand U16422 (N_16422,N_15603,N_15615);
nor U16423 (N_16423,N_15977,N_15926);
and U16424 (N_16424,N_15637,N_15561);
xor U16425 (N_16425,N_15697,N_15564);
and U16426 (N_16426,N_15793,N_15929);
or U16427 (N_16427,N_15971,N_15927);
nand U16428 (N_16428,N_15694,N_15979);
nand U16429 (N_16429,N_15896,N_15582);
or U16430 (N_16430,N_15979,N_15607);
nor U16431 (N_16431,N_15690,N_15624);
or U16432 (N_16432,N_15831,N_15577);
nor U16433 (N_16433,N_15801,N_15612);
nor U16434 (N_16434,N_15664,N_15716);
nand U16435 (N_16435,N_15788,N_15627);
nor U16436 (N_16436,N_15962,N_15504);
nand U16437 (N_16437,N_15709,N_15578);
or U16438 (N_16438,N_15714,N_15602);
nand U16439 (N_16439,N_15966,N_15673);
and U16440 (N_16440,N_15981,N_15576);
xor U16441 (N_16441,N_15892,N_15686);
or U16442 (N_16442,N_15707,N_15994);
or U16443 (N_16443,N_15639,N_15841);
and U16444 (N_16444,N_15879,N_15518);
or U16445 (N_16445,N_15846,N_15551);
xor U16446 (N_16446,N_15721,N_15587);
or U16447 (N_16447,N_15851,N_15709);
or U16448 (N_16448,N_15758,N_15527);
and U16449 (N_16449,N_15737,N_15599);
and U16450 (N_16450,N_15567,N_15796);
nor U16451 (N_16451,N_15864,N_15531);
xnor U16452 (N_16452,N_15750,N_15949);
xor U16453 (N_16453,N_15582,N_15730);
or U16454 (N_16454,N_15515,N_15551);
nor U16455 (N_16455,N_15646,N_15644);
and U16456 (N_16456,N_15794,N_15619);
or U16457 (N_16457,N_15645,N_15591);
xor U16458 (N_16458,N_15569,N_15608);
or U16459 (N_16459,N_15965,N_15707);
nor U16460 (N_16460,N_15620,N_15994);
and U16461 (N_16461,N_15705,N_15812);
xnor U16462 (N_16462,N_15546,N_15590);
and U16463 (N_16463,N_15787,N_15900);
xor U16464 (N_16464,N_15519,N_15571);
nand U16465 (N_16465,N_15975,N_15621);
nand U16466 (N_16466,N_15983,N_15592);
and U16467 (N_16467,N_15907,N_15626);
xor U16468 (N_16468,N_15561,N_15628);
nand U16469 (N_16469,N_15786,N_15673);
or U16470 (N_16470,N_15590,N_15673);
and U16471 (N_16471,N_15702,N_15562);
nand U16472 (N_16472,N_15660,N_15777);
nor U16473 (N_16473,N_15595,N_15926);
nand U16474 (N_16474,N_15627,N_15941);
and U16475 (N_16475,N_15770,N_15797);
and U16476 (N_16476,N_15697,N_15856);
xnor U16477 (N_16477,N_15893,N_15684);
and U16478 (N_16478,N_15873,N_15972);
or U16479 (N_16479,N_15574,N_15562);
xor U16480 (N_16480,N_15955,N_15666);
nand U16481 (N_16481,N_15525,N_15922);
or U16482 (N_16482,N_15706,N_15820);
xnor U16483 (N_16483,N_15794,N_15930);
nand U16484 (N_16484,N_15661,N_15778);
or U16485 (N_16485,N_15577,N_15837);
nor U16486 (N_16486,N_15560,N_15852);
and U16487 (N_16487,N_15751,N_15577);
nor U16488 (N_16488,N_15778,N_15846);
or U16489 (N_16489,N_15819,N_15510);
nor U16490 (N_16490,N_15723,N_15936);
nor U16491 (N_16491,N_15747,N_15504);
xnor U16492 (N_16492,N_15870,N_15750);
nor U16493 (N_16493,N_15594,N_15509);
or U16494 (N_16494,N_15715,N_15849);
and U16495 (N_16495,N_15792,N_15973);
and U16496 (N_16496,N_15568,N_15597);
nand U16497 (N_16497,N_15558,N_15563);
and U16498 (N_16498,N_15833,N_15965);
xnor U16499 (N_16499,N_15730,N_15605);
and U16500 (N_16500,N_16261,N_16438);
or U16501 (N_16501,N_16467,N_16455);
nor U16502 (N_16502,N_16496,N_16354);
or U16503 (N_16503,N_16017,N_16378);
xor U16504 (N_16504,N_16210,N_16126);
nand U16505 (N_16505,N_16301,N_16183);
and U16506 (N_16506,N_16451,N_16476);
nand U16507 (N_16507,N_16380,N_16386);
and U16508 (N_16508,N_16297,N_16216);
or U16509 (N_16509,N_16286,N_16437);
xnor U16510 (N_16510,N_16322,N_16489);
nor U16511 (N_16511,N_16275,N_16133);
xnor U16512 (N_16512,N_16213,N_16135);
or U16513 (N_16513,N_16440,N_16247);
and U16514 (N_16514,N_16391,N_16242);
or U16515 (N_16515,N_16482,N_16282);
or U16516 (N_16516,N_16016,N_16499);
xnor U16517 (N_16517,N_16112,N_16163);
or U16518 (N_16518,N_16290,N_16232);
or U16519 (N_16519,N_16098,N_16356);
and U16520 (N_16520,N_16346,N_16295);
and U16521 (N_16521,N_16487,N_16044);
and U16522 (N_16522,N_16457,N_16330);
and U16523 (N_16523,N_16161,N_16448);
nor U16524 (N_16524,N_16478,N_16184);
or U16525 (N_16525,N_16074,N_16197);
or U16526 (N_16526,N_16260,N_16004);
xor U16527 (N_16527,N_16283,N_16488);
and U16528 (N_16528,N_16234,N_16195);
and U16529 (N_16529,N_16361,N_16119);
xor U16530 (N_16530,N_16257,N_16079);
nor U16531 (N_16531,N_16370,N_16419);
and U16532 (N_16532,N_16353,N_16060);
nor U16533 (N_16533,N_16095,N_16472);
nand U16534 (N_16534,N_16229,N_16070);
or U16535 (N_16535,N_16086,N_16148);
nor U16536 (N_16536,N_16304,N_16019);
nor U16537 (N_16537,N_16055,N_16340);
nand U16538 (N_16538,N_16453,N_16206);
nor U16539 (N_16539,N_16037,N_16491);
or U16540 (N_16540,N_16108,N_16402);
and U16541 (N_16541,N_16377,N_16165);
nor U16542 (N_16542,N_16403,N_16139);
nor U16543 (N_16543,N_16116,N_16101);
and U16544 (N_16544,N_16387,N_16006);
nand U16545 (N_16545,N_16299,N_16039);
and U16546 (N_16546,N_16199,N_16043);
nor U16547 (N_16547,N_16179,N_16315);
xnor U16548 (N_16548,N_16407,N_16097);
xor U16549 (N_16549,N_16110,N_16463);
nor U16550 (N_16550,N_16347,N_16471);
or U16551 (N_16551,N_16452,N_16464);
nand U16552 (N_16552,N_16316,N_16099);
nor U16553 (N_16553,N_16351,N_16169);
nor U16554 (N_16554,N_16211,N_16233);
or U16555 (N_16555,N_16185,N_16313);
nor U16556 (N_16556,N_16320,N_16011);
and U16557 (N_16557,N_16454,N_16157);
xnor U16558 (N_16558,N_16150,N_16344);
nand U16559 (N_16559,N_16287,N_16468);
xnor U16560 (N_16560,N_16067,N_16032);
nand U16561 (N_16561,N_16420,N_16042);
nand U16562 (N_16562,N_16334,N_16433);
xor U16563 (N_16563,N_16336,N_16240);
nand U16564 (N_16564,N_16125,N_16100);
xnor U16565 (N_16565,N_16397,N_16461);
xnor U16566 (N_16566,N_16432,N_16382);
or U16567 (N_16567,N_16312,N_16328);
xnor U16568 (N_16568,N_16159,N_16020);
nor U16569 (N_16569,N_16372,N_16187);
and U16570 (N_16570,N_16041,N_16052);
nor U16571 (N_16571,N_16379,N_16327);
nand U16572 (N_16572,N_16325,N_16215);
and U16573 (N_16573,N_16141,N_16289);
nand U16574 (N_16574,N_16196,N_16331);
and U16575 (N_16575,N_16271,N_16355);
nor U16576 (N_16576,N_16409,N_16064);
xnor U16577 (N_16577,N_16326,N_16430);
or U16578 (N_16578,N_16046,N_16236);
and U16579 (N_16579,N_16250,N_16214);
and U16580 (N_16580,N_16173,N_16235);
nor U16581 (N_16581,N_16104,N_16404);
nand U16582 (N_16582,N_16113,N_16341);
or U16583 (N_16583,N_16167,N_16300);
xnor U16584 (N_16584,N_16094,N_16492);
or U16585 (N_16585,N_16219,N_16337);
nand U16586 (N_16586,N_16057,N_16027);
nor U16587 (N_16587,N_16127,N_16137);
nor U16588 (N_16588,N_16237,N_16117);
or U16589 (N_16589,N_16134,N_16308);
and U16590 (N_16590,N_16026,N_16462);
xnor U16591 (N_16591,N_16458,N_16049);
or U16592 (N_16592,N_16158,N_16224);
and U16593 (N_16593,N_16256,N_16217);
or U16594 (N_16594,N_16259,N_16352);
nand U16595 (N_16595,N_16193,N_16152);
or U16596 (N_16596,N_16151,N_16318);
and U16597 (N_16597,N_16477,N_16093);
or U16598 (N_16598,N_16246,N_16059);
and U16599 (N_16599,N_16305,N_16441);
nand U16600 (N_16600,N_16121,N_16203);
xor U16601 (N_16601,N_16460,N_16083);
nand U16602 (N_16602,N_16238,N_16385);
nor U16603 (N_16603,N_16040,N_16288);
nand U16604 (N_16604,N_16479,N_16263);
and U16605 (N_16605,N_16075,N_16009);
nand U16606 (N_16606,N_16400,N_16048);
or U16607 (N_16607,N_16221,N_16178);
or U16608 (N_16608,N_16031,N_16084);
and U16609 (N_16609,N_16231,N_16294);
nor U16610 (N_16610,N_16002,N_16091);
nor U16611 (N_16611,N_16138,N_16474);
and U16612 (N_16612,N_16000,N_16191);
or U16613 (N_16613,N_16324,N_16005);
nor U16614 (N_16614,N_16359,N_16124);
and U16615 (N_16615,N_16106,N_16089);
or U16616 (N_16616,N_16025,N_16285);
and U16617 (N_16617,N_16072,N_16003);
nand U16618 (N_16618,N_16146,N_16349);
xor U16619 (N_16619,N_16014,N_16303);
nand U16620 (N_16620,N_16245,N_16473);
or U16621 (N_16621,N_16367,N_16088);
nor U16622 (N_16622,N_16228,N_16045);
nor U16623 (N_16623,N_16068,N_16241);
and U16624 (N_16624,N_16076,N_16033);
or U16625 (N_16625,N_16053,N_16298);
and U16626 (N_16626,N_16481,N_16333);
and U16627 (N_16627,N_16147,N_16227);
nand U16628 (N_16628,N_16415,N_16202);
or U16629 (N_16629,N_16155,N_16388);
xnor U16630 (N_16630,N_16248,N_16309);
nor U16631 (N_16631,N_16480,N_16495);
xnor U16632 (N_16632,N_16425,N_16439);
nor U16633 (N_16633,N_16485,N_16080);
nor U16634 (N_16634,N_16434,N_16443);
xor U16635 (N_16635,N_16058,N_16396);
nand U16636 (N_16636,N_16281,N_16024);
nor U16637 (N_16637,N_16450,N_16066);
nand U16638 (N_16638,N_16456,N_16272);
and U16639 (N_16639,N_16278,N_16369);
and U16640 (N_16640,N_16291,N_16062);
nor U16641 (N_16641,N_16343,N_16149);
or U16642 (N_16642,N_16436,N_16047);
nor U16643 (N_16643,N_16253,N_16426);
or U16644 (N_16644,N_16270,N_16408);
xnor U16645 (N_16645,N_16130,N_16244);
or U16646 (N_16646,N_16174,N_16390);
nand U16647 (N_16647,N_16366,N_16389);
or U16648 (N_16648,N_16252,N_16265);
and U16649 (N_16649,N_16394,N_16310);
or U16650 (N_16650,N_16345,N_16063);
or U16651 (N_16651,N_16118,N_16411);
or U16652 (N_16652,N_16249,N_16077);
nor U16653 (N_16653,N_16268,N_16189);
nand U16654 (N_16654,N_16225,N_16494);
or U16655 (N_16655,N_16383,N_16144);
or U16656 (N_16656,N_16132,N_16267);
or U16657 (N_16657,N_16162,N_16358);
and U16658 (N_16658,N_16273,N_16056);
nor U16659 (N_16659,N_16170,N_16103);
or U16660 (N_16660,N_16414,N_16131);
xnor U16661 (N_16661,N_16306,N_16405);
nand U16662 (N_16662,N_16096,N_16470);
or U16663 (N_16663,N_16384,N_16128);
and U16664 (N_16664,N_16164,N_16081);
or U16665 (N_16665,N_16207,N_16090);
and U16666 (N_16666,N_16483,N_16194);
or U16667 (N_16667,N_16412,N_16065);
or U16668 (N_16668,N_16204,N_16406);
and U16669 (N_16669,N_16010,N_16007);
nor U16670 (N_16670,N_16442,N_16449);
xor U16671 (N_16671,N_16251,N_16444);
nand U16672 (N_16672,N_16092,N_16078);
nand U16673 (N_16673,N_16348,N_16319);
nand U16674 (N_16674,N_16218,N_16277);
nand U16675 (N_16675,N_16381,N_16314);
xor U16676 (N_16676,N_16395,N_16051);
nor U16677 (N_16677,N_16226,N_16317);
xor U16678 (N_16678,N_16362,N_16279);
nand U16679 (N_16679,N_16114,N_16435);
xnor U16680 (N_16680,N_16373,N_16469);
xor U16681 (N_16681,N_16422,N_16190);
nor U16682 (N_16682,N_16365,N_16012);
nor U16683 (N_16683,N_16208,N_16028);
xor U16684 (N_16684,N_16311,N_16035);
xnor U16685 (N_16685,N_16357,N_16200);
and U16686 (N_16686,N_16156,N_16030);
and U16687 (N_16687,N_16486,N_16085);
xnor U16688 (N_16688,N_16364,N_16160);
or U16689 (N_16689,N_16129,N_16182);
nand U16690 (N_16690,N_16175,N_16363);
and U16691 (N_16691,N_16050,N_16177);
xnor U16692 (N_16692,N_16493,N_16446);
or U16693 (N_16693,N_16198,N_16323);
or U16694 (N_16694,N_16071,N_16153);
xnor U16695 (N_16695,N_16416,N_16418);
xnor U16696 (N_16696,N_16209,N_16262);
and U16697 (N_16697,N_16168,N_16201);
or U16698 (N_16698,N_16484,N_16109);
nand U16699 (N_16699,N_16181,N_16143);
nand U16700 (N_16700,N_16284,N_16061);
and U16701 (N_16701,N_16447,N_16023);
nand U16702 (N_16702,N_16398,N_16421);
nor U16703 (N_16703,N_16102,N_16293);
xnor U16704 (N_16704,N_16166,N_16417);
nand U16705 (N_16705,N_16008,N_16498);
nor U16706 (N_16706,N_16401,N_16222);
and U16707 (N_16707,N_16223,N_16329);
and U16708 (N_16708,N_16029,N_16038);
or U16709 (N_16709,N_16392,N_16212);
xnor U16710 (N_16710,N_16332,N_16136);
nor U16711 (N_16711,N_16339,N_16368);
or U16712 (N_16712,N_16034,N_16497);
nand U16713 (N_16713,N_16021,N_16274);
or U16714 (N_16714,N_16423,N_16192);
xor U16715 (N_16715,N_16475,N_16082);
and U16716 (N_16716,N_16054,N_16360);
and U16717 (N_16717,N_16427,N_16073);
nor U16718 (N_16718,N_16255,N_16429);
xnor U16719 (N_16719,N_16376,N_16410);
nor U16720 (N_16720,N_16445,N_16269);
or U16721 (N_16721,N_16266,N_16375);
or U16722 (N_16722,N_16015,N_16230);
and U16723 (N_16723,N_16171,N_16205);
or U16724 (N_16724,N_16254,N_16280);
xnor U16725 (N_16725,N_16466,N_16431);
and U16726 (N_16726,N_16239,N_16107);
xor U16727 (N_16727,N_16154,N_16018);
xor U16728 (N_16728,N_16307,N_16292);
xnor U16729 (N_16729,N_16145,N_16276);
xnor U16730 (N_16730,N_16123,N_16176);
nor U16731 (N_16731,N_16321,N_16399);
or U16732 (N_16732,N_16264,N_16374);
xnor U16733 (N_16733,N_16188,N_16022);
nor U16734 (N_16734,N_16180,N_16001);
xnor U16735 (N_16735,N_16490,N_16122);
or U16736 (N_16736,N_16465,N_16342);
xnor U16737 (N_16737,N_16302,N_16413);
nor U16738 (N_16738,N_16105,N_16350);
nand U16739 (N_16739,N_16140,N_16296);
nand U16740 (N_16740,N_16036,N_16186);
nor U16741 (N_16741,N_16115,N_16335);
nor U16742 (N_16742,N_16111,N_16371);
nand U16743 (N_16743,N_16258,N_16172);
and U16744 (N_16744,N_16459,N_16243);
xor U16745 (N_16745,N_16013,N_16393);
or U16746 (N_16746,N_16087,N_16338);
nor U16747 (N_16747,N_16069,N_16142);
nand U16748 (N_16748,N_16120,N_16428);
or U16749 (N_16749,N_16424,N_16220);
and U16750 (N_16750,N_16200,N_16280);
nor U16751 (N_16751,N_16175,N_16484);
nand U16752 (N_16752,N_16033,N_16304);
nand U16753 (N_16753,N_16274,N_16105);
xor U16754 (N_16754,N_16004,N_16377);
nor U16755 (N_16755,N_16203,N_16070);
and U16756 (N_16756,N_16373,N_16097);
nand U16757 (N_16757,N_16378,N_16355);
and U16758 (N_16758,N_16061,N_16161);
xnor U16759 (N_16759,N_16202,N_16493);
xor U16760 (N_16760,N_16072,N_16183);
nor U16761 (N_16761,N_16113,N_16099);
nor U16762 (N_16762,N_16414,N_16028);
or U16763 (N_16763,N_16116,N_16243);
and U16764 (N_16764,N_16018,N_16193);
nand U16765 (N_16765,N_16284,N_16275);
nand U16766 (N_16766,N_16022,N_16355);
xor U16767 (N_16767,N_16211,N_16493);
or U16768 (N_16768,N_16328,N_16462);
or U16769 (N_16769,N_16304,N_16083);
nor U16770 (N_16770,N_16289,N_16273);
nor U16771 (N_16771,N_16155,N_16406);
or U16772 (N_16772,N_16314,N_16462);
xor U16773 (N_16773,N_16311,N_16141);
nor U16774 (N_16774,N_16265,N_16384);
or U16775 (N_16775,N_16197,N_16214);
or U16776 (N_16776,N_16343,N_16456);
and U16777 (N_16777,N_16307,N_16140);
and U16778 (N_16778,N_16483,N_16222);
and U16779 (N_16779,N_16046,N_16080);
or U16780 (N_16780,N_16339,N_16329);
xnor U16781 (N_16781,N_16053,N_16224);
xnor U16782 (N_16782,N_16028,N_16009);
and U16783 (N_16783,N_16197,N_16268);
and U16784 (N_16784,N_16328,N_16425);
and U16785 (N_16785,N_16450,N_16388);
and U16786 (N_16786,N_16088,N_16398);
and U16787 (N_16787,N_16172,N_16155);
nand U16788 (N_16788,N_16305,N_16169);
xnor U16789 (N_16789,N_16300,N_16018);
nor U16790 (N_16790,N_16001,N_16286);
or U16791 (N_16791,N_16162,N_16135);
xnor U16792 (N_16792,N_16262,N_16004);
nand U16793 (N_16793,N_16040,N_16074);
nor U16794 (N_16794,N_16158,N_16094);
nor U16795 (N_16795,N_16393,N_16031);
or U16796 (N_16796,N_16459,N_16269);
and U16797 (N_16797,N_16439,N_16113);
and U16798 (N_16798,N_16125,N_16090);
xnor U16799 (N_16799,N_16344,N_16278);
xor U16800 (N_16800,N_16371,N_16076);
nand U16801 (N_16801,N_16203,N_16449);
or U16802 (N_16802,N_16269,N_16277);
xnor U16803 (N_16803,N_16330,N_16270);
nand U16804 (N_16804,N_16069,N_16054);
or U16805 (N_16805,N_16029,N_16362);
nand U16806 (N_16806,N_16359,N_16206);
nand U16807 (N_16807,N_16381,N_16446);
and U16808 (N_16808,N_16048,N_16356);
nor U16809 (N_16809,N_16000,N_16474);
or U16810 (N_16810,N_16095,N_16458);
nand U16811 (N_16811,N_16431,N_16090);
xnor U16812 (N_16812,N_16300,N_16064);
nand U16813 (N_16813,N_16285,N_16492);
xnor U16814 (N_16814,N_16106,N_16484);
nor U16815 (N_16815,N_16497,N_16127);
nor U16816 (N_16816,N_16232,N_16075);
xor U16817 (N_16817,N_16321,N_16380);
nand U16818 (N_16818,N_16494,N_16274);
xnor U16819 (N_16819,N_16447,N_16202);
xnor U16820 (N_16820,N_16056,N_16383);
or U16821 (N_16821,N_16019,N_16102);
nand U16822 (N_16822,N_16199,N_16225);
or U16823 (N_16823,N_16481,N_16076);
xnor U16824 (N_16824,N_16058,N_16341);
nor U16825 (N_16825,N_16171,N_16103);
nand U16826 (N_16826,N_16435,N_16098);
or U16827 (N_16827,N_16354,N_16158);
nor U16828 (N_16828,N_16273,N_16378);
xnor U16829 (N_16829,N_16186,N_16173);
and U16830 (N_16830,N_16411,N_16450);
nor U16831 (N_16831,N_16085,N_16480);
or U16832 (N_16832,N_16481,N_16235);
or U16833 (N_16833,N_16250,N_16206);
and U16834 (N_16834,N_16394,N_16266);
and U16835 (N_16835,N_16341,N_16338);
nor U16836 (N_16836,N_16416,N_16076);
xor U16837 (N_16837,N_16438,N_16491);
xor U16838 (N_16838,N_16258,N_16495);
nand U16839 (N_16839,N_16482,N_16409);
nor U16840 (N_16840,N_16157,N_16288);
xnor U16841 (N_16841,N_16092,N_16000);
and U16842 (N_16842,N_16210,N_16166);
nor U16843 (N_16843,N_16198,N_16146);
or U16844 (N_16844,N_16498,N_16201);
and U16845 (N_16845,N_16271,N_16388);
xor U16846 (N_16846,N_16263,N_16273);
and U16847 (N_16847,N_16319,N_16453);
and U16848 (N_16848,N_16401,N_16337);
and U16849 (N_16849,N_16435,N_16056);
nor U16850 (N_16850,N_16034,N_16398);
nand U16851 (N_16851,N_16073,N_16316);
and U16852 (N_16852,N_16173,N_16017);
nand U16853 (N_16853,N_16123,N_16314);
or U16854 (N_16854,N_16338,N_16334);
nand U16855 (N_16855,N_16308,N_16211);
and U16856 (N_16856,N_16037,N_16142);
nand U16857 (N_16857,N_16018,N_16249);
and U16858 (N_16858,N_16137,N_16094);
xor U16859 (N_16859,N_16338,N_16342);
and U16860 (N_16860,N_16187,N_16026);
xor U16861 (N_16861,N_16456,N_16222);
and U16862 (N_16862,N_16228,N_16011);
xor U16863 (N_16863,N_16186,N_16323);
nor U16864 (N_16864,N_16037,N_16072);
xor U16865 (N_16865,N_16196,N_16185);
nor U16866 (N_16866,N_16374,N_16410);
or U16867 (N_16867,N_16185,N_16388);
nor U16868 (N_16868,N_16203,N_16054);
nand U16869 (N_16869,N_16197,N_16048);
or U16870 (N_16870,N_16344,N_16414);
or U16871 (N_16871,N_16182,N_16082);
nand U16872 (N_16872,N_16217,N_16144);
nand U16873 (N_16873,N_16069,N_16491);
nand U16874 (N_16874,N_16484,N_16146);
or U16875 (N_16875,N_16031,N_16095);
or U16876 (N_16876,N_16489,N_16361);
nand U16877 (N_16877,N_16000,N_16324);
nor U16878 (N_16878,N_16487,N_16160);
xor U16879 (N_16879,N_16466,N_16176);
and U16880 (N_16880,N_16156,N_16058);
nand U16881 (N_16881,N_16136,N_16312);
nand U16882 (N_16882,N_16039,N_16450);
xor U16883 (N_16883,N_16314,N_16493);
xor U16884 (N_16884,N_16492,N_16082);
xnor U16885 (N_16885,N_16308,N_16083);
xnor U16886 (N_16886,N_16354,N_16079);
and U16887 (N_16887,N_16145,N_16013);
nor U16888 (N_16888,N_16060,N_16223);
xor U16889 (N_16889,N_16399,N_16140);
or U16890 (N_16890,N_16148,N_16239);
xnor U16891 (N_16891,N_16038,N_16008);
nor U16892 (N_16892,N_16025,N_16417);
nor U16893 (N_16893,N_16447,N_16083);
or U16894 (N_16894,N_16145,N_16333);
nand U16895 (N_16895,N_16000,N_16294);
or U16896 (N_16896,N_16492,N_16231);
and U16897 (N_16897,N_16359,N_16087);
xor U16898 (N_16898,N_16302,N_16369);
nor U16899 (N_16899,N_16369,N_16069);
nand U16900 (N_16900,N_16418,N_16474);
xnor U16901 (N_16901,N_16404,N_16339);
and U16902 (N_16902,N_16178,N_16205);
nand U16903 (N_16903,N_16281,N_16368);
nor U16904 (N_16904,N_16001,N_16093);
nor U16905 (N_16905,N_16396,N_16146);
xnor U16906 (N_16906,N_16167,N_16132);
or U16907 (N_16907,N_16178,N_16249);
nand U16908 (N_16908,N_16450,N_16331);
or U16909 (N_16909,N_16487,N_16332);
nor U16910 (N_16910,N_16297,N_16275);
nor U16911 (N_16911,N_16134,N_16097);
nand U16912 (N_16912,N_16044,N_16135);
and U16913 (N_16913,N_16249,N_16273);
or U16914 (N_16914,N_16465,N_16258);
and U16915 (N_16915,N_16413,N_16273);
nor U16916 (N_16916,N_16045,N_16237);
nor U16917 (N_16917,N_16114,N_16025);
and U16918 (N_16918,N_16445,N_16436);
xor U16919 (N_16919,N_16127,N_16276);
and U16920 (N_16920,N_16164,N_16373);
or U16921 (N_16921,N_16473,N_16356);
nand U16922 (N_16922,N_16109,N_16171);
nor U16923 (N_16923,N_16182,N_16106);
or U16924 (N_16924,N_16134,N_16061);
nand U16925 (N_16925,N_16125,N_16412);
and U16926 (N_16926,N_16315,N_16060);
nand U16927 (N_16927,N_16031,N_16112);
nor U16928 (N_16928,N_16451,N_16465);
nand U16929 (N_16929,N_16091,N_16289);
nand U16930 (N_16930,N_16123,N_16378);
nor U16931 (N_16931,N_16494,N_16219);
nand U16932 (N_16932,N_16053,N_16463);
nor U16933 (N_16933,N_16434,N_16216);
and U16934 (N_16934,N_16258,N_16048);
xor U16935 (N_16935,N_16061,N_16405);
nand U16936 (N_16936,N_16372,N_16159);
nor U16937 (N_16937,N_16464,N_16478);
or U16938 (N_16938,N_16070,N_16176);
and U16939 (N_16939,N_16355,N_16302);
nor U16940 (N_16940,N_16227,N_16102);
xnor U16941 (N_16941,N_16163,N_16381);
xor U16942 (N_16942,N_16477,N_16250);
nand U16943 (N_16943,N_16257,N_16318);
nor U16944 (N_16944,N_16120,N_16047);
or U16945 (N_16945,N_16118,N_16431);
xor U16946 (N_16946,N_16433,N_16366);
nor U16947 (N_16947,N_16177,N_16340);
xnor U16948 (N_16948,N_16459,N_16068);
nand U16949 (N_16949,N_16087,N_16052);
and U16950 (N_16950,N_16043,N_16324);
and U16951 (N_16951,N_16084,N_16237);
and U16952 (N_16952,N_16116,N_16077);
nor U16953 (N_16953,N_16427,N_16096);
and U16954 (N_16954,N_16004,N_16216);
and U16955 (N_16955,N_16499,N_16068);
nor U16956 (N_16956,N_16440,N_16441);
and U16957 (N_16957,N_16001,N_16051);
nor U16958 (N_16958,N_16463,N_16441);
and U16959 (N_16959,N_16285,N_16387);
nand U16960 (N_16960,N_16267,N_16170);
nor U16961 (N_16961,N_16235,N_16127);
or U16962 (N_16962,N_16086,N_16019);
nor U16963 (N_16963,N_16321,N_16085);
nand U16964 (N_16964,N_16130,N_16387);
or U16965 (N_16965,N_16459,N_16195);
or U16966 (N_16966,N_16134,N_16339);
xnor U16967 (N_16967,N_16124,N_16158);
nor U16968 (N_16968,N_16414,N_16493);
nand U16969 (N_16969,N_16116,N_16053);
or U16970 (N_16970,N_16348,N_16361);
and U16971 (N_16971,N_16407,N_16101);
or U16972 (N_16972,N_16317,N_16431);
and U16973 (N_16973,N_16130,N_16458);
and U16974 (N_16974,N_16490,N_16267);
and U16975 (N_16975,N_16110,N_16052);
xor U16976 (N_16976,N_16420,N_16291);
nand U16977 (N_16977,N_16184,N_16139);
xor U16978 (N_16978,N_16410,N_16101);
or U16979 (N_16979,N_16114,N_16472);
xor U16980 (N_16980,N_16346,N_16188);
xnor U16981 (N_16981,N_16459,N_16194);
nand U16982 (N_16982,N_16251,N_16223);
and U16983 (N_16983,N_16406,N_16416);
and U16984 (N_16984,N_16026,N_16155);
nor U16985 (N_16985,N_16409,N_16109);
and U16986 (N_16986,N_16147,N_16049);
or U16987 (N_16987,N_16340,N_16370);
and U16988 (N_16988,N_16115,N_16151);
nor U16989 (N_16989,N_16247,N_16337);
and U16990 (N_16990,N_16430,N_16080);
and U16991 (N_16991,N_16136,N_16293);
and U16992 (N_16992,N_16463,N_16001);
nor U16993 (N_16993,N_16324,N_16075);
nor U16994 (N_16994,N_16110,N_16439);
nand U16995 (N_16995,N_16049,N_16369);
nor U16996 (N_16996,N_16242,N_16268);
xnor U16997 (N_16997,N_16349,N_16142);
and U16998 (N_16998,N_16023,N_16152);
xnor U16999 (N_16999,N_16372,N_16368);
xnor U17000 (N_17000,N_16674,N_16988);
nor U17001 (N_17001,N_16881,N_16862);
nand U17002 (N_17002,N_16591,N_16773);
and U17003 (N_17003,N_16909,N_16868);
nor U17004 (N_17004,N_16621,N_16893);
or U17005 (N_17005,N_16628,N_16701);
or U17006 (N_17006,N_16923,N_16627);
and U17007 (N_17007,N_16814,N_16839);
xnor U17008 (N_17008,N_16683,N_16896);
nand U17009 (N_17009,N_16960,N_16800);
xor U17010 (N_17010,N_16920,N_16759);
xor U17011 (N_17011,N_16999,N_16757);
nand U17012 (N_17012,N_16594,N_16662);
and U17013 (N_17013,N_16753,N_16581);
or U17014 (N_17014,N_16982,N_16520);
nand U17015 (N_17015,N_16687,N_16637);
and U17016 (N_17016,N_16981,N_16825);
xnor U17017 (N_17017,N_16643,N_16663);
and U17018 (N_17018,N_16842,N_16978);
or U17019 (N_17019,N_16721,N_16714);
and U17020 (N_17020,N_16750,N_16776);
or U17021 (N_17021,N_16866,N_16899);
or U17022 (N_17022,N_16613,N_16538);
or U17023 (N_17023,N_16642,N_16877);
or U17024 (N_17024,N_16994,N_16617);
and U17025 (N_17025,N_16871,N_16578);
xnor U17026 (N_17026,N_16552,N_16908);
and U17027 (N_17027,N_16506,N_16824);
nand U17028 (N_17028,N_16681,N_16857);
nand U17029 (N_17029,N_16522,N_16525);
nor U17030 (N_17030,N_16571,N_16883);
nand U17031 (N_17031,N_16537,N_16992);
nor U17032 (N_17032,N_16837,N_16726);
and U17033 (N_17033,N_16927,N_16751);
nand U17034 (N_17034,N_16943,N_16577);
nand U17035 (N_17035,N_16963,N_16924);
and U17036 (N_17036,N_16508,N_16942);
xor U17037 (N_17037,N_16616,N_16641);
or U17038 (N_17038,N_16954,N_16778);
xor U17039 (N_17039,N_16730,N_16622);
nand U17040 (N_17040,N_16534,N_16772);
and U17041 (N_17041,N_16907,N_16712);
or U17042 (N_17042,N_16809,N_16579);
nand U17043 (N_17043,N_16848,N_16610);
xnor U17044 (N_17044,N_16567,N_16802);
and U17045 (N_17045,N_16900,N_16913);
nor U17046 (N_17046,N_16922,N_16715);
or U17047 (N_17047,N_16931,N_16740);
or U17048 (N_17048,N_16859,N_16786);
nand U17049 (N_17049,N_16647,N_16864);
nand U17050 (N_17050,N_16636,N_16638);
or U17051 (N_17051,N_16890,N_16820);
nor U17052 (N_17052,N_16656,N_16554);
nor U17053 (N_17053,N_16729,N_16706);
or U17054 (N_17054,N_16659,N_16555);
and U17055 (N_17055,N_16665,N_16504);
xnor U17056 (N_17056,N_16798,N_16744);
nand U17057 (N_17057,N_16535,N_16523);
nand U17058 (N_17058,N_16971,N_16546);
and U17059 (N_17059,N_16669,N_16884);
nand U17060 (N_17060,N_16606,N_16852);
or U17061 (N_17061,N_16598,N_16704);
nand U17062 (N_17062,N_16791,N_16697);
or U17063 (N_17063,N_16536,N_16965);
xnor U17064 (N_17064,N_16664,N_16716);
xor U17065 (N_17065,N_16768,N_16856);
or U17066 (N_17066,N_16583,N_16836);
nor U17067 (N_17067,N_16724,N_16689);
xor U17068 (N_17068,N_16516,N_16782);
and U17069 (N_17069,N_16911,N_16765);
xor U17070 (N_17070,N_16833,N_16897);
and U17071 (N_17071,N_16929,N_16692);
xor U17072 (N_17072,N_16671,N_16595);
or U17073 (N_17073,N_16544,N_16708);
and U17074 (N_17074,N_16901,N_16898);
xnor U17075 (N_17075,N_16763,N_16645);
or U17076 (N_17076,N_16758,N_16957);
or U17077 (N_17077,N_16530,N_16733);
nand U17078 (N_17078,N_16737,N_16804);
and U17079 (N_17079,N_16964,N_16873);
or U17080 (N_17080,N_16743,N_16815);
or U17081 (N_17081,N_16570,N_16604);
and U17082 (N_17082,N_16834,N_16531);
or U17083 (N_17083,N_16686,N_16983);
xor U17084 (N_17084,N_16962,N_16853);
nand U17085 (N_17085,N_16514,N_16867);
or U17086 (N_17086,N_16625,N_16783);
xnor U17087 (N_17087,N_16817,N_16756);
nor U17088 (N_17088,N_16799,N_16949);
and U17089 (N_17089,N_16831,N_16886);
or U17090 (N_17090,N_16549,N_16989);
and U17091 (N_17091,N_16912,N_16958);
or U17092 (N_17092,N_16934,N_16775);
xor U17093 (N_17093,N_16917,N_16905);
nand U17094 (N_17094,N_16832,N_16592);
or U17095 (N_17095,N_16707,N_16533);
and U17096 (N_17096,N_16600,N_16736);
and U17097 (N_17097,N_16795,N_16559);
nor U17098 (N_17098,N_16878,N_16543);
and U17099 (N_17099,N_16967,N_16792);
or U17100 (N_17100,N_16532,N_16602);
and U17101 (N_17101,N_16585,N_16780);
and U17102 (N_17102,N_16705,N_16847);
nor U17103 (N_17103,N_16588,N_16888);
or U17104 (N_17104,N_16560,N_16657);
and U17105 (N_17105,N_16572,N_16732);
nor U17106 (N_17106,N_16891,N_16822);
nand U17107 (N_17107,N_16630,N_16972);
nor U17108 (N_17108,N_16937,N_16614);
xor U17109 (N_17109,N_16728,N_16894);
and U17110 (N_17110,N_16823,N_16915);
nand U17111 (N_17111,N_16906,N_16882);
or U17112 (N_17112,N_16722,N_16648);
nor U17113 (N_17113,N_16690,N_16698);
nand U17114 (N_17114,N_16797,N_16626);
and U17115 (N_17115,N_16519,N_16688);
nand U17116 (N_17116,N_16518,N_16904);
or U17117 (N_17117,N_16762,N_16609);
nand U17118 (N_17118,N_16528,N_16974);
or U17119 (N_17119,N_16682,N_16841);
or U17120 (N_17120,N_16826,N_16968);
nand U17121 (N_17121,N_16576,N_16945);
or U17122 (N_17122,N_16872,N_16580);
and U17123 (N_17123,N_16670,N_16819);
nand U17124 (N_17124,N_16653,N_16774);
xnor U17125 (N_17125,N_16589,N_16603);
nor U17126 (N_17126,N_16785,N_16874);
nor U17127 (N_17127,N_16869,N_16876);
xnor U17128 (N_17128,N_16887,N_16961);
xnor U17129 (N_17129,N_16747,N_16649);
nand U17130 (N_17130,N_16755,N_16738);
xnor U17131 (N_17131,N_16505,N_16952);
or U17132 (N_17132,N_16524,N_16562);
nor U17133 (N_17133,N_16540,N_16879);
nand U17134 (N_17134,N_16838,N_16527);
and U17135 (N_17135,N_16749,N_16752);
nand U17136 (N_17136,N_16955,N_16608);
nand U17137 (N_17137,N_16517,N_16655);
and U17138 (N_17138,N_16596,N_16510);
and U17139 (N_17139,N_16851,N_16921);
and U17140 (N_17140,N_16644,N_16928);
or U17141 (N_17141,N_16620,N_16634);
xor U17142 (N_17142,N_16807,N_16599);
xor U17143 (N_17143,N_16850,N_16590);
and U17144 (N_17144,N_16702,N_16902);
and U17145 (N_17145,N_16816,N_16813);
or U17146 (N_17146,N_16830,N_16985);
nand U17147 (N_17147,N_16631,N_16991);
nor U17148 (N_17148,N_16569,N_16574);
xnor U17149 (N_17149,N_16582,N_16511);
or U17150 (N_17150,N_16501,N_16639);
nor U17151 (N_17151,N_16684,N_16710);
or U17152 (N_17152,N_16863,N_16548);
xnor U17153 (N_17153,N_16916,N_16997);
nand U17154 (N_17154,N_16660,N_16935);
or U17155 (N_17155,N_16623,N_16512);
and U17156 (N_17156,N_16810,N_16844);
or U17157 (N_17157,N_16784,N_16561);
nand U17158 (N_17158,N_16742,N_16767);
nand U17159 (N_17159,N_16564,N_16885);
or U17160 (N_17160,N_16746,N_16666);
or U17161 (N_17161,N_16933,N_16880);
and U17162 (N_17162,N_16969,N_16950);
nand U17163 (N_17163,N_16845,N_16947);
and U17164 (N_17164,N_16547,N_16612);
xor U17165 (N_17165,N_16938,N_16858);
or U17166 (N_17166,N_16761,N_16607);
nor U17167 (N_17167,N_16805,N_16860);
and U17168 (N_17168,N_16727,N_16551);
xnor U17169 (N_17169,N_16586,N_16948);
nor U17170 (N_17170,N_16593,N_16629);
nor U17171 (N_17171,N_16951,N_16875);
or U17172 (N_17172,N_16731,N_16640);
or U17173 (N_17173,N_16944,N_16781);
nor U17174 (N_17174,N_16624,N_16667);
xnor U17175 (N_17175,N_16529,N_16801);
and U17176 (N_17176,N_16500,N_16717);
xor U17177 (N_17177,N_16793,N_16679);
nand U17178 (N_17178,N_16652,N_16680);
nor U17179 (N_17179,N_16827,N_16846);
or U17180 (N_17180,N_16998,N_16502);
xnor U17181 (N_17181,N_16696,N_16914);
or U17182 (N_17182,N_16711,N_16691);
or U17183 (N_17183,N_16796,N_16986);
or U17184 (N_17184,N_16700,N_16840);
nand U17185 (N_17185,N_16849,N_16658);
nor U17186 (N_17186,N_16777,N_16760);
nor U17187 (N_17187,N_16587,N_16632);
nand U17188 (N_17188,N_16790,N_16789);
xnor U17189 (N_17189,N_16720,N_16995);
nand U17190 (N_17190,N_16668,N_16558);
or U17191 (N_17191,N_16745,N_16990);
nand U17192 (N_17192,N_16723,N_16739);
or U17193 (N_17193,N_16672,N_16806);
or U17194 (N_17194,N_16936,N_16787);
xor U17195 (N_17195,N_16811,N_16771);
or U17196 (N_17196,N_16584,N_16557);
and U17197 (N_17197,N_16503,N_16829);
or U17198 (N_17198,N_16970,N_16735);
and U17199 (N_17199,N_16979,N_16966);
or U17200 (N_17200,N_16939,N_16910);
xor U17201 (N_17201,N_16895,N_16977);
and U17202 (N_17202,N_16889,N_16993);
or U17203 (N_17203,N_16940,N_16946);
nand U17204 (N_17204,N_16521,N_16654);
xor U17205 (N_17205,N_16861,N_16821);
nand U17206 (N_17206,N_16605,N_16694);
nand U17207 (N_17207,N_16892,N_16925);
or U17208 (N_17208,N_16545,N_16601);
nand U17209 (N_17209,N_16812,N_16828);
and U17210 (N_17210,N_16865,N_16918);
xor U17211 (N_17211,N_16741,N_16646);
xnor U17212 (N_17212,N_16926,N_16513);
nand U17213 (N_17213,N_16676,N_16855);
xnor U17214 (N_17214,N_16854,N_16734);
nand U17215 (N_17215,N_16615,N_16770);
or U17216 (N_17216,N_16673,N_16973);
or U17217 (N_17217,N_16987,N_16542);
nor U17218 (N_17218,N_16541,N_16699);
nor U17219 (N_17219,N_16769,N_16633);
nor U17220 (N_17220,N_16685,N_16651);
or U17221 (N_17221,N_16553,N_16930);
or U17222 (N_17222,N_16843,N_16619);
xnor U17223 (N_17223,N_16803,N_16718);
and U17224 (N_17224,N_16919,N_16515);
and U17225 (N_17225,N_16635,N_16566);
nor U17226 (N_17226,N_16788,N_16748);
xor U17227 (N_17227,N_16611,N_16941);
nand U17228 (N_17228,N_16563,N_16509);
and U17229 (N_17229,N_16956,N_16932);
or U17230 (N_17230,N_16678,N_16835);
xor U17231 (N_17231,N_16675,N_16975);
xnor U17232 (N_17232,N_16808,N_16539);
xor U17233 (N_17233,N_16996,N_16764);
xor U17234 (N_17234,N_16779,N_16695);
and U17235 (N_17235,N_16976,N_16794);
or U17236 (N_17236,N_16984,N_16713);
xor U17237 (N_17237,N_16903,N_16618);
or U17238 (N_17238,N_16677,N_16959);
or U17239 (N_17239,N_16568,N_16507);
and U17240 (N_17240,N_16597,N_16693);
or U17241 (N_17241,N_16650,N_16980);
nor U17242 (N_17242,N_16818,N_16709);
and U17243 (N_17243,N_16526,N_16556);
nor U17244 (N_17244,N_16870,N_16766);
and U17245 (N_17245,N_16550,N_16661);
nand U17246 (N_17246,N_16725,N_16719);
or U17247 (N_17247,N_16703,N_16575);
nand U17248 (N_17248,N_16953,N_16573);
and U17249 (N_17249,N_16754,N_16565);
xnor U17250 (N_17250,N_16838,N_16871);
and U17251 (N_17251,N_16915,N_16564);
or U17252 (N_17252,N_16978,N_16640);
nor U17253 (N_17253,N_16515,N_16816);
or U17254 (N_17254,N_16675,N_16591);
or U17255 (N_17255,N_16745,N_16700);
or U17256 (N_17256,N_16788,N_16877);
and U17257 (N_17257,N_16537,N_16603);
or U17258 (N_17258,N_16865,N_16979);
nand U17259 (N_17259,N_16547,N_16961);
or U17260 (N_17260,N_16548,N_16596);
xor U17261 (N_17261,N_16781,N_16799);
or U17262 (N_17262,N_16622,N_16925);
xnor U17263 (N_17263,N_16618,N_16670);
nor U17264 (N_17264,N_16740,N_16581);
nor U17265 (N_17265,N_16644,N_16773);
nand U17266 (N_17266,N_16736,N_16560);
nor U17267 (N_17267,N_16585,N_16704);
xor U17268 (N_17268,N_16868,N_16836);
nand U17269 (N_17269,N_16562,N_16885);
xor U17270 (N_17270,N_16598,N_16543);
nand U17271 (N_17271,N_16869,N_16843);
or U17272 (N_17272,N_16908,N_16981);
xnor U17273 (N_17273,N_16774,N_16582);
and U17274 (N_17274,N_16560,N_16809);
nor U17275 (N_17275,N_16661,N_16668);
xor U17276 (N_17276,N_16680,N_16962);
or U17277 (N_17277,N_16876,N_16757);
nand U17278 (N_17278,N_16602,N_16820);
or U17279 (N_17279,N_16804,N_16758);
nor U17280 (N_17280,N_16703,N_16777);
xnor U17281 (N_17281,N_16924,N_16835);
and U17282 (N_17282,N_16582,N_16911);
nand U17283 (N_17283,N_16710,N_16819);
nand U17284 (N_17284,N_16983,N_16601);
and U17285 (N_17285,N_16793,N_16596);
and U17286 (N_17286,N_16596,N_16648);
xor U17287 (N_17287,N_16560,N_16891);
or U17288 (N_17288,N_16638,N_16803);
nor U17289 (N_17289,N_16948,N_16850);
and U17290 (N_17290,N_16846,N_16857);
nor U17291 (N_17291,N_16664,N_16646);
nor U17292 (N_17292,N_16878,N_16506);
or U17293 (N_17293,N_16750,N_16747);
and U17294 (N_17294,N_16631,N_16553);
and U17295 (N_17295,N_16885,N_16963);
nand U17296 (N_17296,N_16625,N_16927);
or U17297 (N_17297,N_16911,N_16549);
or U17298 (N_17298,N_16569,N_16957);
xnor U17299 (N_17299,N_16724,N_16631);
xor U17300 (N_17300,N_16875,N_16532);
and U17301 (N_17301,N_16556,N_16899);
nor U17302 (N_17302,N_16915,N_16894);
xnor U17303 (N_17303,N_16876,N_16867);
and U17304 (N_17304,N_16878,N_16660);
xor U17305 (N_17305,N_16754,N_16637);
xor U17306 (N_17306,N_16915,N_16682);
nand U17307 (N_17307,N_16697,N_16795);
or U17308 (N_17308,N_16562,N_16635);
and U17309 (N_17309,N_16966,N_16629);
nor U17310 (N_17310,N_16977,N_16952);
xnor U17311 (N_17311,N_16630,N_16914);
nand U17312 (N_17312,N_16718,N_16604);
nor U17313 (N_17313,N_16828,N_16738);
nor U17314 (N_17314,N_16990,N_16840);
and U17315 (N_17315,N_16657,N_16805);
nand U17316 (N_17316,N_16779,N_16842);
nand U17317 (N_17317,N_16637,N_16557);
nor U17318 (N_17318,N_16916,N_16649);
nor U17319 (N_17319,N_16767,N_16828);
and U17320 (N_17320,N_16896,N_16703);
nand U17321 (N_17321,N_16987,N_16596);
and U17322 (N_17322,N_16722,N_16596);
nor U17323 (N_17323,N_16562,N_16508);
nand U17324 (N_17324,N_16566,N_16584);
nand U17325 (N_17325,N_16564,N_16844);
and U17326 (N_17326,N_16674,N_16710);
nor U17327 (N_17327,N_16665,N_16689);
nand U17328 (N_17328,N_16900,N_16670);
nand U17329 (N_17329,N_16688,N_16742);
and U17330 (N_17330,N_16892,N_16968);
and U17331 (N_17331,N_16931,N_16980);
nand U17332 (N_17332,N_16826,N_16691);
nor U17333 (N_17333,N_16843,N_16671);
xor U17334 (N_17334,N_16774,N_16573);
and U17335 (N_17335,N_16813,N_16829);
nand U17336 (N_17336,N_16698,N_16931);
nor U17337 (N_17337,N_16630,N_16564);
and U17338 (N_17338,N_16901,N_16605);
nand U17339 (N_17339,N_16563,N_16654);
nand U17340 (N_17340,N_16518,N_16993);
or U17341 (N_17341,N_16972,N_16891);
or U17342 (N_17342,N_16942,N_16616);
nor U17343 (N_17343,N_16655,N_16938);
or U17344 (N_17344,N_16916,N_16646);
and U17345 (N_17345,N_16663,N_16897);
or U17346 (N_17346,N_16939,N_16782);
nand U17347 (N_17347,N_16686,N_16733);
and U17348 (N_17348,N_16912,N_16673);
or U17349 (N_17349,N_16638,N_16613);
or U17350 (N_17350,N_16589,N_16838);
nand U17351 (N_17351,N_16563,N_16613);
nor U17352 (N_17352,N_16651,N_16989);
nor U17353 (N_17353,N_16792,N_16945);
nand U17354 (N_17354,N_16802,N_16652);
xor U17355 (N_17355,N_16871,N_16687);
xnor U17356 (N_17356,N_16708,N_16745);
xnor U17357 (N_17357,N_16908,N_16809);
or U17358 (N_17358,N_16759,N_16872);
and U17359 (N_17359,N_16812,N_16721);
or U17360 (N_17360,N_16679,N_16714);
or U17361 (N_17361,N_16610,N_16520);
nor U17362 (N_17362,N_16820,N_16628);
and U17363 (N_17363,N_16767,N_16686);
or U17364 (N_17364,N_16723,N_16908);
nand U17365 (N_17365,N_16527,N_16913);
xnor U17366 (N_17366,N_16933,N_16924);
xor U17367 (N_17367,N_16872,N_16507);
nand U17368 (N_17368,N_16630,N_16735);
xnor U17369 (N_17369,N_16514,N_16946);
nand U17370 (N_17370,N_16588,N_16640);
nand U17371 (N_17371,N_16642,N_16505);
and U17372 (N_17372,N_16700,N_16585);
xor U17373 (N_17373,N_16626,N_16789);
and U17374 (N_17374,N_16703,N_16721);
xor U17375 (N_17375,N_16781,N_16890);
xnor U17376 (N_17376,N_16748,N_16835);
nor U17377 (N_17377,N_16791,N_16962);
nand U17378 (N_17378,N_16882,N_16792);
nand U17379 (N_17379,N_16753,N_16993);
nand U17380 (N_17380,N_16755,N_16742);
nand U17381 (N_17381,N_16997,N_16874);
nor U17382 (N_17382,N_16948,N_16751);
or U17383 (N_17383,N_16637,N_16768);
or U17384 (N_17384,N_16514,N_16565);
nand U17385 (N_17385,N_16744,N_16948);
nand U17386 (N_17386,N_16554,N_16918);
or U17387 (N_17387,N_16892,N_16651);
or U17388 (N_17388,N_16650,N_16685);
and U17389 (N_17389,N_16776,N_16781);
nor U17390 (N_17390,N_16547,N_16893);
nor U17391 (N_17391,N_16929,N_16948);
xnor U17392 (N_17392,N_16583,N_16916);
nor U17393 (N_17393,N_16955,N_16851);
and U17394 (N_17394,N_16570,N_16534);
or U17395 (N_17395,N_16849,N_16785);
and U17396 (N_17396,N_16756,N_16920);
and U17397 (N_17397,N_16801,N_16686);
and U17398 (N_17398,N_16931,N_16861);
nor U17399 (N_17399,N_16858,N_16924);
nand U17400 (N_17400,N_16750,N_16737);
xor U17401 (N_17401,N_16560,N_16803);
nand U17402 (N_17402,N_16699,N_16808);
or U17403 (N_17403,N_16922,N_16899);
and U17404 (N_17404,N_16876,N_16678);
nor U17405 (N_17405,N_16810,N_16690);
xor U17406 (N_17406,N_16817,N_16560);
nor U17407 (N_17407,N_16693,N_16604);
xor U17408 (N_17408,N_16948,N_16613);
xnor U17409 (N_17409,N_16856,N_16675);
and U17410 (N_17410,N_16753,N_16878);
xnor U17411 (N_17411,N_16512,N_16601);
or U17412 (N_17412,N_16500,N_16913);
nor U17413 (N_17413,N_16635,N_16591);
or U17414 (N_17414,N_16893,N_16620);
or U17415 (N_17415,N_16860,N_16883);
nor U17416 (N_17416,N_16944,N_16645);
nor U17417 (N_17417,N_16936,N_16650);
nor U17418 (N_17418,N_16871,N_16888);
nand U17419 (N_17419,N_16538,N_16655);
xor U17420 (N_17420,N_16798,N_16902);
and U17421 (N_17421,N_16896,N_16818);
nor U17422 (N_17422,N_16966,N_16814);
nor U17423 (N_17423,N_16796,N_16556);
xor U17424 (N_17424,N_16678,N_16562);
nor U17425 (N_17425,N_16736,N_16519);
nor U17426 (N_17426,N_16789,N_16694);
and U17427 (N_17427,N_16575,N_16908);
nor U17428 (N_17428,N_16669,N_16952);
nand U17429 (N_17429,N_16750,N_16937);
nand U17430 (N_17430,N_16964,N_16668);
nor U17431 (N_17431,N_16758,N_16887);
and U17432 (N_17432,N_16831,N_16836);
nor U17433 (N_17433,N_16900,N_16663);
nor U17434 (N_17434,N_16891,N_16734);
nor U17435 (N_17435,N_16937,N_16913);
and U17436 (N_17436,N_16701,N_16608);
xnor U17437 (N_17437,N_16906,N_16657);
or U17438 (N_17438,N_16769,N_16772);
xnor U17439 (N_17439,N_16734,N_16678);
nand U17440 (N_17440,N_16682,N_16773);
nand U17441 (N_17441,N_16698,N_16855);
nand U17442 (N_17442,N_16764,N_16538);
nor U17443 (N_17443,N_16684,N_16660);
and U17444 (N_17444,N_16971,N_16956);
nand U17445 (N_17445,N_16660,N_16940);
or U17446 (N_17446,N_16809,N_16878);
xnor U17447 (N_17447,N_16728,N_16669);
or U17448 (N_17448,N_16658,N_16843);
nand U17449 (N_17449,N_16804,N_16510);
or U17450 (N_17450,N_16536,N_16854);
and U17451 (N_17451,N_16716,N_16529);
nor U17452 (N_17452,N_16860,N_16890);
or U17453 (N_17453,N_16514,N_16988);
nand U17454 (N_17454,N_16566,N_16961);
nand U17455 (N_17455,N_16738,N_16613);
or U17456 (N_17456,N_16630,N_16915);
nor U17457 (N_17457,N_16805,N_16727);
or U17458 (N_17458,N_16961,N_16689);
xor U17459 (N_17459,N_16901,N_16964);
or U17460 (N_17460,N_16552,N_16659);
and U17461 (N_17461,N_16840,N_16955);
xor U17462 (N_17462,N_16938,N_16643);
and U17463 (N_17463,N_16770,N_16838);
nor U17464 (N_17464,N_16565,N_16941);
nand U17465 (N_17465,N_16937,N_16696);
or U17466 (N_17466,N_16974,N_16764);
or U17467 (N_17467,N_16938,N_16781);
and U17468 (N_17468,N_16837,N_16723);
nand U17469 (N_17469,N_16898,N_16744);
and U17470 (N_17470,N_16568,N_16804);
and U17471 (N_17471,N_16546,N_16773);
nand U17472 (N_17472,N_16871,N_16659);
and U17473 (N_17473,N_16963,N_16803);
or U17474 (N_17474,N_16613,N_16602);
or U17475 (N_17475,N_16612,N_16764);
or U17476 (N_17476,N_16569,N_16945);
and U17477 (N_17477,N_16808,N_16797);
nor U17478 (N_17478,N_16714,N_16560);
and U17479 (N_17479,N_16562,N_16857);
xor U17480 (N_17480,N_16773,N_16757);
and U17481 (N_17481,N_16652,N_16801);
or U17482 (N_17482,N_16724,N_16526);
nor U17483 (N_17483,N_16614,N_16774);
or U17484 (N_17484,N_16630,N_16572);
nor U17485 (N_17485,N_16590,N_16706);
and U17486 (N_17486,N_16857,N_16651);
or U17487 (N_17487,N_16697,N_16932);
and U17488 (N_17488,N_16873,N_16629);
nand U17489 (N_17489,N_16724,N_16829);
or U17490 (N_17490,N_16990,N_16581);
xor U17491 (N_17491,N_16594,N_16629);
and U17492 (N_17492,N_16678,N_16811);
nand U17493 (N_17493,N_16903,N_16790);
nand U17494 (N_17494,N_16953,N_16889);
nor U17495 (N_17495,N_16535,N_16940);
nor U17496 (N_17496,N_16771,N_16984);
nor U17497 (N_17497,N_16816,N_16536);
or U17498 (N_17498,N_16990,N_16601);
nand U17499 (N_17499,N_16723,N_16893);
xor U17500 (N_17500,N_17424,N_17400);
nor U17501 (N_17501,N_17045,N_17370);
nor U17502 (N_17502,N_17461,N_17005);
nor U17503 (N_17503,N_17310,N_17335);
and U17504 (N_17504,N_17295,N_17163);
nand U17505 (N_17505,N_17206,N_17173);
or U17506 (N_17506,N_17152,N_17377);
nor U17507 (N_17507,N_17275,N_17352);
nand U17508 (N_17508,N_17149,N_17083);
and U17509 (N_17509,N_17479,N_17313);
or U17510 (N_17510,N_17399,N_17175);
xnor U17511 (N_17511,N_17344,N_17081);
and U17512 (N_17512,N_17358,N_17095);
or U17513 (N_17513,N_17302,N_17017);
nor U17514 (N_17514,N_17248,N_17270);
or U17515 (N_17515,N_17201,N_17453);
nand U17516 (N_17516,N_17343,N_17192);
and U17517 (N_17517,N_17429,N_17218);
nor U17518 (N_17518,N_17378,N_17405);
xor U17519 (N_17519,N_17126,N_17334);
nand U17520 (N_17520,N_17187,N_17182);
xnor U17521 (N_17521,N_17008,N_17019);
and U17522 (N_17522,N_17298,N_17268);
and U17523 (N_17523,N_17035,N_17465);
or U17524 (N_17524,N_17483,N_17020);
and U17525 (N_17525,N_17274,N_17109);
and U17526 (N_17526,N_17407,N_17261);
nand U17527 (N_17527,N_17062,N_17427);
nand U17528 (N_17528,N_17203,N_17022);
or U17529 (N_17529,N_17188,N_17354);
or U17530 (N_17530,N_17039,N_17200);
and U17531 (N_17531,N_17194,N_17044);
and U17532 (N_17532,N_17099,N_17070);
or U17533 (N_17533,N_17094,N_17169);
nor U17534 (N_17534,N_17452,N_17100);
and U17535 (N_17535,N_17214,N_17164);
nand U17536 (N_17536,N_17172,N_17260);
and U17537 (N_17537,N_17469,N_17403);
nand U17538 (N_17538,N_17337,N_17167);
xnor U17539 (N_17539,N_17108,N_17107);
xor U17540 (N_17540,N_17345,N_17224);
and U17541 (N_17541,N_17191,N_17307);
nand U17542 (N_17542,N_17208,N_17114);
nand U17543 (N_17543,N_17454,N_17292);
nand U17544 (N_17544,N_17480,N_17135);
nor U17545 (N_17545,N_17066,N_17369);
xnor U17546 (N_17546,N_17332,N_17048);
nand U17547 (N_17547,N_17280,N_17415);
xor U17548 (N_17548,N_17381,N_17490);
xor U17549 (N_17549,N_17336,N_17103);
or U17550 (N_17550,N_17486,N_17477);
nor U17551 (N_17551,N_17087,N_17340);
or U17552 (N_17552,N_17177,N_17325);
and U17553 (N_17553,N_17080,N_17246);
xor U17554 (N_17554,N_17279,N_17142);
xor U17555 (N_17555,N_17009,N_17255);
nand U17556 (N_17556,N_17414,N_17141);
nor U17557 (N_17557,N_17139,N_17096);
or U17558 (N_17558,N_17316,N_17385);
nand U17559 (N_17559,N_17349,N_17320);
xnor U17560 (N_17560,N_17197,N_17168);
xnor U17561 (N_17561,N_17092,N_17195);
nor U17562 (N_17562,N_17140,N_17128);
and U17563 (N_17563,N_17371,N_17386);
or U17564 (N_17564,N_17374,N_17338);
xnor U17565 (N_17565,N_17402,N_17211);
nand U17566 (N_17566,N_17301,N_17283);
nor U17567 (N_17567,N_17365,N_17276);
and U17568 (N_17568,N_17122,N_17217);
or U17569 (N_17569,N_17159,N_17263);
or U17570 (N_17570,N_17321,N_17312);
nor U17571 (N_17571,N_17055,N_17226);
nand U17572 (N_17572,N_17053,N_17382);
xnor U17573 (N_17573,N_17034,N_17420);
xor U17574 (N_17574,N_17278,N_17038);
nand U17575 (N_17575,N_17216,N_17106);
and U17576 (N_17576,N_17129,N_17198);
nand U17577 (N_17577,N_17183,N_17498);
or U17578 (N_17578,N_17499,N_17487);
and U17579 (N_17579,N_17137,N_17131);
nand U17580 (N_17580,N_17079,N_17394);
nor U17581 (N_17581,N_17372,N_17071);
and U17582 (N_17582,N_17445,N_17076);
and U17583 (N_17583,N_17286,N_17303);
and U17584 (N_17584,N_17431,N_17239);
xor U17585 (N_17585,N_17236,N_17488);
and U17586 (N_17586,N_17401,N_17121);
nor U17587 (N_17587,N_17077,N_17267);
or U17588 (N_17588,N_17375,N_17254);
or U17589 (N_17589,N_17388,N_17161);
nor U17590 (N_17590,N_17379,N_17311);
or U17591 (N_17591,N_17481,N_17018);
and U17592 (N_17592,N_17288,N_17281);
or U17593 (N_17593,N_17342,N_17051);
nand U17594 (N_17594,N_17470,N_17266);
nand U17595 (N_17595,N_17457,N_17423);
or U17596 (N_17596,N_17025,N_17392);
nor U17597 (N_17597,N_17015,N_17130);
nor U17598 (N_17598,N_17251,N_17398);
xnor U17599 (N_17599,N_17024,N_17212);
nand U17600 (N_17600,N_17115,N_17496);
nor U17601 (N_17601,N_17491,N_17190);
xnor U17602 (N_17602,N_17240,N_17433);
nor U17603 (N_17603,N_17287,N_17075);
nand U17604 (N_17604,N_17117,N_17213);
xor U17605 (N_17605,N_17178,N_17442);
xnor U17606 (N_17606,N_17444,N_17012);
or U17607 (N_17607,N_17146,N_17492);
and U17608 (N_17608,N_17359,N_17404);
and U17609 (N_17609,N_17348,N_17258);
nor U17610 (N_17610,N_17319,N_17324);
or U17611 (N_17611,N_17184,N_17305);
and U17612 (N_17612,N_17458,N_17223);
nor U17613 (N_17613,N_17351,N_17418);
or U17614 (N_17614,N_17186,N_17339);
nor U17615 (N_17615,N_17489,N_17057);
xnor U17616 (N_17616,N_17027,N_17028);
nand U17617 (N_17617,N_17361,N_17228);
nand U17618 (N_17618,N_17067,N_17315);
nand U17619 (N_17619,N_17450,N_17393);
nor U17620 (N_17620,N_17265,N_17383);
nor U17621 (N_17621,N_17373,N_17277);
and U17622 (N_17622,N_17410,N_17043);
or U17623 (N_17623,N_17185,N_17065);
nand U17624 (N_17624,N_17082,N_17396);
xnor U17625 (N_17625,N_17170,N_17180);
or U17626 (N_17626,N_17189,N_17150);
nand U17627 (N_17627,N_17237,N_17259);
xor U17628 (N_17628,N_17001,N_17063);
and U17629 (N_17629,N_17026,N_17304);
or U17630 (N_17630,N_17437,N_17143);
nor U17631 (N_17631,N_17322,N_17000);
or U17632 (N_17632,N_17293,N_17422);
nor U17633 (N_17633,N_17032,N_17448);
nor U17634 (N_17634,N_17390,N_17368);
nor U17635 (N_17635,N_17089,N_17033);
nor U17636 (N_17636,N_17451,N_17078);
xor U17637 (N_17637,N_17329,N_17074);
nand U17638 (N_17638,N_17171,N_17272);
nor U17639 (N_17639,N_17050,N_17456);
xnor U17640 (N_17640,N_17289,N_17419);
nand U17641 (N_17641,N_17475,N_17196);
and U17642 (N_17642,N_17157,N_17459);
nand U17643 (N_17643,N_17238,N_17367);
nor U17644 (N_17644,N_17314,N_17417);
and U17645 (N_17645,N_17284,N_17412);
xor U17646 (N_17646,N_17006,N_17125);
nor U17647 (N_17647,N_17341,N_17235);
nand U17648 (N_17648,N_17257,N_17040);
nor U17649 (N_17649,N_17269,N_17347);
or U17650 (N_17650,N_17124,N_17306);
nor U17651 (N_17651,N_17064,N_17209);
nand U17652 (N_17652,N_17318,N_17440);
nor U17653 (N_17653,N_17123,N_17256);
nand U17654 (N_17654,N_17250,N_17273);
xnor U17655 (N_17655,N_17030,N_17085);
and U17656 (N_17656,N_17068,N_17473);
nor U17657 (N_17657,N_17430,N_17007);
and U17658 (N_17658,N_17363,N_17253);
xnor U17659 (N_17659,N_17059,N_17029);
nor U17660 (N_17660,N_17148,N_17154);
and U17661 (N_17661,N_17054,N_17013);
or U17662 (N_17662,N_17447,N_17482);
and U17663 (N_17663,N_17432,N_17136);
nand U17664 (N_17664,N_17225,N_17326);
and U17665 (N_17665,N_17478,N_17247);
xor U17666 (N_17666,N_17449,N_17041);
nand U17667 (N_17667,N_17290,N_17147);
nand U17668 (N_17668,N_17158,N_17144);
and U17669 (N_17669,N_17497,N_17474);
and U17670 (N_17670,N_17090,N_17476);
nor U17671 (N_17671,N_17021,N_17436);
and U17672 (N_17672,N_17389,N_17357);
nor U17673 (N_17673,N_17471,N_17110);
nor U17674 (N_17674,N_17134,N_17016);
nand U17675 (N_17675,N_17252,N_17221);
nor U17676 (N_17676,N_17468,N_17127);
and U17677 (N_17677,N_17297,N_17317);
or U17678 (N_17678,N_17036,N_17262);
or U17679 (N_17679,N_17084,N_17485);
or U17680 (N_17680,N_17362,N_17160);
or U17681 (N_17681,N_17463,N_17384);
nor U17682 (N_17682,N_17181,N_17133);
nand U17683 (N_17683,N_17439,N_17413);
nand U17684 (N_17684,N_17309,N_17495);
nor U17685 (N_17685,N_17004,N_17222);
xnor U17686 (N_17686,N_17231,N_17409);
and U17687 (N_17687,N_17132,N_17219);
and U17688 (N_17688,N_17434,N_17031);
nand U17689 (N_17689,N_17176,N_17072);
xor U17690 (N_17690,N_17119,N_17091);
nand U17691 (N_17691,N_17460,N_17162);
nor U17692 (N_17692,N_17355,N_17230);
xnor U17693 (N_17693,N_17042,N_17155);
or U17694 (N_17694,N_17330,N_17138);
nor U17695 (N_17695,N_17294,N_17056);
and U17696 (N_17696,N_17353,N_17174);
xor U17697 (N_17697,N_17073,N_17421);
xor U17698 (N_17698,N_17300,N_17153);
nor U17699 (N_17699,N_17333,N_17202);
nor U17700 (N_17700,N_17364,N_17443);
nor U17701 (N_17701,N_17455,N_17233);
and U17702 (N_17702,N_17210,N_17244);
nor U17703 (N_17703,N_17484,N_17060);
xnor U17704 (N_17704,N_17111,N_17299);
or U17705 (N_17705,N_17058,N_17166);
or U17706 (N_17706,N_17003,N_17098);
and U17707 (N_17707,N_17199,N_17291);
nor U17708 (N_17708,N_17061,N_17088);
xnor U17709 (N_17709,N_17296,N_17446);
or U17710 (N_17710,N_17380,N_17052);
and U17711 (N_17711,N_17086,N_17493);
and U17712 (N_17712,N_17494,N_17113);
nand U17713 (N_17713,N_17102,N_17408);
or U17714 (N_17714,N_17411,N_17112);
nor U17715 (N_17715,N_17438,N_17328);
nand U17716 (N_17716,N_17425,N_17014);
xor U17717 (N_17717,N_17428,N_17387);
or U17718 (N_17718,N_17145,N_17069);
or U17719 (N_17719,N_17366,N_17151);
nand U17720 (N_17720,N_17205,N_17243);
and U17721 (N_17721,N_17323,N_17207);
or U17722 (N_17722,N_17331,N_17245);
or U17723 (N_17723,N_17232,N_17441);
xor U17724 (N_17724,N_17093,N_17464);
or U17725 (N_17725,N_17120,N_17467);
or U17726 (N_17726,N_17327,N_17118);
or U17727 (N_17727,N_17397,N_17010);
xnor U17728 (N_17728,N_17047,N_17229);
and U17729 (N_17729,N_17011,N_17241);
nand U17730 (N_17730,N_17376,N_17360);
and U17731 (N_17731,N_17104,N_17356);
xnor U17732 (N_17732,N_17116,N_17308);
xnor U17733 (N_17733,N_17234,N_17466);
or U17734 (N_17734,N_17350,N_17165);
nor U17735 (N_17735,N_17156,N_17193);
nand U17736 (N_17736,N_17406,N_17220);
nor U17737 (N_17737,N_17204,N_17416);
and U17738 (N_17738,N_17282,N_17264);
nand U17739 (N_17739,N_17462,N_17242);
and U17740 (N_17740,N_17037,N_17391);
xnor U17741 (N_17741,N_17049,N_17179);
nand U17742 (N_17742,N_17346,N_17395);
xor U17743 (N_17743,N_17227,N_17101);
nand U17744 (N_17744,N_17097,N_17426);
xnor U17745 (N_17745,N_17105,N_17472);
nand U17746 (N_17746,N_17285,N_17435);
and U17747 (N_17747,N_17002,N_17271);
nor U17748 (N_17748,N_17215,N_17249);
nand U17749 (N_17749,N_17023,N_17046);
and U17750 (N_17750,N_17048,N_17014);
or U17751 (N_17751,N_17046,N_17126);
or U17752 (N_17752,N_17259,N_17474);
xnor U17753 (N_17753,N_17355,N_17363);
nor U17754 (N_17754,N_17010,N_17246);
or U17755 (N_17755,N_17001,N_17115);
xor U17756 (N_17756,N_17456,N_17166);
and U17757 (N_17757,N_17030,N_17392);
nor U17758 (N_17758,N_17164,N_17270);
xnor U17759 (N_17759,N_17410,N_17348);
nor U17760 (N_17760,N_17258,N_17425);
or U17761 (N_17761,N_17353,N_17469);
nor U17762 (N_17762,N_17233,N_17144);
and U17763 (N_17763,N_17458,N_17461);
nor U17764 (N_17764,N_17151,N_17123);
or U17765 (N_17765,N_17297,N_17433);
nand U17766 (N_17766,N_17139,N_17067);
or U17767 (N_17767,N_17037,N_17371);
and U17768 (N_17768,N_17446,N_17106);
or U17769 (N_17769,N_17260,N_17479);
nand U17770 (N_17770,N_17314,N_17068);
nand U17771 (N_17771,N_17080,N_17103);
xor U17772 (N_17772,N_17423,N_17194);
or U17773 (N_17773,N_17210,N_17006);
or U17774 (N_17774,N_17447,N_17097);
nor U17775 (N_17775,N_17151,N_17247);
nand U17776 (N_17776,N_17031,N_17159);
xnor U17777 (N_17777,N_17001,N_17253);
xor U17778 (N_17778,N_17356,N_17488);
nor U17779 (N_17779,N_17125,N_17009);
or U17780 (N_17780,N_17192,N_17275);
or U17781 (N_17781,N_17126,N_17295);
and U17782 (N_17782,N_17329,N_17252);
nor U17783 (N_17783,N_17430,N_17084);
nand U17784 (N_17784,N_17371,N_17403);
and U17785 (N_17785,N_17326,N_17177);
or U17786 (N_17786,N_17255,N_17170);
nand U17787 (N_17787,N_17469,N_17233);
or U17788 (N_17788,N_17201,N_17038);
and U17789 (N_17789,N_17391,N_17076);
and U17790 (N_17790,N_17128,N_17324);
and U17791 (N_17791,N_17365,N_17480);
nand U17792 (N_17792,N_17195,N_17387);
xnor U17793 (N_17793,N_17152,N_17292);
nor U17794 (N_17794,N_17339,N_17267);
and U17795 (N_17795,N_17026,N_17309);
nor U17796 (N_17796,N_17326,N_17405);
xor U17797 (N_17797,N_17257,N_17094);
and U17798 (N_17798,N_17103,N_17124);
nand U17799 (N_17799,N_17132,N_17442);
or U17800 (N_17800,N_17117,N_17450);
nand U17801 (N_17801,N_17155,N_17153);
or U17802 (N_17802,N_17134,N_17247);
xnor U17803 (N_17803,N_17474,N_17046);
xor U17804 (N_17804,N_17031,N_17060);
and U17805 (N_17805,N_17120,N_17351);
and U17806 (N_17806,N_17195,N_17439);
nand U17807 (N_17807,N_17108,N_17280);
or U17808 (N_17808,N_17366,N_17415);
or U17809 (N_17809,N_17071,N_17217);
nor U17810 (N_17810,N_17079,N_17149);
or U17811 (N_17811,N_17079,N_17047);
or U17812 (N_17812,N_17116,N_17112);
nor U17813 (N_17813,N_17004,N_17456);
or U17814 (N_17814,N_17029,N_17403);
and U17815 (N_17815,N_17029,N_17275);
and U17816 (N_17816,N_17214,N_17104);
and U17817 (N_17817,N_17210,N_17317);
or U17818 (N_17818,N_17358,N_17470);
nor U17819 (N_17819,N_17380,N_17154);
nand U17820 (N_17820,N_17084,N_17044);
nor U17821 (N_17821,N_17488,N_17093);
and U17822 (N_17822,N_17221,N_17093);
nor U17823 (N_17823,N_17252,N_17043);
and U17824 (N_17824,N_17397,N_17455);
nand U17825 (N_17825,N_17315,N_17496);
or U17826 (N_17826,N_17333,N_17329);
and U17827 (N_17827,N_17181,N_17382);
or U17828 (N_17828,N_17383,N_17211);
or U17829 (N_17829,N_17231,N_17016);
xnor U17830 (N_17830,N_17375,N_17367);
or U17831 (N_17831,N_17222,N_17310);
nor U17832 (N_17832,N_17271,N_17344);
or U17833 (N_17833,N_17404,N_17329);
nor U17834 (N_17834,N_17010,N_17434);
and U17835 (N_17835,N_17457,N_17187);
or U17836 (N_17836,N_17480,N_17063);
nand U17837 (N_17837,N_17270,N_17144);
nor U17838 (N_17838,N_17084,N_17281);
and U17839 (N_17839,N_17467,N_17201);
or U17840 (N_17840,N_17290,N_17437);
and U17841 (N_17841,N_17476,N_17357);
xor U17842 (N_17842,N_17307,N_17267);
nor U17843 (N_17843,N_17347,N_17253);
xor U17844 (N_17844,N_17436,N_17190);
nand U17845 (N_17845,N_17033,N_17314);
and U17846 (N_17846,N_17030,N_17459);
and U17847 (N_17847,N_17160,N_17145);
nand U17848 (N_17848,N_17080,N_17303);
or U17849 (N_17849,N_17073,N_17066);
xor U17850 (N_17850,N_17319,N_17334);
nand U17851 (N_17851,N_17485,N_17299);
nor U17852 (N_17852,N_17201,N_17100);
xnor U17853 (N_17853,N_17237,N_17169);
xnor U17854 (N_17854,N_17399,N_17432);
xnor U17855 (N_17855,N_17046,N_17294);
nor U17856 (N_17856,N_17482,N_17130);
or U17857 (N_17857,N_17118,N_17399);
or U17858 (N_17858,N_17404,N_17240);
nor U17859 (N_17859,N_17458,N_17182);
xnor U17860 (N_17860,N_17090,N_17340);
nand U17861 (N_17861,N_17143,N_17317);
nor U17862 (N_17862,N_17273,N_17086);
xor U17863 (N_17863,N_17476,N_17450);
or U17864 (N_17864,N_17292,N_17103);
xor U17865 (N_17865,N_17007,N_17300);
nand U17866 (N_17866,N_17210,N_17051);
and U17867 (N_17867,N_17390,N_17188);
and U17868 (N_17868,N_17391,N_17045);
and U17869 (N_17869,N_17435,N_17482);
and U17870 (N_17870,N_17121,N_17017);
xor U17871 (N_17871,N_17316,N_17005);
and U17872 (N_17872,N_17478,N_17110);
nor U17873 (N_17873,N_17204,N_17098);
nor U17874 (N_17874,N_17448,N_17332);
or U17875 (N_17875,N_17220,N_17310);
nand U17876 (N_17876,N_17460,N_17325);
and U17877 (N_17877,N_17300,N_17130);
and U17878 (N_17878,N_17388,N_17393);
nor U17879 (N_17879,N_17284,N_17007);
or U17880 (N_17880,N_17438,N_17092);
nor U17881 (N_17881,N_17359,N_17095);
xnor U17882 (N_17882,N_17182,N_17097);
and U17883 (N_17883,N_17430,N_17145);
nor U17884 (N_17884,N_17107,N_17382);
or U17885 (N_17885,N_17454,N_17287);
xor U17886 (N_17886,N_17347,N_17170);
and U17887 (N_17887,N_17045,N_17066);
nor U17888 (N_17888,N_17252,N_17370);
or U17889 (N_17889,N_17102,N_17242);
or U17890 (N_17890,N_17409,N_17121);
nor U17891 (N_17891,N_17453,N_17469);
nor U17892 (N_17892,N_17486,N_17463);
nand U17893 (N_17893,N_17423,N_17022);
or U17894 (N_17894,N_17091,N_17084);
nand U17895 (N_17895,N_17105,N_17262);
xnor U17896 (N_17896,N_17220,N_17272);
or U17897 (N_17897,N_17028,N_17293);
or U17898 (N_17898,N_17201,N_17207);
nand U17899 (N_17899,N_17258,N_17066);
xor U17900 (N_17900,N_17337,N_17036);
xor U17901 (N_17901,N_17396,N_17169);
xnor U17902 (N_17902,N_17106,N_17116);
nor U17903 (N_17903,N_17266,N_17302);
or U17904 (N_17904,N_17293,N_17096);
or U17905 (N_17905,N_17102,N_17332);
or U17906 (N_17906,N_17243,N_17083);
nand U17907 (N_17907,N_17157,N_17160);
nor U17908 (N_17908,N_17303,N_17271);
nor U17909 (N_17909,N_17077,N_17458);
nor U17910 (N_17910,N_17126,N_17022);
and U17911 (N_17911,N_17465,N_17098);
xor U17912 (N_17912,N_17075,N_17015);
nor U17913 (N_17913,N_17455,N_17089);
nand U17914 (N_17914,N_17227,N_17089);
xnor U17915 (N_17915,N_17418,N_17087);
xor U17916 (N_17916,N_17313,N_17032);
nor U17917 (N_17917,N_17199,N_17393);
and U17918 (N_17918,N_17323,N_17064);
nor U17919 (N_17919,N_17146,N_17276);
xnor U17920 (N_17920,N_17477,N_17101);
or U17921 (N_17921,N_17327,N_17192);
or U17922 (N_17922,N_17375,N_17255);
xor U17923 (N_17923,N_17382,N_17066);
nand U17924 (N_17924,N_17206,N_17259);
and U17925 (N_17925,N_17334,N_17246);
nor U17926 (N_17926,N_17024,N_17008);
nand U17927 (N_17927,N_17112,N_17394);
nand U17928 (N_17928,N_17343,N_17340);
nand U17929 (N_17929,N_17126,N_17246);
nor U17930 (N_17930,N_17326,N_17367);
and U17931 (N_17931,N_17059,N_17472);
nand U17932 (N_17932,N_17280,N_17048);
and U17933 (N_17933,N_17316,N_17234);
nand U17934 (N_17934,N_17410,N_17259);
and U17935 (N_17935,N_17207,N_17016);
xor U17936 (N_17936,N_17042,N_17025);
and U17937 (N_17937,N_17261,N_17485);
nor U17938 (N_17938,N_17186,N_17411);
xnor U17939 (N_17939,N_17004,N_17034);
nand U17940 (N_17940,N_17318,N_17192);
xnor U17941 (N_17941,N_17430,N_17429);
nor U17942 (N_17942,N_17379,N_17019);
or U17943 (N_17943,N_17206,N_17440);
and U17944 (N_17944,N_17144,N_17294);
nand U17945 (N_17945,N_17309,N_17367);
or U17946 (N_17946,N_17075,N_17130);
nor U17947 (N_17947,N_17000,N_17188);
xor U17948 (N_17948,N_17054,N_17197);
or U17949 (N_17949,N_17314,N_17375);
nand U17950 (N_17950,N_17262,N_17054);
or U17951 (N_17951,N_17004,N_17033);
and U17952 (N_17952,N_17104,N_17236);
and U17953 (N_17953,N_17162,N_17035);
xnor U17954 (N_17954,N_17474,N_17321);
nor U17955 (N_17955,N_17150,N_17426);
nand U17956 (N_17956,N_17117,N_17252);
nor U17957 (N_17957,N_17239,N_17035);
xor U17958 (N_17958,N_17268,N_17145);
or U17959 (N_17959,N_17226,N_17188);
and U17960 (N_17960,N_17130,N_17054);
nor U17961 (N_17961,N_17285,N_17040);
nand U17962 (N_17962,N_17292,N_17148);
xor U17963 (N_17963,N_17066,N_17475);
nor U17964 (N_17964,N_17478,N_17307);
xor U17965 (N_17965,N_17266,N_17113);
or U17966 (N_17966,N_17398,N_17236);
and U17967 (N_17967,N_17292,N_17355);
nor U17968 (N_17968,N_17008,N_17440);
xor U17969 (N_17969,N_17199,N_17030);
or U17970 (N_17970,N_17248,N_17165);
nand U17971 (N_17971,N_17310,N_17232);
xor U17972 (N_17972,N_17236,N_17329);
or U17973 (N_17973,N_17060,N_17343);
nor U17974 (N_17974,N_17193,N_17415);
and U17975 (N_17975,N_17365,N_17336);
or U17976 (N_17976,N_17064,N_17412);
or U17977 (N_17977,N_17266,N_17188);
nor U17978 (N_17978,N_17309,N_17137);
nand U17979 (N_17979,N_17432,N_17152);
nand U17980 (N_17980,N_17470,N_17346);
nand U17981 (N_17981,N_17275,N_17113);
and U17982 (N_17982,N_17046,N_17396);
or U17983 (N_17983,N_17106,N_17386);
nor U17984 (N_17984,N_17350,N_17425);
or U17985 (N_17985,N_17056,N_17470);
nand U17986 (N_17986,N_17100,N_17478);
nand U17987 (N_17987,N_17222,N_17343);
or U17988 (N_17988,N_17270,N_17259);
nand U17989 (N_17989,N_17069,N_17368);
and U17990 (N_17990,N_17261,N_17187);
nor U17991 (N_17991,N_17419,N_17206);
or U17992 (N_17992,N_17172,N_17383);
nand U17993 (N_17993,N_17263,N_17223);
xor U17994 (N_17994,N_17475,N_17136);
xnor U17995 (N_17995,N_17103,N_17441);
and U17996 (N_17996,N_17427,N_17070);
nand U17997 (N_17997,N_17019,N_17252);
or U17998 (N_17998,N_17357,N_17438);
and U17999 (N_17999,N_17388,N_17168);
nand U18000 (N_18000,N_17597,N_17853);
nor U18001 (N_18001,N_17596,N_17518);
and U18002 (N_18002,N_17774,N_17550);
and U18003 (N_18003,N_17538,N_17714);
or U18004 (N_18004,N_17587,N_17789);
xor U18005 (N_18005,N_17666,N_17971);
xor U18006 (N_18006,N_17546,N_17558);
nor U18007 (N_18007,N_17740,N_17870);
xor U18008 (N_18008,N_17645,N_17904);
and U18009 (N_18009,N_17808,N_17547);
or U18010 (N_18010,N_17926,N_17748);
nor U18011 (N_18011,N_17905,N_17728);
nand U18012 (N_18012,N_17986,N_17946);
xnor U18013 (N_18013,N_17694,N_17802);
nand U18014 (N_18014,N_17651,N_17586);
nand U18015 (N_18015,N_17729,N_17626);
nor U18016 (N_18016,N_17648,N_17697);
and U18017 (N_18017,N_17901,N_17701);
nor U18018 (N_18018,N_17842,N_17511);
xnor U18019 (N_18019,N_17762,N_17973);
and U18020 (N_18020,N_17929,N_17617);
nand U18021 (N_18021,N_17799,N_17878);
nand U18022 (N_18022,N_17744,N_17852);
xor U18023 (N_18023,N_17532,N_17997);
nor U18024 (N_18024,N_17541,N_17578);
and U18025 (N_18025,N_17646,N_17838);
or U18026 (N_18026,N_17724,N_17994);
nand U18027 (N_18027,N_17938,N_17579);
or U18028 (N_18028,N_17529,N_17640);
xnor U18029 (N_18029,N_17784,N_17979);
nor U18030 (N_18030,N_17663,N_17805);
xnor U18031 (N_18031,N_17862,N_17741);
or U18032 (N_18032,N_17897,N_17711);
nand U18033 (N_18033,N_17869,N_17871);
nor U18034 (N_18034,N_17603,N_17957);
nand U18035 (N_18035,N_17860,N_17567);
nor U18036 (N_18036,N_17618,N_17730);
and U18037 (N_18037,N_17914,N_17857);
xor U18038 (N_18038,N_17809,N_17900);
or U18039 (N_18039,N_17710,N_17670);
nand U18040 (N_18040,N_17516,N_17721);
or U18041 (N_18041,N_17936,N_17912);
nand U18042 (N_18042,N_17874,N_17580);
or U18043 (N_18043,N_17656,N_17713);
xor U18044 (N_18044,N_17557,N_17828);
xor U18045 (N_18045,N_17850,N_17998);
nor U18046 (N_18046,N_17611,N_17826);
and U18047 (N_18047,N_17898,N_17715);
xor U18048 (N_18048,N_17562,N_17664);
xnor U18049 (N_18049,N_17556,N_17595);
nand U18050 (N_18050,N_17833,N_17680);
or U18051 (N_18051,N_17781,N_17782);
nand U18052 (N_18052,N_17847,N_17954);
and U18053 (N_18053,N_17768,N_17693);
xnor U18054 (N_18054,N_17976,N_17636);
nor U18055 (N_18055,N_17948,N_17739);
xor U18056 (N_18056,N_17980,N_17778);
nand U18057 (N_18057,N_17812,N_17820);
or U18058 (N_18058,N_17819,N_17633);
and U18059 (N_18059,N_17968,N_17872);
and U18060 (N_18060,N_17987,N_17671);
nand U18061 (N_18061,N_17644,N_17771);
nor U18062 (N_18062,N_17615,N_17628);
xnor U18063 (N_18063,N_17890,N_17930);
nand U18064 (N_18064,N_17554,N_17803);
nand U18065 (N_18065,N_17876,N_17982);
or U18066 (N_18066,N_17649,N_17502);
xor U18067 (N_18067,N_17524,N_17577);
and U18068 (N_18068,N_17821,N_17638);
nor U18069 (N_18069,N_17773,N_17612);
or U18070 (N_18070,N_17574,N_17704);
or U18071 (N_18071,N_17955,N_17951);
or U18072 (N_18072,N_17725,N_17756);
and U18073 (N_18073,N_17661,N_17927);
nand U18074 (N_18074,N_17760,N_17848);
nand U18075 (N_18075,N_17689,N_17829);
or U18076 (N_18076,N_17944,N_17747);
or U18077 (N_18077,N_17967,N_17952);
xor U18078 (N_18078,N_17960,N_17563);
or U18079 (N_18079,N_17984,N_17537);
nor U18080 (N_18080,N_17703,N_17632);
and U18081 (N_18081,N_17947,N_17528);
nand U18082 (N_18082,N_17736,N_17877);
nand U18083 (N_18083,N_17561,N_17508);
nand U18084 (N_18084,N_17500,N_17896);
nor U18085 (N_18085,N_17983,N_17705);
xor U18086 (N_18086,N_17919,N_17962);
nand U18087 (N_18087,N_17893,N_17950);
xor U18088 (N_18088,N_17514,N_17504);
and U18089 (N_18089,N_17868,N_17683);
or U18090 (N_18090,N_17551,N_17684);
xor U18091 (N_18091,N_17902,N_17681);
xnor U18092 (N_18092,N_17840,N_17765);
xnor U18093 (N_18093,N_17759,N_17629);
xnor U18094 (N_18094,N_17658,N_17506);
and U18095 (N_18095,N_17916,N_17698);
or U18096 (N_18096,N_17583,N_17770);
xnor U18097 (N_18097,N_17501,N_17515);
nand U18098 (N_18098,N_17772,N_17956);
and U18099 (N_18099,N_17750,N_17702);
or U18100 (N_18100,N_17953,N_17575);
or U18101 (N_18101,N_17513,N_17841);
and U18102 (N_18102,N_17972,N_17882);
nor U18103 (N_18103,N_17534,N_17751);
xor U18104 (N_18104,N_17667,N_17717);
nor U18105 (N_18105,N_17610,N_17593);
and U18106 (N_18106,N_17922,N_17552);
and U18107 (N_18107,N_17837,N_17881);
or U18108 (N_18108,N_17723,N_17627);
nand U18109 (N_18109,N_17525,N_17544);
nor U18110 (N_18110,N_17619,N_17609);
nand U18111 (N_18111,N_17969,N_17700);
nand U18112 (N_18112,N_17676,N_17920);
nor U18113 (N_18113,N_17915,N_17637);
nand U18114 (N_18114,N_17565,N_17572);
nor U18115 (N_18115,N_17776,N_17908);
xor U18116 (N_18116,N_17801,N_17855);
xnor U18117 (N_18117,N_17849,N_17737);
nor U18118 (N_18118,N_17581,N_17709);
nor U18119 (N_18119,N_17788,N_17790);
nand U18120 (N_18120,N_17553,N_17527);
or U18121 (N_18121,N_17815,N_17607);
and U18122 (N_18122,N_17811,N_17845);
xnor U18123 (N_18123,N_17669,N_17906);
nor U18124 (N_18124,N_17526,N_17793);
or U18125 (N_18125,N_17941,N_17641);
nor U18126 (N_18126,N_17732,N_17530);
or U18127 (N_18127,N_17932,N_17797);
xor U18128 (N_18128,N_17978,N_17832);
and U18129 (N_18129,N_17854,N_17995);
or U18130 (N_18130,N_17807,N_17923);
or U18131 (N_18131,N_17659,N_17660);
and U18132 (N_18132,N_17974,N_17889);
xor U18133 (N_18133,N_17549,N_17894);
nand U18134 (N_18134,N_17509,N_17623);
nand U18135 (N_18135,N_17682,N_17767);
nor U18136 (N_18136,N_17754,N_17522);
or U18137 (N_18137,N_17712,N_17576);
xor U18138 (N_18138,N_17743,N_17591);
and U18139 (N_18139,N_17911,N_17753);
or U18140 (N_18140,N_17865,N_17935);
and U18141 (N_18141,N_17794,N_17787);
xnor U18142 (N_18142,N_17888,N_17699);
or U18143 (N_18143,N_17589,N_17718);
or U18144 (N_18144,N_17824,N_17695);
and U18145 (N_18145,N_17825,N_17545);
or U18146 (N_18146,N_17909,N_17517);
xor U18147 (N_18147,N_17687,N_17861);
and U18148 (N_18148,N_17616,N_17566);
or U18149 (N_18149,N_17599,N_17662);
nand U18150 (N_18150,N_17726,N_17839);
and U18151 (N_18151,N_17925,N_17884);
nand U18152 (N_18152,N_17672,N_17937);
and U18153 (N_18153,N_17548,N_17866);
nor U18154 (N_18154,N_17813,N_17654);
nor U18155 (N_18155,N_17961,N_17688);
nand U18156 (N_18156,N_17569,N_17691);
nand U18157 (N_18157,N_17505,N_17903);
nand U18158 (N_18158,N_17798,N_17592);
xor U18159 (N_18159,N_17988,N_17720);
and U18160 (N_18160,N_17796,N_17823);
or U18161 (N_18161,N_17622,N_17598);
nor U18162 (N_18162,N_17677,N_17523);
and U18163 (N_18163,N_17542,N_17605);
nand U18164 (N_18164,N_17958,N_17634);
nor U18165 (N_18165,N_17835,N_17560);
or U18166 (N_18166,N_17875,N_17873);
nor U18167 (N_18167,N_17650,N_17647);
xor U18168 (N_18168,N_17945,N_17746);
nand U18169 (N_18169,N_17891,N_17928);
nand U18170 (N_18170,N_17999,N_17559);
xnor U18171 (N_18171,N_17921,N_17943);
and U18172 (N_18172,N_17910,N_17512);
nor U18173 (N_18173,N_17630,N_17734);
and U18174 (N_18174,N_17727,N_17814);
nand U18175 (N_18175,N_17886,N_17692);
nand U18176 (N_18176,N_17604,N_17758);
nand U18177 (N_18177,N_17613,N_17779);
xnor U18178 (N_18178,N_17844,N_17696);
xor U18179 (N_18179,N_17863,N_17883);
nand U18180 (N_18180,N_17993,N_17752);
xnor U18181 (N_18181,N_17570,N_17675);
xnor U18182 (N_18182,N_17975,N_17585);
and U18183 (N_18183,N_17964,N_17678);
or U18184 (N_18184,N_17851,N_17965);
xnor U18185 (N_18185,N_17846,N_17867);
xor U18186 (N_18186,N_17786,N_17989);
or U18187 (N_18187,N_17708,N_17738);
nand U18188 (N_18188,N_17584,N_17843);
and U18189 (N_18189,N_17918,N_17764);
xor U18190 (N_18190,N_17913,N_17977);
or U18191 (N_18191,N_17543,N_17970);
or U18192 (N_18192,N_17836,N_17831);
nor U18193 (N_18193,N_17981,N_17933);
nand U18194 (N_18194,N_17571,N_17766);
xnor U18195 (N_18195,N_17657,N_17521);
nor U18196 (N_18196,N_17745,N_17742);
or U18197 (N_18197,N_17939,N_17707);
nand U18198 (N_18198,N_17880,N_17635);
xor U18199 (N_18199,N_17749,N_17555);
xnor U18200 (N_18200,N_17755,N_17931);
nand U18201 (N_18201,N_17674,N_17540);
nor U18202 (N_18202,N_17519,N_17777);
nand U18203 (N_18203,N_17887,N_17639);
and U18204 (N_18204,N_17539,N_17963);
xnor U18205 (N_18205,N_17792,N_17827);
nor U18206 (N_18206,N_17722,N_17594);
or U18207 (N_18207,N_17966,N_17690);
and U18208 (N_18208,N_17783,N_17934);
and U18209 (N_18209,N_17520,N_17685);
and U18210 (N_18210,N_17568,N_17631);
and U18211 (N_18211,N_17735,N_17818);
and U18212 (N_18212,N_17625,N_17757);
nand U18213 (N_18213,N_17806,N_17573);
xnor U18214 (N_18214,N_17991,N_17533);
xor U18215 (N_18215,N_17856,N_17942);
nand U18216 (N_18216,N_17892,N_17621);
nand U18217 (N_18217,N_17769,N_17924);
nor U18218 (N_18218,N_17719,N_17785);
nand U18219 (N_18219,N_17907,N_17822);
or U18220 (N_18220,N_17795,N_17679);
or U18221 (N_18221,N_17655,N_17601);
xor U18222 (N_18222,N_17564,N_17940);
nand U18223 (N_18223,N_17668,N_17864);
and U18224 (N_18224,N_17885,N_17996);
nor U18225 (N_18225,N_17643,N_17642);
or U18226 (N_18226,N_17531,N_17665);
or U18227 (N_18227,N_17582,N_17590);
and U18228 (N_18228,N_17899,N_17949);
nand U18229 (N_18229,N_17830,N_17810);
nor U18230 (N_18230,N_17673,N_17653);
nand U18231 (N_18231,N_17606,N_17895);
nor U18232 (N_18232,N_17763,N_17775);
nand U18233 (N_18233,N_17858,N_17614);
or U18234 (N_18234,N_17507,N_17834);
and U18235 (N_18235,N_17817,N_17990);
nor U18236 (N_18236,N_17608,N_17686);
and U18237 (N_18237,N_17652,N_17992);
and U18238 (N_18238,N_17791,N_17624);
xnor U18239 (N_18239,N_17859,N_17716);
or U18240 (N_18240,N_17588,N_17535);
or U18241 (N_18241,N_17761,N_17731);
nand U18242 (N_18242,N_17602,N_17733);
or U18243 (N_18243,N_17510,N_17917);
or U18244 (N_18244,N_17503,N_17800);
nor U18245 (N_18245,N_17536,N_17780);
nand U18246 (N_18246,N_17816,N_17600);
nor U18247 (N_18247,N_17804,N_17959);
xor U18248 (N_18248,N_17620,N_17985);
and U18249 (N_18249,N_17879,N_17706);
nor U18250 (N_18250,N_17509,N_17555);
nor U18251 (N_18251,N_17694,N_17614);
or U18252 (N_18252,N_17945,N_17970);
nor U18253 (N_18253,N_17640,N_17749);
and U18254 (N_18254,N_17586,N_17941);
nand U18255 (N_18255,N_17699,N_17939);
and U18256 (N_18256,N_17592,N_17570);
nand U18257 (N_18257,N_17871,N_17690);
nand U18258 (N_18258,N_17571,N_17746);
nand U18259 (N_18259,N_17728,N_17570);
xor U18260 (N_18260,N_17963,N_17721);
or U18261 (N_18261,N_17999,N_17739);
and U18262 (N_18262,N_17644,N_17580);
and U18263 (N_18263,N_17656,N_17526);
nor U18264 (N_18264,N_17946,N_17745);
nor U18265 (N_18265,N_17866,N_17565);
or U18266 (N_18266,N_17558,N_17929);
or U18267 (N_18267,N_17758,N_17776);
nor U18268 (N_18268,N_17834,N_17592);
or U18269 (N_18269,N_17834,N_17685);
or U18270 (N_18270,N_17674,N_17987);
or U18271 (N_18271,N_17853,N_17961);
or U18272 (N_18272,N_17531,N_17830);
xnor U18273 (N_18273,N_17590,N_17850);
or U18274 (N_18274,N_17643,N_17531);
xnor U18275 (N_18275,N_17645,N_17750);
nand U18276 (N_18276,N_17730,N_17777);
xor U18277 (N_18277,N_17955,N_17654);
or U18278 (N_18278,N_17580,N_17757);
and U18279 (N_18279,N_17945,N_17928);
nor U18280 (N_18280,N_17657,N_17743);
or U18281 (N_18281,N_17786,N_17681);
and U18282 (N_18282,N_17795,N_17732);
xor U18283 (N_18283,N_17742,N_17975);
or U18284 (N_18284,N_17607,N_17526);
or U18285 (N_18285,N_17596,N_17988);
and U18286 (N_18286,N_17666,N_17669);
or U18287 (N_18287,N_17901,N_17780);
xnor U18288 (N_18288,N_17812,N_17526);
nor U18289 (N_18289,N_17969,N_17987);
or U18290 (N_18290,N_17658,N_17883);
nor U18291 (N_18291,N_17682,N_17652);
and U18292 (N_18292,N_17526,N_17701);
and U18293 (N_18293,N_17591,N_17896);
xor U18294 (N_18294,N_17612,N_17794);
and U18295 (N_18295,N_17738,N_17881);
nand U18296 (N_18296,N_17756,N_17820);
xor U18297 (N_18297,N_17749,N_17772);
nor U18298 (N_18298,N_17568,N_17989);
and U18299 (N_18299,N_17728,N_17819);
and U18300 (N_18300,N_17609,N_17694);
nor U18301 (N_18301,N_17789,N_17788);
xor U18302 (N_18302,N_17726,N_17722);
and U18303 (N_18303,N_17987,N_17822);
xor U18304 (N_18304,N_17907,N_17522);
nand U18305 (N_18305,N_17518,N_17762);
nand U18306 (N_18306,N_17649,N_17553);
nor U18307 (N_18307,N_17606,N_17561);
xor U18308 (N_18308,N_17681,N_17944);
and U18309 (N_18309,N_17782,N_17814);
xnor U18310 (N_18310,N_17784,N_17894);
nor U18311 (N_18311,N_17903,N_17933);
xor U18312 (N_18312,N_17998,N_17768);
nand U18313 (N_18313,N_17704,N_17715);
xor U18314 (N_18314,N_17553,N_17520);
nor U18315 (N_18315,N_17571,N_17805);
nand U18316 (N_18316,N_17518,N_17737);
nand U18317 (N_18317,N_17998,N_17814);
xnor U18318 (N_18318,N_17629,N_17787);
nor U18319 (N_18319,N_17880,N_17940);
xor U18320 (N_18320,N_17646,N_17854);
xnor U18321 (N_18321,N_17925,N_17518);
nand U18322 (N_18322,N_17607,N_17840);
xor U18323 (N_18323,N_17656,N_17834);
nand U18324 (N_18324,N_17959,N_17692);
nor U18325 (N_18325,N_17770,N_17970);
nand U18326 (N_18326,N_17840,N_17550);
or U18327 (N_18327,N_17608,N_17800);
nand U18328 (N_18328,N_17780,N_17841);
or U18329 (N_18329,N_17576,N_17709);
nand U18330 (N_18330,N_17976,N_17660);
xnor U18331 (N_18331,N_17831,N_17964);
and U18332 (N_18332,N_17868,N_17822);
or U18333 (N_18333,N_17575,N_17932);
nor U18334 (N_18334,N_17687,N_17997);
nand U18335 (N_18335,N_17904,N_17680);
or U18336 (N_18336,N_17634,N_17540);
xor U18337 (N_18337,N_17726,N_17585);
nor U18338 (N_18338,N_17693,N_17988);
and U18339 (N_18339,N_17730,N_17830);
and U18340 (N_18340,N_17847,N_17734);
nor U18341 (N_18341,N_17945,N_17583);
or U18342 (N_18342,N_17595,N_17708);
or U18343 (N_18343,N_17640,N_17926);
xnor U18344 (N_18344,N_17648,N_17934);
xor U18345 (N_18345,N_17898,N_17758);
nand U18346 (N_18346,N_17575,N_17781);
xor U18347 (N_18347,N_17721,N_17694);
and U18348 (N_18348,N_17544,N_17518);
or U18349 (N_18349,N_17556,N_17621);
nand U18350 (N_18350,N_17553,N_17849);
or U18351 (N_18351,N_17637,N_17741);
xnor U18352 (N_18352,N_17712,N_17730);
or U18353 (N_18353,N_17575,N_17592);
nor U18354 (N_18354,N_17794,N_17951);
and U18355 (N_18355,N_17742,N_17651);
or U18356 (N_18356,N_17916,N_17808);
and U18357 (N_18357,N_17772,N_17606);
nand U18358 (N_18358,N_17753,N_17735);
nor U18359 (N_18359,N_17787,N_17534);
nand U18360 (N_18360,N_17944,N_17728);
nor U18361 (N_18361,N_17784,N_17883);
nor U18362 (N_18362,N_17709,N_17858);
nand U18363 (N_18363,N_17567,N_17749);
or U18364 (N_18364,N_17937,N_17998);
xor U18365 (N_18365,N_17929,N_17614);
nand U18366 (N_18366,N_17957,N_17513);
and U18367 (N_18367,N_17584,N_17648);
or U18368 (N_18368,N_17785,N_17821);
xnor U18369 (N_18369,N_17709,N_17904);
and U18370 (N_18370,N_17686,N_17566);
and U18371 (N_18371,N_17962,N_17993);
nor U18372 (N_18372,N_17580,N_17514);
nand U18373 (N_18373,N_17551,N_17988);
nand U18374 (N_18374,N_17964,N_17648);
or U18375 (N_18375,N_17633,N_17719);
xnor U18376 (N_18376,N_17700,N_17919);
nor U18377 (N_18377,N_17703,N_17579);
or U18378 (N_18378,N_17962,N_17527);
xor U18379 (N_18379,N_17921,N_17717);
xor U18380 (N_18380,N_17697,N_17936);
and U18381 (N_18381,N_17736,N_17708);
or U18382 (N_18382,N_17775,N_17693);
and U18383 (N_18383,N_17725,N_17629);
nor U18384 (N_18384,N_17909,N_17723);
xor U18385 (N_18385,N_17502,N_17592);
nand U18386 (N_18386,N_17712,N_17802);
nand U18387 (N_18387,N_17877,N_17797);
xnor U18388 (N_18388,N_17506,N_17601);
nor U18389 (N_18389,N_17678,N_17958);
or U18390 (N_18390,N_17935,N_17897);
or U18391 (N_18391,N_17890,N_17611);
and U18392 (N_18392,N_17583,N_17899);
nor U18393 (N_18393,N_17951,N_17969);
nand U18394 (N_18394,N_17546,N_17579);
xnor U18395 (N_18395,N_17805,N_17906);
xor U18396 (N_18396,N_17623,N_17833);
xor U18397 (N_18397,N_17947,N_17517);
or U18398 (N_18398,N_17987,N_17594);
nor U18399 (N_18399,N_17812,N_17642);
xor U18400 (N_18400,N_17636,N_17737);
nand U18401 (N_18401,N_17517,N_17596);
or U18402 (N_18402,N_17703,N_17944);
and U18403 (N_18403,N_17540,N_17556);
or U18404 (N_18404,N_17600,N_17640);
xor U18405 (N_18405,N_17744,N_17654);
or U18406 (N_18406,N_17748,N_17741);
xnor U18407 (N_18407,N_17549,N_17693);
nand U18408 (N_18408,N_17762,N_17645);
nand U18409 (N_18409,N_17947,N_17712);
nor U18410 (N_18410,N_17535,N_17540);
nand U18411 (N_18411,N_17806,N_17943);
nand U18412 (N_18412,N_17540,N_17790);
and U18413 (N_18413,N_17617,N_17765);
nand U18414 (N_18414,N_17779,N_17791);
nor U18415 (N_18415,N_17694,N_17985);
nand U18416 (N_18416,N_17702,N_17953);
or U18417 (N_18417,N_17826,N_17751);
xnor U18418 (N_18418,N_17651,N_17605);
nor U18419 (N_18419,N_17658,N_17535);
xnor U18420 (N_18420,N_17552,N_17604);
or U18421 (N_18421,N_17950,N_17867);
xor U18422 (N_18422,N_17706,N_17692);
xor U18423 (N_18423,N_17661,N_17766);
and U18424 (N_18424,N_17919,N_17994);
nor U18425 (N_18425,N_17810,N_17770);
or U18426 (N_18426,N_17750,N_17912);
nand U18427 (N_18427,N_17574,N_17910);
nor U18428 (N_18428,N_17837,N_17551);
nand U18429 (N_18429,N_17818,N_17516);
or U18430 (N_18430,N_17810,N_17938);
and U18431 (N_18431,N_17965,N_17946);
xnor U18432 (N_18432,N_17892,N_17673);
and U18433 (N_18433,N_17691,N_17543);
xor U18434 (N_18434,N_17701,N_17863);
and U18435 (N_18435,N_17933,N_17555);
or U18436 (N_18436,N_17676,N_17922);
and U18437 (N_18437,N_17908,N_17875);
nand U18438 (N_18438,N_17931,N_17989);
or U18439 (N_18439,N_17508,N_17620);
xor U18440 (N_18440,N_17534,N_17606);
and U18441 (N_18441,N_17697,N_17927);
or U18442 (N_18442,N_17837,N_17960);
xor U18443 (N_18443,N_17642,N_17510);
nor U18444 (N_18444,N_17984,N_17951);
and U18445 (N_18445,N_17976,N_17643);
nand U18446 (N_18446,N_17501,N_17584);
xor U18447 (N_18447,N_17823,N_17555);
or U18448 (N_18448,N_17507,N_17616);
and U18449 (N_18449,N_17874,N_17757);
nand U18450 (N_18450,N_17843,N_17935);
nor U18451 (N_18451,N_17768,N_17996);
and U18452 (N_18452,N_17702,N_17837);
nand U18453 (N_18453,N_17980,N_17659);
and U18454 (N_18454,N_17988,N_17914);
nor U18455 (N_18455,N_17959,N_17689);
and U18456 (N_18456,N_17608,N_17544);
xor U18457 (N_18457,N_17815,N_17945);
nor U18458 (N_18458,N_17966,N_17981);
nor U18459 (N_18459,N_17693,N_17855);
or U18460 (N_18460,N_17862,N_17825);
nand U18461 (N_18461,N_17922,N_17512);
or U18462 (N_18462,N_17516,N_17820);
and U18463 (N_18463,N_17693,N_17965);
and U18464 (N_18464,N_17645,N_17686);
nor U18465 (N_18465,N_17662,N_17634);
nand U18466 (N_18466,N_17742,N_17955);
nand U18467 (N_18467,N_17596,N_17592);
and U18468 (N_18468,N_17516,N_17876);
nand U18469 (N_18469,N_17951,N_17985);
or U18470 (N_18470,N_17833,N_17639);
xnor U18471 (N_18471,N_17963,N_17642);
xnor U18472 (N_18472,N_17938,N_17855);
nor U18473 (N_18473,N_17881,N_17507);
nor U18474 (N_18474,N_17904,N_17591);
nand U18475 (N_18475,N_17960,N_17540);
xnor U18476 (N_18476,N_17854,N_17754);
nand U18477 (N_18477,N_17955,N_17504);
xnor U18478 (N_18478,N_17653,N_17820);
xnor U18479 (N_18479,N_17826,N_17518);
or U18480 (N_18480,N_17931,N_17992);
or U18481 (N_18481,N_17898,N_17668);
or U18482 (N_18482,N_17708,N_17661);
and U18483 (N_18483,N_17858,N_17891);
or U18484 (N_18484,N_17748,N_17625);
nor U18485 (N_18485,N_17578,N_17694);
nand U18486 (N_18486,N_17505,N_17750);
xnor U18487 (N_18487,N_17530,N_17587);
xor U18488 (N_18488,N_17849,N_17546);
xor U18489 (N_18489,N_17875,N_17952);
or U18490 (N_18490,N_17543,N_17633);
xor U18491 (N_18491,N_17541,N_17863);
nor U18492 (N_18492,N_17778,N_17632);
or U18493 (N_18493,N_17753,N_17558);
or U18494 (N_18494,N_17568,N_17681);
or U18495 (N_18495,N_17765,N_17708);
and U18496 (N_18496,N_17801,N_17637);
nor U18497 (N_18497,N_17907,N_17585);
nand U18498 (N_18498,N_17636,N_17867);
nor U18499 (N_18499,N_17846,N_17647);
nor U18500 (N_18500,N_18081,N_18391);
nor U18501 (N_18501,N_18035,N_18366);
xor U18502 (N_18502,N_18483,N_18087);
xor U18503 (N_18503,N_18061,N_18362);
nor U18504 (N_18504,N_18312,N_18481);
xnor U18505 (N_18505,N_18418,N_18268);
xor U18506 (N_18506,N_18271,N_18135);
and U18507 (N_18507,N_18376,N_18461);
nand U18508 (N_18508,N_18170,N_18046);
xnor U18509 (N_18509,N_18319,N_18279);
nand U18510 (N_18510,N_18371,N_18244);
nand U18511 (N_18511,N_18079,N_18356);
nand U18512 (N_18512,N_18198,N_18097);
and U18513 (N_18513,N_18113,N_18395);
xor U18514 (N_18514,N_18055,N_18430);
xnor U18515 (N_18515,N_18092,N_18377);
and U18516 (N_18516,N_18153,N_18161);
or U18517 (N_18517,N_18260,N_18400);
xnor U18518 (N_18518,N_18223,N_18259);
nand U18519 (N_18519,N_18293,N_18382);
xnor U18520 (N_18520,N_18007,N_18424);
or U18521 (N_18521,N_18297,N_18242);
and U18522 (N_18522,N_18166,N_18266);
or U18523 (N_18523,N_18108,N_18020);
or U18524 (N_18524,N_18155,N_18291);
and U18525 (N_18525,N_18167,N_18299);
xnor U18526 (N_18526,N_18445,N_18329);
nand U18527 (N_18527,N_18157,N_18335);
nand U18528 (N_18528,N_18407,N_18453);
and U18529 (N_18529,N_18273,N_18317);
xor U18530 (N_18530,N_18488,N_18475);
xor U18531 (N_18531,N_18011,N_18287);
or U18532 (N_18532,N_18158,N_18363);
nand U18533 (N_18533,N_18015,N_18443);
or U18534 (N_18534,N_18422,N_18197);
and U18535 (N_18535,N_18368,N_18338);
nor U18536 (N_18536,N_18429,N_18220);
xnor U18537 (N_18537,N_18148,N_18369);
nor U18538 (N_18538,N_18272,N_18406);
nand U18539 (N_18539,N_18386,N_18474);
xnor U18540 (N_18540,N_18387,N_18129);
and U18541 (N_18541,N_18265,N_18094);
and U18542 (N_18542,N_18428,N_18193);
and U18543 (N_18543,N_18328,N_18385);
and U18544 (N_18544,N_18064,N_18245);
nand U18545 (N_18545,N_18458,N_18044);
nor U18546 (N_18546,N_18337,N_18436);
nand U18547 (N_18547,N_18334,N_18002);
and U18548 (N_18548,N_18082,N_18039);
or U18549 (N_18549,N_18303,N_18004);
nor U18550 (N_18550,N_18173,N_18309);
xnor U18551 (N_18551,N_18137,N_18147);
and U18552 (N_18552,N_18016,N_18225);
xnor U18553 (N_18553,N_18058,N_18486);
or U18554 (N_18554,N_18304,N_18402);
nor U18555 (N_18555,N_18459,N_18254);
and U18556 (N_18556,N_18238,N_18141);
or U18557 (N_18557,N_18447,N_18469);
or U18558 (N_18558,N_18205,N_18188);
nand U18559 (N_18559,N_18175,N_18003);
nor U18560 (N_18560,N_18359,N_18460);
and U18561 (N_18561,N_18066,N_18036);
xnor U18562 (N_18562,N_18209,N_18345);
nor U18563 (N_18563,N_18292,N_18256);
xor U18564 (N_18564,N_18091,N_18103);
and U18565 (N_18565,N_18229,N_18285);
xor U18566 (N_18566,N_18326,N_18399);
and U18567 (N_18567,N_18029,N_18479);
or U18568 (N_18568,N_18107,N_18180);
xnor U18569 (N_18569,N_18380,N_18408);
xor U18570 (N_18570,N_18189,N_18218);
nand U18571 (N_18571,N_18243,N_18057);
xnor U18572 (N_18572,N_18276,N_18080);
or U18573 (N_18573,N_18423,N_18361);
nand U18574 (N_18574,N_18125,N_18085);
or U18575 (N_18575,N_18263,N_18116);
and U18576 (N_18576,N_18446,N_18373);
or U18577 (N_18577,N_18143,N_18330);
or U18578 (N_18578,N_18000,N_18405);
and U18579 (N_18579,N_18093,N_18340);
and U18580 (N_18580,N_18019,N_18195);
nand U18581 (N_18581,N_18232,N_18301);
or U18582 (N_18582,N_18347,N_18327);
or U18583 (N_18583,N_18182,N_18201);
xnor U18584 (N_18584,N_18110,N_18247);
and U18585 (N_18585,N_18040,N_18230);
xor U18586 (N_18586,N_18455,N_18496);
nor U18587 (N_18587,N_18012,N_18117);
nand U18588 (N_18588,N_18096,N_18250);
xnor U18589 (N_18589,N_18315,N_18289);
or U18590 (N_18590,N_18439,N_18420);
xnor U18591 (N_18591,N_18352,N_18492);
and U18592 (N_18592,N_18191,N_18257);
and U18593 (N_18593,N_18465,N_18401);
or U18594 (N_18594,N_18476,N_18121);
nor U18595 (N_18595,N_18025,N_18417);
nand U18596 (N_18596,N_18199,N_18313);
xnor U18597 (N_18597,N_18028,N_18030);
xnor U18598 (N_18598,N_18236,N_18346);
or U18599 (N_18599,N_18126,N_18069);
nor U18600 (N_18600,N_18294,N_18183);
and U18601 (N_18601,N_18466,N_18332);
or U18602 (N_18602,N_18295,N_18296);
nor U18603 (N_18603,N_18374,N_18045);
and U18604 (N_18604,N_18211,N_18302);
xnor U18605 (N_18605,N_18421,N_18043);
nand U18606 (N_18606,N_18151,N_18450);
nand U18607 (N_18607,N_18398,N_18033);
and U18608 (N_18608,N_18397,N_18112);
nand U18609 (N_18609,N_18214,N_18270);
or U18610 (N_18610,N_18084,N_18095);
nand U18611 (N_18611,N_18278,N_18413);
and U18612 (N_18612,N_18318,N_18073);
nor U18613 (N_18613,N_18231,N_18163);
nor U18614 (N_18614,N_18431,N_18308);
and U18615 (N_18615,N_18001,N_18288);
nor U18616 (N_18616,N_18145,N_18306);
and U18617 (N_18617,N_18241,N_18215);
and U18618 (N_18618,N_18324,N_18381);
or U18619 (N_18619,N_18495,N_18343);
xnor U18620 (N_18620,N_18307,N_18115);
xnor U18621 (N_18621,N_18282,N_18017);
and U18622 (N_18622,N_18300,N_18111);
nand U18623 (N_18623,N_18222,N_18493);
nand U18624 (N_18624,N_18485,N_18419);
and U18625 (N_18625,N_18454,N_18109);
nand U18626 (N_18626,N_18412,N_18342);
xor U18627 (N_18627,N_18379,N_18440);
xor U18628 (N_18628,N_18264,N_18005);
nor U18629 (N_18629,N_18133,N_18498);
nor U18630 (N_18630,N_18206,N_18470);
or U18631 (N_18631,N_18203,N_18261);
xor U18632 (N_18632,N_18118,N_18280);
nor U18633 (N_18633,N_18100,N_18383);
or U18634 (N_18634,N_18070,N_18037);
and U18635 (N_18635,N_18228,N_18441);
or U18636 (N_18636,N_18438,N_18298);
nand U18637 (N_18637,N_18403,N_18196);
nor U18638 (N_18638,N_18089,N_18353);
or U18639 (N_18639,N_18048,N_18122);
xor U18640 (N_18640,N_18047,N_18204);
or U18641 (N_18641,N_18160,N_18022);
or U18642 (N_18642,N_18171,N_18451);
and U18643 (N_18643,N_18212,N_18442);
xnor U18644 (N_18644,N_18491,N_18184);
or U18645 (N_18645,N_18349,N_18364);
xnor U18646 (N_18646,N_18494,N_18456);
nor U18647 (N_18647,N_18393,N_18384);
nor U18648 (N_18648,N_18165,N_18357);
and U18649 (N_18649,N_18034,N_18310);
xor U18650 (N_18650,N_18258,N_18388);
nand U18651 (N_18651,N_18192,N_18119);
nor U18652 (N_18652,N_18339,N_18065);
and U18653 (N_18653,N_18038,N_18255);
or U18654 (N_18654,N_18372,N_18344);
nor U18655 (N_18655,N_18426,N_18086);
nor U18656 (N_18656,N_18168,N_18176);
nand U18657 (N_18657,N_18252,N_18389);
xnor U18658 (N_18658,N_18159,N_18414);
and U18659 (N_18659,N_18060,N_18360);
nand U18660 (N_18660,N_18367,N_18009);
xor U18661 (N_18661,N_18144,N_18437);
nand U18662 (N_18662,N_18051,N_18178);
nor U18663 (N_18663,N_18311,N_18290);
or U18664 (N_18664,N_18416,N_18177);
nor U18665 (N_18665,N_18365,N_18156);
nor U18666 (N_18666,N_18042,N_18008);
nor U18667 (N_18667,N_18006,N_18026);
and U18668 (N_18668,N_18072,N_18078);
nand U18669 (N_18669,N_18262,N_18275);
and U18670 (N_18670,N_18208,N_18234);
and U18671 (N_18671,N_18323,N_18240);
nor U18672 (N_18672,N_18444,N_18425);
nor U18673 (N_18673,N_18233,N_18194);
xnor U18674 (N_18674,N_18321,N_18139);
nand U18675 (N_18675,N_18056,N_18179);
and U18676 (N_18676,N_18127,N_18013);
xor U18677 (N_18677,N_18305,N_18489);
or U18678 (N_18678,N_18409,N_18071);
or U18679 (N_18679,N_18049,N_18142);
and U18680 (N_18680,N_18210,N_18253);
and U18681 (N_18681,N_18120,N_18227);
nand U18682 (N_18682,N_18463,N_18181);
or U18683 (N_18683,N_18370,N_18248);
nand U18684 (N_18684,N_18267,N_18123);
or U18685 (N_18685,N_18131,N_18076);
xor U18686 (N_18686,N_18348,N_18226);
xor U18687 (N_18687,N_18134,N_18471);
or U18688 (N_18688,N_18490,N_18331);
nor U18689 (N_18689,N_18152,N_18050);
and U18690 (N_18690,N_18202,N_18041);
or U18691 (N_18691,N_18411,N_18138);
or U18692 (N_18692,N_18077,N_18106);
or U18693 (N_18693,N_18185,N_18325);
xnor U18694 (N_18694,N_18336,N_18164);
nand U18695 (N_18695,N_18472,N_18031);
and U18696 (N_18696,N_18286,N_18224);
and U18697 (N_18697,N_18448,N_18021);
and U18698 (N_18698,N_18088,N_18477);
xor U18699 (N_18699,N_18102,N_18172);
nor U18700 (N_18700,N_18067,N_18075);
nand U18701 (N_18701,N_18219,N_18154);
xor U18702 (N_18702,N_18316,N_18467);
and U18703 (N_18703,N_18105,N_18378);
and U18704 (N_18704,N_18281,N_18239);
and U18705 (N_18705,N_18136,N_18174);
nand U18706 (N_18706,N_18018,N_18435);
nor U18707 (N_18707,N_18396,N_18054);
nand U18708 (N_18708,N_18200,N_18090);
nor U18709 (N_18709,N_18149,N_18462);
nor U18710 (N_18710,N_18333,N_18432);
nand U18711 (N_18711,N_18283,N_18014);
nand U18712 (N_18712,N_18213,N_18187);
xor U18713 (N_18713,N_18216,N_18499);
or U18714 (N_18714,N_18274,N_18062);
xnor U18715 (N_18715,N_18392,N_18169);
nand U18716 (N_18716,N_18341,N_18053);
and U18717 (N_18717,N_18358,N_18434);
nand U18718 (N_18718,N_18068,N_18027);
and U18719 (N_18719,N_18251,N_18355);
or U18720 (N_18720,N_18246,N_18063);
and U18721 (N_18721,N_18487,N_18322);
nand U18722 (N_18722,N_18249,N_18217);
xnor U18723 (N_18723,N_18052,N_18150);
nor U18724 (N_18724,N_18269,N_18478);
xnor U18725 (N_18725,N_18410,N_18098);
nand U18726 (N_18726,N_18140,N_18024);
and U18727 (N_18727,N_18433,N_18101);
or U18728 (N_18728,N_18074,N_18186);
nor U18729 (N_18729,N_18207,N_18023);
and U18730 (N_18730,N_18314,N_18375);
or U18731 (N_18731,N_18132,N_18235);
or U18732 (N_18732,N_18104,N_18277);
nor U18733 (N_18733,N_18415,N_18480);
xor U18734 (N_18734,N_18114,N_18354);
and U18735 (N_18735,N_18010,N_18099);
and U18736 (N_18736,N_18351,N_18083);
xor U18737 (N_18737,N_18468,N_18473);
xnor U18738 (N_18738,N_18449,N_18390);
or U18739 (N_18739,N_18162,N_18394);
nor U18740 (N_18740,N_18190,N_18482);
or U18741 (N_18741,N_18484,N_18464);
and U18742 (N_18742,N_18457,N_18497);
nand U18743 (N_18743,N_18284,N_18427);
or U18744 (N_18744,N_18350,N_18032);
xor U18745 (N_18745,N_18320,N_18128);
xor U18746 (N_18746,N_18146,N_18124);
and U18747 (N_18747,N_18059,N_18221);
nand U18748 (N_18748,N_18130,N_18237);
nor U18749 (N_18749,N_18452,N_18404);
or U18750 (N_18750,N_18312,N_18268);
xnor U18751 (N_18751,N_18273,N_18475);
or U18752 (N_18752,N_18016,N_18379);
nand U18753 (N_18753,N_18215,N_18431);
and U18754 (N_18754,N_18052,N_18183);
nand U18755 (N_18755,N_18391,N_18227);
xor U18756 (N_18756,N_18055,N_18131);
nor U18757 (N_18757,N_18111,N_18341);
nand U18758 (N_18758,N_18028,N_18187);
xor U18759 (N_18759,N_18158,N_18358);
nor U18760 (N_18760,N_18068,N_18422);
or U18761 (N_18761,N_18111,N_18227);
or U18762 (N_18762,N_18377,N_18302);
or U18763 (N_18763,N_18051,N_18109);
nand U18764 (N_18764,N_18340,N_18411);
and U18765 (N_18765,N_18431,N_18485);
xor U18766 (N_18766,N_18189,N_18495);
xnor U18767 (N_18767,N_18266,N_18313);
or U18768 (N_18768,N_18139,N_18484);
nand U18769 (N_18769,N_18113,N_18272);
and U18770 (N_18770,N_18381,N_18162);
xnor U18771 (N_18771,N_18132,N_18299);
xor U18772 (N_18772,N_18001,N_18209);
xnor U18773 (N_18773,N_18487,N_18319);
nand U18774 (N_18774,N_18043,N_18442);
and U18775 (N_18775,N_18127,N_18317);
or U18776 (N_18776,N_18052,N_18130);
nor U18777 (N_18777,N_18355,N_18366);
or U18778 (N_18778,N_18124,N_18355);
nor U18779 (N_18779,N_18487,N_18001);
and U18780 (N_18780,N_18342,N_18207);
nor U18781 (N_18781,N_18155,N_18493);
xor U18782 (N_18782,N_18280,N_18166);
nor U18783 (N_18783,N_18040,N_18326);
nand U18784 (N_18784,N_18015,N_18058);
nand U18785 (N_18785,N_18371,N_18002);
nor U18786 (N_18786,N_18000,N_18483);
xnor U18787 (N_18787,N_18036,N_18285);
or U18788 (N_18788,N_18480,N_18463);
nand U18789 (N_18789,N_18252,N_18333);
nor U18790 (N_18790,N_18368,N_18323);
xnor U18791 (N_18791,N_18299,N_18432);
nand U18792 (N_18792,N_18262,N_18202);
nor U18793 (N_18793,N_18454,N_18124);
nand U18794 (N_18794,N_18384,N_18172);
nor U18795 (N_18795,N_18128,N_18134);
or U18796 (N_18796,N_18041,N_18217);
and U18797 (N_18797,N_18084,N_18246);
and U18798 (N_18798,N_18382,N_18007);
or U18799 (N_18799,N_18248,N_18019);
and U18800 (N_18800,N_18089,N_18473);
and U18801 (N_18801,N_18333,N_18115);
nor U18802 (N_18802,N_18042,N_18344);
nand U18803 (N_18803,N_18233,N_18035);
nor U18804 (N_18804,N_18359,N_18445);
or U18805 (N_18805,N_18262,N_18133);
nor U18806 (N_18806,N_18182,N_18365);
xor U18807 (N_18807,N_18336,N_18419);
nor U18808 (N_18808,N_18022,N_18420);
nand U18809 (N_18809,N_18317,N_18039);
xor U18810 (N_18810,N_18425,N_18323);
or U18811 (N_18811,N_18144,N_18038);
xnor U18812 (N_18812,N_18189,N_18028);
xor U18813 (N_18813,N_18147,N_18372);
or U18814 (N_18814,N_18144,N_18235);
xnor U18815 (N_18815,N_18347,N_18190);
xnor U18816 (N_18816,N_18362,N_18052);
and U18817 (N_18817,N_18193,N_18109);
nand U18818 (N_18818,N_18241,N_18354);
or U18819 (N_18819,N_18323,N_18335);
or U18820 (N_18820,N_18062,N_18123);
nand U18821 (N_18821,N_18179,N_18037);
and U18822 (N_18822,N_18352,N_18457);
nand U18823 (N_18823,N_18449,N_18416);
nor U18824 (N_18824,N_18445,N_18241);
xor U18825 (N_18825,N_18229,N_18082);
nand U18826 (N_18826,N_18251,N_18376);
xor U18827 (N_18827,N_18007,N_18011);
or U18828 (N_18828,N_18155,N_18160);
nor U18829 (N_18829,N_18412,N_18083);
nand U18830 (N_18830,N_18069,N_18444);
or U18831 (N_18831,N_18193,N_18162);
or U18832 (N_18832,N_18423,N_18083);
and U18833 (N_18833,N_18083,N_18337);
or U18834 (N_18834,N_18423,N_18052);
nor U18835 (N_18835,N_18035,N_18300);
nand U18836 (N_18836,N_18398,N_18214);
xnor U18837 (N_18837,N_18055,N_18286);
nor U18838 (N_18838,N_18398,N_18295);
xor U18839 (N_18839,N_18056,N_18446);
or U18840 (N_18840,N_18152,N_18019);
or U18841 (N_18841,N_18260,N_18192);
xnor U18842 (N_18842,N_18438,N_18088);
nand U18843 (N_18843,N_18060,N_18103);
and U18844 (N_18844,N_18349,N_18256);
or U18845 (N_18845,N_18019,N_18425);
nand U18846 (N_18846,N_18138,N_18432);
nor U18847 (N_18847,N_18153,N_18489);
and U18848 (N_18848,N_18018,N_18129);
nand U18849 (N_18849,N_18279,N_18306);
and U18850 (N_18850,N_18486,N_18267);
xor U18851 (N_18851,N_18468,N_18278);
or U18852 (N_18852,N_18187,N_18171);
nor U18853 (N_18853,N_18326,N_18441);
xnor U18854 (N_18854,N_18436,N_18357);
or U18855 (N_18855,N_18396,N_18126);
nand U18856 (N_18856,N_18253,N_18307);
xor U18857 (N_18857,N_18023,N_18393);
and U18858 (N_18858,N_18401,N_18325);
nand U18859 (N_18859,N_18005,N_18358);
xor U18860 (N_18860,N_18002,N_18249);
xnor U18861 (N_18861,N_18356,N_18485);
and U18862 (N_18862,N_18136,N_18212);
nand U18863 (N_18863,N_18357,N_18242);
and U18864 (N_18864,N_18301,N_18273);
xnor U18865 (N_18865,N_18218,N_18433);
nand U18866 (N_18866,N_18048,N_18440);
and U18867 (N_18867,N_18180,N_18093);
and U18868 (N_18868,N_18413,N_18088);
or U18869 (N_18869,N_18304,N_18345);
nand U18870 (N_18870,N_18381,N_18436);
nand U18871 (N_18871,N_18083,N_18399);
or U18872 (N_18872,N_18397,N_18143);
xor U18873 (N_18873,N_18447,N_18023);
or U18874 (N_18874,N_18140,N_18344);
and U18875 (N_18875,N_18354,N_18098);
nand U18876 (N_18876,N_18184,N_18052);
nand U18877 (N_18877,N_18081,N_18487);
nor U18878 (N_18878,N_18078,N_18212);
xor U18879 (N_18879,N_18338,N_18319);
or U18880 (N_18880,N_18014,N_18441);
nor U18881 (N_18881,N_18215,N_18213);
xor U18882 (N_18882,N_18394,N_18385);
and U18883 (N_18883,N_18425,N_18329);
nor U18884 (N_18884,N_18333,N_18442);
or U18885 (N_18885,N_18324,N_18144);
and U18886 (N_18886,N_18463,N_18451);
or U18887 (N_18887,N_18133,N_18166);
and U18888 (N_18888,N_18447,N_18383);
nor U18889 (N_18889,N_18208,N_18150);
nor U18890 (N_18890,N_18035,N_18208);
nand U18891 (N_18891,N_18060,N_18330);
or U18892 (N_18892,N_18271,N_18011);
or U18893 (N_18893,N_18076,N_18343);
and U18894 (N_18894,N_18234,N_18000);
nand U18895 (N_18895,N_18026,N_18380);
xor U18896 (N_18896,N_18393,N_18138);
or U18897 (N_18897,N_18026,N_18246);
nand U18898 (N_18898,N_18139,N_18187);
and U18899 (N_18899,N_18232,N_18272);
or U18900 (N_18900,N_18102,N_18141);
xor U18901 (N_18901,N_18078,N_18304);
or U18902 (N_18902,N_18395,N_18001);
nor U18903 (N_18903,N_18340,N_18001);
nor U18904 (N_18904,N_18339,N_18270);
nor U18905 (N_18905,N_18096,N_18440);
xnor U18906 (N_18906,N_18023,N_18128);
nor U18907 (N_18907,N_18106,N_18253);
nor U18908 (N_18908,N_18472,N_18006);
xnor U18909 (N_18909,N_18152,N_18121);
or U18910 (N_18910,N_18385,N_18225);
xor U18911 (N_18911,N_18114,N_18301);
xor U18912 (N_18912,N_18035,N_18365);
or U18913 (N_18913,N_18175,N_18215);
nor U18914 (N_18914,N_18344,N_18129);
nor U18915 (N_18915,N_18281,N_18023);
nand U18916 (N_18916,N_18053,N_18346);
xor U18917 (N_18917,N_18135,N_18464);
nand U18918 (N_18918,N_18464,N_18258);
xnor U18919 (N_18919,N_18250,N_18113);
or U18920 (N_18920,N_18060,N_18066);
and U18921 (N_18921,N_18077,N_18434);
or U18922 (N_18922,N_18192,N_18472);
nor U18923 (N_18923,N_18298,N_18489);
nand U18924 (N_18924,N_18389,N_18184);
and U18925 (N_18925,N_18041,N_18190);
and U18926 (N_18926,N_18095,N_18415);
nor U18927 (N_18927,N_18337,N_18313);
or U18928 (N_18928,N_18016,N_18288);
xnor U18929 (N_18929,N_18134,N_18374);
nor U18930 (N_18930,N_18120,N_18376);
or U18931 (N_18931,N_18188,N_18451);
nand U18932 (N_18932,N_18477,N_18495);
xor U18933 (N_18933,N_18136,N_18106);
nand U18934 (N_18934,N_18347,N_18079);
xnor U18935 (N_18935,N_18465,N_18388);
or U18936 (N_18936,N_18275,N_18244);
nor U18937 (N_18937,N_18123,N_18315);
xnor U18938 (N_18938,N_18309,N_18081);
nand U18939 (N_18939,N_18222,N_18110);
nand U18940 (N_18940,N_18022,N_18020);
nor U18941 (N_18941,N_18479,N_18494);
nor U18942 (N_18942,N_18185,N_18118);
nor U18943 (N_18943,N_18164,N_18294);
or U18944 (N_18944,N_18276,N_18110);
nor U18945 (N_18945,N_18143,N_18171);
and U18946 (N_18946,N_18334,N_18157);
or U18947 (N_18947,N_18418,N_18047);
and U18948 (N_18948,N_18390,N_18043);
or U18949 (N_18949,N_18277,N_18487);
nor U18950 (N_18950,N_18053,N_18426);
nand U18951 (N_18951,N_18471,N_18049);
xor U18952 (N_18952,N_18163,N_18429);
nor U18953 (N_18953,N_18482,N_18144);
nor U18954 (N_18954,N_18352,N_18288);
or U18955 (N_18955,N_18470,N_18318);
xor U18956 (N_18956,N_18467,N_18176);
nor U18957 (N_18957,N_18257,N_18110);
or U18958 (N_18958,N_18015,N_18103);
nand U18959 (N_18959,N_18289,N_18163);
or U18960 (N_18960,N_18212,N_18482);
xor U18961 (N_18961,N_18076,N_18420);
nor U18962 (N_18962,N_18202,N_18394);
nand U18963 (N_18963,N_18149,N_18495);
nor U18964 (N_18964,N_18087,N_18214);
xor U18965 (N_18965,N_18491,N_18018);
and U18966 (N_18966,N_18364,N_18495);
nand U18967 (N_18967,N_18200,N_18179);
nand U18968 (N_18968,N_18391,N_18238);
nand U18969 (N_18969,N_18190,N_18035);
nand U18970 (N_18970,N_18082,N_18097);
nor U18971 (N_18971,N_18239,N_18484);
xnor U18972 (N_18972,N_18132,N_18475);
nand U18973 (N_18973,N_18499,N_18259);
xnor U18974 (N_18974,N_18449,N_18042);
nand U18975 (N_18975,N_18499,N_18162);
and U18976 (N_18976,N_18088,N_18182);
xnor U18977 (N_18977,N_18297,N_18334);
xnor U18978 (N_18978,N_18242,N_18095);
and U18979 (N_18979,N_18041,N_18441);
nor U18980 (N_18980,N_18183,N_18011);
xor U18981 (N_18981,N_18041,N_18115);
xor U18982 (N_18982,N_18326,N_18464);
nor U18983 (N_18983,N_18379,N_18497);
nand U18984 (N_18984,N_18283,N_18214);
or U18985 (N_18985,N_18185,N_18035);
nand U18986 (N_18986,N_18052,N_18471);
and U18987 (N_18987,N_18439,N_18430);
nand U18988 (N_18988,N_18062,N_18014);
or U18989 (N_18989,N_18121,N_18141);
or U18990 (N_18990,N_18416,N_18312);
or U18991 (N_18991,N_18225,N_18490);
or U18992 (N_18992,N_18432,N_18214);
nor U18993 (N_18993,N_18197,N_18177);
nand U18994 (N_18994,N_18063,N_18046);
nand U18995 (N_18995,N_18064,N_18014);
nor U18996 (N_18996,N_18407,N_18459);
and U18997 (N_18997,N_18496,N_18196);
and U18998 (N_18998,N_18032,N_18451);
and U18999 (N_18999,N_18253,N_18284);
xor U19000 (N_19000,N_18839,N_18818);
nor U19001 (N_19001,N_18817,N_18815);
nand U19002 (N_19002,N_18510,N_18523);
nor U19003 (N_19003,N_18658,N_18674);
nand U19004 (N_19004,N_18760,N_18643);
or U19005 (N_19005,N_18686,N_18528);
or U19006 (N_19006,N_18948,N_18979);
nand U19007 (N_19007,N_18929,N_18729);
and U19008 (N_19008,N_18507,N_18649);
xor U19009 (N_19009,N_18675,N_18834);
and U19010 (N_19010,N_18813,N_18707);
nand U19011 (N_19011,N_18776,N_18984);
or U19012 (N_19012,N_18607,N_18541);
and U19013 (N_19013,N_18787,N_18924);
or U19014 (N_19014,N_18986,N_18841);
and U19015 (N_19015,N_18951,N_18705);
nor U19016 (N_19016,N_18520,N_18808);
or U19017 (N_19017,N_18862,N_18608);
xnor U19018 (N_19018,N_18648,N_18881);
nand U19019 (N_19019,N_18676,N_18930);
nand U19020 (N_19020,N_18718,N_18927);
or U19021 (N_19021,N_18548,N_18756);
xnor U19022 (N_19022,N_18857,N_18645);
and U19023 (N_19023,N_18698,N_18701);
nand U19024 (N_19024,N_18856,N_18590);
nor U19025 (N_19025,N_18672,N_18943);
nand U19026 (N_19026,N_18653,N_18614);
and U19027 (N_19027,N_18942,N_18646);
and U19028 (N_19028,N_18662,N_18552);
nor U19029 (N_19029,N_18990,N_18956);
nand U19030 (N_19030,N_18636,N_18556);
nor U19031 (N_19031,N_18560,N_18812);
or U19032 (N_19032,N_18750,N_18960);
or U19033 (N_19033,N_18723,N_18621);
xor U19034 (N_19034,N_18780,N_18714);
nand U19035 (N_19035,N_18522,N_18823);
nor U19036 (N_19036,N_18702,N_18761);
xor U19037 (N_19037,N_18816,N_18605);
nand U19038 (N_19038,N_18603,N_18897);
nand U19039 (N_19039,N_18858,N_18850);
xor U19040 (N_19040,N_18641,N_18545);
and U19041 (N_19041,N_18872,N_18525);
nor U19042 (N_19042,N_18963,N_18696);
nand U19043 (N_19043,N_18503,N_18855);
xnor U19044 (N_19044,N_18715,N_18810);
nor U19045 (N_19045,N_18562,N_18952);
and U19046 (N_19046,N_18684,N_18907);
and U19047 (N_19047,N_18671,N_18501);
nand U19048 (N_19048,N_18721,N_18814);
and U19049 (N_19049,N_18728,N_18921);
nand U19050 (N_19050,N_18667,N_18974);
nand U19051 (N_19051,N_18518,N_18690);
or U19052 (N_19052,N_18802,N_18789);
nor U19053 (N_19053,N_18772,N_18899);
nand U19054 (N_19054,N_18546,N_18688);
nand U19055 (N_19055,N_18898,N_18682);
and U19056 (N_19056,N_18766,N_18708);
nand U19057 (N_19057,N_18679,N_18628);
xnor U19058 (N_19058,N_18759,N_18773);
or U19059 (N_19059,N_18741,N_18629);
and U19060 (N_19060,N_18807,N_18875);
and U19061 (N_19061,N_18797,N_18947);
or U19062 (N_19062,N_18865,N_18526);
and U19063 (N_19063,N_18642,N_18965);
and U19064 (N_19064,N_18745,N_18835);
nand U19065 (N_19065,N_18803,N_18615);
xnor U19066 (N_19066,N_18829,N_18717);
nand U19067 (N_19067,N_18555,N_18731);
xor U19068 (N_19068,N_18844,N_18925);
xor U19069 (N_19069,N_18632,N_18508);
nor U19070 (N_19070,N_18768,N_18999);
or U19071 (N_19071,N_18704,N_18763);
and U19072 (N_19072,N_18650,N_18864);
xor U19073 (N_19073,N_18587,N_18551);
xnor U19074 (N_19074,N_18976,N_18524);
or U19075 (N_19075,N_18738,N_18683);
nor U19076 (N_19076,N_18962,N_18565);
xnor U19077 (N_19077,N_18680,N_18712);
nor U19078 (N_19078,N_18842,N_18874);
or U19079 (N_19079,N_18693,N_18668);
or U19080 (N_19080,N_18692,N_18536);
nor U19081 (N_19081,N_18740,N_18700);
xnor U19082 (N_19082,N_18509,N_18737);
nor U19083 (N_19083,N_18877,N_18901);
or U19084 (N_19084,N_18957,N_18848);
nand U19085 (N_19085,N_18977,N_18845);
nor U19086 (N_19086,N_18847,N_18594);
and U19087 (N_19087,N_18549,N_18946);
or U19088 (N_19088,N_18982,N_18846);
xnor U19089 (N_19089,N_18840,N_18611);
nand U19090 (N_19090,N_18869,N_18609);
nor U19091 (N_19091,N_18623,N_18697);
nor U19092 (N_19092,N_18695,N_18935);
nor U19093 (N_19093,N_18751,N_18970);
or U19094 (N_19094,N_18997,N_18767);
xor U19095 (N_19095,N_18870,N_18588);
and U19096 (N_19096,N_18863,N_18900);
and U19097 (N_19097,N_18581,N_18861);
and U19098 (N_19098,N_18585,N_18755);
or U19099 (N_19099,N_18833,N_18558);
nor U19100 (N_19100,N_18639,N_18804);
or U19101 (N_19101,N_18617,N_18630);
nor U19102 (N_19102,N_18533,N_18905);
xor U19103 (N_19103,N_18891,N_18544);
nand U19104 (N_19104,N_18795,N_18706);
or U19105 (N_19105,N_18537,N_18564);
xnor U19106 (N_19106,N_18996,N_18506);
and U19107 (N_19107,N_18961,N_18867);
or U19108 (N_19108,N_18973,N_18655);
and U19109 (N_19109,N_18580,N_18878);
and U19110 (N_19110,N_18792,N_18566);
xor U19111 (N_19111,N_18993,N_18687);
xor U19112 (N_19112,N_18988,N_18915);
xnor U19113 (N_19113,N_18757,N_18589);
nor U19114 (N_19114,N_18866,N_18519);
or U19115 (N_19115,N_18868,N_18652);
or U19116 (N_19116,N_18527,N_18644);
or U19117 (N_19117,N_18681,N_18828);
and U19118 (N_19118,N_18592,N_18955);
xnor U19119 (N_19119,N_18547,N_18719);
or U19120 (N_19120,N_18659,N_18570);
or U19121 (N_19121,N_18673,N_18651);
or U19122 (N_19122,N_18784,N_18601);
nand U19123 (N_19123,N_18599,N_18742);
or U19124 (N_19124,N_18876,N_18666);
xor U19125 (N_19125,N_18620,N_18578);
xor U19126 (N_19126,N_18618,N_18554);
nor U19127 (N_19127,N_18725,N_18710);
and U19128 (N_19128,N_18910,N_18516);
and U19129 (N_19129,N_18535,N_18663);
xnor U19130 (N_19130,N_18969,N_18783);
nor U19131 (N_19131,N_18656,N_18769);
and U19132 (N_19132,N_18532,N_18975);
nor U19133 (N_19133,N_18511,N_18699);
nand U19134 (N_19134,N_18906,N_18604);
or U19135 (N_19135,N_18794,N_18916);
nor U19136 (N_19136,N_18531,N_18574);
nand U19137 (N_19137,N_18933,N_18782);
xor U19138 (N_19138,N_18597,N_18972);
or U19139 (N_19139,N_18515,N_18568);
nand U19140 (N_19140,N_18538,N_18572);
and U19141 (N_19141,N_18980,N_18851);
nor U19142 (N_19142,N_18805,N_18770);
nor U19143 (N_19143,N_18911,N_18923);
xor U19144 (N_19144,N_18938,N_18934);
nand U19145 (N_19145,N_18665,N_18716);
or U19146 (N_19146,N_18920,N_18600);
nand U19147 (N_19147,N_18966,N_18514);
nand U19148 (N_19148,N_18824,N_18879);
nor U19149 (N_19149,N_18912,N_18678);
nand U19150 (N_19150,N_18799,N_18624);
xor U19151 (N_19151,N_18854,N_18837);
nor U19152 (N_19152,N_18557,N_18638);
and U19153 (N_19153,N_18932,N_18550);
nand U19154 (N_19154,N_18529,N_18567);
and U19155 (N_19155,N_18894,N_18505);
and U19156 (N_19156,N_18762,N_18513);
or U19157 (N_19157,N_18918,N_18949);
xnor U19158 (N_19158,N_18827,N_18853);
and U19159 (N_19159,N_18904,N_18991);
xnor U19160 (N_19160,N_18754,N_18909);
or U19161 (N_19161,N_18998,N_18595);
and U19162 (N_19162,N_18749,N_18664);
and U19163 (N_19163,N_18553,N_18753);
and U19164 (N_19164,N_18633,N_18809);
and U19165 (N_19165,N_18896,N_18945);
xor U19166 (N_19166,N_18978,N_18563);
xnor U19167 (N_19167,N_18832,N_18826);
nand U19168 (N_19168,N_18720,N_18631);
nand U19169 (N_19169,N_18542,N_18882);
and U19170 (N_19170,N_18724,N_18661);
and U19171 (N_19171,N_18886,N_18821);
nor U19172 (N_19172,N_18627,N_18579);
xnor U19173 (N_19173,N_18959,N_18625);
xnor U19174 (N_19174,N_18774,N_18781);
nor U19175 (N_19175,N_18722,N_18994);
or U19176 (N_19176,N_18791,N_18540);
and U19177 (N_19177,N_18936,N_18939);
and U19178 (N_19178,N_18559,N_18836);
or U19179 (N_19179,N_18747,N_18602);
and U19180 (N_19180,N_18591,N_18806);
or U19181 (N_19181,N_18670,N_18902);
nand U19182 (N_19182,N_18765,N_18941);
xnor U19183 (N_19183,N_18634,N_18968);
or U19184 (N_19184,N_18539,N_18576);
nor U19185 (N_19185,N_18786,N_18606);
or U19186 (N_19186,N_18831,N_18596);
xnor U19187 (N_19187,N_18657,N_18711);
and U19188 (N_19188,N_18793,N_18830);
nand U19189 (N_19189,N_18852,N_18800);
xor U19190 (N_19190,N_18888,N_18612);
nor U19191 (N_19191,N_18992,N_18859);
xnor U19192 (N_19192,N_18732,N_18796);
nand U19193 (N_19193,N_18801,N_18640);
nor U19194 (N_19194,N_18903,N_18504);
or U19195 (N_19195,N_18619,N_18825);
nor U19196 (N_19196,N_18713,N_18889);
nor U19197 (N_19197,N_18521,N_18569);
xor U19198 (N_19198,N_18953,N_18798);
nor U19199 (N_19199,N_18727,N_18735);
and U19200 (N_19200,N_18860,N_18985);
and U19201 (N_19201,N_18571,N_18981);
and U19202 (N_19202,N_18779,N_18622);
xnor U19203 (N_19203,N_18635,N_18892);
nor U19204 (N_19204,N_18843,N_18733);
xor U19205 (N_19205,N_18734,N_18928);
nor U19206 (N_19206,N_18995,N_18694);
nor U19207 (N_19207,N_18983,N_18512);
xor U19208 (N_19208,N_18849,N_18613);
or U19209 (N_19209,N_18744,N_18880);
xor U19210 (N_19210,N_18883,N_18575);
xnor U19211 (N_19211,N_18616,N_18660);
and U19212 (N_19212,N_18730,N_18967);
xnor U19213 (N_19213,N_18954,N_18819);
nand U19214 (N_19214,N_18873,N_18530);
and U19215 (N_19215,N_18736,N_18626);
nor U19216 (N_19216,N_18777,N_18598);
nor U19217 (N_19217,N_18987,N_18669);
nand U19218 (N_19218,N_18950,N_18940);
xor U19219 (N_19219,N_18726,N_18914);
xnor U19220 (N_19220,N_18913,N_18677);
and U19221 (N_19221,N_18637,N_18790);
nand U19222 (N_19222,N_18778,N_18893);
xor U19223 (N_19223,N_18811,N_18517);
xor U19224 (N_19224,N_18654,N_18890);
or U19225 (N_19225,N_18593,N_18771);
or U19226 (N_19226,N_18647,N_18871);
nand U19227 (N_19227,N_18746,N_18944);
nor U19228 (N_19228,N_18917,N_18764);
or U19229 (N_19229,N_18788,N_18820);
or U19230 (N_19230,N_18691,N_18887);
nor U19231 (N_19231,N_18919,N_18610);
nor U19232 (N_19232,N_18895,N_18752);
or U19233 (N_19233,N_18931,N_18838);
or U19234 (N_19234,N_18926,N_18577);
or U19235 (N_19235,N_18582,N_18586);
xor U19236 (N_19236,N_18971,N_18937);
nor U19237 (N_19237,N_18908,N_18785);
nand U19238 (N_19238,N_18502,N_18743);
and U19239 (N_19239,N_18775,N_18758);
or U19240 (N_19240,N_18709,N_18703);
xnor U19241 (N_19241,N_18822,N_18561);
or U19242 (N_19242,N_18885,N_18748);
nor U19243 (N_19243,N_18884,N_18584);
nor U19244 (N_19244,N_18739,N_18958);
nor U19245 (N_19245,N_18534,N_18500);
and U19246 (N_19246,N_18964,N_18685);
xor U19247 (N_19247,N_18689,N_18922);
nand U19248 (N_19248,N_18543,N_18573);
nand U19249 (N_19249,N_18989,N_18583);
and U19250 (N_19250,N_18523,N_18564);
nand U19251 (N_19251,N_18740,N_18842);
or U19252 (N_19252,N_18634,N_18684);
and U19253 (N_19253,N_18963,N_18583);
xnor U19254 (N_19254,N_18808,N_18511);
nor U19255 (N_19255,N_18544,N_18843);
and U19256 (N_19256,N_18823,N_18921);
xnor U19257 (N_19257,N_18683,N_18531);
nor U19258 (N_19258,N_18913,N_18708);
nor U19259 (N_19259,N_18809,N_18865);
nand U19260 (N_19260,N_18560,N_18867);
or U19261 (N_19261,N_18740,N_18985);
xnor U19262 (N_19262,N_18515,N_18890);
xor U19263 (N_19263,N_18645,N_18548);
xor U19264 (N_19264,N_18832,N_18648);
xnor U19265 (N_19265,N_18584,N_18887);
and U19266 (N_19266,N_18833,N_18658);
nand U19267 (N_19267,N_18565,N_18574);
or U19268 (N_19268,N_18813,N_18857);
nand U19269 (N_19269,N_18752,N_18563);
or U19270 (N_19270,N_18677,N_18610);
nor U19271 (N_19271,N_18628,N_18857);
xor U19272 (N_19272,N_18891,N_18984);
and U19273 (N_19273,N_18700,N_18648);
and U19274 (N_19274,N_18561,N_18961);
and U19275 (N_19275,N_18551,N_18813);
nor U19276 (N_19276,N_18835,N_18588);
or U19277 (N_19277,N_18864,N_18882);
xor U19278 (N_19278,N_18741,N_18838);
nand U19279 (N_19279,N_18827,N_18577);
xor U19280 (N_19280,N_18667,N_18787);
xnor U19281 (N_19281,N_18990,N_18967);
xor U19282 (N_19282,N_18507,N_18522);
nand U19283 (N_19283,N_18562,N_18536);
nand U19284 (N_19284,N_18710,N_18803);
xnor U19285 (N_19285,N_18976,N_18886);
xor U19286 (N_19286,N_18795,N_18554);
nand U19287 (N_19287,N_18690,N_18516);
and U19288 (N_19288,N_18951,N_18618);
or U19289 (N_19289,N_18882,N_18581);
nor U19290 (N_19290,N_18809,N_18648);
nand U19291 (N_19291,N_18875,N_18666);
nor U19292 (N_19292,N_18878,N_18657);
nor U19293 (N_19293,N_18563,N_18557);
and U19294 (N_19294,N_18631,N_18898);
nand U19295 (N_19295,N_18681,N_18867);
xor U19296 (N_19296,N_18850,N_18560);
nor U19297 (N_19297,N_18699,N_18949);
nand U19298 (N_19298,N_18928,N_18730);
or U19299 (N_19299,N_18611,N_18592);
nor U19300 (N_19300,N_18889,N_18894);
nor U19301 (N_19301,N_18574,N_18622);
or U19302 (N_19302,N_18683,N_18934);
xor U19303 (N_19303,N_18996,N_18565);
or U19304 (N_19304,N_18972,N_18511);
xnor U19305 (N_19305,N_18870,N_18872);
nand U19306 (N_19306,N_18898,N_18716);
xnor U19307 (N_19307,N_18923,N_18516);
nand U19308 (N_19308,N_18713,N_18840);
nand U19309 (N_19309,N_18793,N_18611);
or U19310 (N_19310,N_18548,N_18888);
nor U19311 (N_19311,N_18921,N_18969);
xor U19312 (N_19312,N_18786,N_18668);
xor U19313 (N_19313,N_18768,N_18893);
or U19314 (N_19314,N_18860,N_18535);
and U19315 (N_19315,N_18684,N_18860);
and U19316 (N_19316,N_18615,N_18890);
xnor U19317 (N_19317,N_18639,N_18613);
nand U19318 (N_19318,N_18979,N_18937);
nand U19319 (N_19319,N_18590,N_18796);
nand U19320 (N_19320,N_18614,N_18578);
or U19321 (N_19321,N_18862,N_18972);
and U19322 (N_19322,N_18867,N_18502);
nor U19323 (N_19323,N_18744,N_18894);
nor U19324 (N_19324,N_18673,N_18502);
or U19325 (N_19325,N_18551,N_18989);
or U19326 (N_19326,N_18944,N_18943);
nand U19327 (N_19327,N_18544,N_18932);
or U19328 (N_19328,N_18564,N_18968);
nor U19329 (N_19329,N_18770,N_18976);
or U19330 (N_19330,N_18754,N_18569);
nand U19331 (N_19331,N_18747,N_18928);
nor U19332 (N_19332,N_18956,N_18977);
xnor U19333 (N_19333,N_18954,N_18875);
and U19334 (N_19334,N_18663,N_18639);
or U19335 (N_19335,N_18705,N_18764);
and U19336 (N_19336,N_18926,N_18994);
nor U19337 (N_19337,N_18914,N_18832);
xnor U19338 (N_19338,N_18980,N_18522);
or U19339 (N_19339,N_18809,N_18787);
or U19340 (N_19340,N_18921,N_18511);
or U19341 (N_19341,N_18701,N_18702);
xnor U19342 (N_19342,N_18991,N_18503);
nand U19343 (N_19343,N_18907,N_18950);
nor U19344 (N_19344,N_18705,N_18659);
and U19345 (N_19345,N_18917,N_18541);
and U19346 (N_19346,N_18567,N_18821);
or U19347 (N_19347,N_18671,N_18967);
and U19348 (N_19348,N_18880,N_18909);
or U19349 (N_19349,N_18769,N_18954);
or U19350 (N_19350,N_18931,N_18722);
xor U19351 (N_19351,N_18675,N_18809);
xor U19352 (N_19352,N_18829,N_18848);
and U19353 (N_19353,N_18979,N_18814);
xnor U19354 (N_19354,N_18930,N_18728);
and U19355 (N_19355,N_18949,N_18991);
nand U19356 (N_19356,N_18988,N_18919);
nor U19357 (N_19357,N_18639,N_18865);
xnor U19358 (N_19358,N_18576,N_18561);
nor U19359 (N_19359,N_18625,N_18508);
xnor U19360 (N_19360,N_18835,N_18995);
nand U19361 (N_19361,N_18558,N_18838);
nand U19362 (N_19362,N_18784,N_18877);
xor U19363 (N_19363,N_18787,N_18973);
and U19364 (N_19364,N_18514,N_18951);
xnor U19365 (N_19365,N_18796,N_18714);
nor U19366 (N_19366,N_18573,N_18747);
nand U19367 (N_19367,N_18921,N_18560);
or U19368 (N_19368,N_18728,N_18617);
nor U19369 (N_19369,N_18665,N_18749);
or U19370 (N_19370,N_18909,N_18621);
nand U19371 (N_19371,N_18661,N_18960);
nor U19372 (N_19372,N_18876,N_18576);
nand U19373 (N_19373,N_18631,N_18646);
nor U19374 (N_19374,N_18985,N_18780);
or U19375 (N_19375,N_18565,N_18539);
nor U19376 (N_19376,N_18695,N_18612);
or U19377 (N_19377,N_18735,N_18601);
and U19378 (N_19378,N_18717,N_18573);
xor U19379 (N_19379,N_18959,N_18730);
and U19380 (N_19380,N_18948,N_18724);
or U19381 (N_19381,N_18654,N_18773);
and U19382 (N_19382,N_18599,N_18530);
xnor U19383 (N_19383,N_18620,N_18659);
or U19384 (N_19384,N_18771,N_18861);
xor U19385 (N_19385,N_18691,N_18537);
nor U19386 (N_19386,N_18864,N_18740);
and U19387 (N_19387,N_18802,N_18656);
xnor U19388 (N_19388,N_18760,N_18729);
and U19389 (N_19389,N_18754,N_18696);
or U19390 (N_19390,N_18730,N_18831);
nand U19391 (N_19391,N_18932,N_18978);
xor U19392 (N_19392,N_18661,N_18859);
nor U19393 (N_19393,N_18878,N_18992);
nor U19394 (N_19394,N_18872,N_18615);
nand U19395 (N_19395,N_18928,N_18564);
and U19396 (N_19396,N_18757,N_18839);
nand U19397 (N_19397,N_18731,N_18919);
or U19398 (N_19398,N_18856,N_18847);
xor U19399 (N_19399,N_18902,N_18596);
nor U19400 (N_19400,N_18950,N_18830);
nor U19401 (N_19401,N_18857,N_18808);
xor U19402 (N_19402,N_18665,N_18603);
nor U19403 (N_19403,N_18622,N_18951);
xnor U19404 (N_19404,N_18624,N_18772);
nor U19405 (N_19405,N_18597,N_18625);
or U19406 (N_19406,N_18984,N_18744);
nor U19407 (N_19407,N_18690,N_18898);
xor U19408 (N_19408,N_18866,N_18803);
or U19409 (N_19409,N_18643,N_18968);
nand U19410 (N_19410,N_18881,N_18954);
nand U19411 (N_19411,N_18739,N_18906);
nor U19412 (N_19412,N_18617,N_18898);
and U19413 (N_19413,N_18916,N_18966);
nand U19414 (N_19414,N_18671,N_18731);
nand U19415 (N_19415,N_18633,N_18502);
nor U19416 (N_19416,N_18501,N_18707);
xor U19417 (N_19417,N_18887,N_18894);
nand U19418 (N_19418,N_18828,N_18699);
or U19419 (N_19419,N_18727,N_18537);
and U19420 (N_19420,N_18936,N_18923);
or U19421 (N_19421,N_18740,N_18980);
nor U19422 (N_19422,N_18651,N_18961);
and U19423 (N_19423,N_18734,N_18853);
nand U19424 (N_19424,N_18681,N_18561);
nand U19425 (N_19425,N_18990,N_18800);
and U19426 (N_19426,N_18582,N_18944);
nand U19427 (N_19427,N_18760,N_18879);
nor U19428 (N_19428,N_18839,N_18582);
xnor U19429 (N_19429,N_18845,N_18603);
and U19430 (N_19430,N_18971,N_18975);
nand U19431 (N_19431,N_18922,N_18818);
nor U19432 (N_19432,N_18813,N_18664);
nor U19433 (N_19433,N_18788,N_18921);
nand U19434 (N_19434,N_18908,N_18657);
xor U19435 (N_19435,N_18721,N_18937);
nor U19436 (N_19436,N_18775,N_18780);
or U19437 (N_19437,N_18750,N_18550);
or U19438 (N_19438,N_18851,N_18728);
and U19439 (N_19439,N_18764,N_18582);
nor U19440 (N_19440,N_18937,N_18610);
nor U19441 (N_19441,N_18871,N_18849);
xor U19442 (N_19442,N_18593,N_18841);
xor U19443 (N_19443,N_18923,N_18895);
xor U19444 (N_19444,N_18857,N_18991);
or U19445 (N_19445,N_18984,N_18903);
nand U19446 (N_19446,N_18860,N_18796);
xor U19447 (N_19447,N_18996,N_18731);
nand U19448 (N_19448,N_18864,N_18912);
xnor U19449 (N_19449,N_18849,N_18580);
nand U19450 (N_19450,N_18932,N_18853);
nand U19451 (N_19451,N_18634,N_18572);
xor U19452 (N_19452,N_18511,N_18546);
nor U19453 (N_19453,N_18758,N_18576);
xor U19454 (N_19454,N_18822,N_18966);
and U19455 (N_19455,N_18659,N_18906);
or U19456 (N_19456,N_18521,N_18594);
nand U19457 (N_19457,N_18618,N_18674);
nand U19458 (N_19458,N_18942,N_18543);
nor U19459 (N_19459,N_18517,N_18820);
or U19460 (N_19460,N_18624,N_18669);
or U19461 (N_19461,N_18791,N_18905);
nor U19462 (N_19462,N_18722,N_18886);
and U19463 (N_19463,N_18578,N_18905);
nor U19464 (N_19464,N_18500,N_18531);
nor U19465 (N_19465,N_18537,N_18626);
or U19466 (N_19466,N_18545,N_18975);
xor U19467 (N_19467,N_18606,N_18542);
and U19468 (N_19468,N_18711,N_18803);
nand U19469 (N_19469,N_18681,N_18928);
and U19470 (N_19470,N_18524,N_18789);
and U19471 (N_19471,N_18516,N_18522);
nand U19472 (N_19472,N_18544,N_18533);
or U19473 (N_19473,N_18944,N_18677);
and U19474 (N_19474,N_18591,N_18590);
and U19475 (N_19475,N_18699,N_18505);
nand U19476 (N_19476,N_18619,N_18943);
or U19477 (N_19477,N_18865,N_18515);
xor U19478 (N_19478,N_18722,N_18570);
and U19479 (N_19479,N_18809,N_18543);
nand U19480 (N_19480,N_18679,N_18912);
nand U19481 (N_19481,N_18796,N_18622);
and U19482 (N_19482,N_18725,N_18944);
xor U19483 (N_19483,N_18980,N_18565);
or U19484 (N_19484,N_18509,N_18947);
nand U19485 (N_19485,N_18837,N_18797);
xor U19486 (N_19486,N_18872,N_18771);
or U19487 (N_19487,N_18757,N_18749);
xnor U19488 (N_19488,N_18597,N_18680);
or U19489 (N_19489,N_18730,N_18972);
and U19490 (N_19490,N_18883,N_18545);
xnor U19491 (N_19491,N_18744,N_18614);
and U19492 (N_19492,N_18847,N_18910);
nand U19493 (N_19493,N_18811,N_18528);
and U19494 (N_19494,N_18726,N_18711);
and U19495 (N_19495,N_18605,N_18726);
xor U19496 (N_19496,N_18948,N_18631);
or U19497 (N_19497,N_18563,N_18999);
xnor U19498 (N_19498,N_18531,N_18820);
nor U19499 (N_19499,N_18896,N_18566);
nor U19500 (N_19500,N_19183,N_19245);
or U19501 (N_19501,N_19468,N_19222);
or U19502 (N_19502,N_19034,N_19057);
xnor U19503 (N_19503,N_19168,N_19139);
or U19504 (N_19504,N_19163,N_19375);
nor U19505 (N_19505,N_19001,N_19033);
nand U19506 (N_19506,N_19206,N_19293);
nand U19507 (N_19507,N_19195,N_19210);
nor U19508 (N_19508,N_19241,N_19008);
xor U19509 (N_19509,N_19219,N_19157);
and U19510 (N_19510,N_19031,N_19134);
nor U19511 (N_19511,N_19388,N_19410);
nand U19512 (N_19512,N_19082,N_19327);
nor U19513 (N_19513,N_19071,N_19449);
or U19514 (N_19514,N_19416,N_19488);
and U19515 (N_19515,N_19489,N_19428);
and U19516 (N_19516,N_19102,N_19283);
and U19517 (N_19517,N_19151,N_19326);
xor U19518 (N_19518,N_19097,N_19341);
xor U19519 (N_19519,N_19421,N_19119);
and U19520 (N_19520,N_19485,N_19440);
nor U19521 (N_19521,N_19443,N_19147);
or U19522 (N_19522,N_19072,N_19135);
nor U19523 (N_19523,N_19237,N_19038);
xor U19524 (N_19524,N_19412,N_19209);
xor U19525 (N_19525,N_19382,N_19403);
and U19526 (N_19526,N_19073,N_19251);
or U19527 (N_19527,N_19286,N_19360);
and U19528 (N_19528,N_19013,N_19109);
or U19529 (N_19529,N_19215,N_19471);
xor U19530 (N_19530,N_19310,N_19491);
or U19531 (N_19531,N_19110,N_19088);
or U19532 (N_19532,N_19445,N_19002);
and U19533 (N_19533,N_19264,N_19302);
xnor U19534 (N_19534,N_19108,N_19056);
or U19535 (N_19535,N_19374,N_19256);
nor U19536 (N_19536,N_19340,N_19337);
and U19537 (N_19537,N_19091,N_19344);
nand U19538 (N_19538,N_19446,N_19395);
or U19539 (N_19539,N_19462,N_19419);
xnor U19540 (N_19540,N_19339,N_19441);
nor U19541 (N_19541,N_19007,N_19361);
nand U19542 (N_19542,N_19173,N_19390);
nor U19543 (N_19543,N_19265,N_19333);
nor U19544 (N_19544,N_19188,N_19164);
or U19545 (N_19545,N_19036,N_19058);
and U19546 (N_19546,N_19354,N_19185);
nor U19547 (N_19547,N_19044,N_19100);
nor U19548 (N_19548,N_19418,N_19414);
nand U19549 (N_19549,N_19363,N_19211);
xor U19550 (N_19550,N_19325,N_19282);
xnor U19551 (N_19551,N_19121,N_19127);
and U19552 (N_19552,N_19432,N_19045);
or U19553 (N_19553,N_19204,N_19153);
or U19554 (N_19554,N_19423,N_19208);
or U19555 (N_19555,N_19317,N_19150);
nand U19556 (N_19556,N_19186,N_19331);
xnor U19557 (N_19557,N_19125,N_19004);
or U19558 (N_19558,N_19272,N_19247);
nand U19559 (N_19559,N_19404,N_19010);
nand U19560 (N_19560,N_19483,N_19379);
or U19561 (N_19561,N_19285,N_19296);
and U19562 (N_19562,N_19156,N_19218);
or U19563 (N_19563,N_19328,N_19187);
xnor U19564 (N_19564,N_19378,N_19026);
or U19565 (N_19565,N_19053,N_19242);
and U19566 (N_19566,N_19311,N_19452);
nand U19567 (N_19567,N_19233,N_19112);
xnor U19568 (N_19568,N_19380,N_19131);
or U19569 (N_19569,N_19235,N_19323);
nand U19570 (N_19570,N_19267,N_19435);
xor U19571 (N_19571,N_19466,N_19142);
xnor U19572 (N_19572,N_19075,N_19065);
and U19573 (N_19573,N_19025,N_19394);
nand U19574 (N_19574,N_19154,N_19298);
and U19575 (N_19575,N_19236,N_19230);
nand U19576 (N_19576,N_19175,N_19133);
xnor U19577 (N_19577,N_19258,N_19301);
and U19578 (N_19578,N_19292,N_19043);
or U19579 (N_19579,N_19226,N_19113);
nor U19580 (N_19580,N_19227,N_19278);
or U19581 (N_19581,N_19303,N_19397);
nor U19582 (N_19582,N_19406,N_19312);
nand U19583 (N_19583,N_19129,N_19136);
or U19584 (N_19584,N_19478,N_19063);
and U19585 (N_19585,N_19261,N_19146);
xnor U19586 (N_19586,N_19409,N_19308);
or U19587 (N_19587,N_19366,N_19243);
nand U19588 (N_19588,N_19476,N_19239);
nand U19589 (N_19589,N_19262,N_19259);
nor U19590 (N_19590,N_19207,N_19284);
nor U19591 (N_19591,N_19138,N_19212);
and U19592 (N_19592,N_19266,N_19117);
nor U19593 (N_19593,N_19269,N_19047);
or U19594 (N_19594,N_19181,N_19196);
nand U19595 (N_19595,N_19094,N_19042);
and U19596 (N_19596,N_19442,N_19324);
nor U19597 (N_19597,N_19155,N_19407);
or U19598 (N_19598,N_19455,N_19015);
nand U19599 (N_19599,N_19068,N_19376);
nor U19600 (N_19600,N_19429,N_19371);
nor U19601 (N_19601,N_19123,N_19430);
xor U19602 (N_19602,N_19297,N_19077);
or U19603 (N_19603,N_19143,N_19335);
or U19604 (N_19604,N_19448,N_19456);
or U19605 (N_19605,N_19046,N_19049);
nand U19606 (N_19606,N_19161,N_19271);
nor U19607 (N_19607,N_19062,N_19465);
or U19608 (N_19608,N_19257,N_19014);
nor U19609 (N_19609,N_19149,N_19070);
nor U19610 (N_19610,N_19373,N_19064);
nor U19611 (N_19611,N_19289,N_19336);
or U19612 (N_19612,N_19051,N_19166);
nor U19613 (N_19613,N_19497,N_19249);
and U19614 (N_19614,N_19248,N_19330);
or U19615 (N_19615,N_19022,N_19030);
and U19616 (N_19616,N_19069,N_19048);
nor U19617 (N_19617,N_19176,N_19089);
and U19618 (N_19618,N_19370,N_19194);
xor U19619 (N_19619,N_19385,N_19221);
nor U19620 (N_19620,N_19451,N_19334);
nor U19621 (N_19621,N_19329,N_19454);
or U19622 (N_19622,N_19294,N_19021);
nand U19623 (N_19623,N_19486,N_19314);
nor U19624 (N_19624,N_19061,N_19383);
and U19625 (N_19625,N_19052,N_19120);
or U19626 (N_19626,N_19319,N_19316);
or U19627 (N_19627,N_19126,N_19306);
nor U19628 (N_19628,N_19229,N_19377);
or U19629 (N_19629,N_19169,N_19343);
and U19630 (N_19630,N_19040,N_19253);
or U19631 (N_19631,N_19422,N_19162);
and U19632 (N_19632,N_19232,N_19463);
xnor U19633 (N_19633,N_19420,N_19160);
and U19634 (N_19634,N_19305,N_19224);
nor U19635 (N_19635,N_19205,N_19411);
xnor U19636 (N_19636,N_19368,N_19299);
nand U19637 (N_19637,N_19413,N_19480);
nand U19638 (N_19638,N_19074,N_19487);
nor U19639 (N_19639,N_19114,N_19436);
or U19640 (N_19640,N_19009,N_19364);
and U19641 (N_19641,N_19493,N_19039);
nand U19642 (N_19642,N_19392,N_19148);
nor U19643 (N_19643,N_19193,N_19165);
nand U19644 (N_19644,N_19000,N_19355);
or U19645 (N_19645,N_19460,N_19349);
nand U19646 (N_19646,N_19273,N_19450);
nor U19647 (N_19647,N_19059,N_19198);
nand U19648 (N_19648,N_19434,N_19482);
or U19649 (N_19649,N_19470,N_19079);
xor U19650 (N_19650,N_19203,N_19287);
nand U19651 (N_19651,N_19191,N_19346);
nand U19652 (N_19652,N_19159,N_19172);
xor U19653 (N_19653,N_19473,N_19467);
nor U19654 (N_19654,N_19228,N_19122);
xnor U19655 (N_19655,N_19220,N_19260);
nor U19656 (N_19656,N_19495,N_19246);
xnor U19657 (N_19657,N_19137,N_19281);
or U19658 (N_19658,N_19342,N_19178);
or U19659 (N_19659,N_19037,N_19050);
nand U19660 (N_19660,N_19358,N_19274);
nand U19661 (N_19661,N_19288,N_19291);
nand U19662 (N_19662,N_19141,N_19268);
xnor U19663 (N_19663,N_19105,N_19494);
xnor U19664 (N_19664,N_19399,N_19111);
nand U19665 (N_19665,N_19029,N_19098);
xor U19666 (N_19666,N_19469,N_19213);
xor U19667 (N_19667,N_19332,N_19152);
and U19668 (N_19668,N_19101,N_19096);
or U19669 (N_19669,N_19279,N_19372);
nor U19670 (N_19670,N_19200,N_19365);
or U19671 (N_19671,N_19398,N_19118);
xnor U19672 (N_19672,N_19477,N_19225);
nor U19673 (N_19673,N_19167,N_19457);
or U19674 (N_19674,N_19490,N_19367);
nor U19675 (N_19675,N_19234,N_19318);
or U19676 (N_19676,N_19087,N_19402);
or U19677 (N_19677,N_19263,N_19484);
and U19678 (N_19678,N_19369,N_19060);
xnor U19679 (N_19679,N_19090,N_19067);
xnor U19680 (N_19680,N_19499,N_19307);
xnor U19681 (N_19681,N_19081,N_19086);
nor U19682 (N_19682,N_19084,N_19240);
or U19683 (N_19683,N_19359,N_19275);
nor U19684 (N_19684,N_19351,N_19439);
xor U19685 (N_19685,N_19132,N_19458);
xnor U19686 (N_19686,N_19405,N_19199);
or U19687 (N_19687,N_19177,N_19309);
xnor U19688 (N_19688,N_19400,N_19348);
nand U19689 (N_19689,N_19417,N_19016);
xnor U19690 (N_19690,N_19254,N_19444);
xor U19691 (N_19691,N_19214,N_19028);
and U19692 (N_19692,N_19145,N_19158);
and U19693 (N_19693,N_19217,N_19427);
or U19694 (N_19694,N_19391,N_19171);
nand U19695 (N_19695,N_19066,N_19017);
xor U19696 (N_19696,N_19174,N_19280);
and U19697 (N_19697,N_19431,N_19080);
xnor U19698 (N_19698,N_19447,N_19362);
and U19699 (N_19699,N_19252,N_19461);
nor U19700 (N_19700,N_19023,N_19350);
and U19701 (N_19701,N_19464,N_19018);
and U19702 (N_19702,N_19003,N_19475);
nor U19703 (N_19703,N_19216,N_19300);
xor U19704 (N_19704,N_19496,N_19353);
nand U19705 (N_19705,N_19433,N_19180);
nor U19706 (N_19706,N_19315,N_19322);
xnor U19707 (N_19707,N_19093,N_19345);
nand U19708 (N_19708,N_19425,N_19438);
xor U19709 (N_19709,N_19250,N_19115);
nor U19710 (N_19710,N_19347,N_19019);
nand U19711 (N_19711,N_19277,N_19387);
nand U19712 (N_19712,N_19124,N_19190);
xnor U19713 (N_19713,N_19005,N_19386);
nand U19714 (N_19714,N_19116,N_19130);
or U19715 (N_19715,N_19415,N_19276);
nor U19716 (N_19716,N_19083,N_19459);
xnor U19717 (N_19717,N_19192,N_19408);
nand U19718 (N_19718,N_19356,N_19184);
or U19719 (N_19719,N_19492,N_19270);
or U19720 (N_19720,N_19313,N_19011);
or U19721 (N_19721,N_19197,N_19201);
xnor U19722 (N_19722,N_19027,N_19338);
or U19723 (N_19723,N_19170,N_19006);
nand U19724 (N_19724,N_19352,N_19290);
or U19725 (N_19725,N_19384,N_19103);
or U19726 (N_19726,N_19099,N_19055);
and U19727 (N_19727,N_19424,N_19396);
nand U19728 (N_19728,N_19231,N_19401);
nor U19729 (N_19729,N_19223,N_19295);
nand U19730 (N_19730,N_19393,N_19092);
nor U19731 (N_19731,N_19032,N_19182);
and U19732 (N_19732,N_19481,N_19078);
xnor U19733 (N_19733,N_19076,N_19321);
or U19734 (N_19734,N_19389,N_19304);
and U19735 (N_19735,N_19479,N_19255);
xnor U19736 (N_19736,N_19189,N_19140);
xor U19737 (N_19737,N_19095,N_19179);
nor U19738 (N_19738,N_19357,N_19472);
or U19739 (N_19739,N_19106,N_19104);
nor U19740 (N_19740,N_19012,N_19085);
nor U19741 (N_19741,N_19041,N_19381);
nand U19742 (N_19742,N_19144,N_19202);
and U19743 (N_19743,N_19128,N_19474);
nand U19744 (N_19744,N_19238,N_19107);
xor U19745 (N_19745,N_19024,N_19437);
nor U19746 (N_19746,N_19035,N_19320);
or U19747 (N_19747,N_19244,N_19054);
or U19748 (N_19748,N_19020,N_19426);
xor U19749 (N_19749,N_19453,N_19498);
nand U19750 (N_19750,N_19428,N_19311);
and U19751 (N_19751,N_19093,N_19485);
nor U19752 (N_19752,N_19034,N_19260);
nand U19753 (N_19753,N_19173,N_19152);
xor U19754 (N_19754,N_19311,N_19198);
nand U19755 (N_19755,N_19318,N_19385);
or U19756 (N_19756,N_19323,N_19262);
or U19757 (N_19757,N_19356,N_19375);
or U19758 (N_19758,N_19089,N_19302);
nor U19759 (N_19759,N_19373,N_19043);
and U19760 (N_19760,N_19044,N_19102);
and U19761 (N_19761,N_19401,N_19281);
or U19762 (N_19762,N_19032,N_19210);
xor U19763 (N_19763,N_19422,N_19171);
or U19764 (N_19764,N_19048,N_19171);
or U19765 (N_19765,N_19269,N_19090);
xnor U19766 (N_19766,N_19330,N_19433);
and U19767 (N_19767,N_19123,N_19044);
and U19768 (N_19768,N_19373,N_19140);
nand U19769 (N_19769,N_19316,N_19352);
nand U19770 (N_19770,N_19387,N_19268);
nor U19771 (N_19771,N_19105,N_19347);
nor U19772 (N_19772,N_19312,N_19091);
or U19773 (N_19773,N_19000,N_19492);
nand U19774 (N_19774,N_19006,N_19091);
or U19775 (N_19775,N_19223,N_19377);
nor U19776 (N_19776,N_19004,N_19449);
nor U19777 (N_19777,N_19431,N_19489);
and U19778 (N_19778,N_19409,N_19481);
nor U19779 (N_19779,N_19463,N_19166);
nand U19780 (N_19780,N_19191,N_19277);
nand U19781 (N_19781,N_19035,N_19326);
nand U19782 (N_19782,N_19349,N_19144);
xnor U19783 (N_19783,N_19117,N_19328);
or U19784 (N_19784,N_19438,N_19230);
and U19785 (N_19785,N_19077,N_19170);
nor U19786 (N_19786,N_19255,N_19146);
nor U19787 (N_19787,N_19027,N_19267);
nor U19788 (N_19788,N_19335,N_19157);
xor U19789 (N_19789,N_19276,N_19357);
or U19790 (N_19790,N_19164,N_19472);
or U19791 (N_19791,N_19463,N_19302);
nor U19792 (N_19792,N_19176,N_19058);
xor U19793 (N_19793,N_19305,N_19240);
and U19794 (N_19794,N_19167,N_19324);
xor U19795 (N_19795,N_19127,N_19445);
and U19796 (N_19796,N_19070,N_19388);
nand U19797 (N_19797,N_19445,N_19379);
and U19798 (N_19798,N_19015,N_19155);
and U19799 (N_19799,N_19280,N_19033);
and U19800 (N_19800,N_19463,N_19235);
and U19801 (N_19801,N_19174,N_19385);
or U19802 (N_19802,N_19004,N_19188);
nand U19803 (N_19803,N_19069,N_19374);
or U19804 (N_19804,N_19257,N_19378);
or U19805 (N_19805,N_19352,N_19132);
nor U19806 (N_19806,N_19225,N_19284);
nor U19807 (N_19807,N_19060,N_19276);
nand U19808 (N_19808,N_19235,N_19044);
or U19809 (N_19809,N_19472,N_19108);
nand U19810 (N_19810,N_19051,N_19354);
or U19811 (N_19811,N_19291,N_19419);
and U19812 (N_19812,N_19474,N_19074);
xor U19813 (N_19813,N_19081,N_19004);
nor U19814 (N_19814,N_19378,N_19260);
xor U19815 (N_19815,N_19306,N_19090);
or U19816 (N_19816,N_19139,N_19468);
and U19817 (N_19817,N_19448,N_19148);
and U19818 (N_19818,N_19015,N_19405);
nand U19819 (N_19819,N_19033,N_19383);
xor U19820 (N_19820,N_19163,N_19069);
nand U19821 (N_19821,N_19213,N_19319);
nor U19822 (N_19822,N_19213,N_19286);
nor U19823 (N_19823,N_19226,N_19181);
xnor U19824 (N_19824,N_19262,N_19253);
nand U19825 (N_19825,N_19269,N_19391);
nor U19826 (N_19826,N_19095,N_19167);
and U19827 (N_19827,N_19170,N_19207);
nand U19828 (N_19828,N_19028,N_19373);
and U19829 (N_19829,N_19356,N_19498);
nor U19830 (N_19830,N_19004,N_19126);
and U19831 (N_19831,N_19232,N_19256);
nor U19832 (N_19832,N_19112,N_19011);
nand U19833 (N_19833,N_19416,N_19478);
or U19834 (N_19834,N_19144,N_19142);
or U19835 (N_19835,N_19029,N_19178);
and U19836 (N_19836,N_19438,N_19109);
nor U19837 (N_19837,N_19232,N_19107);
or U19838 (N_19838,N_19284,N_19078);
and U19839 (N_19839,N_19061,N_19241);
xor U19840 (N_19840,N_19325,N_19372);
and U19841 (N_19841,N_19084,N_19483);
or U19842 (N_19842,N_19459,N_19361);
xnor U19843 (N_19843,N_19372,N_19024);
nand U19844 (N_19844,N_19097,N_19184);
and U19845 (N_19845,N_19302,N_19497);
and U19846 (N_19846,N_19035,N_19120);
xor U19847 (N_19847,N_19484,N_19145);
xnor U19848 (N_19848,N_19080,N_19291);
nor U19849 (N_19849,N_19213,N_19177);
or U19850 (N_19850,N_19065,N_19042);
xor U19851 (N_19851,N_19241,N_19474);
nand U19852 (N_19852,N_19413,N_19338);
or U19853 (N_19853,N_19083,N_19444);
nand U19854 (N_19854,N_19093,N_19383);
or U19855 (N_19855,N_19269,N_19285);
and U19856 (N_19856,N_19453,N_19144);
nand U19857 (N_19857,N_19424,N_19301);
xor U19858 (N_19858,N_19152,N_19094);
and U19859 (N_19859,N_19101,N_19371);
or U19860 (N_19860,N_19006,N_19140);
nor U19861 (N_19861,N_19325,N_19109);
xor U19862 (N_19862,N_19227,N_19178);
or U19863 (N_19863,N_19063,N_19438);
or U19864 (N_19864,N_19378,N_19329);
nor U19865 (N_19865,N_19232,N_19335);
or U19866 (N_19866,N_19413,N_19201);
xnor U19867 (N_19867,N_19232,N_19350);
nand U19868 (N_19868,N_19218,N_19382);
and U19869 (N_19869,N_19295,N_19250);
or U19870 (N_19870,N_19061,N_19086);
xnor U19871 (N_19871,N_19388,N_19408);
nor U19872 (N_19872,N_19098,N_19386);
or U19873 (N_19873,N_19292,N_19045);
and U19874 (N_19874,N_19209,N_19418);
xor U19875 (N_19875,N_19256,N_19237);
or U19876 (N_19876,N_19365,N_19232);
nand U19877 (N_19877,N_19495,N_19155);
or U19878 (N_19878,N_19256,N_19123);
nor U19879 (N_19879,N_19191,N_19234);
and U19880 (N_19880,N_19112,N_19360);
and U19881 (N_19881,N_19084,N_19017);
nand U19882 (N_19882,N_19363,N_19122);
and U19883 (N_19883,N_19248,N_19352);
or U19884 (N_19884,N_19078,N_19322);
nor U19885 (N_19885,N_19026,N_19401);
or U19886 (N_19886,N_19041,N_19014);
and U19887 (N_19887,N_19321,N_19042);
nor U19888 (N_19888,N_19076,N_19364);
and U19889 (N_19889,N_19138,N_19405);
nand U19890 (N_19890,N_19120,N_19075);
nor U19891 (N_19891,N_19368,N_19430);
and U19892 (N_19892,N_19125,N_19210);
nand U19893 (N_19893,N_19185,N_19432);
nand U19894 (N_19894,N_19262,N_19006);
nand U19895 (N_19895,N_19330,N_19233);
nor U19896 (N_19896,N_19284,N_19406);
and U19897 (N_19897,N_19213,N_19253);
nor U19898 (N_19898,N_19170,N_19465);
and U19899 (N_19899,N_19175,N_19465);
and U19900 (N_19900,N_19218,N_19135);
xnor U19901 (N_19901,N_19032,N_19171);
or U19902 (N_19902,N_19349,N_19443);
and U19903 (N_19903,N_19291,N_19245);
or U19904 (N_19904,N_19311,N_19039);
xnor U19905 (N_19905,N_19347,N_19455);
and U19906 (N_19906,N_19039,N_19419);
and U19907 (N_19907,N_19271,N_19068);
or U19908 (N_19908,N_19333,N_19061);
nor U19909 (N_19909,N_19351,N_19272);
or U19910 (N_19910,N_19203,N_19401);
nor U19911 (N_19911,N_19427,N_19033);
xnor U19912 (N_19912,N_19062,N_19122);
nand U19913 (N_19913,N_19017,N_19150);
xor U19914 (N_19914,N_19191,N_19354);
xor U19915 (N_19915,N_19133,N_19193);
nor U19916 (N_19916,N_19296,N_19077);
or U19917 (N_19917,N_19127,N_19307);
xnor U19918 (N_19918,N_19006,N_19271);
nor U19919 (N_19919,N_19125,N_19464);
nand U19920 (N_19920,N_19031,N_19347);
nor U19921 (N_19921,N_19374,N_19075);
nand U19922 (N_19922,N_19096,N_19019);
nand U19923 (N_19923,N_19351,N_19278);
xnor U19924 (N_19924,N_19496,N_19323);
and U19925 (N_19925,N_19328,N_19497);
xor U19926 (N_19926,N_19322,N_19459);
and U19927 (N_19927,N_19121,N_19462);
or U19928 (N_19928,N_19486,N_19003);
nand U19929 (N_19929,N_19336,N_19027);
nor U19930 (N_19930,N_19128,N_19062);
and U19931 (N_19931,N_19169,N_19382);
nand U19932 (N_19932,N_19067,N_19343);
and U19933 (N_19933,N_19232,N_19043);
nand U19934 (N_19934,N_19125,N_19097);
nor U19935 (N_19935,N_19318,N_19188);
nand U19936 (N_19936,N_19361,N_19037);
or U19937 (N_19937,N_19122,N_19121);
xnor U19938 (N_19938,N_19107,N_19195);
and U19939 (N_19939,N_19293,N_19171);
nor U19940 (N_19940,N_19336,N_19400);
or U19941 (N_19941,N_19431,N_19121);
nor U19942 (N_19942,N_19110,N_19108);
and U19943 (N_19943,N_19358,N_19397);
nand U19944 (N_19944,N_19203,N_19105);
nand U19945 (N_19945,N_19159,N_19044);
nand U19946 (N_19946,N_19135,N_19077);
or U19947 (N_19947,N_19035,N_19367);
and U19948 (N_19948,N_19444,N_19482);
or U19949 (N_19949,N_19374,N_19231);
xor U19950 (N_19950,N_19329,N_19296);
nand U19951 (N_19951,N_19484,N_19035);
xnor U19952 (N_19952,N_19250,N_19288);
or U19953 (N_19953,N_19213,N_19188);
or U19954 (N_19954,N_19436,N_19457);
nand U19955 (N_19955,N_19087,N_19395);
xor U19956 (N_19956,N_19073,N_19293);
or U19957 (N_19957,N_19447,N_19309);
nand U19958 (N_19958,N_19017,N_19171);
and U19959 (N_19959,N_19209,N_19179);
or U19960 (N_19960,N_19478,N_19293);
nand U19961 (N_19961,N_19404,N_19485);
nand U19962 (N_19962,N_19245,N_19163);
xnor U19963 (N_19963,N_19372,N_19250);
and U19964 (N_19964,N_19432,N_19174);
nor U19965 (N_19965,N_19448,N_19310);
nor U19966 (N_19966,N_19002,N_19046);
and U19967 (N_19967,N_19266,N_19059);
or U19968 (N_19968,N_19024,N_19398);
xnor U19969 (N_19969,N_19211,N_19165);
xnor U19970 (N_19970,N_19422,N_19175);
or U19971 (N_19971,N_19143,N_19474);
xor U19972 (N_19972,N_19344,N_19007);
nor U19973 (N_19973,N_19485,N_19167);
and U19974 (N_19974,N_19429,N_19206);
nand U19975 (N_19975,N_19096,N_19458);
and U19976 (N_19976,N_19411,N_19029);
xnor U19977 (N_19977,N_19127,N_19400);
nor U19978 (N_19978,N_19090,N_19160);
xor U19979 (N_19979,N_19346,N_19018);
nor U19980 (N_19980,N_19379,N_19324);
xor U19981 (N_19981,N_19376,N_19244);
xnor U19982 (N_19982,N_19438,N_19163);
and U19983 (N_19983,N_19153,N_19216);
xnor U19984 (N_19984,N_19033,N_19195);
nor U19985 (N_19985,N_19426,N_19100);
xor U19986 (N_19986,N_19477,N_19481);
or U19987 (N_19987,N_19194,N_19372);
nor U19988 (N_19988,N_19138,N_19300);
nor U19989 (N_19989,N_19480,N_19408);
and U19990 (N_19990,N_19282,N_19090);
nor U19991 (N_19991,N_19133,N_19427);
nor U19992 (N_19992,N_19016,N_19047);
nor U19993 (N_19993,N_19443,N_19211);
and U19994 (N_19994,N_19251,N_19353);
xor U19995 (N_19995,N_19331,N_19044);
or U19996 (N_19996,N_19255,N_19211);
or U19997 (N_19997,N_19284,N_19402);
or U19998 (N_19998,N_19432,N_19238);
xor U19999 (N_19999,N_19332,N_19162);
nor U20000 (N_20000,N_19909,N_19624);
nand U20001 (N_20001,N_19816,N_19694);
xnor U20002 (N_20002,N_19794,N_19729);
nor U20003 (N_20003,N_19839,N_19769);
and U20004 (N_20004,N_19786,N_19539);
and U20005 (N_20005,N_19831,N_19675);
nand U20006 (N_20006,N_19500,N_19876);
nor U20007 (N_20007,N_19832,N_19900);
xor U20008 (N_20008,N_19751,N_19682);
or U20009 (N_20009,N_19978,N_19796);
nor U20010 (N_20010,N_19591,N_19771);
nor U20011 (N_20011,N_19578,N_19582);
or U20012 (N_20012,N_19757,N_19838);
nor U20013 (N_20013,N_19603,N_19532);
and U20014 (N_20014,N_19705,N_19898);
nand U20015 (N_20015,N_19570,N_19933);
and U20016 (N_20016,N_19560,N_19809);
nor U20017 (N_20017,N_19706,N_19897);
xnor U20018 (N_20018,N_19581,N_19674);
or U20019 (N_20019,N_19892,N_19995);
or U20020 (N_20020,N_19587,N_19653);
or U20021 (N_20021,N_19661,N_19529);
xor U20022 (N_20022,N_19584,N_19770);
or U20023 (N_20023,N_19704,N_19616);
or U20024 (N_20024,N_19689,N_19760);
nor U20025 (N_20025,N_19501,N_19576);
xor U20026 (N_20026,N_19976,N_19505);
or U20027 (N_20027,N_19939,N_19709);
nor U20028 (N_20028,N_19609,N_19556);
nor U20029 (N_20029,N_19620,N_19766);
nand U20030 (N_20030,N_19647,N_19993);
xor U20031 (N_20031,N_19519,N_19716);
nor U20032 (N_20032,N_19802,N_19657);
xor U20033 (N_20033,N_19905,N_19652);
nand U20034 (N_20034,N_19807,N_19827);
nor U20035 (N_20035,N_19793,N_19861);
nand U20036 (N_20036,N_19670,N_19684);
nand U20037 (N_20037,N_19872,N_19859);
nand U20038 (N_20038,N_19640,N_19884);
and U20039 (N_20039,N_19602,N_19799);
nand U20040 (N_20040,N_19561,N_19812);
xnor U20041 (N_20041,N_19690,N_19870);
nor U20042 (N_20042,N_19969,N_19946);
xnor U20043 (N_20043,N_19862,N_19922);
or U20044 (N_20044,N_19540,N_19887);
or U20045 (N_20045,N_19901,N_19753);
nor U20046 (N_20046,N_19719,N_19549);
or U20047 (N_20047,N_19542,N_19818);
nor U20048 (N_20048,N_19878,N_19881);
nor U20049 (N_20049,N_19586,N_19658);
xnor U20050 (N_20050,N_19625,N_19509);
nand U20051 (N_20051,N_19655,N_19554);
and U20052 (N_20052,N_19575,N_19747);
and U20053 (N_20053,N_19646,N_19514);
or U20054 (N_20054,N_19994,N_19511);
xor U20055 (N_20055,N_19848,N_19502);
nor U20056 (N_20056,N_19685,N_19913);
or U20057 (N_20057,N_19768,N_19999);
or U20058 (N_20058,N_19547,N_19621);
nand U20059 (N_20059,N_19804,N_19577);
or U20060 (N_20060,N_19643,N_19672);
and U20061 (N_20061,N_19638,N_19918);
nor U20062 (N_20062,N_19541,N_19951);
nand U20063 (N_20063,N_19808,N_19854);
nor U20064 (N_20064,N_19671,N_19772);
nor U20065 (N_20065,N_19846,N_19977);
xnor U20066 (N_20066,N_19960,N_19991);
and U20067 (N_20067,N_19911,N_19545);
nor U20068 (N_20068,N_19619,N_19851);
xnor U20069 (N_20069,N_19571,N_19798);
nor U20070 (N_20070,N_19527,N_19773);
and U20071 (N_20071,N_19943,N_19886);
or U20072 (N_20072,N_19622,N_19633);
nand U20073 (N_20073,N_19656,N_19522);
nor U20074 (N_20074,N_19654,N_19634);
and U20075 (N_20075,N_19593,N_19718);
nor U20076 (N_20076,N_19610,N_19919);
xnor U20077 (N_20077,N_19728,N_19681);
nand U20078 (N_20078,N_19596,N_19907);
nor U20079 (N_20079,N_19789,N_19845);
nand U20080 (N_20080,N_19597,N_19936);
xor U20081 (N_20081,N_19651,N_19820);
or U20082 (N_20082,N_19612,N_19930);
and U20083 (N_20083,N_19662,N_19598);
nor U20084 (N_20084,N_19917,N_19959);
and U20085 (N_20085,N_19756,N_19929);
and U20086 (N_20086,N_19567,N_19844);
or U20087 (N_20087,N_19923,N_19693);
nand U20088 (N_20088,N_19891,N_19528);
xnor U20089 (N_20089,N_19955,N_19781);
xnor U20090 (N_20090,N_19776,N_19692);
nor U20091 (N_20091,N_19623,N_19592);
or U20092 (N_20092,N_19941,N_19686);
nor U20093 (N_20093,N_19710,N_19890);
or U20094 (N_20094,N_19687,N_19821);
and U20095 (N_20095,N_19664,N_19665);
nor U20096 (N_20096,N_19834,N_19795);
xnor U20097 (N_20097,N_19660,N_19937);
and U20098 (N_20098,N_19695,N_19608);
and U20099 (N_20099,N_19703,N_19927);
or U20100 (N_20100,N_19948,N_19516);
nor U20101 (N_20101,N_19644,N_19715);
xor U20102 (N_20102,N_19910,N_19850);
xnor U20103 (N_20103,N_19828,N_19521);
and U20104 (N_20104,N_19722,N_19889);
nor U20105 (N_20105,N_19618,N_19787);
nor U20106 (N_20106,N_19829,N_19860);
and U20107 (N_20107,N_19996,N_19797);
or U20108 (N_20108,N_19589,N_19894);
xor U20109 (N_20109,N_19968,N_19880);
or U20110 (N_20110,N_19750,N_19548);
nor U20111 (N_20111,N_19855,N_19814);
nor U20112 (N_20112,N_19767,N_19611);
or U20113 (N_20113,N_19680,N_19600);
xor U20114 (N_20114,N_19701,N_19510);
xnor U20115 (N_20115,N_19924,N_19720);
nor U20116 (N_20116,N_19835,N_19815);
and U20117 (N_20117,N_19906,N_19688);
or U20118 (N_20118,N_19746,N_19745);
and U20119 (N_20119,N_19883,N_19761);
and U20120 (N_20120,N_19607,N_19678);
and U20121 (N_20121,N_19920,N_19819);
xnor U20122 (N_20122,N_19824,N_19931);
xnor U20123 (N_20123,N_19895,N_19837);
or U20124 (N_20124,N_19817,N_19735);
and U20125 (N_20125,N_19712,N_19732);
nand U20126 (N_20126,N_19559,N_19962);
nor U20127 (N_20127,N_19974,N_19721);
nand U20128 (N_20128,N_19617,N_19741);
xnor U20129 (N_20129,N_19928,N_19806);
nor U20130 (N_20130,N_19744,N_19988);
xor U20131 (N_20131,N_19533,N_19736);
nand U20132 (N_20132,N_19515,N_19949);
nor U20133 (N_20133,N_19507,N_19588);
xor U20134 (N_20134,N_19950,N_19535);
or U20135 (N_20135,N_19879,N_19667);
xor U20136 (N_20136,N_19520,N_19604);
or U20137 (N_20137,N_19967,N_19723);
nor U20138 (N_20138,N_19983,N_19645);
and U20139 (N_20139,N_19800,N_19724);
and U20140 (N_20140,N_19987,N_19963);
xnor U20141 (N_20141,N_19626,N_19572);
and U20142 (N_20142,N_19964,N_19822);
xnor U20143 (N_20143,N_19961,N_19874);
and U20144 (N_20144,N_19863,N_19537);
nor U20145 (N_20145,N_19659,N_19777);
and U20146 (N_20146,N_19873,N_19754);
nand U20147 (N_20147,N_19606,N_19613);
or U20148 (N_20148,N_19546,N_19649);
and U20149 (N_20149,N_19912,N_19614);
and U20150 (N_20150,N_19975,N_19915);
nor U20151 (N_20151,N_19791,N_19632);
nor U20152 (N_20152,N_19893,N_19574);
and U20153 (N_20153,N_19877,N_19811);
nand U20154 (N_20154,N_19737,N_19984);
nand U20155 (N_20155,N_19849,N_19708);
nor U20156 (N_20156,N_19641,N_19785);
or U20157 (N_20157,N_19508,N_19595);
nor U20158 (N_20158,N_19947,N_19934);
and U20159 (N_20159,N_19957,N_19569);
xor U20160 (N_20160,N_19579,N_19568);
nand U20161 (N_20161,N_19666,N_19982);
nor U20162 (N_20162,N_19759,N_19629);
nand U20163 (N_20163,N_19864,N_19774);
nor U20164 (N_20164,N_19601,N_19573);
or U20165 (N_20165,N_19740,N_19833);
xor U20166 (N_20166,N_19858,N_19525);
or U20167 (N_20167,N_19867,N_19717);
and U20168 (N_20168,N_19538,N_19702);
nand U20169 (N_20169,N_19630,N_19635);
nor U20170 (N_20170,N_19564,N_19944);
and U20171 (N_20171,N_19868,N_19531);
xnor U20172 (N_20172,N_19792,N_19902);
nor U20173 (N_20173,N_19707,N_19973);
xor U20174 (N_20174,N_19990,N_19734);
nor U20175 (N_20175,N_19783,N_19557);
or U20176 (N_20176,N_19903,N_19544);
nor U20177 (N_20177,N_19826,N_19758);
or U20178 (N_20178,N_19605,N_19823);
and U20179 (N_20179,N_19932,N_19550);
nand U20180 (N_20180,N_19669,N_19765);
and U20181 (N_20181,N_19752,N_19841);
nor U20182 (N_20182,N_19954,N_19530);
xor U20183 (N_20183,N_19583,N_19875);
and U20184 (N_20184,N_19790,N_19524);
xor U20185 (N_20185,N_19840,N_19739);
and U20186 (N_20186,N_19697,N_19989);
nor U20187 (N_20187,N_19585,N_19857);
nor U20188 (N_20188,N_19642,N_19513);
and U20189 (N_20189,N_19801,N_19566);
xor U20190 (N_20190,N_19726,N_19518);
or U20191 (N_20191,N_19725,N_19504);
and U20192 (N_20192,N_19896,N_19805);
or U20193 (N_20193,N_19942,N_19971);
nand U20194 (N_20194,N_19594,N_19981);
nor U20195 (N_20195,N_19637,N_19972);
nand U20196 (N_20196,N_19700,N_19782);
and U20197 (N_20197,N_19985,N_19553);
xor U20198 (N_20198,N_19997,N_19925);
or U20199 (N_20199,N_19543,N_19885);
nand U20200 (N_20200,N_19580,N_19749);
or U20201 (N_20201,N_19940,N_19506);
xnor U20202 (N_20202,N_19888,N_19953);
nand U20203 (N_20203,N_19558,N_19788);
and U20204 (N_20204,N_19679,N_19599);
or U20205 (N_20205,N_19945,N_19738);
nand U20206 (N_20206,N_19866,N_19778);
xnor U20207 (N_20207,N_19908,N_19551);
xor U20208 (N_20208,N_19965,N_19748);
xnor U20209 (N_20209,N_19730,N_19810);
nand U20210 (N_20210,N_19763,N_19636);
nor U20211 (N_20211,N_19631,N_19847);
nor U20212 (N_20212,N_19628,N_19836);
nand U20213 (N_20213,N_19779,N_19935);
nor U20214 (N_20214,N_19565,N_19865);
nor U20215 (N_20215,N_19762,N_19825);
nand U20216 (N_20216,N_19882,N_19727);
or U20217 (N_20217,N_19552,N_19813);
nor U20218 (N_20218,N_19986,N_19938);
xor U20219 (N_20219,N_19843,N_19650);
xnor U20220 (N_20220,N_19830,N_19916);
or U20221 (N_20221,N_19711,N_19966);
nor U20222 (N_20222,N_19523,N_19956);
xor U20223 (N_20223,N_19517,N_19713);
nand U20224 (N_20224,N_19926,N_19733);
or U20225 (N_20225,N_19696,N_19714);
and U20226 (N_20226,N_19555,N_19503);
or U20227 (N_20227,N_19755,N_19803);
or U20228 (N_20228,N_19698,N_19899);
nor U20229 (N_20229,N_19784,N_19871);
nor U20230 (N_20230,N_19677,N_19869);
and U20231 (N_20231,N_19980,N_19699);
or U20232 (N_20232,N_19526,N_19663);
nor U20233 (N_20233,N_19615,N_19731);
nand U20234 (N_20234,N_19780,N_19998);
or U20235 (N_20235,N_19852,N_19764);
nand U20236 (N_20236,N_19921,N_19673);
and U20237 (N_20237,N_19992,N_19563);
nor U20238 (N_20238,N_19952,N_19691);
nor U20239 (N_20239,N_19590,N_19958);
nand U20240 (N_20240,N_19683,N_19914);
or U20241 (N_20241,N_19775,N_19853);
xnor U20242 (N_20242,N_19534,N_19512);
xnor U20243 (N_20243,N_19676,N_19639);
xnor U20244 (N_20244,N_19904,N_19648);
nand U20245 (N_20245,N_19742,N_19562);
nand U20246 (N_20246,N_19856,N_19970);
nor U20247 (N_20247,N_19979,N_19627);
and U20248 (N_20248,N_19668,N_19536);
nor U20249 (N_20249,N_19842,N_19743);
and U20250 (N_20250,N_19983,N_19540);
nand U20251 (N_20251,N_19769,N_19868);
or U20252 (N_20252,N_19782,N_19536);
nand U20253 (N_20253,N_19899,N_19934);
and U20254 (N_20254,N_19932,N_19666);
xnor U20255 (N_20255,N_19780,N_19891);
nor U20256 (N_20256,N_19843,N_19774);
nor U20257 (N_20257,N_19575,N_19613);
nor U20258 (N_20258,N_19633,N_19742);
nor U20259 (N_20259,N_19613,N_19717);
and U20260 (N_20260,N_19909,N_19906);
xor U20261 (N_20261,N_19862,N_19760);
and U20262 (N_20262,N_19759,N_19893);
and U20263 (N_20263,N_19639,N_19898);
or U20264 (N_20264,N_19512,N_19716);
or U20265 (N_20265,N_19742,N_19761);
nand U20266 (N_20266,N_19527,N_19592);
nand U20267 (N_20267,N_19903,N_19825);
nand U20268 (N_20268,N_19609,N_19770);
nand U20269 (N_20269,N_19565,N_19667);
nand U20270 (N_20270,N_19629,N_19583);
and U20271 (N_20271,N_19628,N_19770);
nand U20272 (N_20272,N_19926,N_19734);
and U20273 (N_20273,N_19804,N_19830);
and U20274 (N_20274,N_19886,N_19570);
nand U20275 (N_20275,N_19723,N_19605);
and U20276 (N_20276,N_19671,N_19686);
or U20277 (N_20277,N_19650,N_19764);
xnor U20278 (N_20278,N_19562,N_19991);
and U20279 (N_20279,N_19807,N_19626);
or U20280 (N_20280,N_19909,N_19913);
and U20281 (N_20281,N_19875,N_19908);
and U20282 (N_20282,N_19942,N_19691);
xor U20283 (N_20283,N_19623,N_19859);
and U20284 (N_20284,N_19871,N_19540);
nand U20285 (N_20285,N_19653,N_19658);
and U20286 (N_20286,N_19609,N_19790);
xor U20287 (N_20287,N_19898,N_19973);
or U20288 (N_20288,N_19605,N_19592);
xnor U20289 (N_20289,N_19970,N_19881);
nor U20290 (N_20290,N_19717,N_19773);
nor U20291 (N_20291,N_19624,N_19821);
nand U20292 (N_20292,N_19509,N_19952);
and U20293 (N_20293,N_19567,N_19668);
nand U20294 (N_20294,N_19562,N_19709);
nand U20295 (N_20295,N_19894,N_19936);
nor U20296 (N_20296,N_19609,N_19798);
or U20297 (N_20297,N_19623,N_19885);
or U20298 (N_20298,N_19676,N_19548);
nand U20299 (N_20299,N_19819,N_19653);
nor U20300 (N_20300,N_19713,N_19786);
or U20301 (N_20301,N_19830,N_19611);
and U20302 (N_20302,N_19746,N_19676);
nor U20303 (N_20303,N_19524,N_19780);
xor U20304 (N_20304,N_19948,N_19825);
xnor U20305 (N_20305,N_19668,N_19947);
nand U20306 (N_20306,N_19812,N_19927);
xor U20307 (N_20307,N_19768,N_19706);
or U20308 (N_20308,N_19963,N_19794);
xor U20309 (N_20309,N_19948,N_19849);
xnor U20310 (N_20310,N_19740,N_19511);
nor U20311 (N_20311,N_19910,N_19830);
or U20312 (N_20312,N_19517,N_19752);
xnor U20313 (N_20313,N_19560,N_19774);
and U20314 (N_20314,N_19652,N_19821);
or U20315 (N_20315,N_19676,N_19641);
nand U20316 (N_20316,N_19735,N_19833);
and U20317 (N_20317,N_19765,N_19605);
and U20318 (N_20318,N_19802,N_19760);
or U20319 (N_20319,N_19847,N_19750);
nand U20320 (N_20320,N_19987,N_19930);
nor U20321 (N_20321,N_19960,N_19967);
and U20322 (N_20322,N_19786,N_19984);
nand U20323 (N_20323,N_19527,N_19643);
nor U20324 (N_20324,N_19770,N_19831);
and U20325 (N_20325,N_19642,N_19719);
nor U20326 (N_20326,N_19899,N_19838);
xnor U20327 (N_20327,N_19633,N_19732);
and U20328 (N_20328,N_19736,N_19925);
nand U20329 (N_20329,N_19602,N_19752);
xnor U20330 (N_20330,N_19887,N_19534);
xor U20331 (N_20331,N_19859,N_19735);
nor U20332 (N_20332,N_19867,N_19911);
nor U20333 (N_20333,N_19671,N_19599);
nand U20334 (N_20334,N_19514,N_19506);
xnor U20335 (N_20335,N_19547,N_19719);
xnor U20336 (N_20336,N_19661,N_19549);
and U20337 (N_20337,N_19850,N_19711);
nor U20338 (N_20338,N_19677,N_19872);
or U20339 (N_20339,N_19518,N_19822);
nand U20340 (N_20340,N_19884,N_19837);
and U20341 (N_20341,N_19606,N_19736);
or U20342 (N_20342,N_19999,N_19733);
and U20343 (N_20343,N_19592,N_19704);
xor U20344 (N_20344,N_19704,N_19932);
or U20345 (N_20345,N_19696,N_19818);
or U20346 (N_20346,N_19639,N_19642);
nor U20347 (N_20347,N_19637,N_19708);
xor U20348 (N_20348,N_19558,N_19950);
xor U20349 (N_20349,N_19584,N_19540);
xor U20350 (N_20350,N_19570,N_19895);
nand U20351 (N_20351,N_19671,N_19709);
and U20352 (N_20352,N_19594,N_19891);
nand U20353 (N_20353,N_19918,N_19749);
or U20354 (N_20354,N_19956,N_19538);
or U20355 (N_20355,N_19887,N_19615);
xor U20356 (N_20356,N_19635,N_19751);
xor U20357 (N_20357,N_19942,N_19576);
or U20358 (N_20358,N_19537,N_19890);
xnor U20359 (N_20359,N_19647,N_19518);
or U20360 (N_20360,N_19675,N_19945);
and U20361 (N_20361,N_19736,N_19752);
and U20362 (N_20362,N_19558,N_19870);
and U20363 (N_20363,N_19922,N_19639);
xor U20364 (N_20364,N_19506,N_19597);
xnor U20365 (N_20365,N_19842,N_19813);
nand U20366 (N_20366,N_19740,N_19771);
nand U20367 (N_20367,N_19795,N_19700);
nor U20368 (N_20368,N_19626,N_19976);
nand U20369 (N_20369,N_19561,N_19696);
and U20370 (N_20370,N_19994,N_19663);
and U20371 (N_20371,N_19527,N_19582);
nand U20372 (N_20372,N_19950,N_19812);
nand U20373 (N_20373,N_19885,N_19622);
nor U20374 (N_20374,N_19639,N_19798);
xor U20375 (N_20375,N_19724,N_19832);
and U20376 (N_20376,N_19785,N_19860);
nor U20377 (N_20377,N_19922,N_19506);
nand U20378 (N_20378,N_19747,N_19888);
nor U20379 (N_20379,N_19907,N_19646);
xnor U20380 (N_20380,N_19935,N_19641);
nor U20381 (N_20381,N_19980,N_19873);
xor U20382 (N_20382,N_19658,N_19973);
and U20383 (N_20383,N_19635,N_19532);
or U20384 (N_20384,N_19505,N_19941);
nand U20385 (N_20385,N_19918,N_19671);
nor U20386 (N_20386,N_19710,N_19570);
nand U20387 (N_20387,N_19540,N_19647);
and U20388 (N_20388,N_19503,N_19964);
nand U20389 (N_20389,N_19850,N_19871);
or U20390 (N_20390,N_19634,N_19512);
or U20391 (N_20391,N_19676,N_19772);
nand U20392 (N_20392,N_19546,N_19584);
xnor U20393 (N_20393,N_19751,N_19855);
nand U20394 (N_20394,N_19741,N_19692);
and U20395 (N_20395,N_19743,N_19733);
or U20396 (N_20396,N_19915,N_19737);
nand U20397 (N_20397,N_19908,N_19634);
and U20398 (N_20398,N_19698,N_19820);
nand U20399 (N_20399,N_19549,N_19909);
or U20400 (N_20400,N_19610,N_19606);
or U20401 (N_20401,N_19961,N_19753);
nor U20402 (N_20402,N_19855,N_19595);
and U20403 (N_20403,N_19964,N_19778);
nand U20404 (N_20404,N_19965,N_19867);
nor U20405 (N_20405,N_19685,N_19773);
xnor U20406 (N_20406,N_19846,N_19754);
and U20407 (N_20407,N_19742,N_19971);
and U20408 (N_20408,N_19800,N_19636);
or U20409 (N_20409,N_19581,N_19717);
xor U20410 (N_20410,N_19667,N_19956);
nor U20411 (N_20411,N_19687,N_19698);
nor U20412 (N_20412,N_19741,N_19507);
xor U20413 (N_20413,N_19894,N_19904);
or U20414 (N_20414,N_19507,N_19675);
xnor U20415 (N_20415,N_19953,N_19653);
nand U20416 (N_20416,N_19656,N_19927);
nor U20417 (N_20417,N_19725,N_19994);
nor U20418 (N_20418,N_19832,N_19998);
xor U20419 (N_20419,N_19799,N_19635);
and U20420 (N_20420,N_19745,N_19547);
or U20421 (N_20421,N_19992,N_19870);
nor U20422 (N_20422,N_19933,N_19506);
xnor U20423 (N_20423,N_19712,N_19835);
xor U20424 (N_20424,N_19534,N_19908);
nand U20425 (N_20425,N_19771,N_19888);
or U20426 (N_20426,N_19569,N_19772);
and U20427 (N_20427,N_19989,N_19671);
nand U20428 (N_20428,N_19833,N_19986);
or U20429 (N_20429,N_19994,N_19664);
and U20430 (N_20430,N_19582,N_19622);
or U20431 (N_20431,N_19535,N_19791);
xnor U20432 (N_20432,N_19933,N_19992);
xnor U20433 (N_20433,N_19658,N_19569);
or U20434 (N_20434,N_19703,N_19781);
nor U20435 (N_20435,N_19728,N_19586);
nand U20436 (N_20436,N_19638,N_19636);
or U20437 (N_20437,N_19911,N_19515);
or U20438 (N_20438,N_19863,N_19590);
nand U20439 (N_20439,N_19772,N_19526);
and U20440 (N_20440,N_19596,N_19534);
nand U20441 (N_20441,N_19784,N_19594);
nand U20442 (N_20442,N_19778,N_19934);
nand U20443 (N_20443,N_19579,N_19537);
xnor U20444 (N_20444,N_19869,N_19644);
xor U20445 (N_20445,N_19664,N_19832);
nand U20446 (N_20446,N_19789,N_19599);
or U20447 (N_20447,N_19660,N_19613);
xnor U20448 (N_20448,N_19675,N_19664);
or U20449 (N_20449,N_19594,N_19593);
xor U20450 (N_20450,N_19737,N_19910);
and U20451 (N_20451,N_19723,N_19631);
or U20452 (N_20452,N_19880,N_19695);
xor U20453 (N_20453,N_19564,N_19612);
xor U20454 (N_20454,N_19765,N_19804);
xnor U20455 (N_20455,N_19881,N_19742);
and U20456 (N_20456,N_19674,N_19896);
and U20457 (N_20457,N_19835,N_19923);
nor U20458 (N_20458,N_19992,N_19756);
nor U20459 (N_20459,N_19838,N_19968);
and U20460 (N_20460,N_19629,N_19971);
and U20461 (N_20461,N_19824,N_19832);
or U20462 (N_20462,N_19815,N_19618);
nand U20463 (N_20463,N_19980,N_19673);
nor U20464 (N_20464,N_19664,N_19821);
nor U20465 (N_20465,N_19713,N_19908);
and U20466 (N_20466,N_19691,N_19992);
or U20467 (N_20467,N_19972,N_19962);
or U20468 (N_20468,N_19953,N_19711);
nor U20469 (N_20469,N_19907,N_19991);
and U20470 (N_20470,N_19566,N_19862);
xnor U20471 (N_20471,N_19718,N_19959);
nor U20472 (N_20472,N_19596,N_19687);
xor U20473 (N_20473,N_19838,N_19615);
and U20474 (N_20474,N_19673,N_19853);
and U20475 (N_20475,N_19794,N_19649);
xor U20476 (N_20476,N_19867,N_19704);
xnor U20477 (N_20477,N_19936,N_19695);
nand U20478 (N_20478,N_19768,N_19802);
and U20479 (N_20479,N_19631,N_19741);
and U20480 (N_20480,N_19778,N_19666);
nor U20481 (N_20481,N_19758,N_19887);
or U20482 (N_20482,N_19648,N_19955);
and U20483 (N_20483,N_19979,N_19695);
nor U20484 (N_20484,N_19709,N_19693);
xnor U20485 (N_20485,N_19978,N_19939);
nand U20486 (N_20486,N_19709,N_19672);
xor U20487 (N_20487,N_19804,N_19700);
nand U20488 (N_20488,N_19907,N_19777);
and U20489 (N_20489,N_19986,N_19848);
and U20490 (N_20490,N_19943,N_19992);
nor U20491 (N_20491,N_19981,N_19810);
or U20492 (N_20492,N_19711,N_19626);
nand U20493 (N_20493,N_19729,N_19590);
xor U20494 (N_20494,N_19802,N_19817);
xnor U20495 (N_20495,N_19743,N_19857);
and U20496 (N_20496,N_19950,N_19512);
and U20497 (N_20497,N_19500,N_19801);
nor U20498 (N_20498,N_19708,N_19558);
nand U20499 (N_20499,N_19995,N_19896);
and U20500 (N_20500,N_20482,N_20003);
or U20501 (N_20501,N_20066,N_20440);
and U20502 (N_20502,N_20158,N_20087);
xor U20503 (N_20503,N_20307,N_20364);
xor U20504 (N_20504,N_20162,N_20314);
and U20505 (N_20505,N_20035,N_20232);
or U20506 (N_20506,N_20292,N_20411);
nor U20507 (N_20507,N_20115,N_20049);
nor U20508 (N_20508,N_20337,N_20370);
or U20509 (N_20509,N_20446,N_20209);
or U20510 (N_20510,N_20227,N_20156);
xor U20511 (N_20511,N_20101,N_20058);
xor U20512 (N_20512,N_20461,N_20075);
xor U20513 (N_20513,N_20404,N_20044);
nor U20514 (N_20514,N_20006,N_20384);
xnor U20515 (N_20515,N_20221,N_20485);
or U20516 (N_20516,N_20431,N_20183);
nand U20517 (N_20517,N_20332,N_20286);
nor U20518 (N_20518,N_20192,N_20185);
xor U20519 (N_20519,N_20095,N_20022);
nor U20520 (N_20520,N_20243,N_20424);
nand U20521 (N_20521,N_20420,N_20248);
nor U20522 (N_20522,N_20477,N_20353);
nand U20523 (N_20523,N_20447,N_20074);
xnor U20524 (N_20524,N_20208,N_20394);
and U20525 (N_20525,N_20426,N_20236);
or U20526 (N_20526,N_20050,N_20112);
nor U20527 (N_20527,N_20105,N_20055);
or U20528 (N_20528,N_20172,N_20310);
xnor U20529 (N_20529,N_20182,N_20407);
nand U20530 (N_20530,N_20423,N_20285);
nand U20531 (N_20531,N_20177,N_20282);
nor U20532 (N_20532,N_20478,N_20422);
and U20533 (N_20533,N_20359,N_20316);
nor U20534 (N_20534,N_20122,N_20257);
xnor U20535 (N_20535,N_20202,N_20492);
or U20536 (N_20536,N_20311,N_20439);
xor U20537 (N_20537,N_20014,N_20067);
xor U20538 (N_20538,N_20076,N_20081);
xor U20539 (N_20539,N_20457,N_20261);
nand U20540 (N_20540,N_20358,N_20263);
or U20541 (N_20541,N_20296,N_20387);
xnor U20542 (N_20542,N_20019,N_20334);
or U20543 (N_20543,N_20152,N_20442);
or U20544 (N_20544,N_20195,N_20175);
nand U20545 (N_20545,N_20487,N_20252);
nor U20546 (N_20546,N_20275,N_20323);
xnor U20547 (N_20547,N_20024,N_20166);
nand U20548 (N_20548,N_20410,N_20110);
and U20549 (N_20549,N_20028,N_20490);
or U20550 (N_20550,N_20373,N_20325);
nand U20551 (N_20551,N_20378,N_20348);
and U20552 (N_20552,N_20349,N_20454);
nor U20553 (N_20553,N_20231,N_20381);
xnor U20554 (N_20554,N_20142,N_20109);
and U20555 (N_20555,N_20377,N_20124);
xnor U20556 (N_20556,N_20057,N_20456);
nor U20557 (N_20557,N_20015,N_20437);
nor U20558 (N_20558,N_20472,N_20097);
xnor U20559 (N_20559,N_20179,N_20059);
or U20560 (N_20560,N_20056,N_20294);
nand U20561 (N_20561,N_20464,N_20123);
and U20562 (N_20562,N_20386,N_20260);
xnor U20563 (N_20563,N_20086,N_20465);
xor U20564 (N_20564,N_20018,N_20368);
nor U20565 (N_20565,N_20379,N_20374);
xor U20566 (N_20566,N_20321,N_20107);
nand U20567 (N_20567,N_20299,N_20499);
nand U20568 (N_20568,N_20238,N_20395);
nor U20569 (N_20569,N_20388,N_20168);
xor U20570 (N_20570,N_20144,N_20428);
xnor U20571 (N_20571,N_20119,N_20229);
nor U20572 (N_20572,N_20127,N_20191);
nor U20573 (N_20573,N_20204,N_20020);
or U20574 (N_20574,N_20392,N_20397);
nand U20575 (N_20575,N_20079,N_20017);
or U20576 (N_20576,N_20013,N_20295);
nor U20577 (N_20577,N_20133,N_20154);
nand U20578 (N_20578,N_20201,N_20355);
nand U20579 (N_20579,N_20190,N_20145);
xnor U20580 (N_20580,N_20429,N_20458);
and U20581 (N_20581,N_20432,N_20371);
and U20582 (N_20582,N_20489,N_20106);
xor U20583 (N_20583,N_20413,N_20093);
xnor U20584 (N_20584,N_20290,N_20491);
or U20585 (N_20585,N_20302,N_20343);
or U20586 (N_20586,N_20161,N_20433);
or U20587 (N_20587,N_20047,N_20137);
nor U20588 (N_20588,N_20138,N_20249);
or U20589 (N_20589,N_20148,N_20289);
nand U20590 (N_20590,N_20210,N_20273);
or U20591 (N_20591,N_20130,N_20244);
nor U20592 (N_20592,N_20046,N_20329);
nand U20593 (N_20593,N_20441,N_20063);
or U20594 (N_20594,N_20279,N_20000);
and U20595 (N_20595,N_20459,N_20308);
nor U20596 (N_20596,N_20467,N_20113);
nor U20597 (N_20597,N_20409,N_20463);
or U20598 (N_20598,N_20002,N_20088);
nor U20599 (N_20599,N_20488,N_20254);
and U20600 (N_20600,N_20198,N_20449);
or U20601 (N_20601,N_20274,N_20320);
and U20602 (N_20602,N_20470,N_20346);
nand U20603 (N_20603,N_20434,N_20258);
and U20604 (N_20604,N_20205,N_20425);
xnor U20605 (N_20605,N_20186,N_20230);
nor U20606 (N_20606,N_20139,N_20116);
xnor U20607 (N_20607,N_20173,N_20473);
and U20608 (N_20608,N_20288,N_20197);
nor U20609 (N_20609,N_20284,N_20027);
xor U20610 (N_20610,N_20151,N_20178);
nor U20611 (N_20611,N_20222,N_20398);
nand U20612 (N_20612,N_20268,N_20400);
or U20613 (N_20613,N_20469,N_20300);
and U20614 (N_20614,N_20012,N_20207);
nor U20615 (N_20615,N_20008,N_20427);
nand U20616 (N_20616,N_20167,N_20132);
nand U20617 (N_20617,N_20150,N_20025);
or U20618 (N_20618,N_20077,N_20141);
xnor U20619 (N_20619,N_20318,N_20042);
nor U20620 (N_20620,N_20453,N_20474);
and U20621 (N_20621,N_20234,N_20073);
nor U20622 (N_20622,N_20089,N_20224);
xnor U20623 (N_20623,N_20496,N_20078);
and U20624 (N_20624,N_20096,N_20324);
or U20625 (N_20625,N_20217,N_20389);
xnor U20626 (N_20626,N_20341,N_20436);
nand U20627 (N_20627,N_20125,N_20111);
and U20628 (N_20628,N_20351,N_20365);
nand U20629 (N_20629,N_20216,N_20497);
xnor U20630 (N_20630,N_20354,N_20196);
and U20631 (N_20631,N_20493,N_20445);
nand U20632 (N_20632,N_20038,N_20328);
xor U20633 (N_20633,N_20287,N_20401);
nand U20634 (N_20634,N_20091,N_20382);
or U20635 (N_20635,N_20291,N_20233);
or U20636 (N_20636,N_20468,N_20034);
or U20637 (N_20637,N_20303,N_20357);
xnor U20638 (N_20638,N_20266,N_20312);
and U20639 (N_20639,N_20061,N_20011);
xnor U20640 (N_20640,N_20481,N_20309);
and U20641 (N_20641,N_20272,N_20235);
xnor U20642 (N_20642,N_20180,N_20418);
and U20643 (N_20643,N_20475,N_20242);
xor U20644 (N_20644,N_20052,N_20054);
nor U20645 (N_20645,N_20301,N_20016);
nand U20646 (N_20646,N_20147,N_20246);
and U20647 (N_20647,N_20188,N_20265);
and U20648 (N_20648,N_20170,N_20149);
nand U20649 (N_20649,N_20072,N_20251);
xnor U20650 (N_20650,N_20225,N_20319);
xor U20651 (N_20651,N_20065,N_20080);
and U20652 (N_20652,N_20444,N_20356);
nor U20653 (N_20653,N_20108,N_20193);
xor U20654 (N_20654,N_20062,N_20476);
or U20655 (N_20655,N_20206,N_20339);
and U20656 (N_20656,N_20450,N_20250);
or U20657 (N_20657,N_20462,N_20102);
and U20658 (N_20658,N_20118,N_20369);
and U20659 (N_20659,N_20283,N_20333);
xnor U20660 (N_20660,N_20304,N_20114);
and U20661 (N_20661,N_20160,N_20281);
and U20662 (N_20662,N_20406,N_20376);
xnor U20663 (N_20663,N_20211,N_20181);
xor U20664 (N_20664,N_20347,N_20099);
nand U20665 (N_20665,N_20345,N_20455);
nor U20666 (N_20666,N_20494,N_20342);
xnor U20667 (N_20667,N_20043,N_20435);
and U20668 (N_20668,N_20200,N_20270);
or U20669 (N_20669,N_20070,N_20448);
xnor U20670 (N_20670,N_20094,N_20245);
xnor U20671 (N_20671,N_20335,N_20452);
and U20672 (N_20672,N_20164,N_20327);
and U20673 (N_20673,N_20103,N_20082);
and U20674 (N_20674,N_20001,N_20483);
or U20675 (N_20675,N_20240,N_20068);
or U20676 (N_20676,N_20129,N_20215);
nand U20677 (N_20677,N_20253,N_20030);
nor U20678 (N_20678,N_20412,N_20479);
or U20679 (N_20679,N_20048,N_20415);
or U20680 (N_20680,N_20135,N_20009);
xor U20681 (N_20681,N_20029,N_20298);
nand U20682 (N_20682,N_20220,N_20414);
nor U20683 (N_20683,N_20471,N_20344);
or U20684 (N_20684,N_20226,N_20331);
xor U20685 (N_20685,N_20120,N_20023);
nand U20686 (N_20686,N_20367,N_20187);
and U20687 (N_20687,N_20495,N_20143);
or U20688 (N_20688,N_20053,N_20383);
xnor U20689 (N_20689,N_20098,N_20189);
xnor U20690 (N_20690,N_20010,N_20443);
and U20691 (N_20691,N_20498,N_20218);
nor U20692 (N_20692,N_20360,N_20363);
nand U20693 (N_20693,N_20159,N_20163);
xnor U20694 (N_20694,N_20361,N_20203);
or U20695 (N_20695,N_20267,N_20060);
nor U20696 (N_20696,N_20037,N_20280);
and U20697 (N_20697,N_20085,N_20402);
xor U20698 (N_20698,N_20033,N_20092);
xnor U20699 (N_20699,N_20199,N_20326);
or U20700 (N_20700,N_20297,N_20071);
or U20701 (N_20701,N_20100,N_20486);
or U20702 (N_20702,N_20157,N_20064);
nor U20703 (N_20703,N_20338,N_20126);
nor U20704 (N_20704,N_20480,N_20090);
and U20705 (N_20705,N_20391,N_20393);
and U20706 (N_20706,N_20223,N_20131);
nand U20707 (N_20707,N_20399,N_20390);
nand U20708 (N_20708,N_20277,N_20278);
xor U20709 (N_20709,N_20219,N_20237);
and U20710 (N_20710,N_20315,N_20362);
or U20711 (N_20711,N_20269,N_20069);
and U20712 (N_20712,N_20134,N_20262);
nand U20713 (N_20713,N_20184,N_20031);
and U20714 (N_20714,N_20430,N_20405);
nor U20715 (N_20715,N_20239,N_20313);
xnor U20716 (N_20716,N_20336,N_20032);
nor U20717 (N_20717,N_20104,N_20128);
xnor U20718 (N_20718,N_20256,N_20438);
nor U20719 (N_20719,N_20375,N_20350);
nor U20720 (N_20720,N_20212,N_20174);
and U20721 (N_20721,N_20322,N_20271);
nor U20722 (N_20722,N_20408,N_20293);
nor U20723 (N_20723,N_20039,N_20004);
nor U20724 (N_20724,N_20045,N_20146);
nor U20725 (N_20725,N_20121,N_20380);
nand U20726 (N_20726,N_20255,N_20385);
nand U20727 (N_20727,N_20194,N_20317);
nor U20728 (N_20728,N_20007,N_20466);
nand U20729 (N_20729,N_20306,N_20026);
nand U20730 (N_20730,N_20451,N_20330);
nor U20731 (N_20731,N_20136,N_20084);
nor U20732 (N_20732,N_20340,N_20228);
or U20733 (N_20733,N_20171,N_20247);
or U20734 (N_20734,N_20051,N_20484);
xnor U20735 (N_20735,N_20421,N_20176);
xnor U20736 (N_20736,N_20366,N_20153);
xor U20737 (N_20737,N_20241,N_20040);
nand U20738 (N_20738,N_20372,N_20140);
nor U20739 (N_20739,N_20460,N_20169);
and U20740 (N_20740,N_20264,N_20214);
and U20741 (N_20741,N_20352,N_20419);
xor U20742 (N_20742,N_20036,N_20213);
nand U20743 (N_20743,N_20276,N_20165);
nor U20744 (N_20744,N_20259,N_20417);
or U20745 (N_20745,N_20021,N_20305);
nand U20746 (N_20746,N_20155,N_20416);
and U20747 (N_20747,N_20396,N_20005);
and U20748 (N_20748,N_20403,N_20117);
and U20749 (N_20749,N_20083,N_20041);
nor U20750 (N_20750,N_20162,N_20390);
and U20751 (N_20751,N_20401,N_20453);
and U20752 (N_20752,N_20335,N_20490);
nor U20753 (N_20753,N_20090,N_20288);
nor U20754 (N_20754,N_20454,N_20312);
or U20755 (N_20755,N_20272,N_20229);
nor U20756 (N_20756,N_20052,N_20091);
or U20757 (N_20757,N_20291,N_20021);
and U20758 (N_20758,N_20304,N_20270);
xnor U20759 (N_20759,N_20137,N_20278);
and U20760 (N_20760,N_20399,N_20424);
nand U20761 (N_20761,N_20443,N_20344);
and U20762 (N_20762,N_20095,N_20114);
xor U20763 (N_20763,N_20090,N_20107);
nor U20764 (N_20764,N_20391,N_20483);
nand U20765 (N_20765,N_20311,N_20383);
xor U20766 (N_20766,N_20210,N_20126);
nand U20767 (N_20767,N_20298,N_20178);
nor U20768 (N_20768,N_20433,N_20233);
xnor U20769 (N_20769,N_20267,N_20376);
and U20770 (N_20770,N_20011,N_20093);
or U20771 (N_20771,N_20123,N_20209);
nand U20772 (N_20772,N_20083,N_20095);
nand U20773 (N_20773,N_20310,N_20340);
xor U20774 (N_20774,N_20340,N_20281);
nor U20775 (N_20775,N_20457,N_20098);
nand U20776 (N_20776,N_20161,N_20219);
and U20777 (N_20777,N_20054,N_20313);
and U20778 (N_20778,N_20235,N_20362);
or U20779 (N_20779,N_20413,N_20216);
nor U20780 (N_20780,N_20214,N_20450);
nand U20781 (N_20781,N_20276,N_20448);
and U20782 (N_20782,N_20137,N_20403);
nor U20783 (N_20783,N_20200,N_20452);
or U20784 (N_20784,N_20106,N_20252);
xor U20785 (N_20785,N_20357,N_20355);
nor U20786 (N_20786,N_20357,N_20347);
xor U20787 (N_20787,N_20183,N_20258);
nor U20788 (N_20788,N_20343,N_20051);
nand U20789 (N_20789,N_20397,N_20454);
xor U20790 (N_20790,N_20015,N_20250);
nor U20791 (N_20791,N_20027,N_20127);
nand U20792 (N_20792,N_20385,N_20145);
nor U20793 (N_20793,N_20460,N_20065);
and U20794 (N_20794,N_20246,N_20054);
or U20795 (N_20795,N_20001,N_20346);
nand U20796 (N_20796,N_20196,N_20244);
and U20797 (N_20797,N_20298,N_20187);
xor U20798 (N_20798,N_20338,N_20311);
nand U20799 (N_20799,N_20229,N_20074);
or U20800 (N_20800,N_20235,N_20242);
nand U20801 (N_20801,N_20038,N_20211);
nand U20802 (N_20802,N_20019,N_20192);
and U20803 (N_20803,N_20405,N_20193);
xnor U20804 (N_20804,N_20445,N_20478);
or U20805 (N_20805,N_20125,N_20229);
nand U20806 (N_20806,N_20320,N_20225);
nor U20807 (N_20807,N_20071,N_20467);
xnor U20808 (N_20808,N_20478,N_20130);
xor U20809 (N_20809,N_20207,N_20263);
or U20810 (N_20810,N_20210,N_20272);
nor U20811 (N_20811,N_20170,N_20134);
or U20812 (N_20812,N_20040,N_20102);
xor U20813 (N_20813,N_20069,N_20077);
nor U20814 (N_20814,N_20095,N_20412);
xnor U20815 (N_20815,N_20267,N_20075);
and U20816 (N_20816,N_20262,N_20098);
and U20817 (N_20817,N_20130,N_20305);
xor U20818 (N_20818,N_20036,N_20257);
and U20819 (N_20819,N_20078,N_20104);
xor U20820 (N_20820,N_20273,N_20307);
or U20821 (N_20821,N_20084,N_20467);
or U20822 (N_20822,N_20206,N_20359);
and U20823 (N_20823,N_20369,N_20382);
nor U20824 (N_20824,N_20392,N_20489);
or U20825 (N_20825,N_20474,N_20276);
and U20826 (N_20826,N_20154,N_20355);
or U20827 (N_20827,N_20390,N_20108);
nand U20828 (N_20828,N_20466,N_20058);
xor U20829 (N_20829,N_20225,N_20348);
nor U20830 (N_20830,N_20495,N_20313);
and U20831 (N_20831,N_20019,N_20287);
nand U20832 (N_20832,N_20392,N_20277);
or U20833 (N_20833,N_20269,N_20106);
nand U20834 (N_20834,N_20009,N_20465);
nand U20835 (N_20835,N_20110,N_20129);
nor U20836 (N_20836,N_20451,N_20492);
nand U20837 (N_20837,N_20049,N_20195);
or U20838 (N_20838,N_20057,N_20406);
nand U20839 (N_20839,N_20162,N_20326);
xnor U20840 (N_20840,N_20406,N_20266);
nand U20841 (N_20841,N_20002,N_20410);
and U20842 (N_20842,N_20141,N_20489);
nor U20843 (N_20843,N_20178,N_20451);
or U20844 (N_20844,N_20025,N_20050);
nand U20845 (N_20845,N_20207,N_20431);
nand U20846 (N_20846,N_20440,N_20439);
and U20847 (N_20847,N_20039,N_20003);
nand U20848 (N_20848,N_20255,N_20023);
nor U20849 (N_20849,N_20321,N_20227);
nor U20850 (N_20850,N_20359,N_20062);
nand U20851 (N_20851,N_20057,N_20169);
and U20852 (N_20852,N_20178,N_20425);
and U20853 (N_20853,N_20135,N_20286);
or U20854 (N_20854,N_20269,N_20487);
xor U20855 (N_20855,N_20175,N_20299);
nor U20856 (N_20856,N_20462,N_20345);
nand U20857 (N_20857,N_20105,N_20063);
nand U20858 (N_20858,N_20196,N_20222);
or U20859 (N_20859,N_20189,N_20175);
and U20860 (N_20860,N_20084,N_20348);
nand U20861 (N_20861,N_20241,N_20078);
xor U20862 (N_20862,N_20115,N_20330);
and U20863 (N_20863,N_20203,N_20282);
nand U20864 (N_20864,N_20391,N_20131);
or U20865 (N_20865,N_20160,N_20221);
and U20866 (N_20866,N_20446,N_20191);
nor U20867 (N_20867,N_20309,N_20138);
and U20868 (N_20868,N_20142,N_20216);
nand U20869 (N_20869,N_20357,N_20247);
xnor U20870 (N_20870,N_20159,N_20404);
or U20871 (N_20871,N_20011,N_20007);
nand U20872 (N_20872,N_20400,N_20137);
and U20873 (N_20873,N_20274,N_20260);
and U20874 (N_20874,N_20271,N_20443);
or U20875 (N_20875,N_20387,N_20375);
or U20876 (N_20876,N_20453,N_20112);
nor U20877 (N_20877,N_20409,N_20241);
xor U20878 (N_20878,N_20448,N_20285);
nand U20879 (N_20879,N_20344,N_20163);
nand U20880 (N_20880,N_20180,N_20242);
xnor U20881 (N_20881,N_20467,N_20410);
and U20882 (N_20882,N_20411,N_20238);
or U20883 (N_20883,N_20119,N_20436);
xnor U20884 (N_20884,N_20368,N_20426);
nand U20885 (N_20885,N_20353,N_20297);
nand U20886 (N_20886,N_20325,N_20329);
xor U20887 (N_20887,N_20416,N_20011);
or U20888 (N_20888,N_20106,N_20043);
xnor U20889 (N_20889,N_20349,N_20310);
nor U20890 (N_20890,N_20312,N_20270);
or U20891 (N_20891,N_20241,N_20364);
xor U20892 (N_20892,N_20274,N_20453);
nor U20893 (N_20893,N_20230,N_20438);
and U20894 (N_20894,N_20283,N_20047);
nand U20895 (N_20895,N_20465,N_20343);
or U20896 (N_20896,N_20354,N_20035);
or U20897 (N_20897,N_20473,N_20062);
or U20898 (N_20898,N_20485,N_20088);
nor U20899 (N_20899,N_20033,N_20119);
nor U20900 (N_20900,N_20071,N_20104);
and U20901 (N_20901,N_20226,N_20063);
or U20902 (N_20902,N_20258,N_20177);
or U20903 (N_20903,N_20218,N_20291);
or U20904 (N_20904,N_20229,N_20305);
xor U20905 (N_20905,N_20493,N_20061);
nor U20906 (N_20906,N_20214,N_20020);
and U20907 (N_20907,N_20269,N_20358);
and U20908 (N_20908,N_20104,N_20025);
or U20909 (N_20909,N_20224,N_20189);
nor U20910 (N_20910,N_20108,N_20495);
and U20911 (N_20911,N_20147,N_20131);
and U20912 (N_20912,N_20139,N_20424);
xor U20913 (N_20913,N_20105,N_20044);
and U20914 (N_20914,N_20008,N_20279);
nor U20915 (N_20915,N_20063,N_20210);
nand U20916 (N_20916,N_20233,N_20486);
and U20917 (N_20917,N_20284,N_20323);
xor U20918 (N_20918,N_20178,N_20407);
xor U20919 (N_20919,N_20029,N_20366);
and U20920 (N_20920,N_20355,N_20160);
or U20921 (N_20921,N_20260,N_20335);
nor U20922 (N_20922,N_20261,N_20372);
and U20923 (N_20923,N_20211,N_20064);
or U20924 (N_20924,N_20126,N_20345);
nand U20925 (N_20925,N_20111,N_20354);
or U20926 (N_20926,N_20420,N_20344);
or U20927 (N_20927,N_20108,N_20409);
and U20928 (N_20928,N_20413,N_20466);
or U20929 (N_20929,N_20255,N_20019);
nor U20930 (N_20930,N_20000,N_20189);
nand U20931 (N_20931,N_20013,N_20389);
xor U20932 (N_20932,N_20173,N_20208);
and U20933 (N_20933,N_20382,N_20448);
xor U20934 (N_20934,N_20094,N_20419);
and U20935 (N_20935,N_20308,N_20148);
nand U20936 (N_20936,N_20032,N_20490);
nor U20937 (N_20937,N_20032,N_20015);
or U20938 (N_20938,N_20222,N_20075);
nor U20939 (N_20939,N_20170,N_20010);
and U20940 (N_20940,N_20319,N_20009);
or U20941 (N_20941,N_20348,N_20236);
nand U20942 (N_20942,N_20018,N_20364);
nand U20943 (N_20943,N_20351,N_20273);
nand U20944 (N_20944,N_20081,N_20482);
or U20945 (N_20945,N_20119,N_20444);
xor U20946 (N_20946,N_20480,N_20252);
nor U20947 (N_20947,N_20178,N_20404);
or U20948 (N_20948,N_20442,N_20291);
and U20949 (N_20949,N_20455,N_20476);
nor U20950 (N_20950,N_20373,N_20116);
nor U20951 (N_20951,N_20148,N_20128);
nand U20952 (N_20952,N_20477,N_20423);
or U20953 (N_20953,N_20474,N_20297);
nand U20954 (N_20954,N_20126,N_20467);
nand U20955 (N_20955,N_20402,N_20408);
nor U20956 (N_20956,N_20421,N_20090);
or U20957 (N_20957,N_20165,N_20091);
nor U20958 (N_20958,N_20475,N_20144);
nand U20959 (N_20959,N_20118,N_20278);
nor U20960 (N_20960,N_20035,N_20037);
nor U20961 (N_20961,N_20263,N_20454);
nor U20962 (N_20962,N_20094,N_20374);
or U20963 (N_20963,N_20034,N_20363);
or U20964 (N_20964,N_20005,N_20238);
xor U20965 (N_20965,N_20048,N_20159);
and U20966 (N_20966,N_20193,N_20112);
xnor U20967 (N_20967,N_20334,N_20090);
nand U20968 (N_20968,N_20415,N_20114);
xor U20969 (N_20969,N_20355,N_20438);
xnor U20970 (N_20970,N_20095,N_20449);
nor U20971 (N_20971,N_20457,N_20320);
and U20972 (N_20972,N_20255,N_20286);
and U20973 (N_20973,N_20189,N_20137);
or U20974 (N_20974,N_20474,N_20205);
nand U20975 (N_20975,N_20230,N_20200);
xnor U20976 (N_20976,N_20427,N_20455);
nor U20977 (N_20977,N_20126,N_20360);
and U20978 (N_20978,N_20180,N_20002);
xor U20979 (N_20979,N_20319,N_20015);
or U20980 (N_20980,N_20443,N_20113);
and U20981 (N_20981,N_20209,N_20258);
or U20982 (N_20982,N_20476,N_20008);
nand U20983 (N_20983,N_20377,N_20311);
or U20984 (N_20984,N_20435,N_20031);
nand U20985 (N_20985,N_20249,N_20367);
and U20986 (N_20986,N_20022,N_20397);
and U20987 (N_20987,N_20093,N_20234);
and U20988 (N_20988,N_20293,N_20354);
xor U20989 (N_20989,N_20158,N_20216);
xor U20990 (N_20990,N_20438,N_20445);
and U20991 (N_20991,N_20304,N_20324);
and U20992 (N_20992,N_20271,N_20323);
or U20993 (N_20993,N_20194,N_20336);
xnor U20994 (N_20994,N_20064,N_20468);
or U20995 (N_20995,N_20097,N_20116);
xnor U20996 (N_20996,N_20285,N_20194);
nand U20997 (N_20997,N_20181,N_20480);
nor U20998 (N_20998,N_20217,N_20325);
xor U20999 (N_20999,N_20238,N_20016);
or U21000 (N_21000,N_20991,N_20824);
nor U21001 (N_21001,N_20626,N_20630);
or U21002 (N_21002,N_20948,N_20549);
xor U21003 (N_21003,N_20953,N_20585);
xnor U21004 (N_21004,N_20998,N_20665);
nor U21005 (N_21005,N_20971,N_20992);
nand U21006 (N_21006,N_20691,N_20523);
and U21007 (N_21007,N_20961,N_20956);
or U21008 (N_21008,N_20543,N_20818);
and U21009 (N_21009,N_20724,N_20726);
xor U21010 (N_21010,N_20879,N_20624);
or U21011 (N_21011,N_20609,N_20955);
nor U21012 (N_21012,N_20976,N_20872);
and U21013 (N_21013,N_20914,N_20932);
xor U21014 (N_21014,N_20968,N_20615);
and U21015 (N_21015,N_20735,N_20988);
nor U21016 (N_21016,N_20973,N_20518);
xnor U21017 (N_21017,N_20690,N_20892);
nand U21018 (N_21018,N_20516,N_20551);
xor U21019 (N_21019,N_20531,N_20591);
nand U21020 (N_21020,N_20693,N_20538);
nand U21021 (N_21021,N_20852,N_20838);
and U21022 (N_21022,N_20813,N_20781);
nor U21023 (N_21023,N_20667,N_20946);
nor U21024 (N_21024,N_20796,N_20598);
or U21025 (N_21025,N_20696,N_20515);
nand U21026 (N_21026,N_20773,N_20808);
nand U21027 (N_21027,N_20895,N_20700);
nor U21028 (N_21028,N_20997,N_20625);
nor U21029 (N_21029,N_20705,N_20736);
and U21030 (N_21030,N_20703,N_20763);
xnor U21031 (N_21031,N_20754,N_20602);
nand U21032 (N_21032,N_20534,N_20850);
and U21033 (N_21033,N_20556,N_20827);
nand U21034 (N_21034,N_20897,N_20521);
nand U21035 (N_21035,N_20651,N_20588);
xor U21036 (N_21036,N_20654,N_20788);
nand U21037 (N_21037,N_20981,N_20682);
and U21038 (N_21038,N_20987,N_20554);
and U21039 (N_21039,N_20837,N_20980);
xor U21040 (N_21040,N_20566,N_20666);
nand U21041 (N_21041,N_20923,N_20712);
xor U21042 (N_21042,N_20775,N_20964);
and U21043 (N_21043,N_20590,N_20727);
nand U21044 (N_21044,N_20740,N_20799);
and U21045 (N_21045,N_20750,N_20883);
xor U21046 (N_21046,N_20878,N_20568);
or U21047 (N_21047,N_20650,N_20848);
or U21048 (N_21048,N_20701,N_20795);
xnor U21049 (N_21049,N_20996,N_20683);
nor U21050 (N_21050,N_20755,N_20600);
or U21051 (N_21051,N_20637,N_20919);
nand U21052 (N_21052,N_20714,N_20890);
nand U21053 (N_21053,N_20513,N_20634);
or U21054 (N_21054,N_20839,N_20863);
or U21055 (N_21055,N_20702,N_20514);
or U21056 (N_21056,N_20884,N_20594);
nor U21057 (N_21057,N_20698,N_20849);
nor U21058 (N_21058,N_20765,N_20669);
or U21059 (N_21059,N_20542,N_20752);
xor U21060 (N_21060,N_20638,N_20584);
xor U21061 (N_21061,N_20743,N_20871);
nand U21062 (N_21062,N_20989,N_20966);
xor U21063 (N_21063,N_20646,N_20592);
nor U21064 (N_21064,N_20934,N_20774);
xor U21065 (N_21065,N_20718,N_20512);
nor U21066 (N_21066,N_20560,N_20915);
or U21067 (N_21067,N_20668,N_20604);
or U21068 (N_21068,N_20757,N_20832);
nand U21069 (N_21069,N_20678,N_20741);
xnor U21070 (N_21070,N_20957,N_20937);
and U21071 (N_21071,N_20672,N_20815);
nor U21072 (N_21072,N_20572,N_20503);
xnor U21073 (N_21073,N_20901,N_20906);
and U21074 (N_21074,N_20939,N_20975);
xnor U21075 (N_21075,N_20797,N_20717);
and U21076 (N_21076,N_20926,N_20661);
and U21077 (N_21077,N_20504,N_20784);
or U21078 (N_21078,N_20771,N_20685);
nor U21079 (N_21079,N_20739,N_20697);
or U21080 (N_21080,N_20607,N_20835);
xnor U21081 (N_21081,N_20532,N_20864);
nor U21082 (N_21082,N_20894,N_20836);
nor U21083 (N_21083,N_20876,N_20561);
nand U21084 (N_21084,N_20927,N_20681);
and U21085 (N_21085,N_20785,N_20649);
nor U21086 (N_21086,N_20655,N_20579);
and U21087 (N_21087,N_20911,N_20574);
nor U21088 (N_21088,N_20645,N_20621);
nor U21089 (N_21089,N_20880,N_20967);
nand U21090 (N_21090,N_20522,N_20870);
or U21091 (N_21091,N_20898,N_20581);
nand U21092 (N_21092,N_20641,N_20575);
or U21093 (N_21093,N_20858,N_20627);
or U21094 (N_21094,N_20760,N_20546);
nand U21095 (N_21095,N_20840,N_20605);
or U21096 (N_21096,N_20845,N_20644);
nand U21097 (N_21097,N_20935,N_20983);
nor U21098 (N_21098,N_20722,N_20569);
nand U21099 (N_21099,N_20817,N_20768);
xor U21100 (N_21100,N_20707,N_20558);
nand U21101 (N_21101,N_20555,N_20606);
nand U21102 (N_21102,N_20586,N_20986);
xnor U21103 (N_21103,N_20648,N_20677);
xor U21104 (N_21104,N_20629,N_20943);
nor U21105 (N_21105,N_20704,N_20954);
xor U21106 (N_21106,N_20804,N_20596);
and U21107 (N_21107,N_20676,N_20947);
and U21108 (N_21108,N_20982,N_20603);
nor U21109 (N_21109,N_20933,N_20821);
or U21110 (N_21110,N_20559,N_20731);
nor U21111 (N_21111,N_20732,N_20951);
xnor U21112 (N_21112,N_20537,N_20619);
xnor U21113 (N_21113,N_20814,N_20689);
nor U21114 (N_21114,N_20793,N_20944);
xor U21115 (N_21115,N_20580,N_20995);
and U21116 (N_21116,N_20803,N_20656);
or U21117 (N_21117,N_20830,N_20801);
nor U21118 (N_21118,N_20610,N_20636);
or U21119 (N_21119,N_20847,N_20779);
xor U21120 (N_21120,N_20553,N_20529);
xnor U21121 (N_21121,N_20900,N_20563);
xor U21122 (N_21122,N_20823,N_20974);
nand U21123 (N_21123,N_20660,N_20709);
or U21124 (N_21124,N_20857,N_20859);
and U21125 (N_21125,N_20776,N_20965);
nor U21126 (N_21126,N_20524,N_20977);
xor U21127 (N_21127,N_20545,N_20940);
or U21128 (N_21128,N_20907,N_20684);
and U21129 (N_21129,N_20969,N_20652);
nand U21130 (N_21130,N_20608,N_20505);
nand U21131 (N_21131,N_20647,N_20548);
nor U21132 (N_21132,N_20922,N_20936);
xor U21133 (N_21133,N_20544,N_20786);
and U21134 (N_21134,N_20861,N_20908);
nand U21135 (N_21135,N_20787,N_20500);
or U21136 (N_21136,N_20766,N_20674);
and U21137 (N_21137,N_20846,N_20749);
nand U21138 (N_21138,N_20659,N_20843);
or U21139 (N_21139,N_20924,N_20806);
xnor U21140 (N_21140,N_20893,N_20541);
xnor U21141 (N_21141,N_20885,N_20753);
xor U21142 (N_21142,N_20565,N_20782);
and U21143 (N_21143,N_20509,N_20931);
and U21144 (N_21144,N_20737,N_20868);
or U21145 (N_21145,N_20617,N_20562);
and U21146 (N_21146,N_20962,N_20730);
nor U21147 (N_21147,N_20589,N_20738);
or U21148 (N_21148,N_20734,N_20611);
xor U21149 (N_21149,N_20673,N_20970);
and U21150 (N_21150,N_20886,N_20770);
nand U21151 (N_21151,N_20517,N_20820);
nor U21152 (N_21152,N_20819,N_20903);
nand U21153 (N_21153,N_20519,N_20834);
or U21154 (N_21154,N_20816,N_20692);
and U21155 (N_21155,N_20728,N_20622);
nand U21156 (N_21156,N_20597,N_20599);
or U21157 (N_21157,N_20929,N_20904);
or U21158 (N_21158,N_20642,N_20822);
nand U21159 (N_21159,N_20710,N_20751);
nor U21160 (N_21160,N_20688,N_20985);
or U21161 (N_21161,N_20881,N_20916);
and U21162 (N_21162,N_20950,N_20960);
nor U21163 (N_21163,N_20664,N_20557);
or U21164 (N_21164,N_20745,N_20587);
nand U21165 (N_21165,N_20811,N_20748);
nor U21166 (N_21166,N_20530,N_20866);
and U21167 (N_21167,N_20875,N_20792);
nand U21168 (N_21168,N_20632,N_20789);
and U21169 (N_21169,N_20525,N_20826);
xor U21170 (N_21170,N_20720,N_20620);
nand U21171 (N_21171,N_20507,N_20829);
nor U21172 (N_21172,N_20662,N_20595);
or U21173 (N_21173,N_20733,N_20899);
nor U21174 (N_21174,N_20547,N_20759);
or U21175 (N_21175,N_20680,N_20614);
and U21176 (N_21176,N_20582,N_20510);
xor U21177 (N_21177,N_20536,N_20601);
or U21178 (N_21178,N_20993,N_20844);
or U21179 (N_21179,N_20540,N_20912);
nor U21180 (N_21180,N_20984,N_20888);
or U21181 (N_21181,N_20508,N_20670);
nor U21182 (N_21182,N_20851,N_20723);
or U21183 (N_21183,N_20952,N_20764);
nand U21184 (N_21184,N_20708,N_20694);
nor U21185 (N_21185,N_20772,N_20635);
and U21186 (N_21186,N_20618,N_20778);
nand U21187 (N_21187,N_20856,N_20925);
and U21188 (N_21188,N_20941,N_20695);
xor U21189 (N_21189,N_20887,N_20972);
or U21190 (N_21190,N_20616,N_20913);
xnor U21191 (N_21191,N_20860,N_20828);
nand U21192 (N_21192,N_20794,N_20767);
nand U21193 (N_21193,N_20631,N_20833);
nand U21194 (N_21194,N_20959,N_20721);
and U21195 (N_21195,N_20713,N_20841);
xor U21196 (N_21196,N_20699,N_20949);
and U21197 (N_21197,N_20653,N_20658);
and U21198 (N_21198,N_20831,N_20675);
nor U21199 (N_21199,N_20896,N_20756);
nor U21200 (N_21200,N_20663,N_20533);
and U21201 (N_21201,N_20657,N_20577);
and U21202 (N_21202,N_20891,N_20716);
and U21203 (N_21203,N_20938,N_20853);
and U21204 (N_21204,N_20873,N_20506);
and U21205 (N_21205,N_20910,N_20612);
and U21206 (N_21206,N_20882,N_20628);
xor U21207 (N_21207,N_20769,N_20746);
nand U21208 (N_21208,N_20945,N_20855);
or U21209 (N_21209,N_20578,N_20791);
nand U21210 (N_21210,N_20725,N_20918);
nor U21211 (N_21211,N_20999,N_20990);
nand U21212 (N_21212,N_20550,N_20928);
xnor U21213 (N_21213,N_20686,N_20715);
or U21214 (N_21214,N_20958,N_20744);
nor U21215 (N_21215,N_20706,N_20790);
and U21216 (N_21216,N_20942,N_20729);
or U21217 (N_21217,N_20762,N_20679);
or U21218 (N_21218,N_20576,N_20874);
xor U21219 (N_21219,N_20978,N_20570);
xor U21220 (N_21220,N_20633,N_20719);
xnor U21221 (N_21221,N_20711,N_20930);
nor U21222 (N_21222,N_20501,N_20800);
xor U21223 (N_21223,N_20777,N_20527);
nand U21224 (N_21224,N_20623,N_20535);
and U21225 (N_21225,N_20573,N_20889);
or U21226 (N_21226,N_20511,N_20502);
nand U21227 (N_21227,N_20780,N_20810);
or U21228 (N_21228,N_20809,N_20687);
nor U21229 (N_21229,N_20909,N_20761);
or U21230 (N_21230,N_20920,N_20807);
or U21231 (N_21231,N_20613,N_20805);
nand U21232 (N_21232,N_20643,N_20747);
and U21233 (N_21233,N_20798,N_20867);
nand U21234 (N_21234,N_20593,N_20552);
nor U21235 (N_21235,N_20902,N_20528);
or U21236 (N_21236,N_20921,N_20905);
nor U21237 (N_21237,N_20640,N_20854);
nand U21238 (N_21238,N_20994,N_20865);
xor U21239 (N_21239,N_20869,N_20758);
or U21240 (N_21240,N_20877,N_20917);
or U21241 (N_21241,N_20825,N_20862);
or U21242 (N_21242,N_20783,N_20583);
nand U21243 (N_21243,N_20842,N_20639);
nor U21244 (N_21244,N_20963,N_20571);
or U21245 (N_21245,N_20567,N_20802);
or U21246 (N_21246,N_20520,N_20671);
nor U21247 (N_21247,N_20526,N_20564);
nor U21248 (N_21248,N_20539,N_20979);
xor U21249 (N_21249,N_20812,N_20742);
nor U21250 (N_21250,N_20793,N_20955);
or U21251 (N_21251,N_20590,N_20705);
nand U21252 (N_21252,N_20923,N_20517);
xnor U21253 (N_21253,N_20537,N_20698);
nor U21254 (N_21254,N_20619,N_20604);
nor U21255 (N_21255,N_20631,N_20523);
nand U21256 (N_21256,N_20612,N_20883);
or U21257 (N_21257,N_20513,N_20638);
or U21258 (N_21258,N_20649,N_20606);
nor U21259 (N_21259,N_20875,N_20516);
and U21260 (N_21260,N_20762,N_20770);
xnor U21261 (N_21261,N_20994,N_20985);
nand U21262 (N_21262,N_20630,N_20896);
nor U21263 (N_21263,N_20990,N_20581);
nand U21264 (N_21264,N_20779,N_20759);
or U21265 (N_21265,N_20526,N_20579);
nor U21266 (N_21266,N_20645,N_20618);
xor U21267 (N_21267,N_20861,N_20825);
nor U21268 (N_21268,N_20665,N_20801);
and U21269 (N_21269,N_20788,N_20663);
or U21270 (N_21270,N_20512,N_20567);
xnor U21271 (N_21271,N_20903,N_20947);
or U21272 (N_21272,N_20554,N_20936);
and U21273 (N_21273,N_20835,N_20522);
or U21274 (N_21274,N_20998,N_20995);
and U21275 (N_21275,N_20969,N_20723);
nand U21276 (N_21276,N_20987,N_20996);
xnor U21277 (N_21277,N_20997,N_20909);
nand U21278 (N_21278,N_20699,N_20692);
xnor U21279 (N_21279,N_20978,N_20869);
nor U21280 (N_21280,N_20869,N_20648);
nor U21281 (N_21281,N_20590,N_20756);
xor U21282 (N_21282,N_20654,N_20760);
nand U21283 (N_21283,N_20933,N_20898);
and U21284 (N_21284,N_20749,N_20606);
and U21285 (N_21285,N_20943,N_20827);
nand U21286 (N_21286,N_20878,N_20753);
xnor U21287 (N_21287,N_20880,N_20560);
nor U21288 (N_21288,N_20945,N_20863);
nor U21289 (N_21289,N_20547,N_20646);
nand U21290 (N_21290,N_20680,N_20669);
nand U21291 (N_21291,N_20656,N_20892);
xnor U21292 (N_21292,N_20806,N_20801);
nor U21293 (N_21293,N_20750,N_20697);
and U21294 (N_21294,N_20959,N_20984);
or U21295 (N_21295,N_20959,N_20791);
and U21296 (N_21296,N_20920,N_20826);
nand U21297 (N_21297,N_20571,N_20781);
or U21298 (N_21298,N_20813,N_20629);
xor U21299 (N_21299,N_20627,N_20730);
nor U21300 (N_21300,N_20976,N_20547);
nor U21301 (N_21301,N_20889,N_20884);
xor U21302 (N_21302,N_20781,N_20861);
nor U21303 (N_21303,N_20866,N_20573);
nand U21304 (N_21304,N_20874,N_20926);
xor U21305 (N_21305,N_20862,N_20937);
or U21306 (N_21306,N_20684,N_20953);
or U21307 (N_21307,N_20670,N_20770);
and U21308 (N_21308,N_20947,N_20912);
nand U21309 (N_21309,N_20757,N_20930);
nor U21310 (N_21310,N_20580,N_20544);
nand U21311 (N_21311,N_20746,N_20814);
nand U21312 (N_21312,N_20873,N_20664);
nor U21313 (N_21313,N_20621,N_20779);
or U21314 (N_21314,N_20636,N_20699);
or U21315 (N_21315,N_20661,N_20888);
xor U21316 (N_21316,N_20742,N_20824);
and U21317 (N_21317,N_20862,N_20765);
nand U21318 (N_21318,N_20851,N_20776);
xnor U21319 (N_21319,N_20719,N_20607);
or U21320 (N_21320,N_20816,N_20706);
and U21321 (N_21321,N_20754,N_20685);
and U21322 (N_21322,N_20532,N_20950);
nor U21323 (N_21323,N_20809,N_20583);
nand U21324 (N_21324,N_20630,N_20573);
xnor U21325 (N_21325,N_20685,N_20913);
xnor U21326 (N_21326,N_20804,N_20731);
or U21327 (N_21327,N_20501,N_20903);
nand U21328 (N_21328,N_20860,N_20686);
nand U21329 (N_21329,N_20820,N_20937);
nor U21330 (N_21330,N_20639,N_20891);
xor U21331 (N_21331,N_20684,N_20753);
nor U21332 (N_21332,N_20890,N_20964);
nor U21333 (N_21333,N_20522,N_20847);
nand U21334 (N_21334,N_20801,N_20884);
xor U21335 (N_21335,N_20508,N_20818);
xor U21336 (N_21336,N_20668,N_20878);
and U21337 (N_21337,N_20925,N_20737);
and U21338 (N_21338,N_20517,N_20954);
nor U21339 (N_21339,N_20941,N_20889);
and U21340 (N_21340,N_20965,N_20594);
nor U21341 (N_21341,N_20780,N_20907);
nand U21342 (N_21342,N_20656,N_20798);
or U21343 (N_21343,N_20811,N_20806);
nand U21344 (N_21344,N_20753,N_20517);
and U21345 (N_21345,N_20766,N_20692);
xnor U21346 (N_21346,N_20590,N_20699);
xor U21347 (N_21347,N_20766,N_20511);
xnor U21348 (N_21348,N_20835,N_20662);
or U21349 (N_21349,N_20530,N_20554);
or U21350 (N_21350,N_20539,N_20559);
and U21351 (N_21351,N_20768,N_20856);
and U21352 (N_21352,N_20829,N_20798);
and U21353 (N_21353,N_20878,N_20800);
xnor U21354 (N_21354,N_20871,N_20817);
or U21355 (N_21355,N_20611,N_20842);
and U21356 (N_21356,N_20567,N_20866);
or U21357 (N_21357,N_20908,N_20521);
xnor U21358 (N_21358,N_20808,N_20670);
nor U21359 (N_21359,N_20516,N_20624);
nand U21360 (N_21360,N_20963,N_20759);
xor U21361 (N_21361,N_20693,N_20504);
and U21362 (N_21362,N_20961,N_20890);
nand U21363 (N_21363,N_20559,N_20872);
nand U21364 (N_21364,N_20763,N_20986);
and U21365 (N_21365,N_20534,N_20702);
or U21366 (N_21366,N_20922,N_20564);
and U21367 (N_21367,N_20593,N_20940);
or U21368 (N_21368,N_20526,N_20948);
and U21369 (N_21369,N_20685,N_20831);
nor U21370 (N_21370,N_20582,N_20808);
nand U21371 (N_21371,N_20864,N_20686);
xor U21372 (N_21372,N_20654,N_20900);
and U21373 (N_21373,N_20564,N_20991);
and U21374 (N_21374,N_20751,N_20841);
xnor U21375 (N_21375,N_20900,N_20835);
and U21376 (N_21376,N_20691,N_20827);
nor U21377 (N_21377,N_20856,N_20991);
and U21378 (N_21378,N_20621,N_20504);
xor U21379 (N_21379,N_20638,N_20806);
nor U21380 (N_21380,N_20771,N_20655);
or U21381 (N_21381,N_20640,N_20685);
nor U21382 (N_21382,N_20857,N_20946);
nand U21383 (N_21383,N_20776,N_20970);
and U21384 (N_21384,N_20890,N_20814);
nand U21385 (N_21385,N_20975,N_20804);
xnor U21386 (N_21386,N_20569,N_20890);
nand U21387 (N_21387,N_20765,N_20611);
or U21388 (N_21388,N_20915,N_20806);
or U21389 (N_21389,N_20764,N_20890);
xnor U21390 (N_21390,N_20931,N_20999);
or U21391 (N_21391,N_20794,N_20703);
and U21392 (N_21392,N_20520,N_20945);
xnor U21393 (N_21393,N_20781,N_20640);
xor U21394 (N_21394,N_20676,N_20955);
xnor U21395 (N_21395,N_20707,N_20502);
nor U21396 (N_21396,N_20964,N_20999);
and U21397 (N_21397,N_20549,N_20933);
nor U21398 (N_21398,N_20653,N_20963);
nand U21399 (N_21399,N_20922,N_20679);
xor U21400 (N_21400,N_20740,N_20824);
nand U21401 (N_21401,N_20796,N_20699);
xnor U21402 (N_21402,N_20785,N_20881);
nor U21403 (N_21403,N_20967,N_20847);
nand U21404 (N_21404,N_20950,N_20573);
xor U21405 (N_21405,N_20928,N_20833);
xnor U21406 (N_21406,N_20828,N_20600);
nand U21407 (N_21407,N_20955,N_20561);
or U21408 (N_21408,N_20687,N_20728);
nor U21409 (N_21409,N_20925,N_20903);
xor U21410 (N_21410,N_20980,N_20526);
or U21411 (N_21411,N_20905,N_20827);
nand U21412 (N_21412,N_20893,N_20797);
nand U21413 (N_21413,N_20907,N_20572);
or U21414 (N_21414,N_20851,N_20788);
and U21415 (N_21415,N_20730,N_20694);
xor U21416 (N_21416,N_20772,N_20514);
and U21417 (N_21417,N_20863,N_20546);
xor U21418 (N_21418,N_20769,N_20693);
and U21419 (N_21419,N_20749,N_20900);
or U21420 (N_21420,N_20804,N_20689);
or U21421 (N_21421,N_20827,N_20854);
and U21422 (N_21422,N_20673,N_20820);
xor U21423 (N_21423,N_20882,N_20790);
or U21424 (N_21424,N_20604,N_20959);
and U21425 (N_21425,N_20854,N_20868);
or U21426 (N_21426,N_20815,N_20977);
or U21427 (N_21427,N_20980,N_20550);
or U21428 (N_21428,N_20788,N_20580);
and U21429 (N_21429,N_20538,N_20831);
xnor U21430 (N_21430,N_20622,N_20914);
and U21431 (N_21431,N_20536,N_20901);
nand U21432 (N_21432,N_20869,N_20576);
nor U21433 (N_21433,N_20705,N_20638);
nor U21434 (N_21434,N_20863,N_20566);
nand U21435 (N_21435,N_20804,N_20524);
and U21436 (N_21436,N_20547,N_20552);
nand U21437 (N_21437,N_20762,N_20732);
nand U21438 (N_21438,N_20888,N_20696);
xnor U21439 (N_21439,N_20717,N_20820);
nor U21440 (N_21440,N_20771,N_20848);
nand U21441 (N_21441,N_20978,N_20703);
xor U21442 (N_21442,N_20856,N_20792);
and U21443 (N_21443,N_20888,N_20665);
xor U21444 (N_21444,N_20546,N_20559);
or U21445 (N_21445,N_20612,N_20943);
xor U21446 (N_21446,N_20623,N_20695);
nand U21447 (N_21447,N_20953,N_20780);
and U21448 (N_21448,N_20980,N_20865);
or U21449 (N_21449,N_20730,N_20509);
and U21450 (N_21450,N_20616,N_20583);
or U21451 (N_21451,N_20825,N_20800);
or U21452 (N_21452,N_20951,N_20665);
nand U21453 (N_21453,N_20701,N_20641);
nor U21454 (N_21454,N_20533,N_20924);
xor U21455 (N_21455,N_20773,N_20919);
and U21456 (N_21456,N_20796,N_20856);
xor U21457 (N_21457,N_20794,N_20640);
nand U21458 (N_21458,N_20702,N_20964);
and U21459 (N_21459,N_20541,N_20636);
or U21460 (N_21460,N_20814,N_20880);
nand U21461 (N_21461,N_20687,N_20846);
nor U21462 (N_21462,N_20635,N_20930);
and U21463 (N_21463,N_20909,N_20680);
xnor U21464 (N_21464,N_20825,N_20537);
xnor U21465 (N_21465,N_20694,N_20912);
nor U21466 (N_21466,N_20611,N_20708);
xor U21467 (N_21467,N_20541,N_20545);
and U21468 (N_21468,N_20819,N_20689);
nor U21469 (N_21469,N_20565,N_20716);
or U21470 (N_21470,N_20765,N_20671);
xor U21471 (N_21471,N_20909,N_20652);
nor U21472 (N_21472,N_20995,N_20534);
and U21473 (N_21473,N_20512,N_20888);
xnor U21474 (N_21474,N_20966,N_20944);
nor U21475 (N_21475,N_20822,N_20868);
and U21476 (N_21476,N_20998,N_20875);
xnor U21477 (N_21477,N_20660,N_20858);
xor U21478 (N_21478,N_20701,N_20554);
and U21479 (N_21479,N_20633,N_20877);
and U21480 (N_21480,N_20643,N_20715);
or U21481 (N_21481,N_20589,N_20583);
or U21482 (N_21482,N_20995,N_20504);
nor U21483 (N_21483,N_20798,N_20542);
or U21484 (N_21484,N_20576,N_20955);
xor U21485 (N_21485,N_20871,N_20749);
xor U21486 (N_21486,N_20639,N_20858);
xnor U21487 (N_21487,N_20675,N_20723);
xnor U21488 (N_21488,N_20926,N_20554);
and U21489 (N_21489,N_20535,N_20748);
nand U21490 (N_21490,N_20813,N_20677);
xnor U21491 (N_21491,N_20767,N_20550);
nor U21492 (N_21492,N_20879,N_20651);
and U21493 (N_21493,N_20942,N_20716);
xor U21494 (N_21494,N_20813,N_20697);
xnor U21495 (N_21495,N_20950,N_20759);
nor U21496 (N_21496,N_20948,N_20513);
and U21497 (N_21497,N_20743,N_20918);
or U21498 (N_21498,N_20961,N_20570);
nor U21499 (N_21499,N_20706,N_20909);
or U21500 (N_21500,N_21054,N_21391);
and U21501 (N_21501,N_21000,N_21324);
xor U21502 (N_21502,N_21295,N_21006);
or U21503 (N_21503,N_21291,N_21181);
nor U21504 (N_21504,N_21489,N_21029);
or U21505 (N_21505,N_21214,N_21436);
xor U21506 (N_21506,N_21071,N_21281);
nand U21507 (N_21507,N_21103,N_21338);
nand U21508 (N_21508,N_21130,N_21135);
nor U21509 (N_21509,N_21495,N_21067);
or U21510 (N_21510,N_21199,N_21139);
and U21511 (N_21511,N_21227,N_21266);
and U21512 (N_21512,N_21129,N_21403);
nand U21513 (N_21513,N_21346,N_21083);
nand U21514 (N_21514,N_21073,N_21142);
xnor U21515 (N_21515,N_21137,N_21268);
and U21516 (N_21516,N_21269,N_21310);
xor U21517 (N_21517,N_21074,N_21407);
and U21518 (N_21518,N_21461,N_21410);
and U21519 (N_21519,N_21069,N_21010);
or U21520 (N_21520,N_21233,N_21359);
nand U21521 (N_21521,N_21177,N_21123);
nand U21522 (N_21522,N_21134,N_21484);
or U21523 (N_21523,N_21307,N_21483);
or U21524 (N_21524,N_21144,N_21470);
xor U21525 (N_21525,N_21487,N_21302);
xnor U21526 (N_21526,N_21131,N_21229);
or U21527 (N_21527,N_21241,N_21235);
or U21528 (N_21528,N_21301,N_21476);
xor U21529 (N_21529,N_21136,N_21340);
nor U21530 (N_21530,N_21039,N_21044);
nor U21531 (N_21531,N_21242,N_21011);
or U21532 (N_21532,N_21122,N_21151);
or U21533 (N_21533,N_21368,N_21237);
and U21534 (N_21534,N_21018,N_21399);
xor U21535 (N_21535,N_21111,N_21325);
and U21536 (N_21536,N_21166,N_21202);
nand U21537 (N_21537,N_21027,N_21234);
or U21538 (N_21538,N_21100,N_21133);
nor U21539 (N_21539,N_21298,N_21249);
nand U21540 (N_21540,N_21285,N_21224);
nor U21541 (N_21541,N_21185,N_21005);
xor U21542 (N_21542,N_21211,N_21042);
and U21543 (N_21543,N_21183,N_21383);
nand U21544 (N_21544,N_21104,N_21426);
nor U21545 (N_21545,N_21366,N_21198);
or U21546 (N_21546,N_21394,N_21272);
nor U21547 (N_21547,N_21466,N_21221);
or U21548 (N_21548,N_21244,N_21112);
or U21549 (N_21549,N_21464,N_21297);
or U21550 (N_21550,N_21097,N_21070);
nor U21551 (N_21551,N_21363,N_21022);
xor U21552 (N_21552,N_21287,N_21016);
xnor U21553 (N_21553,N_21456,N_21396);
xnor U21554 (N_21554,N_21007,N_21335);
and U21555 (N_21555,N_21493,N_21056);
xnor U21556 (N_21556,N_21382,N_21173);
xor U21557 (N_21557,N_21036,N_21347);
nor U21558 (N_21558,N_21333,N_21274);
xnor U21559 (N_21559,N_21077,N_21430);
xnor U21560 (N_21560,N_21299,N_21480);
and U21561 (N_21561,N_21058,N_21253);
nor U21562 (N_21562,N_21465,N_21270);
and U21563 (N_21563,N_21479,N_21093);
xnor U21564 (N_21564,N_21095,N_21154);
nor U21565 (N_21565,N_21343,N_21446);
nand U21566 (N_21566,N_21348,N_21458);
nand U21567 (N_21567,N_21259,N_21362);
nand U21568 (N_21568,N_21425,N_21317);
or U21569 (N_21569,N_21390,N_21162);
xor U21570 (N_21570,N_21002,N_21024);
xnor U21571 (N_21571,N_21200,N_21176);
nand U21572 (N_21572,N_21048,N_21365);
or U21573 (N_21573,N_21388,N_21159);
nor U21574 (N_21574,N_21116,N_21296);
xnor U21575 (N_21575,N_21459,N_21252);
nor U21576 (N_21576,N_21157,N_21273);
nor U21577 (N_21577,N_21001,N_21078);
or U21578 (N_21578,N_21498,N_21276);
and U21579 (N_21579,N_21217,N_21125);
and U21580 (N_21580,N_21212,N_21098);
nand U21581 (N_21581,N_21127,N_21280);
or U21582 (N_21582,N_21258,N_21089);
nor U21583 (N_21583,N_21179,N_21444);
xnor U21584 (N_21584,N_21378,N_21328);
xnor U21585 (N_21585,N_21353,N_21230);
or U21586 (N_21586,N_21402,N_21424);
xnor U21587 (N_21587,N_21367,N_21423);
xnor U21588 (N_21588,N_21389,N_21087);
nor U21589 (N_21589,N_21254,N_21448);
and U21590 (N_21590,N_21114,N_21305);
and U21591 (N_21591,N_21192,N_21277);
nor U21592 (N_21592,N_21207,N_21439);
xor U21593 (N_21593,N_21020,N_21431);
and U21594 (N_21594,N_21197,N_21032);
or U21595 (N_21595,N_21442,N_21372);
nor U21596 (N_21596,N_21226,N_21477);
xor U21597 (N_21597,N_21409,N_21014);
xor U21598 (N_21598,N_21469,N_21437);
nor U21599 (N_21599,N_21380,N_21246);
and U21600 (N_21600,N_21395,N_21311);
or U21601 (N_21601,N_21398,N_21428);
nand U21602 (N_21602,N_21141,N_21326);
nor U21603 (N_21603,N_21393,N_21286);
or U21604 (N_21604,N_21496,N_21263);
and U21605 (N_21605,N_21164,N_21292);
and U21606 (N_21606,N_21228,N_21356);
or U21607 (N_21607,N_21499,N_21293);
or U21608 (N_21608,N_21206,N_21321);
and U21609 (N_21609,N_21243,N_21262);
nand U21610 (N_21610,N_21195,N_21117);
or U21611 (N_21611,N_21113,N_21490);
nor U21612 (N_21612,N_21432,N_21146);
or U21613 (N_21613,N_21445,N_21438);
nor U21614 (N_21614,N_21337,N_21386);
xnor U21615 (N_21615,N_21047,N_21161);
and U21616 (N_21616,N_21205,N_21012);
xnor U21617 (N_21617,N_21163,N_21289);
and U21618 (N_21618,N_21160,N_21349);
and U21619 (N_21619,N_21090,N_21381);
or U21620 (N_21620,N_21255,N_21031);
or U21621 (N_21621,N_21481,N_21482);
nand U21622 (N_21622,N_21354,N_21474);
nand U21623 (N_21623,N_21171,N_21015);
nand U21624 (N_21624,N_21057,N_21052);
nand U21625 (N_21625,N_21019,N_21434);
nand U21626 (N_21626,N_21413,N_21025);
nand U21627 (N_21627,N_21361,N_21066);
and U21628 (N_21628,N_21322,N_21061);
and U21629 (N_21629,N_21303,N_21441);
or U21630 (N_21630,N_21472,N_21216);
or U21631 (N_21631,N_21043,N_21455);
or U21632 (N_21632,N_21251,N_21486);
and U21633 (N_21633,N_21319,N_21419);
or U21634 (N_21634,N_21189,N_21165);
and U21635 (N_21635,N_21334,N_21318);
nand U21636 (N_21636,N_21473,N_21488);
and U21637 (N_21637,N_21172,N_21420);
or U21638 (N_21638,N_21284,N_21193);
or U21639 (N_21639,N_21449,N_21222);
nor U21640 (N_21640,N_21110,N_21312);
nand U21641 (N_21641,N_21106,N_21247);
nand U21642 (N_21642,N_21219,N_21101);
xnor U21643 (N_21643,N_21376,N_21148);
and U21644 (N_21644,N_21256,N_21352);
xor U21645 (N_21645,N_21119,N_21447);
xnor U21646 (N_21646,N_21497,N_21187);
xnor U21647 (N_21647,N_21421,N_21245);
xnor U21648 (N_21648,N_21308,N_21231);
xor U21649 (N_21649,N_21451,N_21055);
nand U21650 (N_21650,N_21264,N_21339);
or U21651 (N_21651,N_21492,N_21084);
nand U21652 (N_21652,N_21062,N_21405);
nor U21653 (N_21653,N_21115,N_21240);
nor U21654 (N_21654,N_21046,N_21275);
nor U21655 (N_21655,N_21204,N_21126);
nand U21656 (N_21656,N_21201,N_21467);
or U21657 (N_21657,N_21105,N_21485);
or U21658 (N_21658,N_21037,N_21118);
xnor U21659 (N_21659,N_21081,N_21279);
xnor U21660 (N_21660,N_21239,N_21267);
or U21661 (N_21661,N_21373,N_21099);
and U21662 (N_21662,N_21040,N_21294);
nor U21663 (N_21663,N_21411,N_21282);
nand U21664 (N_21664,N_21248,N_21316);
and U21665 (N_21665,N_21218,N_21250);
xor U21666 (N_21666,N_21153,N_21158);
nand U21667 (N_21667,N_21180,N_21360);
or U21668 (N_21668,N_21208,N_21491);
or U21669 (N_21669,N_21330,N_21190);
xor U21670 (N_21670,N_21320,N_21355);
nor U21671 (N_21671,N_21236,N_21082);
xor U21672 (N_21672,N_21375,N_21138);
nand U21673 (N_21673,N_21315,N_21418);
nand U21674 (N_21674,N_21124,N_21167);
nand U21675 (N_21675,N_21350,N_21152);
nor U21676 (N_21676,N_21435,N_21045);
and U21677 (N_21677,N_21345,N_21351);
nor U21678 (N_21678,N_21076,N_21306);
xnor U21679 (N_21679,N_21463,N_21327);
and U21680 (N_21680,N_21290,N_21049);
xor U21681 (N_21681,N_21102,N_21041);
or U21682 (N_21682,N_21028,N_21358);
nor U21683 (N_21683,N_21387,N_21030);
and U21684 (N_21684,N_21300,N_21026);
and U21685 (N_21685,N_21427,N_21401);
xor U21686 (N_21686,N_21143,N_21452);
and U21687 (N_21687,N_21288,N_21091);
nor U21688 (N_21688,N_21150,N_21120);
nand U21689 (N_21689,N_21009,N_21384);
or U21690 (N_21690,N_21203,N_21213);
or U21691 (N_21691,N_21433,N_21170);
and U21692 (N_21692,N_21454,N_21370);
nand U21693 (N_21693,N_21080,N_21008);
or U21694 (N_21694,N_21034,N_21379);
nor U21695 (N_21695,N_21475,N_21344);
nand U21696 (N_21696,N_21478,N_21086);
xnor U21697 (N_21697,N_21232,N_21023);
xor U21698 (N_21698,N_21323,N_21168);
or U21699 (N_21699,N_21050,N_21184);
nand U21700 (N_21700,N_21017,N_21149);
or U21701 (N_21701,N_21238,N_21404);
or U21702 (N_21702,N_21457,N_21013);
nor U21703 (N_21703,N_21471,N_21145);
nand U21704 (N_21704,N_21265,N_21147);
nand U21705 (N_21705,N_21053,N_21092);
or U21706 (N_21706,N_21215,N_21443);
or U21707 (N_21707,N_21156,N_21038);
or U21708 (N_21708,N_21068,N_21094);
and U21709 (N_21709,N_21453,N_21196);
xnor U21710 (N_21710,N_21175,N_21304);
and U21711 (N_21711,N_21096,N_21412);
nor U21712 (N_21712,N_21342,N_21085);
nor U21713 (N_21713,N_21064,N_21169);
nor U21714 (N_21714,N_21278,N_21257);
nor U21715 (N_21715,N_21035,N_21065);
and U21716 (N_21716,N_21440,N_21210);
xor U21717 (N_21717,N_21063,N_21406);
nand U21718 (N_21718,N_21072,N_21088);
and U21719 (N_21719,N_21108,N_21079);
nand U21720 (N_21720,N_21416,N_21132);
and U21721 (N_21721,N_21186,N_21174);
or U21722 (N_21722,N_21468,N_21225);
xor U21723 (N_21723,N_21429,N_21209);
nor U21724 (N_21724,N_21385,N_21331);
nor U21725 (N_21725,N_21462,N_21494);
nand U21726 (N_21726,N_21004,N_21060);
xnor U21727 (N_21727,N_21140,N_21357);
and U21728 (N_21728,N_21400,N_21450);
and U21729 (N_21729,N_21283,N_21314);
nor U21730 (N_21730,N_21408,N_21194);
nor U21731 (N_21731,N_21309,N_21332);
nor U21732 (N_21732,N_21377,N_21336);
and U21733 (N_21733,N_21341,N_21059);
and U21734 (N_21734,N_21414,N_21392);
and U21735 (N_21735,N_21397,N_21313);
nand U21736 (N_21736,N_21033,N_21107);
xnor U21737 (N_21737,N_21271,N_21220);
and U21738 (N_21738,N_21021,N_21075);
or U21739 (N_21739,N_21260,N_21374);
or U21740 (N_21740,N_21003,N_21178);
nor U21741 (N_21741,N_21191,N_21223);
or U21742 (N_21742,N_21109,N_21415);
or U21743 (N_21743,N_21371,N_21182);
nor U21744 (N_21744,N_21128,N_21422);
and U21745 (N_21745,N_21369,N_21188);
or U21746 (N_21746,N_21261,N_21051);
nand U21747 (N_21747,N_21460,N_21329);
and U21748 (N_21748,N_21364,N_21417);
nor U21749 (N_21749,N_21121,N_21155);
nor U21750 (N_21750,N_21334,N_21428);
or U21751 (N_21751,N_21369,N_21308);
nor U21752 (N_21752,N_21442,N_21054);
xor U21753 (N_21753,N_21087,N_21312);
nand U21754 (N_21754,N_21221,N_21013);
nor U21755 (N_21755,N_21399,N_21217);
nor U21756 (N_21756,N_21104,N_21090);
xnor U21757 (N_21757,N_21306,N_21185);
or U21758 (N_21758,N_21078,N_21405);
nor U21759 (N_21759,N_21329,N_21008);
and U21760 (N_21760,N_21301,N_21126);
nor U21761 (N_21761,N_21361,N_21200);
and U21762 (N_21762,N_21394,N_21192);
xor U21763 (N_21763,N_21112,N_21311);
or U21764 (N_21764,N_21353,N_21189);
nand U21765 (N_21765,N_21475,N_21095);
nor U21766 (N_21766,N_21381,N_21128);
xor U21767 (N_21767,N_21332,N_21471);
nand U21768 (N_21768,N_21191,N_21216);
nand U21769 (N_21769,N_21135,N_21459);
or U21770 (N_21770,N_21126,N_21007);
or U21771 (N_21771,N_21401,N_21334);
and U21772 (N_21772,N_21111,N_21387);
nand U21773 (N_21773,N_21064,N_21035);
xor U21774 (N_21774,N_21220,N_21295);
and U21775 (N_21775,N_21219,N_21479);
nand U21776 (N_21776,N_21058,N_21357);
or U21777 (N_21777,N_21056,N_21307);
xor U21778 (N_21778,N_21473,N_21230);
or U21779 (N_21779,N_21264,N_21097);
xnor U21780 (N_21780,N_21212,N_21211);
and U21781 (N_21781,N_21030,N_21009);
and U21782 (N_21782,N_21263,N_21296);
or U21783 (N_21783,N_21249,N_21007);
nor U21784 (N_21784,N_21142,N_21263);
nand U21785 (N_21785,N_21352,N_21298);
nor U21786 (N_21786,N_21000,N_21466);
or U21787 (N_21787,N_21092,N_21034);
or U21788 (N_21788,N_21175,N_21311);
nor U21789 (N_21789,N_21426,N_21090);
xnor U21790 (N_21790,N_21006,N_21113);
and U21791 (N_21791,N_21226,N_21358);
or U21792 (N_21792,N_21136,N_21130);
xor U21793 (N_21793,N_21034,N_21483);
xor U21794 (N_21794,N_21384,N_21045);
xnor U21795 (N_21795,N_21353,N_21297);
xnor U21796 (N_21796,N_21418,N_21185);
xnor U21797 (N_21797,N_21094,N_21294);
or U21798 (N_21798,N_21171,N_21289);
and U21799 (N_21799,N_21112,N_21193);
and U21800 (N_21800,N_21179,N_21082);
nand U21801 (N_21801,N_21081,N_21351);
nand U21802 (N_21802,N_21361,N_21318);
nor U21803 (N_21803,N_21412,N_21284);
and U21804 (N_21804,N_21302,N_21194);
or U21805 (N_21805,N_21264,N_21338);
or U21806 (N_21806,N_21212,N_21484);
xor U21807 (N_21807,N_21235,N_21151);
nand U21808 (N_21808,N_21210,N_21388);
nor U21809 (N_21809,N_21439,N_21129);
or U21810 (N_21810,N_21456,N_21000);
nor U21811 (N_21811,N_21204,N_21371);
and U21812 (N_21812,N_21103,N_21086);
or U21813 (N_21813,N_21070,N_21306);
nor U21814 (N_21814,N_21351,N_21342);
xor U21815 (N_21815,N_21013,N_21242);
nor U21816 (N_21816,N_21351,N_21461);
nand U21817 (N_21817,N_21332,N_21331);
xnor U21818 (N_21818,N_21021,N_21272);
nor U21819 (N_21819,N_21022,N_21297);
and U21820 (N_21820,N_21345,N_21310);
nand U21821 (N_21821,N_21153,N_21046);
nor U21822 (N_21822,N_21366,N_21056);
and U21823 (N_21823,N_21339,N_21128);
or U21824 (N_21824,N_21057,N_21453);
or U21825 (N_21825,N_21439,N_21117);
nor U21826 (N_21826,N_21343,N_21027);
nand U21827 (N_21827,N_21499,N_21010);
nand U21828 (N_21828,N_21351,N_21375);
or U21829 (N_21829,N_21240,N_21450);
xor U21830 (N_21830,N_21403,N_21061);
nor U21831 (N_21831,N_21262,N_21005);
nand U21832 (N_21832,N_21070,N_21418);
nor U21833 (N_21833,N_21248,N_21243);
and U21834 (N_21834,N_21472,N_21358);
xnor U21835 (N_21835,N_21006,N_21150);
xnor U21836 (N_21836,N_21199,N_21402);
xor U21837 (N_21837,N_21384,N_21265);
nor U21838 (N_21838,N_21447,N_21497);
xnor U21839 (N_21839,N_21211,N_21023);
and U21840 (N_21840,N_21022,N_21185);
nand U21841 (N_21841,N_21150,N_21032);
and U21842 (N_21842,N_21246,N_21290);
nand U21843 (N_21843,N_21151,N_21219);
nor U21844 (N_21844,N_21059,N_21410);
and U21845 (N_21845,N_21428,N_21189);
or U21846 (N_21846,N_21076,N_21130);
nor U21847 (N_21847,N_21374,N_21091);
and U21848 (N_21848,N_21125,N_21393);
and U21849 (N_21849,N_21377,N_21013);
xor U21850 (N_21850,N_21180,N_21389);
or U21851 (N_21851,N_21226,N_21414);
and U21852 (N_21852,N_21020,N_21081);
xor U21853 (N_21853,N_21151,N_21420);
or U21854 (N_21854,N_21453,N_21067);
and U21855 (N_21855,N_21408,N_21246);
and U21856 (N_21856,N_21417,N_21317);
xnor U21857 (N_21857,N_21006,N_21329);
nor U21858 (N_21858,N_21369,N_21410);
xnor U21859 (N_21859,N_21362,N_21325);
and U21860 (N_21860,N_21468,N_21114);
or U21861 (N_21861,N_21187,N_21383);
or U21862 (N_21862,N_21264,N_21310);
and U21863 (N_21863,N_21147,N_21149);
or U21864 (N_21864,N_21437,N_21083);
and U21865 (N_21865,N_21146,N_21354);
or U21866 (N_21866,N_21345,N_21095);
xnor U21867 (N_21867,N_21262,N_21213);
and U21868 (N_21868,N_21287,N_21002);
and U21869 (N_21869,N_21387,N_21357);
or U21870 (N_21870,N_21317,N_21150);
or U21871 (N_21871,N_21299,N_21297);
or U21872 (N_21872,N_21286,N_21223);
nand U21873 (N_21873,N_21332,N_21358);
or U21874 (N_21874,N_21148,N_21309);
and U21875 (N_21875,N_21148,N_21387);
or U21876 (N_21876,N_21066,N_21112);
nor U21877 (N_21877,N_21130,N_21047);
or U21878 (N_21878,N_21095,N_21145);
nor U21879 (N_21879,N_21420,N_21205);
and U21880 (N_21880,N_21257,N_21343);
nor U21881 (N_21881,N_21187,N_21287);
or U21882 (N_21882,N_21402,N_21117);
and U21883 (N_21883,N_21401,N_21372);
nor U21884 (N_21884,N_21108,N_21105);
and U21885 (N_21885,N_21490,N_21366);
or U21886 (N_21886,N_21242,N_21372);
nor U21887 (N_21887,N_21047,N_21395);
nor U21888 (N_21888,N_21382,N_21490);
nand U21889 (N_21889,N_21152,N_21384);
nor U21890 (N_21890,N_21315,N_21383);
nor U21891 (N_21891,N_21313,N_21201);
nand U21892 (N_21892,N_21272,N_21281);
nor U21893 (N_21893,N_21488,N_21190);
nand U21894 (N_21894,N_21016,N_21477);
and U21895 (N_21895,N_21173,N_21426);
xnor U21896 (N_21896,N_21287,N_21301);
nor U21897 (N_21897,N_21074,N_21423);
xnor U21898 (N_21898,N_21106,N_21205);
nand U21899 (N_21899,N_21184,N_21147);
nand U21900 (N_21900,N_21128,N_21434);
nor U21901 (N_21901,N_21478,N_21465);
nand U21902 (N_21902,N_21332,N_21038);
and U21903 (N_21903,N_21276,N_21267);
nor U21904 (N_21904,N_21285,N_21195);
or U21905 (N_21905,N_21199,N_21163);
nand U21906 (N_21906,N_21429,N_21339);
xor U21907 (N_21907,N_21397,N_21011);
nand U21908 (N_21908,N_21328,N_21460);
or U21909 (N_21909,N_21030,N_21210);
and U21910 (N_21910,N_21096,N_21133);
nor U21911 (N_21911,N_21019,N_21456);
nand U21912 (N_21912,N_21210,N_21016);
xnor U21913 (N_21913,N_21261,N_21016);
xor U21914 (N_21914,N_21285,N_21425);
xor U21915 (N_21915,N_21089,N_21233);
or U21916 (N_21916,N_21170,N_21139);
or U21917 (N_21917,N_21190,N_21007);
and U21918 (N_21918,N_21454,N_21453);
nor U21919 (N_21919,N_21284,N_21088);
and U21920 (N_21920,N_21209,N_21106);
nand U21921 (N_21921,N_21162,N_21408);
nand U21922 (N_21922,N_21363,N_21291);
nand U21923 (N_21923,N_21067,N_21172);
nand U21924 (N_21924,N_21224,N_21136);
or U21925 (N_21925,N_21171,N_21269);
nor U21926 (N_21926,N_21205,N_21208);
xnor U21927 (N_21927,N_21217,N_21434);
xnor U21928 (N_21928,N_21160,N_21461);
nand U21929 (N_21929,N_21375,N_21423);
xnor U21930 (N_21930,N_21049,N_21175);
nand U21931 (N_21931,N_21329,N_21022);
nor U21932 (N_21932,N_21448,N_21133);
nor U21933 (N_21933,N_21042,N_21083);
nand U21934 (N_21934,N_21397,N_21216);
or U21935 (N_21935,N_21316,N_21036);
and U21936 (N_21936,N_21257,N_21441);
xnor U21937 (N_21937,N_21028,N_21094);
nor U21938 (N_21938,N_21049,N_21384);
and U21939 (N_21939,N_21065,N_21095);
or U21940 (N_21940,N_21029,N_21203);
nor U21941 (N_21941,N_21116,N_21173);
or U21942 (N_21942,N_21129,N_21134);
nor U21943 (N_21943,N_21119,N_21356);
and U21944 (N_21944,N_21227,N_21040);
nand U21945 (N_21945,N_21449,N_21253);
nand U21946 (N_21946,N_21338,N_21486);
or U21947 (N_21947,N_21173,N_21225);
nand U21948 (N_21948,N_21354,N_21488);
xnor U21949 (N_21949,N_21335,N_21126);
nand U21950 (N_21950,N_21298,N_21308);
nand U21951 (N_21951,N_21131,N_21482);
xnor U21952 (N_21952,N_21157,N_21051);
and U21953 (N_21953,N_21171,N_21038);
or U21954 (N_21954,N_21265,N_21104);
xor U21955 (N_21955,N_21208,N_21376);
and U21956 (N_21956,N_21078,N_21455);
or U21957 (N_21957,N_21465,N_21359);
xor U21958 (N_21958,N_21337,N_21235);
or U21959 (N_21959,N_21181,N_21183);
or U21960 (N_21960,N_21460,N_21092);
nor U21961 (N_21961,N_21249,N_21494);
xor U21962 (N_21962,N_21443,N_21074);
nand U21963 (N_21963,N_21211,N_21137);
and U21964 (N_21964,N_21175,N_21313);
or U21965 (N_21965,N_21320,N_21306);
nand U21966 (N_21966,N_21062,N_21058);
or U21967 (N_21967,N_21247,N_21092);
or U21968 (N_21968,N_21372,N_21342);
nand U21969 (N_21969,N_21401,N_21320);
and U21970 (N_21970,N_21469,N_21162);
xnor U21971 (N_21971,N_21232,N_21391);
nor U21972 (N_21972,N_21017,N_21246);
or U21973 (N_21973,N_21126,N_21462);
nand U21974 (N_21974,N_21477,N_21182);
nor U21975 (N_21975,N_21175,N_21366);
or U21976 (N_21976,N_21217,N_21440);
and U21977 (N_21977,N_21219,N_21301);
xnor U21978 (N_21978,N_21443,N_21157);
and U21979 (N_21979,N_21356,N_21114);
xnor U21980 (N_21980,N_21400,N_21360);
or U21981 (N_21981,N_21489,N_21390);
nand U21982 (N_21982,N_21241,N_21183);
xnor U21983 (N_21983,N_21093,N_21484);
or U21984 (N_21984,N_21469,N_21149);
or U21985 (N_21985,N_21046,N_21491);
nand U21986 (N_21986,N_21022,N_21271);
xor U21987 (N_21987,N_21409,N_21038);
nor U21988 (N_21988,N_21304,N_21408);
or U21989 (N_21989,N_21023,N_21273);
or U21990 (N_21990,N_21408,N_21133);
xor U21991 (N_21991,N_21467,N_21244);
and U21992 (N_21992,N_21118,N_21031);
nand U21993 (N_21993,N_21322,N_21050);
xor U21994 (N_21994,N_21203,N_21138);
nor U21995 (N_21995,N_21096,N_21376);
and U21996 (N_21996,N_21447,N_21015);
or U21997 (N_21997,N_21465,N_21378);
and U21998 (N_21998,N_21493,N_21440);
nor U21999 (N_21999,N_21395,N_21238);
nor U22000 (N_22000,N_21756,N_21922);
nand U22001 (N_22001,N_21744,N_21851);
nor U22002 (N_22002,N_21545,N_21547);
nor U22003 (N_22003,N_21674,N_21880);
nor U22004 (N_22004,N_21883,N_21646);
or U22005 (N_22005,N_21732,N_21524);
xnor U22006 (N_22006,N_21997,N_21872);
xnor U22007 (N_22007,N_21560,N_21840);
nand U22008 (N_22008,N_21553,N_21668);
xor U22009 (N_22009,N_21625,N_21613);
nand U22010 (N_22010,N_21643,N_21861);
xnor U22011 (N_22011,N_21768,N_21663);
nor U22012 (N_22012,N_21957,N_21666);
nor U22013 (N_22013,N_21822,N_21517);
or U22014 (N_22014,N_21838,N_21915);
nand U22015 (N_22015,N_21817,N_21600);
xor U22016 (N_22016,N_21672,N_21877);
xnor U22017 (N_22017,N_21991,N_21684);
or U22018 (N_22018,N_21729,N_21692);
or U22019 (N_22019,N_21733,N_21626);
or U22020 (N_22020,N_21814,N_21824);
and U22021 (N_22021,N_21942,N_21725);
or U22022 (N_22022,N_21970,N_21763);
nand U22023 (N_22023,N_21783,N_21933);
nor U22024 (N_22024,N_21774,N_21571);
xnor U22025 (N_22025,N_21850,N_21607);
xnor U22026 (N_22026,N_21809,N_21631);
xnor U22027 (N_22027,N_21644,N_21971);
and U22028 (N_22028,N_21939,N_21538);
or U22029 (N_22029,N_21887,N_21727);
nand U22030 (N_22030,N_21864,N_21515);
and U22031 (N_22031,N_21664,N_21582);
xnor U22032 (N_22032,N_21953,N_21717);
nor U22033 (N_22033,N_21540,N_21926);
and U22034 (N_22034,N_21941,N_21779);
nand U22035 (N_22035,N_21669,N_21742);
and U22036 (N_22036,N_21903,N_21653);
xor U22037 (N_22037,N_21583,N_21645);
xnor U22038 (N_22038,N_21514,N_21748);
and U22039 (N_22039,N_21827,N_21771);
nor U22040 (N_22040,N_21906,N_21740);
or U22041 (N_22041,N_21723,N_21776);
and U22042 (N_22042,N_21982,N_21893);
xor U22043 (N_22043,N_21879,N_21534);
nor U22044 (N_22044,N_21966,N_21686);
nor U22045 (N_22045,N_21843,N_21705);
nor U22046 (N_22046,N_21988,N_21777);
nor U22047 (N_22047,N_21633,N_21753);
nor U22048 (N_22048,N_21846,N_21802);
nor U22049 (N_22049,N_21696,N_21619);
xnor U22050 (N_22050,N_21932,N_21782);
and U22051 (N_22051,N_21617,N_21606);
nand U22052 (N_22052,N_21876,N_21701);
nand U22053 (N_22053,N_21572,N_21722);
and U22054 (N_22054,N_21813,N_21761);
or U22055 (N_22055,N_21847,N_21637);
nor U22056 (N_22056,N_21839,N_21720);
xor U22057 (N_22057,N_21676,N_21825);
nor U22058 (N_22058,N_21781,N_21796);
and U22059 (N_22059,N_21741,N_21652);
nand U22060 (N_22060,N_21591,N_21803);
nand U22061 (N_22061,N_21946,N_21909);
nand U22062 (N_22062,N_21897,N_21757);
nand U22063 (N_22063,N_21875,N_21972);
and U22064 (N_22064,N_21918,N_21518);
nand U22065 (N_22065,N_21986,N_21920);
or U22066 (N_22066,N_21863,N_21649);
nor U22067 (N_22067,N_21921,N_21647);
xor U22068 (N_22068,N_21690,N_21566);
xor U22069 (N_22069,N_21913,N_21573);
nor U22070 (N_22070,N_21831,N_21820);
nor U22071 (N_22071,N_21541,N_21948);
or U22072 (N_22072,N_21816,N_21849);
nor U22073 (N_22073,N_21503,N_21818);
nor U22074 (N_22074,N_21501,N_21700);
nand U22075 (N_22075,N_21602,N_21559);
xnor U22076 (N_22076,N_21955,N_21789);
or U22077 (N_22077,N_21629,N_21958);
xnor U22078 (N_22078,N_21520,N_21737);
xnor U22079 (N_22079,N_21574,N_21975);
xor U22080 (N_22080,N_21616,N_21758);
and U22081 (N_22081,N_21892,N_21799);
xor U22082 (N_22082,N_21807,N_21521);
xor U22083 (N_22083,N_21829,N_21959);
or U22084 (N_22084,N_21550,N_21685);
nand U22085 (N_22085,N_21739,N_21707);
nor U22086 (N_22086,N_21806,N_21578);
and U22087 (N_22087,N_21724,N_21904);
xor U22088 (N_22088,N_21551,N_21624);
and U22089 (N_22089,N_21593,N_21750);
nand U22090 (N_22090,N_21568,N_21506);
nor U22091 (N_22091,N_21882,N_21622);
and U22092 (N_22092,N_21712,N_21589);
or U22093 (N_22093,N_21635,N_21665);
and U22094 (N_22094,N_21539,N_21549);
and U22095 (N_22095,N_21938,N_21638);
nand U22096 (N_22096,N_21931,N_21639);
nand U22097 (N_22097,N_21759,N_21730);
nor U22098 (N_22098,N_21798,N_21603);
or U22099 (N_22099,N_21765,N_21576);
or U22100 (N_22100,N_21710,N_21731);
or U22101 (N_22101,N_21532,N_21556);
and U22102 (N_22102,N_21785,N_21661);
and U22103 (N_22103,N_21592,N_21841);
or U22104 (N_22104,N_21721,N_21516);
nand U22105 (N_22105,N_21580,N_21762);
nor U22106 (N_22106,N_21916,N_21734);
nor U22107 (N_22107,N_21670,N_21680);
or U22108 (N_22108,N_21659,N_21570);
or U22109 (N_22109,N_21735,N_21947);
xnor U22110 (N_22110,N_21977,N_21787);
and U22111 (N_22111,N_21969,N_21956);
nand U22112 (N_22112,N_21963,N_21858);
xnor U22113 (N_22113,N_21702,N_21962);
or U22114 (N_22114,N_21967,N_21558);
nand U22115 (N_22115,N_21775,N_21786);
and U22116 (N_22116,N_21844,N_21888);
xnor U22117 (N_22117,N_21862,N_21585);
nor U22118 (N_22118,N_21992,N_21793);
nand U22119 (N_22119,N_21673,N_21527);
nand U22120 (N_22120,N_21509,N_21715);
and U22121 (N_22121,N_21687,N_21682);
xor U22122 (N_22122,N_21679,N_21642);
xnor U22123 (N_22123,N_21905,N_21927);
and U22124 (N_22124,N_21562,N_21934);
and U22125 (N_22125,N_21743,N_21859);
nor U22126 (N_22126,N_21772,N_21749);
nand U22127 (N_22127,N_21978,N_21819);
nand U22128 (N_22128,N_21821,N_21792);
nand U22129 (N_22129,N_21899,N_21608);
and U22130 (N_22130,N_21990,N_21878);
and U22131 (N_22131,N_21908,N_21854);
and U22132 (N_22132,N_21584,N_21885);
nor U22133 (N_22133,N_21871,N_21699);
xor U22134 (N_22134,N_21678,N_21598);
xnor U22135 (N_22135,N_21627,N_21675);
nand U22136 (N_22136,N_21836,N_21853);
or U22137 (N_22137,N_21718,N_21565);
and U22138 (N_22138,N_21693,N_21577);
or U22139 (N_22139,N_21529,N_21830);
nor U22140 (N_22140,N_21979,N_21508);
xnor U22141 (N_22141,N_21581,N_21755);
nor U22142 (N_22142,N_21900,N_21834);
nand U22143 (N_22143,N_21531,N_21930);
xnor U22144 (N_22144,N_21944,N_21528);
xnor U22145 (N_22145,N_21951,N_21695);
xnor U22146 (N_22146,N_21995,N_21703);
nand U22147 (N_22147,N_21985,N_21569);
nand U22148 (N_22148,N_21597,N_21842);
xnor U22149 (N_22149,N_21848,N_21736);
and U22150 (N_22150,N_21869,N_21530);
or U22151 (N_22151,N_21780,N_21891);
nand U22152 (N_22152,N_21615,N_21697);
nor U22153 (N_22153,N_21586,N_21974);
and U22154 (N_22154,N_21950,N_21940);
nand U22155 (N_22155,N_21949,N_21898);
nor U22156 (N_22156,N_21901,N_21914);
xor U22157 (N_22157,N_21812,N_21655);
nand U22158 (N_22158,N_21605,N_21618);
xnor U22159 (N_22159,N_21594,N_21552);
nand U22160 (N_22160,N_21925,N_21567);
and U22161 (N_22161,N_21533,N_21996);
nor U22162 (N_22162,N_21620,N_21691);
or U22163 (N_22163,N_21614,N_21632);
or U22164 (N_22164,N_21512,N_21952);
nand U22165 (N_22165,N_21714,N_21601);
nand U22166 (N_22166,N_21865,N_21561);
and U22167 (N_22167,N_21505,N_21630);
and U22168 (N_22168,N_21706,N_21935);
xor U22169 (N_22169,N_21596,N_21965);
xor U22170 (N_22170,N_21579,N_21535);
xnor U22171 (N_22171,N_21555,N_21747);
xnor U22172 (N_22172,N_21791,N_21987);
or U22173 (N_22173,N_21945,N_21677);
and U22174 (N_22174,N_21778,N_21658);
or U22175 (N_22175,N_21867,N_21623);
and U22176 (N_22176,N_21890,N_21857);
nand U22177 (N_22177,N_21751,N_21800);
nand U22178 (N_22178,N_21640,N_21689);
and U22179 (N_22179,N_21557,N_21548);
nand U22180 (N_22180,N_21587,N_21968);
and U22181 (N_22181,N_21896,N_21683);
xnor U22182 (N_22182,N_21808,N_21745);
and U22183 (N_22183,N_21788,N_21973);
nor U22184 (N_22184,N_21911,N_21954);
and U22185 (N_22185,N_21797,N_21998);
xor U22186 (N_22186,N_21924,N_21575);
nand U22187 (N_22187,N_21826,N_21886);
or U22188 (N_22188,N_21976,N_21599);
and U22189 (N_22189,N_21636,N_21804);
nand U22190 (N_22190,N_21828,N_21989);
or U22191 (N_22191,N_21855,N_21912);
nand U22192 (N_22192,N_21667,N_21544);
or U22193 (N_22193,N_21654,N_21656);
or U22194 (N_22194,N_21500,N_21960);
and U22195 (N_22195,N_21523,N_21917);
xnor U22196 (N_22196,N_21907,N_21889);
nor U22197 (N_22197,N_21815,N_21525);
nand U22198 (N_22198,N_21766,N_21628);
nand U22199 (N_22199,N_21641,N_21704);
nor U22200 (N_22200,N_21852,N_21590);
or U22201 (N_22201,N_21764,N_21713);
nand U22202 (N_22202,N_21564,N_21651);
nor U22203 (N_22203,N_21502,N_21794);
nand U22204 (N_22204,N_21795,N_21964);
nand U22205 (N_22205,N_21719,N_21770);
and U22206 (N_22206,N_21536,N_21919);
nor U22207 (N_22207,N_21981,N_21522);
xnor U22208 (N_22208,N_21688,N_21928);
and U22209 (N_22209,N_21833,N_21621);
xnor U22210 (N_22210,N_21961,N_21769);
xor U22211 (N_22211,N_21983,N_21728);
or U22212 (N_22212,N_21588,N_21860);
nor U22213 (N_22213,N_21543,N_21546);
xnor U22214 (N_22214,N_21595,N_21610);
and U22215 (N_22215,N_21835,N_21856);
nor U22216 (N_22216,N_21870,N_21910);
or U22217 (N_22217,N_21604,N_21511);
and U22218 (N_22218,N_21754,N_21716);
and U22219 (N_22219,N_21648,N_21510);
nor U22220 (N_22220,N_21513,N_21752);
xor U22221 (N_22221,N_21563,N_21837);
xnor U22222 (N_22222,N_21507,N_21760);
nor U22223 (N_22223,N_21832,N_21810);
xor U22224 (N_22224,N_21519,N_21980);
xor U22225 (N_22225,N_21504,N_21650);
xnor U22226 (N_22226,N_21537,N_21554);
xor U22227 (N_22227,N_21866,N_21611);
or U22228 (N_22228,N_21868,N_21923);
xnor U22229 (N_22229,N_21784,N_21694);
or U22230 (N_22230,N_21811,N_21999);
or U22231 (N_22231,N_21936,N_21657);
or U22232 (N_22232,N_21708,N_21609);
xnor U22233 (N_22233,N_21767,N_21895);
xor U22234 (N_22234,N_21823,N_21681);
and U22235 (N_22235,N_21902,N_21612);
nand U22236 (N_22236,N_21874,N_21805);
xor U22237 (N_22237,N_21801,N_21711);
nand U22238 (N_22238,N_21773,N_21634);
and U22239 (N_22239,N_21660,N_21845);
xnor U22240 (N_22240,N_21746,N_21937);
or U22241 (N_22241,N_21709,N_21726);
or U22242 (N_22242,N_21526,N_21929);
nand U22243 (N_22243,N_21881,N_21993);
and U22244 (N_22244,N_21884,N_21662);
nor U22245 (N_22245,N_21994,N_21790);
xor U22246 (N_22246,N_21698,N_21943);
or U22247 (N_22247,N_21894,N_21873);
or U22248 (N_22248,N_21984,N_21542);
nor U22249 (N_22249,N_21671,N_21738);
nand U22250 (N_22250,N_21614,N_21808);
nor U22251 (N_22251,N_21671,N_21565);
and U22252 (N_22252,N_21510,N_21740);
nor U22253 (N_22253,N_21920,N_21747);
nor U22254 (N_22254,N_21605,N_21533);
or U22255 (N_22255,N_21670,N_21737);
xor U22256 (N_22256,N_21894,N_21532);
nor U22257 (N_22257,N_21936,N_21765);
and U22258 (N_22258,N_21850,N_21899);
xor U22259 (N_22259,N_21566,N_21782);
and U22260 (N_22260,N_21739,N_21919);
nor U22261 (N_22261,N_21503,N_21764);
xnor U22262 (N_22262,N_21763,N_21809);
and U22263 (N_22263,N_21577,N_21509);
and U22264 (N_22264,N_21598,N_21808);
nand U22265 (N_22265,N_21515,N_21740);
or U22266 (N_22266,N_21812,N_21578);
xnor U22267 (N_22267,N_21611,N_21680);
nand U22268 (N_22268,N_21792,N_21545);
xnor U22269 (N_22269,N_21830,N_21644);
xnor U22270 (N_22270,N_21819,N_21839);
xor U22271 (N_22271,N_21875,N_21934);
xor U22272 (N_22272,N_21726,N_21559);
or U22273 (N_22273,N_21665,N_21594);
nand U22274 (N_22274,N_21942,N_21565);
or U22275 (N_22275,N_21912,N_21798);
and U22276 (N_22276,N_21931,N_21820);
nor U22277 (N_22277,N_21661,N_21595);
and U22278 (N_22278,N_21975,N_21934);
nand U22279 (N_22279,N_21779,N_21511);
nor U22280 (N_22280,N_21863,N_21509);
and U22281 (N_22281,N_21839,N_21627);
and U22282 (N_22282,N_21922,N_21561);
and U22283 (N_22283,N_21951,N_21644);
nor U22284 (N_22284,N_21596,N_21631);
xor U22285 (N_22285,N_21950,N_21574);
or U22286 (N_22286,N_21542,N_21624);
nand U22287 (N_22287,N_21600,N_21782);
or U22288 (N_22288,N_21847,N_21981);
or U22289 (N_22289,N_21523,N_21673);
or U22290 (N_22290,N_21500,N_21528);
and U22291 (N_22291,N_21771,N_21789);
nand U22292 (N_22292,N_21623,N_21567);
or U22293 (N_22293,N_21809,N_21812);
or U22294 (N_22294,N_21591,N_21739);
xor U22295 (N_22295,N_21607,N_21803);
xnor U22296 (N_22296,N_21513,N_21594);
xor U22297 (N_22297,N_21577,N_21674);
nor U22298 (N_22298,N_21566,N_21965);
or U22299 (N_22299,N_21689,N_21508);
nand U22300 (N_22300,N_21827,N_21510);
nand U22301 (N_22301,N_21629,N_21658);
nor U22302 (N_22302,N_21797,N_21875);
nand U22303 (N_22303,N_21993,N_21995);
or U22304 (N_22304,N_21625,N_21538);
nand U22305 (N_22305,N_21812,N_21752);
nand U22306 (N_22306,N_21535,N_21768);
or U22307 (N_22307,N_21923,N_21700);
or U22308 (N_22308,N_21874,N_21979);
xnor U22309 (N_22309,N_21500,N_21876);
nor U22310 (N_22310,N_21642,N_21566);
nand U22311 (N_22311,N_21597,N_21721);
nand U22312 (N_22312,N_21814,N_21686);
or U22313 (N_22313,N_21605,N_21543);
nand U22314 (N_22314,N_21782,N_21772);
nand U22315 (N_22315,N_21601,N_21982);
nand U22316 (N_22316,N_21752,N_21930);
and U22317 (N_22317,N_21975,N_21768);
and U22318 (N_22318,N_21861,N_21591);
xnor U22319 (N_22319,N_21681,N_21818);
and U22320 (N_22320,N_21923,N_21637);
nand U22321 (N_22321,N_21575,N_21838);
nand U22322 (N_22322,N_21737,N_21642);
or U22323 (N_22323,N_21906,N_21549);
or U22324 (N_22324,N_21997,N_21904);
and U22325 (N_22325,N_21906,N_21675);
and U22326 (N_22326,N_21661,N_21540);
and U22327 (N_22327,N_21754,N_21968);
or U22328 (N_22328,N_21782,N_21896);
or U22329 (N_22329,N_21916,N_21942);
nand U22330 (N_22330,N_21767,N_21905);
or U22331 (N_22331,N_21982,N_21653);
and U22332 (N_22332,N_21867,N_21576);
and U22333 (N_22333,N_21818,N_21600);
and U22334 (N_22334,N_21838,N_21730);
or U22335 (N_22335,N_21509,N_21524);
nand U22336 (N_22336,N_21932,N_21599);
and U22337 (N_22337,N_21786,N_21826);
xor U22338 (N_22338,N_21648,N_21921);
and U22339 (N_22339,N_21932,N_21825);
nand U22340 (N_22340,N_21920,N_21850);
and U22341 (N_22341,N_21767,N_21760);
and U22342 (N_22342,N_21551,N_21679);
or U22343 (N_22343,N_21641,N_21593);
or U22344 (N_22344,N_21603,N_21639);
nand U22345 (N_22345,N_21503,N_21602);
xor U22346 (N_22346,N_21649,N_21639);
xor U22347 (N_22347,N_21764,N_21564);
nor U22348 (N_22348,N_21792,N_21772);
or U22349 (N_22349,N_21798,N_21591);
xnor U22350 (N_22350,N_21818,N_21743);
and U22351 (N_22351,N_21962,N_21663);
nor U22352 (N_22352,N_21997,N_21894);
and U22353 (N_22353,N_21914,N_21934);
and U22354 (N_22354,N_21989,N_21768);
and U22355 (N_22355,N_21712,N_21757);
nor U22356 (N_22356,N_21865,N_21721);
nor U22357 (N_22357,N_21582,N_21948);
nor U22358 (N_22358,N_21600,N_21833);
nand U22359 (N_22359,N_21694,N_21958);
and U22360 (N_22360,N_21575,N_21510);
and U22361 (N_22361,N_21928,N_21792);
nor U22362 (N_22362,N_21815,N_21654);
and U22363 (N_22363,N_21848,N_21815);
nand U22364 (N_22364,N_21500,N_21956);
or U22365 (N_22365,N_21805,N_21716);
xnor U22366 (N_22366,N_21942,N_21987);
and U22367 (N_22367,N_21853,N_21561);
or U22368 (N_22368,N_21599,N_21809);
nor U22369 (N_22369,N_21703,N_21940);
or U22370 (N_22370,N_21926,N_21778);
xnor U22371 (N_22371,N_21588,N_21721);
or U22372 (N_22372,N_21542,N_21902);
xnor U22373 (N_22373,N_21835,N_21560);
or U22374 (N_22374,N_21591,N_21661);
xnor U22375 (N_22375,N_21584,N_21550);
or U22376 (N_22376,N_21679,N_21985);
and U22377 (N_22377,N_21885,N_21684);
nor U22378 (N_22378,N_21806,N_21853);
or U22379 (N_22379,N_21743,N_21967);
and U22380 (N_22380,N_21665,N_21781);
or U22381 (N_22381,N_21822,N_21562);
or U22382 (N_22382,N_21908,N_21655);
xor U22383 (N_22383,N_21668,N_21628);
xnor U22384 (N_22384,N_21698,N_21860);
or U22385 (N_22385,N_21973,N_21946);
nand U22386 (N_22386,N_21927,N_21714);
or U22387 (N_22387,N_21849,N_21564);
or U22388 (N_22388,N_21879,N_21934);
nand U22389 (N_22389,N_21654,N_21863);
nand U22390 (N_22390,N_21594,N_21704);
and U22391 (N_22391,N_21623,N_21751);
and U22392 (N_22392,N_21653,N_21829);
nand U22393 (N_22393,N_21864,N_21821);
and U22394 (N_22394,N_21796,N_21869);
nand U22395 (N_22395,N_21616,N_21605);
nor U22396 (N_22396,N_21929,N_21979);
or U22397 (N_22397,N_21519,N_21586);
nor U22398 (N_22398,N_21922,N_21527);
and U22399 (N_22399,N_21508,N_21770);
nand U22400 (N_22400,N_21616,N_21939);
nand U22401 (N_22401,N_21644,N_21932);
nor U22402 (N_22402,N_21592,N_21518);
nor U22403 (N_22403,N_21987,N_21781);
xor U22404 (N_22404,N_21765,N_21753);
nand U22405 (N_22405,N_21928,N_21938);
nor U22406 (N_22406,N_21932,N_21632);
nor U22407 (N_22407,N_21857,N_21838);
nand U22408 (N_22408,N_21974,N_21567);
nand U22409 (N_22409,N_21844,N_21982);
or U22410 (N_22410,N_21751,N_21820);
xnor U22411 (N_22411,N_21620,N_21582);
or U22412 (N_22412,N_21751,N_21567);
xor U22413 (N_22413,N_21754,N_21554);
and U22414 (N_22414,N_21918,N_21627);
xnor U22415 (N_22415,N_21753,N_21728);
nor U22416 (N_22416,N_21638,N_21907);
nand U22417 (N_22417,N_21971,N_21585);
xnor U22418 (N_22418,N_21715,N_21567);
xor U22419 (N_22419,N_21888,N_21548);
and U22420 (N_22420,N_21795,N_21502);
or U22421 (N_22421,N_21605,N_21798);
xnor U22422 (N_22422,N_21605,N_21728);
and U22423 (N_22423,N_21997,N_21639);
nand U22424 (N_22424,N_21845,N_21818);
nor U22425 (N_22425,N_21806,N_21744);
nor U22426 (N_22426,N_21866,N_21689);
nor U22427 (N_22427,N_21680,N_21840);
or U22428 (N_22428,N_21860,N_21803);
nor U22429 (N_22429,N_21858,N_21747);
or U22430 (N_22430,N_21708,N_21884);
or U22431 (N_22431,N_21752,N_21528);
xnor U22432 (N_22432,N_21649,N_21599);
nor U22433 (N_22433,N_21614,N_21899);
nor U22434 (N_22434,N_21549,N_21810);
or U22435 (N_22435,N_21806,N_21766);
or U22436 (N_22436,N_21776,N_21500);
nor U22437 (N_22437,N_21552,N_21586);
and U22438 (N_22438,N_21758,N_21781);
nor U22439 (N_22439,N_21911,N_21566);
xnor U22440 (N_22440,N_21860,N_21768);
or U22441 (N_22441,N_21690,N_21950);
nor U22442 (N_22442,N_21829,N_21918);
and U22443 (N_22443,N_21890,N_21911);
xor U22444 (N_22444,N_21845,N_21526);
or U22445 (N_22445,N_21830,N_21787);
and U22446 (N_22446,N_21589,N_21754);
nand U22447 (N_22447,N_21612,N_21778);
and U22448 (N_22448,N_21533,N_21685);
nor U22449 (N_22449,N_21595,N_21854);
nand U22450 (N_22450,N_21930,N_21674);
nand U22451 (N_22451,N_21568,N_21917);
nand U22452 (N_22452,N_21738,N_21928);
xor U22453 (N_22453,N_21626,N_21680);
nor U22454 (N_22454,N_21757,N_21763);
nor U22455 (N_22455,N_21980,N_21836);
or U22456 (N_22456,N_21919,N_21647);
xor U22457 (N_22457,N_21791,N_21608);
xor U22458 (N_22458,N_21514,N_21500);
xnor U22459 (N_22459,N_21694,N_21899);
xnor U22460 (N_22460,N_21637,N_21887);
or U22461 (N_22461,N_21902,N_21593);
nand U22462 (N_22462,N_21835,N_21962);
and U22463 (N_22463,N_21656,N_21914);
nor U22464 (N_22464,N_21933,N_21630);
or U22465 (N_22465,N_21805,N_21518);
xnor U22466 (N_22466,N_21621,N_21710);
and U22467 (N_22467,N_21620,N_21688);
nor U22468 (N_22468,N_21870,N_21732);
and U22469 (N_22469,N_21527,N_21572);
nor U22470 (N_22470,N_21844,N_21555);
xor U22471 (N_22471,N_21838,N_21749);
nor U22472 (N_22472,N_21569,N_21708);
and U22473 (N_22473,N_21666,N_21541);
and U22474 (N_22474,N_21793,N_21525);
and U22475 (N_22475,N_21640,N_21973);
and U22476 (N_22476,N_21751,N_21729);
or U22477 (N_22477,N_21897,N_21728);
xnor U22478 (N_22478,N_21857,N_21635);
and U22479 (N_22479,N_21659,N_21939);
and U22480 (N_22480,N_21839,N_21906);
nand U22481 (N_22481,N_21986,N_21620);
nor U22482 (N_22482,N_21554,N_21643);
xnor U22483 (N_22483,N_21809,N_21767);
or U22484 (N_22484,N_21514,N_21867);
xnor U22485 (N_22485,N_21840,N_21806);
xor U22486 (N_22486,N_21865,N_21684);
nand U22487 (N_22487,N_21914,N_21567);
or U22488 (N_22488,N_21513,N_21922);
and U22489 (N_22489,N_21729,N_21994);
nor U22490 (N_22490,N_21784,N_21713);
nor U22491 (N_22491,N_21718,N_21626);
nor U22492 (N_22492,N_21854,N_21850);
nor U22493 (N_22493,N_21797,N_21528);
nand U22494 (N_22494,N_21830,N_21866);
and U22495 (N_22495,N_21537,N_21799);
xor U22496 (N_22496,N_21961,N_21522);
and U22497 (N_22497,N_21686,N_21964);
and U22498 (N_22498,N_21718,N_21548);
and U22499 (N_22499,N_21915,N_21794);
xnor U22500 (N_22500,N_22379,N_22128);
and U22501 (N_22501,N_22484,N_22031);
nand U22502 (N_22502,N_22327,N_22049);
nand U22503 (N_22503,N_22374,N_22483);
nor U22504 (N_22504,N_22365,N_22094);
or U22505 (N_22505,N_22352,N_22410);
nor U22506 (N_22506,N_22239,N_22170);
xor U22507 (N_22507,N_22281,N_22441);
and U22508 (N_22508,N_22419,N_22383);
nand U22509 (N_22509,N_22032,N_22443);
or U22510 (N_22510,N_22320,N_22323);
or U22511 (N_22511,N_22378,N_22103);
nand U22512 (N_22512,N_22226,N_22356);
and U22513 (N_22513,N_22242,N_22291);
and U22514 (N_22514,N_22305,N_22053);
nand U22515 (N_22515,N_22423,N_22440);
xor U22516 (N_22516,N_22260,N_22150);
nand U22517 (N_22517,N_22045,N_22208);
nor U22518 (N_22518,N_22171,N_22288);
xor U22519 (N_22519,N_22360,N_22283);
nand U22520 (N_22520,N_22039,N_22401);
or U22521 (N_22521,N_22185,N_22349);
nand U22522 (N_22522,N_22167,N_22308);
nor U22523 (N_22523,N_22263,N_22471);
nor U22524 (N_22524,N_22033,N_22013);
or U22525 (N_22525,N_22102,N_22057);
nand U22526 (N_22526,N_22119,N_22001);
nor U22527 (N_22527,N_22165,N_22160);
nor U22528 (N_22528,N_22307,N_22386);
nor U22529 (N_22529,N_22331,N_22144);
xor U22530 (N_22530,N_22442,N_22458);
nor U22531 (N_22531,N_22496,N_22205);
xnor U22532 (N_22532,N_22136,N_22427);
xor U22533 (N_22533,N_22491,N_22285);
or U22534 (N_22534,N_22002,N_22355);
xnor U22535 (N_22535,N_22137,N_22181);
or U22536 (N_22536,N_22343,N_22490);
or U22537 (N_22537,N_22473,N_22451);
or U22538 (N_22538,N_22147,N_22105);
nor U22539 (N_22539,N_22123,N_22130);
nor U22540 (N_22540,N_22418,N_22061);
nand U22541 (N_22541,N_22209,N_22309);
nor U22542 (N_22542,N_22151,N_22254);
xnor U22543 (N_22543,N_22248,N_22408);
xor U22544 (N_22544,N_22036,N_22395);
and U22545 (N_22545,N_22329,N_22158);
nor U22546 (N_22546,N_22044,N_22078);
and U22547 (N_22547,N_22012,N_22085);
nand U22548 (N_22548,N_22186,N_22413);
or U22549 (N_22549,N_22474,N_22172);
xnor U22550 (N_22550,N_22030,N_22071);
or U22551 (N_22551,N_22026,N_22357);
nor U22552 (N_22552,N_22231,N_22269);
or U22553 (N_22553,N_22475,N_22354);
or U22554 (N_22554,N_22138,N_22194);
xnor U22555 (N_22555,N_22425,N_22249);
and U22556 (N_22556,N_22132,N_22081);
nor U22557 (N_22557,N_22051,N_22481);
and U22558 (N_22558,N_22371,N_22113);
nand U22559 (N_22559,N_22019,N_22008);
nand U22560 (N_22560,N_22361,N_22325);
and U22561 (N_22561,N_22224,N_22333);
nand U22562 (N_22562,N_22162,N_22237);
nand U22563 (N_22563,N_22096,N_22328);
nand U22564 (N_22564,N_22430,N_22313);
or U22565 (N_22565,N_22477,N_22214);
nor U22566 (N_22566,N_22256,N_22411);
and U22567 (N_22567,N_22335,N_22017);
nand U22568 (N_22568,N_22042,N_22211);
nor U22569 (N_22569,N_22275,N_22429);
nand U22570 (N_22570,N_22337,N_22197);
and U22571 (N_22571,N_22265,N_22290);
nor U22572 (N_22572,N_22083,N_22048);
nor U22573 (N_22573,N_22052,N_22054);
and U22574 (N_22574,N_22183,N_22225);
and U22575 (N_22575,N_22180,N_22292);
nand U22576 (N_22576,N_22375,N_22005);
xnor U22577 (N_22577,N_22279,N_22227);
nor U22578 (N_22578,N_22196,N_22041);
or U22579 (N_22579,N_22240,N_22212);
or U22580 (N_22580,N_22424,N_22121);
nand U22581 (N_22581,N_22255,N_22312);
and U22582 (N_22582,N_22278,N_22306);
nor U22583 (N_22583,N_22345,N_22038);
nor U22584 (N_22584,N_22104,N_22101);
and U22585 (N_22585,N_22079,N_22216);
or U22586 (N_22586,N_22110,N_22220);
nand U22587 (N_22587,N_22184,N_22022);
or U22588 (N_22588,N_22493,N_22339);
nand U22589 (N_22589,N_22326,N_22348);
nand U22590 (N_22590,N_22107,N_22011);
or U22591 (N_22591,N_22295,N_22176);
nor U22592 (N_22592,N_22407,N_22006);
and U22593 (N_22593,N_22402,N_22193);
and U22594 (N_22594,N_22015,N_22095);
nor U22595 (N_22595,N_22399,N_22433);
xor U22596 (N_22596,N_22029,N_22392);
nor U22597 (N_22597,N_22297,N_22228);
nand U22598 (N_22598,N_22321,N_22222);
and U22599 (N_22599,N_22479,N_22449);
nor U22600 (N_22600,N_22494,N_22060);
or U22601 (N_22601,N_22201,N_22416);
or U22602 (N_22602,N_22446,N_22245);
nand U22603 (N_22603,N_22089,N_22190);
nand U22604 (N_22604,N_22252,N_22324);
and U22605 (N_22605,N_22341,N_22210);
and U22606 (N_22606,N_22109,N_22420);
nor U22607 (N_22607,N_22223,N_22422);
or U22608 (N_22608,N_22065,N_22134);
nand U22609 (N_22609,N_22404,N_22097);
and U22610 (N_22610,N_22298,N_22043);
nor U22611 (N_22611,N_22315,N_22236);
nand U22612 (N_22612,N_22142,N_22317);
or U22613 (N_22613,N_22489,N_22164);
xor U22614 (N_22614,N_22463,N_22334);
and U22615 (N_22615,N_22319,N_22131);
nor U22616 (N_22616,N_22247,N_22367);
xor U22617 (N_22617,N_22100,N_22445);
xor U22618 (N_22618,N_22074,N_22232);
nor U22619 (N_22619,N_22314,N_22466);
nand U22620 (N_22620,N_22221,N_22090);
xor U22621 (N_22621,N_22372,N_22086);
or U22622 (N_22622,N_22262,N_22387);
nand U22623 (N_22623,N_22124,N_22431);
and U22624 (N_22624,N_22120,N_22056);
and U22625 (N_22625,N_22310,N_22390);
nand U22626 (N_22626,N_22362,N_22447);
or U22627 (N_22627,N_22116,N_22351);
or U22628 (N_22628,N_22454,N_22082);
nand U22629 (N_22629,N_22296,N_22139);
and U22630 (N_22630,N_22462,N_22087);
or U22631 (N_22631,N_22125,N_22182);
nor U22632 (N_22632,N_22280,N_22485);
xnor U22633 (N_22633,N_22117,N_22385);
and U22634 (N_22634,N_22173,N_22482);
xor U22635 (N_22635,N_22108,N_22099);
nor U22636 (N_22636,N_22301,N_22289);
nor U22637 (N_22637,N_22270,N_22072);
xor U22638 (N_22638,N_22020,N_22047);
or U22639 (N_22639,N_22338,N_22114);
nor U22640 (N_22640,N_22010,N_22456);
or U22641 (N_22641,N_22293,N_22003);
xnor U22642 (N_22642,N_22267,N_22322);
nand U22643 (N_22643,N_22219,N_22203);
or U22644 (N_22644,N_22344,N_22303);
or U22645 (N_22645,N_22217,N_22187);
or U22646 (N_22646,N_22480,N_22486);
and U22647 (N_22647,N_22432,N_22068);
nor U22648 (N_22648,N_22453,N_22340);
or U22649 (N_22649,N_22073,N_22257);
or U22650 (N_22650,N_22455,N_22396);
xnor U22651 (N_22651,N_22406,N_22055);
and U22652 (N_22652,N_22014,N_22177);
nand U22653 (N_22653,N_22369,N_22204);
xor U22654 (N_22654,N_22188,N_22088);
nand U22655 (N_22655,N_22435,N_22023);
and U22656 (N_22656,N_22215,N_22464);
nand U22657 (N_22657,N_22330,N_22364);
nor U22658 (N_22658,N_22145,N_22436);
and U22659 (N_22659,N_22034,N_22381);
nor U22660 (N_22660,N_22403,N_22168);
or U22661 (N_22661,N_22389,N_22342);
xnor U22662 (N_22662,N_22066,N_22311);
or U22663 (N_22663,N_22428,N_22046);
or U22664 (N_22664,N_22159,N_22253);
nor U22665 (N_22665,N_22206,N_22476);
nor U22666 (N_22666,N_22370,N_22492);
nor U22667 (N_22667,N_22273,N_22450);
or U22668 (N_22668,N_22300,N_22016);
xnor U22669 (N_22669,N_22282,N_22274);
or U22670 (N_22670,N_22202,N_22487);
nand U22671 (N_22671,N_22111,N_22318);
nor U22672 (N_22672,N_22037,N_22118);
nor U22673 (N_22673,N_22135,N_22200);
or U22674 (N_22674,N_22398,N_22112);
nor U22675 (N_22675,N_22470,N_22434);
nor U22676 (N_22676,N_22384,N_22098);
nor U22677 (N_22677,N_22021,N_22175);
nor U22678 (N_22678,N_22478,N_22394);
nor U22679 (N_22679,N_22437,N_22163);
or U22680 (N_22680,N_22472,N_22353);
xor U22681 (N_22681,N_22400,N_22141);
and U22682 (N_22682,N_22009,N_22152);
or U22683 (N_22683,N_22234,N_22235);
or U22684 (N_22684,N_22063,N_22122);
xnor U22685 (N_22685,N_22488,N_22213);
nand U22686 (N_22686,N_22148,N_22092);
nand U22687 (N_22687,N_22391,N_22178);
xor U22688 (N_22688,N_22380,N_22294);
nor U22689 (N_22689,N_22363,N_22018);
or U22690 (N_22690,N_22166,N_22457);
xor U22691 (N_22691,N_22241,N_22229);
nor U22692 (N_22692,N_22316,N_22149);
nand U22693 (N_22693,N_22459,N_22258);
xor U22694 (N_22694,N_22373,N_22077);
and U22695 (N_22695,N_22075,N_22304);
xor U22696 (N_22696,N_22040,N_22233);
or U22697 (N_22697,N_22497,N_22004);
nand U22698 (N_22698,N_22465,N_22069);
nor U22699 (N_22699,N_22126,N_22452);
or U22700 (N_22700,N_22080,N_22024);
xor U22701 (N_22701,N_22007,N_22093);
xor U22702 (N_22702,N_22251,N_22115);
nor U22703 (N_22703,N_22062,N_22243);
and U22704 (N_22704,N_22091,N_22161);
nand U22705 (N_22705,N_22332,N_22460);
nor U22706 (N_22706,N_22358,N_22264);
or U22707 (N_22707,N_22439,N_22246);
and U22708 (N_22708,N_22405,N_22347);
and U22709 (N_22709,N_22271,N_22143);
or U22710 (N_22710,N_22058,N_22146);
nor U22711 (N_22711,N_22426,N_22415);
xnor U22712 (N_22712,N_22027,N_22189);
nor U22713 (N_22713,N_22421,N_22025);
xor U22714 (N_22714,N_22250,N_22414);
nor U22715 (N_22715,N_22127,N_22174);
xor U22716 (N_22716,N_22268,N_22388);
nor U22717 (N_22717,N_22498,N_22140);
nor U22718 (N_22718,N_22359,N_22153);
nor U22719 (N_22719,N_22000,N_22438);
nand U22720 (N_22720,N_22035,N_22238);
nand U22721 (N_22721,N_22299,N_22409);
nor U22722 (N_22722,N_22050,N_22286);
xor U22723 (N_22723,N_22284,N_22192);
or U22724 (N_22724,N_22397,N_22495);
xnor U22725 (N_22725,N_22261,N_22366);
nor U22726 (N_22726,N_22302,N_22412);
or U22727 (N_22727,N_22154,N_22417);
xnor U22728 (N_22728,N_22266,N_22377);
nor U22729 (N_22729,N_22157,N_22198);
nand U22730 (N_22730,N_22067,N_22230);
nand U22731 (N_22731,N_22277,N_22133);
xor U22732 (N_22732,N_22444,N_22084);
nor U22733 (N_22733,N_22028,N_22156);
xor U22734 (N_22734,N_22179,N_22287);
and U22735 (N_22735,N_22272,N_22199);
nand U22736 (N_22736,N_22376,N_22059);
and U22737 (N_22737,N_22468,N_22169);
xnor U22738 (N_22738,N_22350,N_22191);
nor U22739 (N_22739,N_22336,N_22499);
nor U22740 (N_22740,N_22195,N_22218);
nor U22741 (N_22741,N_22448,N_22106);
or U22742 (N_22742,N_22070,N_22346);
or U22743 (N_22743,N_22129,N_22244);
and U22744 (N_22744,N_22469,N_22368);
xor U22745 (N_22745,N_22207,N_22155);
and U22746 (N_22746,N_22259,N_22467);
nor U22747 (N_22747,N_22076,N_22393);
nor U22748 (N_22748,N_22276,N_22461);
or U22749 (N_22749,N_22382,N_22064);
xnor U22750 (N_22750,N_22348,N_22110);
xnor U22751 (N_22751,N_22212,N_22425);
and U22752 (N_22752,N_22200,N_22406);
nand U22753 (N_22753,N_22498,N_22334);
or U22754 (N_22754,N_22295,N_22306);
nor U22755 (N_22755,N_22449,N_22155);
nand U22756 (N_22756,N_22277,N_22058);
nand U22757 (N_22757,N_22206,N_22248);
or U22758 (N_22758,N_22368,N_22221);
and U22759 (N_22759,N_22213,N_22134);
and U22760 (N_22760,N_22000,N_22235);
nor U22761 (N_22761,N_22301,N_22287);
nor U22762 (N_22762,N_22075,N_22384);
nor U22763 (N_22763,N_22321,N_22208);
xor U22764 (N_22764,N_22410,N_22097);
nor U22765 (N_22765,N_22341,N_22153);
nor U22766 (N_22766,N_22419,N_22373);
nor U22767 (N_22767,N_22050,N_22101);
and U22768 (N_22768,N_22246,N_22220);
nor U22769 (N_22769,N_22204,N_22366);
nor U22770 (N_22770,N_22321,N_22141);
or U22771 (N_22771,N_22037,N_22350);
nand U22772 (N_22772,N_22311,N_22420);
xor U22773 (N_22773,N_22223,N_22236);
xnor U22774 (N_22774,N_22146,N_22111);
nand U22775 (N_22775,N_22373,N_22291);
and U22776 (N_22776,N_22279,N_22169);
and U22777 (N_22777,N_22128,N_22295);
or U22778 (N_22778,N_22044,N_22218);
or U22779 (N_22779,N_22365,N_22078);
nor U22780 (N_22780,N_22449,N_22153);
and U22781 (N_22781,N_22083,N_22463);
xor U22782 (N_22782,N_22164,N_22276);
nor U22783 (N_22783,N_22320,N_22078);
nand U22784 (N_22784,N_22342,N_22283);
nor U22785 (N_22785,N_22254,N_22330);
or U22786 (N_22786,N_22496,N_22004);
nand U22787 (N_22787,N_22434,N_22037);
and U22788 (N_22788,N_22111,N_22211);
nand U22789 (N_22789,N_22045,N_22246);
or U22790 (N_22790,N_22087,N_22281);
or U22791 (N_22791,N_22390,N_22263);
xor U22792 (N_22792,N_22239,N_22425);
or U22793 (N_22793,N_22184,N_22360);
xor U22794 (N_22794,N_22355,N_22197);
xnor U22795 (N_22795,N_22026,N_22231);
and U22796 (N_22796,N_22342,N_22458);
or U22797 (N_22797,N_22013,N_22309);
and U22798 (N_22798,N_22358,N_22476);
and U22799 (N_22799,N_22419,N_22347);
nand U22800 (N_22800,N_22174,N_22120);
nor U22801 (N_22801,N_22012,N_22490);
xnor U22802 (N_22802,N_22279,N_22186);
nand U22803 (N_22803,N_22079,N_22066);
nor U22804 (N_22804,N_22443,N_22366);
xnor U22805 (N_22805,N_22059,N_22013);
xor U22806 (N_22806,N_22093,N_22495);
nand U22807 (N_22807,N_22465,N_22419);
xnor U22808 (N_22808,N_22203,N_22407);
xor U22809 (N_22809,N_22455,N_22035);
xnor U22810 (N_22810,N_22366,N_22491);
nand U22811 (N_22811,N_22072,N_22018);
nand U22812 (N_22812,N_22390,N_22132);
nor U22813 (N_22813,N_22077,N_22294);
and U22814 (N_22814,N_22383,N_22373);
or U22815 (N_22815,N_22290,N_22168);
and U22816 (N_22816,N_22095,N_22068);
nand U22817 (N_22817,N_22225,N_22210);
nor U22818 (N_22818,N_22343,N_22015);
nor U22819 (N_22819,N_22162,N_22015);
and U22820 (N_22820,N_22476,N_22007);
nand U22821 (N_22821,N_22192,N_22077);
nor U22822 (N_22822,N_22124,N_22277);
nand U22823 (N_22823,N_22419,N_22319);
nor U22824 (N_22824,N_22092,N_22399);
xor U22825 (N_22825,N_22272,N_22248);
nor U22826 (N_22826,N_22064,N_22094);
and U22827 (N_22827,N_22093,N_22004);
or U22828 (N_22828,N_22191,N_22063);
nor U22829 (N_22829,N_22087,N_22469);
nand U22830 (N_22830,N_22223,N_22198);
nand U22831 (N_22831,N_22395,N_22391);
and U22832 (N_22832,N_22219,N_22474);
nand U22833 (N_22833,N_22473,N_22178);
and U22834 (N_22834,N_22382,N_22019);
xor U22835 (N_22835,N_22348,N_22154);
nor U22836 (N_22836,N_22065,N_22059);
nor U22837 (N_22837,N_22121,N_22490);
xor U22838 (N_22838,N_22327,N_22326);
nand U22839 (N_22839,N_22396,N_22026);
nand U22840 (N_22840,N_22070,N_22341);
xor U22841 (N_22841,N_22018,N_22055);
and U22842 (N_22842,N_22359,N_22177);
nand U22843 (N_22843,N_22204,N_22239);
xor U22844 (N_22844,N_22489,N_22121);
nand U22845 (N_22845,N_22249,N_22196);
nand U22846 (N_22846,N_22437,N_22465);
nor U22847 (N_22847,N_22025,N_22400);
nand U22848 (N_22848,N_22024,N_22042);
xnor U22849 (N_22849,N_22246,N_22388);
xnor U22850 (N_22850,N_22099,N_22464);
nor U22851 (N_22851,N_22012,N_22024);
or U22852 (N_22852,N_22041,N_22370);
or U22853 (N_22853,N_22022,N_22056);
or U22854 (N_22854,N_22451,N_22394);
nor U22855 (N_22855,N_22487,N_22329);
nor U22856 (N_22856,N_22360,N_22217);
nor U22857 (N_22857,N_22115,N_22245);
nor U22858 (N_22858,N_22422,N_22324);
nand U22859 (N_22859,N_22102,N_22252);
or U22860 (N_22860,N_22233,N_22000);
or U22861 (N_22861,N_22068,N_22303);
xor U22862 (N_22862,N_22019,N_22403);
xor U22863 (N_22863,N_22060,N_22455);
or U22864 (N_22864,N_22461,N_22290);
xor U22865 (N_22865,N_22339,N_22001);
and U22866 (N_22866,N_22157,N_22484);
xor U22867 (N_22867,N_22298,N_22127);
xor U22868 (N_22868,N_22289,N_22292);
nor U22869 (N_22869,N_22171,N_22035);
nor U22870 (N_22870,N_22129,N_22319);
or U22871 (N_22871,N_22236,N_22482);
xnor U22872 (N_22872,N_22189,N_22381);
nor U22873 (N_22873,N_22025,N_22104);
nand U22874 (N_22874,N_22001,N_22335);
or U22875 (N_22875,N_22135,N_22113);
or U22876 (N_22876,N_22344,N_22234);
xor U22877 (N_22877,N_22340,N_22346);
or U22878 (N_22878,N_22424,N_22082);
or U22879 (N_22879,N_22249,N_22481);
or U22880 (N_22880,N_22355,N_22026);
nor U22881 (N_22881,N_22207,N_22355);
or U22882 (N_22882,N_22075,N_22487);
nand U22883 (N_22883,N_22108,N_22048);
nor U22884 (N_22884,N_22009,N_22428);
nand U22885 (N_22885,N_22111,N_22407);
or U22886 (N_22886,N_22101,N_22468);
and U22887 (N_22887,N_22127,N_22231);
nor U22888 (N_22888,N_22031,N_22069);
nor U22889 (N_22889,N_22277,N_22375);
and U22890 (N_22890,N_22294,N_22176);
xnor U22891 (N_22891,N_22023,N_22053);
nand U22892 (N_22892,N_22010,N_22482);
xnor U22893 (N_22893,N_22335,N_22124);
xnor U22894 (N_22894,N_22055,N_22100);
or U22895 (N_22895,N_22196,N_22348);
or U22896 (N_22896,N_22369,N_22424);
xor U22897 (N_22897,N_22355,N_22333);
xor U22898 (N_22898,N_22136,N_22248);
and U22899 (N_22899,N_22199,N_22045);
nand U22900 (N_22900,N_22058,N_22334);
nor U22901 (N_22901,N_22177,N_22158);
and U22902 (N_22902,N_22097,N_22153);
nand U22903 (N_22903,N_22173,N_22273);
and U22904 (N_22904,N_22490,N_22241);
nor U22905 (N_22905,N_22256,N_22179);
or U22906 (N_22906,N_22268,N_22066);
xor U22907 (N_22907,N_22408,N_22460);
xor U22908 (N_22908,N_22256,N_22301);
or U22909 (N_22909,N_22060,N_22390);
xor U22910 (N_22910,N_22178,N_22181);
or U22911 (N_22911,N_22203,N_22237);
nand U22912 (N_22912,N_22298,N_22355);
or U22913 (N_22913,N_22081,N_22298);
and U22914 (N_22914,N_22056,N_22256);
nand U22915 (N_22915,N_22061,N_22113);
and U22916 (N_22916,N_22205,N_22309);
xor U22917 (N_22917,N_22072,N_22441);
nor U22918 (N_22918,N_22298,N_22350);
xor U22919 (N_22919,N_22447,N_22204);
xor U22920 (N_22920,N_22111,N_22252);
or U22921 (N_22921,N_22100,N_22385);
nand U22922 (N_22922,N_22363,N_22414);
and U22923 (N_22923,N_22318,N_22254);
xor U22924 (N_22924,N_22024,N_22283);
xnor U22925 (N_22925,N_22121,N_22236);
and U22926 (N_22926,N_22329,N_22461);
nand U22927 (N_22927,N_22436,N_22462);
or U22928 (N_22928,N_22296,N_22197);
nand U22929 (N_22929,N_22069,N_22271);
and U22930 (N_22930,N_22052,N_22247);
nand U22931 (N_22931,N_22092,N_22433);
xnor U22932 (N_22932,N_22471,N_22139);
and U22933 (N_22933,N_22040,N_22161);
nor U22934 (N_22934,N_22191,N_22044);
nand U22935 (N_22935,N_22286,N_22301);
and U22936 (N_22936,N_22267,N_22427);
or U22937 (N_22937,N_22394,N_22460);
nor U22938 (N_22938,N_22459,N_22362);
nor U22939 (N_22939,N_22434,N_22241);
xor U22940 (N_22940,N_22237,N_22097);
or U22941 (N_22941,N_22428,N_22467);
or U22942 (N_22942,N_22011,N_22134);
and U22943 (N_22943,N_22194,N_22171);
nand U22944 (N_22944,N_22058,N_22218);
nor U22945 (N_22945,N_22079,N_22137);
nor U22946 (N_22946,N_22445,N_22294);
nand U22947 (N_22947,N_22070,N_22061);
nand U22948 (N_22948,N_22182,N_22419);
and U22949 (N_22949,N_22361,N_22483);
xnor U22950 (N_22950,N_22291,N_22015);
or U22951 (N_22951,N_22177,N_22220);
nand U22952 (N_22952,N_22343,N_22417);
and U22953 (N_22953,N_22414,N_22434);
and U22954 (N_22954,N_22455,N_22158);
or U22955 (N_22955,N_22440,N_22056);
nor U22956 (N_22956,N_22164,N_22270);
nor U22957 (N_22957,N_22347,N_22221);
nand U22958 (N_22958,N_22137,N_22499);
or U22959 (N_22959,N_22065,N_22472);
nand U22960 (N_22960,N_22114,N_22474);
nor U22961 (N_22961,N_22108,N_22207);
nor U22962 (N_22962,N_22473,N_22427);
and U22963 (N_22963,N_22375,N_22148);
or U22964 (N_22964,N_22046,N_22058);
and U22965 (N_22965,N_22260,N_22269);
xor U22966 (N_22966,N_22141,N_22153);
and U22967 (N_22967,N_22252,N_22047);
or U22968 (N_22968,N_22423,N_22160);
or U22969 (N_22969,N_22401,N_22465);
and U22970 (N_22970,N_22239,N_22002);
nand U22971 (N_22971,N_22387,N_22452);
nor U22972 (N_22972,N_22257,N_22328);
and U22973 (N_22973,N_22297,N_22390);
or U22974 (N_22974,N_22453,N_22094);
or U22975 (N_22975,N_22418,N_22298);
nand U22976 (N_22976,N_22277,N_22331);
or U22977 (N_22977,N_22434,N_22139);
nor U22978 (N_22978,N_22153,N_22240);
xor U22979 (N_22979,N_22417,N_22241);
or U22980 (N_22980,N_22413,N_22341);
and U22981 (N_22981,N_22220,N_22012);
and U22982 (N_22982,N_22348,N_22100);
nand U22983 (N_22983,N_22277,N_22328);
nand U22984 (N_22984,N_22484,N_22144);
nor U22985 (N_22985,N_22404,N_22256);
nor U22986 (N_22986,N_22353,N_22277);
nor U22987 (N_22987,N_22321,N_22364);
and U22988 (N_22988,N_22493,N_22264);
nand U22989 (N_22989,N_22474,N_22373);
and U22990 (N_22990,N_22171,N_22446);
and U22991 (N_22991,N_22367,N_22178);
nor U22992 (N_22992,N_22461,N_22322);
or U22993 (N_22993,N_22296,N_22391);
and U22994 (N_22994,N_22489,N_22344);
xnor U22995 (N_22995,N_22382,N_22198);
and U22996 (N_22996,N_22021,N_22317);
xor U22997 (N_22997,N_22430,N_22097);
or U22998 (N_22998,N_22475,N_22119);
xnor U22999 (N_22999,N_22203,N_22310);
xor U23000 (N_23000,N_22760,N_22977);
nor U23001 (N_23001,N_22592,N_22913);
or U23002 (N_23002,N_22656,N_22584);
nand U23003 (N_23003,N_22882,N_22520);
nand U23004 (N_23004,N_22859,N_22537);
or U23005 (N_23005,N_22790,N_22660);
or U23006 (N_23006,N_22665,N_22690);
and U23007 (N_23007,N_22762,N_22826);
and U23008 (N_23008,N_22595,N_22582);
or U23009 (N_23009,N_22551,N_22532);
nand U23010 (N_23010,N_22625,N_22563);
nand U23011 (N_23011,N_22650,N_22905);
or U23012 (N_23012,N_22804,N_22755);
and U23013 (N_23013,N_22587,N_22978);
or U23014 (N_23014,N_22854,N_22529);
xnor U23015 (N_23015,N_22813,N_22961);
nor U23016 (N_23016,N_22597,N_22632);
and U23017 (N_23017,N_22679,N_22929);
nand U23018 (N_23018,N_22623,N_22748);
nor U23019 (N_23019,N_22766,N_22526);
nor U23020 (N_23020,N_22709,N_22674);
or U23021 (N_23021,N_22543,N_22620);
or U23022 (N_23022,N_22522,N_22899);
nand U23023 (N_23023,N_22993,N_22586);
nor U23024 (N_23024,N_22682,N_22821);
and U23025 (N_23025,N_22874,N_22606);
and U23026 (N_23026,N_22744,N_22856);
xor U23027 (N_23027,N_22910,N_22718);
nand U23028 (N_23028,N_22548,N_22628);
or U23029 (N_23029,N_22895,N_22521);
and U23030 (N_23030,N_22873,N_22825);
or U23031 (N_23031,N_22667,N_22735);
and U23032 (N_23032,N_22773,N_22917);
nor U23033 (N_23033,N_22890,N_22759);
nor U23034 (N_23034,N_22765,N_22539);
nor U23035 (N_23035,N_22603,N_22731);
xnor U23036 (N_23036,N_22888,N_22875);
or U23037 (N_23037,N_22538,N_22997);
and U23038 (N_23038,N_22750,N_22732);
and U23039 (N_23039,N_22953,N_22823);
xor U23040 (N_23040,N_22542,N_22545);
and U23041 (N_23041,N_22962,N_22878);
xnor U23042 (N_23042,N_22747,N_22619);
xnor U23043 (N_23043,N_22872,N_22559);
nor U23044 (N_23044,N_22915,N_22906);
nand U23045 (N_23045,N_22975,N_22992);
and U23046 (N_23046,N_22863,N_22883);
xor U23047 (N_23047,N_22843,N_22796);
or U23048 (N_23048,N_22830,N_22786);
nor U23049 (N_23049,N_22585,N_22635);
xnor U23050 (N_23050,N_22810,N_22927);
nand U23051 (N_23051,N_22970,N_22662);
nor U23052 (N_23052,N_22552,N_22835);
nor U23053 (N_23053,N_22651,N_22904);
nand U23054 (N_23054,N_22562,N_22787);
nand U23055 (N_23055,N_22955,N_22911);
and U23056 (N_23056,N_22699,N_22653);
xnor U23057 (N_23057,N_22643,N_22509);
nor U23058 (N_23058,N_22837,N_22842);
nand U23059 (N_23059,N_22897,N_22633);
nand U23060 (N_23060,N_22921,N_22641);
nand U23061 (N_23061,N_22969,N_22518);
or U23062 (N_23062,N_22935,N_22968);
nor U23063 (N_23063,N_22776,N_22946);
nor U23064 (N_23064,N_22885,N_22546);
or U23065 (N_23065,N_22881,N_22999);
nand U23066 (N_23066,N_22805,N_22980);
xor U23067 (N_23067,N_22752,N_22788);
or U23068 (N_23068,N_22892,N_22986);
xor U23069 (N_23069,N_22549,N_22743);
and U23070 (N_23070,N_22500,N_22964);
xnor U23071 (N_23071,N_22951,N_22852);
xor U23072 (N_23072,N_22928,N_22506);
and U23073 (N_23073,N_22612,N_22954);
nor U23074 (N_23074,N_22700,N_22754);
or U23075 (N_23075,N_22753,N_22907);
nand U23076 (N_23076,N_22801,N_22864);
and U23077 (N_23077,N_22893,N_22689);
or U23078 (N_23078,N_22916,N_22507);
xnor U23079 (N_23079,N_22624,N_22841);
or U23080 (N_23080,N_22886,N_22716);
and U23081 (N_23081,N_22581,N_22794);
and U23082 (N_23082,N_22741,N_22902);
nand U23083 (N_23083,N_22965,N_22615);
or U23084 (N_23084,N_22503,N_22909);
or U23085 (N_23085,N_22621,N_22678);
xor U23086 (N_23086,N_22736,N_22827);
nand U23087 (N_23087,N_22574,N_22703);
or U23088 (N_23088,N_22914,N_22833);
nand U23089 (N_23089,N_22922,N_22933);
nand U23090 (N_23090,N_22555,N_22779);
xor U23091 (N_23091,N_22894,N_22880);
or U23092 (N_23092,N_22834,N_22816);
nand U23093 (N_23093,N_22636,N_22756);
or U23094 (N_23094,N_22535,N_22676);
nor U23095 (N_23095,N_22565,N_22793);
or U23096 (N_23096,N_22634,N_22695);
or U23097 (N_23097,N_22711,N_22717);
and U23098 (N_23098,N_22956,N_22784);
or U23099 (N_23099,N_22647,N_22848);
nor U23100 (N_23100,N_22761,N_22818);
and U23101 (N_23101,N_22569,N_22661);
nand U23102 (N_23102,N_22558,N_22819);
nor U23103 (N_23103,N_22663,N_22560);
xor U23104 (N_23104,N_22683,N_22723);
xnor U23105 (N_23105,N_22722,N_22797);
or U23106 (N_23106,N_22697,N_22926);
nand U23107 (N_23107,N_22573,N_22828);
nand U23108 (N_23108,N_22846,N_22767);
or U23109 (N_23109,N_22831,N_22778);
and U23110 (N_23110,N_22959,N_22727);
xnor U23111 (N_23111,N_22795,N_22578);
xor U23112 (N_23112,N_22877,N_22508);
and U23113 (N_23113,N_22769,N_22939);
or U23114 (N_23114,N_22958,N_22630);
or U23115 (N_23115,N_22824,N_22685);
nand U23116 (N_23116,N_22714,N_22626);
and U23117 (N_23117,N_22698,N_22629);
nand U23118 (N_23118,N_22639,N_22853);
nor U23119 (N_23119,N_22668,N_22822);
nor U23120 (N_23120,N_22594,N_22862);
and U23121 (N_23121,N_22931,N_22974);
nor U23122 (N_23122,N_22687,N_22601);
xnor U23123 (N_23123,N_22912,N_22791);
and U23124 (N_23124,N_22807,N_22572);
or U23125 (N_23125,N_22947,N_22949);
or U23126 (N_23126,N_22940,N_22729);
and U23127 (N_23127,N_22876,N_22941);
nand U23128 (N_23128,N_22829,N_22996);
and U23129 (N_23129,N_22780,N_22924);
nand U23130 (N_23130,N_22884,N_22995);
and U23131 (N_23131,N_22934,N_22513);
nor U23132 (N_23132,N_22589,N_22879);
xor U23133 (N_23133,N_22920,N_22950);
nand U23134 (N_23134,N_22814,N_22596);
or U23135 (N_23135,N_22600,N_22708);
nand U23136 (N_23136,N_22945,N_22739);
nor U23137 (N_23137,N_22903,N_22638);
xor U23138 (N_23138,N_22775,N_22806);
nand U23139 (N_23139,N_22836,N_22654);
nand U23140 (N_23140,N_22745,N_22608);
nor U23141 (N_23141,N_22868,N_22771);
and U23142 (N_23142,N_22900,N_22936);
or U23143 (N_23143,N_22751,N_22789);
nand U23144 (N_23144,N_22571,N_22887);
or U23145 (N_23145,N_22607,N_22870);
nor U23146 (N_23146,N_22901,N_22557);
xnor U23147 (N_23147,N_22865,N_22764);
and U23148 (N_23148,N_22749,N_22757);
and U23149 (N_23149,N_22618,N_22737);
xnor U23150 (N_23150,N_22855,N_22800);
nor U23151 (N_23151,N_22983,N_22967);
nand U23152 (N_23152,N_22817,N_22923);
and U23153 (N_23153,N_22740,N_22631);
xnor U23154 (N_23154,N_22966,N_22721);
nand U23155 (N_23155,N_22525,N_22547);
nor U23156 (N_23156,N_22659,N_22501);
nand U23157 (N_23157,N_22658,N_22847);
nor U23158 (N_23158,N_22990,N_22567);
nor U23159 (N_23159,N_22815,N_22719);
xnor U23160 (N_23160,N_22693,N_22580);
and U23161 (N_23161,N_22564,N_22527);
and U23162 (N_23162,N_22541,N_22785);
nor U23163 (N_23163,N_22918,N_22973);
nand U23164 (N_23164,N_22994,N_22963);
or U23165 (N_23165,N_22561,N_22861);
nor U23166 (N_23166,N_22534,N_22728);
or U23167 (N_23167,N_22556,N_22982);
nor U23168 (N_23168,N_22531,N_22648);
and U23169 (N_23169,N_22715,N_22649);
or U23170 (N_23170,N_22688,N_22701);
xnor U23171 (N_23171,N_22669,N_22512);
or U23172 (N_23172,N_22839,N_22932);
nand U23173 (N_23173,N_22925,N_22707);
nand U23174 (N_23174,N_22979,N_22942);
xnor U23175 (N_23175,N_22763,N_22891);
and U23176 (N_23176,N_22738,N_22981);
or U23177 (N_23177,N_22998,N_22976);
or U23178 (N_23178,N_22577,N_22536);
and U23179 (N_23179,N_22889,N_22799);
nor U23180 (N_23180,N_22664,N_22777);
xor U23181 (N_23181,N_22684,N_22583);
nor U23182 (N_23182,N_22504,N_22742);
nor U23183 (N_23183,N_22972,N_22782);
and U23184 (N_23184,N_22971,N_22733);
nor U23185 (N_23185,N_22808,N_22524);
nand U23186 (N_23186,N_22591,N_22726);
nor U23187 (N_23187,N_22613,N_22919);
or U23188 (N_23188,N_22655,N_22730);
xor U23189 (N_23189,N_22640,N_22576);
and U23190 (N_23190,N_22937,N_22944);
and U23191 (N_23191,N_22991,N_22724);
nand U23192 (N_23192,N_22602,N_22812);
xnor U23193 (N_23193,N_22908,N_22988);
xnor U23194 (N_23194,N_22850,N_22938);
and U23195 (N_23195,N_22867,N_22948);
nor U23196 (N_23196,N_22666,N_22609);
nand U23197 (N_23197,N_22645,N_22519);
and U23198 (N_23198,N_22599,N_22798);
xnor U23199 (N_23199,N_22671,N_22866);
or U23200 (N_23200,N_22898,N_22691);
nand U23201 (N_23201,N_22517,N_22984);
xor U23202 (N_23202,N_22616,N_22811);
nor U23203 (N_23203,N_22725,N_22851);
xor U23204 (N_23204,N_22734,N_22670);
and U23205 (N_23205,N_22987,N_22675);
nor U23206 (N_23206,N_22832,N_22985);
or U23207 (N_23207,N_22590,N_22652);
nor U23208 (N_23208,N_22502,N_22960);
or U23209 (N_23209,N_22845,N_22696);
nand U23210 (N_23210,N_22792,N_22511);
xnor U23211 (N_23211,N_22702,N_22774);
and U23212 (N_23212,N_22781,N_22644);
nand U23213 (N_23213,N_22713,N_22720);
nand U23214 (N_23214,N_22627,N_22515);
and U23215 (N_23215,N_22869,N_22530);
or U23216 (N_23216,N_22989,N_22554);
nor U23217 (N_23217,N_22871,N_22553);
and U23218 (N_23218,N_22943,N_22622);
nand U23219 (N_23219,N_22579,N_22692);
nand U23220 (N_23220,N_22746,N_22657);
nand U23221 (N_23221,N_22505,N_22604);
and U23222 (N_23222,N_22610,N_22772);
nor U23223 (N_23223,N_22849,N_22857);
xnor U23224 (N_23224,N_22930,N_22704);
and U23225 (N_23225,N_22611,N_22598);
xor U23226 (N_23226,N_22566,N_22694);
xor U23227 (N_23227,N_22710,N_22770);
and U23228 (N_23228,N_22860,N_22705);
or U23229 (N_23229,N_22605,N_22896);
and U23230 (N_23230,N_22768,N_22809);
and U23231 (N_23231,N_22840,N_22544);
nor U23232 (N_23232,N_22952,N_22614);
nand U23233 (N_23233,N_22588,N_22712);
xor U23234 (N_23234,N_22540,N_22838);
and U23235 (N_23235,N_22844,N_22677);
xnor U23236 (N_23236,N_22637,N_22516);
nand U23237 (N_23237,N_22523,N_22706);
and U23238 (N_23238,N_22957,N_22686);
nand U23239 (N_23239,N_22642,N_22802);
nor U23240 (N_23240,N_22858,N_22570);
nor U23241 (N_23241,N_22575,N_22568);
and U23242 (N_23242,N_22528,N_22593);
nor U23243 (N_23243,N_22550,N_22803);
xor U23244 (N_23244,N_22680,N_22681);
nand U23245 (N_23245,N_22820,N_22533);
xnor U23246 (N_23246,N_22758,N_22510);
nand U23247 (N_23247,N_22673,N_22672);
nand U23248 (N_23248,N_22514,N_22783);
nand U23249 (N_23249,N_22617,N_22646);
or U23250 (N_23250,N_22782,N_22519);
nor U23251 (N_23251,N_22595,N_22853);
nand U23252 (N_23252,N_22574,N_22861);
and U23253 (N_23253,N_22847,N_22802);
and U23254 (N_23254,N_22701,N_22858);
nor U23255 (N_23255,N_22529,N_22968);
xnor U23256 (N_23256,N_22560,N_22941);
xor U23257 (N_23257,N_22779,N_22758);
or U23258 (N_23258,N_22915,N_22579);
xnor U23259 (N_23259,N_22726,N_22974);
and U23260 (N_23260,N_22749,N_22955);
nand U23261 (N_23261,N_22910,N_22780);
nor U23262 (N_23262,N_22631,N_22993);
xnor U23263 (N_23263,N_22837,N_22975);
nand U23264 (N_23264,N_22626,N_22957);
or U23265 (N_23265,N_22965,N_22628);
or U23266 (N_23266,N_22944,N_22875);
nand U23267 (N_23267,N_22951,N_22602);
xnor U23268 (N_23268,N_22885,N_22841);
xor U23269 (N_23269,N_22638,N_22605);
nor U23270 (N_23270,N_22697,N_22701);
or U23271 (N_23271,N_22533,N_22553);
and U23272 (N_23272,N_22922,N_22525);
xor U23273 (N_23273,N_22820,N_22601);
or U23274 (N_23274,N_22687,N_22932);
and U23275 (N_23275,N_22788,N_22746);
nand U23276 (N_23276,N_22935,N_22545);
nand U23277 (N_23277,N_22604,N_22575);
xnor U23278 (N_23278,N_22941,N_22804);
nor U23279 (N_23279,N_22662,N_22609);
nand U23280 (N_23280,N_22699,N_22743);
nor U23281 (N_23281,N_22731,N_22559);
or U23282 (N_23282,N_22971,N_22617);
or U23283 (N_23283,N_22518,N_22907);
xor U23284 (N_23284,N_22868,N_22731);
or U23285 (N_23285,N_22967,N_22593);
xnor U23286 (N_23286,N_22547,N_22689);
nand U23287 (N_23287,N_22782,N_22533);
nand U23288 (N_23288,N_22677,N_22627);
xnor U23289 (N_23289,N_22591,N_22796);
and U23290 (N_23290,N_22823,N_22579);
and U23291 (N_23291,N_22515,N_22900);
nor U23292 (N_23292,N_22797,N_22542);
and U23293 (N_23293,N_22560,N_22674);
xnor U23294 (N_23294,N_22623,N_22939);
xor U23295 (N_23295,N_22763,N_22564);
nand U23296 (N_23296,N_22793,N_22573);
nand U23297 (N_23297,N_22862,N_22962);
or U23298 (N_23298,N_22683,N_22976);
nor U23299 (N_23299,N_22975,N_22939);
nand U23300 (N_23300,N_22951,N_22853);
or U23301 (N_23301,N_22688,N_22994);
nand U23302 (N_23302,N_22840,N_22669);
nor U23303 (N_23303,N_22637,N_22687);
nand U23304 (N_23304,N_22620,N_22958);
nand U23305 (N_23305,N_22839,N_22829);
nor U23306 (N_23306,N_22542,N_22531);
nor U23307 (N_23307,N_22980,N_22731);
nor U23308 (N_23308,N_22535,N_22908);
nand U23309 (N_23309,N_22715,N_22636);
xnor U23310 (N_23310,N_22739,N_22835);
nor U23311 (N_23311,N_22825,N_22703);
and U23312 (N_23312,N_22591,N_22526);
nand U23313 (N_23313,N_22995,N_22532);
and U23314 (N_23314,N_22840,N_22784);
nor U23315 (N_23315,N_22828,N_22917);
or U23316 (N_23316,N_22920,N_22834);
xnor U23317 (N_23317,N_22881,N_22540);
xnor U23318 (N_23318,N_22557,N_22821);
xor U23319 (N_23319,N_22747,N_22978);
nor U23320 (N_23320,N_22681,N_22514);
and U23321 (N_23321,N_22563,N_22772);
nand U23322 (N_23322,N_22579,N_22996);
nand U23323 (N_23323,N_22852,N_22541);
xor U23324 (N_23324,N_22641,N_22752);
and U23325 (N_23325,N_22741,N_22882);
nand U23326 (N_23326,N_22591,N_22688);
or U23327 (N_23327,N_22723,N_22697);
and U23328 (N_23328,N_22537,N_22663);
and U23329 (N_23329,N_22552,N_22722);
nand U23330 (N_23330,N_22560,N_22709);
and U23331 (N_23331,N_22648,N_22733);
nor U23332 (N_23332,N_22564,N_22972);
or U23333 (N_23333,N_22972,N_22947);
and U23334 (N_23334,N_22868,N_22928);
nand U23335 (N_23335,N_22507,N_22557);
nor U23336 (N_23336,N_22836,N_22650);
and U23337 (N_23337,N_22662,N_22750);
and U23338 (N_23338,N_22911,N_22917);
or U23339 (N_23339,N_22830,N_22722);
and U23340 (N_23340,N_22711,N_22530);
nand U23341 (N_23341,N_22798,N_22767);
and U23342 (N_23342,N_22873,N_22950);
xor U23343 (N_23343,N_22854,N_22756);
xnor U23344 (N_23344,N_22759,N_22732);
nor U23345 (N_23345,N_22966,N_22796);
nand U23346 (N_23346,N_22558,N_22781);
nand U23347 (N_23347,N_22667,N_22578);
xor U23348 (N_23348,N_22779,N_22813);
and U23349 (N_23349,N_22795,N_22758);
xnor U23350 (N_23350,N_22748,N_22960);
and U23351 (N_23351,N_22841,N_22670);
nor U23352 (N_23352,N_22875,N_22687);
or U23353 (N_23353,N_22846,N_22916);
or U23354 (N_23354,N_22648,N_22975);
nand U23355 (N_23355,N_22669,N_22777);
nand U23356 (N_23356,N_22697,N_22656);
or U23357 (N_23357,N_22694,N_22878);
xnor U23358 (N_23358,N_22687,N_22929);
xor U23359 (N_23359,N_22595,N_22752);
nor U23360 (N_23360,N_22687,N_22827);
nand U23361 (N_23361,N_22618,N_22975);
and U23362 (N_23362,N_22812,N_22690);
xor U23363 (N_23363,N_22808,N_22654);
nor U23364 (N_23364,N_22785,N_22710);
nand U23365 (N_23365,N_22667,N_22950);
xnor U23366 (N_23366,N_22800,N_22941);
and U23367 (N_23367,N_22682,N_22593);
nand U23368 (N_23368,N_22605,N_22779);
xnor U23369 (N_23369,N_22937,N_22976);
or U23370 (N_23370,N_22570,N_22578);
xnor U23371 (N_23371,N_22959,N_22849);
nand U23372 (N_23372,N_22977,N_22915);
nand U23373 (N_23373,N_22612,N_22859);
xor U23374 (N_23374,N_22584,N_22652);
and U23375 (N_23375,N_22815,N_22771);
or U23376 (N_23376,N_22925,N_22689);
or U23377 (N_23377,N_22757,N_22616);
nand U23378 (N_23378,N_22577,N_22982);
xnor U23379 (N_23379,N_22568,N_22810);
and U23380 (N_23380,N_22520,N_22552);
nor U23381 (N_23381,N_22672,N_22799);
xnor U23382 (N_23382,N_22598,N_22580);
nor U23383 (N_23383,N_22847,N_22890);
or U23384 (N_23384,N_22707,N_22559);
nand U23385 (N_23385,N_22711,N_22729);
xnor U23386 (N_23386,N_22766,N_22504);
and U23387 (N_23387,N_22566,N_22802);
nor U23388 (N_23388,N_22532,N_22671);
and U23389 (N_23389,N_22695,N_22576);
nor U23390 (N_23390,N_22935,N_22528);
nand U23391 (N_23391,N_22906,N_22863);
and U23392 (N_23392,N_22923,N_22765);
xor U23393 (N_23393,N_22903,N_22692);
and U23394 (N_23394,N_22975,N_22559);
or U23395 (N_23395,N_22726,N_22573);
nor U23396 (N_23396,N_22979,N_22582);
xnor U23397 (N_23397,N_22659,N_22944);
nor U23398 (N_23398,N_22642,N_22632);
nand U23399 (N_23399,N_22764,N_22528);
xnor U23400 (N_23400,N_22553,N_22537);
nand U23401 (N_23401,N_22523,N_22507);
xnor U23402 (N_23402,N_22948,N_22849);
nand U23403 (N_23403,N_22869,N_22652);
nand U23404 (N_23404,N_22611,N_22872);
or U23405 (N_23405,N_22942,N_22712);
nor U23406 (N_23406,N_22542,N_22751);
or U23407 (N_23407,N_22866,N_22885);
nor U23408 (N_23408,N_22750,N_22623);
nand U23409 (N_23409,N_22545,N_22810);
or U23410 (N_23410,N_22642,N_22816);
nand U23411 (N_23411,N_22535,N_22994);
nor U23412 (N_23412,N_22894,N_22578);
or U23413 (N_23413,N_22618,N_22907);
nand U23414 (N_23414,N_22542,N_22692);
nor U23415 (N_23415,N_22700,N_22738);
nor U23416 (N_23416,N_22693,N_22601);
and U23417 (N_23417,N_22875,N_22605);
xor U23418 (N_23418,N_22636,N_22832);
and U23419 (N_23419,N_22868,N_22547);
xor U23420 (N_23420,N_22840,N_22947);
nor U23421 (N_23421,N_22881,N_22996);
nor U23422 (N_23422,N_22888,N_22629);
and U23423 (N_23423,N_22915,N_22858);
nand U23424 (N_23424,N_22637,N_22758);
or U23425 (N_23425,N_22645,N_22886);
or U23426 (N_23426,N_22884,N_22924);
and U23427 (N_23427,N_22546,N_22512);
or U23428 (N_23428,N_22511,N_22771);
nand U23429 (N_23429,N_22544,N_22800);
nor U23430 (N_23430,N_22840,N_22793);
nor U23431 (N_23431,N_22585,N_22583);
nand U23432 (N_23432,N_22555,N_22695);
nand U23433 (N_23433,N_22840,N_22526);
and U23434 (N_23434,N_22635,N_22815);
nand U23435 (N_23435,N_22696,N_22669);
nand U23436 (N_23436,N_22984,N_22709);
or U23437 (N_23437,N_22898,N_22573);
and U23438 (N_23438,N_22783,N_22654);
or U23439 (N_23439,N_22607,N_22806);
nor U23440 (N_23440,N_22684,N_22525);
or U23441 (N_23441,N_22894,N_22503);
nor U23442 (N_23442,N_22833,N_22952);
nor U23443 (N_23443,N_22787,N_22950);
or U23444 (N_23444,N_22975,N_22581);
and U23445 (N_23445,N_22541,N_22841);
or U23446 (N_23446,N_22820,N_22778);
and U23447 (N_23447,N_22612,N_22966);
or U23448 (N_23448,N_22880,N_22814);
nor U23449 (N_23449,N_22757,N_22572);
nor U23450 (N_23450,N_22768,N_22825);
nand U23451 (N_23451,N_22969,N_22616);
or U23452 (N_23452,N_22753,N_22801);
nor U23453 (N_23453,N_22887,N_22529);
xor U23454 (N_23454,N_22540,N_22939);
and U23455 (N_23455,N_22624,N_22631);
or U23456 (N_23456,N_22682,N_22568);
nand U23457 (N_23457,N_22856,N_22713);
nand U23458 (N_23458,N_22566,N_22612);
nor U23459 (N_23459,N_22734,N_22895);
xor U23460 (N_23460,N_22930,N_22993);
xnor U23461 (N_23461,N_22982,N_22818);
nor U23462 (N_23462,N_22551,N_22949);
nor U23463 (N_23463,N_22584,N_22826);
and U23464 (N_23464,N_22906,N_22771);
and U23465 (N_23465,N_22639,N_22537);
and U23466 (N_23466,N_22547,N_22570);
and U23467 (N_23467,N_22766,N_22847);
and U23468 (N_23468,N_22807,N_22896);
nor U23469 (N_23469,N_22871,N_22857);
nor U23470 (N_23470,N_22834,N_22693);
nor U23471 (N_23471,N_22896,N_22797);
xor U23472 (N_23472,N_22987,N_22652);
or U23473 (N_23473,N_22923,N_22684);
nor U23474 (N_23474,N_22955,N_22986);
or U23475 (N_23475,N_22859,N_22794);
nor U23476 (N_23476,N_22928,N_22851);
or U23477 (N_23477,N_22893,N_22831);
xnor U23478 (N_23478,N_22616,N_22863);
nand U23479 (N_23479,N_22854,N_22882);
nor U23480 (N_23480,N_22871,N_22671);
or U23481 (N_23481,N_22605,N_22943);
and U23482 (N_23482,N_22917,N_22585);
xnor U23483 (N_23483,N_22707,N_22976);
nand U23484 (N_23484,N_22907,N_22739);
nand U23485 (N_23485,N_22880,N_22951);
xor U23486 (N_23486,N_22983,N_22898);
or U23487 (N_23487,N_22670,N_22749);
nand U23488 (N_23488,N_22591,N_22636);
and U23489 (N_23489,N_22659,N_22598);
nand U23490 (N_23490,N_22696,N_22600);
xor U23491 (N_23491,N_22603,N_22728);
xor U23492 (N_23492,N_22629,N_22900);
nor U23493 (N_23493,N_22678,N_22979);
nor U23494 (N_23494,N_22725,N_22687);
xor U23495 (N_23495,N_22571,N_22741);
or U23496 (N_23496,N_22619,N_22654);
xor U23497 (N_23497,N_22781,N_22516);
nor U23498 (N_23498,N_22622,N_22554);
nand U23499 (N_23499,N_22584,N_22913);
or U23500 (N_23500,N_23287,N_23219);
or U23501 (N_23501,N_23323,N_23116);
or U23502 (N_23502,N_23083,N_23076);
and U23503 (N_23503,N_23129,N_23303);
nor U23504 (N_23504,N_23145,N_23274);
nor U23505 (N_23505,N_23078,N_23049);
nand U23506 (N_23506,N_23086,N_23029);
nor U23507 (N_23507,N_23241,N_23342);
or U23508 (N_23508,N_23189,N_23109);
and U23509 (N_23509,N_23305,N_23120);
nand U23510 (N_23510,N_23061,N_23039);
xnor U23511 (N_23511,N_23392,N_23420);
xnor U23512 (N_23512,N_23495,N_23073);
nand U23513 (N_23513,N_23258,N_23063);
nand U23514 (N_23514,N_23020,N_23385);
nand U23515 (N_23515,N_23113,N_23164);
and U23516 (N_23516,N_23177,N_23101);
nor U23517 (N_23517,N_23438,N_23325);
and U23518 (N_23518,N_23348,N_23494);
xor U23519 (N_23519,N_23004,N_23077);
and U23520 (N_23520,N_23210,N_23140);
or U23521 (N_23521,N_23288,N_23005);
xor U23522 (N_23522,N_23341,N_23463);
xor U23523 (N_23523,N_23355,N_23103);
nand U23524 (N_23524,N_23184,N_23472);
or U23525 (N_23525,N_23409,N_23406);
and U23526 (N_23526,N_23006,N_23315);
nand U23527 (N_23527,N_23448,N_23011);
xnor U23528 (N_23528,N_23285,N_23293);
and U23529 (N_23529,N_23460,N_23324);
and U23530 (N_23530,N_23070,N_23334);
nand U23531 (N_23531,N_23223,N_23379);
and U23532 (N_23532,N_23474,N_23021);
and U23533 (N_23533,N_23319,N_23253);
nor U23534 (N_23534,N_23405,N_23037);
xor U23535 (N_23535,N_23138,N_23097);
and U23536 (N_23536,N_23298,N_23117);
or U23537 (N_23537,N_23336,N_23008);
xnor U23538 (N_23538,N_23240,N_23060);
and U23539 (N_23539,N_23173,N_23216);
or U23540 (N_23540,N_23407,N_23374);
nor U23541 (N_23541,N_23149,N_23125);
xnor U23542 (N_23542,N_23382,N_23032);
xor U23543 (N_23543,N_23304,N_23176);
or U23544 (N_23544,N_23003,N_23330);
nor U23545 (N_23545,N_23200,N_23335);
and U23546 (N_23546,N_23014,N_23433);
and U23547 (N_23547,N_23134,N_23136);
xnor U23548 (N_23548,N_23419,N_23050);
nor U23549 (N_23549,N_23269,N_23312);
nand U23550 (N_23550,N_23192,N_23318);
or U23551 (N_23551,N_23111,N_23390);
or U23552 (N_23552,N_23168,N_23194);
nand U23553 (N_23553,N_23163,N_23297);
or U23554 (N_23554,N_23327,N_23175);
xor U23555 (N_23555,N_23126,N_23055);
and U23556 (N_23556,N_23443,N_23337);
nor U23557 (N_23557,N_23350,N_23244);
nand U23558 (N_23558,N_23371,N_23208);
or U23559 (N_23559,N_23262,N_23307);
xnor U23560 (N_23560,N_23224,N_23453);
xor U23561 (N_23561,N_23493,N_23442);
nor U23562 (N_23562,N_23461,N_23480);
and U23563 (N_23563,N_23127,N_23187);
and U23564 (N_23564,N_23038,N_23378);
and U23565 (N_23565,N_23071,N_23267);
and U23566 (N_23566,N_23256,N_23081);
nand U23567 (N_23567,N_23423,N_23190);
or U23568 (N_23568,N_23230,N_23326);
and U23569 (N_23569,N_23166,N_23376);
nor U23570 (N_23570,N_23220,N_23135);
nand U23571 (N_23571,N_23024,N_23012);
xor U23572 (N_23572,N_23377,N_23479);
or U23573 (N_23573,N_23048,N_23380);
or U23574 (N_23574,N_23273,N_23051);
nand U23575 (N_23575,N_23160,N_23246);
or U23576 (N_23576,N_23046,N_23308);
xnor U23577 (N_23577,N_23485,N_23491);
and U23578 (N_23578,N_23096,N_23345);
xnor U23579 (N_23579,N_23291,N_23232);
nor U23580 (N_23580,N_23384,N_23344);
xnor U23581 (N_23581,N_23432,N_23064);
xor U23582 (N_23582,N_23088,N_23434);
nand U23583 (N_23583,N_23393,N_23496);
and U23584 (N_23584,N_23261,N_23186);
nand U23585 (N_23585,N_23375,N_23180);
nor U23586 (N_23586,N_23457,N_23114);
nand U23587 (N_23587,N_23248,N_23497);
and U23588 (N_23588,N_23047,N_23358);
xnor U23589 (N_23589,N_23475,N_23022);
nor U23590 (N_23590,N_23027,N_23329);
and U23591 (N_23591,N_23320,N_23229);
or U23592 (N_23592,N_23306,N_23132);
xnor U23593 (N_23593,N_23042,N_23389);
and U23594 (N_23594,N_23452,N_23340);
and U23595 (N_23595,N_23013,N_23123);
nor U23596 (N_23596,N_23483,N_23310);
xor U23597 (N_23597,N_23359,N_23015);
nand U23598 (N_23598,N_23299,N_23365);
nor U23599 (N_23599,N_23399,N_23473);
xor U23600 (N_23600,N_23467,N_23322);
nand U23601 (N_23601,N_23338,N_23198);
xor U23602 (N_23602,N_23281,N_23417);
xnor U23603 (N_23603,N_23272,N_23143);
nor U23604 (N_23604,N_23002,N_23105);
and U23605 (N_23605,N_23162,N_23201);
nand U23606 (N_23606,N_23155,N_23196);
xnor U23607 (N_23607,N_23362,N_23440);
xnor U23608 (N_23608,N_23498,N_23130);
nor U23609 (N_23609,N_23209,N_23302);
and U23610 (N_23610,N_23279,N_23346);
and U23611 (N_23611,N_23441,N_23300);
nand U23612 (N_23612,N_23368,N_23489);
or U23613 (N_23613,N_23301,N_23482);
or U23614 (N_23614,N_23481,N_23159);
nor U23615 (N_23615,N_23041,N_23369);
nor U23616 (N_23616,N_23152,N_23429);
xnor U23617 (N_23617,N_23094,N_23199);
nor U23618 (N_23618,N_23424,N_23131);
nand U23619 (N_23619,N_23028,N_23079);
and U23620 (N_23620,N_23144,N_23353);
nand U23621 (N_23621,N_23314,N_23215);
xor U23622 (N_23622,N_23084,N_23275);
nor U23623 (N_23623,N_23148,N_23197);
and U23624 (N_23624,N_23099,N_23454);
xor U23625 (N_23625,N_23373,N_23328);
nand U23626 (N_23626,N_23278,N_23431);
nand U23627 (N_23627,N_23062,N_23477);
nand U23628 (N_23628,N_23191,N_23107);
and U23629 (N_23629,N_23091,N_23309);
nor U23630 (N_23630,N_23052,N_23234);
nand U23631 (N_23631,N_23255,N_23277);
xnor U23632 (N_23632,N_23360,N_23182);
nand U23633 (N_23633,N_23231,N_23030);
nor U23634 (N_23634,N_23110,N_23239);
nand U23635 (N_23635,N_23435,N_23263);
nor U23636 (N_23636,N_23124,N_23080);
or U23637 (N_23637,N_23236,N_23331);
xor U23638 (N_23638,N_23218,N_23252);
and U23639 (N_23639,N_23092,N_23391);
xor U23640 (N_23640,N_23415,N_23413);
and U23641 (N_23641,N_23235,N_23017);
and U23642 (N_23642,N_23311,N_23068);
xor U23643 (N_23643,N_23188,N_23313);
xnor U23644 (N_23644,N_23082,N_23447);
nand U23645 (N_23645,N_23221,N_23490);
xor U23646 (N_23646,N_23402,N_23150);
xor U23647 (N_23647,N_23427,N_23464);
xor U23648 (N_23648,N_23400,N_23458);
nand U23649 (N_23649,N_23478,N_23364);
or U23650 (N_23650,N_23172,N_23245);
or U23651 (N_23651,N_23466,N_23445);
nand U23652 (N_23652,N_23260,N_23025);
or U23653 (N_23653,N_23167,N_23247);
or U23654 (N_23654,N_23403,N_23211);
xnor U23655 (N_23655,N_23207,N_23054);
nand U23656 (N_23656,N_23156,N_23356);
or U23657 (N_23657,N_23171,N_23492);
or U23658 (N_23658,N_23087,N_23339);
and U23659 (N_23659,N_23225,N_23426);
or U23660 (N_23660,N_23372,N_23268);
xnor U23661 (N_23661,N_23100,N_23286);
nand U23662 (N_23662,N_23000,N_23416);
or U23663 (N_23663,N_23459,N_23456);
xnor U23664 (N_23664,N_23462,N_23161);
xor U23665 (N_23665,N_23465,N_23468);
nand U23666 (N_23666,N_23106,N_23007);
and U23667 (N_23667,N_23398,N_23238);
nor U23668 (N_23668,N_23271,N_23095);
nor U23669 (N_23669,N_23059,N_23137);
or U23670 (N_23670,N_23093,N_23251);
and U23671 (N_23671,N_23284,N_23031);
nor U23672 (N_23672,N_23484,N_23072);
xnor U23673 (N_23673,N_23019,N_23089);
and U23674 (N_23674,N_23254,N_23292);
nor U23675 (N_23675,N_23226,N_23469);
xor U23676 (N_23676,N_23488,N_23009);
and U23677 (N_23677,N_23410,N_23001);
nor U23678 (N_23678,N_23090,N_23455);
nand U23679 (N_23679,N_23316,N_23058);
nand U23680 (N_23680,N_23499,N_23010);
and U23681 (N_23681,N_23444,N_23411);
xor U23682 (N_23682,N_23449,N_23151);
xnor U23683 (N_23683,N_23035,N_23446);
nor U23684 (N_23684,N_23233,N_23056);
and U23685 (N_23685,N_23066,N_23396);
or U23686 (N_23686,N_23178,N_23237);
xor U23687 (N_23687,N_23053,N_23158);
nand U23688 (N_23688,N_23264,N_23206);
and U23689 (N_23689,N_23205,N_23425);
nand U23690 (N_23690,N_23487,N_23265);
nand U23691 (N_23691,N_23193,N_23295);
or U23692 (N_23692,N_23098,N_23257);
xor U23693 (N_23693,N_23115,N_23333);
xor U23694 (N_23694,N_23141,N_23227);
xnor U23695 (N_23695,N_23486,N_23352);
or U23696 (N_23696,N_23383,N_23276);
nor U23697 (N_23697,N_23033,N_23034);
nor U23698 (N_23698,N_23283,N_23018);
nand U23699 (N_23699,N_23397,N_23289);
or U23700 (N_23700,N_23386,N_23119);
or U23701 (N_23701,N_23349,N_23065);
xor U23702 (N_23702,N_23153,N_23204);
nand U23703 (N_23703,N_23451,N_23418);
nand U23704 (N_23704,N_23112,N_23074);
and U23705 (N_23705,N_23351,N_23170);
nor U23706 (N_23706,N_23183,N_23361);
or U23707 (N_23707,N_23118,N_23450);
xnor U23708 (N_23708,N_23179,N_23213);
and U23709 (N_23709,N_23354,N_23147);
nand U23710 (N_23710,N_23282,N_23228);
xnor U23711 (N_23711,N_23057,N_23470);
xor U23712 (N_23712,N_23214,N_23102);
or U23713 (N_23713,N_23357,N_23243);
nor U23714 (N_23714,N_23154,N_23185);
or U23715 (N_23715,N_23121,N_23174);
and U23716 (N_23716,N_23157,N_23045);
or U23717 (N_23717,N_23040,N_23142);
nor U23718 (N_23718,N_23067,N_23044);
xor U23719 (N_23719,N_23290,N_23439);
xnor U23720 (N_23720,N_23343,N_23133);
nand U23721 (N_23721,N_23169,N_23075);
xnor U23722 (N_23722,N_23165,N_23404);
or U23723 (N_23723,N_23395,N_23437);
xnor U23724 (N_23724,N_23266,N_23036);
or U23725 (N_23725,N_23128,N_23394);
nor U23726 (N_23726,N_23222,N_23436);
and U23727 (N_23727,N_23367,N_23321);
xor U23728 (N_23728,N_23270,N_23069);
nor U23729 (N_23729,N_23408,N_23043);
nand U23730 (N_23730,N_23250,N_23412);
or U23731 (N_23731,N_23217,N_23108);
and U23732 (N_23732,N_23422,N_23122);
nand U23733 (N_23733,N_23026,N_23249);
and U23734 (N_23734,N_23366,N_23414);
and U23735 (N_23735,N_23317,N_23181);
nor U23736 (N_23736,N_23202,N_23085);
nand U23737 (N_23737,N_23370,N_23139);
nand U23738 (N_23738,N_23296,N_23388);
nor U23739 (N_23739,N_23104,N_23387);
nand U23740 (N_23740,N_23347,N_23428);
nor U23741 (N_23741,N_23146,N_23476);
or U23742 (N_23742,N_23332,N_23259);
and U23743 (N_23743,N_23421,N_23203);
or U23744 (N_23744,N_23381,N_23242);
xor U23745 (N_23745,N_23280,N_23016);
xor U23746 (N_23746,N_23195,N_23471);
or U23747 (N_23747,N_23023,N_23294);
xnor U23748 (N_23748,N_23430,N_23401);
nor U23749 (N_23749,N_23363,N_23212);
and U23750 (N_23750,N_23118,N_23142);
xor U23751 (N_23751,N_23071,N_23080);
xor U23752 (N_23752,N_23281,N_23025);
xor U23753 (N_23753,N_23278,N_23181);
nor U23754 (N_23754,N_23324,N_23307);
xnor U23755 (N_23755,N_23300,N_23001);
nor U23756 (N_23756,N_23357,N_23201);
nor U23757 (N_23757,N_23198,N_23008);
and U23758 (N_23758,N_23338,N_23381);
and U23759 (N_23759,N_23199,N_23490);
or U23760 (N_23760,N_23254,N_23052);
nor U23761 (N_23761,N_23161,N_23281);
or U23762 (N_23762,N_23497,N_23090);
or U23763 (N_23763,N_23023,N_23362);
nand U23764 (N_23764,N_23147,N_23291);
nand U23765 (N_23765,N_23147,N_23267);
or U23766 (N_23766,N_23264,N_23473);
xnor U23767 (N_23767,N_23228,N_23362);
xnor U23768 (N_23768,N_23138,N_23108);
or U23769 (N_23769,N_23336,N_23357);
or U23770 (N_23770,N_23488,N_23281);
nand U23771 (N_23771,N_23464,N_23100);
nand U23772 (N_23772,N_23171,N_23037);
nand U23773 (N_23773,N_23456,N_23234);
or U23774 (N_23774,N_23195,N_23028);
or U23775 (N_23775,N_23293,N_23072);
xor U23776 (N_23776,N_23082,N_23380);
nand U23777 (N_23777,N_23022,N_23127);
or U23778 (N_23778,N_23399,N_23120);
xor U23779 (N_23779,N_23401,N_23050);
or U23780 (N_23780,N_23175,N_23362);
nand U23781 (N_23781,N_23159,N_23164);
xor U23782 (N_23782,N_23380,N_23229);
nand U23783 (N_23783,N_23469,N_23000);
or U23784 (N_23784,N_23088,N_23278);
xor U23785 (N_23785,N_23094,N_23305);
xnor U23786 (N_23786,N_23206,N_23237);
and U23787 (N_23787,N_23346,N_23331);
nand U23788 (N_23788,N_23193,N_23145);
or U23789 (N_23789,N_23272,N_23238);
or U23790 (N_23790,N_23307,N_23068);
nor U23791 (N_23791,N_23389,N_23062);
and U23792 (N_23792,N_23023,N_23351);
xor U23793 (N_23793,N_23392,N_23486);
xnor U23794 (N_23794,N_23369,N_23099);
nor U23795 (N_23795,N_23139,N_23158);
nand U23796 (N_23796,N_23029,N_23066);
or U23797 (N_23797,N_23398,N_23133);
and U23798 (N_23798,N_23033,N_23427);
nor U23799 (N_23799,N_23219,N_23496);
nor U23800 (N_23800,N_23231,N_23452);
nand U23801 (N_23801,N_23441,N_23308);
xnor U23802 (N_23802,N_23251,N_23082);
xnor U23803 (N_23803,N_23349,N_23347);
nor U23804 (N_23804,N_23147,N_23130);
xnor U23805 (N_23805,N_23178,N_23458);
xnor U23806 (N_23806,N_23138,N_23070);
xnor U23807 (N_23807,N_23424,N_23427);
or U23808 (N_23808,N_23480,N_23212);
and U23809 (N_23809,N_23102,N_23424);
or U23810 (N_23810,N_23144,N_23406);
or U23811 (N_23811,N_23438,N_23369);
nor U23812 (N_23812,N_23342,N_23367);
and U23813 (N_23813,N_23470,N_23347);
nand U23814 (N_23814,N_23236,N_23460);
and U23815 (N_23815,N_23404,N_23074);
nand U23816 (N_23816,N_23077,N_23068);
xnor U23817 (N_23817,N_23310,N_23037);
nand U23818 (N_23818,N_23189,N_23202);
or U23819 (N_23819,N_23018,N_23177);
xor U23820 (N_23820,N_23496,N_23006);
xnor U23821 (N_23821,N_23064,N_23119);
or U23822 (N_23822,N_23269,N_23418);
and U23823 (N_23823,N_23446,N_23029);
and U23824 (N_23824,N_23497,N_23264);
nand U23825 (N_23825,N_23059,N_23105);
or U23826 (N_23826,N_23064,N_23006);
and U23827 (N_23827,N_23033,N_23277);
xnor U23828 (N_23828,N_23068,N_23408);
and U23829 (N_23829,N_23047,N_23326);
nand U23830 (N_23830,N_23459,N_23342);
nor U23831 (N_23831,N_23457,N_23379);
xor U23832 (N_23832,N_23061,N_23282);
nor U23833 (N_23833,N_23433,N_23372);
nor U23834 (N_23834,N_23461,N_23232);
and U23835 (N_23835,N_23030,N_23169);
nor U23836 (N_23836,N_23145,N_23120);
nor U23837 (N_23837,N_23477,N_23029);
and U23838 (N_23838,N_23140,N_23226);
xnor U23839 (N_23839,N_23319,N_23242);
or U23840 (N_23840,N_23445,N_23437);
nor U23841 (N_23841,N_23281,N_23268);
xnor U23842 (N_23842,N_23064,N_23226);
nand U23843 (N_23843,N_23323,N_23095);
nor U23844 (N_23844,N_23235,N_23495);
nand U23845 (N_23845,N_23029,N_23226);
and U23846 (N_23846,N_23366,N_23342);
nand U23847 (N_23847,N_23351,N_23365);
or U23848 (N_23848,N_23235,N_23146);
and U23849 (N_23849,N_23420,N_23097);
nand U23850 (N_23850,N_23029,N_23273);
xnor U23851 (N_23851,N_23073,N_23023);
xnor U23852 (N_23852,N_23111,N_23219);
nand U23853 (N_23853,N_23383,N_23051);
xnor U23854 (N_23854,N_23166,N_23454);
and U23855 (N_23855,N_23246,N_23149);
nor U23856 (N_23856,N_23049,N_23120);
nand U23857 (N_23857,N_23152,N_23045);
nand U23858 (N_23858,N_23165,N_23191);
and U23859 (N_23859,N_23016,N_23070);
nor U23860 (N_23860,N_23259,N_23049);
or U23861 (N_23861,N_23307,N_23425);
and U23862 (N_23862,N_23157,N_23490);
or U23863 (N_23863,N_23232,N_23478);
nand U23864 (N_23864,N_23059,N_23335);
or U23865 (N_23865,N_23459,N_23057);
xor U23866 (N_23866,N_23075,N_23285);
or U23867 (N_23867,N_23154,N_23067);
nor U23868 (N_23868,N_23459,N_23174);
or U23869 (N_23869,N_23259,N_23199);
and U23870 (N_23870,N_23209,N_23330);
or U23871 (N_23871,N_23492,N_23286);
nand U23872 (N_23872,N_23302,N_23495);
xnor U23873 (N_23873,N_23132,N_23271);
xnor U23874 (N_23874,N_23297,N_23014);
xnor U23875 (N_23875,N_23406,N_23389);
xor U23876 (N_23876,N_23185,N_23121);
nand U23877 (N_23877,N_23136,N_23237);
or U23878 (N_23878,N_23161,N_23249);
xor U23879 (N_23879,N_23359,N_23324);
and U23880 (N_23880,N_23096,N_23056);
xnor U23881 (N_23881,N_23442,N_23007);
or U23882 (N_23882,N_23061,N_23430);
nor U23883 (N_23883,N_23253,N_23413);
nor U23884 (N_23884,N_23471,N_23315);
or U23885 (N_23885,N_23478,N_23318);
and U23886 (N_23886,N_23434,N_23445);
xnor U23887 (N_23887,N_23098,N_23350);
or U23888 (N_23888,N_23444,N_23099);
nand U23889 (N_23889,N_23450,N_23079);
nand U23890 (N_23890,N_23324,N_23123);
nand U23891 (N_23891,N_23084,N_23165);
nor U23892 (N_23892,N_23456,N_23274);
and U23893 (N_23893,N_23031,N_23053);
or U23894 (N_23894,N_23085,N_23329);
and U23895 (N_23895,N_23148,N_23129);
xnor U23896 (N_23896,N_23462,N_23094);
xnor U23897 (N_23897,N_23090,N_23491);
xnor U23898 (N_23898,N_23402,N_23188);
xor U23899 (N_23899,N_23421,N_23147);
or U23900 (N_23900,N_23239,N_23274);
nor U23901 (N_23901,N_23236,N_23498);
nor U23902 (N_23902,N_23080,N_23275);
xnor U23903 (N_23903,N_23042,N_23256);
nor U23904 (N_23904,N_23441,N_23266);
and U23905 (N_23905,N_23034,N_23250);
or U23906 (N_23906,N_23436,N_23006);
and U23907 (N_23907,N_23446,N_23360);
or U23908 (N_23908,N_23074,N_23202);
and U23909 (N_23909,N_23447,N_23361);
nand U23910 (N_23910,N_23057,N_23333);
nand U23911 (N_23911,N_23252,N_23057);
nor U23912 (N_23912,N_23427,N_23060);
nor U23913 (N_23913,N_23074,N_23118);
nand U23914 (N_23914,N_23044,N_23434);
nand U23915 (N_23915,N_23310,N_23244);
or U23916 (N_23916,N_23310,N_23025);
nand U23917 (N_23917,N_23336,N_23074);
xor U23918 (N_23918,N_23270,N_23300);
and U23919 (N_23919,N_23170,N_23091);
or U23920 (N_23920,N_23347,N_23006);
nor U23921 (N_23921,N_23124,N_23359);
xor U23922 (N_23922,N_23031,N_23291);
xor U23923 (N_23923,N_23393,N_23286);
and U23924 (N_23924,N_23348,N_23126);
xnor U23925 (N_23925,N_23473,N_23133);
or U23926 (N_23926,N_23253,N_23338);
or U23927 (N_23927,N_23497,N_23318);
nor U23928 (N_23928,N_23372,N_23412);
xor U23929 (N_23929,N_23165,N_23371);
nor U23930 (N_23930,N_23478,N_23052);
xor U23931 (N_23931,N_23225,N_23193);
and U23932 (N_23932,N_23043,N_23273);
or U23933 (N_23933,N_23340,N_23146);
and U23934 (N_23934,N_23069,N_23213);
and U23935 (N_23935,N_23384,N_23094);
nand U23936 (N_23936,N_23178,N_23109);
nand U23937 (N_23937,N_23195,N_23025);
nand U23938 (N_23938,N_23440,N_23153);
nand U23939 (N_23939,N_23368,N_23100);
nor U23940 (N_23940,N_23269,N_23338);
nand U23941 (N_23941,N_23278,N_23332);
xor U23942 (N_23942,N_23079,N_23193);
nor U23943 (N_23943,N_23426,N_23150);
xor U23944 (N_23944,N_23413,N_23464);
and U23945 (N_23945,N_23399,N_23274);
nor U23946 (N_23946,N_23313,N_23243);
or U23947 (N_23947,N_23104,N_23027);
and U23948 (N_23948,N_23266,N_23173);
xnor U23949 (N_23949,N_23206,N_23137);
or U23950 (N_23950,N_23139,N_23197);
nor U23951 (N_23951,N_23465,N_23398);
or U23952 (N_23952,N_23451,N_23296);
nor U23953 (N_23953,N_23210,N_23112);
nor U23954 (N_23954,N_23394,N_23163);
nor U23955 (N_23955,N_23055,N_23239);
and U23956 (N_23956,N_23273,N_23190);
nand U23957 (N_23957,N_23155,N_23331);
and U23958 (N_23958,N_23150,N_23337);
nor U23959 (N_23959,N_23412,N_23247);
nor U23960 (N_23960,N_23150,N_23129);
xnor U23961 (N_23961,N_23475,N_23498);
or U23962 (N_23962,N_23164,N_23226);
nor U23963 (N_23963,N_23314,N_23323);
and U23964 (N_23964,N_23362,N_23407);
and U23965 (N_23965,N_23164,N_23452);
or U23966 (N_23966,N_23018,N_23198);
nand U23967 (N_23967,N_23486,N_23109);
and U23968 (N_23968,N_23273,N_23260);
or U23969 (N_23969,N_23253,N_23062);
and U23970 (N_23970,N_23107,N_23415);
nor U23971 (N_23971,N_23013,N_23112);
and U23972 (N_23972,N_23484,N_23307);
xor U23973 (N_23973,N_23475,N_23126);
or U23974 (N_23974,N_23223,N_23318);
xnor U23975 (N_23975,N_23324,N_23136);
nor U23976 (N_23976,N_23346,N_23408);
and U23977 (N_23977,N_23220,N_23312);
and U23978 (N_23978,N_23352,N_23319);
nand U23979 (N_23979,N_23387,N_23368);
xor U23980 (N_23980,N_23354,N_23488);
nor U23981 (N_23981,N_23115,N_23391);
xor U23982 (N_23982,N_23491,N_23436);
or U23983 (N_23983,N_23475,N_23292);
nand U23984 (N_23984,N_23469,N_23337);
and U23985 (N_23985,N_23172,N_23192);
nor U23986 (N_23986,N_23298,N_23064);
and U23987 (N_23987,N_23281,N_23153);
and U23988 (N_23988,N_23183,N_23014);
xor U23989 (N_23989,N_23150,N_23458);
and U23990 (N_23990,N_23462,N_23459);
xor U23991 (N_23991,N_23261,N_23456);
or U23992 (N_23992,N_23251,N_23278);
nor U23993 (N_23993,N_23486,N_23444);
xnor U23994 (N_23994,N_23306,N_23151);
nor U23995 (N_23995,N_23303,N_23262);
or U23996 (N_23996,N_23366,N_23438);
and U23997 (N_23997,N_23441,N_23470);
nand U23998 (N_23998,N_23115,N_23492);
nand U23999 (N_23999,N_23496,N_23132);
xor U24000 (N_24000,N_23699,N_23783);
and U24001 (N_24001,N_23752,N_23883);
nor U24002 (N_24002,N_23858,N_23599);
or U24003 (N_24003,N_23618,N_23712);
nor U24004 (N_24004,N_23585,N_23732);
or U24005 (N_24005,N_23506,N_23844);
nor U24006 (N_24006,N_23760,N_23645);
nand U24007 (N_24007,N_23744,N_23688);
xor U24008 (N_24008,N_23829,N_23847);
and U24009 (N_24009,N_23721,N_23836);
or U24010 (N_24010,N_23708,N_23541);
xor U24011 (N_24011,N_23930,N_23872);
xor U24012 (N_24012,N_23984,N_23603);
and U24013 (N_24013,N_23908,N_23670);
nor U24014 (N_24014,N_23894,N_23631);
or U24015 (N_24015,N_23826,N_23980);
nor U24016 (N_24016,N_23500,N_23580);
xor U24017 (N_24017,N_23607,N_23503);
and U24018 (N_24018,N_23716,N_23881);
nor U24019 (N_24019,N_23973,N_23907);
nand U24020 (N_24020,N_23632,N_23562);
or U24021 (N_24021,N_23935,N_23625);
nand U24022 (N_24022,N_23568,N_23684);
and U24023 (N_24023,N_23681,N_23547);
and U24024 (N_24024,N_23651,N_23777);
xor U24025 (N_24025,N_23975,N_23751);
and U24026 (N_24026,N_23917,N_23658);
nor U24027 (N_24027,N_23834,N_23579);
and U24028 (N_24028,N_23793,N_23910);
nand U24029 (N_24029,N_23835,N_23637);
nor U24030 (N_24030,N_23617,N_23630);
nand U24031 (N_24031,N_23545,N_23671);
nand U24032 (N_24032,N_23601,N_23685);
nand U24033 (N_24033,N_23564,N_23683);
xnor U24034 (N_24034,N_23700,N_23968);
or U24035 (N_24035,N_23841,N_23845);
and U24036 (N_24036,N_23602,N_23522);
nand U24037 (N_24037,N_23556,N_23669);
nand U24038 (N_24038,N_23900,N_23635);
nand U24039 (N_24039,N_23848,N_23742);
xnor U24040 (N_24040,N_23866,N_23843);
or U24041 (N_24041,N_23726,N_23567);
nand U24042 (N_24042,N_23813,N_23689);
nor U24043 (N_24043,N_23596,N_23927);
or U24044 (N_24044,N_23513,N_23924);
nand U24045 (N_24045,N_23842,N_23583);
nor U24046 (N_24046,N_23796,N_23737);
nor U24047 (N_24047,N_23736,N_23807);
nand U24048 (N_24048,N_23855,N_23821);
nor U24049 (N_24049,N_23864,N_23548);
or U24050 (N_24050,N_23905,N_23825);
or U24051 (N_24051,N_23703,N_23901);
nor U24052 (N_24052,N_23990,N_23882);
or U24053 (N_24053,N_23823,N_23920);
and U24054 (N_24054,N_23867,N_23928);
xnor U24055 (N_24055,N_23997,N_23952);
nor U24056 (N_24056,N_23974,N_23949);
nand U24057 (N_24057,N_23819,N_23587);
xnor U24058 (N_24058,N_23717,N_23809);
nand U24059 (N_24059,N_23851,N_23509);
nor U24060 (N_24060,N_23918,N_23878);
and U24061 (N_24061,N_23730,N_23660);
nor U24062 (N_24062,N_23538,N_23902);
nand U24063 (N_24063,N_23750,N_23971);
nand U24064 (N_24064,N_23840,N_23891);
nand U24065 (N_24065,N_23923,N_23831);
and U24066 (N_24066,N_23765,N_23914);
nand U24067 (N_24067,N_23898,N_23507);
xnor U24068 (N_24068,N_23789,N_23776);
or U24069 (N_24069,N_23916,N_23536);
and U24070 (N_24070,N_23824,N_23537);
and U24071 (N_24071,N_23704,N_23856);
nand U24072 (N_24072,N_23666,N_23615);
or U24073 (N_24073,N_23738,N_23687);
and U24074 (N_24074,N_23691,N_23767);
nand U24075 (N_24075,N_23741,N_23994);
nand U24076 (N_24076,N_23609,N_23578);
nor U24077 (N_24077,N_23680,N_23868);
xnor U24078 (N_24078,N_23652,N_23711);
xor U24079 (N_24079,N_23925,N_23722);
nor U24080 (N_24080,N_23889,N_23523);
nor U24081 (N_24081,N_23991,N_23566);
xnor U24082 (N_24082,N_23644,N_23511);
nor U24083 (N_24083,N_23985,N_23954);
or U24084 (N_24084,N_23964,N_23502);
and U24085 (N_24085,N_23938,N_23701);
nor U24086 (N_24086,N_23871,N_23739);
or U24087 (N_24087,N_23664,N_23890);
nor U24088 (N_24088,N_23791,N_23608);
and U24089 (N_24089,N_23501,N_23965);
and U24090 (N_24090,N_23880,N_23944);
or U24091 (N_24091,N_23932,N_23720);
or U24092 (N_24092,N_23774,N_23758);
or U24093 (N_24093,N_23863,N_23921);
xor U24094 (N_24094,N_23960,N_23981);
and U24095 (N_24095,N_23859,N_23888);
or U24096 (N_24096,N_23621,N_23544);
or U24097 (N_24097,N_23527,N_23636);
nand U24098 (N_24098,N_23521,N_23761);
or U24099 (N_24099,N_23628,N_23942);
or U24100 (N_24100,N_23622,N_23565);
and U24101 (N_24101,N_23639,N_23860);
nand U24102 (N_24102,N_23557,N_23572);
nor U24103 (N_24103,N_23514,N_23873);
nand U24104 (N_24104,N_23972,N_23801);
xor U24105 (N_24105,N_23724,N_23592);
nor U24106 (N_24106,N_23504,N_23633);
xnor U24107 (N_24107,N_23811,N_23673);
nor U24108 (N_24108,N_23757,N_23626);
nand U24109 (N_24109,N_23728,N_23904);
nand U24110 (N_24110,N_23946,N_23933);
or U24111 (N_24111,N_23613,N_23586);
or U24112 (N_24112,N_23540,N_23674);
nand U24113 (N_24113,N_23803,N_23754);
and U24114 (N_24114,N_23852,N_23668);
and U24115 (N_24115,N_23931,N_23763);
nand U24116 (N_24116,N_23550,N_23869);
nand U24117 (N_24117,N_23837,N_23582);
or U24118 (N_24118,N_23654,N_23698);
nor U24119 (N_24119,N_23505,N_23812);
or U24120 (N_24120,N_23672,N_23525);
or U24121 (N_24121,N_23551,N_23542);
and U24122 (N_24122,N_23573,N_23899);
or U24123 (N_24123,N_23675,N_23715);
nand U24124 (N_24124,N_23978,N_23679);
and U24125 (N_24125,N_23595,N_23589);
nand U24126 (N_24126,N_23749,N_23945);
or U24127 (N_24127,N_23814,N_23828);
or U24128 (N_24128,N_23510,N_23643);
nor U24129 (N_24129,N_23766,N_23528);
or U24130 (N_24130,N_23559,N_23913);
xnor U24131 (N_24131,N_23695,N_23934);
nor U24132 (N_24132,N_23784,N_23970);
or U24133 (N_24133,N_23667,N_23771);
nor U24134 (N_24134,N_23787,N_23552);
nand U24135 (N_24135,N_23966,N_23957);
nand U24136 (N_24136,N_23958,N_23570);
or U24137 (N_24137,N_23517,N_23770);
nand U24138 (N_24138,N_23950,N_23802);
nor U24139 (N_24139,N_23804,N_23690);
xor U24140 (N_24140,N_23940,N_23977);
or U24141 (N_24141,N_23629,N_23555);
nor U24142 (N_24142,N_23561,N_23947);
and U24143 (N_24143,N_23533,N_23729);
nor U24144 (N_24144,N_23764,N_23815);
xor U24145 (N_24145,N_23919,N_23591);
and U24146 (N_24146,N_23976,N_23773);
nor U24147 (N_24147,N_23982,N_23929);
nor U24148 (N_24148,N_23598,N_23939);
or U24149 (N_24149,N_23623,N_23647);
xnor U24150 (N_24150,N_23986,N_23576);
nor U24151 (N_24151,N_23584,N_23969);
or U24152 (N_24152,N_23792,N_23549);
and U24153 (N_24153,N_23951,N_23659);
nand U24154 (N_24154,N_23850,N_23612);
nor U24155 (N_24155,N_23747,N_23820);
or U24156 (N_24156,N_23912,N_23862);
xor U24157 (N_24157,N_23948,N_23646);
nand U24158 (N_24158,N_23718,N_23581);
or U24159 (N_24159,N_23854,N_23988);
or U24160 (N_24160,N_23605,N_23884);
or U24161 (N_24161,N_23606,N_23624);
xnor U24162 (N_24162,N_23650,N_23686);
nand U24163 (N_24163,N_23554,N_23759);
xor U24164 (N_24164,N_23619,N_23661);
xor U24165 (N_24165,N_23531,N_23817);
xnor U24166 (N_24166,N_23656,N_23861);
or U24167 (N_24167,N_23775,N_23909);
nor U24168 (N_24168,N_23853,N_23707);
nand U24169 (N_24169,N_23682,N_23956);
or U24170 (N_24170,N_23719,N_23516);
nor U24171 (N_24171,N_23778,N_23941);
or U24172 (N_24172,N_23723,N_23530);
and U24173 (N_24173,N_23508,N_23588);
nand U24174 (N_24174,N_23896,N_23857);
xnor U24175 (N_24175,N_23953,N_23512);
nor U24176 (N_24176,N_23830,N_23534);
and U24177 (N_24177,N_23999,N_23745);
nand U24178 (N_24178,N_23577,N_23865);
nand U24179 (N_24179,N_23518,N_23702);
or U24180 (N_24180,N_23616,N_23755);
or U24181 (N_24181,N_23876,N_23897);
xnor U24182 (N_24182,N_23519,N_23893);
nor U24183 (N_24183,N_23705,N_23962);
nor U24184 (N_24184,N_23655,N_23906);
and U24185 (N_24185,N_23676,N_23887);
and U24186 (N_24186,N_23590,N_23627);
xnor U24187 (N_24187,N_23779,N_23653);
nand U24188 (N_24188,N_23526,N_23979);
xor U24189 (N_24189,N_23786,N_23714);
nand U24190 (N_24190,N_23553,N_23780);
xnor U24191 (N_24191,N_23725,N_23998);
nor U24192 (N_24192,N_23696,N_23795);
xor U24193 (N_24193,N_23665,N_23838);
or U24194 (N_24194,N_23768,N_23993);
nor U24195 (N_24195,N_23713,N_23515);
and U24196 (N_24196,N_23877,N_23943);
and U24197 (N_24197,N_23710,N_23911);
xor U24198 (N_24198,N_23571,N_23546);
nand U24199 (N_24199,N_23532,N_23604);
or U24200 (N_24200,N_23794,N_23892);
and U24201 (N_24201,N_23611,N_23937);
nand U24202 (N_24202,N_23808,N_23657);
nor U24203 (N_24203,N_23756,N_23753);
or U24204 (N_24204,N_23805,N_23959);
nand U24205 (N_24205,N_23800,N_23885);
xnor U24206 (N_24206,N_23593,N_23799);
nor U24207 (N_24207,N_23693,N_23833);
and U24208 (N_24208,N_23535,N_23879);
xor U24209 (N_24209,N_23569,N_23524);
xnor U24210 (N_24210,N_23827,N_23963);
and U24211 (N_24211,N_23575,N_23886);
nor U24212 (N_24212,N_23903,N_23790);
or U24213 (N_24213,N_23640,N_23594);
nor U24214 (N_24214,N_23740,N_23563);
and U24215 (N_24215,N_23967,N_23772);
or U24216 (N_24216,N_23936,N_23798);
nand U24217 (N_24217,N_23610,N_23574);
and U24218 (N_24218,N_23983,N_23762);
nor U24219 (N_24219,N_23748,N_23694);
and U24220 (N_24220,N_23846,N_23806);
nand U24221 (N_24221,N_23614,N_23926);
nand U24222 (N_24222,N_23849,N_23733);
nor U24223 (N_24223,N_23642,N_23987);
xor U24224 (N_24224,N_23706,N_23663);
and U24225 (N_24225,N_23529,N_23649);
xor U24226 (N_24226,N_23678,N_23597);
xnor U24227 (N_24227,N_23539,N_23677);
nand U24228 (N_24228,N_23961,N_23955);
and U24229 (N_24229,N_23543,N_23727);
and U24230 (N_24230,N_23746,N_23895);
or U24231 (N_24231,N_23989,N_23839);
nor U24232 (N_24232,N_23634,N_23832);
or U24233 (N_24233,N_23620,N_23782);
xor U24234 (N_24234,N_23648,N_23996);
or U24235 (N_24235,N_23870,N_23785);
nor U24236 (N_24236,N_23816,N_23600);
xor U24237 (N_24237,N_23743,N_23822);
and U24238 (N_24238,N_23818,N_23638);
or U24239 (N_24239,N_23810,N_23520);
nor U24240 (N_24240,N_23781,N_23560);
xor U24241 (N_24241,N_23875,N_23874);
nand U24242 (N_24242,N_23769,N_23692);
nor U24243 (N_24243,N_23697,N_23662);
nand U24244 (N_24244,N_23797,N_23922);
xor U24245 (N_24245,N_23992,N_23731);
or U24246 (N_24246,N_23734,N_23995);
and U24247 (N_24247,N_23558,N_23788);
xor U24248 (N_24248,N_23735,N_23709);
and U24249 (N_24249,N_23641,N_23915);
nor U24250 (N_24250,N_23816,N_23880);
nor U24251 (N_24251,N_23931,N_23981);
xnor U24252 (N_24252,N_23525,N_23934);
xnor U24253 (N_24253,N_23684,N_23767);
or U24254 (N_24254,N_23922,N_23636);
nand U24255 (N_24255,N_23794,N_23965);
nor U24256 (N_24256,N_23964,N_23639);
and U24257 (N_24257,N_23809,N_23852);
xor U24258 (N_24258,N_23896,N_23575);
or U24259 (N_24259,N_23801,N_23771);
nand U24260 (N_24260,N_23823,N_23736);
and U24261 (N_24261,N_23736,N_23733);
or U24262 (N_24262,N_23890,N_23991);
nand U24263 (N_24263,N_23653,N_23954);
or U24264 (N_24264,N_23582,N_23980);
or U24265 (N_24265,N_23774,N_23815);
nand U24266 (N_24266,N_23897,N_23927);
and U24267 (N_24267,N_23608,N_23792);
nor U24268 (N_24268,N_23884,N_23931);
xor U24269 (N_24269,N_23750,N_23605);
or U24270 (N_24270,N_23794,N_23562);
or U24271 (N_24271,N_23637,N_23669);
xnor U24272 (N_24272,N_23775,N_23663);
xnor U24273 (N_24273,N_23769,N_23651);
xor U24274 (N_24274,N_23972,N_23686);
nand U24275 (N_24275,N_23807,N_23716);
and U24276 (N_24276,N_23819,N_23789);
nor U24277 (N_24277,N_23942,N_23962);
nand U24278 (N_24278,N_23908,N_23552);
nor U24279 (N_24279,N_23973,N_23916);
nor U24280 (N_24280,N_23763,N_23942);
nand U24281 (N_24281,N_23743,N_23685);
xnor U24282 (N_24282,N_23978,N_23576);
nand U24283 (N_24283,N_23803,N_23700);
or U24284 (N_24284,N_23611,N_23799);
or U24285 (N_24285,N_23548,N_23755);
nand U24286 (N_24286,N_23949,N_23576);
and U24287 (N_24287,N_23980,N_23774);
nor U24288 (N_24288,N_23948,N_23624);
nand U24289 (N_24289,N_23648,N_23817);
or U24290 (N_24290,N_23934,N_23993);
and U24291 (N_24291,N_23934,N_23739);
or U24292 (N_24292,N_23991,N_23904);
nor U24293 (N_24293,N_23609,N_23613);
or U24294 (N_24294,N_23620,N_23773);
and U24295 (N_24295,N_23953,N_23668);
and U24296 (N_24296,N_23749,N_23695);
nor U24297 (N_24297,N_23742,N_23612);
xnor U24298 (N_24298,N_23740,N_23921);
nor U24299 (N_24299,N_23640,N_23917);
or U24300 (N_24300,N_23602,N_23562);
or U24301 (N_24301,N_23590,N_23669);
or U24302 (N_24302,N_23972,N_23744);
or U24303 (N_24303,N_23895,N_23818);
nand U24304 (N_24304,N_23906,N_23651);
and U24305 (N_24305,N_23948,N_23923);
nand U24306 (N_24306,N_23818,N_23752);
xor U24307 (N_24307,N_23747,N_23936);
or U24308 (N_24308,N_23526,N_23788);
or U24309 (N_24309,N_23871,N_23629);
xnor U24310 (N_24310,N_23547,N_23933);
xnor U24311 (N_24311,N_23553,N_23900);
nor U24312 (N_24312,N_23617,N_23506);
nor U24313 (N_24313,N_23546,N_23694);
nand U24314 (N_24314,N_23952,N_23994);
nor U24315 (N_24315,N_23617,N_23934);
nand U24316 (N_24316,N_23770,N_23977);
nand U24317 (N_24317,N_23678,N_23955);
xnor U24318 (N_24318,N_23934,N_23598);
or U24319 (N_24319,N_23617,N_23533);
and U24320 (N_24320,N_23511,N_23924);
nand U24321 (N_24321,N_23924,N_23505);
and U24322 (N_24322,N_23865,N_23591);
nor U24323 (N_24323,N_23646,N_23611);
nand U24324 (N_24324,N_23986,N_23929);
and U24325 (N_24325,N_23663,N_23795);
xor U24326 (N_24326,N_23895,N_23991);
nand U24327 (N_24327,N_23762,N_23879);
and U24328 (N_24328,N_23599,N_23551);
xor U24329 (N_24329,N_23506,N_23820);
xor U24330 (N_24330,N_23868,N_23935);
nand U24331 (N_24331,N_23903,N_23555);
or U24332 (N_24332,N_23912,N_23995);
or U24333 (N_24333,N_23607,N_23715);
and U24334 (N_24334,N_23976,N_23748);
or U24335 (N_24335,N_23558,N_23985);
and U24336 (N_24336,N_23878,N_23695);
and U24337 (N_24337,N_23832,N_23960);
xor U24338 (N_24338,N_23515,N_23512);
and U24339 (N_24339,N_23901,N_23567);
or U24340 (N_24340,N_23819,N_23510);
xnor U24341 (N_24341,N_23977,N_23829);
nand U24342 (N_24342,N_23629,N_23561);
nor U24343 (N_24343,N_23680,N_23548);
nor U24344 (N_24344,N_23520,N_23787);
nand U24345 (N_24345,N_23538,N_23944);
or U24346 (N_24346,N_23844,N_23920);
nand U24347 (N_24347,N_23682,N_23647);
or U24348 (N_24348,N_23894,N_23571);
or U24349 (N_24349,N_23846,N_23988);
and U24350 (N_24350,N_23687,N_23637);
and U24351 (N_24351,N_23627,N_23913);
or U24352 (N_24352,N_23619,N_23800);
nor U24353 (N_24353,N_23723,N_23711);
or U24354 (N_24354,N_23794,N_23815);
and U24355 (N_24355,N_23824,N_23671);
nor U24356 (N_24356,N_23744,N_23888);
nor U24357 (N_24357,N_23618,N_23726);
or U24358 (N_24358,N_23849,N_23760);
or U24359 (N_24359,N_23536,N_23604);
nor U24360 (N_24360,N_23650,N_23586);
xnor U24361 (N_24361,N_23942,N_23869);
xor U24362 (N_24362,N_23836,N_23945);
nand U24363 (N_24363,N_23761,N_23980);
nor U24364 (N_24364,N_23870,N_23830);
xor U24365 (N_24365,N_23832,N_23985);
and U24366 (N_24366,N_23804,N_23863);
xnor U24367 (N_24367,N_23920,N_23675);
and U24368 (N_24368,N_23741,N_23660);
nand U24369 (N_24369,N_23565,N_23507);
xnor U24370 (N_24370,N_23915,N_23919);
or U24371 (N_24371,N_23960,N_23769);
nor U24372 (N_24372,N_23531,N_23814);
nor U24373 (N_24373,N_23975,N_23995);
and U24374 (N_24374,N_23868,N_23819);
xnor U24375 (N_24375,N_23808,N_23850);
xnor U24376 (N_24376,N_23777,N_23838);
nor U24377 (N_24377,N_23509,N_23693);
nor U24378 (N_24378,N_23581,N_23651);
xnor U24379 (N_24379,N_23776,N_23570);
nand U24380 (N_24380,N_23833,N_23658);
nor U24381 (N_24381,N_23779,N_23862);
nor U24382 (N_24382,N_23853,N_23890);
nor U24383 (N_24383,N_23608,N_23645);
or U24384 (N_24384,N_23956,N_23882);
or U24385 (N_24385,N_23538,N_23827);
and U24386 (N_24386,N_23652,N_23653);
nand U24387 (N_24387,N_23826,N_23854);
nor U24388 (N_24388,N_23896,N_23957);
or U24389 (N_24389,N_23621,N_23608);
nand U24390 (N_24390,N_23956,N_23830);
nand U24391 (N_24391,N_23688,N_23518);
nor U24392 (N_24392,N_23904,N_23756);
xor U24393 (N_24393,N_23886,N_23908);
nor U24394 (N_24394,N_23557,N_23626);
xor U24395 (N_24395,N_23689,N_23553);
or U24396 (N_24396,N_23699,N_23768);
nand U24397 (N_24397,N_23982,N_23799);
or U24398 (N_24398,N_23942,N_23769);
nand U24399 (N_24399,N_23848,N_23928);
nor U24400 (N_24400,N_23722,N_23943);
or U24401 (N_24401,N_23553,N_23802);
nand U24402 (N_24402,N_23731,N_23691);
or U24403 (N_24403,N_23988,N_23990);
and U24404 (N_24404,N_23859,N_23671);
or U24405 (N_24405,N_23760,N_23665);
nor U24406 (N_24406,N_23837,N_23664);
nand U24407 (N_24407,N_23545,N_23531);
nor U24408 (N_24408,N_23643,N_23747);
or U24409 (N_24409,N_23540,N_23972);
and U24410 (N_24410,N_23501,N_23876);
xnor U24411 (N_24411,N_23763,N_23715);
or U24412 (N_24412,N_23737,N_23979);
nand U24413 (N_24413,N_23708,N_23542);
nand U24414 (N_24414,N_23770,N_23998);
and U24415 (N_24415,N_23902,N_23542);
nand U24416 (N_24416,N_23605,N_23668);
nand U24417 (N_24417,N_23655,N_23804);
nand U24418 (N_24418,N_23958,N_23603);
or U24419 (N_24419,N_23622,N_23763);
nor U24420 (N_24420,N_23948,N_23724);
nand U24421 (N_24421,N_23528,N_23735);
nor U24422 (N_24422,N_23734,N_23708);
xor U24423 (N_24423,N_23607,N_23903);
nor U24424 (N_24424,N_23957,N_23774);
nor U24425 (N_24425,N_23964,N_23723);
and U24426 (N_24426,N_23720,N_23845);
nor U24427 (N_24427,N_23504,N_23975);
or U24428 (N_24428,N_23526,N_23878);
or U24429 (N_24429,N_23947,N_23904);
nor U24430 (N_24430,N_23908,N_23672);
and U24431 (N_24431,N_23589,N_23620);
nand U24432 (N_24432,N_23935,N_23589);
xnor U24433 (N_24433,N_23895,N_23579);
nor U24434 (N_24434,N_23941,N_23594);
nor U24435 (N_24435,N_23523,N_23654);
nand U24436 (N_24436,N_23971,N_23804);
nor U24437 (N_24437,N_23524,N_23681);
nor U24438 (N_24438,N_23502,N_23595);
xnor U24439 (N_24439,N_23595,N_23650);
nand U24440 (N_24440,N_23762,N_23900);
xor U24441 (N_24441,N_23518,N_23608);
nor U24442 (N_24442,N_23916,N_23908);
xnor U24443 (N_24443,N_23533,N_23674);
xor U24444 (N_24444,N_23880,N_23976);
nand U24445 (N_24445,N_23550,N_23700);
or U24446 (N_24446,N_23545,N_23968);
nor U24447 (N_24447,N_23714,N_23979);
xor U24448 (N_24448,N_23764,N_23716);
xor U24449 (N_24449,N_23658,N_23983);
nand U24450 (N_24450,N_23960,N_23915);
or U24451 (N_24451,N_23696,N_23963);
nor U24452 (N_24452,N_23974,N_23897);
nand U24453 (N_24453,N_23520,N_23963);
or U24454 (N_24454,N_23966,N_23891);
xor U24455 (N_24455,N_23511,N_23530);
xnor U24456 (N_24456,N_23990,N_23931);
and U24457 (N_24457,N_23875,N_23664);
nor U24458 (N_24458,N_23920,N_23781);
nor U24459 (N_24459,N_23575,N_23639);
nor U24460 (N_24460,N_23767,N_23596);
or U24461 (N_24461,N_23868,N_23729);
nand U24462 (N_24462,N_23918,N_23814);
nand U24463 (N_24463,N_23530,N_23913);
or U24464 (N_24464,N_23667,N_23613);
nand U24465 (N_24465,N_23847,N_23788);
or U24466 (N_24466,N_23649,N_23581);
nand U24467 (N_24467,N_23814,N_23651);
xor U24468 (N_24468,N_23807,N_23583);
nand U24469 (N_24469,N_23709,N_23685);
and U24470 (N_24470,N_23697,N_23909);
and U24471 (N_24471,N_23526,N_23633);
xnor U24472 (N_24472,N_23895,N_23704);
nand U24473 (N_24473,N_23972,N_23958);
nand U24474 (N_24474,N_23744,N_23675);
xnor U24475 (N_24475,N_23514,N_23576);
and U24476 (N_24476,N_23518,N_23532);
xor U24477 (N_24477,N_23776,N_23656);
or U24478 (N_24478,N_23730,N_23712);
and U24479 (N_24479,N_23961,N_23901);
nor U24480 (N_24480,N_23688,N_23554);
xor U24481 (N_24481,N_23880,N_23885);
nor U24482 (N_24482,N_23977,N_23886);
or U24483 (N_24483,N_23723,N_23807);
nand U24484 (N_24484,N_23956,N_23668);
nand U24485 (N_24485,N_23721,N_23826);
nand U24486 (N_24486,N_23655,N_23778);
or U24487 (N_24487,N_23600,N_23582);
nand U24488 (N_24488,N_23984,N_23783);
and U24489 (N_24489,N_23702,N_23692);
or U24490 (N_24490,N_23771,N_23625);
nor U24491 (N_24491,N_23512,N_23636);
and U24492 (N_24492,N_23555,N_23615);
nand U24493 (N_24493,N_23724,N_23660);
xnor U24494 (N_24494,N_23831,N_23553);
and U24495 (N_24495,N_23615,N_23698);
nor U24496 (N_24496,N_23887,N_23729);
nor U24497 (N_24497,N_23745,N_23903);
or U24498 (N_24498,N_23670,N_23741);
nor U24499 (N_24499,N_23697,N_23991);
nor U24500 (N_24500,N_24467,N_24307);
and U24501 (N_24501,N_24324,N_24426);
nor U24502 (N_24502,N_24270,N_24365);
nor U24503 (N_24503,N_24078,N_24011);
nand U24504 (N_24504,N_24394,N_24013);
nand U24505 (N_24505,N_24395,N_24456);
nor U24506 (N_24506,N_24271,N_24001);
nand U24507 (N_24507,N_24290,N_24184);
xnor U24508 (N_24508,N_24172,N_24058);
and U24509 (N_24509,N_24299,N_24083);
and U24510 (N_24510,N_24152,N_24225);
and U24511 (N_24511,N_24375,N_24416);
and U24512 (N_24512,N_24059,N_24351);
nand U24513 (N_24513,N_24476,N_24391);
nand U24514 (N_24514,N_24255,N_24355);
nor U24515 (N_24515,N_24433,N_24200);
and U24516 (N_24516,N_24010,N_24085);
nor U24517 (N_24517,N_24114,N_24260);
xnor U24518 (N_24518,N_24331,N_24428);
nor U24519 (N_24519,N_24376,N_24396);
and U24520 (N_24520,N_24107,N_24095);
xnor U24521 (N_24521,N_24047,N_24491);
nand U24522 (N_24522,N_24398,N_24486);
nand U24523 (N_24523,N_24070,N_24026);
and U24524 (N_24524,N_24481,N_24357);
xor U24525 (N_24525,N_24474,N_24303);
and U24526 (N_24526,N_24234,N_24262);
nand U24527 (N_24527,N_24119,N_24419);
xnor U24528 (N_24528,N_24090,N_24320);
nand U24529 (N_24529,N_24215,N_24148);
or U24530 (N_24530,N_24492,N_24199);
nand U24531 (N_24531,N_24111,N_24342);
xnor U24532 (N_24532,N_24166,N_24319);
nor U24533 (N_24533,N_24084,N_24359);
xnor U24534 (N_24534,N_24462,N_24191);
or U24535 (N_24535,N_24240,N_24141);
nor U24536 (N_24536,N_24005,N_24473);
nor U24537 (N_24537,N_24366,N_24062);
and U24538 (N_24538,N_24449,N_24310);
or U24539 (N_24539,N_24427,N_24160);
nor U24540 (N_24540,N_24325,N_24499);
xnor U24541 (N_24541,N_24381,N_24096);
and U24542 (N_24542,N_24444,N_24135);
nand U24543 (N_24543,N_24393,N_24293);
or U24544 (N_24544,N_24168,N_24201);
xor U24545 (N_24545,N_24109,N_24007);
and U24546 (N_24546,N_24175,N_24251);
nand U24547 (N_24547,N_24280,N_24340);
and U24548 (N_24548,N_24347,N_24269);
and U24549 (N_24549,N_24131,N_24284);
and U24550 (N_24550,N_24003,N_24134);
or U24551 (N_24551,N_24079,N_24432);
and U24552 (N_24552,N_24489,N_24086);
nor U24553 (N_24553,N_24438,N_24032);
or U24554 (N_24554,N_24401,N_24214);
nand U24555 (N_24555,N_24480,N_24328);
nand U24556 (N_24556,N_24371,N_24350);
xor U24557 (N_24557,N_24036,N_24336);
nor U24558 (N_24558,N_24445,N_24226);
xor U24559 (N_24559,N_24322,N_24118);
and U24560 (N_24560,N_24144,N_24126);
xor U24561 (N_24561,N_24165,N_24469);
xnor U24562 (N_24562,N_24498,N_24495);
nand U24563 (N_24563,N_24222,N_24281);
or U24564 (N_24564,N_24441,N_24430);
nand U24565 (N_24565,N_24389,N_24023);
xnor U24566 (N_24566,N_24117,N_24051);
xnor U24567 (N_24567,N_24143,N_24087);
xnor U24568 (N_24568,N_24493,N_24202);
xnor U24569 (N_24569,N_24294,N_24415);
xnor U24570 (N_24570,N_24162,N_24248);
or U24571 (N_24571,N_24470,N_24037);
nand U24572 (N_24572,N_24334,N_24203);
and U24573 (N_24573,N_24156,N_24309);
nor U24574 (N_24574,N_24247,N_24439);
nor U24575 (N_24575,N_24257,N_24400);
or U24576 (N_24576,N_24127,N_24031);
or U24577 (N_24577,N_24386,N_24478);
or U24578 (N_24578,N_24313,N_24335);
and U24579 (N_24579,N_24088,N_24291);
nand U24580 (N_24580,N_24420,N_24329);
xnor U24581 (N_24581,N_24108,N_24170);
nand U24582 (N_24582,N_24435,N_24140);
and U24583 (N_24583,N_24345,N_24139);
and U24584 (N_24584,N_24460,N_24112);
and U24585 (N_24585,N_24124,N_24224);
and U24586 (N_24586,N_24150,N_24380);
or U24587 (N_24587,N_24128,N_24061);
and U24588 (N_24588,N_24276,N_24060);
nor U24589 (N_24589,N_24264,N_24154);
and U24590 (N_24590,N_24110,N_24198);
xnor U24591 (N_24591,N_24102,N_24443);
xor U24592 (N_24592,N_24197,N_24372);
nand U24593 (N_24593,N_24423,N_24158);
and U24594 (N_24594,N_24490,N_24362);
or U24595 (N_24595,N_24116,N_24465);
nand U24596 (N_24596,N_24179,N_24341);
nor U24597 (N_24597,N_24487,N_24193);
and U24598 (N_24598,N_24073,N_24295);
nand U24599 (N_24599,N_24403,N_24074);
or U24600 (N_24600,N_24475,N_24223);
or U24601 (N_24601,N_24397,N_24015);
and U24602 (N_24602,N_24321,N_24218);
nand U24603 (N_24603,N_24055,N_24122);
or U24604 (N_24604,N_24315,N_24043);
or U24605 (N_24605,N_24318,N_24067);
nor U24606 (N_24606,N_24369,N_24268);
and U24607 (N_24607,N_24016,N_24301);
nor U24608 (N_24608,N_24233,N_24004);
and U24609 (N_24609,N_24330,N_24408);
or U24610 (N_24610,N_24113,N_24298);
xor U24611 (N_24611,N_24132,N_24275);
nand U24612 (N_24612,N_24206,N_24285);
xnor U24613 (N_24613,N_24484,N_24354);
nand U24614 (N_24614,N_24077,N_24064);
nor U24615 (N_24615,N_24093,N_24250);
xnor U24616 (N_24616,N_24219,N_24000);
xor U24617 (N_24617,N_24136,N_24384);
nor U24618 (N_24618,N_24072,N_24425);
nor U24619 (N_24619,N_24254,N_24065);
and U24620 (N_24620,N_24305,N_24429);
or U24621 (N_24621,N_24306,N_24497);
or U24622 (N_24622,N_24056,N_24496);
xor U24623 (N_24623,N_24069,N_24451);
xor U24624 (N_24624,N_24022,N_24244);
xnor U24625 (N_24625,N_24287,N_24187);
nand U24626 (N_24626,N_24195,N_24379);
nand U24627 (N_24627,N_24446,N_24133);
nand U24628 (N_24628,N_24289,N_24304);
nand U24629 (N_24629,N_24123,N_24263);
xor U24630 (N_24630,N_24146,N_24453);
nor U24631 (N_24631,N_24209,N_24349);
xor U24632 (N_24632,N_24405,N_24387);
and U24633 (N_24633,N_24259,N_24171);
nand U24634 (N_24634,N_24044,N_24228);
nand U24635 (N_24635,N_24180,N_24278);
nand U24636 (N_24636,N_24190,N_24245);
or U24637 (N_24637,N_24314,N_24272);
nor U24638 (N_24638,N_24482,N_24008);
or U24639 (N_24639,N_24185,N_24327);
nand U24640 (N_24640,N_24368,N_24027);
or U24641 (N_24641,N_24018,N_24174);
or U24642 (N_24642,N_24358,N_24188);
nand U24643 (N_24643,N_24409,N_24207);
nand U24644 (N_24644,N_24390,N_24485);
xnor U24645 (N_24645,N_24436,N_24377);
nand U24646 (N_24646,N_24300,N_24103);
xor U24647 (N_24647,N_24242,N_24297);
nand U24648 (N_24648,N_24232,N_24494);
xor U24649 (N_24649,N_24054,N_24477);
and U24650 (N_24650,N_24045,N_24002);
nand U24651 (N_24651,N_24081,N_24472);
xor U24652 (N_24652,N_24479,N_24343);
and U24653 (N_24653,N_24283,N_24367);
xnor U24654 (N_24654,N_24217,N_24080);
and U24655 (N_24655,N_24265,N_24361);
nor U24656 (N_24656,N_24249,N_24266);
xor U24657 (N_24657,N_24411,N_24053);
xnor U24658 (N_24658,N_24035,N_24099);
nand U24659 (N_24659,N_24137,N_24040);
xor U24660 (N_24660,N_24373,N_24286);
and U24661 (N_24661,N_24458,N_24292);
nor U24662 (N_24662,N_24344,N_24332);
and U24663 (N_24663,N_24147,N_24189);
xor U24664 (N_24664,N_24014,N_24075);
nand U24665 (N_24665,N_24076,N_24104);
or U24666 (N_24666,N_24048,N_24006);
or U24667 (N_24667,N_24155,N_24145);
and U24668 (N_24668,N_24421,N_24089);
and U24669 (N_24669,N_24049,N_24177);
nand U24670 (N_24670,N_24461,N_24352);
or U24671 (N_24671,N_24282,N_24100);
nor U24672 (N_24672,N_24063,N_24196);
and U24673 (N_24673,N_24442,N_24235);
nand U24674 (N_24674,N_24360,N_24316);
xor U24675 (N_24675,N_24192,N_24459);
and U24676 (N_24676,N_24399,N_24012);
nand U24677 (N_24677,N_24169,N_24106);
nor U24678 (N_24678,N_24452,N_24238);
and U24679 (N_24679,N_24082,N_24221);
and U24680 (N_24680,N_24237,N_24097);
nor U24681 (N_24681,N_24382,N_24378);
and U24682 (N_24682,N_24092,N_24216);
and U24683 (N_24683,N_24211,N_24370);
or U24684 (N_24684,N_24213,N_24431);
or U24685 (N_24685,N_24440,N_24273);
nand U24686 (N_24686,N_24464,N_24437);
nor U24687 (N_24687,N_24447,N_24205);
and U24688 (N_24688,N_24455,N_24178);
or U24689 (N_24689,N_24153,N_24253);
and U24690 (N_24690,N_24230,N_24346);
xnor U24691 (N_24691,N_24034,N_24138);
or U24692 (N_24692,N_24279,N_24021);
or U24693 (N_24693,N_24167,N_24115);
or U24694 (N_24694,N_24227,N_24164);
nand U24695 (N_24695,N_24392,N_24039);
or U24696 (N_24696,N_24050,N_24186);
or U24697 (N_24697,N_24448,N_24017);
and U24698 (N_24698,N_24038,N_24413);
and U24699 (N_24699,N_24068,N_24157);
nand U24700 (N_24700,N_24418,N_24353);
and U24701 (N_24701,N_24161,N_24091);
or U24702 (N_24702,N_24434,N_24338);
nand U24703 (N_24703,N_24277,N_24312);
nand U24704 (N_24704,N_24057,N_24274);
xnor U24705 (N_24705,N_24422,N_24406);
nand U24706 (N_24706,N_24258,N_24457);
and U24707 (N_24707,N_24066,N_24046);
nand U24708 (N_24708,N_24468,N_24163);
and U24709 (N_24709,N_24414,N_24348);
nor U24710 (N_24710,N_24019,N_24302);
nand U24711 (N_24711,N_24388,N_24383);
or U24712 (N_24712,N_24364,N_24121);
xor U24713 (N_24713,N_24308,N_24471);
xor U24714 (N_24714,N_24488,N_24105);
nand U24715 (N_24715,N_24220,N_24009);
nand U24716 (N_24716,N_24071,N_24424);
nand U24717 (N_24717,N_24024,N_24101);
or U24718 (N_24718,N_24317,N_24407);
or U24719 (N_24719,N_24208,N_24098);
and U24720 (N_24720,N_24323,N_24120);
and U24721 (N_24721,N_24033,N_24311);
nor U24722 (N_24722,N_24410,N_24151);
nand U24723 (N_24723,N_24129,N_24463);
xnor U24724 (N_24724,N_24212,N_24149);
nand U24725 (N_24725,N_24030,N_24229);
nor U24726 (N_24726,N_24041,N_24337);
xor U24727 (N_24727,N_24020,N_24246);
xor U24728 (N_24728,N_24385,N_24450);
nor U24729 (N_24729,N_24194,N_24239);
nor U24730 (N_24730,N_24231,N_24130);
and U24731 (N_24731,N_24159,N_24094);
nor U24732 (N_24732,N_24028,N_24173);
or U24733 (N_24733,N_24029,N_24256);
nand U24734 (N_24734,N_24042,N_24204);
nand U24735 (N_24735,N_24267,N_24288);
and U24736 (N_24736,N_24142,N_24182);
and U24737 (N_24737,N_24402,N_24181);
nand U24738 (N_24738,N_24356,N_24404);
nand U24739 (N_24739,N_24252,N_24236);
xnor U24740 (N_24740,N_24210,N_24176);
and U24741 (N_24741,N_24454,N_24363);
xor U24742 (N_24742,N_24483,N_24261);
or U24743 (N_24743,N_24243,N_24125);
xnor U24744 (N_24744,N_24025,N_24339);
or U24745 (N_24745,N_24296,N_24374);
and U24746 (N_24746,N_24412,N_24417);
or U24747 (N_24747,N_24183,N_24333);
and U24748 (N_24748,N_24052,N_24466);
and U24749 (N_24749,N_24241,N_24326);
or U24750 (N_24750,N_24018,N_24497);
or U24751 (N_24751,N_24260,N_24181);
or U24752 (N_24752,N_24206,N_24221);
or U24753 (N_24753,N_24352,N_24484);
nor U24754 (N_24754,N_24399,N_24060);
and U24755 (N_24755,N_24052,N_24276);
or U24756 (N_24756,N_24257,N_24304);
nand U24757 (N_24757,N_24325,N_24244);
or U24758 (N_24758,N_24032,N_24157);
or U24759 (N_24759,N_24238,N_24270);
and U24760 (N_24760,N_24279,N_24146);
nand U24761 (N_24761,N_24488,N_24071);
nor U24762 (N_24762,N_24386,N_24437);
xor U24763 (N_24763,N_24386,N_24251);
and U24764 (N_24764,N_24184,N_24050);
xor U24765 (N_24765,N_24490,N_24131);
or U24766 (N_24766,N_24296,N_24419);
or U24767 (N_24767,N_24108,N_24232);
nand U24768 (N_24768,N_24388,N_24483);
nand U24769 (N_24769,N_24054,N_24134);
nor U24770 (N_24770,N_24430,N_24058);
and U24771 (N_24771,N_24381,N_24322);
nand U24772 (N_24772,N_24240,N_24493);
nor U24773 (N_24773,N_24386,N_24197);
and U24774 (N_24774,N_24128,N_24312);
nor U24775 (N_24775,N_24340,N_24411);
nand U24776 (N_24776,N_24397,N_24220);
nand U24777 (N_24777,N_24443,N_24451);
xnor U24778 (N_24778,N_24491,N_24281);
xnor U24779 (N_24779,N_24420,N_24390);
nand U24780 (N_24780,N_24053,N_24152);
nor U24781 (N_24781,N_24465,N_24217);
nor U24782 (N_24782,N_24116,N_24345);
nand U24783 (N_24783,N_24127,N_24402);
nor U24784 (N_24784,N_24311,N_24236);
and U24785 (N_24785,N_24458,N_24392);
nand U24786 (N_24786,N_24126,N_24422);
nor U24787 (N_24787,N_24212,N_24476);
nand U24788 (N_24788,N_24121,N_24459);
or U24789 (N_24789,N_24381,N_24373);
nor U24790 (N_24790,N_24288,N_24067);
nor U24791 (N_24791,N_24310,N_24038);
nor U24792 (N_24792,N_24235,N_24308);
nand U24793 (N_24793,N_24362,N_24233);
nor U24794 (N_24794,N_24154,N_24139);
and U24795 (N_24795,N_24318,N_24420);
nor U24796 (N_24796,N_24470,N_24338);
xnor U24797 (N_24797,N_24234,N_24288);
or U24798 (N_24798,N_24148,N_24257);
nand U24799 (N_24799,N_24199,N_24425);
and U24800 (N_24800,N_24389,N_24415);
nor U24801 (N_24801,N_24157,N_24198);
and U24802 (N_24802,N_24030,N_24102);
nor U24803 (N_24803,N_24413,N_24124);
xor U24804 (N_24804,N_24382,N_24186);
nor U24805 (N_24805,N_24493,N_24319);
or U24806 (N_24806,N_24339,N_24037);
or U24807 (N_24807,N_24462,N_24276);
and U24808 (N_24808,N_24488,N_24476);
nand U24809 (N_24809,N_24442,N_24348);
xnor U24810 (N_24810,N_24322,N_24264);
and U24811 (N_24811,N_24057,N_24379);
nor U24812 (N_24812,N_24292,N_24365);
nand U24813 (N_24813,N_24060,N_24428);
xnor U24814 (N_24814,N_24383,N_24282);
nand U24815 (N_24815,N_24176,N_24066);
and U24816 (N_24816,N_24218,N_24384);
nand U24817 (N_24817,N_24385,N_24499);
or U24818 (N_24818,N_24060,N_24042);
or U24819 (N_24819,N_24065,N_24235);
xor U24820 (N_24820,N_24241,N_24170);
nor U24821 (N_24821,N_24240,N_24225);
nor U24822 (N_24822,N_24487,N_24370);
and U24823 (N_24823,N_24428,N_24313);
nor U24824 (N_24824,N_24414,N_24488);
nor U24825 (N_24825,N_24041,N_24366);
nand U24826 (N_24826,N_24284,N_24438);
and U24827 (N_24827,N_24334,N_24361);
or U24828 (N_24828,N_24122,N_24384);
or U24829 (N_24829,N_24027,N_24418);
nor U24830 (N_24830,N_24305,N_24353);
or U24831 (N_24831,N_24220,N_24325);
and U24832 (N_24832,N_24091,N_24172);
or U24833 (N_24833,N_24476,N_24137);
and U24834 (N_24834,N_24047,N_24391);
or U24835 (N_24835,N_24485,N_24017);
or U24836 (N_24836,N_24179,N_24476);
xnor U24837 (N_24837,N_24219,N_24349);
nand U24838 (N_24838,N_24136,N_24445);
or U24839 (N_24839,N_24121,N_24061);
or U24840 (N_24840,N_24145,N_24237);
xor U24841 (N_24841,N_24403,N_24051);
nor U24842 (N_24842,N_24301,N_24401);
or U24843 (N_24843,N_24453,N_24084);
and U24844 (N_24844,N_24237,N_24154);
xnor U24845 (N_24845,N_24317,N_24212);
or U24846 (N_24846,N_24306,N_24327);
nor U24847 (N_24847,N_24219,N_24032);
and U24848 (N_24848,N_24439,N_24263);
and U24849 (N_24849,N_24292,N_24286);
nor U24850 (N_24850,N_24020,N_24017);
nand U24851 (N_24851,N_24497,N_24189);
nand U24852 (N_24852,N_24393,N_24094);
or U24853 (N_24853,N_24367,N_24126);
and U24854 (N_24854,N_24468,N_24383);
or U24855 (N_24855,N_24396,N_24189);
nor U24856 (N_24856,N_24059,N_24396);
or U24857 (N_24857,N_24473,N_24105);
and U24858 (N_24858,N_24035,N_24289);
or U24859 (N_24859,N_24283,N_24470);
nand U24860 (N_24860,N_24311,N_24255);
and U24861 (N_24861,N_24098,N_24045);
and U24862 (N_24862,N_24213,N_24285);
and U24863 (N_24863,N_24056,N_24480);
and U24864 (N_24864,N_24235,N_24381);
nor U24865 (N_24865,N_24439,N_24214);
and U24866 (N_24866,N_24244,N_24493);
or U24867 (N_24867,N_24415,N_24380);
and U24868 (N_24868,N_24355,N_24078);
nand U24869 (N_24869,N_24068,N_24447);
or U24870 (N_24870,N_24139,N_24093);
or U24871 (N_24871,N_24351,N_24427);
nand U24872 (N_24872,N_24308,N_24050);
and U24873 (N_24873,N_24327,N_24377);
and U24874 (N_24874,N_24207,N_24106);
nor U24875 (N_24875,N_24001,N_24387);
or U24876 (N_24876,N_24486,N_24459);
or U24877 (N_24877,N_24313,N_24215);
and U24878 (N_24878,N_24210,N_24250);
and U24879 (N_24879,N_24388,N_24195);
and U24880 (N_24880,N_24208,N_24166);
and U24881 (N_24881,N_24313,N_24223);
nor U24882 (N_24882,N_24178,N_24384);
and U24883 (N_24883,N_24450,N_24441);
nand U24884 (N_24884,N_24276,N_24246);
or U24885 (N_24885,N_24401,N_24038);
xnor U24886 (N_24886,N_24124,N_24498);
and U24887 (N_24887,N_24406,N_24181);
and U24888 (N_24888,N_24480,N_24104);
or U24889 (N_24889,N_24299,N_24119);
or U24890 (N_24890,N_24261,N_24014);
xor U24891 (N_24891,N_24129,N_24031);
nor U24892 (N_24892,N_24429,N_24200);
nor U24893 (N_24893,N_24349,N_24309);
xor U24894 (N_24894,N_24445,N_24287);
and U24895 (N_24895,N_24172,N_24158);
xor U24896 (N_24896,N_24032,N_24233);
or U24897 (N_24897,N_24388,N_24091);
nor U24898 (N_24898,N_24378,N_24355);
and U24899 (N_24899,N_24457,N_24241);
nand U24900 (N_24900,N_24469,N_24145);
nor U24901 (N_24901,N_24018,N_24485);
and U24902 (N_24902,N_24336,N_24097);
nand U24903 (N_24903,N_24245,N_24359);
or U24904 (N_24904,N_24238,N_24222);
nand U24905 (N_24905,N_24337,N_24491);
or U24906 (N_24906,N_24385,N_24315);
or U24907 (N_24907,N_24141,N_24198);
and U24908 (N_24908,N_24228,N_24071);
nor U24909 (N_24909,N_24402,N_24025);
nor U24910 (N_24910,N_24338,N_24144);
xor U24911 (N_24911,N_24469,N_24493);
nor U24912 (N_24912,N_24081,N_24285);
or U24913 (N_24913,N_24308,N_24179);
or U24914 (N_24914,N_24099,N_24236);
nor U24915 (N_24915,N_24423,N_24247);
nor U24916 (N_24916,N_24438,N_24396);
nor U24917 (N_24917,N_24045,N_24493);
or U24918 (N_24918,N_24287,N_24318);
and U24919 (N_24919,N_24285,N_24300);
xor U24920 (N_24920,N_24393,N_24270);
nor U24921 (N_24921,N_24302,N_24319);
and U24922 (N_24922,N_24185,N_24371);
xor U24923 (N_24923,N_24098,N_24369);
or U24924 (N_24924,N_24288,N_24292);
xor U24925 (N_24925,N_24136,N_24376);
nor U24926 (N_24926,N_24213,N_24295);
or U24927 (N_24927,N_24367,N_24481);
nor U24928 (N_24928,N_24114,N_24054);
or U24929 (N_24929,N_24308,N_24000);
or U24930 (N_24930,N_24166,N_24059);
xnor U24931 (N_24931,N_24297,N_24374);
and U24932 (N_24932,N_24317,N_24037);
and U24933 (N_24933,N_24240,N_24457);
or U24934 (N_24934,N_24127,N_24296);
and U24935 (N_24935,N_24323,N_24394);
nor U24936 (N_24936,N_24394,N_24301);
nor U24937 (N_24937,N_24396,N_24206);
nand U24938 (N_24938,N_24139,N_24297);
and U24939 (N_24939,N_24433,N_24462);
or U24940 (N_24940,N_24243,N_24081);
and U24941 (N_24941,N_24324,N_24264);
nand U24942 (N_24942,N_24336,N_24170);
nand U24943 (N_24943,N_24013,N_24399);
xnor U24944 (N_24944,N_24366,N_24114);
xor U24945 (N_24945,N_24316,N_24013);
nor U24946 (N_24946,N_24276,N_24217);
nand U24947 (N_24947,N_24379,N_24325);
and U24948 (N_24948,N_24470,N_24310);
or U24949 (N_24949,N_24236,N_24018);
or U24950 (N_24950,N_24079,N_24458);
nand U24951 (N_24951,N_24496,N_24094);
xnor U24952 (N_24952,N_24409,N_24382);
and U24953 (N_24953,N_24100,N_24426);
and U24954 (N_24954,N_24348,N_24498);
or U24955 (N_24955,N_24196,N_24392);
xnor U24956 (N_24956,N_24364,N_24386);
and U24957 (N_24957,N_24052,N_24272);
or U24958 (N_24958,N_24161,N_24014);
and U24959 (N_24959,N_24286,N_24427);
nand U24960 (N_24960,N_24414,N_24354);
and U24961 (N_24961,N_24106,N_24179);
nand U24962 (N_24962,N_24300,N_24496);
and U24963 (N_24963,N_24265,N_24151);
and U24964 (N_24964,N_24483,N_24235);
or U24965 (N_24965,N_24314,N_24277);
or U24966 (N_24966,N_24058,N_24317);
nor U24967 (N_24967,N_24269,N_24007);
nor U24968 (N_24968,N_24228,N_24317);
xnor U24969 (N_24969,N_24459,N_24420);
nor U24970 (N_24970,N_24419,N_24162);
or U24971 (N_24971,N_24430,N_24196);
or U24972 (N_24972,N_24237,N_24100);
nand U24973 (N_24973,N_24261,N_24242);
nand U24974 (N_24974,N_24239,N_24466);
and U24975 (N_24975,N_24247,N_24328);
and U24976 (N_24976,N_24324,N_24066);
nand U24977 (N_24977,N_24023,N_24322);
nand U24978 (N_24978,N_24454,N_24267);
nand U24979 (N_24979,N_24437,N_24254);
xor U24980 (N_24980,N_24236,N_24409);
and U24981 (N_24981,N_24255,N_24429);
xor U24982 (N_24982,N_24392,N_24053);
and U24983 (N_24983,N_24107,N_24227);
and U24984 (N_24984,N_24242,N_24332);
nand U24985 (N_24985,N_24424,N_24096);
or U24986 (N_24986,N_24053,N_24186);
nor U24987 (N_24987,N_24415,N_24405);
xnor U24988 (N_24988,N_24441,N_24411);
nor U24989 (N_24989,N_24457,N_24284);
nor U24990 (N_24990,N_24211,N_24471);
nand U24991 (N_24991,N_24241,N_24472);
and U24992 (N_24992,N_24344,N_24166);
or U24993 (N_24993,N_24458,N_24347);
nand U24994 (N_24994,N_24006,N_24342);
nor U24995 (N_24995,N_24135,N_24103);
or U24996 (N_24996,N_24263,N_24156);
nor U24997 (N_24997,N_24053,N_24266);
or U24998 (N_24998,N_24216,N_24429);
nor U24999 (N_24999,N_24156,N_24066);
nand U25000 (N_25000,N_24577,N_24701);
and U25001 (N_25001,N_24695,N_24608);
nand U25002 (N_25002,N_24958,N_24794);
nand U25003 (N_25003,N_24938,N_24592);
nand U25004 (N_25004,N_24635,N_24541);
or U25005 (N_25005,N_24530,N_24925);
and U25006 (N_25006,N_24671,N_24884);
nor U25007 (N_25007,N_24900,N_24786);
xnor U25008 (N_25008,N_24706,N_24791);
nand U25009 (N_25009,N_24994,N_24922);
and U25010 (N_25010,N_24961,N_24683);
or U25011 (N_25011,N_24979,N_24563);
xnor U25012 (N_25012,N_24949,N_24647);
nand U25013 (N_25013,N_24525,N_24948);
or U25014 (N_25014,N_24677,N_24595);
xor U25015 (N_25015,N_24660,N_24777);
nor U25016 (N_25016,N_24669,N_24590);
nand U25017 (N_25017,N_24687,N_24906);
or U25018 (N_25018,N_24727,N_24553);
and U25019 (N_25019,N_24916,N_24760);
and U25020 (N_25020,N_24616,N_24887);
and U25021 (N_25021,N_24516,N_24555);
xnor U25022 (N_25022,N_24567,N_24703);
nor U25023 (N_25023,N_24575,N_24837);
nor U25024 (N_25024,N_24691,N_24751);
xor U25025 (N_25025,N_24743,N_24593);
xor U25026 (N_25026,N_24766,N_24598);
or U25027 (N_25027,N_24601,N_24679);
xor U25028 (N_25028,N_24972,N_24645);
nor U25029 (N_25029,N_24545,N_24926);
and U25030 (N_25030,N_24845,N_24813);
or U25031 (N_25031,N_24672,N_24615);
nand U25032 (N_25032,N_24842,N_24789);
xor U25033 (N_25033,N_24862,N_24790);
nor U25034 (N_25034,N_24589,N_24977);
xnor U25035 (N_25035,N_24947,N_24664);
nor U25036 (N_25036,N_24769,N_24606);
xnor U25037 (N_25037,N_24620,N_24897);
nand U25038 (N_25038,N_24918,N_24557);
xor U25039 (N_25039,N_24890,N_24982);
nand U25040 (N_25040,N_24819,N_24778);
nor U25041 (N_25041,N_24855,N_24711);
or U25042 (N_25042,N_24886,N_24940);
nand U25043 (N_25043,N_24914,N_24973);
and U25044 (N_25044,N_24936,N_24632);
and U25045 (N_25045,N_24536,N_24854);
xor U25046 (N_25046,N_24623,N_24543);
or U25047 (N_25047,N_24966,N_24882);
xor U25048 (N_25048,N_24740,N_24867);
or U25049 (N_25049,N_24946,N_24821);
or U25050 (N_25050,N_24712,N_24825);
nand U25051 (N_25051,N_24708,N_24907);
and U25052 (N_25052,N_24588,N_24731);
xor U25053 (N_25053,N_24941,N_24534);
and U25054 (N_25054,N_24678,N_24722);
and U25055 (N_25055,N_24501,N_24990);
nor U25056 (N_25056,N_24749,N_24573);
and U25057 (N_25057,N_24866,N_24704);
or U25058 (N_25058,N_24599,N_24657);
nand U25059 (N_25059,N_24604,N_24901);
and U25060 (N_25060,N_24957,N_24986);
and U25061 (N_25061,N_24848,N_24945);
or U25062 (N_25062,N_24630,N_24771);
xnor U25063 (N_25063,N_24646,N_24628);
or U25064 (N_25064,N_24633,N_24617);
nand U25065 (N_25065,N_24509,N_24971);
nor U25066 (N_25066,N_24519,N_24607);
nand U25067 (N_25067,N_24735,N_24962);
nand U25068 (N_25068,N_24725,N_24871);
xnor U25069 (N_25069,N_24547,N_24992);
and U25070 (N_25070,N_24768,N_24603);
and U25071 (N_25071,N_24627,N_24642);
or U25072 (N_25072,N_24767,N_24558);
nand U25073 (N_25073,N_24920,N_24911);
and U25074 (N_25074,N_24934,N_24650);
xnor U25075 (N_25075,N_24734,N_24889);
and U25076 (N_25076,N_24909,N_24591);
or U25077 (N_25077,N_24883,N_24540);
or U25078 (N_25078,N_24960,N_24795);
or U25079 (N_25079,N_24666,N_24629);
and U25080 (N_25080,N_24638,N_24921);
xor U25081 (N_25081,N_24953,N_24805);
nor U25082 (N_25082,N_24748,N_24856);
nand U25083 (N_25083,N_24648,N_24689);
nand U25084 (N_25084,N_24643,N_24718);
nand U25085 (N_25085,N_24637,N_24548);
xor U25086 (N_25086,N_24674,N_24844);
nor U25087 (N_25087,N_24846,N_24552);
nand U25088 (N_25088,N_24828,N_24565);
nand U25089 (N_25089,N_24667,N_24931);
nand U25090 (N_25090,N_24746,N_24763);
nand U25091 (N_25091,N_24991,N_24881);
xnor U25092 (N_25092,N_24798,N_24974);
nor U25093 (N_25093,N_24765,N_24787);
nand U25094 (N_25094,N_24518,N_24823);
xor U25095 (N_25095,N_24728,N_24651);
and U25096 (N_25096,N_24944,N_24585);
or U25097 (N_25097,N_24707,N_24579);
xor U25098 (N_25098,N_24504,N_24562);
and U25099 (N_25099,N_24853,N_24967);
nand U25100 (N_25100,N_24750,N_24843);
xnor U25101 (N_25101,N_24511,N_24661);
and U25102 (N_25102,N_24863,N_24662);
nand U25103 (N_25103,N_24658,N_24736);
xor U25104 (N_25104,N_24759,N_24952);
xnor U25105 (N_25105,N_24685,N_24665);
nand U25106 (N_25106,N_24969,N_24696);
nor U25107 (N_25107,N_24913,N_24564);
or U25108 (N_25108,N_24508,N_24758);
nand U25109 (N_25109,N_24800,N_24517);
nor U25110 (N_25110,N_24716,N_24621);
or U25111 (N_25111,N_24870,N_24717);
nor U25112 (N_25112,N_24928,N_24507);
xor U25113 (N_25113,N_24812,N_24899);
nor U25114 (N_25114,N_24797,N_24705);
and U25115 (N_25115,N_24681,N_24584);
nor U25116 (N_25116,N_24656,N_24514);
or U25117 (N_25117,N_24885,N_24859);
or U25118 (N_25118,N_24818,N_24532);
or U25119 (N_25119,N_24539,N_24675);
nand U25120 (N_25120,N_24876,N_24993);
nand U25121 (N_25121,N_24950,N_24587);
or U25122 (N_25122,N_24522,N_24724);
xor U25123 (N_25123,N_24989,N_24891);
nor U25124 (N_25124,N_24997,N_24723);
nand U25125 (N_25125,N_24506,N_24873);
nor U25126 (N_25126,N_24613,N_24597);
and U25127 (N_25127,N_24773,N_24618);
and U25128 (N_25128,N_24520,N_24738);
and U25129 (N_25129,N_24531,N_24781);
nor U25130 (N_25130,N_24521,N_24880);
or U25131 (N_25131,N_24719,N_24793);
nand U25132 (N_25132,N_24568,N_24850);
xnor U25133 (N_25133,N_24694,N_24903);
and U25134 (N_25134,N_24868,N_24817);
xnor U25135 (N_25135,N_24935,N_24799);
and U25136 (N_25136,N_24614,N_24524);
or U25137 (N_25137,N_24865,N_24513);
nand U25138 (N_25138,N_24753,N_24570);
nor U25139 (N_25139,N_24998,N_24512);
nor U25140 (N_25140,N_24594,N_24860);
or U25141 (N_25141,N_24566,N_24851);
xor U25142 (N_25142,N_24822,N_24976);
or U25143 (N_25143,N_24721,N_24874);
nand U25144 (N_25144,N_24757,N_24849);
or U25145 (N_25145,N_24528,N_24755);
nor U25146 (N_25146,N_24893,N_24908);
and U25147 (N_25147,N_24840,N_24690);
xnor U25148 (N_25148,N_24898,N_24902);
xnor U25149 (N_25149,N_24785,N_24806);
xnor U25150 (N_25150,N_24542,N_24833);
or U25151 (N_25151,N_24634,N_24535);
or U25152 (N_25152,N_24831,N_24838);
xor U25153 (N_25153,N_24611,N_24583);
or U25154 (N_25154,N_24644,N_24640);
xnor U25155 (N_25155,N_24779,N_24861);
nand U25156 (N_25156,N_24747,N_24709);
and U25157 (N_25157,N_24830,N_24754);
nor U25158 (N_25158,N_24698,N_24939);
and U25159 (N_25159,N_24841,N_24919);
xnor U25160 (N_25160,N_24559,N_24737);
nor U25161 (N_25161,N_24804,N_24744);
xor U25162 (N_25162,N_24680,N_24927);
or U25163 (N_25163,N_24730,N_24814);
nand U25164 (N_25164,N_24788,N_24770);
or U25165 (N_25165,N_24796,N_24929);
or U25166 (N_25166,N_24857,N_24636);
xnor U25167 (N_25167,N_24816,N_24801);
or U25168 (N_25168,N_24942,N_24896);
nand U25169 (N_25169,N_24673,N_24905);
nor U25170 (N_25170,N_24985,N_24892);
and U25171 (N_25171,N_24869,N_24659);
and U25172 (N_25172,N_24574,N_24682);
xnor U25173 (N_25173,N_24686,N_24515);
and U25174 (N_25174,N_24839,N_24756);
and U25175 (N_25175,N_24772,N_24820);
or U25176 (N_25176,N_24970,N_24510);
nor U25177 (N_25177,N_24829,N_24631);
nor U25178 (N_25178,N_24752,N_24847);
and U25179 (N_25179,N_24581,N_24888);
or U25180 (N_25180,N_24729,N_24639);
or U25181 (N_25181,N_24984,N_24917);
and U25182 (N_25182,N_24937,N_24954);
or U25183 (N_25183,N_24502,N_24894);
nor U25184 (N_25184,N_24688,N_24742);
xnor U25185 (N_25185,N_24537,N_24626);
nand U25186 (N_25186,N_24503,N_24578);
and U25187 (N_25187,N_24715,N_24605);
nand U25188 (N_25188,N_24999,N_24625);
and U25189 (N_25189,N_24609,N_24784);
or U25190 (N_25190,N_24904,N_24832);
or U25191 (N_25191,N_24964,N_24808);
xnor U25192 (N_25192,N_24872,N_24761);
xor U25193 (N_25193,N_24782,N_24619);
or U25194 (N_25194,N_24933,N_24878);
and U25195 (N_25195,N_24775,N_24943);
and U25196 (N_25196,N_24955,N_24702);
and U25197 (N_25197,N_24963,N_24864);
or U25198 (N_25198,N_24726,N_24692);
xnor U25199 (N_25199,N_24710,N_24923);
and U25200 (N_25200,N_24538,N_24560);
nor U25201 (N_25201,N_24803,N_24783);
nand U25202 (N_25202,N_24714,N_24988);
or U25203 (N_25203,N_24569,N_24877);
nor U25204 (N_25204,N_24995,N_24526);
xor U25205 (N_25205,N_24956,N_24610);
xor U25206 (N_25206,N_24549,N_24527);
and U25207 (N_25207,N_24670,N_24600);
nor U25208 (N_25208,N_24741,N_24807);
and U25209 (N_25209,N_24739,N_24550);
and U25210 (N_25210,N_24596,N_24612);
nor U25211 (N_25211,N_24930,N_24572);
nor U25212 (N_25212,N_24852,N_24505);
or U25213 (N_25213,N_24745,N_24655);
or U25214 (N_25214,N_24975,N_24713);
nor U25215 (N_25215,N_24676,N_24981);
nand U25216 (N_25216,N_24978,N_24529);
nor U25217 (N_25217,N_24551,N_24586);
nand U25218 (N_25218,N_24932,N_24858);
nand U25219 (N_25219,N_24663,N_24693);
or U25220 (N_25220,N_24826,N_24810);
or U25221 (N_25221,N_24762,N_24580);
nor U25222 (N_25222,N_24654,N_24500);
or U25223 (N_25223,N_24951,N_24733);
nand U25224 (N_25224,N_24875,N_24523);
or U25225 (N_25225,N_24576,N_24602);
nand U25226 (N_25226,N_24700,N_24802);
xnor U25227 (N_25227,N_24809,N_24649);
and U25228 (N_25228,N_24697,N_24835);
nand U25229 (N_25229,N_24699,N_24641);
and U25230 (N_25230,N_24912,N_24836);
nor U25231 (N_25231,N_24554,N_24684);
xor U25232 (N_25232,N_24827,N_24965);
nor U25233 (N_25233,N_24652,N_24980);
nand U25234 (N_25234,N_24653,N_24959);
or U25235 (N_25235,N_24546,N_24764);
nand U25236 (N_25236,N_24924,N_24792);
nor U25237 (N_25237,N_24732,N_24561);
or U25238 (N_25238,N_24996,N_24774);
xnor U25239 (N_25239,N_24780,N_24987);
or U25240 (N_25240,N_24624,N_24720);
and U25241 (N_25241,N_24556,N_24983);
and U25242 (N_25242,N_24622,N_24879);
and U25243 (N_25243,N_24910,N_24815);
nand U25244 (N_25244,N_24544,N_24968);
nor U25245 (N_25245,N_24895,N_24776);
xor U25246 (N_25246,N_24811,N_24834);
nor U25247 (N_25247,N_24571,N_24915);
nor U25248 (N_25248,N_24582,N_24668);
and U25249 (N_25249,N_24824,N_24533);
nor U25250 (N_25250,N_24772,N_24996);
or U25251 (N_25251,N_24917,N_24543);
or U25252 (N_25252,N_24900,N_24929);
xor U25253 (N_25253,N_24924,N_24729);
nand U25254 (N_25254,N_24539,N_24898);
or U25255 (N_25255,N_24514,N_24831);
or U25256 (N_25256,N_24645,N_24842);
nand U25257 (N_25257,N_24826,N_24766);
xnor U25258 (N_25258,N_24916,N_24694);
or U25259 (N_25259,N_24539,N_24551);
nor U25260 (N_25260,N_24656,N_24570);
nor U25261 (N_25261,N_24824,N_24858);
nand U25262 (N_25262,N_24566,N_24662);
and U25263 (N_25263,N_24503,N_24671);
nor U25264 (N_25264,N_24806,N_24555);
and U25265 (N_25265,N_24899,N_24968);
or U25266 (N_25266,N_24752,N_24831);
nand U25267 (N_25267,N_24571,N_24623);
nand U25268 (N_25268,N_24721,N_24996);
or U25269 (N_25269,N_24677,N_24599);
xnor U25270 (N_25270,N_24646,N_24840);
nor U25271 (N_25271,N_24516,N_24766);
or U25272 (N_25272,N_24972,N_24779);
nor U25273 (N_25273,N_24705,N_24701);
nor U25274 (N_25274,N_24984,N_24883);
or U25275 (N_25275,N_24553,N_24883);
nand U25276 (N_25276,N_24575,N_24924);
nand U25277 (N_25277,N_24773,N_24691);
xnor U25278 (N_25278,N_24689,N_24752);
and U25279 (N_25279,N_24926,N_24816);
and U25280 (N_25280,N_24654,N_24604);
xor U25281 (N_25281,N_24595,N_24835);
xor U25282 (N_25282,N_24811,N_24852);
nor U25283 (N_25283,N_24506,N_24822);
nor U25284 (N_25284,N_24942,N_24691);
xor U25285 (N_25285,N_24814,N_24888);
or U25286 (N_25286,N_24945,N_24819);
nand U25287 (N_25287,N_24884,N_24907);
or U25288 (N_25288,N_24900,N_24892);
nor U25289 (N_25289,N_24939,N_24988);
nand U25290 (N_25290,N_24698,N_24738);
and U25291 (N_25291,N_24860,N_24622);
xor U25292 (N_25292,N_24786,N_24975);
or U25293 (N_25293,N_24798,N_24629);
xor U25294 (N_25294,N_24868,N_24636);
xor U25295 (N_25295,N_24711,N_24700);
or U25296 (N_25296,N_24897,N_24834);
and U25297 (N_25297,N_24936,N_24831);
nor U25298 (N_25298,N_24758,N_24899);
xor U25299 (N_25299,N_24733,N_24894);
and U25300 (N_25300,N_24975,N_24668);
nand U25301 (N_25301,N_24674,N_24996);
nor U25302 (N_25302,N_24522,N_24971);
or U25303 (N_25303,N_24626,N_24864);
or U25304 (N_25304,N_24910,N_24866);
or U25305 (N_25305,N_24516,N_24667);
nand U25306 (N_25306,N_24508,N_24506);
xor U25307 (N_25307,N_24826,N_24666);
and U25308 (N_25308,N_24758,N_24772);
nor U25309 (N_25309,N_24832,N_24915);
nand U25310 (N_25310,N_24566,N_24579);
and U25311 (N_25311,N_24846,N_24665);
nor U25312 (N_25312,N_24551,N_24559);
xnor U25313 (N_25313,N_24580,N_24912);
nand U25314 (N_25314,N_24567,N_24590);
nor U25315 (N_25315,N_24759,N_24506);
or U25316 (N_25316,N_24621,N_24947);
xnor U25317 (N_25317,N_24653,N_24662);
nand U25318 (N_25318,N_24523,N_24796);
nand U25319 (N_25319,N_24501,N_24581);
and U25320 (N_25320,N_24750,N_24897);
nor U25321 (N_25321,N_24703,N_24921);
and U25322 (N_25322,N_24518,N_24865);
or U25323 (N_25323,N_24726,N_24857);
nand U25324 (N_25324,N_24737,N_24526);
nand U25325 (N_25325,N_24935,N_24689);
nand U25326 (N_25326,N_24886,N_24629);
and U25327 (N_25327,N_24532,N_24693);
and U25328 (N_25328,N_24959,N_24687);
or U25329 (N_25329,N_24992,N_24823);
xor U25330 (N_25330,N_24948,N_24996);
xnor U25331 (N_25331,N_24733,N_24634);
or U25332 (N_25332,N_24600,N_24895);
and U25333 (N_25333,N_24901,N_24641);
and U25334 (N_25334,N_24614,N_24914);
nor U25335 (N_25335,N_24719,N_24506);
xor U25336 (N_25336,N_24522,N_24728);
nand U25337 (N_25337,N_24710,N_24696);
and U25338 (N_25338,N_24864,N_24825);
and U25339 (N_25339,N_24995,N_24961);
nand U25340 (N_25340,N_24545,N_24731);
nor U25341 (N_25341,N_24522,N_24663);
nand U25342 (N_25342,N_24894,N_24992);
and U25343 (N_25343,N_24675,N_24828);
and U25344 (N_25344,N_24600,N_24840);
nand U25345 (N_25345,N_24962,N_24949);
xnor U25346 (N_25346,N_24729,N_24666);
nand U25347 (N_25347,N_24523,N_24825);
and U25348 (N_25348,N_24803,N_24503);
or U25349 (N_25349,N_24601,N_24650);
nand U25350 (N_25350,N_24780,N_24578);
and U25351 (N_25351,N_24646,N_24558);
nor U25352 (N_25352,N_24729,N_24896);
nor U25353 (N_25353,N_24913,N_24724);
nor U25354 (N_25354,N_24987,N_24773);
nand U25355 (N_25355,N_24553,N_24780);
or U25356 (N_25356,N_24818,N_24644);
nor U25357 (N_25357,N_24767,N_24937);
and U25358 (N_25358,N_24650,N_24839);
nand U25359 (N_25359,N_24764,N_24666);
and U25360 (N_25360,N_24579,N_24995);
and U25361 (N_25361,N_24656,N_24753);
and U25362 (N_25362,N_24956,N_24970);
xnor U25363 (N_25363,N_24690,N_24952);
and U25364 (N_25364,N_24673,N_24912);
nor U25365 (N_25365,N_24720,N_24698);
nor U25366 (N_25366,N_24861,N_24892);
or U25367 (N_25367,N_24617,N_24840);
nor U25368 (N_25368,N_24837,N_24516);
nand U25369 (N_25369,N_24942,N_24793);
and U25370 (N_25370,N_24723,N_24978);
nor U25371 (N_25371,N_24693,N_24700);
xnor U25372 (N_25372,N_24970,N_24928);
and U25373 (N_25373,N_24780,N_24696);
and U25374 (N_25374,N_24762,N_24830);
or U25375 (N_25375,N_24967,N_24568);
and U25376 (N_25376,N_24798,N_24973);
nor U25377 (N_25377,N_24705,N_24956);
xor U25378 (N_25378,N_24592,N_24559);
or U25379 (N_25379,N_24607,N_24798);
nor U25380 (N_25380,N_24953,N_24606);
and U25381 (N_25381,N_24513,N_24924);
or U25382 (N_25382,N_24578,N_24734);
xor U25383 (N_25383,N_24700,N_24671);
or U25384 (N_25384,N_24914,N_24581);
nor U25385 (N_25385,N_24688,N_24850);
or U25386 (N_25386,N_24513,N_24798);
nand U25387 (N_25387,N_24825,N_24999);
nor U25388 (N_25388,N_24959,N_24627);
nor U25389 (N_25389,N_24769,N_24635);
nor U25390 (N_25390,N_24799,N_24779);
nor U25391 (N_25391,N_24593,N_24633);
nor U25392 (N_25392,N_24930,N_24746);
and U25393 (N_25393,N_24703,N_24757);
or U25394 (N_25394,N_24536,N_24717);
nand U25395 (N_25395,N_24697,N_24587);
or U25396 (N_25396,N_24650,N_24855);
xnor U25397 (N_25397,N_24602,N_24747);
xnor U25398 (N_25398,N_24955,N_24695);
and U25399 (N_25399,N_24631,N_24880);
nor U25400 (N_25400,N_24860,N_24849);
xnor U25401 (N_25401,N_24860,N_24522);
or U25402 (N_25402,N_24624,N_24949);
xnor U25403 (N_25403,N_24861,N_24544);
nand U25404 (N_25404,N_24754,N_24816);
xor U25405 (N_25405,N_24538,N_24596);
and U25406 (N_25406,N_24832,N_24837);
xor U25407 (N_25407,N_24699,N_24872);
xor U25408 (N_25408,N_24973,N_24980);
or U25409 (N_25409,N_24984,N_24959);
nand U25410 (N_25410,N_24836,N_24786);
and U25411 (N_25411,N_24777,N_24645);
and U25412 (N_25412,N_24910,N_24594);
xor U25413 (N_25413,N_24556,N_24766);
nor U25414 (N_25414,N_24533,N_24830);
or U25415 (N_25415,N_24555,N_24517);
and U25416 (N_25416,N_24808,N_24798);
nand U25417 (N_25417,N_24616,N_24744);
nand U25418 (N_25418,N_24663,N_24823);
xor U25419 (N_25419,N_24980,N_24923);
xor U25420 (N_25420,N_24893,N_24811);
nand U25421 (N_25421,N_24800,N_24850);
nor U25422 (N_25422,N_24792,N_24840);
nor U25423 (N_25423,N_24858,N_24868);
xnor U25424 (N_25424,N_24851,N_24597);
xor U25425 (N_25425,N_24864,N_24749);
and U25426 (N_25426,N_24584,N_24635);
nand U25427 (N_25427,N_24888,N_24963);
and U25428 (N_25428,N_24635,N_24659);
and U25429 (N_25429,N_24897,N_24912);
or U25430 (N_25430,N_24531,N_24632);
nand U25431 (N_25431,N_24925,N_24938);
nand U25432 (N_25432,N_24874,N_24719);
nor U25433 (N_25433,N_24609,N_24558);
nor U25434 (N_25434,N_24767,N_24524);
and U25435 (N_25435,N_24593,N_24613);
and U25436 (N_25436,N_24531,N_24877);
nor U25437 (N_25437,N_24659,N_24751);
or U25438 (N_25438,N_24726,N_24809);
or U25439 (N_25439,N_24971,N_24606);
nand U25440 (N_25440,N_24990,N_24667);
xor U25441 (N_25441,N_24912,N_24654);
xnor U25442 (N_25442,N_24816,N_24679);
and U25443 (N_25443,N_24753,N_24931);
or U25444 (N_25444,N_24911,N_24703);
nor U25445 (N_25445,N_24583,N_24508);
nor U25446 (N_25446,N_24605,N_24987);
nand U25447 (N_25447,N_24633,N_24831);
nand U25448 (N_25448,N_24777,N_24735);
xnor U25449 (N_25449,N_24764,N_24564);
or U25450 (N_25450,N_24698,N_24578);
and U25451 (N_25451,N_24717,N_24805);
xor U25452 (N_25452,N_24979,N_24713);
nor U25453 (N_25453,N_24678,N_24693);
nand U25454 (N_25454,N_24874,N_24819);
nand U25455 (N_25455,N_24591,N_24607);
xor U25456 (N_25456,N_24935,N_24605);
or U25457 (N_25457,N_24500,N_24919);
or U25458 (N_25458,N_24543,N_24721);
and U25459 (N_25459,N_24573,N_24889);
nor U25460 (N_25460,N_24644,N_24733);
xor U25461 (N_25461,N_24803,N_24809);
nor U25462 (N_25462,N_24580,N_24505);
xor U25463 (N_25463,N_24754,N_24900);
nor U25464 (N_25464,N_24620,N_24655);
or U25465 (N_25465,N_24652,N_24536);
and U25466 (N_25466,N_24973,N_24666);
nand U25467 (N_25467,N_24635,N_24521);
and U25468 (N_25468,N_24990,N_24838);
nor U25469 (N_25469,N_24968,N_24785);
nor U25470 (N_25470,N_24529,N_24790);
nand U25471 (N_25471,N_24867,N_24683);
xnor U25472 (N_25472,N_24878,N_24975);
xor U25473 (N_25473,N_24799,N_24694);
or U25474 (N_25474,N_24779,N_24874);
and U25475 (N_25475,N_24756,N_24917);
nor U25476 (N_25476,N_24612,N_24721);
xnor U25477 (N_25477,N_24978,N_24972);
nand U25478 (N_25478,N_24940,N_24840);
nand U25479 (N_25479,N_24778,N_24512);
nor U25480 (N_25480,N_24526,N_24509);
xnor U25481 (N_25481,N_24551,N_24732);
and U25482 (N_25482,N_24961,N_24749);
nor U25483 (N_25483,N_24669,N_24657);
nor U25484 (N_25484,N_24741,N_24752);
nand U25485 (N_25485,N_24824,N_24742);
nand U25486 (N_25486,N_24694,N_24633);
nor U25487 (N_25487,N_24732,N_24841);
and U25488 (N_25488,N_24860,N_24646);
or U25489 (N_25489,N_24823,N_24975);
nor U25490 (N_25490,N_24975,N_24901);
nand U25491 (N_25491,N_24515,N_24590);
xnor U25492 (N_25492,N_24773,N_24538);
nor U25493 (N_25493,N_24723,N_24520);
xnor U25494 (N_25494,N_24538,N_24787);
xor U25495 (N_25495,N_24582,N_24629);
and U25496 (N_25496,N_24759,N_24771);
nand U25497 (N_25497,N_24757,N_24586);
nand U25498 (N_25498,N_24516,N_24920);
nor U25499 (N_25499,N_24640,N_24683);
xor U25500 (N_25500,N_25070,N_25479);
xnor U25501 (N_25501,N_25171,N_25452);
nor U25502 (N_25502,N_25419,N_25245);
nand U25503 (N_25503,N_25469,N_25020);
and U25504 (N_25504,N_25300,N_25333);
or U25505 (N_25505,N_25236,N_25373);
or U25506 (N_25506,N_25259,N_25000);
or U25507 (N_25507,N_25191,N_25451);
and U25508 (N_25508,N_25134,N_25340);
nand U25509 (N_25509,N_25278,N_25196);
xor U25510 (N_25510,N_25455,N_25337);
or U25511 (N_25511,N_25012,N_25114);
nand U25512 (N_25512,N_25009,N_25464);
xor U25513 (N_25513,N_25431,N_25332);
or U25514 (N_25514,N_25211,N_25054);
nand U25515 (N_25515,N_25076,N_25263);
nor U25516 (N_25516,N_25166,N_25417);
or U25517 (N_25517,N_25477,N_25237);
nand U25518 (N_25518,N_25446,N_25097);
and U25519 (N_25519,N_25124,N_25405);
or U25520 (N_25520,N_25344,N_25346);
and U25521 (N_25521,N_25163,N_25193);
nor U25522 (N_25522,N_25302,N_25434);
or U25523 (N_25523,N_25383,N_25125);
and U25524 (N_25524,N_25246,N_25024);
nand U25525 (N_25525,N_25198,N_25031);
nand U25526 (N_25526,N_25287,N_25017);
or U25527 (N_25527,N_25232,N_25338);
xor U25528 (N_25528,N_25055,N_25056);
nand U25529 (N_25529,N_25361,N_25286);
nor U25530 (N_25530,N_25248,N_25227);
xnor U25531 (N_25531,N_25242,N_25182);
and U25532 (N_25532,N_25058,N_25436);
and U25533 (N_25533,N_25352,N_25366);
and U25534 (N_25534,N_25268,N_25398);
and U25535 (N_25535,N_25051,N_25129);
and U25536 (N_25536,N_25491,N_25316);
nand U25537 (N_25537,N_25425,N_25084);
nor U25538 (N_25538,N_25450,N_25345);
nor U25539 (N_25539,N_25485,N_25011);
xnor U25540 (N_25540,N_25174,N_25381);
nand U25541 (N_25541,N_25035,N_25492);
or U25542 (N_25542,N_25014,N_25433);
nand U25543 (N_25543,N_25355,N_25325);
and U25544 (N_25544,N_25386,N_25388);
nand U25545 (N_25545,N_25207,N_25402);
nand U25546 (N_25546,N_25271,N_25208);
or U25547 (N_25547,N_25277,N_25162);
xor U25548 (N_25548,N_25112,N_25314);
nand U25549 (N_25549,N_25418,N_25001);
nand U25550 (N_25550,N_25221,N_25487);
nor U25551 (N_25551,N_25224,N_25078);
and U25552 (N_25552,N_25230,N_25247);
nor U25553 (N_25553,N_25336,N_25194);
nand U25554 (N_25554,N_25441,N_25215);
and U25555 (N_25555,N_25362,N_25180);
nor U25556 (N_25556,N_25347,N_25257);
or U25557 (N_25557,N_25132,N_25019);
or U25558 (N_25558,N_25308,N_25157);
and U25559 (N_25559,N_25382,N_25113);
nor U25560 (N_25560,N_25372,N_25497);
nand U25561 (N_25561,N_25251,N_25442);
and U25562 (N_25562,N_25213,N_25266);
nor U25563 (N_25563,N_25393,N_25123);
or U25564 (N_25564,N_25460,N_25034);
or U25565 (N_25565,N_25197,N_25489);
xor U25566 (N_25566,N_25292,N_25092);
and U25567 (N_25567,N_25065,N_25411);
nand U25568 (N_25568,N_25146,N_25149);
or U25569 (N_25569,N_25397,N_25186);
nor U25570 (N_25570,N_25088,N_25407);
nand U25571 (N_25571,N_25470,N_25262);
xor U25572 (N_25572,N_25150,N_25368);
and U25573 (N_25573,N_25404,N_25095);
nand U25574 (N_25574,N_25119,N_25235);
and U25575 (N_25575,N_25281,N_25484);
or U25576 (N_25576,N_25108,N_25323);
nand U25577 (N_25577,N_25151,N_25288);
and U25578 (N_25578,N_25304,N_25253);
nand U25579 (N_25579,N_25170,N_25305);
xor U25580 (N_25580,N_25395,N_25496);
and U25581 (N_25581,N_25106,N_25083);
nor U25582 (N_25582,N_25403,N_25075);
and U25583 (N_25583,N_25053,N_25392);
xnor U25584 (N_25584,N_25057,N_25326);
nor U25585 (N_25585,N_25364,N_25175);
or U25586 (N_25586,N_25309,N_25141);
nand U25587 (N_25587,N_25466,N_25199);
nor U25588 (N_25588,N_25093,N_25423);
nand U25589 (N_25589,N_25110,N_25293);
and U25590 (N_25590,N_25069,N_25426);
nand U25591 (N_25591,N_25152,N_25313);
and U25592 (N_25592,N_25115,N_25252);
xnor U25593 (N_25593,N_25318,N_25006);
and U25594 (N_25594,N_25297,N_25080);
and U25595 (N_25595,N_25026,N_25254);
and U25596 (N_25596,N_25354,N_25087);
or U25597 (N_25597,N_25127,N_25081);
xnor U25598 (N_25598,N_25273,N_25371);
nand U25599 (N_25599,N_25013,N_25463);
and U25600 (N_25600,N_25089,N_25444);
and U25601 (N_25601,N_25155,N_25408);
and U25602 (N_25602,N_25330,N_25234);
and U25603 (N_25603,N_25422,N_25189);
and U25604 (N_25604,N_25212,N_25285);
nor U25605 (N_25605,N_25091,N_25178);
and U25606 (N_25606,N_25401,N_25130);
and U25607 (N_25607,N_25066,N_25409);
nor U25608 (N_25608,N_25317,N_25062);
or U25609 (N_25609,N_25482,N_25439);
or U25610 (N_25610,N_25427,N_25121);
xnor U25611 (N_25611,N_25241,N_25290);
nand U25612 (N_25612,N_25493,N_25499);
and U25613 (N_25613,N_25086,N_25027);
nor U25614 (N_25614,N_25003,N_25226);
xnor U25615 (N_25615,N_25298,N_25320);
xnor U25616 (N_25616,N_25453,N_25424);
and U25617 (N_25617,N_25435,N_25385);
xor U25618 (N_25618,N_25459,N_25188);
nor U25619 (N_25619,N_25265,N_25085);
xor U25620 (N_25620,N_25454,N_25032);
nor U25621 (N_25621,N_25131,N_25465);
xor U25622 (N_25622,N_25160,N_25218);
or U25623 (N_25623,N_25378,N_25339);
xor U25624 (N_25624,N_25445,N_25274);
or U25625 (N_25625,N_25214,N_25486);
nor U25626 (N_25626,N_25359,N_25322);
nor U25627 (N_25627,N_25367,N_25349);
nand U25628 (N_25628,N_25416,N_25190);
nor U25629 (N_25629,N_25147,N_25033);
or U25630 (N_25630,N_25348,N_25467);
xor U25631 (N_25631,N_25156,N_25135);
and U25632 (N_25632,N_25133,N_25279);
nand U25633 (N_25633,N_25261,N_25036);
nand U25634 (N_25634,N_25443,N_25413);
or U25635 (N_25635,N_25100,N_25468);
and U25636 (N_25636,N_25421,N_25018);
xnor U25637 (N_25637,N_25391,N_25449);
and U25638 (N_25638,N_25428,N_25291);
and U25639 (N_25639,N_25143,N_25165);
and U25640 (N_25640,N_25229,N_25406);
and U25641 (N_25641,N_25046,N_25052);
or U25642 (N_25642,N_25329,N_25250);
xor U25643 (N_25643,N_25118,N_25311);
and U25644 (N_25644,N_25415,N_25039);
nand U25645 (N_25645,N_25111,N_25360);
nand U25646 (N_25646,N_25101,N_25310);
xor U25647 (N_25647,N_25374,N_25233);
and U25648 (N_25648,N_25049,N_25181);
or U25649 (N_25649,N_25341,N_25136);
or U25650 (N_25650,N_25267,N_25161);
or U25651 (N_25651,N_25358,N_25475);
nand U25652 (N_25652,N_25357,N_25370);
and U25653 (N_25653,N_25239,N_25353);
xor U25654 (N_25654,N_25447,N_25380);
nand U25655 (N_25655,N_25255,N_25072);
nor U25656 (N_25656,N_25389,N_25045);
xnor U25657 (N_25657,N_25437,N_25016);
xor U25658 (N_25658,N_25047,N_25275);
and U25659 (N_25659,N_25159,N_25327);
xor U25660 (N_25660,N_25041,N_25138);
nor U25661 (N_25661,N_25260,N_25289);
and U25662 (N_25662,N_25264,N_25176);
xnor U25663 (N_25663,N_25420,N_25319);
nand U25664 (N_25664,N_25154,N_25205);
nor U25665 (N_25665,N_25128,N_25270);
and U25666 (N_25666,N_25042,N_25328);
nor U25667 (N_25667,N_25394,N_25210);
and U25668 (N_25668,N_25167,N_25342);
and U25669 (N_25669,N_25483,N_25272);
nand U25670 (N_25670,N_25117,N_25022);
nand U25671 (N_25671,N_25010,N_25387);
or U25672 (N_25672,N_25312,N_25356);
or U25673 (N_25673,N_25140,N_25334);
xnor U25674 (N_25674,N_25096,N_25461);
xnor U25675 (N_25675,N_25158,N_25025);
xor U25676 (N_25676,N_25144,N_25172);
and U25677 (N_25677,N_25220,N_25480);
nor U25678 (N_25678,N_25440,N_25094);
and U25679 (N_25679,N_25050,N_25412);
xnor U25680 (N_25680,N_25063,N_25153);
xor U25681 (N_25681,N_25185,N_25021);
xnor U25682 (N_25682,N_25490,N_25369);
nor U25683 (N_25683,N_25216,N_25301);
and U25684 (N_25684,N_25145,N_25122);
or U25685 (N_25685,N_25195,N_25282);
nand U25686 (N_25686,N_25296,N_25201);
nand U25687 (N_25687,N_25476,N_25116);
nor U25688 (N_25688,N_25177,N_25284);
nand U25689 (N_25689,N_25432,N_25200);
nand U25690 (N_25690,N_25410,N_25377);
nor U25691 (N_25691,N_25375,N_25472);
xor U25692 (N_25692,N_25462,N_25139);
nand U25693 (N_25693,N_25228,N_25044);
nor U25694 (N_25694,N_25067,N_25028);
nand U25695 (N_25695,N_25007,N_25074);
xnor U25696 (N_25696,N_25280,N_25038);
nand U25697 (N_25697,N_25495,N_25498);
xnor U25698 (N_25698,N_25457,N_25098);
or U25699 (N_25699,N_25306,N_25077);
nor U25700 (N_25700,N_25004,N_25494);
or U25701 (N_25701,N_25448,N_25064);
and U25702 (N_25702,N_25202,N_25090);
nor U25703 (N_25703,N_25008,N_25040);
or U25704 (N_25704,N_25335,N_25473);
or U25705 (N_25705,N_25376,N_25183);
xnor U25706 (N_25706,N_25294,N_25184);
nor U25707 (N_25707,N_25071,N_25488);
and U25708 (N_25708,N_25173,N_25206);
and U25709 (N_25709,N_25225,N_25363);
or U25710 (N_25710,N_25307,N_25192);
or U25711 (N_25711,N_25379,N_25179);
nand U25712 (N_25712,N_25295,N_25283);
nor U25713 (N_25713,N_25299,N_25037);
nor U25714 (N_25714,N_25209,N_25429);
and U25715 (N_25715,N_25105,N_25082);
nand U25716 (N_25716,N_25169,N_25438);
and U25717 (N_25717,N_25243,N_25148);
nand U25718 (N_25718,N_25474,N_25456);
nor U25719 (N_25719,N_25244,N_25269);
and U25720 (N_25720,N_25217,N_25126);
xor U25721 (N_25721,N_25390,N_25331);
and U25722 (N_25722,N_25399,N_25015);
or U25723 (N_25723,N_25079,N_25107);
nand U25724 (N_25724,N_25073,N_25023);
or U25725 (N_25725,N_25137,N_25481);
nor U25726 (N_25726,N_25168,N_25396);
nor U25727 (N_25727,N_25231,N_25164);
nand U25728 (N_25728,N_25030,N_25458);
and U25729 (N_25729,N_25276,N_25099);
and U25730 (N_25730,N_25222,N_25256);
and U25731 (N_25731,N_25187,N_25384);
xor U25732 (N_25732,N_25043,N_25343);
xnor U25733 (N_25733,N_25059,N_25061);
nor U25734 (N_25734,N_25400,N_25350);
xor U25735 (N_25735,N_25414,N_25471);
nand U25736 (N_25736,N_25238,N_25321);
xor U25737 (N_25737,N_25223,N_25478);
and U25738 (N_25738,N_25068,N_25103);
xnor U25739 (N_25739,N_25048,N_25029);
nand U25740 (N_25740,N_25005,N_25351);
or U25741 (N_25741,N_25365,N_25324);
and U25742 (N_25742,N_25249,N_25203);
nor U25743 (N_25743,N_25104,N_25102);
or U25744 (N_25744,N_25120,N_25142);
nand U25745 (N_25745,N_25002,N_25109);
nand U25746 (N_25746,N_25219,N_25060);
nand U25747 (N_25747,N_25315,N_25303);
and U25748 (N_25748,N_25258,N_25240);
and U25749 (N_25749,N_25430,N_25204);
or U25750 (N_25750,N_25154,N_25238);
xor U25751 (N_25751,N_25049,N_25385);
and U25752 (N_25752,N_25311,N_25175);
xnor U25753 (N_25753,N_25247,N_25193);
nor U25754 (N_25754,N_25317,N_25045);
nor U25755 (N_25755,N_25143,N_25170);
and U25756 (N_25756,N_25131,N_25216);
nand U25757 (N_25757,N_25122,N_25483);
xor U25758 (N_25758,N_25039,N_25459);
nor U25759 (N_25759,N_25232,N_25161);
and U25760 (N_25760,N_25359,N_25353);
xor U25761 (N_25761,N_25015,N_25473);
nand U25762 (N_25762,N_25301,N_25284);
and U25763 (N_25763,N_25390,N_25306);
nor U25764 (N_25764,N_25484,N_25255);
nor U25765 (N_25765,N_25164,N_25135);
and U25766 (N_25766,N_25417,N_25215);
or U25767 (N_25767,N_25386,N_25470);
or U25768 (N_25768,N_25223,N_25312);
nor U25769 (N_25769,N_25378,N_25001);
nand U25770 (N_25770,N_25090,N_25149);
nor U25771 (N_25771,N_25386,N_25462);
xnor U25772 (N_25772,N_25325,N_25344);
or U25773 (N_25773,N_25208,N_25174);
and U25774 (N_25774,N_25317,N_25371);
nor U25775 (N_25775,N_25315,N_25335);
or U25776 (N_25776,N_25205,N_25168);
nor U25777 (N_25777,N_25299,N_25338);
nand U25778 (N_25778,N_25495,N_25289);
xor U25779 (N_25779,N_25030,N_25452);
or U25780 (N_25780,N_25224,N_25350);
xor U25781 (N_25781,N_25217,N_25472);
and U25782 (N_25782,N_25275,N_25009);
nand U25783 (N_25783,N_25224,N_25097);
and U25784 (N_25784,N_25220,N_25248);
nand U25785 (N_25785,N_25455,N_25284);
xnor U25786 (N_25786,N_25354,N_25080);
nor U25787 (N_25787,N_25182,N_25358);
xor U25788 (N_25788,N_25349,N_25425);
nor U25789 (N_25789,N_25154,N_25380);
xnor U25790 (N_25790,N_25051,N_25366);
and U25791 (N_25791,N_25209,N_25359);
and U25792 (N_25792,N_25181,N_25111);
nor U25793 (N_25793,N_25400,N_25099);
nor U25794 (N_25794,N_25160,N_25277);
nor U25795 (N_25795,N_25104,N_25141);
or U25796 (N_25796,N_25496,N_25017);
nor U25797 (N_25797,N_25232,N_25063);
nor U25798 (N_25798,N_25295,N_25066);
and U25799 (N_25799,N_25420,N_25269);
nor U25800 (N_25800,N_25383,N_25319);
nor U25801 (N_25801,N_25201,N_25034);
nor U25802 (N_25802,N_25409,N_25204);
xor U25803 (N_25803,N_25118,N_25419);
xnor U25804 (N_25804,N_25211,N_25207);
nor U25805 (N_25805,N_25284,N_25139);
nand U25806 (N_25806,N_25408,N_25252);
nor U25807 (N_25807,N_25250,N_25159);
nor U25808 (N_25808,N_25370,N_25312);
xor U25809 (N_25809,N_25042,N_25437);
nand U25810 (N_25810,N_25300,N_25341);
xnor U25811 (N_25811,N_25240,N_25101);
xor U25812 (N_25812,N_25170,N_25081);
nand U25813 (N_25813,N_25103,N_25209);
and U25814 (N_25814,N_25390,N_25273);
nand U25815 (N_25815,N_25166,N_25180);
nor U25816 (N_25816,N_25125,N_25084);
nor U25817 (N_25817,N_25216,N_25333);
nor U25818 (N_25818,N_25246,N_25288);
or U25819 (N_25819,N_25220,N_25388);
or U25820 (N_25820,N_25325,N_25153);
nand U25821 (N_25821,N_25041,N_25442);
nor U25822 (N_25822,N_25024,N_25346);
nand U25823 (N_25823,N_25481,N_25476);
and U25824 (N_25824,N_25240,N_25304);
and U25825 (N_25825,N_25232,N_25402);
nand U25826 (N_25826,N_25147,N_25344);
and U25827 (N_25827,N_25210,N_25136);
nand U25828 (N_25828,N_25471,N_25349);
nand U25829 (N_25829,N_25196,N_25192);
or U25830 (N_25830,N_25379,N_25461);
xnor U25831 (N_25831,N_25077,N_25273);
or U25832 (N_25832,N_25121,N_25323);
and U25833 (N_25833,N_25070,N_25058);
and U25834 (N_25834,N_25366,N_25264);
and U25835 (N_25835,N_25088,N_25026);
xor U25836 (N_25836,N_25352,N_25084);
xnor U25837 (N_25837,N_25250,N_25476);
nor U25838 (N_25838,N_25189,N_25385);
and U25839 (N_25839,N_25020,N_25101);
nor U25840 (N_25840,N_25268,N_25127);
xnor U25841 (N_25841,N_25330,N_25379);
nor U25842 (N_25842,N_25147,N_25423);
xnor U25843 (N_25843,N_25309,N_25195);
nand U25844 (N_25844,N_25289,N_25436);
or U25845 (N_25845,N_25099,N_25268);
and U25846 (N_25846,N_25202,N_25070);
and U25847 (N_25847,N_25000,N_25065);
or U25848 (N_25848,N_25354,N_25153);
xor U25849 (N_25849,N_25090,N_25074);
xnor U25850 (N_25850,N_25378,N_25357);
nor U25851 (N_25851,N_25431,N_25182);
or U25852 (N_25852,N_25338,N_25186);
or U25853 (N_25853,N_25274,N_25248);
nand U25854 (N_25854,N_25460,N_25298);
nand U25855 (N_25855,N_25103,N_25129);
xnor U25856 (N_25856,N_25074,N_25274);
or U25857 (N_25857,N_25491,N_25068);
and U25858 (N_25858,N_25394,N_25396);
xnor U25859 (N_25859,N_25032,N_25449);
and U25860 (N_25860,N_25365,N_25347);
nand U25861 (N_25861,N_25098,N_25160);
or U25862 (N_25862,N_25319,N_25251);
nor U25863 (N_25863,N_25324,N_25474);
xor U25864 (N_25864,N_25209,N_25305);
nand U25865 (N_25865,N_25065,N_25485);
nand U25866 (N_25866,N_25455,N_25333);
or U25867 (N_25867,N_25014,N_25027);
nand U25868 (N_25868,N_25132,N_25446);
or U25869 (N_25869,N_25226,N_25066);
nand U25870 (N_25870,N_25099,N_25424);
nand U25871 (N_25871,N_25220,N_25451);
and U25872 (N_25872,N_25054,N_25032);
nand U25873 (N_25873,N_25031,N_25158);
or U25874 (N_25874,N_25494,N_25083);
xor U25875 (N_25875,N_25161,N_25033);
or U25876 (N_25876,N_25138,N_25021);
nor U25877 (N_25877,N_25343,N_25183);
or U25878 (N_25878,N_25271,N_25293);
nand U25879 (N_25879,N_25049,N_25497);
and U25880 (N_25880,N_25142,N_25051);
nor U25881 (N_25881,N_25165,N_25169);
nor U25882 (N_25882,N_25361,N_25335);
nor U25883 (N_25883,N_25456,N_25429);
nand U25884 (N_25884,N_25087,N_25237);
nand U25885 (N_25885,N_25207,N_25171);
or U25886 (N_25886,N_25338,N_25268);
and U25887 (N_25887,N_25402,N_25228);
nor U25888 (N_25888,N_25334,N_25343);
xor U25889 (N_25889,N_25464,N_25207);
nand U25890 (N_25890,N_25209,N_25082);
or U25891 (N_25891,N_25028,N_25047);
nor U25892 (N_25892,N_25232,N_25340);
or U25893 (N_25893,N_25239,N_25452);
and U25894 (N_25894,N_25467,N_25388);
nor U25895 (N_25895,N_25163,N_25206);
or U25896 (N_25896,N_25307,N_25238);
or U25897 (N_25897,N_25051,N_25425);
or U25898 (N_25898,N_25021,N_25032);
nand U25899 (N_25899,N_25497,N_25228);
nor U25900 (N_25900,N_25210,N_25032);
or U25901 (N_25901,N_25062,N_25009);
xor U25902 (N_25902,N_25133,N_25041);
nand U25903 (N_25903,N_25441,N_25197);
and U25904 (N_25904,N_25436,N_25294);
nand U25905 (N_25905,N_25467,N_25034);
xnor U25906 (N_25906,N_25336,N_25438);
xnor U25907 (N_25907,N_25206,N_25211);
nand U25908 (N_25908,N_25405,N_25495);
and U25909 (N_25909,N_25205,N_25148);
nor U25910 (N_25910,N_25420,N_25035);
xor U25911 (N_25911,N_25286,N_25189);
or U25912 (N_25912,N_25087,N_25449);
and U25913 (N_25913,N_25461,N_25155);
or U25914 (N_25914,N_25180,N_25463);
nand U25915 (N_25915,N_25191,N_25342);
xor U25916 (N_25916,N_25165,N_25402);
and U25917 (N_25917,N_25313,N_25361);
xor U25918 (N_25918,N_25140,N_25141);
xnor U25919 (N_25919,N_25386,N_25490);
or U25920 (N_25920,N_25112,N_25154);
or U25921 (N_25921,N_25064,N_25089);
or U25922 (N_25922,N_25348,N_25108);
and U25923 (N_25923,N_25300,N_25376);
or U25924 (N_25924,N_25391,N_25381);
xnor U25925 (N_25925,N_25128,N_25337);
or U25926 (N_25926,N_25224,N_25080);
and U25927 (N_25927,N_25190,N_25075);
nor U25928 (N_25928,N_25377,N_25071);
or U25929 (N_25929,N_25075,N_25426);
xnor U25930 (N_25930,N_25197,N_25180);
xor U25931 (N_25931,N_25006,N_25174);
xnor U25932 (N_25932,N_25132,N_25450);
xor U25933 (N_25933,N_25407,N_25290);
and U25934 (N_25934,N_25485,N_25070);
nor U25935 (N_25935,N_25375,N_25102);
nand U25936 (N_25936,N_25028,N_25452);
xor U25937 (N_25937,N_25257,N_25309);
nand U25938 (N_25938,N_25220,N_25046);
nor U25939 (N_25939,N_25245,N_25242);
and U25940 (N_25940,N_25085,N_25325);
xnor U25941 (N_25941,N_25152,N_25071);
nor U25942 (N_25942,N_25481,N_25252);
nand U25943 (N_25943,N_25128,N_25364);
or U25944 (N_25944,N_25244,N_25247);
or U25945 (N_25945,N_25438,N_25092);
xor U25946 (N_25946,N_25009,N_25078);
or U25947 (N_25947,N_25359,N_25308);
or U25948 (N_25948,N_25036,N_25093);
or U25949 (N_25949,N_25067,N_25340);
and U25950 (N_25950,N_25234,N_25117);
and U25951 (N_25951,N_25196,N_25380);
nand U25952 (N_25952,N_25462,N_25495);
nand U25953 (N_25953,N_25419,N_25308);
and U25954 (N_25954,N_25119,N_25067);
nand U25955 (N_25955,N_25011,N_25391);
nand U25956 (N_25956,N_25205,N_25250);
nor U25957 (N_25957,N_25063,N_25322);
or U25958 (N_25958,N_25029,N_25018);
nor U25959 (N_25959,N_25029,N_25167);
nand U25960 (N_25960,N_25271,N_25240);
xnor U25961 (N_25961,N_25468,N_25165);
nor U25962 (N_25962,N_25463,N_25093);
xor U25963 (N_25963,N_25041,N_25433);
nand U25964 (N_25964,N_25177,N_25148);
nand U25965 (N_25965,N_25393,N_25492);
and U25966 (N_25966,N_25440,N_25313);
and U25967 (N_25967,N_25474,N_25195);
xnor U25968 (N_25968,N_25246,N_25415);
nor U25969 (N_25969,N_25000,N_25155);
nor U25970 (N_25970,N_25314,N_25394);
and U25971 (N_25971,N_25333,N_25290);
nand U25972 (N_25972,N_25314,N_25007);
and U25973 (N_25973,N_25215,N_25283);
and U25974 (N_25974,N_25347,N_25081);
or U25975 (N_25975,N_25437,N_25234);
nor U25976 (N_25976,N_25085,N_25329);
nand U25977 (N_25977,N_25044,N_25035);
nand U25978 (N_25978,N_25350,N_25454);
nand U25979 (N_25979,N_25241,N_25376);
xor U25980 (N_25980,N_25214,N_25464);
nor U25981 (N_25981,N_25128,N_25084);
nor U25982 (N_25982,N_25071,N_25240);
and U25983 (N_25983,N_25163,N_25018);
nand U25984 (N_25984,N_25425,N_25240);
nor U25985 (N_25985,N_25277,N_25132);
xnor U25986 (N_25986,N_25082,N_25303);
nor U25987 (N_25987,N_25443,N_25261);
nor U25988 (N_25988,N_25084,N_25133);
nor U25989 (N_25989,N_25351,N_25410);
and U25990 (N_25990,N_25282,N_25074);
xor U25991 (N_25991,N_25487,N_25330);
and U25992 (N_25992,N_25242,N_25263);
and U25993 (N_25993,N_25484,N_25058);
or U25994 (N_25994,N_25080,N_25095);
nand U25995 (N_25995,N_25341,N_25145);
nand U25996 (N_25996,N_25014,N_25098);
and U25997 (N_25997,N_25235,N_25327);
or U25998 (N_25998,N_25480,N_25453);
and U25999 (N_25999,N_25146,N_25207);
and U26000 (N_26000,N_25577,N_25642);
and U26001 (N_26001,N_25819,N_25894);
xor U26002 (N_26002,N_25922,N_25941);
nand U26003 (N_26003,N_25571,N_25964);
xor U26004 (N_26004,N_25679,N_25666);
and U26005 (N_26005,N_25982,N_25880);
and U26006 (N_26006,N_25847,N_25920);
nor U26007 (N_26007,N_25669,N_25948);
nand U26008 (N_26008,N_25971,N_25755);
xor U26009 (N_26009,N_25912,N_25639);
xor U26010 (N_26010,N_25973,N_25520);
nand U26011 (N_26011,N_25717,N_25711);
nor U26012 (N_26012,N_25690,N_25745);
and U26013 (N_26013,N_25836,N_25828);
and U26014 (N_26014,N_25817,N_25584);
nand U26015 (N_26015,N_25528,N_25953);
xnor U26016 (N_26016,N_25968,N_25879);
nor U26017 (N_26017,N_25565,N_25995);
or U26018 (N_26018,N_25949,N_25574);
nand U26019 (N_26019,N_25709,N_25606);
and U26020 (N_26020,N_25849,N_25903);
nor U26021 (N_26021,N_25857,N_25511);
nand U26022 (N_26022,N_25805,N_25656);
or U26023 (N_26023,N_25659,N_25604);
and U26024 (N_26024,N_25631,N_25594);
xor U26025 (N_26025,N_25815,N_25811);
xor U26026 (N_26026,N_25977,N_25750);
xnor U26027 (N_26027,N_25535,N_25615);
and U26028 (N_26028,N_25617,N_25713);
xor U26029 (N_26029,N_25766,N_25914);
nor U26030 (N_26030,N_25944,N_25579);
and U26031 (N_26031,N_25911,N_25865);
xor U26032 (N_26032,N_25600,N_25583);
and U26033 (N_26033,N_25746,N_25887);
nand U26034 (N_26034,N_25681,N_25599);
nand U26035 (N_26035,N_25800,N_25969);
or U26036 (N_26036,N_25798,N_25785);
and U26037 (N_26037,N_25705,N_25742);
xnor U26038 (N_26038,N_25706,N_25649);
or U26039 (N_26039,N_25844,N_25657);
xnor U26040 (N_26040,N_25626,N_25931);
xnor U26041 (N_26041,N_25508,N_25622);
nand U26042 (N_26042,N_25648,N_25881);
or U26043 (N_26043,N_25760,N_25651);
or U26044 (N_26044,N_25667,N_25888);
and U26045 (N_26045,N_25719,N_25981);
nor U26046 (N_26046,N_25856,N_25509);
xnor U26047 (N_26047,N_25588,N_25562);
nand U26048 (N_26048,N_25616,N_25807);
nand U26049 (N_26049,N_25665,N_25989);
or U26050 (N_26050,N_25947,N_25915);
and U26051 (N_26051,N_25878,N_25591);
nor U26052 (N_26052,N_25547,N_25826);
or U26053 (N_26053,N_25543,N_25806);
nand U26054 (N_26054,N_25563,N_25897);
and U26055 (N_26055,N_25741,N_25675);
xor U26056 (N_26056,N_25647,N_25824);
nor U26057 (N_26057,N_25635,N_25998);
and U26058 (N_26058,N_25768,N_25788);
xor U26059 (N_26059,N_25598,N_25646);
xnor U26060 (N_26060,N_25929,N_25852);
or U26061 (N_26061,N_25814,N_25875);
xnor U26062 (N_26062,N_25960,N_25688);
or U26063 (N_26063,N_25792,N_25560);
nor U26064 (N_26064,N_25994,N_25672);
nor U26065 (N_26065,N_25595,N_25862);
and U26066 (N_26066,N_25634,N_25506);
nor U26067 (N_26067,N_25654,N_25553);
nand U26068 (N_26068,N_25812,N_25791);
or U26069 (N_26069,N_25658,N_25939);
or U26070 (N_26070,N_25629,N_25951);
or U26071 (N_26071,N_25582,N_25820);
xnor U26072 (N_26072,N_25728,N_25702);
nand U26073 (N_26073,N_25533,N_25794);
and U26074 (N_26074,N_25732,N_25809);
nand U26075 (N_26075,N_25696,N_25924);
nand U26076 (N_26076,N_25692,N_25896);
or U26077 (N_26077,N_25943,N_25796);
xor U26078 (N_26078,N_25945,N_25860);
nand U26079 (N_26079,N_25925,N_25933);
or U26080 (N_26080,N_25913,N_25942);
xnor U26081 (N_26081,N_25540,N_25715);
or U26082 (N_26082,N_25641,N_25673);
nor U26083 (N_26083,N_25686,N_25593);
and U26084 (N_26084,N_25883,N_25640);
or U26085 (N_26085,N_25627,N_25858);
and U26086 (N_26086,N_25778,N_25633);
nand U26087 (N_26087,N_25567,N_25992);
or U26088 (N_26088,N_25988,N_25611);
nand U26089 (N_26089,N_25699,N_25714);
and U26090 (N_26090,N_25930,N_25892);
nand U26091 (N_26091,N_25572,N_25843);
and U26092 (N_26092,N_25643,N_25740);
xor U26093 (N_26093,N_25605,N_25851);
nor U26094 (N_26094,N_25570,N_25764);
nand U26095 (N_26095,N_25845,N_25561);
nand U26096 (N_26096,N_25674,N_25730);
and U26097 (N_26097,N_25687,N_25777);
and U26098 (N_26098,N_25813,N_25661);
and U26099 (N_26099,N_25774,N_25697);
xnor U26100 (N_26100,N_25979,N_25756);
nand U26101 (N_26101,N_25884,N_25795);
xor U26102 (N_26102,N_25905,N_25564);
nand U26103 (N_26103,N_25872,N_25590);
and U26104 (N_26104,N_25923,N_25628);
and U26105 (N_26105,N_25581,N_25753);
nor U26106 (N_26106,N_25996,N_25921);
or U26107 (N_26107,N_25762,N_25891);
and U26108 (N_26108,N_25952,N_25830);
and U26109 (N_26109,N_25662,N_25551);
xor U26110 (N_26110,N_25818,N_25735);
xor U26111 (N_26111,N_25899,N_25799);
nand U26112 (N_26112,N_25636,N_25703);
and U26113 (N_26113,N_25737,N_25691);
xor U26114 (N_26114,N_25693,N_25603);
nor U26115 (N_26115,N_25816,N_25609);
nand U26116 (N_26116,N_25576,N_25502);
or U26117 (N_26117,N_25985,N_25873);
nor U26118 (N_26118,N_25866,N_25840);
nand U26119 (N_26119,N_25548,N_25987);
xnor U26120 (N_26120,N_25909,N_25829);
nor U26121 (N_26121,N_25644,N_25682);
nor U26122 (N_26122,N_25664,N_25578);
xor U26123 (N_26123,N_25680,N_25573);
nor U26124 (N_26124,N_25904,N_25505);
xor U26125 (N_26125,N_25868,N_25918);
nor U26126 (N_26126,N_25784,N_25864);
nor U26127 (N_26127,N_25550,N_25575);
nand U26128 (N_26128,N_25779,N_25676);
nand U26129 (N_26129,N_25978,N_25838);
and U26130 (N_26130,N_25630,N_25723);
and U26131 (N_26131,N_25650,N_25527);
or U26132 (N_26132,N_25712,N_25835);
and U26133 (N_26133,N_25801,N_25965);
and U26134 (N_26134,N_25698,N_25782);
or U26135 (N_26135,N_25776,N_25504);
or U26136 (N_26136,N_25513,N_25514);
nor U26137 (N_26137,N_25769,N_25708);
or U26138 (N_26138,N_25739,N_25957);
nor U26139 (N_26139,N_25962,N_25638);
or U26140 (N_26140,N_25602,N_25773);
and U26141 (N_26141,N_25793,N_25542);
nor U26142 (N_26142,N_25585,N_25889);
nand U26143 (N_26143,N_25910,N_25874);
and U26144 (N_26144,N_25775,N_25991);
nand U26145 (N_26145,N_25652,N_25521);
or U26146 (N_26146,N_25980,N_25932);
and U26147 (N_26147,N_25526,N_25855);
xnor U26148 (N_26148,N_25751,N_25767);
xor U26149 (N_26149,N_25954,N_25886);
nor U26150 (N_26150,N_25823,N_25902);
nand U26151 (N_26151,N_25545,N_25592);
xnor U26152 (N_26152,N_25853,N_25919);
or U26153 (N_26153,N_25736,N_25601);
nand U26154 (N_26154,N_25790,N_25938);
and U26155 (N_26155,N_25976,N_25833);
nand U26156 (N_26156,N_25786,N_25937);
xor U26157 (N_26157,N_25958,N_25695);
nor U26158 (N_26158,N_25519,N_25621);
nand U26159 (N_26159,N_25901,N_25770);
xnor U26160 (N_26160,N_25780,N_25534);
nand U26161 (N_26161,N_25710,N_25848);
nor U26162 (N_26162,N_25789,N_25597);
xnor U26163 (N_26163,N_25733,N_25803);
and U26164 (N_26164,N_25907,N_25832);
and U26165 (N_26165,N_25936,N_25683);
xor U26166 (N_26166,N_25906,N_25761);
or U26167 (N_26167,N_25677,N_25678);
and U26168 (N_26168,N_25757,N_25694);
or U26169 (N_26169,N_25983,N_25546);
or U26170 (N_26170,N_25926,N_25701);
nand U26171 (N_26171,N_25620,N_25895);
and U26172 (N_26172,N_25744,N_25765);
nand U26173 (N_26173,N_25810,N_25787);
xnor U26174 (N_26174,N_25781,N_25890);
nor U26175 (N_26175,N_25607,N_25928);
and U26176 (N_26176,N_25975,N_25722);
nand U26177 (N_26177,N_25934,N_25625);
nor U26178 (N_26178,N_25552,N_25518);
nor U26179 (N_26179,N_25839,N_25935);
nor U26180 (N_26180,N_25908,N_25608);
or U26181 (N_26181,N_25725,N_25716);
xor U26182 (N_26182,N_25704,N_25808);
and U26183 (N_26183,N_25993,N_25729);
or U26184 (N_26184,N_25821,N_25645);
nand U26185 (N_26185,N_25893,N_25556);
nand U26186 (N_26186,N_25940,N_25731);
nor U26187 (N_26187,N_25950,N_25885);
nand U26188 (N_26188,N_25772,N_25738);
and U26189 (N_26189,N_25869,N_25963);
nand U26190 (N_26190,N_25580,N_25589);
or U26191 (N_26191,N_25537,N_25822);
and U26192 (N_26192,N_25530,N_25554);
or U26193 (N_26193,N_25623,N_25999);
xnor U26194 (N_26194,N_25707,N_25524);
or U26195 (N_26195,N_25538,N_25671);
and U26196 (N_26196,N_25837,N_25917);
xor U26197 (N_26197,N_25846,N_25670);
or U26198 (N_26198,N_25689,N_25825);
xnor U26199 (N_26199,N_25668,N_25586);
xor U26200 (N_26200,N_25900,N_25539);
or U26201 (N_26201,N_25967,N_25587);
or U26202 (N_26202,N_25804,N_25842);
xnor U26203 (N_26203,N_25566,N_25632);
xor U26204 (N_26204,N_25700,N_25559);
or U26205 (N_26205,N_25959,N_25684);
xor U26206 (N_26206,N_25834,N_25850);
nand U26207 (N_26207,N_25758,N_25618);
or U26208 (N_26208,N_25541,N_25759);
nor U26209 (N_26209,N_25596,N_25763);
nor U26210 (N_26210,N_25721,N_25997);
xnor U26211 (N_26211,N_25984,N_25624);
xor U26212 (N_26212,N_25685,N_25557);
nor U26213 (N_26213,N_25720,N_25536);
nor U26214 (N_26214,N_25529,N_25507);
nor U26215 (N_26215,N_25544,N_25863);
or U26216 (N_26216,N_25749,N_25955);
and U26217 (N_26217,N_25516,N_25966);
and U26218 (N_26218,N_25771,N_25990);
and U26219 (N_26219,N_25802,N_25956);
nand U26220 (N_26220,N_25523,N_25974);
and U26221 (N_26221,N_25946,N_25653);
xor U26222 (N_26222,N_25517,N_25501);
xor U26223 (N_26223,N_25827,N_25568);
and U26224 (N_26224,N_25916,N_25871);
and U26225 (N_26225,N_25726,N_25512);
xor U26226 (N_26226,N_25870,N_25797);
xnor U26227 (N_26227,N_25510,N_25754);
nor U26228 (N_26228,N_25558,N_25748);
or U26229 (N_26229,N_25531,N_25555);
xor U26230 (N_26230,N_25532,N_25613);
or U26231 (N_26231,N_25637,N_25663);
and U26232 (N_26232,N_25841,N_25747);
and U26233 (N_26233,N_25970,N_25861);
xor U26234 (N_26234,N_25500,N_25660);
nor U26235 (N_26235,N_25503,N_25752);
xor U26236 (N_26236,N_25718,N_25734);
and U26237 (N_26237,N_25867,N_25783);
nand U26238 (N_26238,N_25727,N_25961);
nand U26239 (N_26239,N_25882,N_25877);
nand U26240 (N_26240,N_25724,N_25898);
or U26241 (N_26241,N_25612,N_25522);
and U26242 (N_26242,N_25876,N_25614);
nor U26243 (N_26243,N_25610,N_25569);
xnor U26244 (N_26244,N_25986,N_25549);
nor U26245 (N_26245,N_25515,N_25859);
xnor U26246 (N_26246,N_25972,N_25831);
xnor U26247 (N_26247,N_25619,N_25743);
xor U26248 (N_26248,N_25927,N_25525);
nor U26249 (N_26249,N_25854,N_25655);
xor U26250 (N_26250,N_25643,N_25663);
and U26251 (N_26251,N_25532,N_25542);
nand U26252 (N_26252,N_25634,N_25765);
nand U26253 (N_26253,N_25633,N_25528);
nand U26254 (N_26254,N_25514,N_25996);
and U26255 (N_26255,N_25588,N_25658);
xor U26256 (N_26256,N_25790,N_25606);
xor U26257 (N_26257,N_25854,N_25744);
xnor U26258 (N_26258,N_25718,N_25842);
nor U26259 (N_26259,N_25879,N_25747);
and U26260 (N_26260,N_25790,N_25691);
xnor U26261 (N_26261,N_25962,N_25791);
nand U26262 (N_26262,N_25769,N_25983);
xnor U26263 (N_26263,N_25733,N_25736);
or U26264 (N_26264,N_25664,N_25731);
or U26265 (N_26265,N_25686,N_25513);
xnor U26266 (N_26266,N_25780,N_25872);
nor U26267 (N_26267,N_25692,N_25819);
nor U26268 (N_26268,N_25688,N_25797);
xnor U26269 (N_26269,N_25530,N_25754);
and U26270 (N_26270,N_25522,N_25802);
or U26271 (N_26271,N_25811,N_25832);
and U26272 (N_26272,N_25757,N_25529);
or U26273 (N_26273,N_25610,N_25527);
and U26274 (N_26274,N_25635,N_25700);
or U26275 (N_26275,N_25783,N_25660);
xnor U26276 (N_26276,N_25951,N_25841);
nand U26277 (N_26277,N_25934,N_25703);
xor U26278 (N_26278,N_25556,N_25774);
or U26279 (N_26279,N_25567,N_25769);
nand U26280 (N_26280,N_25868,N_25849);
xor U26281 (N_26281,N_25821,N_25874);
or U26282 (N_26282,N_25898,N_25877);
xnor U26283 (N_26283,N_25894,N_25785);
nand U26284 (N_26284,N_25760,N_25933);
nand U26285 (N_26285,N_25666,N_25526);
nand U26286 (N_26286,N_25766,N_25572);
and U26287 (N_26287,N_25779,N_25791);
xor U26288 (N_26288,N_25788,N_25705);
and U26289 (N_26289,N_25716,N_25794);
nor U26290 (N_26290,N_25975,N_25618);
xor U26291 (N_26291,N_25910,N_25649);
nor U26292 (N_26292,N_25699,N_25842);
nand U26293 (N_26293,N_25887,N_25586);
xor U26294 (N_26294,N_25525,N_25737);
xor U26295 (N_26295,N_25594,N_25625);
nor U26296 (N_26296,N_25597,N_25740);
and U26297 (N_26297,N_25512,N_25861);
and U26298 (N_26298,N_25686,N_25737);
nor U26299 (N_26299,N_25785,N_25636);
nor U26300 (N_26300,N_25530,N_25948);
xor U26301 (N_26301,N_25699,N_25986);
xor U26302 (N_26302,N_25636,N_25782);
and U26303 (N_26303,N_25558,N_25717);
nor U26304 (N_26304,N_25955,N_25615);
nand U26305 (N_26305,N_25900,N_25806);
xnor U26306 (N_26306,N_25527,N_25829);
nand U26307 (N_26307,N_25528,N_25727);
or U26308 (N_26308,N_25712,N_25758);
xor U26309 (N_26309,N_25922,N_25973);
nor U26310 (N_26310,N_25995,N_25527);
and U26311 (N_26311,N_25948,N_25684);
xnor U26312 (N_26312,N_25635,N_25935);
nand U26313 (N_26313,N_25612,N_25549);
and U26314 (N_26314,N_25923,N_25921);
or U26315 (N_26315,N_25786,N_25854);
nor U26316 (N_26316,N_25941,N_25547);
nand U26317 (N_26317,N_25861,N_25966);
xor U26318 (N_26318,N_25553,N_25528);
nand U26319 (N_26319,N_25606,N_25690);
or U26320 (N_26320,N_25789,N_25996);
xnor U26321 (N_26321,N_25639,N_25979);
xor U26322 (N_26322,N_25528,N_25524);
nor U26323 (N_26323,N_25614,N_25924);
or U26324 (N_26324,N_25821,N_25891);
xor U26325 (N_26325,N_25713,N_25583);
xnor U26326 (N_26326,N_25644,N_25697);
nor U26327 (N_26327,N_25502,N_25788);
nor U26328 (N_26328,N_25930,N_25572);
nand U26329 (N_26329,N_25711,N_25628);
nor U26330 (N_26330,N_25852,N_25898);
xnor U26331 (N_26331,N_25881,N_25617);
nor U26332 (N_26332,N_25654,N_25661);
nor U26333 (N_26333,N_25949,N_25894);
xnor U26334 (N_26334,N_25656,N_25885);
or U26335 (N_26335,N_25821,N_25667);
xor U26336 (N_26336,N_25594,N_25884);
nand U26337 (N_26337,N_25743,N_25795);
nand U26338 (N_26338,N_25613,N_25985);
xor U26339 (N_26339,N_25810,N_25790);
nor U26340 (N_26340,N_25703,N_25766);
or U26341 (N_26341,N_25678,N_25940);
nand U26342 (N_26342,N_25676,N_25904);
xor U26343 (N_26343,N_25649,N_25970);
xor U26344 (N_26344,N_25687,N_25957);
and U26345 (N_26345,N_25773,N_25617);
or U26346 (N_26346,N_25514,N_25948);
nand U26347 (N_26347,N_25752,N_25685);
and U26348 (N_26348,N_25777,N_25813);
or U26349 (N_26349,N_25813,N_25770);
nand U26350 (N_26350,N_25767,N_25523);
or U26351 (N_26351,N_25555,N_25784);
xor U26352 (N_26352,N_25873,N_25738);
nor U26353 (N_26353,N_25857,N_25730);
nand U26354 (N_26354,N_25548,N_25742);
and U26355 (N_26355,N_25930,N_25964);
xnor U26356 (N_26356,N_25786,N_25808);
nor U26357 (N_26357,N_25765,N_25762);
nor U26358 (N_26358,N_25662,N_25866);
nor U26359 (N_26359,N_25835,N_25703);
xor U26360 (N_26360,N_25764,N_25559);
xor U26361 (N_26361,N_25571,N_25788);
nand U26362 (N_26362,N_25834,N_25526);
or U26363 (N_26363,N_25645,N_25598);
nor U26364 (N_26364,N_25834,N_25862);
nor U26365 (N_26365,N_25810,N_25770);
nand U26366 (N_26366,N_25720,N_25962);
or U26367 (N_26367,N_25557,N_25673);
nand U26368 (N_26368,N_25852,N_25850);
nand U26369 (N_26369,N_25525,N_25580);
or U26370 (N_26370,N_25766,N_25540);
nor U26371 (N_26371,N_25880,N_25858);
and U26372 (N_26372,N_25895,N_25859);
xnor U26373 (N_26373,N_25734,N_25737);
nor U26374 (N_26374,N_25675,N_25673);
nor U26375 (N_26375,N_25900,N_25580);
or U26376 (N_26376,N_25943,N_25615);
or U26377 (N_26377,N_25914,N_25925);
nor U26378 (N_26378,N_25899,N_25693);
nor U26379 (N_26379,N_25770,N_25750);
or U26380 (N_26380,N_25959,N_25610);
nand U26381 (N_26381,N_25655,N_25730);
xor U26382 (N_26382,N_25686,N_25747);
xor U26383 (N_26383,N_25873,N_25932);
nor U26384 (N_26384,N_25660,N_25708);
and U26385 (N_26385,N_25742,N_25972);
or U26386 (N_26386,N_25751,N_25829);
xor U26387 (N_26387,N_25573,N_25647);
or U26388 (N_26388,N_25598,N_25997);
nand U26389 (N_26389,N_25741,N_25824);
xor U26390 (N_26390,N_25628,N_25610);
nand U26391 (N_26391,N_25956,N_25662);
and U26392 (N_26392,N_25841,N_25511);
and U26393 (N_26393,N_25845,N_25804);
or U26394 (N_26394,N_25581,N_25999);
and U26395 (N_26395,N_25819,N_25768);
and U26396 (N_26396,N_25893,N_25937);
nand U26397 (N_26397,N_25852,N_25882);
or U26398 (N_26398,N_25733,N_25524);
nand U26399 (N_26399,N_25737,N_25585);
nor U26400 (N_26400,N_25849,N_25807);
xnor U26401 (N_26401,N_25802,N_25691);
and U26402 (N_26402,N_25938,N_25629);
nor U26403 (N_26403,N_25782,N_25718);
nor U26404 (N_26404,N_25900,N_25688);
xor U26405 (N_26405,N_25787,N_25822);
or U26406 (N_26406,N_25969,N_25839);
or U26407 (N_26407,N_25979,N_25635);
nand U26408 (N_26408,N_25550,N_25697);
nand U26409 (N_26409,N_25816,N_25560);
or U26410 (N_26410,N_25714,N_25990);
nand U26411 (N_26411,N_25762,N_25632);
nand U26412 (N_26412,N_25548,N_25890);
and U26413 (N_26413,N_25755,N_25934);
nand U26414 (N_26414,N_25675,N_25541);
nor U26415 (N_26415,N_25787,N_25832);
and U26416 (N_26416,N_25732,N_25607);
or U26417 (N_26417,N_25623,N_25871);
xnor U26418 (N_26418,N_25626,N_25667);
xnor U26419 (N_26419,N_25832,N_25660);
xor U26420 (N_26420,N_25545,N_25817);
nor U26421 (N_26421,N_25767,N_25595);
xnor U26422 (N_26422,N_25719,N_25980);
and U26423 (N_26423,N_25997,N_25848);
nand U26424 (N_26424,N_25828,N_25941);
and U26425 (N_26425,N_25785,N_25654);
xor U26426 (N_26426,N_25747,N_25702);
nor U26427 (N_26427,N_25855,N_25919);
nand U26428 (N_26428,N_25938,N_25587);
and U26429 (N_26429,N_25556,N_25728);
nor U26430 (N_26430,N_25951,N_25638);
xor U26431 (N_26431,N_25569,N_25787);
or U26432 (N_26432,N_25777,N_25830);
nand U26433 (N_26433,N_25967,N_25841);
xnor U26434 (N_26434,N_25964,N_25514);
xnor U26435 (N_26435,N_25832,N_25586);
nand U26436 (N_26436,N_25905,N_25628);
xnor U26437 (N_26437,N_25510,N_25836);
nand U26438 (N_26438,N_25815,N_25705);
or U26439 (N_26439,N_25532,N_25943);
xor U26440 (N_26440,N_25868,N_25966);
nor U26441 (N_26441,N_25903,N_25675);
xor U26442 (N_26442,N_25889,N_25900);
xnor U26443 (N_26443,N_25591,N_25627);
nand U26444 (N_26444,N_25758,N_25768);
nor U26445 (N_26445,N_25935,N_25594);
nor U26446 (N_26446,N_25969,N_25602);
and U26447 (N_26447,N_25914,N_25813);
xor U26448 (N_26448,N_25882,N_25553);
or U26449 (N_26449,N_25634,N_25931);
xnor U26450 (N_26450,N_25713,N_25644);
xnor U26451 (N_26451,N_25714,N_25787);
and U26452 (N_26452,N_25602,N_25890);
nor U26453 (N_26453,N_25778,N_25729);
nor U26454 (N_26454,N_25559,N_25789);
or U26455 (N_26455,N_25803,N_25504);
xnor U26456 (N_26456,N_25682,N_25766);
and U26457 (N_26457,N_25597,N_25750);
nand U26458 (N_26458,N_25959,N_25576);
or U26459 (N_26459,N_25792,N_25786);
nand U26460 (N_26460,N_25635,N_25865);
and U26461 (N_26461,N_25992,N_25813);
xnor U26462 (N_26462,N_25645,N_25925);
nand U26463 (N_26463,N_25988,N_25922);
nor U26464 (N_26464,N_25903,N_25942);
and U26465 (N_26465,N_25602,N_25639);
xor U26466 (N_26466,N_25678,N_25927);
nand U26467 (N_26467,N_25745,N_25924);
nor U26468 (N_26468,N_25996,N_25738);
or U26469 (N_26469,N_25582,N_25594);
and U26470 (N_26470,N_25928,N_25750);
xnor U26471 (N_26471,N_25884,N_25530);
xnor U26472 (N_26472,N_25835,N_25933);
nor U26473 (N_26473,N_25680,N_25675);
and U26474 (N_26474,N_25684,N_25735);
nor U26475 (N_26475,N_25544,N_25967);
xnor U26476 (N_26476,N_25997,N_25673);
xor U26477 (N_26477,N_25970,N_25574);
and U26478 (N_26478,N_25748,N_25502);
nand U26479 (N_26479,N_25889,N_25814);
nor U26480 (N_26480,N_25816,N_25770);
and U26481 (N_26481,N_25801,N_25701);
xnor U26482 (N_26482,N_25682,N_25994);
nand U26483 (N_26483,N_25989,N_25731);
nand U26484 (N_26484,N_25797,N_25743);
and U26485 (N_26485,N_25807,N_25970);
nand U26486 (N_26486,N_25997,N_25912);
or U26487 (N_26487,N_25901,N_25990);
xor U26488 (N_26488,N_25699,N_25800);
xor U26489 (N_26489,N_25958,N_25572);
xor U26490 (N_26490,N_25967,N_25595);
and U26491 (N_26491,N_25737,N_25913);
and U26492 (N_26492,N_25699,N_25887);
nor U26493 (N_26493,N_25603,N_25668);
nor U26494 (N_26494,N_25946,N_25976);
nor U26495 (N_26495,N_25769,N_25705);
nand U26496 (N_26496,N_25579,N_25864);
or U26497 (N_26497,N_25781,N_25675);
or U26498 (N_26498,N_25810,N_25734);
nor U26499 (N_26499,N_25613,N_25543);
or U26500 (N_26500,N_26041,N_26336);
or U26501 (N_26501,N_26250,N_26039);
nor U26502 (N_26502,N_26284,N_26311);
xor U26503 (N_26503,N_26204,N_26075);
xor U26504 (N_26504,N_26397,N_26053);
xor U26505 (N_26505,N_26224,N_26038);
and U26506 (N_26506,N_26316,N_26168);
nor U26507 (N_26507,N_26062,N_26273);
or U26508 (N_26508,N_26322,N_26127);
xnor U26509 (N_26509,N_26431,N_26118);
nor U26510 (N_26510,N_26134,N_26049);
or U26511 (N_26511,N_26028,N_26324);
xor U26512 (N_26512,N_26415,N_26402);
nand U26513 (N_26513,N_26436,N_26132);
xor U26514 (N_26514,N_26492,N_26223);
nor U26515 (N_26515,N_26111,N_26275);
nand U26516 (N_26516,N_26435,N_26234);
nand U26517 (N_26517,N_26023,N_26044);
and U26518 (N_26518,N_26280,N_26084);
or U26519 (N_26519,N_26155,N_26129);
nand U26520 (N_26520,N_26298,N_26177);
and U26521 (N_26521,N_26115,N_26192);
or U26522 (N_26522,N_26248,N_26110);
or U26523 (N_26523,N_26025,N_26011);
and U26524 (N_26524,N_26088,N_26003);
nor U26525 (N_26525,N_26063,N_26413);
or U26526 (N_26526,N_26007,N_26477);
nand U26527 (N_26527,N_26403,N_26405);
nand U26528 (N_26528,N_26335,N_26164);
xnor U26529 (N_26529,N_26200,N_26065);
and U26530 (N_26530,N_26101,N_26312);
nor U26531 (N_26531,N_26434,N_26462);
and U26532 (N_26532,N_26125,N_26342);
xnor U26533 (N_26533,N_26404,N_26314);
nand U26534 (N_26534,N_26212,N_26352);
or U26535 (N_26535,N_26099,N_26207);
xor U26536 (N_26536,N_26292,N_26407);
nand U26537 (N_26537,N_26203,N_26499);
xor U26538 (N_26538,N_26114,N_26349);
xor U26539 (N_26539,N_26024,N_26343);
nor U26540 (N_26540,N_26429,N_26359);
and U26541 (N_26541,N_26152,N_26108);
nand U26542 (N_26542,N_26165,N_26470);
xnor U26543 (N_26543,N_26411,N_26332);
and U26544 (N_26544,N_26031,N_26387);
nand U26545 (N_26545,N_26082,N_26150);
and U26546 (N_26546,N_26338,N_26458);
nor U26547 (N_26547,N_26206,N_26498);
nor U26548 (N_26548,N_26293,N_26399);
nor U26549 (N_26549,N_26214,N_26201);
nand U26550 (N_26550,N_26267,N_26231);
or U26551 (N_26551,N_26488,N_26469);
nand U26552 (N_26552,N_26090,N_26472);
nor U26553 (N_26553,N_26363,N_26162);
nand U26554 (N_26554,N_26307,N_26466);
nand U26555 (N_26555,N_26457,N_26339);
nor U26556 (N_26556,N_26179,N_26002);
xnor U26557 (N_26557,N_26046,N_26116);
xor U26558 (N_26558,N_26061,N_26442);
nand U26559 (N_26559,N_26306,N_26210);
nand U26560 (N_26560,N_26334,N_26133);
or U26561 (N_26561,N_26083,N_26058);
and U26562 (N_26562,N_26015,N_26167);
or U26563 (N_26563,N_26222,N_26260);
and U26564 (N_26564,N_26193,N_26093);
xnor U26565 (N_26565,N_26493,N_26228);
nor U26566 (N_26566,N_26050,N_26047);
and U26567 (N_26567,N_26253,N_26256);
nand U26568 (N_26568,N_26425,N_26045);
or U26569 (N_26569,N_26030,N_26244);
and U26570 (N_26570,N_26016,N_26019);
xnor U26571 (N_26571,N_26421,N_26227);
xnor U26572 (N_26572,N_26455,N_26364);
nor U26573 (N_26573,N_26296,N_26313);
nand U26574 (N_26574,N_26022,N_26281);
nor U26575 (N_26575,N_26128,N_26422);
and U26576 (N_26576,N_26416,N_26277);
or U26577 (N_26577,N_26361,N_26265);
nor U26578 (N_26578,N_26173,N_26271);
xor U26579 (N_26579,N_26305,N_26219);
or U26580 (N_26580,N_26299,N_26372);
nor U26581 (N_26581,N_26395,N_26189);
or U26582 (N_26582,N_26430,N_26471);
and U26583 (N_26583,N_26018,N_26287);
and U26584 (N_26584,N_26368,N_26444);
or U26585 (N_26585,N_26278,N_26414);
and U26586 (N_26586,N_26027,N_26274);
and U26587 (N_26587,N_26104,N_26072);
xnor U26588 (N_26588,N_26383,N_26329);
nor U26589 (N_26589,N_26318,N_26282);
or U26590 (N_26590,N_26379,N_26406);
and U26591 (N_26591,N_26366,N_26448);
and U26592 (N_26592,N_26000,N_26220);
nor U26593 (N_26593,N_26239,N_26191);
xnor U26594 (N_26594,N_26428,N_26303);
or U26595 (N_26595,N_26170,N_26034);
xnor U26596 (N_26596,N_26350,N_26323);
nand U26597 (N_26597,N_26137,N_26085);
nand U26598 (N_26598,N_26400,N_26198);
nor U26599 (N_26599,N_26057,N_26348);
nand U26600 (N_26600,N_26295,N_26255);
nand U26601 (N_26601,N_26266,N_26480);
and U26602 (N_26602,N_26320,N_26123);
and U26603 (N_26603,N_26355,N_26183);
nor U26604 (N_26604,N_26490,N_26051);
or U26605 (N_26605,N_26396,N_26229);
nand U26606 (N_26606,N_26095,N_26145);
nor U26607 (N_26607,N_26106,N_26308);
xnor U26608 (N_26608,N_26136,N_26241);
xnor U26609 (N_26609,N_26494,N_26094);
nand U26610 (N_26610,N_26008,N_26059);
and U26611 (N_26611,N_26496,N_26365);
nand U26612 (N_26612,N_26432,N_26158);
or U26613 (N_26613,N_26160,N_26393);
nor U26614 (N_26614,N_26197,N_26238);
xor U26615 (N_26615,N_26196,N_26163);
and U26616 (N_26616,N_26237,N_26139);
or U26617 (N_26617,N_26330,N_26454);
nand U26618 (N_26618,N_26412,N_26426);
and U26619 (N_26619,N_26309,N_26463);
or U26620 (N_26620,N_26195,N_26447);
nor U26621 (N_26621,N_26317,N_26438);
and U26622 (N_26622,N_26124,N_26424);
nor U26623 (N_26623,N_26004,N_26186);
nand U26624 (N_26624,N_26122,N_26262);
or U26625 (N_26625,N_26140,N_26087);
nand U26626 (N_26626,N_26378,N_26489);
or U26627 (N_26627,N_26357,N_26091);
nor U26628 (N_26628,N_26290,N_26117);
and U26629 (N_26629,N_26441,N_26473);
nand U26630 (N_26630,N_26240,N_26269);
or U26631 (N_26631,N_26048,N_26138);
nand U26632 (N_26632,N_26130,N_26070);
nor U26633 (N_26633,N_26433,N_26181);
nand U26634 (N_26634,N_26009,N_26279);
and U26635 (N_26635,N_26209,N_26199);
or U26636 (N_26636,N_26386,N_26385);
or U26637 (N_26637,N_26495,N_26076);
or U26638 (N_26638,N_26390,N_26077);
and U26639 (N_26639,N_26325,N_26449);
nor U26640 (N_26640,N_26391,N_26036);
or U26641 (N_26641,N_26235,N_26345);
nand U26642 (N_26642,N_26254,N_26142);
or U26643 (N_26643,N_26474,N_26258);
or U26644 (N_26644,N_26100,N_26144);
xnor U26645 (N_26645,N_26465,N_26467);
or U26646 (N_26646,N_26079,N_26180);
or U26647 (N_26647,N_26109,N_26456);
nor U26648 (N_26648,N_26172,N_26486);
xor U26649 (N_26649,N_26071,N_26182);
or U26650 (N_26650,N_26042,N_26301);
xor U26651 (N_26651,N_26382,N_26013);
xor U26652 (N_26652,N_26190,N_26131);
nand U26653 (N_26653,N_26141,N_26340);
nand U26654 (N_26654,N_26001,N_26178);
nor U26655 (N_26655,N_26147,N_26389);
nand U26656 (N_26656,N_26344,N_26261);
and U26657 (N_26657,N_26326,N_26113);
nand U26658 (N_26658,N_26175,N_26052);
nor U26659 (N_26659,N_26302,N_26020);
xnor U26660 (N_26660,N_26069,N_26242);
xnor U26661 (N_26661,N_26270,N_26394);
xor U26662 (N_26662,N_26217,N_26156);
or U26663 (N_26663,N_26102,N_26373);
and U26664 (N_26664,N_26362,N_26066);
and U26665 (N_26665,N_26054,N_26021);
nor U26666 (N_26666,N_26064,N_26475);
nor U26667 (N_26667,N_26126,N_26353);
and U26668 (N_26668,N_26478,N_26423);
or U26669 (N_26669,N_26371,N_26450);
nand U26670 (N_26670,N_26184,N_26067);
nand U26671 (N_26671,N_26452,N_26010);
xnor U26672 (N_26672,N_26300,N_26263);
and U26673 (N_26673,N_26294,N_26211);
nor U26674 (N_26674,N_26153,N_26377);
xor U26675 (N_26675,N_26376,N_26439);
and U26676 (N_26676,N_26483,N_26208);
xor U26677 (N_26677,N_26367,N_26086);
xnor U26678 (N_26678,N_26297,N_26040);
nor U26679 (N_26679,N_26485,N_26187);
xor U26680 (N_26680,N_26068,N_26257);
and U26681 (N_26681,N_26148,N_26119);
and U26682 (N_26682,N_26374,N_26218);
xor U26683 (N_26683,N_26446,N_26171);
xor U26684 (N_26684,N_26096,N_26327);
xnor U26685 (N_26685,N_26440,N_26460);
nand U26686 (N_26686,N_26249,N_26443);
nand U26687 (N_26687,N_26169,N_26017);
nor U26688 (N_26688,N_26026,N_26328);
and U26689 (N_26689,N_26437,N_26230);
nor U26690 (N_26690,N_26252,N_26286);
or U26691 (N_26691,N_26243,N_26451);
and U26692 (N_26692,N_26259,N_26081);
and U26693 (N_26693,N_26285,N_26321);
and U26694 (N_26694,N_26112,N_26236);
nand U26695 (N_26695,N_26418,N_26232);
nand U26696 (N_26696,N_26103,N_26331);
xor U26697 (N_26697,N_26417,N_26149);
and U26698 (N_26698,N_26157,N_26035);
nor U26699 (N_26699,N_26226,N_26225);
nor U26700 (N_26700,N_26161,N_26484);
nand U26701 (N_26701,N_26121,N_26408);
nor U26702 (N_26702,N_26360,N_26333);
nor U26703 (N_26703,N_26380,N_26098);
xnor U26704 (N_26704,N_26319,N_26151);
xnor U26705 (N_26705,N_26251,N_26388);
and U26706 (N_26706,N_26245,N_26398);
nor U26707 (N_26707,N_26143,N_26176);
and U26708 (N_26708,N_26341,N_26268);
and U26709 (N_26709,N_26105,N_26089);
nor U26710 (N_26710,N_26185,N_26246);
xor U26711 (N_26711,N_26107,N_26351);
and U26712 (N_26712,N_26188,N_26247);
xor U26713 (N_26713,N_26056,N_26445);
xnor U26714 (N_26714,N_26491,N_26487);
or U26715 (N_26715,N_26346,N_26221);
nor U26716 (N_26716,N_26006,N_26005);
and U26717 (N_26717,N_26481,N_26419);
nor U26718 (N_26718,N_26012,N_26356);
xor U26719 (N_26719,N_26154,N_26453);
nor U26720 (N_26720,N_26464,N_26304);
and U26721 (N_26721,N_26120,N_26205);
nand U26722 (N_26722,N_26315,N_26014);
xnor U26723 (N_26723,N_26337,N_26288);
nand U26724 (N_26724,N_26370,N_26055);
and U26725 (N_26725,N_26215,N_26410);
nand U26726 (N_26726,N_26497,N_26078);
and U26727 (N_26727,N_26461,N_26216);
nand U26728 (N_26728,N_26401,N_26092);
and U26729 (N_26729,N_26074,N_26202);
nor U26730 (N_26730,N_26032,N_26384);
xnor U26731 (N_26731,N_26159,N_26381);
nand U26732 (N_26732,N_26043,N_26459);
or U26733 (N_26733,N_26073,N_26420);
nor U26734 (N_26734,N_26479,N_26358);
and U26735 (N_26735,N_26427,N_26310);
nand U26736 (N_26736,N_26264,N_26213);
xnor U26737 (N_26737,N_26135,N_26369);
or U26738 (N_26738,N_26482,N_26409);
or U26739 (N_26739,N_26354,N_26468);
nand U26740 (N_26740,N_26194,N_26272);
and U26741 (N_26741,N_26291,N_26060);
nand U26742 (N_26742,N_26276,N_26392);
nor U26743 (N_26743,N_26146,N_26097);
and U26744 (N_26744,N_26283,N_26033);
nand U26745 (N_26745,N_26375,N_26476);
or U26746 (N_26746,N_26029,N_26166);
nand U26747 (N_26747,N_26174,N_26037);
xor U26748 (N_26748,N_26233,N_26289);
nand U26749 (N_26749,N_26080,N_26347);
xnor U26750 (N_26750,N_26456,N_26107);
nand U26751 (N_26751,N_26231,N_26213);
nor U26752 (N_26752,N_26437,N_26069);
nor U26753 (N_26753,N_26019,N_26360);
nand U26754 (N_26754,N_26025,N_26048);
nand U26755 (N_26755,N_26480,N_26446);
xnor U26756 (N_26756,N_26144,N_26294);
nor U26757 (N_26757,N_26377,N_26276);
nand U26758 (N_26758,N_26108,N_26271);
or U26759 (N_26759,N_26377,N_26233);
xnor U26760 (N_26760,N_26173,N_26355);
or U26761 (N_26761,N_26237,N_26179);
and U26762 (N_26762,N_26259,N_26490);
or U26763 (N_26763,N_26199,N_26344);
xor U26764 (N_26764,N_26311,N_26094);
nand U26765 (N_26765,N_26252,N_26258);
or U26766 (N_26766,N_26399,N_26078);
nor U26767 (N_26767,N_26198,N_26242);
and U26768 (N_26768,N_26214,N_26267);
xor U26769 (N_26769,N_26118,N_26251);
and U26770 (N_26770,N_26289,N_26456);
nand U26771 (N_26771,N_26415,N_26493);
and U26772 (N_26772,N_26156,N_26223);
nand U26773 (N_26773,N_26060,N_26464);
xnor U26774 (N_26774,N_26372,N_26042);
and U26775 (N_26775,N_26328,N_26300);
nand U26776 (N_26776,N_26105,N_26029);
and U26777 (N_26777,N_26247,N_26305);
or U26778 (N_26778,N_26491,N_26007);
nand U26779 (N_26779,N_26006,N_26321);
xor U26780 (N_26780,N_26082,N_26016);
nand U26781 (N_26781,N_26238,N_26245);
xor U26782 (N_26782,N_26192,N_26465);
nand U26783 (N_26783,N_26020,N_26079);
nor U26784 (N_26784,N_26139,N_26034);
nor U26785 (N_26785,N_26436,N_26332);
nor U26786 (N_26786,N_26161,N_26389);
nor U26787 (N_26787,N_26435,N_26233);
nor U26788 (N_26788,N_26444,N_26207);
or U26789 (N_26789,N_26446,N_26002);
and U26790 (N_26790,N_26130,N_26359);
and U26791 (N_26791,N_26497,N_26256);
nand U26792 (N_26792,N_26054,N_26071);
and U26793 (N_26793,N_26225,N_26072);
xnor U26794 (N_26794,N_26104,N_26440);
and U26795 (N_26795,N_26182,N_26369);
nor U26796 (N_26796,N_26010,N_26006);
xor U26797 (N_26797,N_26285,N_26017);
or U26798 (N_26798,N_26005,N_26387);
or U26799 (N_26799,N_26264,N_26063);
and U26800 (N_26800,N_26190,N_26042);
or U26801 (N_26801,N_26438,N_26186);
and U26802 (N_26802,N_26435,N_26157);
or U26803 (N_26803,N_26261,N_26450);
nand U26804 (N_26804,N_26294,N_26354);
nor U26805 (N_26805,N_26369,N_26109);
and U26806 (N_26806,N_26233,N_26057);
nand U26807 (N_26807,N_26057,N_26106);
xnor U26808 (N_26808,N_26051,N_26263);
xor U26809 (N_26809,N_26396,N_26129);
xor U26810 (N_26810,N_26252,N_26294);
and U26811 (N_26811,N_26286,N_26098);
nand U26812 (N_26812,N_26419,N_26115);
nor U26813 (N_26813,N_26257,N_26177);
nor U26814 (N_26814,N_26443,N_26172);
xnor U26815 (N_26815,N_26180,N_26254);
nor U26816 (N_26816,N_26462,N_26246);
and U26817 (N_26817,N_26005,N_26209);
nor U26818 (N_26818,N_26452,N_26092);
or U26819 (N_26819,N_26209,N_26399);
xor U26820 (N_26820,N_26321,N_26061);
and U26821 (N_26821,N_26003,N_26306);
nand U26822 (N_26822,N_26239,N_26177);
and U26823 (N_26823,N_26126,N_26347);
or U26824 (N_26824,N_26155,N_26295);
nand U26825 (N_26825,N_26150,N_26341);
and U26826 (N_26826,N_26098,N_26019);
nor U26827 (N_26827,N_26302,N_26242);
xnor U26828 (N_26828,N_26475,N_26307);
nor U26829 (N_26829,N_26434,N_26231);
or U26830 (N_26830,N_26258,N_26323);
nand U26831 (N_26831,N_26169,N_26016);
nand U26832 (N_26832,N_26433,N_26225);
xnor U26833 (N_26833,N_26466,N_26346);
xor U26834 (N_26834,N_26255,N_26039);
nor U26835 (N_26835,N_26260,N_26221);
and U26836 (N_26836,N_26225,N_26079);
nor U26837 (N_26837,N_26092,N_26431);
xor U26838 (N_26838,N_26344,N_26226);
nand U26839 (N_26839,N_26077,N_26290);
and U26840 (N_26840,N_26172,N_26023);
or U26841 (N_26841,N_26235,N_26254);
or U26842 (N_26842,N_26088,N_26060);
or U26843 (N_26843,N_26062,N_26154);
and U26844 (N_26844,N_26242,N_26478);
nor U26845 (N_26845,N_26089,N_26294);
nor U26846 (N_26846,N_26389,N_26204);
nor U26847 (N_26847,N_26300,N_26481);
nand U26848 (N_26848,N_26389,N_26495);
nor U26849 (N_26849,N_26429,N_26393);
nor U26850 (N_26850,N_26077,N_26021);
xor U26851 (N_26851,N_26213,N_26314);
xor U26852 (N_26852,N_26197,N_26147);
nand U26853 (N_26853,N_26417,N_26327);
or U26854 (N_26854,N_26130,N_26223);
nor U26855 (N_26855,N_26478,N_26025);
and U26856 (N_26856,N_26489,N_26328);
and U26857 (N_26857,N_26474,N_26058);
and U26858 (N_26858,N_26250,N_26465);
nand U26859 (N_26859,N_26153,N_26417);
nor U26860 (N_26860,N_26299,N_26275);
xnor U26861 (N_26861,N_26217,N_26461);
nor U26862 (N_26862,N_26165,N_26406);
or U26863 (N_26863,N_26255,N_26081);
xor U26864 (N_26864,N_26137,N_26405);
and U26865 (N_26865,N_26322,N_26473);
nand U26866 (N_26866,N_26095,N_26039);
or U26867 (N_26867,N_26072,N_26486);
xnor U26868 (N_26868,N_26131,N_26223);
nor U26869 (N_26869,N_26148,N_26410);
or U26870 (N_26870,N_26049,N_26390);
or U26871 (N_26871,N_26254,N_26489);
and U26872 (N_26872,N_26198,N_26356);
nand U26873 (N_26873,N_26153,N_26176);
nand U26874 (N_26874,N_26114,N_26111);
nor U26875 (N_26875,N_26115,N_26276);
or U26876 (N_26876,N_26203,N_26374);
xor U26877 (N_26877,N_26336,N_26124);
nand U26878 (N_26878,N_26136,N_26314);
and U26879 (N_26879,N_26452,N_26217);
or U26880 (N_26880,N_26188,N_26200);
nor U26881 (N_26881,N_26355,N_26440);
xnor U26882 (N_26882,N_26458,N_26481);
xnor U26883 (N_26883,N_26265,N_26302);
or U26884 (N_26884,N_26491,N_26153);
or U26885 (N_26885,N_26294,N_26371);
or U26886 (N_26886,N_26184,N_26476);
nand U26887 (N_26887,N_26216,N_26487);
nor U26888 (N_26888,N_26051,N_26175);
and U26889 (N_26889,N_26428,N_26393);
nand U26890 (N_26890,N_26054,N_26441);
and U26891 (N_26891,N_26361,N_26104);
nor U26892 (N_26892,N_26245,N_26369);
nand U26893 (N_26893,N_26153,N_26361);
xor U26894 (N_26894,N_26039,N_26197);
or U26895 (N_26895,N_26400,N_26172);
nor U26896 (N_26896,N_26050,N_26098);
and U26897 (N_26897,N_26466,N_26138);
or U26898 (N_26898,N_26344,N_26286);
or U26899 (N_26899,N_26396,N_26476);
or U26900 (N_26900,N_26239,N_26089);
and U26901 (N_26901,N_26154,N_26145);
and U26902 (N_26902,N_26423,N_26310);
nor U26903 (N_26903,N_26460,N_26341);
or U26904 (N_26904,N_26034,N_26053);
and U26905 (N_26905,N_26303,N_26457);
nand U26906 (N_26906,N_26201,N_26179);
xor U26907 (N_26907,N_26378,N_26483);
and U26908 (N_26908,N_26466,N_26208);
nand U26909 (N_26909,N_26042,N_26427);
nand U26910 (N_26910,N_26223,N_26277);
nor U26911 (N_26911,N_26333,N_26316);
nor U26912 (N_26912,N_26444,N_26131);
or U26913 (N_26913,N_26051,N_26378);
xnor U26914 (N_26914,N_26345,N_26267);
nor U26915 (N_26915,N_26175,N_26497);
xor U26916 (N_26916,N_26414,N_26025);
nor U26917 (N_26917,N_26246,N_26391);
xor U26918 (N_26918,N_26038,N_26487);
xor U26919 (N_26919,N_26086,N_26018);
nand U26920 (N_26920,N_26489,N_26419);
xnor U26921 (N_26921,N_26046,N_26394);
nor U26922 (N_26922,N_26311,N_26151);
or U26923 (N_26923,N_26378,N_26267);
nor U26924 (N_26924,N_26198,N_26071);
and U26925 (N_26925,N_26195,N_26024);
and U26926 (N_26926,N_26204,N_26404);
or U26927 (N_26927,N_26135,N_26421);
and U26928 (N_26928,N_26477,N_26205);
xor U26929 (N_26929,N_26289,N_26466);
nand U26930 (N_26930,N_26203,N_26063);
or U26931 (N_26931,N_26291,N_26394);
or U26932 (N_26932,N_26062,N_26089);
or U26933 (N_26933,N_26260,N_26212);
xnor U26934 (N_26934,N_26432,N_26111);
nand U26935 (N_26935,N_26336,N_26146);
xor U26936 (N_26936,N_26147,N_26367);
and U26937 (N_26937,N_26214,N_26088);
or U26938 (N_26938,N_26031,N_26448);
xor U26939 (N_26939,N_26036,N_26368);
nor U26940 (N_26940,N_26480,N_26192);
nor U26941 (N_26941,N_26379,N_26089);
or U26942 (N_26942,N_26221,N_26427);
nor U26943 (N_26943,N_26391,N_26255);
nor U26944 (N_26944,N_26422,N_26486);
and U26945 (N_26945,N_26077,N_26215);
or U26946 (N_26946,N_26380,N_26434);
nand U26947 (N_26947,N_26467,N_26477);
or U26948 (N_26948,N_26110,N_26146);
xor U26949 (N_26949,N_26369,N_26442);
xnor U26950 (N_26950,N_26261,N_26386);
nand U26951 (N_26951,N_26200,N_26408);
or U26952 (N_26952,N_26051,N_26317);
or U26953 (N_26953,N_26186,N_26071);
nor U26954 (N_26954,N_26138,N_26136);
or U26955 (N_26955,N_26449,N_26006);
nand U26956 (N_26956,N_26115,N_26443);
nand U26957 (N_26957,N_26496,N_26218);
nor U26958 (N_26958,N_26009,N_26310);
and U26959 (N_26959,N_26092,N_26176);
nand U26960 (N_26960,N_26416,N_26419);
nor U26961 (N_26961,N_26370,N_26033);
and U26962 (N_26962,N_26068,N_26381);
xnor U26963 (N_26963,N_26082,N_26201);
and U26964 (N_26964,N_26211,N_26370);
nand U26965 (N_26965,N_26022,N_26408);
xnor U26966 (N_26966,N_26454,N_26233);
and U26967 (N_26967,N_26423,N_26196);
nor U26968 (N_26968,N_26337,N_26442);
nand U26969 (N_26969,N_26494,N_26091);
xnor U26970 (N_26970,N_26240,N_26394);
and U26971 (N_26971,N_26136,N_26311);
and U26972 (N_26972,N_26139,N_26149);
or U26973 (N_26973,N_26492,N_26378);
xor U26974 (N_26974,N_26138,N_26441);
nor U26975 (N_26975,N_26373,N_26370);
and U26976 (N_26976,N_26372,N_26252);
and U26977 (N_26977,N_26339,N_26493);
or U26978 (N_26978,N_26492,N_26386);
or U26979 (N_26979,N_26306,N_26266);
nand U26980 (N_26980,N_26113,N_26341);
and U26981 (N_26981,N_26420,N_26297);
nor U26982 (N_26982,N_26188,N_26420);
or U26983 (N_26983,N_26348,N_26295);
nor U26984 (N_26984,N_26102,N_26452);
nand U26985 (N_26985,N_26467,N_26325);
nand U26986 (N_26986,N_26200,N_26403);
xor U26987 (N_26987,N_26460,N_26375);
or U26988 (N_26988,N_26135,N_26328);
nor U26989 (N_26989,N_26003,N_26008);
and U26990 (N_26990,N_26386,N_26177);
or U26991 (N_26991,N_26439,N_26227);
or U26992 (N_26992,N_26485,N_26118);
nor U26993 (N_26993,N_26049,N_26394);
nand U26994 (N_26994,N_26219,N_26314);
or U26995 (N_26995,N_26258,N_26392);
nor U26996 (N_26996,N_26291,N_26346);
or U26997 (N_26997,N_26497,N_26225);
nand U26998 (N_26998,N_26297,N_26097);
nor U26999 (N_26999,N_26377,N_26092);
xnor U27000 (N_27000,N_26920,N_26749);
and U27001 (N_27001,N_26794,N_26868);
xor U27002 (N_27002,N_26514,N_26585);
nand U27003 (N_27003,N_26574,N_26958);
and U27004 (N_27004,N_26990,N_26744);
or U27005 (N_27005,N_26583,N_26881);
nor U27006 (N_27006,N_26850,N_26548);
nor U27007 (N_27007,N_26921,N_26773);
and U27008 (N_27008,N_26849,N_26537);
or U27009 (N_27009,N_26598,N_26538);
nand U27010 (N_27010,N_26852,N_26597);
and U27011 (N_27011,N_26542,N_26714);
nor U27012 (N_27012,N_26835,N_26747);
nand U27013 (N_27013,N_26946,N_26563);
or U27014 (N_27014,N_26648,N_26615);
or U27015 (N_27015,N_26971,N_26909);
nor U27016 (N_27016,N_26669,N_26596);
or U27017 (N_27017,N_26664,N_26690);
nor U27018 (N_27018,N_26549,N_26717);
nor U27019 (N_27019,N_26892,N_26612);
and U27020 (N_27020,N_26878,N_26523);
and U27021 (N_27021,N_26711,N_26674);
or U27022 (N_27022,N_26704,N_26680);
nand U27023 (N_27023,N_26983,N_26931);
nand U27024 (N_27024,N_26634,N_26817);
and U27025 (N_27025,N_26684,N_26837);
and U27026 (N_27026,N_26888,N_26687);
nor U27027 (N_27027,N_26956,N_26544);
and U27028 (N_27028,N_26898,N_26871);
nor U27029 (N_27029,N_26936,N_26724);
and U27030 (N_27030,N_26599,N_26654);
or U27031 (N_27031,N_26814,N_26795);
xor U27032 (N_27032,N_26789,N_26541);
xnor U27033 (N_27033,N_26504,N_26527);
nor U27034 (N_27034,N_26531,N_26867);
and U27035 (N_27035,N_26508,N_26735);
and U27036 (N_27036,N_26824,N_26565);
or U27037 (N_27037,N_26534,N_26978);
or U27038 (N_27038,N_26947,N_26670);
xnor U27039 (N_27039,N_26866,N_26944);
nor U27040 (N_27040,N_26792,N_26666);
xnor U27041 (N_27041,N_26839,N_26826);
or U27042 (N_27042,N_26847,N_26556);
and U27043 (N_27043,N_26938,N_26729);
and U27044 (N_27044,N_26708,N_26611);
and U27045 (N_27045,N_26624,N_26859);
xor U27046 (N_27046,N_26891,N_26590);
and U27047 (N_27047,N_26509,N_26753);
xor U27048 (N_27048,N_26778,N_26502);
nand U27049 (N_27049,N_26910,N_26649);
xor U27050 (N_27050,N_26627,N_26780);
or U27051 (N_27051,N_26854,N_26752);
nor U27052 (N_27052,N_26713,N_26526);
or U27053 (N_27053,N_26894,N_26808);
xor U27054 (N_27054,N_26790,N_26896);
or U27055 (N_27055,N_26836,N_26799);
and U27056 (N_27056,N_26614,N_26775);
nor U27057 (N_27057,N_26997,N_26879);
and U27058 (N_27058,N_26766,N_26736);
nor U27059 (N_27059,N_26844,N_26831);
and U27060 (N_27060,N_26846,N_26750);
nand U27061 (N_27061,N_26945,N_26683);
nand U27062 (N_27062,N_26988,N_26884);
xnor U27063 (N_27063,N_26832,N_26791);
nor U27064 (N_27064,N_26626,N_26969);
or U27065 (N_27065,N_26967,N_26906);
nor U27066 (N_27066,N_26700,N_26647);
and U27067 (N_27067,N_26941,N_26511);
or U27068 (N_27068,N_26620,N_26578);
xor U27069 (N_27069,N_26678,N_26676);
xnor U27070 (N_27070,N_26782,N_26591);
xnor U27071 (N_27071,N_26857,N_26830);
xor U27072 (N_27072,N_26918,N_26507);
nand U27073 (N_27073,N_26838,N_26707);
or U27074 (N_27074,N_26730,N_26505);
or U27075 (N_27075,N_26914,N_26812);
and U27076 (N_27076,N_26767,N_26855);
nor U27077 (N_27077,N_26919,N_26963);
nand U27078 (N_27078,N_26672,N_26943);
or U27079 (N_27079,N_26907,N_26746);
or U27080 (N_27080,N_26996,N_26779);
or U27081 (N_27081,N_26719,N_26569);
and U27082 (N_27082,N_26592,N_26632);
nor U27083 (N_27083,N_26821,N_26638);
nand U27084 (N_27084,N_26913,N_26915);
xor U27085 (N_27085,N_26607,N_26706);
and U27086 (N_27086,N_26558,N_26876);
nor U27087 (N_27087,N_26774,N_26805);
xor U27088 (N_27088,N_26555,N_26922);
or U27089 (N_27089,N_26865,N_26581);
xor U27090 (N_27090,N_26692,N_26965);
nand U27091 (N_27091,N_26513,N_26618);
xor U27092 (N_27092,N_26874,N_26681);
or U27093 (N_27093,N_26663,N_26580);
and U27094 (N_27094,N_26725,N_26723);
and U27095 (N_27095,N_26568,N_26842);
and U27096 (N_27096,N_26807,N_26619);
xnor U27097 (N_27097,N_26570,N_26966);
and U27098 (N_27098,N_26543,N_26895);
or U27099 (N_27099,N_26740,N_26893);
xor U27100 (N_27100,N_26986,N_26856);
and U27101 (N_27101,N_26897,N_26933);
nand U27102 (N_27102,N_26950,N_26733);
nand U27103 (N_27103,N_26903,N_26561);
xor U27104 (N_27104,N_26822,N_26977);
nand U27105 (N_27105,N_26751,N_26699);
nor U27106 (N_27106,N_26809,N_26694);
and U27107 (N_27107,N_26829,N_26520);
and U27108 (N_27108,N_26994,N_26688);
nand U27109 (N_27109,N_26501,N_26515);
or U27110 (N_27110,N_26557,N_26551);
nor U27111 (N_27111,N_26677,N_26595);
nand U27112 (N_27112,N_26671,N_26912);
xnor U27113 (N_27113,N_26667,N_26727);
nor U27114 (N_27114,N_26675,N_26639);
nor U27115 (N_27115,N_26816,N_26603);
nand U27116 (N_27116,N_26889,N_26575);
nor U27117 (N_27117,N_26981,N_26658);
xor U27118 (N_27118,N_26579,N_26754);
nand U27119 (N_27119,N_26695,N_26870);
nor U27120 (N_27120,N_26763,N_26640);
nor U27121 (N_27121,N_26629,N_26540);
and U27122 (N_27122,N_26605,N_26552);
and U27123 (N_27123,N_26616,N_26800);
or U27124 (N_27124,N_26972,N_26732);
nor U27125 (N_27125,N_26528,N_26659);
or U27126 (N_27126,N_26848,N_26979);
nor U27127 (N_27127,N_26518,N_26567);
or U27128 (N_27128,N_26962,N_26762);
xnor U27129 (N_27129,N_26742,N_26760);
and U27130 (N_27130,N_26547,N_26572);
or U27131 (N_27131,N_26637,N_26604);
and U27132 (N_27132,N_26940,N_26987);
and U27133 (N_27133,N_26873,N_26989);
nor U27134 (N_27134,N_26784,N_26927);
nand U27135 (N_27135,N_26928,N_26954);
and U27136 (N_27136,N_26715,N_26546);
or U27137 (N_27137,N_26646,N_26872);
nor U27138 (N_27138,N_26880,N_26655);
and U27139 (N_27139,N_26923,N_26609);
xor U27140 (N_27140,N_26693,N_26722);
and U27141 (N_27141,N_26529,N_26970);
xor U27142 (N_27142,N_26818,N_26932);
nand U27143 (N_27143,N_26642,N_26623);
xor U27144 (N_27144,N_26716,N_26517);
nand U27145 (N_27145,N_26522,N_26802);
nand U27146 (N_27146,N_26959,N_26636);
xor U27147 (N_27147,N_26968,N_26925);
nand U27148 (N_27148,N_26576,N_26532);
xor U27149 (N_27149,N_26653,N_26960);
or U27150 (N_27150,N_26863,N_26705);
or U27151 (N_27151,N_26500,N_26562);
or U27152 (N_27152,N_26606,N_26777);
or U27153 (N_27153,N_26617,N_26726);
nor U27154 (N_27154,N_26890,N_26851);
nand U27155 (N_27155,N_26793,N_26902);
nand U27156 (N_27156,N_26524,N_26900);
or U27157 (N_27157,N_26712,N_26682);
and U27158 (N_27158,N_26937,N_26813);
or U27159 (N_27159,N_26901,N_26625);
and U27160 (N_27160,N_26628,N_26761);
and U27161 (N_27161,N_26768,N_26539);
xor U27162 (N_27162,N_26869,N_26765);
or U27163 (N_27163,N_26698,N_26833);
xnor U27164 (N_27164,N_26593,N_26701);
nand U27165 (N_27165,N_26660,N_26709);
or U27166 (N_27166,N_26686,N_26521);
nand U27167 (N_27167,N_26644,N_26827);
xor U27168 (N_27168,N_26991,N_26796);
and U27169 (N_27169,N_26999,N_26608);
xnor U27170 (N_27170,N_26961,N_26545);
nand U27171 (N_27171,N_26955,N_26845);
nor U27172 (N_27172,N_26586,N_26820);
nor U27173 (N_27173,N_26594,N_26843);
nor U27174 (N_27174,N_26926,N_26957);
xnor U27175 (N_27175,N_26622,N_26588);
and U27176 (N_27176,N_26942,N_26939);
nor U27177 (N_27177,N_26982,N_26853);
nand U27178 (N_27178,N_26776,N_26975);
and U27179 (N_27179,N_26720,N_26823);
and U27180 (N_27180,N_26697,N_26691);
nand U27181 (N_27181,N_26573,N_26783);
or U27182 (N_27182,N_26862,N_26984);
or U27183 (N_27183,N_26600,N_26815);
xor U27184 (N_27184,N_26535,N_26657);
nand U27185 (N_27185,N_26566,N_26721);
or U27186 (N_27186,N_26755,N_26702);
or U27187 (N_27187,N_26728,N_26801);
xor U27188 (N_27188,N_26503,N_26743);
and U27189 (N_27189,N_26512,N_26643);
nor U27190 (N_27190,N_26601,N_26916);
nand U27191 (N_27191,N_26748,N_26905);
nand U27192 (N_27192,N_26560,N_26993);
and U27193 (N_27193,N_26788,N_26741);
xor U27194 (N_27194,N_26564,N_26656);
and U27195 (N_27195,N_26980,N_26710);
xor U27196 (N_27196,N_26861,N_26798);
and U27197 (N_27197,N_26759,N_26810);
nor U27198 (N_27198,N_26533,N_26911);
xor U27199 (N_27199,N_26948,N_26992);
nand U27200 (N_27200,N_26734,N_26745);
or U27201 (N_27201,N_26554,N_26651);
nand U27202 (N_27202,N_26875,N_26757);
nor U27203 (N_27203,N_26882,N_26883);
nand U27204 (N_27204,N_26908,N_26976);
and U27205 (N_27205,N_26516,N_26899);
xnor U27206 (N_27206,N_26973,N_26641);
nand U27207 (N_27207,N_26679,N_26673);
xor U27208 (N_27208,N_26985,N_26652);
xnor U27209 (N_27209,N_26731,N_26995);
xor U27210 (N_27210,N_26860,N_26786);
xnor U27211 (N_27211,N_26787,N_26571);
nor U27212 (N_27212,N_26904,N_26696);
and U27213 (N_27213,N_26525,N_26610);
nor U27214 (N_27214,N_26930,N_26739);
and U27215 (N_27215,N_26770,N_26718);
nor U27216 (N_27216,N_26886,N_26650);
or U27217 (N_27217,N_26858,N_26621);
nor U27218 (N_27218,N_26864,N_26553);
or U27219 (N_27219,N_26811,N_26645);
nand U27220 (N_27220,N_26785,N_26769);
and U27221 (N_27221,N_26737,N_26803);
and U27222 (N_27222,N_26877,N_26633);
and U27223 (N_27223,N_26506,N_26613);
nand U27224 (N_27224,N_26530,N_26929);
nor U27225 (N_27225,N_26772,N_26587);
or U27226 (N_27226,N_26584,N_26825);
nand U27227 (N_27227,N_26703,N_26964);
and U27228 (N_27228,N_26834,N_26828);
and U27229 (N_27229,N_26917,N_26559);
nand U27230 (N_27230,N_26631,N_26665);
xnor U27231 (N_27231,N_26953,N_26758);
xnor U27232 (N_27232,N_26949,N_26924);
nor U27233 (N_27233,N_26951,N_26577);
and U27234 (N_27234,N_26841,N_26589);
nand U27235 (N_27235,N_26668,N_26685);
xnor U27236 (N_27236,N_26952,N_26887);
and U27237 (N_27237,N_26661,N_26819);
or U27238 (N_27238,N_26630,N_26550);
xnor U27239 (N_27239,N_26738,N_26934);
nand U27240 (N_27240,N_26974,N_26771);
xor U27241 (N_27241,N_26840,N_26662);
nor U27242 (N_27242,N_26806,N_26935);
nor U27243 (N_27243,N_26510,N_26536);
nor U27244 (N_27244,N_26797,N_26764);
and U27245 (N_27245,N_26885,N_26781);
xnor U27246 (N_27246,N_26602,N_26998);
nand U27247 (N_27247,N_26635,N_26804);
nand U27248 (N_27248,N_26756,N_26582);
nor U27249 (N_27249,N_26689,N_26519);
and U27250 (N_27250,N_26638,N_26873);
xnor U27251 (N_27251,N_26710,N_26842);
or U27252 (N_27252,N_26908,N_26931);
nand U27253 (N_27253,N_26991,N_26741);
and U27254 (N_27254,N_26779,N_26673);
nor U27255 (N_27255,N_26718,N_26885);
nor U27256 (N_27256,N_26962,N_26896);
xor U27257 (N_27257,N_26792,N_26593);
or U27258 (N_27258,N_26615,N_26929);
xnor U27259 (N_27259,N_26959,N_26803);
nor U27260 (N_27260,N_26701,N_26607);
nand U27261 (N_27261,N_26888,N_26523);
and U27262 (N_27262,N_26724,N_26917);
and U27263 (N_27263,N_26872,N_26567);
nor U27264 (N_27264,N_26954,N_26715);
nand U27265 (N_27265,N_26686,N_26976);
xnor U27266 (N_27266,N_26970,N_26898);
and U27267 (N_27267,N_26512,N_26977);
xnor U27268 (N_27268,N_26666,N_26796);
xnor U27269 (N_27269,N_26785,N_26681);
and U27270 (N_27270,N_26658,N_26788);
nand U27271 (N_27271,N_26700,N_26990);
nand U27272 (N_27272,N_26879,N_26883);
xor U27273 (N_27273,N_26608,N_26546);
or U27274 (N_27274,N_26822,N_26820);
xor U27275 (N_27275,N_26758,N_26720);
xor U27276 (N_27276,N_26886,N_26607);
and U27277 (N_27277,N_26700,N_26845);
xor U27278 (N_27278,N_26664,N_26833);
xor U27279 (N_27279,N_26855,N_26950);
or U27280 (N_27280,N_26864,N_26818);
xor U27281 (N_27281,N_26842,N_26984);
and U27282 (N_27282,N_26888,N_26883);
nand U27283 (N_27283,N_26898,N_26511);
nand U27284 (N_27284,N_26541,N_26873);
or U27285 (N_27285,N_26780,N_26929);
or U27286 (N_27286,N_26516,N_26598);
xnor U27287 (N_27287,N_26663,N_26569);
or U27288 (N_27288,N_26749,N_26720);
nand U27289 (N_27289,N_26904,N_26518);
xnor U27290 (N_27290,N_26754,N_26881);
nand U27291 (N_27291,N_26650,N_26834);
or U27292 (N_27292,N_26745,N_26819);
nand U27293 (N_27293,N_26832,N_26659);
nand U27294 (N_27294,N_26647,N_26690);
xor U27295 (N_27295,N_26958,N_26880);
nor U27296 (N_27296,N_26992,N_26554);
or U27297 (N_27297,N_26602,N_26662);
nand U27298 (N_27298,N_26560,N_26555);
xnor U27299 (N_27299,N_26759,N_26646);
xor U27300 (N_27300,N_26600,N_26810);
or U27301 (N_27301,N_26934,N_26762);
and U27302 (N_27302,N_26749,N_26979);
nor U27303 (N_27303,N_26510,N_26668);
xor U27304 (N_27304,N_26919,N_26664);
xor U27305 (N_27305,N_26823,N_26982);
and U27306 (N_27306,N_26928,N_26534);
nand U27307 (N_27307,N_26668,N_26730);
and U27308 (N_27308,N_26899,N_26867);
nand U27309 (N_27309,N_26668,N_26698);
and U27310 (N_27310,N_26793,N_26866);
nand U27311 (N_27311,N_26516,N_26611);
or U27312 (N_27312,N_26793,N_26597);
and U27313 (N_27313,N_26838,N_26779);
nand U27314 (N_27314,N_26574,N_26940);
and U27315 (N_27315,N_26933,N_26630);
nand U27316 (N_27316,N_26993,N_26818);
and U27317 (N_27317,N_26664,N_26710);
or U27318 (N_27318,N_26531,N_26552);
xor U27319 (N_27319,N_26618,N_26946);
or U27320 (N_27320,N_26783,N_26976);
nand U27321 (N_27321,N_26826,N_26577);
nor U27322 (N_27322,N_26650,N_26671);
xor U27323 (N_27323,N_26549,N_26534);
xnor U27324 (N_27324,N_26615,N_26837);
nor U27325 (N_27325,N_26793,N_26816);
or U27326 (N_27326,N_26767,N_26740);
nor U27327 (N_27327,N_26559,N_26939);
and U27328 (N_27328,N_26941,N_26938);
and U27329 (N_27329,N_26961,N_26810);
or U27330 (N_27330,N_26982,N_26770);
or U27331 (N_27331,N_26644,N_26672);
xor U27332 (N_27332,N_26904,N_26703);
xor U27333 (N_27333,N_26702,N_26535);
nor U27334 (N_27334,N_26538,N_26738);
nor U27335 (N_27335,N_26625,N_26980);
nor U27336 (N_27336,N_26740,N_26509);
xor U27337 (N_27337,N_26747,N_26527);
and U27338 (N_27338,N_26648,N_26645);
xnor U27339 (N_27339,N_26587,N_26898);
xor U27340 (N_27340,N_26500,N_26885);
nand U27341 (N_27341,N_26685,N_26620);
xnor U27342 (N_27342,N_26512,N_26692);
xnor U27343 (N_27343,N_26527,N_26559);
and U27344 (N_27344,N_26670,N_26921);
nand U27345 (N_27345,N_26561,N_26868);
or U27346 (N_27346,N_26661,N_26569);
xor U27347 (N_27347,N_26810,N_26642);
nor U27348 (N_27348,N_26642,N_26980);
nor U27349 (N_27349,N_26958,N_26882);
nor U27350 (N_27350,N_26929,N_26793);
and U27351 (N_27351,N_26999,N_26779);
and U27352 (N_27352,N_26696,N_26922);
xnor U27353 (N_27353,N_26791,N_26883);
and U27354 (N_27354,N_26878,N_26630);
nor U27355 (N_27355,N_26955,N_26837);
nor U27356 (N_27356,N_26755,N_26635);
nor U27357 (N_27357,N_26638,N_26544);
nor U27358 (N_27358,N_26796,N_26596);
and U27359 (N_27359,N_26869,N_26535);
nor U27360 (N_27360,N_26882,N_26561);
nand U27361 (N_27361,N_26824,N_26729);
xor U27362 (N_27362,N_26548,N_26746);
and U27363 (N_27363,N_26503,N_26553);
nor U27364 (N_27364,N_26650,N_26581);
and U27365 (N_27365,N_26853,N_26762);
or U27366 (N_27366,N_26668,N_26818);
xnor U27367 (N_27367,N_26848,N_26599);
and U27368 (N_27368,N_26751,N_26624);
nand U27369 (N_27369,N_26745,N_26550);
nand U27370 (N_27370,N_26755,N_26717);
nor U27371 (N_27371,N_26679,N_26766);
or U27372 (N_27372,N_26626,N_26642);
and U27373 (N_27373,N_26976,N_26899);
xor U27374 (N_27374,N_26818,N_26878);
nand U27375 (N_27375,N_26990,N_26979);
and U27376 (N_27376,N_26665,N_26868);
or U27377 (N_27377,N_26970,N_26839);
nand U27378 (N_27378,N_26713,N_26902);
xnor U27379 (N_27379,N_26730,N_26800);
nand U27380 (N_27380,N_26542,N_26851);
or U27381 (N_27381,N_26657,N_26667);
nand U27382 (N_27382,N_26993,N_26913);
and U27383 (N_27383,N_26986,N_26530);
nor U27384 (N_27384,N_26506,N_26799);
xnor U27385 (N_27385,N_26689,N_26914);
and U27386 (N_27386,N_26988,N_26582);
or U27387 (N_27387,N_26972,N_26733);
xor U27388 (N_27388,N_26571,N_26777);
or U27389 (N_27389,N_26511,N_26799);
xnor U27390 (N_27390,N_26548,N_26741);
nor U27391 (N_27391,N_26862,N_26606);
and U27392 (N_27392,N_26655,N_26980);
nand U27393 (N_27393,N_26754,N_26909);
nand U27394 (N_27394,N_26901,N_26943);
or U27395 (N_27395,N_26945,N_26612);
xnor U27396 (N_27396,N_26532,N_26751);
and U27397 (N_27397,N_26720,N_26571);
or U27398 (N_27398,N_26688,N_26818);
xnor U27399 (N_27399,N_26926,N_26884);
and U27400 (N_27400,N_26550,N_26578);
nor U27401 (N_27401,N_26683,N_26634);
nand U27402 (N_27402,N_26975,N_26700);
xnor U27403 (N_27403,N_26792,N_26560);
or U27404 (N_27404,N_26723,N_26599);
nor U27405 (N_27405,N_26643,N_26603);
nand U27406 (N_27406,N_26540,N_26894);
nor U27407 (N_27407,N_26614,N_26603);
nor U27408 (N_27408,N_26982,N_26581);
and U27409 (N_27409,N_26605,N_26506);
and U27410 (N_27410,N_26837,N_26959);
nor U27411 (N_27411,N_26927,N_26619);
or U27412 (N_27412,N_26560,N_26584);
or U27413 (N_27413,N_26979,N_26994);
nand U27414 (N_27414,N_26841,N_26530);
and U27415 (N_27415,N_26751,N_26805);
nor U27416 (N_27416,N_26606,N_26697);
nor U27417 (N_27417,N_26857,N_26701);
and U27418 (N_27418,N_26751,N_26777);
nor U27419 (N_27419,N_26786,N_26934);
or U27420 (N_27420,N_26521,N_26747);
xnor U27421 (N_27421,N_26777,N_26586);
xnor U27422 (N_27422,N_26779,N_26524);
and U27423 (N_27423,N_26872,N_26656);
xnor U27424 (N_27424,N_26860,N_26542);
or U27425 (N_27425,N_26669,N_26768);
xnor U27426 (N_27426,N_26825,N_26952);
or U27427 (N_27427,N_26695,N_26696);
xnor U27428 (N_27428,N_26538,N_26603);
nand U27429 (N_27429,N_26842,N_26748);
nand U27430 (N_27430,N_26907,N_26903);
or U27431 (N_27431,N_26726,N_26985);
nand U27432 (N_27432,N_26703,N_26726);
xnor U27433 (N_27433,N_26695,N_26766);
xnor U27434 (N_27434,N_26528,N_26871);
or U27435 (N_27435,N_26742,N_26991);
and U27436 (N_27436,N_26785,N_26690);
nor U27437 (N_27437,N_26955,N_26603);
nand U27438 (N_27438,N_26698,N_26966);
or U27439 (N_27439,N_26725,N_26651);
or U27440 (N_27440,N_26533,N_26962);
xnor U27441 (N_27441,N_26900,N_26946);
nand U27442 (N_27442,N_26790,N_26888);
nand U27443 (N_27443,N_26560,N_26931);
nand U27444 (N_27444,N_26892,N_26651);
or U27445 (N_27445,N_26709,N_26640);
or U27446 (N_27446,N_26770,N_26974);
nand U27447 (N_27447,N_26862,N_26854);
xor U27448 (N_27448,N_26828,N_26651);
xnor U27449 (N_27449,N_26855,N_26634);
and U27450 (N_27450,N_26937,N_26612);
and U27451 (N_27451,N_26781,N_26745);
and U27452 (N_27452,N_26550,N_26753);
or U27453 (N_27453,N_26597,N_26882);
nand U27454 (N_27454,N_26993,N_26689);
or U27455 (N_27455,N_26806,N_26559);
nor U27456 (N_27456,N_26703,N_26754);
nand U27457 (N_27457,N_26958,N_26798);
nor U27458 (N_27458,N_26667,N_26802);
and U27459 (N_27459,N_26801,N_26892);
nor U27460 (N_27460,N_26690,N_26942);
nand U27461 (N_27461,N_26730,N_26680);
or U27462 (N_27462,N_26509,N_26929);
nor U27463 (N_27463,N_26534,N_26639);
or U27464 (N_27464,N_26970,N_26909);
nor U27465 (N_27465,N_26537,N_26568);
or U27466 (N_27466,N_26925,N_26951);
or U27467 (N_27467,N_26563,N_26926);
and U27468 (N_27468,N_26529,N_26815);
or U27469 (N_27469,N_26581,N_26653);
nor U27470 (N_27470,N_26607,N_26589);
nor U27471 (N_27471,N_26833,N_26944);
nand U27472 (N_27472,N_26636,N_26781);
nand U27473 (N_27473,N_26655,N_26695);
and U27474 (N_27474,N_26725,N_26763);
nor U27475 (N_27475,N_26617,N_26693);
xor U27476 (N_27476,N_26988,N_26876);
and U27477 (N_27477,N_26971,N_26997);
or U27478 (N_27478,N_26698,N_26615);
nor U27479 (N_27479,N_26561,N_26850);
xnor U27480 (N_27480,N_26853,N_26789);
nor U27481 (N_27481,N_26844,N_26505);
xor U27482 (N_27482,N_26737,N_26741);
or U27483 (N_27483,N_26773,N_26566);
nand U27484 (N_27484,N_26611,N_26683);
and U27485 (N_27485,N_26972,N_26816);
nor U27486 (N_27486,N_26699,N_26585);
xor U27487 (N_27487,N_26928,N_26715);
and U27488 (N_27488,N_26957,N_26609);
and U27489 (N_27489,N_26738,N_26658);
nand U27490 (N_27490,N_26597,N_26765);
xor U27491 (N_27491,N_26513,N_26816);
or U27492 (N_27492,N_26773,N_26732);
or U27493 (N_27493,N_26785,N_26550);
or U27494 (N_27494,N_26700,N_26842);
or U27495 (N_27495,N_26950,N_26579);
xnor U27496 (N_27496,N_26514,N_26630);
nand U27497 (N_27497,N_26680,N_26546);
or U27498 (N_27498,N_26983,N_26649);
and U27499 (N_27499,N_26567,N_26930);
or U27500 (N_27500,N_27326,N_27176);
xnor U27501 (N_27501,N_27079,N_27154);
and U27502 (N_27502,N_27467,N_27409);
or U27503 (N_27503,N_27072,N_27076);
and U27504 (N_27504,N_27363,N_27465);
xnor U27505 (N_27505,N_27429,N_27066);
and U27506 (N_27506,N_27395,N_27005);
or U27507 (N_27507,N_27125,N_27400);
xnor U27508 (N_27508,N_27206,N_27373);
nor U27509 (N_27509,N_27362,N_27484);
and U27510 (N_27510,N_27211,N_27290);
or U27511 (N_27511,N_27455,N_27101);
and U27512 (N_27512,N_27388,N_27051);
and U27513 (N_27513,N_27139,N_27311);
and U27514 (N_27514,N_27392,N_27038);
nor U27515 (N_27515,N_27365,N_27452);
and U27516 (N_27516,N_27394,N_27399);
and U27517 (N_27517,N_27445,N_27095);
and U27518 (N_27518,N_27466,N_27314);
nor U27519 (N_27519,N_27093,N_27319);
nor U27520 (N_27520,N_27411,N_27096);
nand U27521 (N_27521,N_27118,N_27396);
nor U27522 (N_27522,N_27062,N_27166);
xor U27523 (N_27523,N_27043,N_27324);
or U27524 (N_27524,N_27121,N_27074);
or U27525 (N_27525,N_27350,N_27247);
and U27526 (N_27526,N_27416,N_27194);
xor U27527 (N_27527,N_27495,N_27011);
nand U27528 (N_27528,N_27190,N_27478);
xor U27529 (N_27529,N_27272,N_27178);
or U27530 (N_27530,N_27420,N_27331);
and U27531 (N_27531,N_27209,N_27286);
nor U27532 (N_27532,N_27345,N_27022);
and U27533 (N_27533,N_27298,N_27262);
nor U27534 (N_27534,N_27199,N_27168);
xor U27535 (N_27535,N_27342,N_27171);
or U27536 (N_27536,N_27320,N_27404);
and U27537 (N_27537,N_27008,N_27481);
nand U27538 (N_27538,N_27431,N_27334);
xor U27539 (N_27539,N_27348,N_27182);
nand U27540 (N_27540,N_27053,N_27160);
xor U27541 (N_27541,N_27110,N_27189);
xor U27542 (N_27542,N_27493,N_27167);
xnor U27543 (N_27543,N_27047,N_27258);
xnor U27544 (N_27544,N_27186,N_27122);
xor U27545 (N_27545,N_27149,N_27418);
or U27546 (N_27546,N_27057,N_27210);
or U27547 (N_27547,N_27475,N_27274);
and U27548 (N_27548,N_27023,N_27035);
or U27549 (N_27549,N_27024,N_27039);
xnor U27550 (N_27550,N_27054,N_27486);
and U27551 (N_27551,N_27260,N_27414);
xor U27552 (N_27552,N_27044,N_27491);
nor U27553 (N_27553,N_27347,N_27236);
nor U27554 (N_27554,N_27150,N_27113);
and U27555 (N_27555,N_27041,N_27198);
nor U27556 (N_27556,N_27461,N_27226);
and U27557 (N_27557,N_27369,N_27317);
nor U27558 (N_27558,N_27257,N_27151);
or U27559 (N_27559,N_27213,N_27378);
nand U27560 (N_27560,N_27059,N_27425);
and U27561 (N_27561,N_27124,N_27427);
and U27562 (N_27562,N_27215,N_27480);
or U27563 (N_27563,N_27380,N_27048);
nor U27564 (N_27564,N_27398,N_27296);
xnor U27565 (N_27565,N_27034,N_27292);
and U27566 (N_27566,N_27437,N_27128);
nand U27567 (N_27567,N_27473,N_27476);
or U27568 (N_27568,N_27126,N_27134);
nor U27569 (N_27569,N_27393,N_27007);
nand U27570 (N_27570,N_27088,N_27438);
or U27571 (N_27571,N_27436,N_27318);
nor U27572 (N_27572,N_27137,N_27158);
xor U27573 (N_27573,N_27338,N_27025);
xnor U27574 (N_27574,N_27141,N_27267);
nand U27575 (N_27575,N_27360,N_27441);
and U27576 (N_27576,N_27100,N_27092);
nand U27577 (N_27577,N_27001,N_27470);
and U27578 (N_27578,N_27401,N_27090);
nand U27579 (N_27579,N_27245,N_27063);
nor U27580 (N_27580,N_27002,N_27143);
or U27581 (N_27581,N_27234,N_27253);
nand U27582 (N_27582,N_27287,N_27197);
nor U27583 (N_27583,N_27387,N_27336);
or U27584 (N_27584,N_27322,N_27289);
or U27585 (N_27585,N_27270,N_27277);
and U27586 (N_27586,N_27312,N_27216);
xor U27587 (N_27587,N_27162,N_27045);
nor U27588 (N_27588,N_27165,N_27083);
and U27589 (N_27589,N_27085,N_27444);
nor U27590 (N_27590,N_27443,N_27228);
and U27591 (N_27591,N_27352,N_27397);
nand U27592 (N_27592,N_27281,N_27372);
and U27593 (N_27593,N_27172,N_27329);
nor U27594 (N_27594,N_27094,N_27152);
nor U27595 (N_27595,N_27303,N_27354);
and U27596 (N_27596,N_27271,N_27227);
nor U27597 (N_27597,N_27114,N_27243);
nand U27598 (N_27598,N_27458,N_27061);
xnor U27599 (N_27599,N_27446,N_27067);
nor U27600 (N_27600,N_27056,N_27408);
nor U27601 (N_27601,N_27340,N_27027);
xnor U27602 (N_27602,N_27159,N_27412);
or U27603 (N_27603,N_27019,N_27136);
nand U27604 (N_27604,N_27081,N_27106);
nor U27605 (N_27605,N_27280,N_27310);
nor U27606 (N_27606,N_27488,N_27265);
and U27607 (N_27607,N_27353,N_27483);
nand U27608 (N_27608,N_27434,N_27084);
and U27609 (N_27609,N_27295,N_27482);
or U27610 (N_27610,N_27423,N_27264);
or U27611 (N_27611,N_27323,N_27077);
or U27612 (N_27612,N_27275,N_27115);
nand U27613 (N_27613,N_27366,N_27021);
and U27614 (N_27614,N_27492,N_27069);
nand U27615 (N_27615,N_27464,N_27435);
or U27616 (N_27616,N_27278,N_27055);
and U27617 (N_27617,N_27407,N_27183);
nor U27618 (N_27618,N_27138,N_27489);
or U27619 (N_27619,N_27391,N_27268);
nor U27620 (N_27620,N_27419,N_27225);
nor U27621 (N_27621,N_27450,N_27117);
nor U27622 (N_27622,N_27107,N_27223);
nand U27623 (N_27623,N_27238,N_27376);
or U27624 (N_27624,N_27367,N_27109);
nand U27625 (N_27625,N_27073,N_27448);
xor U27626 (N_27626,N_27468,N_27357);
xnor U27627 (N_27627,N_27200,N_27358);
nor U27628 (N_27628,N_27191,N_27184);
xor U27629 (N_27629,N_27164,N_27018);
and U27630 (N_27630,N_27327,N_27104);
nor U27631 (N_27631,N_27263,N_27349);
nand U27632 (N_27632,N_27006,N_27294);
nand U27633 (N_27633,N_27193,N_27355);
nand U27634 (N_27634,N_27205,N_27037);
or U27635 (N_27635,N_27413,N_27368);
nor U27636 (N_27636,N_27010,N_27179);
xnor U27637 (N_27637,N_27250,N_27442);
or U27638 (N_27638,N_27089,N_27333);
xor U27639 (N_27639,N_27014,N_27454);
nor U27640 (N_27640,N_27325,N_27246);
xnor U27641 (N_27641,N_27239,N_27221);
nand U27642 (N_27642,N_27487,N_27432);
and U27643 (N_27643,N_27112,N_27147);
or U27644 (N_27644,N_27332,N_27163);
and U27645 (N_27645,N_27224,N_27406);
xor U27646 (N_27646,N_27430,N_27075);
xnor U27647 (N_27647,N_27328,N_27249);
nor U27648 (N_27648,N_27173,N_27098);
nor U27649 (N_27649,N_27012,N_27015);
or U27650 (N_27650,N_27201,N_27175);
or U27651 (N_27651,N_27214,N_27346);
and U27652 (N_27652,N_27030,N_27485);
nor U27653 (N_27653,N_27241,N_27259);
or U27654 (N_27654,N_27299,N_27208);
nor U27655 (N_27655,N_27004,N_27130);
nor U27656 (N_27656,N_27086,N_27305);
nor U27657 (N_27657,N_27082,N_27440);
nand U27658 (N_27658,N_27282,N_27129);
or U27659 (N_27659,N_27049,N_27170);
nand U27660 (N_27660,N_27252,N_27217);
xor U27661 (N_27661,N_27451,N_27251);
or U27662 (N_27662,N_27279,N_27212);
nor U27663 (N_27663,N_27218,N_27091);
nor U27664 (N_27664,N_27181,N_27196);
xnor U27665 (N_27665,N_27422,N_27254);
nor U27666 (N_27666,N_27188,N_27306);
and U27667 (N_27667,N_27140,N_27050);
and U27668 (N_27668,N_27309,N_27403);
xnor U27669 (N_27669,N_27477,N_27060);
and U27670 (N_27670,N_27370,N_27235);
and U27671 (N_27671,N_27374,N_27195);
nand U27672 (N_27672,N_27169,N_27156);
or U27673 (N_27673,N_27105,N_27026);
nand U27674 (N_27674,N_27284,N_27462);
nand U27675 (N_27675,N_27364,N_27233);
and U27676 (N_27676,N_27207,N_27383);
and U27677 (N_27677,N_27269,N_27116);
nor U27678 (N_27678,N_27017,N_27421);
nand U27679 (N_27679,N_27457,N_27231);
and U27680 (N_27680,N_27127,N_27071);
xor U27681 (N_27681,N_27204,N_27261);
nor U27682 (N_27682,N_27029,N_27131);
and U27683 (N_27683,N_27293,N_27174);
or U27684 (N_27684,N_27361,N_27424);
nor U27685 (N_27685,N_27405,N_27285);
nor U27686 (N_27686,N_27145,N_27428);
and U27687 (N_27687,N_27132,N_27490);
nand U27688 (N_27688,N_27237,N_27111);
and U27689 (N_27689,N_27120,N_27315);
and U27690 (N_27690,N_27052,N_27499);
nor U27691 (N_27691,N_27003,N_27087);
or U27692 (N_27692,N_27463,N_27013);
or U27693 (N_27693,N_27185,N_27177);
nand U27694 (N_27694,N_27460,N_27356);
and U27695 (N_27695,N_27375,N_27222);
nor U27696 (N_27696,N_27288,N_27036);
and U27697 (N_27697,N_27449,N_27433);
and U27698 (N_27698,N_27058,N_27135);
and U27699 (N_27699,N_27313,N_27020);
nor U27700 (N_27700,N_27123,N_27273);
or U27701 (N_27701,N_27339,N_27144);
nand U27702 (N_27702,N_27161,N_27351);
nor U27703 (N_27703,N_27343,N_27240);
or U27704 (N_27704,N_27302,N_27078);
nor U27705 (N_27705,N_27080,N_27046);
nor U27706 (N_27706,N_27180,N_27300);
xnor U27707 (N_27707,N_27496,N_27417);
and U27708 (N_27708,N_27479,N_27494);
nor U27709 (N_27709,N_27133,N_27308);
or U27710 (N_27710,N_27384,N_27472);
xnor U27711 (N_27711,N_27377,N_27390);
and U27712 (N_27712,N_27359,N_27065);
xor U27713 (N_27713,N_27297,N_27291);
and U27714 (N_27714,N_27187,N_27382);
xor U27715 (N_27715,N_27456,N_27379);
and U27716 (N_27716,N_27203,N_27341);
or U27717 (N_27717,N_27068,N_27097);
or U27718 (N_27718,N_27344,N_27371);
or U27719 (N_27719,N_27155,N_27229);
xor U27720 (N_27720,N_27148,N_27410);
nor U27721 (N_27721,N_27232,N_27330);
or U27722 (N_27722,N_27402,N_27381);
nor U27723 (N_27723,N_27248,N_27256);
xor U27724 (N_27724,N_27283,N_27386);
nand U27725 (N_27725,N_27244,N_27119);
xnor U27726 (N_27726,N_27103,N_27070);
and U27727 (N_27727,N_27108,N_27192);
nor U27728 (N_27728,N_27471,N_27202);
or U27729 (N_27729,N_27307,N_27453);
nand U27730 (N_27730,N_27157,N_27459);
and U27731 (N_27731,N_27219,N_27276);
and U27732 (N_27732,N_27042,N_27102);
and U27733 (N_27733,N_27439,N_27099);
or U27734 (N_27734,N_27497,N_27031);
and U27735 (N_27735,N_27142,N_27316);
nor U27736 (N_27736,N_27474,N_27469);
or U27737 (N_27737,N_27220,N_27016);
or U27738 (N_27738,N_27498,N_27153);
or U27739 (N_27739,N_27033,N_27009);
xor U27740 (N_27740,N_27337,N_27335);
xor U27741 (N_27741,N_27064,N_27301);
nor U27742 (N_27742,N_27415,N_27000);
nand U27743 (N_27743,N_27447,N_27426);
xor U27744 (N_27744,N_27146,N_27032);
or U27745 (N_27745,N_27255,N_27242);
xnor U27746 (N_27746,N_27304,N_27266);
or U27747 (N_27747,N_27040,N_27230);
nor U27748 (N_27748,N_27321,N_27389);
or U27749 (N_27749,N_27028,N_27385);
xor U27750 (N_27750,N_27434,N_27315);
xnor U27751 (N_27751,N_27285,N_27152);
xor U27752 (N_27752,N_27341,N_27198);
nor U27753 (N_27753,N_27204,N_27391);
nand U27754 (N_27754,N_27347,N_27295);
nand U27755 (N_27755,N_27470,N_27098);
nor U27756 (N_27756,N_27201,N_27160);
nor U27757 (N_27757,N_27453,N_27311);
xor U27758 (N_27758,N_27143,N_27050);
or U27759 (N_27759,N_27022,N_27413);
and U27760 (N_27760,N_27266,N_27451);
nor U27761 (N_27761,N_27053,N_27084);
xnor U27762 (N_27762,N_27116,N_27412);
nor U27763 (N_27763,N_27295,N_27439);
nand U27764 (N_27764,N_27438,N_27211);
xor U27765 (N_27765,N_27140,N_27490);
and U27766 (N_27766,N_27422,N_27185);
nand U27767 (N_27767,N_27207,N_27187);
nor U27768 (N_27768,N_27377,N_27193);
xnor U27769 (N_27769,N_27352,N_27097);
and U27770 (N_27770,N_27415,N_27366);
xor U27771 (N_27771,N_27143,N_27394);
xor U27772 (N_27772,N_27041,N_27293);
xor U27773 (N_27773,N_27296,N_27371);
and U27774 (N_27774,N_27381,N_27431);
xor U27775 (N_27775,N_27290,N_27235);
nor U27776 (N_27776,N_27483,N_27065);
or U27777 (N_27777,N_27125,N_27196);
nor U27778 (N_27778,N_27177,N_27358);
and U27779 (N_27779,N_27422,N_27346);
nand U27780 (N_27780,N_27229,N_27448);
xor U27781 (N_27781,N_27020,N_27426);
or U27782 (N_27782,N_27472,N_27178);
and U27783 (N_27783,N_27073,N_27425);
xor U27784 (N_27784,N_27265,N_27190);
or U27785 (N_27785,N_27443,N_27315);
and U27786 (N_27786,N_27107,N_27318);
xnor U27787 (N_27787,N_27330,N_27341);
xor U27788 (N_27788,N_27251,N_27032);
xor U27789 (N_27789,N_27443,N_27235);
and U27790 (N_27790,N_27043,N_27381);
nor U27791 (N_27791,N_27038,N_27401);
nand U27792 (N_27792,N_27040,N_27165);
or U27793 (N_27793,N_27289,N_27414);
xor U27794 (N_27794,N_27375,N_27472);
nor U27795 (N_27795,N_27059,N_27057);
and U27796 (N_27796,N_27388,N_27369);
xnor U27797 (N_27797,N_27434,N_27470);
nor U27798 (N_27798,N_27256,N_27401);
or U27799 (N_27799,N_27084,N_27057);
xnor U27800 (N_27800,N_27222,N_27429);
nor U27801 (N_27801,N_27130,N_27376);
or U27802 (N_27802,N_27129,N_27076);
or U27803 (N_27803,N_27267,N_27022);
nor U27804 (N_27804,N_27443,N_27088);
nor U27805 (N_27805,N_27192,N_27039);
nor U27806 (N_27806,N_27247,N_27119);
nor U27807 (N_27807,N_27028,N_27309);
xnor U27808 (N_27808,N_27317,N_27366);
or U27809 (N_27809,N_27289,N_27439);
nor U27810 (N_27810,N_27433,N_27136);
xnor U27811 (N_27811,N_27450,N_27143);
xor U27812 (N_27812,N_27493,N_27311);
nor U27813 (N_27813,N_27122,N_27326);
xnor U27814 (N_27814,N_27434,N_27411);
nor U27815 (N_27815,N_27269,N_27067);
xor U27816 (N_27816,N_27055,N_27238);
or U27817 (N_27817,N_27176,N_27317);
nor U27818 (N_27818,N_27488,N_27477);
nor U27819 (N_27819,N_27174,N_27498);
or U27820 (N_27820,N_27416,N_27113);
nand U27821 (N_27821,N_27077,N_27138);
or U27822 (N_27822,N_27481,N_27344);
nand U27823 (N_27823,N_27458,N_27131);
xor U27824 (N_27824,N_27479,N_27445);
nor U27825 (N_27825,N_27325,N_27029);
or U27826 (N_27826,N_27367,N_27456);
nor U27827 (N_27827,N_27041,N_27464);
nand U27828 (N_27828,N_27260,N_27324);
or U27829 (N_27829,N_27022,N_27177);
or U27830 (N_27830,N_27338,N_27484);
xnor U27831 (N_27831,N_27226,N_27294);
and U27832 (N_27832,N_27056,N_27403);
and U27833 (N_27833,N_27313,N_27086);
xor U27834 (N_27834,N_27038,N_27152);
or U27835 (N_27835,N_27490,N_27328);
or U27836 (N_27836,N_27453,N_27195);
nand U27837 (N_27837,N_27479,N_27158);
and U27838 (N_27838,N_27078,N_27394);
nor U27839 (N_27839,N_27304,N_27443);
or U27840 (N_27840,N_27266,N_27202);
nor U27841 (N_27841,N_27168,N_27386);
xor U27842 (N_27842,N_27224,N_27223);
nand U27843 (N_27843,N_27057,N_27455);
nand U27844 (N_27844,N_27202,N_27262);
nor U27845 (N_27845,N_27063,N_27175);
xnor U27846 (N_27846,N_27485,N_27158);
and U27847 (N_27847,N_27303,N_27432);
nor U27848 (N_27848,N_27115,N_27075);
xnor U27849 (N_27849,N_27248,N_27053);
or U27850 (N_27850,N_27339,N_27115);
xnor U27851 (N_27851,N_27038,N_27157);
and U27852 (N_27852,N_27117,N_27440);
xor U27853 (N_27853,N_27007,N_27345);
or U27854 (N_27854,N_27464,N_27190);
nor U27855 (N_27855,N_27101,N_27470);
or U27856 (N_27856,N_27122,N_27421);
nor U27857 (N_27857,N_27065,N_27140);
xor U27858 (N_27858,N_27399,N_27110);
and U27859 (N_27859,N_27397,N_27146);
or U27860 (N_27860,N_27391,N_27161);
nand U27861 (N_27861,N_27168,N_27187);
and U27862 (N_27862,N_27414,N_27431);
xnor U27863 (N_27863,N_27451,N_27051);
nand U27864 (N_27864,N_27204,N_27369);
xor U27865 (N_27865,N_27042,N_27418);
nor U27866 (N_27866,N_27123,N_27497);
xor U27867 (N_27867,N_27017,N_27234);
and U27868 (N_27868,N_27303,N_27333);
xnor U27869 (N_27869,N_27292,N_27260);
or U27870 (N_27870,N_27388,N_27360);
and U27871 (N_27871,N_27489,N_27159);
or U27872 (N_27872,N_27372,N_27390);
nand U27873 (N_27873,N_27053,N_27114);
nor U27874 (N_27874,N_27408,N_27138);
xor U27875 (N_27875,N_27451,N_27123);
nand U27876 (N_27876,N_27424,N_27051);
or U27877 (N_27877,N_27054,N_27202);
or U27878 (N_27878,N_27474,N_27483);
xnor U27879 (N_27879,N_27355,N_27037);
nand U27880 (N_27880,N_27469,N_27292);
nor U27881 (N_27881,N_27234,N_27097);
nor U27882 (N_27882,N_27152,N_27082);
and U27883 (N_27883,N_27273,N_27200);
nor U27884 (N_27884,N_27482,N_27090);
nor U27885 (N_27885,N_27119,N_27376);
or U27886 (N_27886,N_27105,N_27246);
or U27887 (N_27887,N_27154,N_27106);
and U27888 (N_27888,N_27264,N_27416);
and U27889 (N_27889,N_27477,N_27229);
and U27890 (N_27890,N_27038,N_27092);
and U27891 (N_27891,N_27131,N_27159);
nor U27892 (N_27892,N_27493,N_27125);
nor U27893 (N_27893,N_27262,N_27253);
nand U27894 (N_27894,N_27275,N_27305);
and U27895 (N_27895,N_27366,N_27381);
xor U27896 (N_27896,N_27069,N_27152);
and U27897 (N_27897,N_27338,N_27016);
xnor U27898 (N_27898,N_27431,N_27172);
nor U27899 (N_27899,N_27261,N_27002);
or U27900 (N_27900,N_27294,N_27423);
nor U27901 (N_27901,N_27379,N_27435);
nor U27902 (N_27902,N_27073,N_27458);
nor U27903 (N_27903,N_27000,N_27130);
nand U27904 (N_27904,N_27073,N_27352);
or U27905 (N_27905,N_27343,N_27311);
xor U27906 (N_27906,N_27134,N_27337);
nand U27907 (N_27907,N_27060,N_27088);
nor U27908 (N_27908,N_27036,N_27060);
nand U27909 (N_27909,N_27268,N_27166);
xor U27910 (N_27910,N_27458,N_27359);
nor U27911 (N_27911,N_27067,N_27456);
nor U27912 (N_27912,N_27471,N_27333);
or U27913 (N_27913,N_27021,N_27248);
and U27914 (N_27914,N_27182,N_27467);
and U27915 (N_27915,N_27148,N_27294);
nand U27916 (N_27916,N_27113,N_27255);
nand U27917 (N_27917,N_27017,N_27268);
and U27918 (N_27918,N_27430,N_27118);
xnor U27919 (N_27919,N_27420,N_27218);
and U27920 (N_27920,N_27106,N_27355);
nor U27921 (N_27921,N_27084,N_27322);
and U27922 (N_27922,N_27251,N_27495);
xor U27923 (N_27923,N_27131,N_27182);
nor U27924 (N_27924,N_27084,N_27294);
nor U27925 (N_27925,N_27228,N_27499);
and U27926 (N_27926,N_27069,N_27415);
and U27927 (N_27927,N_27433,N_27088);
xor U27928 (N_27928,N_27146,N_27040);
xnor U27929 (N_27929,N_27495,N_27306);
and U27930 (N_27930,N_27123,N_27060);
nor U27931 (N_27931,N_27419,N_27304);
or U27932 (N_27932,N_27457,N_27448);
xor U27933 (N_27933,N_27312,N_27162);
xnor U27934 (N_27934,N_27012,N_27050);
nand U27935 (N_27935,N_27154,N_27195);
nor U27936 (N_27936,N_27171,N_27315);
xnor U27937 (N_27937,N_27419,N_27198);
nor U27938 (N_27938,N_27428,N_27377);
or U27939 (N_27939,N_27472,N_27489);
xor U27940 (N_27940,N_27023,N_27447);
xnor U27941 (N_27941,N_27455,N_27194);
or U27942 (N_27942,N_27305,N_27256);
nor U27943 (N_27943,N_27001,N_27184);
and U27944 (N_27944,N_27163,N_27420);
or U27945 (N_27945,N_27301,N_27142);
nor U27946 (N_27946,N_27422,N_27450);
or U27947 (N_27947,N_27276,N_27055);
nor U27948 (N_27948,N_27307,N_27455);
nor U27949 (N_27949,N_27499,N_27316);
nor U27950 (N_27950,N_27369,N_27282);
nor U27951 (N_27951,N_27458,N_27424);
xor U27952 (N_27952,N_27022,N_27173);
xnor U27953 (N_27953,N_27362,N_27081);
and U27954 (N_27954,N_27380,N_27231);
nand U27955 (N_27955,N_27330,N_27123);
xor U27956 (N_27956,N_27043,N_27282);
or U27957 (N_27957,N_27173,N_27179);
nor U27958 (N_27958,N_27425,N_27105);
or U27959 (N_27959,N_27092,N_27407);
xor U27960 (N_27960,N_27382,N_27314);
nand U27961 (N_27961,N_27345,N_27217);
nor U27962 (N_27962,N_27468,N_27266);
or U27963 (N_27963,N_27271,N_27384);
nor U27964 (N_27964,N_27079,N_27407);
nor U27965 (N_27965,N_27101,N_27305);
and U27966 (N_27966,N_27496,N_27283);
and U27967 (N_27967,N_27443,N_27245);
or U27968 (N_27968,N_27346,N_27171);
nand U27969 (N_27969,N_27120,N_27042);
or U27970 (N_27970,N_27094,N_27496);
nor U27971 (N_27971,N_27142,N_27327);
xnor U27972 (N_27972,N_27160,N_27418);
xor U27973 (N_27973,N_27000,N_27241);
nand U27974 (N_27974,N_27061,N_27213);
nand U27975 (N_27975,N_27460,N_27092);
xnor U27976 (N_27976,N_27124,N_27438);
and U27977 (N_27977,N_27493,N_27452);
nor U27978 (N_27978,N_27466,N_27299);
xor U27979 (N_27979,N_27028,N_27044);
xnor U27980 (N_27980,N_27067,N_27295);
nor U27981 (N_27981,N_27121,N_27327);
xor U27982 (N_27982,N_27191,N_27013);
or U27983 (N_27983,N_27408,N_27160);
or U27984 (N_27984,N_27477,N_27193);
and U27985 (N_27985,N_27479,N_27459);
xnor U27986 (N_27986,N_27354,N_27132);
nor U27987 (N_27987,N_27261,N_27400);
or U27988 (N_27988,N_27385,N_27129);
nand U27989 (N_27989,N_27098,N_27009);
and U27990 (N_27990,N_27053,N_27475);
nor U27991 (N_27991,N_27203,N_27406);
nor U27992 (N_27992,N_27032,N_27091);
nor U27993 (N_27993,N_27234,N_27169);
nand U27994 (N_27994,N_27302,N_27021);
and U27995 (N_27995,N_27419,N_27314);
or U27996 (N_27996,N_27139,N_27276);
nand U27997 (N_27997,N_27190,N_27040);
and U27998 (N_27998,N_27043,N_27489);
xnor U27999 (N_27999,N_27114,N_27046);
and U28000 (N_28000,N_27611,N_27649);
nand U28001 (N_28001,N_27618,N_27853);
nor U28002 (N_28002,N_27986,N_27789);
xor U28003 (N_28003,N_27935,N_27578);
nand U28004 (N_28004,N_27912,N_27902);
or U28005 (N_28005,N_27849,N_27694);
xnor U28006 (N_28006,N_27996,N_27963);
nor U28007 (N_28007,N_27679,N_27857);
xnor U28008 (N_28008,N_27975,N_27998);
or U28009 (N_28009,N_27878,N_27620);
xor U28010 (N_28010,N_27943,N_27865);
nand U28011 (N_28011,N_27826,N_27641);
and U28012 (N_28012,N_27840,N_27901);
or U28013 (N_28013,N_27628,N_27724);
nor U28014 (N_28014,N_27900,N_27699);
nor U28015 (N_28015,N_27562,N_27794);
nor U28016 (N_28016,N_27719,N_27602);
nand U28017 (N_28017,N_27807,N_27927);
nor U28018 (N_28018,N_27730,N_27856);
xor U28019 (N_28019,N_27893,N_27868);
xnor U28020 (N_28020,N_27588,N_27973);
nor U28021 (N_28021,N_27877,N_27586);
xnor U28022 (N_28022,N_27775,N_27977);
or U28023 (N_28023,N_27928,N_27987);
or U28024 (N_28024,N_27929,N_27806);
nand U28025 (N_28025,N_27947,N_27674);
or U28026 (N_28026,N_27559,N_27945);
xor U28027 (N_28027,N_27659,N_27704);
xor U28028 (N_28028,N_27729,N_27899);
and U28029 (N_28029,N_27604,N_27999);
nand U28030 (N_28030,N_27887,N_27886);
nand U28031 (N_28031,N_27520,N_27869);
and U28032 (N_28032,N_27718,N_27573);
nor U28033 (N_28033,N_27872,N_27764);
and U28034 (N_28034,N_27832,N_27818);
and U28035 (N_28035,N_27725,N_27951);
xnor U28036 (N_28036,N_27521,N_27721);
or U28037 (N_28037,N_27985,N_27582);
nand U28038 (N_28038,N_27883,N_27515);
nand U28039 (N_28039,N_27739,N_27575);
and U28040 (N_28040,N_27979,N_27557);
nand U28041 (N_28041,N_27919,N_27926);
xnor U28042 (N_28042,N_27938,N_27599);
nand U28043 (N_28043,N_27579,N_27675);
nor U28044 (N_28044,N_27745,N_27770);
nor U28045 (N_28045,N_27668,N_27522);
nand U28046 (N_28046,N_27629,N_27792);
xor U28047 (N_28047,N_27847,N_27990);
or U28048 (N_28048,N_27690,N_27646);
nor U28049 (N_28049,N_27768,N_27648);
nand U28050 (N_28050,N_27633,N_27962);
or U28051 (N_28051,N_27655,N_27956);
xnor U28052 (N_28052,N_27665,N_27911);
nand U28053 (N_28053,N_27726,N_27898);
xor U28054 (N_28054,N_27795,N_27913);
nand U28055 (N_28055,N_27995,N_27639);
and U28056 (N_28056,N_27744,N_27953);
or U28057 (N_28057,N_27591,N_27761);
nor U28058 (N_28058,N_27689,N_27669);
nand U28059 (N_28059,N_27527,N_27903);
or U28060 (N_28060,N_27624,N_27643);
nand U28061 (N_28061,N_27677,N_27671);
nor U28062 (N_28062,N_27723,N_27703);
nand U28063 (N_28063,N_27771,N_27637);
and U28064 (N_28064,N_27613,N_27571);
nor U28065 (N_28065,N_27653,N_27574);
xnor U28066 (N_28066,N_27686,N_27692);
or U28067 (N_28067,N_27844,N_27933);
and U28068 (N_28068,N_27914,N_27596);
xor U28069 (N_28069,N_27747,N_27866);
nor U28070 (N_28070,N_27864,N_27946);
nor U28071 (N_28071,N_27576,N_27793);
xnor U28072 (N_28072,N_27528,N_27835);
xnor U28073 (N_28073,N_27988,N_27631);
or U28074 (N_28074,N_27852,N_27994);
and U28075 (N_28075,N_27532,N_27905);
or U28076 (N_28076,N_27693,N_27874);
or U28077 (N_28077,N_27920,N_27583);
nand U28078 (N_28078,N_27757,N_27592);
and U28079 (N_28079,N_27802,N_27625);
or U28080 (N_28080,N_27547,N_27682);
nor U28081 (N_28081,N_27627,N_27535);
or U28082 (N_28082,N_27955,N_27566);
nand U28083 (N_28083,N_27676,N_27507);
and U28084 (N_28084,N_27537,N_27940);
or U28085 (N_28085,N_27696,N_27650);
xor U28086 (N_28086,N_27801,N_27838);
and U28087 (N_28087,N_27720,N_27519);
nand U28088 (N_28088,N_27897,N_27969);
xnor U28089 (N_28089,N_27716,N_27743);
or U28090 (N_28090,N_27824,N_27984);
nor U28091 (N_28091,N_27701,N_27558);
nand U28092 (N_28092,N_27820,N_27673);
xor U28093 (N_28093,N_27584,N_27555);
xnor U28094 (N_28094,N_27711,N_27981);
and U28095 (N_28095,N_27556,N_27827);
nor U28096 (N_28096,N_27645,N_27552);
and U28097 (N_28097,N_27765,N_27731);
nor U28098 (N_28098,N_27608,N_27805);
or U28099 (N_28099,N_27722,N_27954);
or U28100 (N_28100,N_27589,N_27819);
or U28101 (N_28101,N_27959,N_27873);
or U28102 (N_28102,N_27958,N_27937);
and U28103 (N_28103,N_27569,N_27691);
nand U28104 (N_28104,N_27523,N_27880);
nor U28105 (N_28105,N_27760,N_27798);
nand U28106 (N_28106,N_27706,N_27755);
nand U28107 (N_28107,N_27910,N_27879);
nand U28108 (N_28108,N_27595,N_27504);
or U28109 (N_28109,N_27585,N_27543);
or U28110 (N_28110,N_27577,N_27567);
nand U28111 (N_28111,N_27823,N_27758);
or U28112 (N_28112,N_27505,N_27888);
nand U28113 (N_28113,N_27836,N_27550);
nand U28114 (N_28114,N_27825,N_27784);
or U28115 (N_28115,N_27967,N_27767);
and U28116 (N_28116,N_27681,N_27907);
or U28117 (N_28117,N_27728,N_27949);
and U28118 (N_28118,N_27525,N_27785);
nand U28119 (N_28119,N_27517,N_27607);
nor U28120 (N_28120,N_27672,N_27980);
nor U28121 (N_28121,N_27597,N_27786);
nand U28122 (N_28122,N_27749,N_27909);
nand U28123 (N_28123,N_27713,N_27509);
nor U28124 (N_28124,N_27539,N_27572);
xnor U28125 (N_28125,N_27875,N_27941);
and U28126 (N_28126,N_27850,N_27553);
xnor U28127 (N_28127,N_27960,N_27833);
xor U28128 (N_28128,N_27972,N_27791);
nor U28129 (N_28129,N_27670,N_27930);
nor U28130 (N_28130,N_27735,N_27830);
or U28131 (N_28131,N_27862,N_27983);
nand U28132 (N_28132,N_27892,N_27514);
xor U28133 (N_28133,N_27621,N_27797);
or U28134 (N_28134,N_27828,N_27727);
xor U28135 (N_28135,N_27976,N_27516);
xor U28136 (N_28136,N_27750,N_27753);
xnor U28137 (N_28137,N_27709,N_27506);
nor U28138 (N_28138,N_27740,N_27815);
or U28139 (N_28139,N_27982,N_27964);
and U28140 (N_28140,N_27950,N_27863);
and U28141 (N_28141,N_27781,N_27560);
nor U28142 (N_28142,N_27884,N_27551);
nor U28143 (N_28143,N_27776,N_27876);
and U28144 (N_28144,N_27510,N_27657);
xor U28145 (N_28145,N_27598,N_27546);
xnor U28146 (N_28146,N_27891,N_27752);
and U28147 (N_28147,N_27896,N_27808);
or U28148 (N_28148,N_27921,N_27993);
nand U28149 (N_28149,N_27904,N_27822);
and U28150 (N_28150,N_27568,N_27617);
or U28151 (N_28151,N_27895,N_27695);
and U28152 (N_28152,N_27630,N_27778);
xnor U28153 (N_28153,N_27906,N_27541);
or U28154 (N_28154,N_27881,N_27997);
xor U28155 (N_28155,N_27612,N_27774);
nand U28156 (N_28156,N_27626,N_27647);
nand U28157 (N_28157,N_27859,N_27564);
and U28158 (N_28158,N_27738,N_27654);
and U28159 (N_28159,N_27762,N_27530);
nand U28160 (N_28160,N_27683,N_27609);
or U28161 (N_28161,N_27538,N_27549);
and U28162 (N_28162,N_27652,N_27748);
and U28163 (N_28163,N_27531,N_27780);
or U28164 (N_28164,N_27788,N_27890);
xor U28165 (N_28165,N_27800,N_27871);
nor U28166 (N_28166,N_27702,N_27763);
nor U28167 (N_28167,N_27534,N_27717);
and U28168 (N_28168,N_27736,N_27854);
or U28169 (N_28169,N_27922,N_27831);
nand U28170 (N_28170,N_27799,N_27554);
xor U28171 (N_28171,N_27772,N_27644);
nor U28172 (N_28172,N_27614,N_27974);
nand U28173 (N_28173,N_27870,N_27658);
nor U28174 (N_28174,N_27513,N_27754);
nor U28175 (N_28175,N_27687,N_27812);
nor U28176 (N_28176,N_27751,N_27606);
nor U28177 (N_28177,N_27587,N_27769);
nand U28178 (N_28178,N_27846,N_27500);
xor U28179 (N_28179,N_27732,N_27707);
xor U28180 (N_28180,N_27581,N_27845);
xor U28181 (N_28181,N_27680,N_27684);
xnor U28182 (N_28182,N_27518,N_27779);
or U28183 (N_28183,N_27660,N_27968);
nor U28184 (N_28184,N_27783,N_27851);
or U28185 (N_28185,N_27508,N_27966);
xor U28186 (N_28186,N_27685,N_27715);
or U28187 (N_28187,N_27813,N_27834);
or U28188 (N_28188,N_27924,N_27811);
nor U28189 (N_28189,N_27616,N_27512);
xnor U28190 (N_28190,N_27570,N_27855);
xnor U28191 (N_28191,N_27734,N_27741);
or U28192 (N_28192,N_27841,N_27957);
xor U28193 (N_28193,N_27858,N_27536);
and U28194 (N_28194,N_27961,N_27894);
nand U28195 (N_28195,N_27638,N_27756);
xnor U28196 (N_28196,N_27803,N_27563);
or U28197 (N_28197,N_27601,N_27810);
nand U28198 (N_28198,N_27839,N_27932);
or U28199 (N_28199,N_27593,N_27759);
or U28200 (N_28200,N_27544,N_27837);
or U28201 (N_28201,N_27622,N_27916);
xor U28202 (N_28202,N_27942,N_27662);
nor U28203 (N_28203,N_27545,N_27978);
or U28204 (N_28204,N_27842,N_27636);
or U28205 (N_28205,N_27918,N_27971);
and U28206 (N_28206,N_27817,N_27540);
or U28207 (N_28207,N_27925,N_27708);
or U28208 (N_28208,N_27623,N_27989);
nor U28209 (N_28209,N_27948,N_27816);
nand U28210 (N_28210,N_27533,N_27733);
nand U28211 (N_28211,N_27700,N_27923);
and U28212 (N_28212,N_27889,N_27640);
nand U28213 (N_28213,N_27790,N_27787);
and U28214 (N_28214,N_27712,N_27663);
or U28215 (N_28215,N_27908,N_27777);
and U28216 (N_28216,N_27632,N_27524);
nand U28217 (N_28217,N_27580,N_27590);
and U28218 (N_28218,N_27773,N_27529);
and U28219 (N_28219,N_27697,N_27698);
and U28220 (N_28220,N_27542,N_27661);
and U28221 (N_28221,N_27934,N_27511);
xnor U28222 (N_28222,N_27634,N_27917);
xnor U28223 (N_28223,N_27861,N_27678);
xnor U28224 (N_28224,N_27561,N_27970);
nand U28225 (N_28225,N_27502,N_27666);
nor U28226 (N_28226,N_27600,N_27991);
or U28227 (N_28227,N_27848,N_27882);
nand U28228 (N_28228,N_27656,N_27526);
xor U28229 (N_28229,N_27915,N_27809);
or U28230 (N_28230,N_27885,N_27501);
nor U28231 (N_28231,N_27635,N_27944);
and U28232 (N_28232,N_27610,N_27737);
xor U28233 (N_28233,N_27936,N_27952);
and U28234 (N_28234,N_27548,N_27503);
xor U28235 (N_28235,N_27821,N_27664);
nand U28236 (N_28236,N_27931,N_27710);
and U28237 (N_28237,N_27605,N_27867);
nand U28238 (N_28238,N_27782,N_27814);
xor U28239 (N_28239,N_27619,N_27843);
nor U28240 (N_28240,N_27766,N_27603);
nor U28241 (N_28241,N_27642,N_27565);
or U28242 (N_28242,N_27804,N_27992);
and U28243 (N_28243,N_27860,N_27796);
nor U28244 (N_28244,N_27742,N_27746);
nand U28245 (N_28245,N_27615,N_27939);
nor U28246 (N_28246,N_27965,N_27688);
xnor U28247 (N_28247,N_27829,N_27651);
and U28248 (N_28248,N_27705,N_27714);
nand U28249 (N_28249,N_27667,N_27594);
nor U28250 (N_28250,N_27695,N_27609);
or U28251 (N_28251,N_27559,N_27626);
nand U28252 (N_28252,N_27998,N_27635);
or U28253 (N_28253,N_27528,N_27778);
or U28254 (N_28254,N_27814,N_27500);
xor U28255 (N_28255,N_27944,N_27610);
nor U28256 (N_28256,N_27609,N_27503);
xnor U28257 (N_28257,N_27768,N_27742);
or U28258 (N_28258,N_27972,N_27636);
and U28259 (N_28259,N_27674,N_27788);
xnor U28260 (N_28260,N_27827,N_27701);
and U28261 (N_28261,N_27965,N_27715);
nand U28262 (N_28262,N_27521,N_27781);
and U28263 (N_28263,N_27673,N_27954);
and U28264 (N_28264,N_27854,N_27652);
xor U28265 (N_28265,N_27612,N_27674);
or U28266 (N_28266,N_27704,N_27983);
xor U28267 (N_28267,N_27936,N_27695);
and U28268 (N_28268,N_27975,N_27759);
nand U28269 (N_28269,N_27696,N_27977);
xnor U28270 (N_28270,N_27915,N_27558);
and U28271 (N_28271,N_27882,N_27791);
nand U28272 (N_28272,N_27580,N_27642);
nand U28273 (N_28273,N_27644,N_27747);
nor U28274 (N_28274,N_27567,N_27807);
and U28275 (N_28275,N_27825,N_27794);
and U28276 (N_28276,N_27760,N_27657);
xor U28277 (N_28277,N_27619,N_27552);
nand U28278 (N_28278,N_27570,N_27945);
nor U28279 (N_28279,N_27959,N_27891);
nand U28280 (N_28280,N_27735,N_27833);
nand U28281 (N_28281,N_27601,N_27557);
nand U28282 (N_28282,N_27676,N_27532);
or U28283 (N_28283,N_27698,N_27871);
nor U28284 (N_28284,N_27966,N_27833);
xnor U28285 (N_28285,N_27741,N_27620);
or U28286 (N_28286,N_27594,N_27950);
nor U28287 (N_28287,N_27771,N_27990);
nor U28288 (N_28288,N_27677,N_27734);
or U28289 (N_28289,N_27534,N_27770);
or U28290 (N_28290,N_27842,N_27873);
and U28291 (N_28291,N_27774,N_27561);
nand U28292 (N_28292,N_27755,N_27777);
and U28293 (N_28293,N_27552,N_27994);
xnor U28294 (N_28294,N_27875,N_27861);
nand U28295 (N_28295,N_27858,N_27903);
nand U28296 (N_28296,N_27573,N_27757);
and U28297 (N_28297,N_27812,N_27564);
or U28298 (N_28298,N_27581,N_27763);
and U28299 (N_28299,N_27775,N_27802);
nand U28300 (N_28300,N_27551,N_27857);
or U28301 (N_28301,N_27502,N_27789);
nor U28302 (N_28302,N_27952,N_27732);
or U28303 (N_28303,N_27700,N_27674);
or U28304 (N_28304,N_27619,N_27963);
nor U28305 (N_28305,N_27821,N_27654);
nor U28306 (N_28306,N_27861,N_27574);
nand U28307 (N_28307,N_27753,N_27997);
nor U28308 (N_28308,N_27584,N_27926);
nor U28309 (N_28309,N_27980,N_27983);
and U28310 (N_28310,N_27874,N_27526);
nor U28311 (N_28311,N_27993,N_27829);
xor U28312 (N_28312,N_27649,N_27677);
nor U28313 (N_28313,N_27529,N_27809);
nand U28314 (N_28314,N_27593,N_27512);
and U28315 (N_28315,N_27681,N_27577);
nand U28316 (N_28316,N_27558,N_27710);
xor U28317 (N_28317,N_27616,N_27733);
nor U28318 (N_28318,N_27545,N_27719);
xnor U28319 (N_28319,N_27681,N_27882);
nor U28320 (N_28320,N_27711,N_27556);
xnor U28321 (N_28321,N_27801,N_27761);
nand U28322 (N_28322,N_27603,N_27622);
or U28323 (N_28323,N_27780,N_27863);
xnor U28324 (N_28324,N_27721,N_27982);
nand U28325 (N_28325,N_27890,N_27645);
or U28326 (N_28326,N_27727,N_27627);
nand U28327 (N_28327,N_27860,N_27868);
xnor U28328 (N_28328,N_27928,N_27983);
nand U28329 (N_28329,N_27852,N_27920);
or U28330 (N_28330,N_27554,N_27681);
nor U28331 (N_28331,N_27572,N_27892);
nand U28332 (N_28332,N_27683,N_27652);
xnor U28333 (N_28333,N_27952,N_27546);
nor U28334 (N_28334,N_27730,N_27524);
nor U28335 (N_28335,N_27741,N_27660);
nor U28336 (N_28336,N_27560,N_27989);
xnor U28337 (N_28337,N_27707,N_27608);
or U28338 (N_28338,N_27569,N_27800);
nor U28339 (N_28339,N_27513,N_27659);
nand U28340 (N_28340,N_27555,N_27843);
and U28341 (N_28341,N_27759,N_27855);
or U28342 (N_28342,N_27624,N_27871);
nor U28343 (N_28343,N_27780,N_27886);
and U28344 (N_28344,N_27825,N_27734);
nor U28345 (N_28345,N_27828,N_27627);
xnor U28346 (N_28346,N_27733,N_27637);
nor U28347 (N_28347,N_27930,N_27872);
xor U28348 (N_28348,N_27755,N_27649);
nand U28349 (N_28349,N_27599,N_27868);
or U28350 (N_28350,N_27731,N_27975);
nor U28351 (N_28351,N_27791,N_27676);
nand U28352 (N_28352,N_27669,N_27773);
or U28353 (N_28353,N_27963,N_27523);
or U28354 (N_28354,N_27912,N_27965);
or U28355 (N_28355,N_27628,N_27872);
nand U28356 (N_28356,N_27890,N_27726);
nor U28357 (N_28357,N_27734,N_27785);
xor U28358 (N_28358,N_27724,N_27814);
and U28359 (N_28359,N_27921,N_27757);
nand U28360 (N_28360,N_27782,N_27578);
nor U28361 (N_28361,N_27931,N_27537);
nand U28362 (N_28362,N_27956,N_27941);
nor U28363 (N_28363,N_27734,N_27577);
or U28364 (N_28364,N_27585,N_27638);
nand U28365 (N_28365,N_27796,N_27878);
nor U28366 (N_28366,N_27705,N_27685);
xor U28367 (N_28367,N_27750,N_27514);
nand U28368 (N_28368,N_27843,N_27635);
nand U28369 (N_28369,N_27545,N_27838);
xnor U28370 (N_28370,N_27620,N_27875);
xor U28371 (N_28371,N_27827,N_27906);
nand U28372 (N_28372,N_27807,N_27951);
and U28373 (N_28373,N_27500,N_27752);
or U28374 (N_28374,N_27656,N_27654);
xor U28375 (N_28375,N_27940,N_27669);
or U28376 (N_28376,N_27967,N_27823);
xnor U28377 (N_28377,N_27544,N_27537);
nor U28378 (N_28378,N_27584,N_27844);
and U28379 (N_28379,N_27604,N_27730);
or U28380 (N_28380,N_27659,N_27668);
nor U28381 (N_28381,N_27504,N_27570);
or U28382 (N_28382,N_27986,N_27610);
xnor U28383 (N_28383,N_27950,N_27768);
nand U28384 (N_28384,N_27819,N_27918);
and U28385 (N_28385,N_27777,N_27617);
or U28386 (N_28386,N_27944,N_27963);
or U28387 (N_28387,N_27560,N_27524);
nand U28388 (N_28388,N_27895,N_27580);
nand U28389 (N_28389,N_27704,N_27852);
and U28390 (N_28390,N_27886,N_27762);
xor U28391 (N_28391,N_27745,N_27557);
nand U28392 (N_28392,N_27623,N_27724);
nand U28393 (N_28393,N_27597,N_27575);
or U28394 (N_28394,N_27568,N_27673);
nor U28395 (N_28395,N_27500,N_27574);
or U28396 (N_28396,N_27783,N_27617);
xor U28397 (N_28397,N_27773,N_27594);
nand U28398 (N_28398,N_27660,N_27970);
or U28399 (N_28399,N_27847,N_27601);
nor U28400 (N_28400,N_27662,N_27548);
nor U28401 (N_28401,N_27910,N_27729);
nand U28402 (N_28402,N_27615,N_27502);
and U28403 (N_28403,N_27515,N_27668);
nand U28404 (N_28404,N_27561,N_27714);
and U28405 (N_28405,N_27798,N_27924);
nor U28406 (N_28406,N_27751,N_27580);
nand U28407 (N_28407,N_27683,N_27627);
or U28408 (N_28408,N_27982,N_27841);
nor U28409 (N_28409,N_27851,N_27860);
or U28410 (N_28410,N_27865,N_27573);
or U28411 (N_28411,N_27744,N_27668);
nand U28412 (N_28412,N_27519,N_27919);
nor U28413 (N_28413,N_27543,N_27689);
and U28414 (N_28414,N_27649,N_27990);
nand U28415 (N_28415,N_27526,N_27981);
or U28416 (N_28416,N_27773,N_27940);
xor U28417 (N_28417,N_27637,N_27983);
xor U28418 (N_28418,N_27837,N_27730);
nor U28419 (N_28419,N_27508,N_27544);
and U28420 (N_28420,N_27925,N_27891);
xor U28421 (N_28421,N_27878,N_27937);
or U28422 (N_28422,N_27980,N_27538);
and U28423 (N_28423,N_27644,N_27902);
or U28424 (N_28424,N_27715,N_27764);
xnor U28425 (N_28425,N_27500,N_27729);
xor U28426 (N_28426,N_27924,N_27834);
xnor U28427 (N_28427,N_27911,N_27513);
nor U28428 (N_28428,N_27592,N_27994);
nor U28429 (N_28429,N_27617,N_27594);
nor U28430 (N_28430,N_27687,N_27952);
and U28431 (N_28431,N_27584,N_27700);
nor U28432 (N_28432,N_27729,N_27633);
nor U28433 (N_28433,N_27627,N_27780);
nand U28434 (N_28434,N_27777,N_27938);
or U28435 (N_28435,N_27796,N_27564);
nand U28436 (N_28436,N_27528,N_27555);
nor U28437 (N_28437,N_27576,N_27748);
nand U28438 (N_28438,N_27865,N_27554);
xnor U28439 (N_28439,N_27831,N_27845);
or U28440 (N_28440,N_27890,N_27629);
nand U28441 (N_28441,N_27669,N_27667);
nand U28442 (N_28442,N_27618,N_27557);
or U28443 (N_28443,N_27881,N_27651);
and U28444 (N_28444,N_27605,N_27866);
and U28445 (N_28445,N_27788,N_27979);
or U28446 (N_28446,N_27733,N_27662);
nand U28447 (N_28447,N_27597,N_27984);
xnor U28448 (N_28448,N_27843,N_27659);
nor U28449 (N_28449,N_27641,N_27740);
xnor U28450 (N_28450,N_27665,N_27782);
nand U28451 (N_28451,N_27868,N_27567);
nor U28452 (N_28452,N_27870,N_27745);
nor U28453 (N_28453,N_27986,N_27585);
or U28454 (N_28454,N_27565,N_27800);
xor U28455 (N_28455,N_27714,N_27958);
nand U28456 (N_28456,N_27914,N_27630);
xnor U28457 (N_28457,N_27604,N_27922);
or U28458 (N_28458,N_27731,N_27565);
or U28459 (N_28459,N_27733,N_27642);
nand U28460 (N_28460,N_27977,N_27697);
xor U28461 (N_28461,N_27985,N_27998);
xor U28462 (N_28462,N_27682,N_27821);
xnor U28463 (N_28463,N_27927,N_27887);
or U28464 (N_28464,N_27674,N_27687);
nor U28465 (N_28465,N_27645,N_27610);
xor U28466 (N_28466,N_27928,N_27678);
or U28467 (N_28467,N_27897,N_27785);
and U28468 (N_28468,N_27969,N_27524);
or U28469 (N_28469,N_27568,N_27643);
nor U28470 (N_28470,N_27741,N_27910);
or U28471 (N_28471,N_27858,N_27833);
or U28472 (N_28472,N_27827,N_27696);
and U28473 (N_28473,N_27615,N_27709);
nor U28474 (N_28474,N_27746,N_27720);
nor U28475 (N_28475,N_27970,N_27540);
or U28476 (N_28476,N_27744,N_27764);
or U28477 (N_28477,N_27726,N_27539);
nand U28478 (N_28478,N_27964,N_27694);
or U28479 (N_28479,N_27977,N_27749);
or U28480 (N_28480,N_27804,N_27976);
nand U28481 (N_28481,N_27856,N_27960);
nor U28482 (N_28482,N_27639,N_27712);
or U28483 (N_28483,N_27641,N_27872);
or U28484 (N_28484,N_27550,N_27835);
xnor U28485 (N_28485,N_27830,N_27795);
nand U28486 (N_28486,N_27679,N_27553);
nor U28487 (N_28487,N_27939,N_27813);
and U28488 (N_28488,N_27910,N_27984);
xnor U28489 (N_28489,N_27874,N_27548);
nor U28490 (N_28490,N_27784,N_27590);
nor U28491 (N_28491,N_27973,N_27856);
or U28492 (N_28492,N_27501,N_27919);
xor U28493 (N_28493,N_27707,N_27658);
or U28494 (N_28494,N_27608,N_27641);
nand U28495 (N_28495,N_27760,N_27527);
and U28496 (N_28496,N_27980,N_27566);
and U28497 (N_28497,N_27894,N_27651);
or U28498 (N_28498,N_27824,N_27712);
nand U28499 (N_28499,N_27834,N_27641);
nand U28500 (N_28500,N_28444,N_28073);
nand U28501 (N_28501,N_28168,N_28325);
nor U28502 (N_28502,N_28180,N_28259);
or U28503 (N_28503,N_28334,N_28327);
and U28504 (N_28504,N_28297,N_28231);
nor U28505 (N_28505,N_28390,N_28447);
or U28506 (N_28506,N_28145,N_28497);
nor U28507 (N_28507,N_28378,N_28467);
nor U28508 (N_28508,N_28037,N_28372);
nand U28509 (N_28509,N_28186,N_28414);
and U28510 (N_28510,N_28094,N_28189);
nor U28511 (N_28511,N_28235,N_28382);
or U28512 (N_28512,N_28004,N_28140);
xnor U28513 (N_28513,N_28277,N_28193);
or U28514 (N_28514,N_28086,N_28465);
and U28515 (N_28515,N_28479,N_28198);
or U28516 (N_28516,N_28379,N_28085);
xnor U28517 (N_28517,N_28391,N_28351);
and U28518 (N_28518,N_28057,N_28438);
nand U28519 (N_28519,N_28044,N_28374);
or U28520 (N_28520,N_28412,N_28081);
nor U28521 (N_28521,N_28339,N_28187);
and U28522 (N_28522,N_28464,N_28255);
and U28523 (N_28523,N_28343,N_28029);
and U28524 (N_28524,N_28034,N_28436);
nand U28525 (N_28525,N_28495,N_28133);
nand U28526 (N_28526,N_28107,N_28370);
or U28527 (N_28527,N_28344,N_28319);
nand U28528 (N_28528,N_28405,N_28125);
or U28529 (N_28529,N_28216,N_28478);
or U28530 (N_28530,N_28234,N_28388);
nor U28531 (N_28531,N_28345,N_28045);
or U28532 (N_28532,N_28402,N_28361);
or U28533 (N_28533,N_28032,N_28244);
nor U28534 (N_28534,N_28445,N_28093);
and U28535 (N_28535,N_28191,N_28322);
or U28536 (N_28536,N_28063,N_28158);
xor U28537 (N_28537,N_28236,N_28272);
or U28538 (N_28538,N_28389,N_28279);
and U28539 (N_28539,N_28080,N_28395);
nand U28540 (N_28540,N_28157,N_28160);
nor U28541 (N_28541,N_28060,N_28172);
nand U28542 (N_28542,N_28058,N_28061);
nor U28543 (N_28543,N_28052,N_28323);
or U28544 (N_28544,N_28201,N_28330);
or U28545 (N_28545,N_28055,N_28408);
xnor U28546 (N_28546,N_28119,N_28011);
and U28547 (N_28547,N_28018,N_28290);
nand U28548 (N_28548,N_28102,N_28144);
xnor U28549 (N_28549,N_28371,N_28127);
or U28550 (N_28550,N_28417,N_28383);
nand U28551 (N_28551,N_28048,N_28240);
nor U28552 (N_28552,N_28273,N_28051);
xnor U28553 (N_28553,N_28104,N_28084);
nand U28554 (N_28554,N_28266,N_28305);
nor U28555 (N_28555,N_28298,N_28350);
nand U28556 (N_28556,N_28090,N_28369);
or U28557 (N_28557,N_28271,N_28488);
nand U28558 (N_28558,N_28178,N_28328);
nand U28559 (N_28559,N_28114,N_28132);
or U28560 (N_28560,N_28110,N_28439);
xor U28561 (N_28561,N_28142,N_28243);
or U28562 (N_28562,N_28059,N_28377);
and U28563 (N_28563,N_28095,N_28123);
xor U28564 (N_28564,N_28264,N_28027);
nand U28565 (N_28565,N_28237,N_28014);
nor U28566 (N_28566,N_28486,N_28311);
xor U28567 (N_28567,N_28270,N_28130);
or U28568 (N_28568,N_28484,N_28326);
or U28569 (N_28569,N_28353,N_28012);
and U28570 (N_28570,N_28210,N_28241);
nand U28571 (N_28571,N_28017,N_28111);
or U28572 (N_28572,N_28415,N_28253);
nand U28573 (N_28573,N_28219,N_28418);
or U28574 (N_28574,N_28005,N_28173);
and U28575 (N_28575,N_28190,N_28098);
or U28576 (N_28576,N_28366,N_28202);
nand U28577 (N_28577,N_28065,N_28092);
and U28578 (N_28578,N_28324,N_28352);
or U28579 (N_28579,N_28209,N_28170);
and U28580 (N_28580,N_28247,N_28089);
xnor U28581 (N_28581,N_28340,N_28028);
or U28582 (N_28582,N_28454,N_28437);
nand U28583 (N_28583,N_28069,N_28221);
nand U28584 (N_28584,N_28101,N_28149);
or U28585 (N_28585,N_28204,N_28078);
xnor U28586 (N_28586,N_28008,N_28200);
or U28587 (N_28587,N_28143,N_28076);
nand U28588 (N_28588,N_28376,N_28294);
or U28589 (N_28589,N_28498,N_28321);
or U28590 (N_28590,N_28346,N_28407);
nand U28591 (N_28591,N_28403,N_28152);
nor U28592 (N_28592,N_28238,N_28167);
nand U28593 (N_28593,N_28226,N_28232);
or U28594 (N_28594,N_28285,N_28473);
and U28595 (N_28595,N_28136,N_28485);
nor U28596 (N_28596,N_28349,N_28096);
xnor U28597 (N_28597,N_28135,N_28248);
xor U28598 (N_28598,N_28306,N_28450);
and U28599 (N_28599,N_28074,N_28062);
xor U28600 (N_28600,N_28254,N_28239);
nor U28601 (N_28601,N_28475,N_28159);
nor U28602 (N_28602,N_28064,N_28121);
nand U28603 (N_28603,N_28177,N_28206);
nand U28604 (N_28604,N_28457,N_28068);
nor U28605 (N_28605,N_28449,N_28263);
and U28606 (N_28606,N_28278,N_28338);
nor U28607 (N_28607,N_28000,N_28252);
xnor U28608 (N_28608,N_28406,N_28458);
and U28609 (N_28609,N_28205,N_28109);
nor U28610 (N_28610,N_28024,N_28033);
nand U28611 (N_28611,N_28286,N_28099);
and U28612 (N_28612,N_28357,N_28347);
nor U28613 (N_28613,N_28106,N_28077);
xnor U28614 (N_28614,N_28316,N_28223);
and U28615 (N_28615,N_28435,N_28208);
or U28616 (N_28616,N_28013,N_28215);
nand U28617 (N_28617,N_28268,N_28434);
nor U28618 (N_28618,N_28117,N_28171);
nor U28619 (N_28619,N_28476,N_28046);
nand U28620 (N_28620,N_28477,N_28282);
and U28621 (N_28621,N_28153,N_28303);
xnor U28622 (N_28622,N_28097,N_28214);
or U28623 (N_28623,N_28251,N_28296);
nand U28624 (N_28624,N_28066,N_28308);
xor U28625 (N_28625,N_28466,N_28267);
or U28626 (N_28626,N_28211,N_28203);
and U28627 (N_28627,N_28363,N_28246);
nand U28628 (N_28628,N_28329,N_28331);
and U28629 (N_28629,N_28228,N_28196);
or U28630 (N_28630,N_28360,N_28399);
nor U28631 (N_28631,N_28103,N_28281);
nor U28632 (N_28632,N_28015,N_28217);
nor U28633 (N_28633,N_28194,N_28087);
nor U28634 (N_28634,N_28075,N_28441);
nor U28635 (N_28635,N_28091,N_28367);
xor U28636 (N_28636,N_28003,N_28242);
xor U28637 (N_28637,N_28487,N_28460);
xnor U28638 (N_28638,N_28416,N_28482);
and U28639 (N_28639,N_28364,N_28494);
nand U28640 (N_28640,N_28373,N_28079);
nor U28641 (N_28641,N_28431,N_28227);
nand U28642 (N_28642,N_28425,N_28420);
nand U28643 (N_28643,N_28195,N_28258);
nor U28644 (N_28644,N_28129,N_28124);
xor U28645 (N_28645,N_28317,N_28164);
xnor U28646 (N_28646,N_28493,N_28468);
nand U28647 (N_28647,N_28197,N_28452);
and U28648 (N_28648,N_28222,N_28150);
and U28649 (N_28649,N_28146,N_28137);
nor U28650 (N_28650,N_28455,N_28175);
xor U28651 (N_28651,N_28312,N_28042);
xor U28652 (N_28652,N_28470,N_28120);
nor U28653 (N_28653,N_28362,N_28481);
nor U28654 (N_28654,N_28006,N_28451);
nand U28655 (N_28655,N_28397,N_28474);
nand U28656 (N_28656,N_28333,N_28499);
and U28657 (N_28657,N_28183,N_28304);
nand U28658 (N_28658,N_28380,N_28147);
or U28659 (N_28659,N_28365,N_28428);
nand U28660 (N_28660,N_28442,N_28315);
or U28661 (N_28661,N_28009,N_28161);
nand U28662 (N_28662,N_28448,N_28422);
or U28663 (N_28663,N_28260,N_28356);
xnor U28664 (N_28664,N_28088,N_28010);
and U28665 (N_28665,N_28100,N_28443);
and U28666 (N_28666,N_28404,N_28398);
nor U28667 (N_28667,N_28245,N_28386);
or U28668 (N_28668,N_28283,N_28050);
nor U28669 (N_28669,N_28348,N_28289);
and U28670 (N_28670,N_28256,N_28396);
or U28671 (N_28671,N_28313,N_28291);
nor U28672 (N_28672,N_28122,N_28047);
nand U28673 (N_28673,N_28413,N_28025);
or U28674 (N_28674,N_28026,N_28218);
xnor U28675 (N_28675,N_28141,N_28128);
xnor U28676 (N_28676,N_28426,N_28368);
nor U28677 (N_28677,N_28179,N_28411);
or U28678 (N_28678,N_28292,N_28393);
xor U28679 (N_28679,N_28118,N_28381);
and U28680 (N_28680,N_28355,N_28269);
xnor U28681 (N_28681,N_28049,N_28332);
xnor U28682 (N_28682,N_28036,N_28038);
or U28683 (N_28683,N_28020,N_28199);
xnor U28684 (N_28684,N_28139,N_28354);
and U28685 (N_28685,N_28113,N_28302);
and U28686 (N_28686,N_28001,N_28480);
nand U28687 (N_28687,N_28453,N_28056);
nor U28688 (N_28688,N_28156,N_28490);
and U28689 (N_28689,N_28023,N_28424);
nand U28690 (N_28690,N_28212,N_28284);
nand U28691 (N_28691,N_28358,N_28131);
nor U28692 (N_28692,N_28262,N_28463);
nor U28693 (N_28693,N_28423,N_28392);
nand U28694 (N_28694,N_28257,N_28421);
and U28695 (N_28695,N_28162,N_28151);
nor U28696 (N_28696,N_28039,N_28280);
or U28697 (N_28697,N_28213,N_28337);
xnor U28698 (N_28698,N_28320,N_28293);
and U28699 (N_28699,N_28394,N_28148);
and U28700 (N_28700,N_28072,N_28385);
nor U28701 (N_28701,N_28419,N_28375);
and U28702 (N_28702,N_28154,N_28318);
nor U28703 (N_28703,N_28054,N_28163);
or U28704 (N_28704,N_28207,N_28176);
nand U28705 (N_28705,N_28400,N_28166);
or U28706 (N_28706,N_28165,N_28030);
nor U28707 (N_28707,N_28261,N_28469);
nor U28708 (N_28708,N_28031,N_28192);
nor U28709 (N_28709,N_28105,N_28265);
nand U28710 (N_28710,N_28430,N_28115);
nor U28711 (N_28711,N_28188,N_28472);
nand U28712 (N_28712,N_28301,N_28300);
xnor U28713 (N_28713,N_28276,N_28310);
or U28714 (N_28714,N_28082,N_28410);
and U28715 (N_28715,N_28112,N_28335);
and U28716 (N_28716,N_28155,N_28288);
and U28717 (N_28717,N_28116,N_28174);
nor U28718 (N_28718,N_28040,N_28384);
or U28719 (N_28719,N_28307,N_28220);
xor U28720 (N_28720,N_28287,N_28336);
nand U28721 (N_28721,N_28409,N_28230);
xnor U28722 (N_28722,N_28432,N_28314);
and U28723 (N_28723,N_28083,N_28492);
xor U28724 (N_28724,N_28471,N_28440);
and U28725 (N_28725,N_28456,N_28070);
nor U28726 (N_28726,N_28007,N_28043);
and U28727 (N_28727,N_28489,N_28250);
nor U28728 (N_28728,N_28229,N_28169);
nor U28729 (N_28729,N_28462,N_28224);
or U28730 (N_28730,N_28401,N_28342);
or U28731 (N_28731,N_28067,N_28233);
nand U28732 (N_28732,N_28249,N_28071);
nand U28733 (N_28733,N_28035,N_28225);
xor U28734 (N_28734,N_28041,N_28459);
nor U28735 (N_28735,N_28274,N_28053);
nor U28736 (N_28736,N_28019,N_28309);
or U28737 (N_28737,N_28181,N_28496);
or U28738 (N_28738,N_28461,N_28433);
nand U28739 (N_28739,N_28295,N_28491);
and U28740 (N_28740,N_28108,N_28184);
nor U28741 (N_28741,N_28341,N_28185);
nand U28742 (N_28742,N_28275,N_28429);
nor U28743 (N_28743,N_28446,N_28359);
nor U28744 (N_28744,N_28299,N_28387);
xor U28745 (N_28745,N_28427,N_28002);
or U28746 (N_28746,N_28483,N_28021);
nand U28747 (N_28747,N_28138,N_28182);
xnor U28748 (N_28748,N_28134,N_28022);
nand U28749 (N_28749,N_28126,N_28016);
and U28750 (N_28750,N_28438,N_28129);
xnor U28751 (N_28751,N_28019,N_28357);
or U28752 (N_28752,N_28271,N_28071);
nor U28753 (N_28753,N_28341,N_28375);
and U28754 (N_28754,N_28011,N_28277);
nand U28755 (N_28755,N_28361,N_28050);
or U28756 (N_28756,N_28222,N_28232);
and U28757 (N_28757,N_28275,N_28237);
nor U28758 (N_28758,N_28293,N_28167);
nand U28759 (N_28759,N_28410,N_28491);
and U28760 (N_28760,N_28169,N_28377);
or U28761 (N_28761,N_28001,N_28391);
or U28762 (N_28762,N_28309,N_28355);
nor U28763 (N_28763,N_28433,N_28365);
and U28764 (N_28764,N_28056,N_28460);
nor U28765 (N_28765,N_28444,N_28330);
or U28766 (N_28766,N_28211,N_28255);
or U28767 (N_28767,N_28146,N_28221);
and U28768 (N_28768,N_28021,N_28217);
nand U28769 (N_28769,N_28148,N_28161);
or U28770 (N_28770,N_28329,N_28251);
nor U28771 (N_28771,N_28400,N_28342);
or U28772 (N_28772,N_28427,N_28439);
and U28773 (N_28773,N_28361,N_28096);
nor U28774 (N_28774,N_28418,N_28479);
xor U28775 (N_28775,N_28148,N_28396);
nand U28776 (N_28776,N_28370,N_28053);
or U28777 (N_28777,N_28142,N_28340);
xor U28778 (N_28778,N_28346,N_28241);
or U28779 (N_28779,N_28277,N_28233);
or U28780 (N_28780,N_28079,N_28048);
nor U28781 (N_28781,N_28473,N_28312);
or U28782 (N_28782,N_28475,N_28093);
and U28783 (N_28783,N_28010,N_28403);
or U28784 (N_28784,N_28211,N_28385);
and U28785 (N_28785,N_28169,N_28479);
nand U28786 (N_28786,N_28047,N_28070);
nand U28787 (N_28787,N_28394,N_28488);
or U28788 (N_28788,N_28077,N_28462);
and U28789 (N_28789,N_28388,N_28218);
or U28790 (N_28790,N_28080,N_28415);
xnor U28791 (N_28791,N_28081,N_28170);
nand U28792 (N_28792,N_28092,N_28467);
nor U28793 (N_28793,N_28318,N_28177);
nor U28794 (N_28794,N_28428,N_28143);
nor U28795 (N_28795,N_28374,N_28364);
and U28796 (N_28796,N_28235,N_28149);
and U28797 (N_28797,N_28111,N_28341);
xnor U28798 (N_28798,N_28178,N_28299);
or U28799 (N_28799,N_28114,N_28021);
or U28800 (N_28800,N_28268,N_28393);
nor U28801 (N_28801,N_28363,N_28178);
and U28802 (N_28802,N_28144,N_28090);
and U28803 (N_28803,N_28328,N_28110);
nor U28804 (N_28804,N_28418,N_28158);
nor U28805 (N_28805,N_28347,N_28264);
nor U28806 (N_28806,N_28119,N_28376);
and U28807 (N_28807,N_28481,N_28079);
nand U28808 (N_28808,N_28370,N_28438);
nor U28809 (N_28809,N_28125,N_28375);
nor U28810 (N_28810,N_28092,N_28338);
nand U28811 (N_28811,N_28370,N_28419);
nor U28812 (N_28812,N_28080,N_28305);
and U28813 (N_28813,N_28325,N_28496);
nor U28814 (N_28814,N_28331,N_28170);
or U28815 (N_28815,N_28428,N_28063);
nand U28816 (N_28816,N_28262,N_28144);
and U28817 (N_28817,N_28375,N_28149);
nand U28818 (N_28818,N_28278,N_28121);
nor U28819 (N_28819,N_28115,N_28442);
nor U28820 (N_28820,N_28005,N_28019);
or U28821 (N_28821,N_28479,N_28249);
or U28822 (N_28822,N_28212,N_28352);
xor U28823 (N_28823,N_28076,N_28492);
xnor U28824 (N_28824,N_28377,N_28443);
or U28825 (N_28825,N_28277,N_28137);
nor U28826 (N_28826,N_28185,N_28058);
xor U28827 (N_28827,N_28276,N_28163);
xnor U28828 (N_28828,N_28373,N_28092);
xor U28829 (N_28829,N_28076,N_28194);
and U28830 (N_28830,N_28459,N_28152);
or U28831 (N_28831,N_28306,N_28384);
nor U28832 (N_28832,N_28335,N_28163);
nand U28833 (N_28833,N_28406,N_28288);
nor U28834 (N_28834,N_28211,N_28233);
xnor U28835 (N_28835,N_28362,N_28405);
nand U28836 (N_28836,N_28376,N_28404);
xnor U28837 (N_28837,N_28214,N_28161);
and U28838 (N_28838,N_28423,N_28015);
xor U28839 (N_28839,N_28113,N_28102);
nand U28840 (N_28840,N_28060,N_28486);
nand U28841 (N_28841,N_28453,N_28341);
nand U28842 (N_28842,N_28083,N_28279);
nand U28843 (N_28843,N_28339,N_28346);
or U28844 (N_28844,N_28201,N_28100);
nor U28845 (N_28845,N_28045,N_28076);
and U28846 (N_28846,N_28253,N_28120);
and U28847 (N_28847,N_28021,N_28490);
or U28848 (N_28848,N_28489,N_28020);
or U28849 (N_28849,N_28445,N_28091);
xnor U28850 (N_28850,N_28150,N_28250);
or U28851 (N_28851,N_28416,N_28078);
xor U28852 (N_28852,N_28458,N_28279);
xor U28853 (N_28853,N_28481,N_28392);
nor U28854 (N_28854,N_28075,N_28108);
or U28855 (N_28855,N_28216,N_28218);
or U28856 (N_28856,N_28366,N_28068);
xnor U28857 (N_28857,N_28273,N_28070);
xnor U28858 (N_28858,N_28236,N_28116);
and U28859 (N_28859,N_28184,N_28360);
or U28860 (N_28860,N_28104,N_28213);
and U28861 (N_28861,N_28061,N_28089);
and U28862 (N_28862,N_28223,N_28295);
xor U28863 (N_28863,N_28097,N_28100);
or U28864 (N_28864,N_28128,N_28244);
nand U28865 (N_28865,N_28475,N_28137);
and U28866 (N_28866,N_28252,N_28323);
xor U28867 (N_28867,N_28271,N_28403);
nand U28868 (N_28868,N_28174,N_28323);
xnor U28869 (N_28869,N_28215,N_28143);
or U28870 (N_28870,N_28305,N_28384);
nor U28871 (N_28871,N_28496,N_28089);
nand U28872 (N_28872,N_28003,N_28020);
or U28873 (N_28873,N_28009,N_28096);
and U28874 (N_28874,N_28306,N_28128);
or U28875 (N_28875,N_28130,N_28263);
or U28876 (N_28876,N_28168,N_28305);
and U28877 (N_28877,N_28006,N_28437);
nor U28878 (N_28878,N_28058,N_28194);
and U28879 (N_28879,N_28001,N_28298);
and U28880 (N_28880,N_28111,N_28261);
or U28881 (N_28881,N_28158,N_28482);
or U28882 (N_28882,N_28066,N_28239);
xor U28883 (N_28883,N_28049,N_28353);
nand U28884 (N_28884,N_28189,N_28111);
and U28885 (N_28885,N_28416,N_28202);
or U28886 (N_28886,N_28326,N_28242);
and U28887 (N_28887,N_28480,N_28439);
nand U28888 (N_28888,N_28334,N_28203);
and U28889 (N_28889,N_28381,N_28189);
xor U28890 (N_28890,N_28022,N_28098);
nor U28891 (N_28891,N_28439,N_28380);
or U28892 (N_28892,N_28374,N_28086);
or U28893 (N_28893,N_28326,N_28026);
nor U28894 (N_28894,N_28177,N_28148);
xnor U28895 (N_28895,N_28274,N_28253);
or U28896 (N_28896,N_28060,N_28478);
and U28897 (N_28897,N_28074,N_28278);
or U28898 (N_28898,N_28300,N_28413);
xnor U28899 (N_28899,N_28394,N_28078);
nand U28900 (N_28900,N_28046,N_28266);
xor U28901 (N_28901,N_28176,N_28460);
nand U28902 (N_28902,N_28048,N_28053);
nand U28903 (N_28903,N_28373,N_28336);
nor U28904 (N_28904,N_28052,N_28376);
or U28905 (N_28905,N_28034,N_28177);
nor U28906 (N_28906,N_28378,N_28322);
nor U28907 (N_28907,N_28410,N_28259);
or U28908 (N_28908,N_28177,N_28159);
nand U28909 (N_28909,N_28365,N_28367);
or U28910 (N_28910,N_28006,N_28278);
nand U28911 (N_28911,N_28409,N_28403);
and U28912 (N_28912,N_28386,N_28096);
nand U28913 (N_28913,N_28467,N_28419);
xnor U28914 (N_28914,N_28222,N_28073);
nand U28915 (N_28915,N_28267,N_28292);
nor U28916 (N_28916,N_28202,N_28115);
nand U28917 (N_28917,N_28443,N_28015);
nor U28918 (N_28918,N_28350,N_28004);
and U28919 (N_28919,N_28437,N_28079);
or U28920 (N_28920,N_28425,N_28291);
and U28921 (N_28921,N_28118,N_28488);
nor U28922 (N_28922,N_28375,N_28414);
or U28923 (N_28923,N_28187,N_28057);
or U28924 (N_28924,N_28328,N_28027);
nand U28925 (N_28925,N_28252,N_28199);
nor U28926 (N_28926,N_28368,N_28494);
xnor U28927 (N_28927,N_28211,N_28446);
xor U28928 (N_28928,N_28049,N_28082);
nor U28929 (N_28929,N_28076,N_28152);
nand U28930 (N_28930,N_28121,N_28157);
nand U28931 (N_28931,N_28272,N_28097);
or U28932 (N_28932,N_28099,N_28343);
and U28933 (N_28933,N_28449,N_28126);
xor U28934 (N_28934,N_28312,N_28446);
and U28935 (N_28935,N_28337,N_28084);
xor U28936 (N_28936,N_28266,N_28262);
and U28937 (N_28937,N_28340,N_28081);
nor U28938 (N_28938,N_28128,N_28341);
and U28939 (N_28939,N_28420,N_28363);
nand U28940 (N_28940,N_28061,N_28018);
nand U28941 (N_28941,N_28406,N_28297);
nand U28942 (N_28942,N_28064,N_28048);
xnor U28943 (N_28943,N_28308,N_28480);
and U28944 (N_28944,N_28189,N_28476);
and U28945 (N_28945,N_28052,N_28250);
nand U28946 (N_28946,N_28388,N_28248);
or U28947 (N_28947,N_28494,N_28469);
and U28948 (N_28948,N_28054,N_28060);
or U28949 (N_28949,N_28283,N_28382);
and U28950 (N_28950,N_28283,N_28374);
and U28951 (N_28951,N_28154,N_28496);
or U28952 (N_28952,N_28215,N_28151);
nor U28953 (N_28953,N_28053,N_28455);
nor U28954 (N_28954,N_28033,N_28074);
xor U28955 (N_28955,N_28116,N_28100);
and U28956 (N_28956,N_28195,N_28461);
and U28957 (N_28957,N_28476,N_28072);
and U28958 (N_28958,N_28117,N_28010);
and U28959 (N_28959,N_28258,N_28104);
and U28960 (N_28960,N_28232,N_28198);
nand U28961 (N_28961,N_28088,N_28341);
and U28962 (N_28962,N_28010,N_28004);
and U28963 (N_28963,N_28028,N_28025);
or U28964 (N_28964,N_28125,N_28128);
nor U28965 (N_28965,N_28151,N_28104);
or U28966 (N_28966,N_28390,N_28338);
or U28967 (N_28967,N_28257,N_28183);
nand U28968 (N_28968,N_28215,N_28006);
and U28969 (N_28969,N_28340,N_28369);
nand U28970 (N_28970,N_28098,N_28095);
xor U28971 (N_28971,N_28205,N_28411);
xor U28972 (N_28972,N_28186,N_28399);
xor U28973 (N_28973,N_28032,N_28189);
nor U28974 (N_28974,N_28292,N_28073);
or U28975 (N_28975,N_28240,N_28024);
nand U28976 (N_28976,N_28410,N_28023);
xnor U28977 (N_28977,N_28079,N_28317);
xor U28978 (N_28978,N_28364,N_28404);
and U28979 (N_28979,N_28133,N_28124);
xnor U28980 (N_28980,N_28195,N_28174);
nor U28981 (N_28981,N_28243,N_28271);
or U28982 (N_28982,N_28373,N_28024);
nor U28983 (N_28983,N_28470,N_28442);
nor U28984 (N_28984,N_28190,N_28150);
nand U28985 (N_28985,N_28053,N_28267);
nand U28986 (N_28986,N_28336,N_28454);
nor U28987 (N_28987,N_28103,N_28457);
or U28988 (N_28988,N_28323,N_28057);
nor U28989 (N_28989,N_28030,N_28381);
xor U28990 (N_28990,N_28322,N_28483);
nand U28991 (N_28991,N_28116,N_28188);
nor U28992 (N_28992,N_28041,N_28248);
and U28993 (N_28993,N_28178,N_28167);
nor U28994 (N_28994,N_28348,N_28330);
or U28995 (N_28995,N_28328,N_28464);
nor U28996 (N_28996,N_28269,N_28301);
or U28997 (N_28997,N_28299,N_28116);
and U28998 (N_28998,N_28284,N_28076);
and U28999 (N_28999,N_28165,N_28319);
nor U29000 (N_29000,N_28695,N_28863);
nand U29001 (N_29001,N_28558,N_28841);
nand U29002 (N_29002,N_28537,N_28619);
xor U29003 (N_29003,N_28797,N_28726);
nand U29004 (N_29004,N_28748,N_28757);
or U29005 (N_29005,N_28515,N_28674);
nand U29006 (N_29006,N_28793,N_28563);
nor U29007 (N_29007,N_28738,N_28668);
or U29008 (N_29008,N_28733,N_28551);
nor U29009 (N_29009,N_28647,N_28538);
and U29010 (N_29010,N_28827,N_28544);
nor U29011 (N_29011,N_28658,N_28582);
xor U29012 (N_29012,N_28547,N_28694);
and U29013 (N_29013,N_28911,N_28833);
or U29014 (N_29014,N_28632,N_28909);
xor U29015 (N_29015,N_28772,N_28795);
or U29016 (N_29016,N_28887,N_28924);
or U29017 (N_29017,N_28705,N_28822);
xor U29018 (N_29018,N_28727,N_28825);
xor U29019 (N_29019,N_28732,N_28831);
or U29020 (N_29020,N_28778,N_28643);
xnor U29021 (N_29021,N_28902,N_28921);
xnor U29022 (N_29022,N_28768,N_28655);
and U29023 (N_29023,N_28665,N_28780);
xnor U29024 (N_29024,N_28503,N_28687);
xor U29025 (N_29025,N_28671,N_28653);
nand U29026 (N_29026,N_28720,N_28814);
nor U29027 (N_29027,N_28667,N_28696);
xor U29028 (N_29028,N_28621,N_28819);
and U29029 (N_29029,N_28791,N_28783);
xnor U29030 (N_29030,N_28517,N_28620);
and U29031 (N_29031,N_28565,N_28991);
xnor U29032 (N_29032,N_28755,N_28860);
nor U29033 (N_29033,N_28800,N_28820);
nor U29034 (N_29034,N_28818,N_28907);
nand U29035 (N_29035,N_28617,N_28927);
and U29036 (N_29036,N_28719,N_28876);
nand U29037 (N_29037,N_28976,N_28714);
nand U29038 (N_29038,N_28746,N_28850);
or U29039 (N_29039,N_28966,N_28903);
and U29040 (N_29040,N_28504,N_28897);
xnor U29041 (N_29041,N_28691,N_28592);
xnor U29042 (N_29042,N_28870,N_28759);
xnor U29043 (N_29043,N_28855,N_28629);
nand U29044 (N_29044,N_28704,N_28996);
or U29045 (N_29045,N_28873,N_28815);
xor U29046 (N_29046,N_28752,N_28523);
or U29047 (N_29047,N_28584,N_28805);
xnor U29048 (N_29048,N_28982,N_28980);
and U29049 (N_29049,N_28939,N_28593);
and U29050 (N_29050,N_28781,N_28846);
nor U29051 (N_29051,N_28634,N_28869);
and U29052 (N_29052,N_28962,N_28555);
and U29053 (N_29053,N_28590,N_28995);
nand U29054 (N_29054,N_28600,N_28811);
nand U29055 (N_29055,N_28735,N_28586);
and U29056 (N_29056,N_28889,N_28960);
or U29057 (N_29057,N_28808,N_28673);
nor U29058 (N_29058,N_28627,N_28968);
or U29059 (N_29059,N_28683,N_28766);
or U29060 (N_29060,N_28946,N_28580);
nor U29061 (N_29061,N_28804,N_28979);
nand U29062 (N_29062,N_28684,N_28882);
xor U29063 (N_29063,N_28510,N_28554);
xor U29064 (N_29064,N_28654,N_28834);
xor U29065 (N_29065,N_28843,N_28874);
or U29066 (N_29066,N_28848,N_28802);
or U29067 (N_29067,N_28926,N_28892);
xnor U29068 (N_29068,N_28830,N_28972);
xor U29069 (N_29069,N_28796,N_28676);
xnor U29070 (N_29070,N_28576,N_28697);
nand U29071 (N_29071,N_28959,N_28711);
and U29072 (N_29072,N_28739,N_28524);
and U29073 (N_29073,N_28568,N_28989);
and U29074 (N_29074,N_28597,N_28708);
xnor U29075 (N_29075,N_28591,N_28905);
xor U29076 (N_29076,N_28669,N_28853);
and U29077 (N_29077,N_28845,N_28685);
nand U29078 (N_29078,N_28541,N_28659);
or U29079 (N_29079,N_28895,N_28965);
and U29080 (N_29080,N_28707,N_28703);
and U29081 (N_29081,N_28957,N_28931);
nor U29082 (N_29082,N_28923,N_28806);
nand U29083 (N_29083,N_28657,N_28531);
xnor U29084 (N_29084,N_28609,N_28749);
nor U29085 (N_29085,N_28777,N_28832);
nor U29086 (N_29086,N_28648,N_28934);
or U29087 (N_29087,N_28813,N_28794);
nand U29088 (N_29088,N_28751,N_28737);
nand U29089 (N_29089,N_28710,N_28680);
nand U29090 (N_29090,N_28978,N_28664);
xor U29091 (N_29091,N_28545,N_28937);
and U29092 (N_29092,N_28809,N_28810);
nand U29093 (N_29093,N_28776,N_28637);
xnor U29094 (N_29094,N_28641,N_28891);
and U29095 (N_29095,N_28828,N_28666);
nor U29096 (N_29096,N_28514,N_28938);
and U29097 (N_29097,N_28508,N_28839);
and U29098 (N_29098,N_28599,N_28894);
or U29099 (N_29099,N_28678,N_28522);
xor U29100 (N_29100,N_28798,N_28816);
xnor U29101 (N_29101,N_28502,N_28856);
xor U29102 (N_29102,N_28606,N_28925);
and U29103 (N_29103,N_28635,N_28518);
nand U29104 (N_29104,N_28579,N_28928);
nor U29105 (N_29105,N_28702,N_28901);
nor U29106 (N_29106,N_28569,N_28570);
xnor U29107 (N_29107,N_28602,N_28725);
or U29108 (N_29108,N_28747,N_28782);
xnor U29109 (N_29109,N_28542,N_28628);
and U29110 (N_29110,N_28525,N_28535);
xor U29111 (N_29111,N_28754,N_28530);
xnor U29112 (N_29112,N_28756,N_28649);
and U29113 (N_29113,N_28589,N_28871);
nand U29114 (N_29114,N_28505,N_28682);
nand U29115 (N_29115,N_28999,N_28500);
nand U29116 (N_29116,N_28595,N_28829);
nor U29117 (N_29117,N_28788,N_28775);
and U29118 (N_29118,N_28573,N_28539);
nand U29119 (N_29119,N_28693,N_28598);
and U29120 (N_29120,N_28662,N_28933);
xor U29121 (N_29121,N_28618,N_28698);
or U29122 (N_29122,N_28556,N_28868);
and U29123 (N_29123,N_28935,N_28859);
xnor U29124 (N_29124,N_28823,N_28724);
xnor U29125 (N_29125,N_28936,N_28663);
nor U29126 (N_29126,N_28753,N_28890);
and U29127 (N_29127,N_28630,N_28742);
or U29128 (N_29128,N_28624,N_28983);
and U29129 (N_29129,N_28528,N_28646);
nand U29130 (N_29130,N_28867,N_28679);
and U29131 (N_29131,N_28571,N_28837);
nand U29132 (N_29132,N_28789,N_28801);
or U29133 (N_29133,N_28516,N_28501);
or U29134 (N_29134,N_28526,N_28849);
nand U29135 (N_29135,N_28826,N_28616);
and U29136 (N_29136,N_28922,N_28852);
nand U29137 (N_29137,N_28987,N_28587);
and U29138 (N_29138,N_28562,N_28779);
nand U29139 (N_29139,N_28631,N_28913);
or U29140 (N_29140,N_28672,N_28608);
and U29141 (N_29141,N_28765,N_28785);
and U29142 (N_29142,N_28633,N_28896);
or U29143 (N_29143,N_28561,N_28984);
and U29144 (N_29144,N_28533,N_28919);
nand U29145 (N_29145,N_28604,N_28821);
nor U29146 (N_29146,N_28842,N_28914);
and U29147 (N_29147,N_28851,N_28854);
xnor U29148 (N_29148,N_28880,N_28650);
xnor U29149 (N_29149,N_28988,N_28799);
xnor U29150 (N_29150,N_28844,N_28949);
nand U29151 (N_29151,N_28709,N_28866);
nand U29152 (N_29152,N_28689,N_28741);
nand U29153 (N_29153,N_28763,N_28540);
nor U29154 (N_29154,N_28520,N_28642);
and U29155 (N_29155,N_28945,N_28686);
and U29156 (N_29156,N_28560,N_28862);
nand U29157 (N_29157,N_28745,N_28534);
nand U29158 (N_29158,N_28638,N_28730);
xnor U29159 (N_29159,N_28917,N_28971);
or U29160 (N_29160,N_28900,N_28567);
nor U29161 (N_29161,N_28888,N_28622);
or U29162 (N_29162,N_28614,N_28997);
nand U29163 (N_29163,N_28993,N_28688);
nor U29164 (N_29164,N_28615,N_28603);
nand U29165 (N_29165,N_28572,N_28761);
or U29166 (N_29166,N_28527,N_28581);
nand U29167 (N_29167,N_28546,N_28881);
nor U29168 (N_29168,N_28951,N_28836);
nor U29169 (N_29169,N_28985,N_28961);
nor U29170 (N_29170,N_28990,N_28929);
and U29171 (N_29171,N_28918,N_28588);
xor U29172 (N_29172,N_28706,N_28920);
nor U29173 (N_29173,N_28625,N_28543);
xnor U29174 (N_29174,N_28875,N_28952);
or U29175 (N_29175,N_28731,N_28877);
and U29176 (N_29176,N_28743,N_28692);
nand U29177 (N_29177,N_28941,N_28986);
nand U29178 (N_29178,N_28723,N_28509);
xnor U29179 (N_29179,N_28564,N_28953);
or U29180 (N_29180,N_28915,N_28908);
nand U29181 (N_29181,N_28660,N_28549);
xor U29182 (N_29182,N_28786,N_28956);
nor U29183 (N_29183,N_28557,N_28601);
xnor U29184 (N_29184,N_28611,N_28612);
and U29185 (N_29185,N_28947,N_28879);
nand U29186 (N_29186,N_28847,N_28840);
xnor U29187 (N_29187,N_28740,N_28607);
nand U29188 (N_29188,N_28942,N_28728);
and U29189 (N_29189,N_28893,N_28940);
and U29190 (N_29190,N_28640,N_28864);
or U29191 (N_29191,N_28906,N_28974);
xnor U29192 (N_29192,N_28596,N_28661);
or U29193 (N_29193,N_28787,N_28977);
nor U29194 (N_29194,N_28729,N_28736);
nand U29195 (N_29195,N_28771,N_28675);
xnor U29196 (N_29196,N_28670,N_28838);
or U29197 (N_29197,N_28700,N_28883);
and U29198 (N_29198,N_28784,N_28944);
or U29199 (N_29199,N_28930,N_28722);
nand U29200 (N_29200,N_28932,N_28812);
or U29201 (N_29201,N_28548,N_28701);
and U29202 (N_29202,N_28718,N_28513);
nand U29203 (N_29203,N_28574,N_28636);
or U29204 (N_29204,N_28750,N_28553);
nor U29205 (N_29205,N_28511,N_28578);
xor U29206 (N_29206,N_28529,N_28566);
or U29207 (N_29207,N_28717,N_28790);
nand U29208 (N_29208,N_28758,N_28769);
nor U29209 (N_29209,N_28699,N_28858);
xor U29210 (N_29210,N_28964,N_28955);
and U29211 (N_29211,N_28992,N_28559);
and U29212 (N_29212,N_28865,N_28885);
xnor U29213 (N_29213,N_28872,N_28521);
nand U29214 (N_29214,N_28712,N_28762);
or U29215 (N_29215,N_28716,N_28734);
nor U29216 (N_29216,N_28898,N_28690);
xor U29217 (N_29217,N_28512,N_28652);
xnor U29218 (N_29218,N_28861,N_28656);
nand U29219 (N_29219,N_28916,N_28981);
or U29220 (N_29220,N_28770,N_28744);
nor U29221 (N_29221,N_28760,N_28681);
xnor U29222 (N_29222,N_28884,N_28950);
xor U29223 (N_29223,N_28575,N_28975);
and U29224 (N_29224,N_28773,N_28943);
nor U29225 (N_29225,N_28970,N_28651);
nor U29226 (N_29226,N_28803,N_28626);
nand U29227 (N_29227,N_28715,N_28764);
nand U29228 (N_29228,N_28948,N_28767);
nor U29229 (N_29229,N_28644,N_28994);
and U29230 (N_29230,N_28639,N_28963);
xnor U29231 (N_29231,N_28958,N_28645);
nor U29232 (N_29232,N_28519,N_28550);
nand U29233 (N_29233,N_28910,N_28585);
or U29234 (N_29234,N_28577,N_28899);
xnor U29235 (N_29235,N_28721,N_28912);
nand U29236 (N_29236,N_28605,N_28507);
nor U29237 (N_29237,N_28824,N_28610);
xnor U29238 (N_29238,N_28954,N_28713);
xnor U29239 (N_29239,N_28506,N_28677);
xnor U29240 (N_29240,N_28774,N_28613);
and U29241 (N_29241,N_28886,N_28835);
or U29242 (N_29242,N_28817,N_28857);
xor U29243 (N_29243,N_28967,N_28536);
nor U29244 (N_29244,N_28594,N_28552);
or U29245 (N_29245,N_28792,N_28532);
xor U29246 (N_29246,N_28583,N_28969);
xor U29247 (N_29247,N_28973,N_28998);
nand U29248 (N_29248,N_28807,N_28904);
nor U29249 (N_29249,N_28878,N_28623);
nand U29250 (N_29250,N_28692,N_28505);
xor U29251 (N_29251,N_28846,N_28857);
or U29252 (N_29252,N_28719,N_28742);
and U29253 (N_29253,N_28662,N_28860);
and U29254 (N_29254,N_28832,N_28944);
nor U29255 (N_29255,N_28522,N_28778);
and U29256 (N_29256,N_28690,N_28611);
or U29257 (N_29257,N_28648,N_28686);
nand U29258 (N_29258,N_28995,N_28854);
or U29259 (N_29259,N_28802,N_28942);
or U29260 (N_29260,N_28930,N_28556);
nand U29261 (N_29261,N_28707,N_28990);
nor U29262 (N_29262,N_28983,N_28773);
xnor U29263 (N_29263,N_28729,N_28695);
or U29264 (N_29264,N_28668,N_28520);
xor U29265 (N_29265,N_28771,N_28667);
and U29266 (N_29266,N_28642,N_28926);
nor U29267 (N_29267,N_28820,N_28585);
nand U29268 (N_29268,N_28982,N_28573);
or U29269 (N_29269,N_28904,N_28801);
and U29270 (N_29270,N_28585,N_28835);
or U29271 (N_29271,N_28547,N_28660);
and U29272 (N_29272,N_28579,N_28672);
nor U29273 (N_29273,N_28866,N_28565);
xor U29274 (N_29274,N_28710,N_28502);
or U29275 (N_29275,N_28549,N_28514);
nand U29276 (N_29276,N_28847,N_28968);
nor U29277 (N_29277,N_28753,N_28515);
or U29278 (N_29278,N_28638,N_28749);
nor U29279 (N_29279,N_28501,N_28943);
nand U29280 (N_29280,N_28860,N_28660);
xnor U29281 (N_29281,N_28878,N_28746);
nor U29282 (N_29282,N_28804,N_28812);
and U29283 (N_29283,N_28880,N_28615);
and U29284 (N_29284,N_28634,N_28916);
or U29285 (N_29285,N_28910,N_28912);
nand U29286 (N_29286,N_28963,N_28551);
nor U29287 (N_29287,N_28778,N_28589);
nand U29288 (N_29288,N_28767,N_28556);
nand U29289 (N_29289,N_28540,N_28980);
nand U29290 (N_29290,N_28606,N_28980);
or U29291 (N_29291,N_28979,N_28566);
xor U29292 (N_29292,N_28575,N_28569);
nand U29293 (N_29293,N_28736,N_28584);
xnor U29294 (N_29294,N_28530,N_28915);
or U29295 (N_29295,N_28946,N_28779);
or U29296 (N_29296,N_28844,N_28973);
nor U29297 (N_29297,N_28511,N_28694);
xor U29298 (N_29298,N_28509,N_28756);
xnor U29299 (N_29299,N_28939,N_28522);
and U29300 (N_29300,N_28579,N_28944);
xnor U29301 (N_29301,N_28509,N_28705);
or U29302 (N_29302,N_28915,N_28848);
or U29303 (N_29303,N_28631,N_28751);
nor U29304 (N_29304,N_28833,N_28569);
and U29305 (N_29305,N_28843,N_28791);
and U29306 (N_29306,N_28576,N_28885);
or U29307 (N_29307,N_28746,N_28803);
xor U29308 (N_29308,N_28567,N_28640);
or U29309 (N_29309,N_28505,N_28918);
nand U29310 (N_29310,N_28906,N_28787);
and U29311 (N_29311,N_28667,N_28567);
xor U29312 (N_29312,N_28547,N_28564);
nor U29313 (N_29313,N_28746,N_28699);
and U29314 (N_29314,N_28535,N_28973);
nor U29315 (N_29315,N_28805,N_28706);
nor U29316 (N_29316,N_28769,N_28633);
nor U29317 (N_29317,N_28890,N_28682);
or U29318 (N_29318,N_28607,N_28975);
nor U29319 (N_29319,N_28645,N_28831);
and U29320 (N_29320,N_28728,N_28535);
or U29321 (N_29321,N_28654,N_28925);
nand U29322 (N_29322,N_28859,N_28746);
nor U29323 (N_29323,N_28635,N_28785);
or U29324 (N_29324,N_28897,N_28964);
nand U29325 (N_29325,N_28610,N_28803);
or U29326 (N_29326,N_28983,N_28886);
nand U29327 (N_29327,N_28627,N_28526);
nor U29328 (N_29328,N_28707,N_28794);
and U29329 (N_29329,N_28604,N_28681);
xor U29330 (N_29330,N_28919,N_28812);
xor U29331 (N_29331,N_28987,N_28535);
xor U29332 (N_29332,N_28984,N_28790);
or U29333 (N_29333,N_28548,N_28549);
nor U29334 (N_29334,N_28695,N_28693);
or U29335 (N_29335,N_28989,N_28786);
nand U29336 (N_29336,N_28670,N_28760);
xor U29337 (N_29337,N_28639,N_28816);
nand U29338 (N_29338,N_28789,N_28579);
and U29339 (N_29339,N_28612,N_28949);
nor U29340 (N_29340,N_28555,N_28583);
xor U29341 (N_29341,N_28519,N_28713);
nor U29342 (N_29342,N_28671,N_28661);
xnor U29343 (N_29343,N_28652,N_28880);
or U29344 (N_29344,N_28595,N_28758);
nand U29345 (N_29345,N_28642,N_28570);
nor U29346 (N_29346,N_28727,N_28917);
and U29347 (N_29347,N_28565,N_28779);
xor U29348 (N_29348,N_28636,N_28759);
nor U29349 (N_29349,N_28793,N_28609);
or U29350 (N_29350,N_28717,N_28868);
xnor U29351 (N_29351,N_28744,N_28868);
and U29352 (N_29352,N_28953,N_28737);
and U29353 (N_29353,N_28681,N_28948);
xnor U29354 (N_29354,N_28630,N_28575);
nor U29355 (N_29355,N_28701,N_28681);
or U29356 (N_29356,N_28875,N_28869);
nand U29357 (N_29357,N_28655,N_28594);
nor U29358 (N_29358,N_28983,N_28941);
nor U29359 (N_29359,N_28639,N_28580);
xor U29360 (N_29360,N_28727,N_28664);
nor U29361 (N_29361,N_28808,N_28561);
nor U29362 (N_29362,N_28689,N_28701);
nor U29363 (N_29363,N_28907,N_28988);
nor U29364 (N_29364,N_28619,N_28630);
nand U29365 (N_29365,N_28734,N_28555);
xor U29366 (N_29366,N_28537,N_28843);
xnor U29367 (N_29367,N_28956,N_28748);
or U29368 (N_29368,N_28539,N_28701);
nand U29369 (N_29369,N_28902,N_28561);
nor U29370 (N_29370,N_28712,N_28928);
or U29371 (N_29371,N_28647,N_28747);
nand U29372 (N_29372,N_28942,N_28937);
or U29373 (N_29373,N_28723,N_28686);
nand U29374 (N_29374,N_28508,N_28915);
nand U29375 (N_29375,N_28997,N_28928);
and U29376 (N_29376,N_28691,N_28642);
or U29377 (N_29377,N_28807,N_28678);
nand U29378 (N_29378,N_28904,N_28616);
nor U29379 (N_29379,N_28608,N_28681);
and U29380 (N_29380,N_28755,N_28865);
and U29381 (N_29381,N_28967,N_28976);
xor U29382 (N_29382,N_28765,N_28633);
nand U29383 (N_29383,N_28657,N_28782);
nand U29384 (N_29384,N_28670,N_28942);
nand U29385 (N_29385,N_28583,N_28802);
xnor U29386 (N_29386,N_28831,N_28634);
or U29387 (N_29387,N_28775,N_28674);
or U29388 (N_29388,N_28860,N_28802);
nand U29389 (N_29389,N_28916,N_28898);
nand U29390 (N_29390,N_28977,N_28668);
or U29391 (N_29391,N_28741,N_28933);
nand U29392 (N_29392,N_28940,N_28591);
xor U29393 (N_29393,N_28685,N_28645);
nand U29394 (N_29394,N_28923,N_28770);
xnor U29395 (N_29395,N_28885,N_28689);
and U29396 (N_29396,N_28851,N_28548);
xor U29397 (N_29397,N_28669,N_28702);
or U29398 (N_29398,N_28950,N_28700);
nor U29399 (N_29399,N_28547,N_28714);
xnor U29400 (N_29400,N_28656,N_28908);
and U29401 (N_29401,N_28582,N_28858);
xor U29402 (N_29402,N_28646,N_28854);
and U29403 (N_29403,N_28907,N_28627);
xnor U29404 (N_29404,N_28580,N_28854);
or U29405 (N_29405,N_28659,N_28877);
and U29406 (N_29406,N_28801,N_28810);
nor U29407 (N_29407,N_28584,N_28620);
xor U29408 (N_29408,N_28536,N_28547);
nor U29409 (N_29409,N_28826,N_28788);
nand U29410 (N_29410,N_28662,N_28753);
or U29411 (N_29411,N_28599,N_28956);
or U29412 (N_29412,N_28571,N_28681);
nand U29413 (N_29413,N_28767,N_28543);
nand U29414 (N_29414,N_28618,N_28918);
nor U29415 (N_29415,N_28876,N_28726);
xor U29416 (N_29416,N_28952,N_28926);
or U29417 (N_29417,N_28693,N_28805);
nand U29418 (N_29418,N_28985,N_28896);
nor U29419 (N_29419,N_28643,N_28976);
nand U29420 (N_29420,N_28575,N_28964);
nand U29421 (N_29421,N_28847,N_28834);
xnor U29422 (N_29422,N_28773,N_28711);
xnor U29423 (N_29423,N_28805,N_28609);
and U29424 (N_29424,N_28841,N_28520);
or U29425 (N_29425,N_28556,N_28908);
nor U29426 (N_29426,N_28892,N_28886);
and U29427 (N_29427,N_28902,N_28560);
nor U29428 (N_29428,N_28603,N_28976);
or U29429 (N_29429,N_28712,N_28656);
or U29430 (N_29430,N_28858,N_28632);
or U29431 (N_29431,N_28882,N_28836);
nand U29432 (N_29432,N_28852,N_28634);
nor U29433 (N_29433,N_28743,N_28535);
nor U29434 (N_29434,N_28662,N_28818);
or U29435 (N_29435,N_28642,N_28534);
nand U29436 (N_29436,N_28745,N_28690);
nand U29437 (N_29437,N_28862,N_28829);
or U29438 (N_29438,N_28805,N_28730);
and U29439 (N_29439,N_28984,N_28773);
xor U29440 (N_29440,N_28654,N_28824);
xor U29441 (N_29441,N_28805,N_28648);
nor U29442 (N_29442,N_28603,N_28580);
nor U29443 (N_29443,N_28816,N_28939);
and U29444 (N_29444,N_28518,N_28848);
nor U29445 (N_29445,N_28822,N_28922);
xor U29446 (N_29446,N_28540,N_28831);
or U29447 (N_29447,N_28520,N_28760);
xnor U29448 (N_29448,N_28837,N_28758);
or U29449 (N_29449,N_28625,N_28558);
or U29450 (N_29450,N_28622,N_28529);
xor U29451 (N_29451,N_28606,N_28755);
or U29452 (N_29452,N_28630,N_28625);
or U29453 (N_29453,N_28521,N_28894);
and U29454 (N_29454,N_28949,N_28917);
xor U29455 (N_29455,N_28603,N_28781);
nand U29456 (N_29456,N_28947,N_28515);
xor U29457 (N_29457,N_28792,N_28630);
xnor U29458 (N_29458,N_28888,N_28641);
nor U29459 (N_29459,N_28548,N_28673);
or U29460 (N_29460,N_28683,N_28902);
nand U29461 (N_29461,N_28903,N_28731);
nand U29462 (N_29462,N_28806,N_28728);
or U29463 (N_29463,N_28744,N_28506);
and U29464 (N_29464,N_28574,N_28745);
nor U29465 (N_29465,N_28751,N_28630);
nand U29466 (N_29466,N_28619,N_28890);
xnor U29467 (N_29467,N_28669,N_28776);
nor U29468 (N_29468,N_28906,N_28986);
or U29469 (N_29469,N_28735,N_28528);
or U29470 (N_29470,N_28631,N_28851);
and U29471 (N_29471,N_28807,N_28782);
or U29472 (N_29472,N_28514,N_28524);
xnor U29473 (N_29473,N_28794,N_28558);
or U29474 (N_29474,N_28582,N_28649);
nor U29475 (N_29475,N_28863,N_28721);
xnor U29476 (N_29476,N_28768,N_28689);
or U29477 (N_29477,N_28694,N_28783);
nor U29478 (N_29478,N_28708,N_28901);
nand U29479 (N_29479,N_28783,N_28601);
xnor U29480 (N_29480,N_28576,N_28528);
or U29481 (N_29481,N_28645,N_28615);
xnor U29482 (N_29482,N_28746,N_28864);
nand U29483 (N_29483,N_28806,N_28880);
and U29484 (N_29484,N_28659,N_28964);
xor U29485 (N_29485,N_28918,N_28846);
xor U29486 (N_29486,N_28514,N_28643);
nand U29487 (N_29487,N_28828,N_28716);
or U29488 (N_29488,N_28770,N_28840);
nand U29489 (N_29489,N_28973,N_28905);
or U29490 (N_29490,N_28819,N_28666);
xor U29491 (N_29491,N_28513,N_28506);
and U29492 (N_29492,N_28688,N_28789);
xor U29493 (N_29493,N_28725,N_28670);
xor U29494 (N_29494,N_28923,N_28508);
and U29495 (N_29495,N_28552,N_28567);
nand U29496 (N_29496,N_28709,N_28653);
nor U29497 (N_29497,N_28649,N_28978);
and U29498 (N_29498,N_28847,N_28589);
and U29499 (N_29499,N_28625,N_28583);
or U29500 (N_29500,N_29482,N_29146);
xor U29501 (N_29501,N_29322,N_29015);
nor U29502 (N_29502,N_29467,N_29068);
xnor U29503 (N_29503,N_29290,N_29084);
nor U29504 (N_29504,N_29405,N_29284);
and U29505 (N_29505,N_29369,N_29077);
or U29506 (N_29506,N_29321,N_29025);
and U29507 (N_29507,N_29493,N_29026);
nor U29508 (N_29508,N_29488,N_29377);
and U29509 (N_29509,N_29186,N_29128);
or U29510 (N_29510,N_29013,N_29009);
and U29511 (N_29511,N_29059,N_29062);
nand U29512 (N_29512,N_29361,N_29315);
nor U29513 (N_29513,N_29384,N_29347);
xnor U29514 (N_29514,N_29253,N_29292);
and U29515 (N_29515,N_29051,N_29298);
and U29516 (N_29516,N_29181,N_29118);
xnor U29517 (N_29517,N_29403,N_29410);
or U29518 (N_29518,N_29358,N_29209);
nand U29519 (N_29519,N_29192,N_29350);
or U29520 (N_29520,N_29173,N_29004);
xor U29521 (N_29521,N_29193,N_29152);
and U29522 (N_29522,N_29497,N_29006);
and U29523 (N_29523,N_29110,N_29466);
xnor U29524 (N_29524,N_29218,N_29188);
nand U29525 (N_29525,N_29221,N_29327);
and U29526 (N_29526,N_29468,N_29450);
nor U29527 (N_29527,N_29324,N_29334);
nor U29528 (N_29528,N_29379,N_29142);
or U29529 (N_29529,N_29308,N_29370);
xnor U29530 (N_29530,N_29237,N_29392);
and U29531 (N_29531,N_29233,N_29312);
xnor U29532 (N_29532,N_29363,N_29258);
and U29533 (N_29533,N_29432,N_29032);
nand U29534 (N_29534,N_29279,N_29338);
nand U29535 (N_29535,N_29293,N_29044);
nor U29536 (N_29536,N_29280,N_29429);
nand U29537 (N_29537,N_29171,N_29356);
or U29538 (N_29538,N_29449,N_29210);
or U29539 (N_29539,N_29232,N_29225);
xnor U29540 (N_29540,N_29072,N_29011);
nor U29541 (N_29541,N_29170,N_29275);
and U29542 (N_29542,N_29409,N_29165);
xnor U29543 (N_29543,N_29163,N_29157);
xor U29544 (N_29544,N_29336,N_29424);
nor U29545 (N_29545,N_29088,N_29477);
xnor U29546 (N_29546,N_29287,N_29436);
xnor U29547 (N_29547,N_29178,N_29273);
xnor U29548 (N_29548,N_29257,N_29398);
nand U29549 (N_29549,N_29082,N_29138);
nand U29550 (N_29550,N_29156,N_29160);
xnor U29551 (N_29551,N_29254,N_29313);
nor U29552 (N_29552,N_29244,N_29199);
and U29553 (N_29553,N_29055,N_29224);
nand U29554 (N_29554,N_29302,N_29462);
xor U29555 (N_29555,N_29387,N_29208);
nor U29556 (N_29556,N_29086,N_29335);
xnor U29557 (N_29557,N_29260,N_29317);
nand U29558 (N_29558,N_29179,N_29019);
xor U29559 (N_29559,N_29437,N_29365);
or U29560 (N_29560,N_29277,N_29164);
nor U29561 (N_29561,N_29113,N_29265);
xor U29562 (N_29562,N_29139,N_29326);
and U29563 (N_29563,N_29373,N_29442);
xnor U29564 (N_29564,N_29214,N_29382);
and U29565 (N_29565,N_29499,N_29033);
xnor U29566 (N_29566,N_29433,N_29031);
and U29567 (N_29567,N_29211,N_29242);
and U29568 (N_29568,N_29487,N_29243);
or U29569 (N_29569,N_29272,N_29155);
nor U29570 (N_29570,N_29268,N_29161);
nor U29571 (N_29571,N_29415,N_29296);
or U29572 (N_29572,N_29318,N_29041);
and U29573 (N_29573,N_29021,N_29485);
nand U29574 (N_29574,N_29459,N_29134);
nor U29575 (N_29575,N_29207,N_29458);
nand U29576 (N_29576,N_29331,N_29291);
nor U29577 (N_29577,N_29039,N_29353);
and U29578 (N_29578,N_29368,N_29071);
nor U29579 (N_29579,N_29271,N_29114);
nand U29580 (N_29580,N_29107,N_29343);
nand U29581 (N_29581,N_29212,N_29469);
xnor U29582 (N_29582,N_29372,N_29337);
and U29583 (N_29583,N_29345,N_29213);
nand U29584 (N_29584,N_29422,N_29129);
and U29585 (N_29585,N_29416,N_29130);
nor U29586 (N_29586,N_29401,N_29095);
xor U29587 (N_29587,N_29256,N_29445);
nand U29588 (N_29588,N_29393,N_29465);
and U29589 (N_29589,N_29119,N_29180);
nand U29590 (N_29590,N_29219,N_29460);
xnor U29591 (N_29591,N_29305,N_29234);
nor U29592 (N_29592,N_29127,N_29255);
or U29593 (N_29593,N_29029,N_29002);
or U29594 (N_29594,N_29215,N_29137);
and U29595 (N_29595,N_29297,N_29200);
nor U29596 (N_29596,N_29120,N_29328);
nand U29597 (N_29597,N_29046,N_29206);
or U29598 (N_29598,N_29201,N_29075);
and U29599 (N_29599,N_29184,N_29235);
xnor U29600 (N_29600,N_29306,N_29177);
xnor U29601 (N_29601,N_29463,N_29252);
and U29602 (N_29602,N_29168,N_29080);
or U29603 (N_29603,N_29310,N_29438);
nand U29604 (N_29604,N_29136,N_29359);
and U29605 (N_29605,N_29319,N_29141);
xnor U29606 (N_29606,N_29223,N_29248);
xnor U29607 (N_29607,N_29230,N_29017);
or U29608 (N_29608,N_29123,N_29109);
and U29609 (N_29609,N_29079,N_29388);
nor U29610 (N_29610,N_29471,N_29117);
nor U29611 (N_29611,N_29351,N_29001);
nor U29612 (N_29612,N_29103,N_29202);
and U29613 (N_29613,N_29150,N_29456);
or U29614 (N_29614,N_29367,N_29263);
nor U29615 (N_29615,N_29143,N_29037);
and U29616 (N_29616,N_29259,N_29311);
nor U29617 (N_29617,N_29380,N_29049);
or U29618 (N_29618,N_29187,N_29111);
and U29619 (N_29619,N_29022,N_29145);
xor U29620 (N_29620,N_29149,N_29042);
nand U29621 (N_29621,N_29116,N_29070);
or U29622 (N_29622,N_29346,N_29288);
and U29623 (N_29623,N_29494,N_29480);
nor U29624 (N_29624,N_29417,N_29175);
nor U29625 (N_29625,N_29355,N_29339);
nor U29626 (N_29626,N_29381,N_29008);
nand U29627 (N_29627,N_29495,N_29091);
or U29628 (N_29628,N_29464,N_29481);
and U29629 (N_29629,N_29435,N_29183);
xnor U29630 (N_29630,N_29089,N_29144);
nor U29631 (N_29631,N_29304,N_29282);
or U29632 (N_29632,N_29301,N_29278);
xnor U29633 (N_29633,N_29198,N_29083);
nor U29634 (N_29634,N_29289,N_29060);
or U29635 (N_29635,N_29245,N_29366);
nand U29636 (N_29636,N_29020,N_29197);
nor U29637 (N_29637,N_29147,N_29362);
or U29638 (N_29638,N_29099,N_29172);
or U29639 (N_29639,N_29154,N_29411);
or U29640 (N_29640,N_29404,N_29283);
and U29641 (N_29641,N_29121,N_29076);
or U29642 (N_29642,N_29090,N_29434);
nor U29643 (N_29643,N_29489,N_29092);
xnor U29644 (N_29644,N_29455,N_29444);
or U29645 (N_29645,N_29389,N_29307);
nand U29646 (N_29646,N_29397,N_29446);
or U29647 (N_29647,N_29182,N_29457);
and U29648 (N_29648,N_29390,N_29461);
and U29649 (N_29649,N_29058,N_29131);
and U29650 (N_29650,N_29126,N_29309);
nor U29651 (N_29651,N_29344,N_29486);
and U29652 (N_29652,N_29196,N_29348);
and U29653 (N_29653,N_29045,N_29217);
nand U29654 (N_29654,N_29040,N_29300);
nand U29655 (N_29655,N_29276,N_29052);
xnor U29656 (N_29656,N_29047,N_29274);
and U29657 (N_29657,N_29240,N_29490);
nand U29658 (N_29658,N_29093,N_29108);
nand U29659 (N_29659,N_29428,N_29010);
nand U29660 (N_29660,N_29431,N_29194);
or U29661 (N_29661,N_29176,N_29453);
nor U29662 (N_29662,N_29492,N_29427);
or U29663 (N_29663,N_29249,N_29426);
or U29664 (N_29664,N_29383,N_29421);
nand U29665 (N_29665,N_29038,N_29447);
or U29666 (N_29666,N_29413,N_29185);
xnor U29667 (N_29667,N_29430,N_29281);
or U29668 (N_29668,N_29478,N_29069);
or U29669 (N_29669,N_29239,N_29078);
and U29670 (N_29670,N_29352,N_29473);
xor U29671 (N_29671,N_29028,N_29267);
nand U29672 (N_29672,N_29316,N_29386);
nor U29673 (N_29673,N_29371,N_29228);
nor U29674 (N_29674,N_29122,N_29053);
xor U29675 (N_29675,N_29231,N_29050);
and U29676 (N_29676,N_29250,N_29101);
nor U29677 (N_29677,N_29262,N_29402);
xor U29678 (N_29678,N_29330,N_29266);
xor U29679 (N_29679,N_29251,N_29323);
and U29680 (N_29680,N_29027,N_29329);
nand U29681 (N_29681,N_29391,N_29098);
nor U29682 (N_29682,N_29203,N_29375);
nand U29683 (N_29683,N_29294,N_29229);
and U29684 (N_29684,N_29132,N_29479);
nand U29685 (N_29685,N_29195,N_29357);
or U29686 (N_29686,N_29066,N_29448);
and U29687 (N_29687,N_29476,N_29412);
nand U29688 (N_29688,N_29498,N_29349);
and U29689 (N_29689,N_29135,N_29007);
or U29690 (N_29690,N_29394,N_29332);
or U29691 (N_29691,N_29005,N_29104);
xnor U29692 (N_29692,N_29423,N_29073);
and U29693 (N_29693,N_29236,N_29354);
or U29694 (N_29694,N_29096,N_29454);
xor U29695 (N_29695,N_29472,N_29102);
xnor U29696 (N_29696,N_29474,N_29148);
xnor U29697 (N_29697,N_29342,N_29261);
nand U29698 (N_29698,N_29320,N_29140);
or U29699 (N_29699,N_29169,N_29241);
nor U29700 (N_29700,N_29425,N_29067);
nor U29701 (N_29701,N_29064,N_29097);
nor U29702 (N_29702,N_29162,N_29125);
xnor U29703 (N_29703,N_29085,N_29191);
and U29704 (N_29704,N_29012,N_29166);
nor U29705 (N_29705,N_29246,N_29419);
nand U29706 (N_29706,N_29023,N_29205);
xnor U29707 (N_29707,N_29000,N_29406);
nand U29708 (N_29708,N_29376,N_29056);
and U29709 (N_29709,N_29451,N_29440);
nand U29710 (N_29710,N_29227,N_29439);
xor U29711 (N_29711,N_29112,N_29303);
or U29712 (N_29712,N_29484,N_29054);
nor U29713 (N_29713,N_29043,N_29408);
nor U29714 (N_29714,N_29189,N_29420);
and U29715 (N_29715,N_29270,N_29470);
nor U29716 (N_29716,N_29333,N_29034);
or U29717 (N_29717,N_29414,N_29061);
nor U29718 (N_29718,N_29314,N_29159);
xnor U29719 (N_29719,N_29299,N_29238);
xor U29720 (N_29720,N_29220,N_29247);
nor U29721 (N_29721,N_29396,N_29216);
nand U29722 (N_29722,N_29094,N_29443);
xnor U29723 (N_29723,N_29204,N_29360);
or U29724 (N_29724,N_29035,N_29222);
or U29725 (N_29725,N_29295,N_29036);
and U29726 (N_29726,N_29378,N_29158);
nor U29727 (N_29727,N_29087,N_29024);
nor U29728 (N_29728,N_29264,N_29407);
nand U29729 (N_29729,N_29030,N_29395);
or U29730 (N_29730,N_29190,N_29074);
or U29731 (N_29731,N_29475,N_29105);
and U29732 (N_29732,N_29048,N_29151);
xor U29733 (N_29733,N_29081,N_29491);
or U29734 (N_29734,N_29286,N_29018);
and U29735 (N_29735,N_29340,N_29167);
and U29736 (N_29736,N_29115,N_29418);
xnor U29737 (N_29737,N_29100,N_29364);
xnor U29738 (N_29738,N_29399,N_29496);
nor U29739 (N_29739,N_29374,N_29124);
or U29740 (N_29740,N_29057,N_29014);
xnor U29741 (N_29741,N_29065,N_29483);
or U29742 (N_29742,N_29441,N_29174);
and U29743 (N_29743,N_29106,N_29016);
xnor U29744 (N_29744,N_29285,N_29400);
and U29745 (N_29745,N_29063,N_29385);
and U29746 (N_29746,N_29226,N_29133);
xnor U29747 (N_29747,N_29269,N_29325);
nand U29748 (N_29748,N_29341,N_29452);
nor U29749 (N_29749,N_29003,N_29153);
and U29750 (N_29750,N_29007,N_29211);
xnor U29751 (N_29751,N_29205,N_29005);
and U29752 (N_29752,N_29318,N_29072);
xor U29753 (N_29753,N_29090,N_29125);
and U29754 (N_29754,N_29498,N_29454);
xnor U29755 (N_29755,N_29475,N_29046);
nand U29756 (N_29756,N_29120,N_29319);
nor U29757 (N_29757,N_29463,N_29372);
or U29758 (N_29758,N_29281,N_29388);
xor U29759 (N_29759,N_29299,N_29036);
nand U29760 (N_29760,N_29319,N_29406);
nand U29761 (N_29761,N_29445,N_29187);
and U29762 (N_29762,N_29423,N_29262);
nand U29763 (N_29763,N_29366,N_29195);
nand U29764 (N_29764,N_29221,N_29115);
nor U29765 (N_29765,N_29155,N_29062);
nor U29766 (N_29766,N_29163,N_29071);
nor U29767 (N_29767,N_29385,N_29305);
nand U29768 (N_29768,N_29362,N_29062);
nand U29769 (N_29769,N_29398,N_29346);
or U29770 (N_29770,N_29095,N_29241);
nor U29771 (N_29771,N_29286,N_29000);
xnor U29772 (N_29772,N_29150,N_29122);
xor U29773 (N_29773,N_29472,N_29349);
xnor U29774 (N_29774,N_29057,N_29294);
or U29775 (N_29775,N_29111,N_29127);
nand U29776 (N_29776,N_29110,N_29396);
and U29777 (N_29777,N_29226,N_29094);
xor U29778 (N_29778,N_29492,N_29225);
nand U29779 (N_29779,N_29430,N_29231);
nor U29780 (N_29780,N_29046,N_29470);
nor U29781 (N_29781,N_29446,N_29366);
or U29782 (N_29782,N_29063,N_29068);
xnor U29783 (N_29783,N_29497,N_29386);
nand U29784 (N_29784,N_29490,N_29382);
nand U29785 (N_29785,N_29202,N_29017);
nand U29786 (N_29786,N_29318,N_29422);
and U29787 (N_29787,N_29153,N_29364);
or U29788 (N_29788,N_29381,N_29462);
xnor U29789 (N_29789,N_29199,N_29253);
or U29790 (N_29790,N_29239,N_29450);
nand U29791 (N_29791,N_29403,N_29374);
xor U29792 (N_29792,N_29070,N_29199);
and U29793 (N_29793,N_29484,N_29041);
nand U29794 (N_29794,N_29482,N_29236);
xor U29795 (N_29795,N_29381,N_29456);
nor U29796 (N_29796,N_29491,N_29217);
or U29797 (N_29797,N_29019,N_29209);
xor U29798 (N_29798,N_29361,N_29235);
or U29799 (N_29799,N_29157,N_29389);
and U29800 (N_29800,N_29447,N_29422);
xnor U29801 (N_29801,N_29195,N_29197);
and U29802 (N_29802,N_29094,N_29367);
nand U29803 (N_29803,N_29346,N_29091);
and U29804 (N_29804,N_29123,N_29133);
nand U29805 (N_29805,N_29188,N_29009);
or U29806 (N_29806,N_29392,N_29023);
and U29807 (N_29807,N_29223,N_29446);
xor U29808 (N_29808,N_29172,N_29459);
or U29809 (N_29809,N_29061,N_29322);
and U29810 (N_29810,N_29250,N_29383);
and U29811 (N_29811,N_29175,N_29420);
and U29812 (N_29812,N_29269,N_29204);
and U29813 (N_29813,N_29285,N_29247);
nand U29814 (N_29814,N_29227,N_29194);
and U29815 (N_29815,N_29225,N_29035);
nand U29816 (N_29816,N_29284,N_29450);
xor U29817 (N_29817,N_29006,N_29030);
or U29818 (N_29818,N_29228,N_29251);
xor U29819 (N_29819,N_29136,N_29118);
and U29820 (N_29820,N_29332,N_29248);
nor U29821 (N_29821,N_29356,N_29291);
nor U29822 (N_29822,N_29186,N_29182);
nand U29823 (N_29823,N_29290,N_29450);
nand U29824 (N_29824,N_29108,N_29137);
and U29825 (N_29825,N_29107,N_29493);
or U29826 (N_29826,N_29111,N_29417);
nand U29827 (N_29827,N_29019,N_29262);
nor U29828 (N_29828,N_29460,N_29062);
nand U29829 (N_29829,N_29279,N_29203);
or U29830 (N_29830,N_29242,N_29328);
or U29831 (N_29831,N_29442,N_29262);
xor U29832 (N_29832,N_29261,N_29371);
or U29833 (N_29833,N_29453,N_29130);
or U29834 (N_29834,N_29103,N_29307);
nor U29835 (N_29835,N_29398,N_29399);
xnor U29836 (N_29836,N_29084,N_29169);
or U29837 (N_29837,N_29135,N_29183);
nand U29838 (N_29838,N_29387,N_29197);
xnor U29839 (N_29839,N_29340,N_29274);
or U29840 (N_29840,N_29030,N_29446);
nand U29841 (N_29841,N_29113,N_29187);
xnor U29842 (N_29842,N_29287,N_29112);
nand U29843 (N_29843,N_29267,N_29202);
or U29844 (N_29844,N_29267,N_29399);
nor U29845 (N_29845,N_29072,N_29497);
or U29846 (N_29846,N_29466,N_29486);
or U29847 (N_29847,N_29496,N_29093);
and U29848 (N_29848,N_29140,N_29260);
xnor U29849 (N_29849,N_29447,N_29430);
xor U29850 (N_29850,N_29159,N_29440);
nand U29851 (N_29851,N_29259,N_29122);
nor U29852 (N_29852,N_29352,N_29226);
xnor U29853 (N_29853,N_29166,N_29113);
or U29854 (N_29854,N_29402,N_29155);
and U29855 (N_29855,N_29353,N_29471);
nor U29856 (N_29856,N_29204,N_29304);
nand U29857 (N_29857,N_29319,N_29163);
nand U29858 (N_29858,N_29075,N_29032);
and U29859 (N_29859,N_29120,N_29022);
and U29860 (N_29860,N_29355,N_29452);
xor U29861 (N_29861,N_29134,N_29360);
xnor U29862 (N_29862,N_29019,N_29196);
nor U29863 (N_29863,N_29208,N_29357);
nand U29864 (N_29864,N_29490,N_29117);
and U29865 (N_29865,N_29161,N_29108);
and U29866 (N_29866,N_29118,N_29187);
nor U29867 (N_29867,N_29104,N_29398);
nor U29868 (N_29868,N_29402,N_29021);
or U29869 (N_29869,N_29169,N_29467);
or U29870 (N_29870,N_29074,N_29427);
and U29871 (N_29871,N_29354,N_29050);
and U29872 (N_29872,N_29232,N_29171);
or U29873 (N_29873,N_29448,N_29077);
and U29874 (N_29874,N_29428,N_29100);
nand U29875 (N_29875,N_29009,N_29116);
and U29876 (N_29876,N_29491,N_29227);
xor U29877 (N_29877,N_29034,N_29390);
nand U29878 (N_29878,N_29405,N_29469);
nor U29879 (N_29879,N_29205,N_29245);
xnor U29880 (N_29880,N_29104,N_29108);
or U29881 (N_29881,N_29318,N_29296);
or U29882 (N_29882,N_29469,N_29210);
xnor U29883 (N_29883,N_29395,N_29213);
or U29884 (N_29884,N_29126,N_29122);
xor U29885 (N_29885,N_29357,N_29191);
nand U29886 (N_29886,N_29008,N_29180);
nor U29887 (N_29887,N_29481,N_29432);
xnor U29888 (N_29888,N_29120,N_29151);
nor U29889 (N_29889,N_29245,N_29488);
or U29890 (N_29890,N_29306,N_29153);
nor U29891 (N_29891,N_29060,N_29496);
or U29892 (N_29892,N_29309,N_29186);
nand U29893 (N_29893,N_29476,N_29173);
nor U29894 (N_29894,N_29078,N_29388);
nor U29895 (N_29895,N_29158,N_29389);
or U29896 (N_29896,N_29115,N_29483);
or U29897 (N_29897,N_29440,N_29108);
xor U29898 (N_29898,N_29243,N_29010);
nor U29899 (N_29899,N_29462,N_29085);
nor U29900 (N_29900,N_29395,N_29439);
or U29901 (N_29901,N_29409,N_29197);
nor U29902 (N_29902,N_29246,N_29330);
or U29903 (N_29903,N_29208,N_29398);
nor U29904 (N_29904,N_29493,N_29270);
xnor U29905 (N_29905,N_29412,N_29202);
and U29906 (N_29906,N_29252,N_29035);
nand U29907 (N_29907,N_29321,N_29333);
xor U29908 (N_29908,N_29123,N_29287);
nand U29909 (N_29909,N_29060,N_29386);
xor U29910 (N_29910,N_29192,N_29461);
or U29911 (N_29911,N_29356,N_29285);
or U29912 (N_29912,N_29431,N_29064);
and U29913 (N_29913,N_29156,N_29031);
xor U29914 (N_29914,N_29223,N_29152);
or U29915 (N_29915,N_29223,N_29373);
nor U29916 (N_29916,N_29191,N_29383);
and U29917 (N_29917,N_29115,N_29413);
or U29918 (N_29918,N_29489,N_29346);
nor U29919 (N_29919,N_29254,N_29100);
nor U29920 (N_29920,N_29426,N_29481);
nor U29921 (N_29921,N_29243,N_29006);
nor U29922 (N_29922,N_29028,N_29214);
nor U29923 (N_29923,N_29432,N_29219);
or U29924 (N_29924,N_29371,N_29237);
xnor U29925 (N_29925,N_29010,N_29022);
nor U29926 (N_29926,N_29498,N_29377);
and U29927 (N_29927,N_29445,N_29421);
and U29928 (N_29928,N_29347,N_29307);
xor U29929 (N_29929,N_29145,N_29175);
or U29930 (N_29930,N_29132,N_29454);
and U29931 (N_29931,N_29373,N_29119);
nor U29932 (N_29932,N_29445,N_29309);
and U29933 (N_29933,N_29224,N_29296);
nand U29934 (N_29934,N_29108,N_29024);
or U29935 (N_29935,N_29036,N_29317);
nor U29936 (N_29936,N_29119,N_29338);
and U29937 (N_29937,N_29351,N_29256);
and U29938 (N_29938,N_29365,N_29230);
or U29939 (N_29939,N_29015,N_29033);
nand U29940 (N_29940,N_29072,N_29177);
xor U29941 (N_29941,N_29374,N_29425);
or U29942 (N_29942,N_29433,N_29136);
xor U29943 (N_29943,N_29151,N_29042);
nand U29944 (N_29944,N_29349,N_29454);
nor U29945 (N_29945,N_29464,N_29088);
nor U29946 (N_29946,N_29306,N_29012);
or U29947 (N_29947,N_29031,N_29480);
nor U29948 (N_29948,N_29070,N_29417);
xnor U29949 (N_29949,N_29165,N_29280);
and U29950 (N_29950,N_29133,N_29326);
or U29951 (N_29951,N_29213,N_29337);
or U29952 (N_29952,N_29280,N_29425);
xnor U29953 (N_29953,N_29056,N_29092);
xnor U29954 (N_29954,N_29106,N_29440);
nand U29955 (N_29955,N_29449,N_29091);
nor U29956 (N_29956,N_29203,N_29166);
xor U29957 (N_29957,N_29452,N_29317);
xnor U29958 (N_29958,N_29184,N_29238);
or U29959 (N_29959,N_29475,N_29356);
and U29960 (N_29960,N_29079,N_29255);
or U29961 (N_29961,N_29377,N_29406);
or U29962 (N_29962,N_29029,N_29474);
and U29963 (N_29963,N_29399,N_29387);
or U29964 (N_29964,N_29259,N_29287);
nand U29965 (N_29965,N_29095,N_29199);
nand U29966 (N_29966,N_29149,N_29023);
nand U29967 (N_29967,N_29283,N_29338);
or U29968 (N_29968,N_29045,N_29306);
xor U29969 (N_29969,N_29100,N_29182);
and U29970 (N_29970,N_29175,N_29468);
nor U29971 (N_29971,N_29488,N_29319);
and U29972 (N_29972,N_29063,N_29333);
and U29973 (N_29973,N_29318,N_29020);
and U29974 (N_29974,N_29084,N_29472);
xnor U29975 (N_29975,N_29131,N_29038);
xor U29976 (N_29976,N_29245,N_29362);
xor U29977 (N_29977,N_29021,N_29167);
xor U29978 (N_29978,N_29179,N_29276);
xor U29979 (N_29979,N_29413,N_29016);
or U29980 (N_29980,N_29389,N_29443);
and U29981 (N_29981,N_29011,N_29270);
xnor U29982 (N_29982,N_29384,N_29305);
xor U29983 (N_29983,N_29189,N_29405);
nor U29984 (N_29984,N_29029,N_29207);
nand U29985 (N_29985,N_29250,N_29400);
or U29986 (N_29986,N_29121,N_29496);
nor U29987 (N_29987,N_29004,N_29065);
or U29988 (N_29988,N_29142,N_29405);
xnor U29989 (N_29989,N_29102,N_29143);
nand U29990 (N_29990,N_29077,N_29243);
nand U29991 (N_29991,N_29140,N_29496);
and U29992 (N_29992,N_29025,N_29303);
and U29993 (N_29993,N_29231,N_29258);
xor U29994 (N_29994,N_29329,N_29186);
nand U29995 (N_29995,N_29144,N_29153);
nor U29996 (N_29996,N_29079,N_29376);
xnor U29997 (N_29997,N_29250,N_29329);
nand U29998 (N_29998,N_29431,N_29069);
nor U29999 (N_29999,N_29112,N_29387);
and UO_0 (O_0,N_29782,N_29924);
or UO_1 (O_1,N_29872,N_29516);
or UO_2 (O_2,N_29860,N_29763);
nor UO_3 (O_3,N_29759,N_29644);
and UO_4 (O_4,N_29737,N_29680);
and UO_5 (O_5,N_29977,N_29593);
and UO_6 (O_6,N_29895,N_29795);
nand UO_7 (O_7,N_29932,N_29538);
nand UO_8 (O_8,N_29767,N_29891);
xnor UO_9 (O_9,N_29546,N_29619);
nor UO_10 (O_10,N_29682,N_29614);
and UO_11 (O_11,N_29637,N_29889);
xnor UO_12 (O_12,N_29804,N_29996);
xor UO_13 (O_13,N_29707,N_29848);
nor UO_14 (O_14,N_29999,N_29567);
or UO_15 (O_15,N_29590,N_29665);
xnor UO_16 (O_16,N_29969,N_29908);
nand UO_17 (O_17,N_29610,N_29942);
nand UO_18 (O_18,N_29608,N_29958);
or UO_19 (O_19,N_29808,N_29881);
nor UO_20 (O_20,N_29612,N_29527);
xor UO_21 (O_21,N_29744,N_29851);
or UO_22 (O_22,N_29943,N_29971);
nor UO_23 (O_23,N_29626,N_29713);
nor UO_24 (O_24,N_29620,N_29653);
nand UO_25 (O_25,N_29831,N_29978);
or UO_26 (O_26,N_29790,N_29915);
or UO_27 (O_27,N_29761,N_29993);
and UO_28 (O_28,N_29687,N_29771);
xnor UO_29 (O_29,N_29894,N_29950);
xnor UO_30 (O_30,N_29903,N_29788);
nand UO_31 (O_31,N_29579,N_29515);
nand UO_32 (O_32,N_29743,N_29921);
nor UO_33 (O_33,N_29602,N_29990);
or UO_34 (O_34,N_29973,N_29754);
or UO_35 (O_35,N_29630,N_29651);
nor UO_36 (O_36,N_29668,N_29575);
nand UO_37 (O_37,N_29883,N_29581);
nand UO_38 (O_38,N_29642,N_29890);
or UO_39 (O_39,N_29641,N_29525);
and UO_40 (O_40,N_29632,N_29721);
or UO_41 (O_41,N_29736,N_29667);
or UO_42 (O_42,N_29805,N_29899);
and UO_43 (O_43,N_29888,N_29607);
and UO_44 (O_44,N_29512,N_29898);
or UO_45 (O_45,N_29726,N_29912);
nor UO_46 (O_46,N_29727,N_29697);
nor UO_47 (O_47,N_29949,N_29542);
nor UO_48 (O_48,N_29529,N_29838);
nand UO_49 (O_49,N_29989,N_29572);
nand UO_50 (O_50,N_29778,N_29933);
and UO_51 (O_51,N_29852,N_29826);
xor UO_52 (O_52,N_29663,N_29959);
or UO_53 (O_53,N_29827,N_29675);
and UO_54 (O_54,N_29998,N_29897);
and UO_55 (O_55,N_29875,N_29649);
xnor UO_56 (O_56,N_29864,N_29750);
nand UO_57 (O_57,N_29829,N_29671);
nand UO_58 (O_58,N_29765,N_29693);
and UO_59 (O_59,N_29659,N_29878);
and UO_60 (O_60,N_29625,N_29601);
nor UO_61 (O_61,N_29640,N_29664);
and UO_62 (O_62,N_29940,N_29725);
nor UO_63 (O_63,N_29749,N_29561);
xor UO_64 (O_64,N_29807,N_29738);
and UO_65 (O_65,N_29967,N_29603);
xor UO_66 (O_66,N_29592,N_29714);
xor UO_67 (O_67,N_29518,N_29972);
or UO_68 (O_68,N_29643,N_29780);
or UO_69 (O_69,N_29700,N_29769);
xnor UO_70 (O_70,N_29683,N_29505);
nor UO_71 (O_71,N_29623,N_29841);
or UO_72 (O_72,N_29957,N_29877);
xnor UO_73 (O_73,N_29655,N_29944);
nand UO_74 (O_74,N_29900,N_29624);
and UO_75 (O_75,N_29728,N_29753);
xor UO_76 (O_76,N_29509,N_29676);
or UO_77 (O_77,N_29656,N_29824);
nor UO_78 (O_78,N_29695,N_29861);
xnor UO_79 (O_79,N_29658,N_29712);
nor UO_80 (O_80,N_29734,N_29660);
or UO_81 (O_81,N_29554,N_29513);
nor UO_82 (O_82,N_29783,N_29735);
or UO_83 (O_83,N_29616,N_29688);
and UO_84 (O_84,N_29965,N_29893);
or UO_85 (O_85,N_29530,N_29885);
or UO_86 (O_86,N_29652,N_29573);
and UO_87 (O_87,N_29715,N_29500);
and UO_88 (O_88,N_29563,N_29634);
nor UO_89 (O_89,N_29822,N_29920);
nand UO_90 (O_90,N_29757,N_29692);
and UO_91 (O_91,N_29504,N_29691);
xnor UO_92 (O_92,N_29834,N_29636);
and UO_93 (O_93,N_29723,N_29540);
or UO_94 (O_94,N_29997,N_29722);
and UO_95 (O_95,N_29785,N_29923);
nor UO_96 (O_96,N_29938,N_29992);
xor UO_97 (O_97,N_29628,N_29947);
and UO_98 (O_98,N_29926,N_29764);
nor UO_99 (O_99,N_29797,N_29814);
xnor UO_100 (O_100,N_29584,N_29528);
xor UO_101 (O_101,N_29589,N_29832);
or UO_102 (O_102,N_29879,N_29657);
or UO_103 (O_103,N_29793,N_29510);
or UO_104 (O_104,N_29919,N_29756);
nor UO_105 (O_105,N_29532,N_29987);
nand UO_106 (O_106,N_29597,N_29719);
and UO_107 (O_107,N_29670,N_29865);
nand UO_108 (O_108,N_29874,N_29842);
nand UO_109 (O_109,N_29577,N_29799);
nand UO_110 (O_110,N_29574,N_29545);
xor UO_111 (O_111,N_29536,N_29913);
or UO_112 (O_112,N_29507,N_29704);
nand UO_113 (O_113,N_29629,N_29552);
and UO_114 (O_114,N_29605,N_29905);
or UO_115 (O_115,N_29806,N_29937);
nand UO_116 (O_116,N_29731,N_29880);
and UO_117 (O_117,N_29741,N_29635);
nand UO_118 (O_118,N_29836,N_29689);
xor UO_119 (O_119,N_29594,N_29720);
xor UO_120 (O_120,N_29907,N_29514);
and UO_121 (O_121,N_29698,N_29857);
nand UO_122 (O_122,N_29850,N_29846);
nor UO_123 (O_123,N_29639,N_29646);
and UO_124 (O_124,N_29758,N_29553);
nand UO_125 (O_125,N_29854,N_29576);
nor UO_126 (O_126,N_29954,N_29777);
and UO_127 (O_127,N_29935,N_29939);
or UO_128 (O_128,N_29746,N_29648);
xnor UO_129 (O_129,N_29729,N_29696);
and UO_130 (O_130,N_29882,N_29855);
xnor UO_131 (O_131,N_29873,N_29781);
nor UO_132 (O_132,N_29568,N_29533);
nor UO_133 (O_133,N_29618,N_29849);
or UO_134 (O_134,N_29730,N_29586);
xor UO_135 (O_135,N_29591,N_29833);
and UO_136 (O_136,N_29869,N_29966);
or UO_137 (O_137,N_29588,N_29747);
nor UO_138 (O_138,N_29535,N_29779);
nor UO_139 (O_139,N_29724,N_29521);
nand UO_140 (O_140,N_29910,N_29548);
or UO_141 (O_141,N_29526,N_29981);
and UO_142 (O_142,N_29776,N_29543);
nand UO_143 (O_143,N_29517,N_29520);
nor UO_144 (O_144,N_29669,N_29925);
nor UO_145 (O_145,N_29703,N_29564);
and UO_146 (O_146,N_29549,N_29887);
xnor UO_147 (O_147,N_29970,N_29839);
and UO_148 (O_148,N_29760,N_29914);
nor UO_149 (O_149,N_29803,N_29968);
nand UO_150 (O_150,N_29708,N_29537);
or UO_151 (O_151,N_29876,N_29884);
and UO_152 (O_152,N_29596,N_29931);
nand UO_153 (O_153,N_29963,N_29558);
nor UO_154 (O_154,N_29627,N_29582);
nor UO_155 (O_155,N_29856,N_29733);
xnor UO_156 (O_156,N_29508,N_29844);
or UO_157 (O_157,N_29952,N_29524);
and UO_158 (O_158,N_29948,N_29916);
nor UO_159 (O_159,N_29816,N_29867);
nor UO_160 (O_160,N_29936,N_29511);
xor UO_161 (O_161,N_29631,N_29709);
xor UO_162 (O_162,N_29995,N_29953);
or UO_163 (O_163,N_29820,N_29661);
and UO_164 (O_164,N_29904,N_29984);
nand UO_165 (O_165,N_29985,N_29858);
nor UO_166 (O_166,N_29927,N_29974);
or UO_167 (O_167,N_29701,N_29633);
nor UO_168 (O_168,N_29565,N_29650);
or UO_169 (O_169,N_29975,N_29599);
xor UO_170 (O_170,N_29569,N_29613);
or UO_171 (O_171,N_29560,N_29845);
or UO_172 (O_172,N_29906,N_29929);
or UO_173 (O_173,N_29994,N_29541);
nand UO_174 (O_174,N_29557,N_29980);
nand UO_175 (O_175,N_29802,N_29621);
nor UO_176 (O_176,N_29611,N_29587);
xnor UO_177 (O_177,N_29911,N_29666);
nand UO_178 (O_178,N_29654,N_29684);
nand UO_179 (O_179,N_29506,N_29732);
and UO_180 (O_180,N_29559,N_29812);
or UO_181 (O_181,N_29868,N_29556);
nor UO_182 (O_182,N_29870,N_29706);
and UO_183 (O_183,N_29951,N_29815);
nor UO_184 (O_184,N_29813,N_29922);
and UO_185 (O_185,N_29681,N_29823);
and UO_186 (O_186,N_29991,N_29555);
or UO_187 (O_187,N_29673,N_29585);
or UO_188 (O_188,N_29794,N_29918);
or UO_189 (O_189,N_29960,N_29501);
nor UO_190 (O_190,N_29818,N_29934);
and UO_191 (O_191,N_29786,N_29672);
or UO_192 (O_192,N_29578,N_29847);
or UO_193 (O_193,N_29745,N_29766);
nand UO_194 (O_194,N_29705,N_29571);
nand UO_195 (O_195,N_29690,N_29828);
nand UO_196 (O_196,N_29717,N_29787);
and UO_197 (O_197,N_29662,N_29566);
nand UO_198 (O_198,N_29762,N_29686);
or UO_199 (O_199,N_29711,N_29604);
xor UO_200 (O_200,N_29755,N_29896);
or UO_201 (O_201,N_29821,N_29819);
nand UO_202 (O_202,N_29674,N_29742);
nor UO_203 (O_203,N_29609,N_29946);
and UO_204 (O_204,N_29941,N_29817);
nand UO_205 (O_205,N_29519,N_29901);
xor UO_206 (O_206,N_29685,N_29774);
or UO_207 (O_207,N_29983,N_29752);
or UO_208 (O_208,N_29716,N_29617);
and UO_209 (O_209,N_29835,N_29956);
xor UO_210 (O_210,N_29909,N_29902);
or UO_211 (O_211,N_29792,N_29570);
nor UO_212 (O_212,N_29964,N_29772);
nand UO_213 (O_213,N_29615,N_29677);
xnor UO_214 (O_214,N_29796,N_29544);
and UO_215 (O_215,N_29988,N_29955);
or UO_216 (O_216,N_29928,N_29801);
or UO_217 (O_217,N_29502,N_29830);
nand UO_218 (O_218,N_29534,N_29595);
or UO_219 (O_219,N_29892,N_29768);
nor UO_220 (O_220,N_29551,N_29751);
xnor UO_221 (O_221,N_29917,N_29694);
and UO_222 (O_222,N_29740,N_29961);
or UO_223 (O_223,N_29982,N_29638);
xnor UO_224 (O_224,N_29945,N_29791);
and UO_225 (O_225,N_29718,N_29583);
and UO_226 (O_226,N_29825,N_29930);
xnor UO_227 (O_227,N_29871,N_29531);
nand UO_228 (O_228,N_29853,N_29739);
nand UO_229 (O_229,N_29789,N_29863);
and UO_230 (O_230,N_29547,N_29798);
and UO_231 (O_231,N_29770,N_29523);
nor UO_232 (O_232,N_29840,N_29710);
nand UO_233 (O_233,N_29645,N_29606);
nor UO_234 (O_234,N_29837,N_29522);
xor UO_235 (O_235,N_29800,N_29809);
nor UO_236 (O_236,N_29647,N_29976);
nand UO_237 (O_237,N_29866,N_29562);
xnor UO_238 (O_238,N_29679,N_29962);
nor UO_239 (O_239,N_29775,N_29859);
or UO_240 (O_240,N_29678,N_29886);
nor UO_241 (O_241,N_29862,N_29843);
xor UO_242 (O_242,N_29539,N_29702);
nand UO_243 (O_243,N_29598,N_29550);
nor UO_244 (O_244,N_29773,N_29748);
and UO_245 (O_245,N_29580,N_29622);
xor UO_246 (O_246,N_29784,N_29810);
xor UO_247 (O_247,N_29979,N_29600);
xnor UO_248 (O_248,N_29503,N_29986);
xnor UO_249 (O_249,N_29699,N_29811);
or UO_250 (O_250,N_29639,N_29596);
or UO_251 (O_251,N_29588,N_29710);
nand UO_252 (O_252,N_29846,N_29670);
nor UO_253 (O_253,N_29618,N_29609);
or UO_254 (O_254,N_29585,N_29732);
and UO_255 (O_255,N_29790,N_29990);
nand UO_256 (O_256,N_29670,N_29671);
nand UO_257 (O_257,N_29705,N_29921);
nand UO_258 (O_258,N_29546,N_29953);
and UO_259 (O_259,N_29780,N_29817);
and UO_260 (O_260,N_29722,N_29729);
nor UO_261 (O_261,N_29508,N_29783);
or UO_262 (O_262,N_29952,N_29965);
or UO_263 (O_263,N_29593,N_29841);
or UO_264 (O_264,N_29970,N_29718);
xnor UO_265 (O_265,N_29826,N_29997);
and UO_266 (O_266,N_29540,N_29944);
nor UO_267 (O_267,N_29612,N_29956);
and UO_268 (O_268,N_29940,N_29981);
nand UO_269 (O_269,N_29579,N_29791);
or UO_270 (O_270,N_29745,N_29849);
xor UO_271 (O_271,N_29546,N_29694);
xor UO_272 (O_272,N_29506,N_29994);
and UO_273 (O_273,N_29809,N_29718);
nor UO_274 (O_274,N_29735,N_29615);
xnor UO_275 (O_275,N_29504,N_29761);
and UO_276 (O_276,N_29652,N_29566);
and UO_277 (O_277,N_29911,N_29898);
nand UO_278 (O_278,N_29678,N_29947);
nor UO_279 (O_279,N_29773,N_29739);
nand UO_280 (O_280,N_29956,N_29831);
or UO_281 (O_281,N_29941,N_29916);
xor UO_282 (O_282,N_29597,N_29948);
nor UO_283 (O_283,N_29520,N_29788);
nor UO_284 (O_284,N_29880,N_29570);
or UO_285 (O_285,N_29983,N_29573);
or UO_286 (O_286,N_29648,N_29759);
nand UO_287 (O_287,N_29506,N_29632);
nor UO_288 (O_288,N_29899,N_29719);
nor UO_289 (O_289,N_29504,N_29933);
nand UO_290 (O_290,N_29502,N_29737);
nand UO_291 (O_291,N_29954,N_29941);
nor UO_292 (O_292,N_29992,N_29819);
xor UO_293 (O_293,N_29911,N_29688);
and UO_294 (O_294,N_29723,N_29677);
nand UO_295 (O_295,N_29839,N_29554);
and UO_296 (O_296,N_29877,N_29875);
nor UO_297 (O_297,N_29539,N_29704);
and UO_298 (O_298,N_29901,N_29671);
or UO_299 (O_299,N_29650,N_29635);
xnor UO_300 (O_300,N_29579,N_29987);
and UO_301 (O_301,N_29702,N_29707);
xnor UO_302 (O_302,N_29669,N_29595);
and UO_303 (O_303,N_29994,N_29606);
and UO_304 (O_304,N_29772,N_29803);
and UO_305 (O_305,N_29987,N_29863);
xor UO_306 (O_306,N_29667,N_29684);
or UO_307 (O_307,N_29973,N_29850);
nand UO_308 (O_308,N_29632,N_29831);
nand UO_309 (O_309,N_29935,N_29807);
and UO_310 (O_310,N_29710,N_29617);
or UO_311 (O_311,N_29759,N_29584);
and UO_312 (O_312,N_29655,N_29862);
xor UO_313 (O_313,N_29619,N_29832);
xor UO_314 (O_314,N_29577,N_29965);
and UO_315 (O_315,N_29943,N_29927);
nand UO_316 (O_316,N_29658,N_29789);
xnor UO_317 (O_317,N_29945,N_29853);
nor UO_318 (O_318,N_29771,N_29659);
nor UO_319 (O_319,N_29537,N_29572);
and UO_320 (O_320,N_29737,N_29725);
xnor UO_321 (O_321,N_29883,N_29874);
xnor UO_322 (O_322,N_29884,N_29595);
nand UO_323 (O_323,N_29632,N_29526);
xor UO_324 (O_324,N_29804,N_29827);
and UO_325 (O_325,N_29651,N_29520);
nor UO_326 (O_326,N_29968,N_29582);
and UO_327 (O_327,N_29870,N_29876);
nor UO_328 (O_328,N_29897,N_29961);
or UO_329 (O_329,N_29888,N_29843);
nor UO_330 (O_330,N_29672,N_29659);
nor UO_331 (O_331,N_29804,N_29684);
xnor UO_332 (O_332,N_29712,N_29964);
and UO_333 (O_333,N_29818,N_29790);
nand UO_334 (O_334,N_29626,N_29788);
xnor UO_335 (O_335,N_29560,N_29693);
nor UO_336 (O_336,N_29711,N_29961);
xor UO_337 (O_337,N_29869,N_29815);
and UO_338 (O_338,N_29621,N_29727);
nand UO_339 (O_339,N_29997,N_29738);
nor UO_340 (O_340,N_29811,N_29710);
and UO_341 (O_341,N_29637,N_29827);
and UO_342 (O_342,N_29879,N_29596);
nor UO_343 (O_343,N_29682,N_29617);
xnor UO_344 (O_344,N_29716,N_29664);
or UO_345 (O_345,N_29848,N_29624);
nor UO_346 (O_346,N_29916,N_29615);
nor UO_347 (O_347,N_29997,N_29650);
xor UO_348 (O_348,N_29996,N_29815);
or UO_349 (O_349,N_29541,N_29957);
and UO_350 (O_350,N_29951,N_29918);
and UO_351 (O_351,N_29512,N_29907);
xor UO_352 (O_352,N_29734,N_29923);
or UO_353 (O_353,N_29986,N_29941);
xor UO_354 (O_354,N_29682,N_29924);
nand UO_355 (O_355,N_29851,N_29575);
and UO_356 (O_356,N_29693,N_29999);
nand UO_357 (O_357,N_29583,N_29592);
and UO_358 (O_358,N_29564,N_29585);
or UO_359 (O_359,N_29766,N_29878);
nand UO_360 (O_360,N_29589,N_29910);
or UO_361 (O_361,N_29761,N_29825);
or UO_362 (O_362,N_29581,N_29809);
xor UO_363 (O_363,N_29658,N_29555);
xor UO_364 (O_364,N_29541,N_29999);
xor UO_365 (O_365,N_29695,N_29810);
xor UO_366 (O_366,N_29892,N_29932);
nor UO_367 (O_367,N_29784,N_29971);
xor UO_368 (O_368,N_29795,N_29861);
or UO_369 (O_369,N_29559,N_29918);
nand UO_370 (O_370,N_29649,N_29538);
xor UO_371 (O_371,N_29746,N_29969);
nor UO_372 (O_372,N_29986,N_29548);
nand UO_373 (O_373,N_29662,N_29750);
nand UO_374 (O_374,N_29974,N_29924);
nor UO_375 (O_375,N_29776,N_29606);
xor UO_376 (O_376,N_29743,N_29673);
or UO_377 (O_377,N_29821,N_29953);
nor UO_378 (O_378,N_29846,N_29613);
nor UO_379 (O_379,N_29914,N_29657);
xor UO_380 (O_380,N_29530,N_29561);
nor UO_381 (O_381,N_29758,N_29607);
nand UO_382 (O_382,N_29683,N_29837);
xnor UO_383 (O_383,N_29523,N_29786);
or UO_384 (O_384,N_29962,N_29878);
xor UO_385 (O_385,N_29783,N_29796);
xor UO_386 (O_386,N_29615,N_29659);
nand UO_387 (O_387,N_29584,N_29601);
and UO_388 (O_388,N_29545,N_29858);
and UO_389 (O_389,N_29877,N_29654);
xnor UO_390 (O_390,N_29973,N_29548);
nor UO_391 (O_391,N_29674,N_29644);
nor UO_392 (O_392,N_29876,N_29898);
nor UO_393 (O_393,N_29958,N_29667);
xnor UO_394 (O_394,N_29551,N_29530);
and UO_395 (O_395,N_29672,N_29635);
and UO_396 (O_396,N_29868,N_29512);
nand UO_397 (O_397,N_29738,N_29745);
and UO_398 (O_398,N_29528,N_29707);
nor UO_399 (O_399,N_29617,N_29936);
or UO_400 (O_400,N_29609,N_29661);
xnor UO_401 (O_401,N_29971,N_29811);
or UO_402 (O_402,N_29635,N_29688);
nor UO_403 (O_403,N_29706,N_29527);
nor UO_404 (O_404,N_29757,N_29954);
xnor UO_405 (O_405,N_29652,N_29929);
nand UO_406 (O_406,N_29616,N_29743);
nor UO_407 (O_407,N_29891,N_29761);
and UO_408 (O_408,N_29852,N_29737);
or UO_409 (O_409,N_29820,N_29986);
xor UO_410 (O_410,N_29828,N_29777);
nor UO_411 (O_411,N_29647,N_29623);
and UO_412 (O_412,N_29739,N_29601);
xor UO_413 (O_413,N_29578,N_29724);
and UO_414 (O_414,N_29765,N_29801);
nand UO_415 (O_415,N_29926,N_29672);
and UO_416 (O_416,N_29973,N_29526);
nor UO_417 (O_417,N_29659,N_29700);
xnor UO_418 (O_418,N_29614,N_29894);
nand UO_419 (O_419,N_29975,N_29526);
or UO_420 (O_420,N_29994,N_29779);
nand UO_421 (O_421,N_29935,N_29770);
or UO_422 (O_422,N_29579,N_29752);
or UO_423 (O_423,N_29846,N_29830);
xor UO_424 (O_424,N_29861,N_29620);
xnor UO_425 (O_425,N_29562,N_29768);
or UO_426 (O_426,N_29652,N_29704);
and UO_427 (O_427,N_29962,N_29880);
nand UO_428 (O_428,N_29901,N_29640);
nand UO_429 (O_429,N_29507,N_29584);
nor UO_430 (O_430,N_29623,N_29528);
nor UO_431 (O_431,N_29949,N_29766);
or UO_432 (O_432,N_29643,N_29943);
xor UO_433 (O_433,N_29929,N_29593);
nor UO_434 (O_434,N_29830,N_29602);
xnor UO_435 (O_435,N_29776,N_29982);
nor UO_436 (O_436,N_29700,N_29832);
nand UO_437 (O_437,N_29515,N_29626);
nand UO_438 (O_438,N_29591,N_29532);
nor UO_439 (O_439,N_29653,N_29668);
xor UO_440 (O_440,N_29932,N_29772);
and UO_441 (O_441,N_29915,N_29886);
nor UO_442 (O_442,N_29866,N_29888);
nor UO_443 (O_443,N_29616,N_29950);
nand UO_444 (O_444,N_29669,N_29979);
and UO_445 (O_445,N_29774,N_29732);
xnor UO_446 (O_446,N_29834,N_29515);
and UO_447 (O_447,N_29511,N_29788);
or UO_448 (O_448,N_29923,N_29625);
nor UO_449 (O_449,N_29875,N_29834);
nand UO_450 (O_450,N_29953,N_29716);
xnor UO_451 (O_451,N_29986,N_29670);
xnor UO_452 (O_452,N_29539,N_29538);
and UO_453 (O_453,N_29798,N_29636);
nor UO_454 (O_454,N_29582,N_29689);
xor UO_455 (O_455,N_29986,N_29709);
nor UO_456 (O_456,N_29581,N_29916);
or UO_457 (O_457,N_29857,N_29602);
nand UO_458 (O_458,N_29777,N_29973);
or UO_459 (O_459,N_29763,N_29855);
or UO_460 (O_460,N_29672,N_29535);
or UO_461 (O_461,N_29600,N_29826);
xnor UO_462 (O_462,N_29614,N_29963);
xnor UO_463 (O_463,N_29927,N_29925);
and UO_464 (O_464,N_29607,N_29943);
nor UO_465 (O_465,N_29901,N_29840);
nand UO_466 (O_466,N_29649,N_29997);
nor UO_467 (O_467,N_29907,N_29952);
and UO_468 (O_468,N_29803,N_29886);
nor UO_469 (O_469,N_29977,N_29766);
and UO_470 (O_470,N_29797,N_29519);
nand UO_471 (O_471,N_29777,N_29541);
or UO_472 (O_472,N_29729,N_29847);
nand UO_473 (O_473,N_29871,N_29961);
or UO_474 (O_474,N_29689,N_29963);
or UO_475 (O_475,N_29863,N_29555);
nand UO_476 (O_476,N_29589,N_29720);
and UO_477 (O_477,N_29587,N_29628);
and UO_478 (O_478,N_29986,N_29928);
nor UO_479 (O_479,N_29533,N_29833);
nand UO_480 (O_480,N_29753,N_29935);
nand UO_481 (O_481,N_29697,N_29880);
and UO_482 (O_482,N_29831,N_29929);
xor UO_483 (O_483,N_29688,N_29904);
nand UO_484 (O_484,N_29912,N_29908);
and UO_485 (O_485,N_29989,N_29752);
nor UO_486 (O_486,N_29724,N_29533);
nor UO_487 (O_487,N_29628,N_29990);
nand UO_488 (O_488,N_29886,N_29535);
and UO_489 (O_489,N_29525,N_29541);
nand UO_490 (O_490,N_29744,N_29530);
and UO_491 (O_491,N_29599,N_29500);
xnor UO_492 (O_492,N_29827,N_29502);
nor UO_493 (O_493,N_29822,N_29906);
and UO_494 (O_494,N_29958,N_29652);
or UO_495 (O_495,N_29844,N_29919);
xor UO_496 (O_496,N_29873,N_29918);
xnor UO_497 (O_497,N_29962,N_29619);
nand UO_498 (O_498,N_29657,N_29809);
xnor UO_499 (O_499,N_29830,N_29698);
nor UO_500 (O_500,N_29934,N_29779);
or UO_501 (O_501,N_29883,N_29612);
or UO_502 (O_502,N_29590,N_29950);
nor UO_503 (O_503,N_29518,N_29603);
or UO_504 (O_504,N_29795,N_29764);
xor UO_505 (O_505,N_29846,N_29868);
nand UO_506 (O_506,N_29539,N_29650);
nor UO_507 (O_507,N_29777,N_29991);
and UO_508 (O_508,N_29799,N_29692);
xor UO_509 (O_509,N_29780,N_29701);
nor UO_510 (O_510,N_29873,N_29504);
or UO_511 (O_511,N_29905,N_29763);
nand UO_512 (O_512,N_29842,N_29728);
xor UO_513 (O_513,N_29617,N_29707);
and UO_514 (O_514,N_29945,N_29576);
nand UO_515 (O_515,N_29749,N_29911);
and UO_516 (O_516,N_29987,N_29715);
nand UO_517 (O_517,N_29976,N_29719);
or UO_518 (O_518,N_29715,N_29511);
nor UO_519 (O_519,N_29822,N_29547);
nor UO_520 (O_520,N_29711,N_29685);
or UO_521 (O_521,N_29568,N_29696);
xor UO_522 (O_522,N_29697,N_29570);
and UO_523 (O_523,N_29885,N_29995);
nor UO_524 (O_524,N_29850,N_29642);
nor UO_525 (O_525,N_29752,N_29938);
or UO_526 (O_526,N_29615,N_29603);
nand UO_527 (O_527,N_29620,N_29602);
xor UO_528 (O_528,N_29925,N_29936);
xnor UO_529 (O_529,N_29661,N_29959);
nor UO_530 (O_530,N_29902,N_29813);
and UO_531 (O_531,N_29741,N_29628);
nor UO_532 (O_532,N_29830,N_29604);
nor UO_533 (O_533,N_29829,N_29765);
or UO_534 (O_534,N_29979,N_29872);
and UO_535 (O_535,N_29644,N_29883);
xnor UO_536 (O_536,N_29861,N_29577);
and UO_537 (O_537,N_29991,N_29594);
and UO_538 (O_538,N_29774,N_29994);
or UO_539 (O_539,N_29696,N_29907);
xnor UO_540 (O_540,N_29949,N_29575);
and UO_541 (O_541,N_29919,N_29808);
xnor UO_542 (O_542,N_29835,N_29827);
nor UO_543 (O_543,N_29566,N_29654);
nand UO_544 (O_544,N_29948,N_29943);
nor UO_545 (O_545,N_29631,N_29767);
xnor UO_546 (O_546,N_29557,N_29956);
or UO_547 (O_547,N_29611,N_29784);
nand UO_548 (O_548,N_29590,N_29942);
and UO_549 (O_549,N_29826,N_29584);
nand UO_550 (O_550,N_29761,N_29715);
and UO_551 (O_551,N_29779,N_29514);
nand UO_552 (O_552,N_29577,N_29721);
nor UO_553 (O_553,N_29681,N_29796);
nor UO_554 (O_554,N_29868,N_29591);
nand UO_555 (O_555,N_29853,N_29682);
and UO_556 (O_556,N_29664,N_29864);
xnor UO_557 (O_557,N_29989,N_29813);
or UO_558 (O_558,N_29681,N_29916);
nand UO_559 (O_559,N_29578,N_29623);
and UO_560 (O_560,N_29987,N_29659);
and UO_561 (O_561,N_29798,N_29912);
nor UO_562 (O_562,N_29865,N_29859);
xor UO_563 (O_563,N_29848,N_29566);
xor UO_564 (O_564,N_29956,N_29567);
and UO_565 (O_565,N_29850,N_29954);
and UO_566 (O_566,N_29831,N_29668);
or UO_567 (O_567,N_29767,N_29757);
or UO_568 (O_568,N_29535,N_29726);
xnor UO_569 (O_569,N_29524,N_29645);
nor UO_570 (O_570,N_29800,N_29774);
nand UO_571 (O_571,N_29896,N_29859);
nor UO_572 (O_572,N_29698,N_29521);
xnor UO_573 (O_573,N_29946,N_29930);
nand UO_574 (O_574,N_29643,N_29638);
or UO_575 (O_575,N_29570,N_29909);
xor UO_576 (O_576,N_29749,N_29521);
xor UO_577 (O_577,N_29836,N_29922);
nand UO_578 (O_578,N_29600,N_29741);
nor UO_579 (O_579,N_29877,N_29781);
nor UO_580 (O_580,N_29845,N_29758);
and UO_581 (O_581,N_29854,N_29691);
nand UO_582 (O_582,N_29622,N_29750);
and UO_583 (O_583,N_29952,N_29731);
nor UO_584 (O_584,N_29817,N_29959);
or UO_585 (O_585,N_29958,N_29925);
or UO_586 (O_586,N_29620,N_29564);
and UO_587 (O_587,N_29895,N_29736);
and UO_588 (O_588,N_29831,N_29700);
and UO_589 (O_589,N_29962,N_29650);
nor UO_590 (O_590,N_29920,N_29540);
and UO_591 (O_591,N_29825,N_29891);
or UO_592 (O_592,N_29842,N_29705);
nor UO_593 (O_593,N_29853,N_29812);
nor UO_594 (O_594,N_29521,N_29861);
or UO_595 (O_595,N_29993,N_29547);
nor UO_596 (O_596,N_29969,N_29873);
nor UO_597 (O_597,N_29944,N_29963);
nor UO_598 (O_598,N_29505,N_29968);
or UO_599 (O_599,N_29945,N_29925);
or UO_600 (O_600,N_29864,N_29589);
or UO_601 (O_601,N_29982,N_29966);
nand UO_602 (O_602,N_29658,N_29948);
nand UO_603 (O_603,N_29882,N_29528);
nand UO_604 (O_604,N_29652,N_29508);
nor UO_605 (O_605,N_29650,N_29641);
nand UO_606 (O_606,N_29907,N_29733);
nand UO_607 (O_607,N_29762,N_29678);
nor UO_608 (O_608,N_29578,N_29680);
nand UO_609 (O_609,N_29819,N_29997);
nand UO_610 (O_610,N_29792,N_29595);
nor UO_611 (O_611,N_29670,N_29769);
nor UO_612 (O_612,N_29566,N_29896);
and UO_613 (O_613,N_29784,N_29735);
xnor UO_614 (O_614,N_29945,N_29834);
nand UO_615 (O_615,N_29665,N_29789);
xor UO_616 (O_616,N_29696,N_29550);
and UO_617 (O_617,N_29892,N_29508);
and UO_618 (O_618,N_29956,N_29903);
xnor UO_619 (O_619,N_29570,N_29645);
or UO_620 (O_620,N_29661,N_29740);
nor UO_621 (O_621,N_29806,N_29797);
xnor UO_622 (O_622,N_29691,N_29525);
or UO_623 (O_623,N_29887,N_29777);
or UO_624 (O_624,N_29698,N_29782);
and UO_625 (O_625,N_29806,N_29830);
xor UO_626 (O_626,N_29556,N_29875);
nand UO_627 (O_627,N_29777,N_29755);
nor UO_628 (O_628,N_29925,N_29745);
xnor UO_629 (O_629,N_29630,N_29683);
nor UO_630 (O_630,N_29631,N_29616);
or UO_631 (O_631,N_29678,N_29575);
and UO_632 (O_632,N_29510,N_29831);
or UO_633 (O_633,N_29763,N_29788);
nor UO_634 (O_634,N_29552,N_29722);
xor UO_635 (O_635,N_29766,N_29664);
nor UO_636 (O_636,N_29651,N_29883);
nor UO_637 (O_637,N_29901,N_29725);
xnor UO_638 (O_638,N_29640,N_29905);
and UO_639 (O_639,N_29635,N_29940);
nand UO_640 (O_640,N_29852,N_29981);
nor UO_641 (O_641,N_29726,N_29943);
xnor UO_642 (O_642,N_29918,N_29972);
and UO_643 (O_643,N_29896,N_29956);
or UO_644 (O_644,N_29761,N_29800);
nor UO_645 (O_645,N_29638,N_29942);
nor UO_646 (O_646,N_29835,N_29953);
nor UO_647 (O_647,N_29555,N_29634);
or UO_648 (O_648,N_29953,N_29529);
nand UO_649 (O_649,N_29827,N_29993);
or UO_650 (O_650,N_29956,N_29913);
xor UO_651 (O_651,N_29585,N_29542);
nand UO_652 (O_652,N_29582,N_29722);
or UO_653 (O_653,N_29589,N_29705);
and UO_654 (O_654,N_29999,N_29983);
nand UO_655 (O_655,N_29719,N_29821);
and UO_656 (O_656,N_29525,N_29573);
nor UO_657 (O_657,N_29517,N_29884);
nor UO_658 (O_658,N_29611,N_29971);
or UO_659 (O_659,N_29682,N_29976);
xnor UO_660 (O_660,N_29808,N_29533);
nor UO_661 (O_661,N_29988,N_29518);
nor UO_662 (O_662,N_29512,N_29954);
xnor UO_663 (O_663,N_29760,N_29628);
or UO_664 (O_664,N_29857,N_29531);
or UO_665 (O_665,N_29566,N_29635);
xnor UO_666 (O_666,N_29729,N_29996);
nor UO_667 (O_667,N_29717,N_29824);
and UO_668 (O_668,N_29833,N_29982);
xor UO_669 (O_669,N_29754,N_29676);
and UO_670 (O_670,N_29959,N_29966);
or UO_671 (O_671,N_29723,N_29991);
or UO_672 (O_672,N_29824,N_29582);
nand UO_673 (O_673,N_29715,N_29769);
nand UO_674 (O_674,N_29688,N_29995);
xnor UO_675 (O_675,N_29916,N_29912);
nor UO_676 (O_676,N_29834,N_29854);
xor UO_677 (O_677,N_29705,N_29526);
and UO_678 (O_678,N_29827,N_29930);
nand UO_679 (O_679,N_29647,N_29856);
nand UO_680 (O_680,N_29790,N_29873);
and UO_681 (O_681,N_29684,N_29782);
nor UO_682 (O_682,N_29920,N_29982);
or UO_683 (O_683,N_29945,N_29821);
nand UO_684 (O_684,N_29583,N_29875);
nand UO_685 (O_685,N_29738,N_29928);
and UO_686 (O_686,N_29814,N_29792);
and UO_687 (O_687,N_29526,N_29675);
or UO_688 (O_688,N_29881,N_29542);
xor UO_689 (O_689,N_29673,N_29964);
or UO_690 (O_690,N_29905,N_29911);
nand UO_691 (O_691,N_29698,N_29553);
nor UO_692 (O_692,N_29832,N_29512);
nand UO_693 (O_693,N_29750,N_29840);
nor UO_694 (O_694,N_29846,N_29701);
nand UO_695 (O_695,N_29891,N_29658);
xor UO_696 (O_696,N_29664,N_29786);
nand UO_697 (O_697,N_29933,N_29623);
xor UO_698 (O_698,N_29600,N_29785);
nor UO_699 (O_699,N_29709,N_29610);
xnor UO_700 (O_700,N_29651,N_29741);
or UO_701 (O_701,N_29707,N_29554);
nor UO_702 (O_702,N_29783,N_29622);
xnor UO_703 (O_703,N_29615,N_29630);
nor UO_704 (O_704,N_29759,N_29502);
nor UO_705 (O_705,N_29852,N_29575);
and UO_706 (O_706,N_29766,N_29534);
xor UO_707 (O_707,N_29560,N_29855);
nand UO_708 (O_708,N_29926,N_29700);
nand UO_709 (O_709,N_29853,N_29696);
nor UO_710 (O_710,N_29993,N_29766);
or UO_711 (O_711,N_29975,N_29741);
nor UO_712 (O_712,N_29983,N_29893);
nand UO_713 (O_713,N_29929,N_29772);
or UO_714 (O_714,N_29563,N_29761);
nand UO_715 (O_715,N_29618,N_29864);
and UO_716 (O_716,N_29526,N_29987);
or UO_717 (O_717,N_29772,N_29718);
and UO_718 (O_718,N_29539,N_29707);
nand UO_719 (O_719,N_29619,N_29935);
nor UO_720 (O_720,N_29521,N_29680);
or UO_721 (O_721,N_29756,N_29698);
or UO_722 (O_722,N_29714,N_29600);
nand UO_723 (O_723,N_29811,N_29725);
or UO_724 (O_724,N_29822,N_29664);
nor UO_725 (O_725,N_29631,N_29941);
or UO_726 (O_726,N_29656,N_29810);
nor UO_727 (O_727,N_29541,N_29877);
and UO_728 (O_728,N_29638,N_29838);
nand UO_729 (O_729,N_29633,N_29598);
and UO_730 (O_730,N_29911,N_29588);
and UO_731 (O_731,N_29782,N_29794);
and UO_732 (O_732,N_29794,N_29606);
and UO_733 (O_733,N_29933,N_29589);
nor UO_734 (O_734,N_29925,N_29543);
nand UO_735 (O_735,N_29947,N_29504);
xor UO_736 (O_736,N_29910,N_29595);
or UO_737 (O_737,N_29880,N_29639);
and UO_738 (O_738,N_29825,N_29688);
nand UO_739 (O_739,N_29726,N_29963);
nand UO_740 (O_740,N_29701,N_29575);
and UO_741 (O_741,N_29707,N_29572);
and UO_742 (O_742,N_29670,N_29823);
or UO_743 (O_743,N_29675,N_29685);
or UO_744 (O_744,N_29586,N_29952);
or UO_745 (O_745,N_29535,N_29928);
and UO_746 (O_746,N_29793,N_29686);
and UO_747 (O_747,N_29823,N_29985);
nor UO_748 (O_748,N_29668,N_29592);
nand UO_749 (O_749,N_29997,N_29696);
nor UO_750 (O_750,N_29953,N_29637);
and UO_751 (O_751,N_29718,N_29524);
or UO_752 (O_752,N_29918,N_29726);
and UO_753 (O_753,N_29598,N_29876);
nor UO_754 (O_754,N_29775,N_29932);
or UO_755 (O_755,N_29602,N_29694);
nor UO_756 (O_756,N_29780,N_29776);
nor UO_757 (O_757,N_29739,N_29656);
nor UO_758 (O_758,N_29849,N_29885);
nand UO_759 (O_759,N_29570,N_29743);
or UO_760 (O_760,N_29564,N_29922);
and UO_761 (O_761,N_29900,N_29742);
and UO_762 (O_762,N_29760,N_29734);
nor UO_763 (O_763,N_29833,N_29950);
xor UO_764 (O_764,N_29787,N_29625);
nand UO_765 (O_765,N_29693,N_29666);
and UO_766 (O_766,N_29658,N_29597);
and UO_767 (O_767,N_29813,N_29895);
and UO_768 (O_768,N_29678,N_29536);
xnor UO_769 (O_769,N_29835,N_29563);
and UO_770 (O_770,N_29917,N_29919);
xor UO_771 (O_771,N_29840,N_29688);
or UO_772 (O_772,N_29857,N_29591);
nor UO_773 (O_773,N_29933,N_29765);
nor UO_774 (O_774,N_29978,N_29802);
or UO_775 (O_775,N_29772,N_29884);
nor UO_776 (O_776,N_29902,N_29523);
nor UO_777 (O_777,N_29681,N_29999);
or UO_778 (O_778,N_29584,N_29605);
xnor UO_779 (O_779,N_29845,N_29533);
and UO_780 (O_780,N_29868,N_29991);
xnor UO_781 (O_781,N_29802,N_29636);
or UO_782 (O_782,N_29808,N_29794);
or UO_783 (O_783,N_29508,N_29653);
nor UO_784 (O_784,N_29969,N_29906);
nor UO_785 (O_785,N_29803,N_29856);
xor UO_786 (O_786,N_29777,N_29628);
nor UO_787 (O_787,N_29607,N_29713);
nor UO_788 (O_788,N_29985,N_29875);
and UO_789 (O_789,N_29967,N_29565);
and UO_790 (O_790,N_29547,N_29773);
nand UO_791 (O_791,N_29766,N_29898);
and UO_792 (O_792,N_29742,N_29943);
and UO_793 (O_793,N_29902,N_29790);
nand UO_794 (O_794,N_29714,N_29544);
and UO_795 (O_795,N_29750,N_29955);
nor UO_796 (O_796,N_29926,N_29712);
xor UO_797 (O_797,N_29529,N_29510);
xnor UO_798 (O_798,N_29616,N_29899);
and UO_799 (O_799,N_29938,N_29940);
nand UO_800 (O_800,N_29877,N_29991);
xnor UO_801 (O_801,N_29654,N_29818);
or UO_802 (O_802,N_29931,N_29741);
xor UO_803 (O_803,N_29654,N_29726);
or UO_804 (O_804,N_29573,N_29575);
nor UO_805 (O_805,N_29948,N_29699);
and UO_806 (O_806,N_29991,N_29834);
or UO_807 (O_807,N_29896,N_29698);
xor UO_808 (O_808,N_29671,N_29632);
and UO_809 (O_809,N_29965,N_29572);
and UO_810 (O_810,N_29612,N_29528);
nand UO_811 (O_811,N_29549,N_29675);
nor UO_812 (O_812,N_29931,N_29610);
nor UO_813 (O_813,N_29997,N_29637);
and UO_814 (O_814,N_29986,N_29963);
xor UO_815 (O_815,N_29747,N_29704);
xor UO_816 (O_816,N_29957,N_29648);
xor UO_817 (O_817,N_29962,N_29934);
or UO_818 (O_818,N_29772,N_29792);
nand UO_819 (O_819,N_29805,N_29778);
nand UO_820 (O_820,N_29627,N_29576);
xor UO_821 (O_821,N_29739,N_29709);
xnor UO_822 (O_822,N_29912,N_29552);
and UO_823 (O_823,N_29910,N_29650);
or UO_824 (O_824,N_29527,N_29820);
and UO_825 (O_825,N_29501,N_29863);
nor UO_826 (O_826,N_29767,N_29922);
or UO_827 (O_827,N_29588,N_29992);
and UO_828 (O_828,N_29766,N_29927);
or UO_829 (O_829,N_29542,N_29624);
nand UO_830 (O_830,N_29507,N_29845);
nand UO_831 (O_831,N_29692,N_29733);
xnor UO_832 (O_832,N_29579,N_29672);
xnor UO_833 (O_833,N_29853,N_29599);
xor UO_834 (O_834,N_29923,N_29896);
xnor UO_835 (O_835,N_29993,N_29842);
or UO_836 (O_836,N_29556,N_29859);
or UO_837 (O_837,N_29919,N_29562);
nand UO_838 (O_838,N_29977,N_29504);
and UO_839 (O_839,N_29912,N_29727);
nor UO_840 (O_840,N_29653,N_29690);
nand UO_841 (O_841,N_29607,N_29996);
nor UO_842 (O_842,N_29702,N_29625);
nor UO_843 (O_843,N_29592,N_29515);
nor UO_844 (O_844,N_29850,N_29823);
xor UO_845 (O_845,N_29773,N_29563);
and UO_846 (O_846,N_29897,N_29515);
nor UO_847 (O_847,N_29794,N_29537);
nor UO_848 (O_848,N_29984,N_29581);
xnor UO_849 (O_849,N_29571,N_29619);
nand UO_850 (O_850,N_29604,N_29535);
and UO_851 (O_851,N_29879,N_29632);
xor UO_852 (O_852,N_29839,N_29621);
and UO_853 (O_853,N_29835,N_29797);
or UO_854 (O_854,N_29989,N_29909);
or UO_855 (O_855,N_29982,N_29932);
or UO_856 (O_856,N_29606,N_29602);
and UO_857 (O_857,N_29919,N_29604);
nand UO_858 (O_858,N_29814,N_29696);
and UO_859 (O_859,N_29586,N_29656);
nand UO_860 (O_860,N_29834,N_29663);
nor UO_861 (O_861,N_29910,N_29999);
nand UO_862 (O_862,N_29878,N_29762);
nor UO_863 (O_863,N_29663,N_29570);
nor UO_864 (O_864,N_29926,N_29575);
xor UO_865 (O_865,N_29987,N_29947);
or UO_866 (O_866,N_29621,N_29581);
nand UO_867 (O_867,N_29771,N_29653);
or UO_868 (O_868,N_29941,N_29704);
nor UO_869 (O_869,N_29915,N_29651);
or UO_870 (O_870,N_29965,N_29903);
and UO_871 (O_871,N_29804,N_29634);
or UO_872 (O_872,N_29828,N_29610);
xnor UO_873 (O_873,N_29536,N_29686);
nor UO_874 (O_874,N_29777,N_29963);
nand UO_875 (O_875,N_29911,N_29785);
or UO_876 (O_876,N_29804,N_29776);
or UO_877 (O_877,N_29701,N_29995);
nor UO_878 (O_878,N_29870,N_29933);
and UO_879 (O_879,N_29972,N_29939);
xnor UO_880 (O_880,N_29825,N_29767);
or UO_881 (O_881,N_29999,N_29628);
or UO_882 (O_882,N_29519,N_29540);
and UO_883 (O_883,N_29523,N_29970);
nor UO_884 (O_884,N_29910,N_29849);
nor UO_885 (O_885,N_29886,N_29822);
or UO_886 (O_886,N_29810,N_29967);
and UO_887 (O_887,N_29751,N_29733);
xor UO_888 (O_888,N_29677,N_29518);
nor UO_889 (O_889,N_29938,N_29560);
and UO_890 (O_890,N_29768,N_29890);
nor UO_891 (O_891,N_29568,N_29517);
xnor UO_892 (O_892,N_29779,N_29970);
nor UO_893 (O_893,N_29964,N_29928);
nor UO_894 (O_894,N_29803,N_29719);
xnor UO_895 (O_895,N_29935,N_29657);
xnor UO_896 (O_896,N_29736,N_29954);
nand UO_897 (O_897,N_29677,N_29604);
xnor UO_898 (O_898,N_29900,N_29832);
or UO_899 (O_899,N_29742,N_29920);
xor UO_900 (O_900,N_29590,N_29952);
or UO_901 (O_901,N_29841,N_29607);
nor UO_902 (O_902,N_29568,N_29868);
xnor UO_903 (O_903,N_29574,N_29613);
nand UO_904 (O_904,N_29648,N_29512);
and UO_905 (O_905,N_29843,N_29714);
or UO_906 (O_906,N_29910,N_29522);
nor UO_907 (O_907,N_29892,N_29839);
or UO_908 (O_908,N_29552,N_29864);
nor UO_909 (O_909,N_29848,N_29954);
xor UO_910 (O_910,N_29785,N_29750);
or UO_911 (O_911,N_29893,N_29976);
or UO_912 (O_912,N_29949,N_29563);
or UO_913 (O_913,N_29521,N_29876);
xor UO_914 (O_914,N_29591,N_29924);
or UO_915 (O_915,N_29727,N_29554);
nor UO_916 (O_916,N_29836,N_29623);
nand UO_917 (O_917,N_29725,N_29698);
nand UO_918 (O_918,N_29627,N_29823);
nand UO_919 (O_919,N_29900,N_29796);
xor UO_920 (O_920,N_29772,N_29626);
or UO_921 (O_921,N_29585,N_29778);
or UO_922 (O_922,N_29612,N_29841);
nand UO_923 (O_923,N_29680,N_29928);
and UO_924 (O_924,N_29941,N_29665);
xnor UO_925 (O_925,N_29709,N_29828);
nor UO_926 (O_926,N_29503,N_29649);
or UO_927 (O_927,N_29686,N_29857);
xor UO_928 (O_928,N_29875,N_29860);
nor UO_929 (O_929,N_29700,N_29974);
xor UO_930 (O_930,N_29825,N_29845);
nand UO_931 (O_931,N_29664,N_29713);
or UO_932 (O_932,N_29713,N_29762);
and UO_933 (O_933,N_29588,N_29741);
or UO_934 (O_934,N_29857,N_29539);
xnor UO_935 (O_935,N_29766,N_29857);
and UO_936 (O_936,N_29794,N_29925);
and UO_937 (O_937,N_29501,N_29884);
xor UO_938 (O_938,N_29741,N_29550);
nor UO_939 (O_939,N_29529,N_29636);
or UO_940 (O_940,N_29715,N_29899);
nand UO_941 (O_941,N_29822,N_29711);
xnor UO_942 (O_942,N_29776,N_29541);
nand UO_943 (O_943,N_29644,N_29910);
nand UO_944 (O_944,N_29928,N_29903);
and UO_945 (O_945,N_29851,N_29722);
nand UO_946 (O_946,N_29710,N_29656);
or UO_947 (O_947,N_29739,N_29973);
xor UO_948 (O_948,N_29562,N_29997);
nand UO_949 (O_949,N_29574,N_29834);
or UO_950 (O_950,N_29714,N_29869);
or UO_951 (O_951,N_29902,N_29720);
xnor UO_952 (O_952,N_29571,N_29813);
and UO_953 (O_953,N_29965,N_29660);
or UO_954 (O_954,N_29577,N_29789);
and UO_955 (O_955,N_29563,N_29580);
xor UO_956 (O_956,N_29949,N_29531);
xor UO_957 (O_957,N_29859,N_29520);
nor UO_958 (O_958,N_29951,N_29827);
or UO_959 (O_959,N_29541,N_29605);
xor UO_960 (O_960,N_29602,N_29752);
or UO_961 (O_961,N_29706,N_29628);
nor UO_962 (O_962,N_29984,N_29588);
and UO_963 (O_963,N_29859,N_29578);
and UO_964 (O_964,N_29532,N_29637);
and UO_965 (O_965,N_29854,N_29584);
nand UO_966 (O_966,N_29805,N_29712);
and UO_967 (O_967,N_29651,N_29736);
nor UO_968 (O_968,N_29696,N_29949);
and UO_969 (O_969,N_29922,N_29910);
xnor UO_970 (O_970,N_29911,N_29833);
xnor UO_971 (O_971,N_29816,N_29709);
xnor UO_972 (O_972,N_29509,N_29738);
xor UO_973 (O_973,N_29814,N_29773);
or UO_974 (O_974,N_29945,N_29716);
or UO_975 (O_975,N_29763,N_29932);
or UO_976 (O_976,N_29712,N_29919);
and UO_977 (O_977,N_29793,N_29601);
nor UO_978 (O_978,N_29732,N_29960);
nand UO_979 (O_979,N_29621,N_29619);
xor UO_980 (O_980,N_29777,N_29884);
xor UO_981 (O_981,N_29556,N_29988);
and UO_982 (O_982,N_29764,N_29640);
nand UO_983 (O_983,N_29665,N_29745);
nand UO_984 (O_984,N_29804,N_29546);
or UO_985 (O_985,N_29518,N_29577);
nor UO_986 (O_986,N_29732,N_29536);
nand UO_987 (O_987,N_29812,N_29674);
nand UO_988 (O_988,N_29526,N_29977);
nand UO_989 (O_989,N_29642,N_29927);
xnor UO_990 (O_990,N_29693,N_29994);
or UO_991 (O_991,N_29764,N_29999);
nand UO_992 (O_992,N_29797,N_29625);
or UO_993 (O_993,N_29605,N_29835);
nand UO_994 (O_994,N_29548,N_29796);
or UO_995 (O_995,N_29742,N_29635);
xor UO_996 (O_996,N_29762,N_29850);
xnor UO_997 (O_997,N_29630,N_29568);
xnor UO_998 (O_998,N_29562,N_29800);
or UO_999 (O_999,N_29718,N_29810);
and UO_1000 (O_1000,N_29882,N_29745);
nor UO_1001 (O_1001,N_29910,N_29784);
nand UO_1002 (O_1002,N_29701,N_29538);
xor UO_1003 (O_1003,N_29610,N_29538);
or UO_1004 (O_1004,N_29704,N_29810);
nand UO_1005 (O_1005,N_29720,N_29638);
nand UO_1006 (O_1006,N_29931,N_29947);
or UO_1007 (O_1007,N_29793,N_29575);
or UO_1008 (O_1008,N_29792,N_29888);
xor UO_1009 (O_1009,N_29716,N_29510);
and UO_1010 (O_1010,N_29933,N_29522);
or UO_1011 (O_1011,N_29681,N_29598);
and UO_1012 (O_1012,N_29873,N_29894);
nor UO_1013 (O_1013,N_29868,N_29606);
or UO_1014 (O_1014,N_29906,N_29691);
and UO_1015 (O_1015,N_29683,N_29961);
xnor UO_1016 (O_1016,N_29521,N_29568);
nand UO_1017 (O_1017,N_29968,N_29592);
or UO_1018 (O_1018,N_29904,N_29662);
and UO_1019 (O_1019,N_29955,N_29861);
or UO_1020 (O_1020,N_29693,N_29951);
xnor UO_1021 (O_1021,N_29806,N_29570);
and UO_1022 (O_1022,N_29817,N_29855);
xor UO_1023 (O_1023,N_29693,N_29690);
and UO_1024 (O_1024,N_29566,N_29702);
or UO_1025 (O_1025,N_29872,N_29886);
or UO_1026 (O_1026,N_29861,N_29678);
nand UO_1027 (O_1027,N_29693,N_29548);
nor UO_1028 (O_1028,N_29543,N_29626);
or UO_1029 (O_1029,N_29508,N_29693);
nand UO_1030 (O_1030,N_29860,N_29687);
or UO_1031 (O_1031,N_29700,N_29680);
xor UO_1032 (O_1032,N_29613,N_29661);
nand UO_1033 (O_1033,N_29511,N_29654);
xnor UO_1034 (O_1034,N_29935,N_29805);
or UO_1035 (O_1035,N_29679,N_29928);
nor UO_1036 (O_1036,N_29575,N_29572);
or UO_1037 (O_1037,N_29663,N_29647);
nand UO_1038 (O_1038,N_29921,N_29785);
xor UO_1039 (O_1039,N_29816,N_29528);
or UO_1040 (O_1040,N_29685,N_29530);
xnor UO_1041 (O_1041,N_29748,N_29825);
or UO_1042 (O_1042,N_29903,N_29979);
xor UO_1043 (O_1043,N_29611,N_29881);
and UO_1044 (O_1044,N_29843,N_29543);
xnor UO_1045 (O_1045,N_29744,N_29612);
nand UO_1046 (O_1046,N_29800,N_29799);
nand UO_1047 (O_1047,N_29864,N_29931);
and UO_1048 (O_1048,N_29996,N_29854);
and UO_1049 (O_1049,N_29638,N_29878);
xor UO_1050 (O_1050,N_29756,N_29630);
xor UO_1051 (O_1051,N_29949,N_29673);
or UO_1052 (O_1052,N_29874,N_29913);
xor UO_1053 (O_1053,N_29772,N_29890);
or UO_1054 (O_1054,N_29997,N_29792);
nand UO_1055 (O_1055,N_29606,N_29876);
nor UO_1056 (O_1056,N_29589,N_29932);
nand UO_1057 (O_1057,N_29920,N_29621);
nor UO_1058 (O_1058,N_29734,N_29600);
xor UO_1059 (O_1059,N_29984,N_29528);
and UO_1060 (O_1060,N_29677,N_29782);
nand UO_1061 (O_1061,N_29804,N_29521);
or UO_1062 (O_1062,N_29761,N_29846);
nand UO_1063 (O_1063,N_29891,N_29965);
xor UO_1064 (O_1064,N_29861,N_29728);
or UO_1065 (O_1065,N_29866,N_29605);
nor UO_1066 (O_1066,N_29996,N_29560);
xor UO_1067 (O_1067,N_29893,N_29776);
xnor UO_1068 (O_1068,N_29815,N_29593);
or UO_1069 (O_1069,N_29598,N_29769);
and UO_1070 (O_1070,N_29718,N_29510);
nor UO_1071 (O_1071,N_29909,N_29765);
or UO_1072 (O_1072,N_29831,N_29804);
and UO_1073 (O_1073,N_29592,N_29986);
xnor UO_1074 (O_1074,N_29520,N_29987);
nand UO_1075 (O_1075,N_29947,N_29627);
and UO_1076 (O_1076,N_29984,N_29761);
xnor UO_1077 (O_1077,N_29932,N_29801);
or UO_1078 (O_1078,N_29700,N_29558);
nand UO_1079 (O_1079,N_29831,N_29538);
or UO_1080 (O_1080,N_29606,N_29982);
nor UO_1081 (O_1081,N_29669,N_29831);
nand UO_1082 (O_1082,N_29759,N_29897);
xor UO_1083 (O_1083,N_29669,N_29747);
xnor UO_1084 (O_1084,N_29513,N_29642);
nand UO_1085 (O_1085,N_29564,N_29670);
and UO_1086 (O_1086,N_29851,N_29682);
nand UO_1087 (O_1087,N_29928,N_29958);
nor UO_1088 (O_1088,N_29692,N_29515);
nor UO_1089 (O_1089,N_29666,N_29532);
or UO_1090 (O_1090,N_29637,N_29623);
nor UO_1091 (O_1091,N_29632,N_29635);
and UO_1092 (O_1092,N_29950,N_29668);
xor UO_1093 (O_1093,N_29776,N_29540);
or UO_1094 (O_1094,N_29887,N_29542);
xnor UO_1095 (O_1095,N_29893,N_29836);
nand UO_1096 (O_1096,N_29917,N_29996);
and UO_1097 (O_1097,N_29585,N_29761);
or UO_1098 (O_1098,N_29604,N_29693);
xnor UO_1099 (O_1099,N_29689,N_29505);
nand UO_1100 (O_1100,N_29711,N_29986);
xnor UO_1101 (O_1101,N_29790,N_29509);
xor UO_1102 (O_1102,N_29855,N_29551);
and UO_1103 (O_1103,N_29552,N_29783);
nor UO_1104 (O_1104,N_29712,N_29977);
and UO_1105 (O_1105,N_29994,N_29715);
nand UO_1106 (O_1106,N_29751,N_29641);
nor UO_1107 (O_1107,N_29812,N_29755);
or UO_1108 (O_1108,N_29694,N_29759);
or UO_1109 (O_1109,N_29627,N_29578);
xor UO_1110 (O_1110,N_29607,N_29629);
xnor UO_1111 (O_1111,N_29968,N_29876);
and UO_1112 (O_1112,N_29632,N_29806);
and UO_1113 (O_1113,N_29989,N_29654);
and UO_1114 (O_1114,N_29735,N_29727);
xor UO_1115 (O_1115,N_29809,N_29544);
nand UO_1116 (O_1116,N_29781,N_29616);
and UO_1117 (O_1117,N_29639,N_29789);
nor UO_1118 (O_1118,N_29791,N_29962);
xor UO_1119 (O_1119,N_29881,N_29857);
or UO_1120 (O_1120,N_29979,N_29623);
nor UO_1121 (O_1121,N_29910,N_29500);
nand UO_1122 (O_1122,N_29665,N_29568);
xnor UO_1123 (O_1123,N_29975,N_29751);
nand UO_1124 (O_1124,N_29886,N_29667);
or UO_1125 (O_1125,N_29945,N_29967);
nand UO_1126 (O_1126,N_29924,N_29624);
and UO_1127 (O_1127,N_29933,N_29869);
nand UO_1128 (O_1128,N_29979,N_29604);
xnor UO_1129 (O_1129,N_29809,N_29923);
nor UO_1130 (O_1130,N_29723,N_29816);
nor UO_1131 (O_1131,N_29869,N_29600);
nand UO_1132 (O_1132,N_29930,N_29784);
xnor UO_1133 (O_1133,N_29681,N_29552);
or UO_1134 (O_1134,N_29592,N_29589);
or UO_1135 (O_1135,N_29763,N_29693);
and UO_1136 (O_1136,N_29652,N_29741);
xnor UO_1137 (O_1137,N_29652,N_29646);
and UO_1138 (O_1138,N_29608,N_29560);
or UO_1139 (O_1139,N_29873,N_29628);
or UO_1140 (O_1140,N_29575,N_29735);
xor UO_1141 (O_1141,N_29752,N_29695);
nand UO_1142 (O_1142,N_29731,N_29675);
nor UO_1143 (O_1143,N_29666,N_29682);
nor UO_1144 (O_1144,N_29653,N_29679);
nand UO_1145 (O_1145,N_29606,N_29541);
xnor UO_1146 (O_1146,N_29719,N_29895);
and UO_1147 (O_1147,N_29665,N_29562);
nor UO_1148 (O_1148,N_29963,N_29643);
and UO_1149 (O_1149,N_29521,N_29553);
and UO_1150 (O_1150,N_29532,N_29519);
nand UO_1151 (O_1151,N_29509,N_29610);
xor UO_1152 (O_1152,N_29919,N_29563);
xnor UO_1153 (O_1153,N_29798,N_29962);
nor UO_1154 (O_1154,N_29682,N_29807);
and UO_1155 (O_1155,N_29879,N_29710);
nor UO_1156 (O_1156,N_29842,N_29932);
and UO_1157 (O_1157,N_29907,N_29541);
and UO_1158 (O_1158,N_29755,N_29527);
or UO_1159 (O_1159,N_29615,N_29713);
nor UO_1160 (O_1160,N_29902,N_29819);
nor UO_1161 (O_1161,N_29558,N_29663);
xnor UO_1162 (O_1162,N_29806,N_29991);
and UO_1163 (O_1163,N_29525,N_29714);
and UO_1164 (O_1164,N_29559,N_29817);
xor UO_1165 (O_1165,N_29688,N_29826);
xnor UO_1166 (O_1166,N_29898,N_29908);
xnor UO_1167 (O_1167,N_29574,N_29936);
nor UO_1168 (O_1168,N_29939,N_29855);
or UO_1169 (O_1169,N_29555,N_29942);
or UO_1170 (O_1170,N_29891,N_29509);
and UO_1171 (O_1171,N_29723,N_29725);
or UO_1172 (O_1172,N_29628,N_29585);
nand UO_1173 (O_1173,N_29810,N_29593);
and UO_1174 (O_1174,N_29577,N_29635);
or UO_1175 (O_1175,N_29982,N_29544);
or UO_1176 (O_1176,N_29545,N_29982);
nor UO_1177 (O_1177,N_29746,N_29673);
xnor UO_1178 (O_1178,N_29780,N_29764);
nand UO_1179 (O_1179,N_29909,N_29655);
nor UO_1180 (O_1180,N_29795,N_29641);
xor UO_1181 (O_1181,N_29509,N_29756);
or UO_1182 (O_1182,N_29966,N_29698);
nand UO_1183 (O_1183,N_29889,N_29669);
xor UO_1184 (O_1184,N_29519,N_29561);
or UO_1185 (O_1185,N_29964,N_29933);
nor UO_1186 (O_1186,N_29796,N_29866);
xor UO_1187 (O_1187,N_29893,N_29736);
or UO_1188 (O_1188,N_29710,N_29864);
nor UO_1189 (O_1189,N_29738,N_29811);
xnor UO_1190 (O_1190,N_29686,N_29811);
nor UO_1191 (O_1191,N_29878,N_29788);
nand UO_1192 (O_1192,N_29855,N_29872);
nor UO_1193 (O_1193,N_29593,N_29867);
and UO_1194 (O_1194,N_29630,N_29554);
nand UO_1195 (O_1195,N_29753,N_29696);
xor UO_1196 (O_1196,N_29589,N_29803);
nor UO_1197 (O_1197,N_29685,N_29651);
or UO_1198 (O_1198,N_29865,N_29611);
or UO_1199 (O_1199,N_29507,N_29585);
nor UO_1200 (O_1200,N_29977,N_29663);
and UO_1201 (O_1201,N_29903,N_29552);
nor UO_1202 (O_1202,N_29741,N_29578);
nor UO_1203 (O_1203,N_29560,N_29859);
and UO_1204 (O_1204,N_29682,N_29723);
xor UO_1205 (O_1205,N_29812,N_29539);
and UO_1206 (O_1206,N_29959,N_29873);
xor UO_1207 (O_1207,N_29861,N_29751);
nand UO_1208 (O_1208,N_29736,N_29555);
and UO_1209 (O_1209,N_29961,N_29990);
or UO_1210 (O_1210,N_29661,N_29517);
nand UO_1211 (O_1211,N_29711,N_29773);
nand UO_1212 (O_1212,N_29731,N_29874);
xor UO_1213 (O_1213,N_29698,N_29700);
and UO_1214 (O_1214,N_29963,N_29813);
or UO_1215 (O_1215,N_29649,N_29688);
and UO_1216 (O_1216,N_29691,N_29668);
or UO_1217 (O_1217,N_29678,N_29510);
or UO_1218 (O_1218,N_29713,N_29845);
nor UO_1219 (O_1219,N_29892,N_29953);
or UO_1220 (O_1220,N_29660,N_29711);
and UO_1221 (O_1221,N_29915,N_29730);
nor UO_1222 (O_1222,N_29514,N_29715);
or UO_1223 (O_1223,N_29773,N_29725);
nand UO_1224 (O_1224,N_29808,N_29769);
or UO_1225 (O_1225,N_29543,N_29579);
or UO_1226 (O_1226,N_29538,N_29752);
and UO_1227 (O_1227,N_29909,N_29507);
nand UO_1228 (O_1228,N_29929,N_29900);
nor UO_1229 (O_1229,N_29560,N_29737);
nand UO_1230 (O_1230,N_29886,N_29764);
nor UO_1231 (O_1231,N_29757,N_29789);
nand UO_1232 (O_1232,N_29656,N_29732);
or UO_1233 (O_1233,N_29951,N_29563);
nand UO_1234 (O_1234,N_29624,N_29926);
nand UO_1235 (O_1235,N_29537,N_29609);
xnor UO_1236 (O_1236,N_29640,N_29635);
nor UO_1237 (O_1237,N_29909,N_29806);
and UO_1238 (O_1238,N_29735,N_29547);
or UO_1239 (O_1239,N_29822,N_29829);
or UO_1240 (O_1240,N_29516,N_29592);
xor UO_1241 (O_1241,N_29617,N_29924);
or UO_1242 (O_1242,N_29717,N_29692);
nand UO_1243 (O_1243,N_29563,N_29622);
xnor UO_1244 (O_1244,N_29809,N_29987);
and UO_1245 (O_1245,N_29588,N_29725);
nand UO_1246 (O_1246,N_29686,N_29898);
and UO_1247 (O_1247,N_29897,N_29962);
or UO_1248 (O_1248,N_29647,N_29862);
nand UO_1249 (O_1249,N_29761,N_29885);
nor UO_1250 (O_1250,N_29723,N_29988);
nand UO_1251 (O_1251,N_29593,N_29909);
nand UO_1252 (O_1252,N_29754,N_29863);
and UO_1253 (O_1253,N_29908,N_29535);
xor UO_1254 (O_1254,N_29919,N_29713);
or UO_1255 (O_1255,N_29799,N_29755);
nor UO_1256 (O_1256,N_29605,N_29758);
xnor UO_1257 (O_1257,N_29579,N_29765);
or UO_1258 (O_1258,N_29727,N_29837);
or UO_1259 (O_1259,N_29534,N_29708);
xnor UO_1260 (O_1260,N_29567,N_29919);
xnor UO_1261 (O_1261,N_29504,N_29789);
or UO_1262 (O_1262,N_29559,N_29914);
nor UO_1263 (O_1263,N_29557,N_29590);
or UO_1264 (O_1264,N_29805,N_29890);
nand UO_1265 (O_1265,N_29950,N_29899);
and UO_1266 (O_1266,N_29825,N_29587);
nand UO_1267 (O_1267,N_29864,N_29950);
nor UO_1268 (O_1268,N_29818,N_29840);
nor UO_1269 (O_1269,N_29546,N_29507);
or UO_1270 (O_1270,N_29835,N_29883);
xor UO_1271 (O_1271,N_29619,N_29646);
or UO_1272 (O_1272,N_29729,N_29584);
xor UO_1273 (O_1273,N_29711,N_29946);
nor UO_1274 (O_1274,N_29938,N_29724);
nor UO_1275 (O_1275,N_29814,N_29939);
nor UO_1276 (O_1276,N_29662,N_29653);
and UO_1277 (O_1277,N_29623,N_29733);
and UO_1278 (O_1278,N_29583,N_29673);
nand UO_1279 (O_1279,N_29897,N_29806);
or UO_1280 (O_1280,N_29651,N_29931);
nand UO_1281 (O_1281,N_29680,N_29587);
nand UO_1282 (O_1282,N_29673,N_29625);
nand UO_1283 (O_1283,N_29891,N_29712);
nor UO_1284 (O_1284,N_29759,N_29835);
or UO_1285 (O_1285,N_29578,N_29792);
nor UO_1286 (O_1286,N_29690,N_29776);
or UO_1287 (O_1287,N_29651,N_29584);
and UO_1288 (O_1288,N_29975,N_29612);
nor UO_1289 (O_1289,N_29610,N_29707);
or UO_1290 (O_1290,N_29610,N_29500);
nor UO_1291 (O_1291,N_29578,N_29895);
nor UO_1292 (O_1292,N_29527,N_29589);
or UO_1293 (O_1293,N_29503,N_29875);
xnor UO_1294 (O_1294,N_29582,N_29700);
or UO_1295 (O_1295,N_29941,N_29543);
nand UO_1296 (O_1296,N_29984,N_29794);
and UO_1297 (O_1297,N_29709,N_29644);
xnor UO_1298 (O_1298,N_29822,N_29891);
and UO_1299 (O_1299,N_29967,N_29515);
or UO_1300 (O_1300,N_29895,N_29584);
and UO_1301 (O_1301,N_29674,N_29525);
nor UO_1302 (O_1302,N_29647,N_29957);
xnor UO_1303 (O_1303,N_29916,N_29730);
xor UO_1304 (O_1304,N_29696,N_29544);
nand UO_1305 (O_1305,N_29805,N_29563);
nor UO_1306 (O_1306,N_29916,N_29589);
nor UO_1307 (O_1307,N_29756,N_29889);
nand UO_1308 (O_1308,N_29611,N_29902);
xor UO_1309 (O_1309,N_29974,N_29770);
nor UO_1310 (O_1310,N_29695,N_29793);
nor UO_1311 (O_1311,N_29569,N_29875);
xor UO_1312 (O_1312,N_29967,N_29750);
nand UO_1313 (O_1313,N_29741,N_29713);
and UO_1314 (O_1314,N_29959,N_29553);
and UO_1315 (O_1315,N_29584,N_29661);
xor UO_1316 (O_1316,N_29727,N_29893);
or UO_1317 (O_1317,N_29795,N_29743);
xor UO_1318 (O_1318,N_29941,N_29675);
nand UO_1319 (O_1319,N_29659,N_29890);
and UO_1320 (O_1320,N_29605,N_29775);
xnor UO_1321 (O_1321,N_29820,N_29978);
and UO_1322 (O_1322,N_29974,N_29504);
xnor UO_1323 (O_1323,N_29912,N_29814);
nand UO_1324 (O_1324,N_29531,N_29509);
nor UO_1325 (O_1325,N_29908,N_29985);
nand UO_1326 (O_1326,N_29995,N_29696);
xnor UO_1327 (O_1327,N_29967,N_29753);
and UO_1328 (O_1328,N_29657,N_29712);
xnor UO_1329 (O_1329,N_29959,N_29902);
or UO_1330 (O_1330,N_29728,N_29561);
nor UO_1331 (O_1331,N_29795,N_29965);
nand UO_1332 (O_1332,N_29989,N_29983);
and UO_1333 (O_1333,N_29672,N_29867);
xor UO_1334 (O_1334,N_29880,N_29805);
nor UO_1335 (O_1335,N_29557,N_29968);
nor UO_1336 (O_1336,N_29728,N_29647);
nand UO_1337 (O_1337,N_29918,N_29553);
xor UO_1338 (O_1338,N_29704,N_29546);
nand UO_1339 (O_1339,N_29859,N_29602);
xor UO_1340 (O_1340,N_29567,N_29583);
xor UO_1341 (O_1341,N_29964,N_29558);
nor UO_1342 (O_1342,N_29967,N_29981);
nand UO_1343 (O_1343,N_29990,N_29605);
nor UO_1344 (O_1344,N_29922,N_29526);
xor UO_1345 (O_1345,N_29508,N_29758);
nor UO_1346 (O_1346,N_29984,N_29818);
and UO_1347 (O_1347,N_29541,N_29590);
nand UO_1348 (O_1348,N_29518,N_29700);
nor UO_1349 (O_1349,N_29774,N_29996);
and UO_1350 (O_1350,N_29639,N_29962);
or UO_1351 (O_1351,N_29704,N_29635);
and UO_1352 (O_1352,N_29980,N_29520);
nand UO_1353 (O_1353,N_29691,N_29596);
or UO_1354 (O_1354,N_29887,N_29511);
nand UO_1355 (O_1355,N_29519,N_29589);
nand UO_1356 (O_1356,N_29743,N_29686);
or UO_1357 (O_1357,N_29729,N_29505);
xor UO_1358 (O_1358,N_29850,N_29715);
or UO_1359 (O_1359,N_29905,N_29896);
nor UO_1360 (O_1360,N_29580,N_29545);
nor UO_1361 (O_1361,N_29511,N_29718);
xnor UO_1362 (O_1362,N_29799,N_29912);
nor UO_1363 (O_1363,N_29922,N_29877);
and UO_1364 (O_1364,N_29635,N_29619);
xnor UO_1365 (O_1365,N_29625,N_29533);
nand UO_1366 (O_1366,N_29877,N_29632);
nor UO_1367 (O_1367,N_29633,N_29534);
and UO_1368 (O_1368,N_29946,N_29697);
and UO_1369 (O_1369,N_29553,N_29626);
and UO_1370 (O_1370,N_29746,N_29535);
nor UO_1371 (O_1371,N_29655,N_29804);
xnor UO_1372 (O_1372,N_29658,N_29641);
or UO_1373 (O_1373,N_29552,N_29507);
xnor UO_1374 (O_1374,N_29836,N_29504);
xnor UO_1375 (O_1375,N_29957,N_29854);
and UO_1376 (O_1376,N_29701,N_29524);
or UO_1377 (O_1377,N_29754,N_29815);
xnor UO_1378 (O_1378,N_29572,N_29838);
nand UO_1379 (O_1379,N_29961,N_29829);
nand UO_1380 (O_1380,N_29526,N_29509);
xnor UO_1381 (O_1381,N_29799,N_29821);
and UO_1382 (O_1382,N_29717,N_29737);
xor UO_1383 (O_1383,N_29712,N_29600);
or UO_1384 (O_1384,N_29877,N_29911);
xnor UO_1385 (O_1385,N_29835,N_29606);
nand UO_1386 (O_1386,N_29529,N_29890);
nor UO_1387 (O_1387,N_29942,N_29955);
nand UO_1388 (O_1388,N_29608,N_29940);
nor UO_1389 (O_1389,N_29502,N_29865);
nor UO_1390 (O_1390,N_29645,N_29631);
or UO_1391 (O_1391,N_29982,N_29678);
xor UO_1392 (O_1392,N_29772,N_29560);
nor UO_1393 (O_1393,N_29681,N_29592);
and UO_1394 (O_1394,N_29772,N_29925);
xnor UO_1395 (O_1395,N_29845,N_29884);
nor UO_1396 (O_1396,N_29843,N_29555);
nand UO_1397 (O_1397,N_29974,N_29644);
and UO_1398 (O_1398,N_29978,N_29895);
and UO_1399 (O_1399,N_29634,N_29853);
nor UO_1400 (O_1400,N_29913,N_29919);
nor UO_1401 (O_1401,N_29842,N_29543);
nor UO_1402 (O_1402,N_29923,N_29689);
or UO_1403 (O_1403,N_29711,N_29823);
or UO_1404 (O_1404,N_29830,N_29758);
or UO_1405 (O_1405,N_29613,N_29653);
and UO_1406 (O_1406,N_29967,N_29815);
xnor UO_1407 (O_1407,N_29705,N_29632);
xor UO_1408 (O_1408,N_29574,N_29912);
xnor UO_1409 (O_1409,N_29708,N_29581);
or UO_1410 (O_1410,N_29879,N_29924);
xor UO_1411 (O_1411,N_29576,N_29846);
or UO_1412 (O_1412,N_29681,N_29593);
nor UO_1413 (O_1413,N_29610,N_29742);
or UO_1414 (O_1414,N_29540,N_29674);
and UO_1415 (O_1415,N_29972,N_29616);
or UO_1416 (O_1416,N_29686,N_29792);
nor UO_1417 (O_1417,N_29828,N_29632);
nand UO_1418 (O_1418,N_29756,N_29949);
and UO_1419 (O_1419,N_29716,N_29980);
and UO_1420 (O_1420,N_29554,N_29671);
nand UO_1421 (O_1421,N_29541,N_29837);
and UO_1422 (O_1422,N_29829,N_29784);
nand UO_1423 (O_1423,N_29811,N_29709);
and UO_1424 (O_1424,N_29564,N_29602);
nor UO_1425 (O_1425,N_29882,N_29878);
nand UO_1426 (O_1426,N_29727,N_29902);
or UO_1427 (O_1427,N_29980,N_29597);
nor UO_1428 (O_1428,N_29949,N_29731);
or UO_1429 (O_1429,N_29734,N_29889);
nor UO_1430 (O_1430,N_29509,N_29913);
nand UO_1431 (O_1431,N_29516,N_29719);
nor UO_1432 (O_1432,N_29674,N_29604);
and UO_1433 (O_1433,N_29500,N_29712);
or UO_1434 (O_1434,N_29521,N_29524);
nand UO_1435 (O_1435,N_29739,N_29906);
nor UO_1436 (O_1436,N_29550,N_29652);
and UO_1437 (O_1437,N_29623,N_29670);
nor UO_1438 (O_1438,N_29742,N_29884);
nand UO_1439 (O_1439,N_29572,N_29700);
nor UO_1440 (O_1440,N_29866,N_29828);
and UO_1441 (O_1441,N_29929,N_29930);
or UO_1442 (O_1442,N_29770,N_29780);
nor UO_1443 (O_1443,N_29695,N_29835);
xnor UO_1444 (O_1444,N_29962,N_29591);
nor UO_1445 (O_1445,N_29918,N_29937);
and UO_1446 (O_1446,N_29966,N_29908);
and UO_1447 (O_1447,N_29804,N_29887);
or UO_1448 (O_1448,N_29969,N_29710);
xor UO_1449 (O_1449,N_29894,N_29533);
nor UO_1450 (O_1450,N_29694,N_29904);
nor UO_1451 (O_1451,N_29863,N_29775);
xnor UO_1452 (O_1452,N_29618,N_29937);
and UO_1453 (O_1453,N_29543,N_29994);
xor UO_1454 (O_1454,N_29883,N_29822);
nor UO_1455 (O_1455,N_29664,N_29800);
or UO_1456 (O_1456,N_29732,N_29599);
nand UO_1457 (O_1457,N_29793,N_29569);
xnor UO_1458 (O_1458,N_29896,N_29546);
nand UO_1459 (O_1459,N_29825,N_29665);
or UO_1460 (O_1460,N_29990,N_29832);
xor UO_1461 (O_1461,N_29665,N_29987);
xnor UO_1462 (O_1462,N_29529,N_29633);
nand UO_1463 (O_1463,N_29912,N_29865);
nor UO_1464 (O_1464,N_29939,N_29505);
nand UO_1465 (O_1465,N_29917,N_29954);
and UO_1466 (O_1466,N_29806,N_29855);
and UO_1467 (O_1467,N_29602,N_29647);
and UO_1468 (O_1468,N_29835,N_29667);
or UO_1469 (O_1469,N_29543,N_29885);
nand UO_1470 (O_1470,N_29917,N_29681);
nand UO_1471 (O_1471,N_29691,N_29590);
or UO_1472 (O_1472,N_29875,N_29983);
xor UO_1473 (O_1473,N_29843,N_29641);
nand UO_1474 (O_1474,N_29826,N_29785);
nand UO_1475 (O_1475,N_29914,N_29955);
and UO_1476 (O_1476,N_29549,N_29625);
nand UO_1477 (O_1477,N_29510,N_29737);
and UO_1478 (O_1478,N_29913,N_29513);
nand UO_1479 (O_1479,N_29693,N_29702);
nand UO_1480 (O_1480,N_29517,N_29791);
nor UO_1481 (O_1481,N_29933,N_29643);
or UO_1482 (O_1482,N_29576,N_29650);
xor UO_1483 (O_1483,N_29888,N_29589);
xor UO_1484 (O_1484,N_29526,N_29658);
or UO_1485 (O_1485,N_29911,N_29551);
or UO_1486 (O_1486,N_29535,N_29643);
nor UO_1487 (O_1487,N_29930,N_29952);
nor UO_1488 (O_1488,N_29918,N_29632);
and UO_1489 (O_1489,N_29773,N_29614);
or UO_1490 (O_1490,N_29568,N_29564);
or UO_1491 (O_1491,N_29541,N_29920);
and UO_1492 (O_1492,N_29872,N_29936);
and UO_1493 (O_1493,N_29593,N_29878);
and UO_1494 (O_1494,N_29540,N_29584);
nor UO_1495 (O_1495,N_29573,N_29599);
xor UO_1496 (O_1496,N_29830,N_29934);
and UO_1497 (O_1497,N_29697,N_29652);
nor UO_1498 (O_1498,N_29822,N_29553);
xor UO_1499 (O_1499,N_29905,N_29973);
or UO_1500 (O_1500,N_29782,N_29754);
or UO_1501 (O_1501,N_29949,N_29518);
xor UO_1502 (O_1502,N_29962,N_29524);
nand UO_1503 (O_1503,N_29993,N_29638);
or UO_1504 (O_1504,N_29987,N_29814);
xnor UO_1505 (O_1505,N_29803,N_29526);
or UO_1506 (O_1506,N_29717,N_29900);
xnor UO_1507 (O_1507,N_29509,N_29613);
or UO_1508 (O_1508,N_29772,N_29578);
and UO_1509 (O_1509,N_29928,N_29732);
xnor UO_1510 (O_1510,N_29930,N_29657);
and UO_1511 (O_1511,N_29907,N_29818);
or UO_1512 (O_1512,N_29899,N_29976);
or UO_1513 (O_1513,N_29665,N_29510);
xnor UO_1514 (O_1514,N_29638,N_29783);
or UO_1515 (O_1515,N_29892,N_29965);
nor UO_1516 (O_1516,N_29678,N_29781);
nor UO_1517 (O_1517,N_29620,N_29835);
nand UO_1518 (O_1518,N_29676,N_29848);
xor UO_1519 (O_1519,N_29643,N_29704);
or UO_1520 (O_1520,N_29825,N_29931);
or UO_1521 (O_1521,N_29909,N_29952);
nor UO_1522 (O_1522,N_29947,N_29975);
nand UO_1523 (O_1523,N_29668,N_29860);
or UO_1524 (O_1524,N_29838,N_29599);
nor UO_1525 (O_1525,N_29660,N_29876);
xor UO_1526 (O_1526,N_29994,N_29652);
nand UO_1527 (O_1527,N_29587,N_29955);
and UO_1528 (O_1528,N_29602,N_29932);
nand UO_1529 (O_1529,N_29784,N_29883);
and UO_1530 (O_1530,N_29835,N_29665);
nor UO_1531 (O_1531,N_29558,N_29900);
nand UO_1532 (O_1532,N_29901,N_29566);
nor UO_1533 (O_1533,N_29722,N_29927);
nor UO_1534 (O_1534,N_29823,N_29878);
nand UO_1535 (O_1535,N_29741,N_29776);
nor UO_1536 (O_1536,N_29923,N_29573);
or UO_1537 (O_1537,N_29858,N_29738);
nor UO_1538 (O_1538,N_29896,N_29893);
nand UO_1539 (O_1539,N_29639,N_29940);
xnor UO_1540 (O_1540,N_29946,N_29608);
and UO_1541 (O_1541,N_29754,N_29970);
nand UO_1542 (O_1542,N_29902,N_29766);
or UO_1543 (O_1543,N_29767,N_29964);
xnor UO_1544 (O_1544,N_29721,N_29888);
xnor UO_1545 (O_1545,N_29545,N_29898);
nand UO_1546 (O_1546,N_29708,N_29982);
and UO_1547 (O_1547,N_29878,N_29722);
nor UO_1548 (O_1548,N_29979,N_29699);
xor UO_1549 (O_1549,N_29986,N_29979);
and UO_1550 (O_1550,N_29763,N_29507);
nand UO_1551 (O_1551,N_29713,N_29579);
or UO_1552 (O_1552,N_29846,N_29836);
nand UO_1553 (O_1553,N_29737,N_29660);
nand UO_1554 (O_1554,N_29838,N_29594);
xor UO_1555 (O_1555,N_29695,N_29649);
nor UO_1556 (O_1556,N_29664,N_29583);
xor UO_1557 (O_1557,N_29990,N_29878);
xnor UO_1558 (O_1558,N_29580,N_29993);
nor UO_1559 (O_1559,N_29854,N_29820);
nor UO_1560 (O_1560,N_29884,N_29671);
or UO_1561 (O_1561,N_29784,N_29965);
nand UO_1562 (O_1562,N_29625,N_29886);
nor UO_1563 (O_1563,N_29603,N_29609);
and UO_1564 (O_1564,N_29950,N_29528);
xnor UO_1565 (O_1565,N_29576,N_29581);
and UO_1566 (O_1566,N_29787,N_29853);
or UO_1567 (O_1567,N_29643,N_29968);
or UO_1568 (O_1568,N_29739,N_29961);
and UO_1569 (O_1569,N_29614,N_29848);
xnor UO_1570 (O_1570,N_29959,N_29518);
nand UO_1571 (O_1571,N_29648,N_29985);
and UO_1572 (O_1572,N_29648,N_29788);
xnor UO_1573 (O_1573,N_29563,N_29620);
or UO_1574 (O_1574,N_29760,N_29501);
nand UO_1575 (O_1575,N_29871,N_29657);
nor UO_1576 (O_1576,N_29790,N_29667);
nor UO_1577 (O_1577,N_29702,N_29737);
nand UO_1578 (O_1578,N_29767,N_29731);
nand UO_1579 (O_1579,N_29552,N_29721);
nand UO_1580 (O_1580,N_29690,N_29628);
xor UO_1581 (O_1581,N_29736,N_29797);
xor UO_1582 (O_1582,N_29923,N_29797);
nor UO_1583 (O_1583,N_29863,N_29826);
and UO_1584 (O_1584,N_29533,N_29692);
nor UO_1585 (O_1585,N_29957,N_29884);
and UO_1586 (O_1586,N_29621,N_29926);
nand UO_1587 (O_1587,N_29801,N_29974);
nor UO_1588 (O_1588,N_29617,N_29983);
or UO_1589 (O_1589,N_29830,N_29650);
or UO_1590 (O_1590,N_29774,N_29876);
or UO_1591 (O_1591,N_29588,N_29882);
nor UO_1592 (O_1592,N_29942,N_29817);
or UO_1593 (O_1593,N_29891,N_29793);
or UO_1594 (O_1594,N_29555,N_29636);
nor UO_1595 (O_1595,N_29617,N_29715);
nand UO_1596 (O_1596,N_29786,N_29649);
nor UO_1597 (O_1597,N_29669,N_29566);
xnor UO_1598 (O_1598,N_29728,N_29837);
nand UO_1599 (O_1599,N_29795,N_29606);
and UO_1600 (O_1600,N_29662,N_29840);
or UO_1601 (O_1601,N_29537,N_29811);
and UO_1602 (O_1602,N_29739,N_29747);
nor UO_1603 (O_1603,N_29888,N_29616);
nor UO_1604 (O_1604,N_29834,N_29738);
nand UO_1605 (O_1605,N_29708,N_29777);
and UO_1606 (O_1606,N_29569,N_29705);
and UO_1607 (O_1607,N_29906,N_29779);
nand UO_1608 (O_1608,N_29794,N_29619);
xor UO_1609 (O_1609,N_29527,N_29610);
nor UO_1610 (O_1610,N_29985,N_29621);
nor UO_1611 (O_1611,N_29515,N_29661);
xnor UO_1612 (O_1612,N_29985,N_29690);
nor UO_1613 (O_1613,N_29627,N_29795);
and UO_1614 (O_1614,N_29859,N_29608);
xnor UO_1615 (O_1615,N_29953,N_29719);
xnor UO_1616 (O_1616,N_29899,N_29645);
nor UO_1617 (O_1617,N_29866,N_29780);
nand UO_1618 (O_1618,N_29638,N_29804);
xor UO_1619 (O_1619,N_29836,N_29841);
nand UO_1620 (O_1620,N_29636,N_29586);
or UO_1621 (O_1621,N_29778,N_29650);
nand UO_1622 (O_1622,N_29508,N_29667);
or UO_1623 (O_1623,N_29965,N_29526);
xnor UO_1624 (O_1624,N_29918,N_29626);
nor UO_1625 (O_1625,N_29647,N_29943);
and UO_1626 (O_1626,N_29879,N_29671);
nor UO_1627 (O_1627,N_29652,N_29614);
nand UO_1628 (O_1628,N_29873,N_29958);
and UO_1629 (O_1629,N_29826,N_29805);
or UO_1630 (O_1630,N_29526,N_29902);
and UO_1631 (O_1631,N_29722,N_29747);
and UO_1632 (O_1632,N_29502,N_29560);
nor UO_1633 (O_1633,N_29789,N_29999);
or UO_1634 (O_1634,N_29842,N_29695);
nor UO_1635 (O_1635,N_29546,N_29968);
or UO_1636 (O_1636,N_29606,N_29851);
and UO_1637 (O_1637,N_29709,N_29818);
nand UO_1638 (O_1638,N_29628,N_29978);
nand UO_1639 (O_1639,N_29873,N_29938);
nand UO_1640 (O_1640,N_29706,N_29746);
nand UO_1641 (O_1641,N_29550,N_29812);
xnor UO_1642 (O_1642,N_29507,N_29748);
and UO_1643 (O_1643,N_29631,N_29918);
and UO_1644 (O_1644,N_29661,N_29742);
nand UO_1645 (O_1645,N_29829,N_29836);
and UO_1646 (O_1646,N_29759,N_29763);
xnor UO_1647 (O_1647,N_29529,N_29816);
and UO_1648 (O_1648,N_29991,N_29894);
nor UO_1649 (O_1649,N_29800,N_29642);
or UO_1650 (O_1650,N_29959,N_29579);
and UO_1651 (O_1651,N_29979,N_29861);
xnor UO_1652 (O_1652,N_29692,N_29583);
nand UO_1653 (O_1653,N_29725,N_29847);
nor UO_1654 (O_1654,N_29700,N_29726);
nand UO_1655 (O_1655,N_29626,N_29988);
nand UO_1656 (O_1656,N_29766,N_29715);
xor UO_1657 (O_1657,N_29633,N_29818);
xnor UO_1658 (O_1658,N_29667,N_29759);
nand UO_1659 (O_1659,N_29550,N_29955);
and UO_1660 (O_1660,N_29688,N_29617);
and UO_1661 (O_1661,N_29773,N_29831);
xor UO_1662 (O_1662,N_29877,N_29702);
nor UO_1663 (O_1663,N_29845,N_29531);
or UO_1664 (O_1664,N_29892,N_29745);
or UO_1665 (O_1665,N_29540,N_29912);
xnor UO_1666 (O_1666,N_29980,N_29997);
xnor UO_1667 (O_1667,N_29896,N_29710);
nand UO_1668 (O_1668,N_29593,N_29790);
nand UO_1669 (O_1669,N_29683,N_29989);
and UO_1670 (O_1670,N_29824,N_29731);
nand UO_1671 (O_1671,N_29610,N_29981);
or UO_1672 (O_1672,N_29803,N_29547);
nor UO_1673 (O_1673,N_29694,N_29743);
nor UO_1674 (O_1674,N_29614,N_29948);
xor UO_1675 (O_1675,N_29581,N_29645);
xnor UO_1676 (O_1676,N_29964,N_29769);
nor UO_1677 (O_1677,N_29698,N_29523);
nand UO_1678 (O_1678,N_29958,N_29602);
or UO_1679 (O_1679,N_29560,N_29812);
or UO_1680 (O_1680,N_29720,N_29549);
or UO_1681 (O_1681,N_29689,N_29958);
nand UO_1682 (O_1682,N_29680,N_29695);
and UO_1683 (O_1683,N_29988,N_29519);
and UO_1684 (O_1684,N_29983,N_29525);
and UO_1685 (O_1685,N_29549,N_29780);
or UO_1686 (O_1686,N_29869,N_29867);
nand UO_1687 (O_1687,N_29862,N_29916);
nand UO_1688 (O_1688,N_29730,N_29760);
nor UO_1689 (O_1689,N_29931,N_29791);
nand UO_1690 (O_1690,N_29917,N_29505);
and UO_1691 (O_1691,N_29891,N_29675);
and UO_1692 (O_1692,N_29918,N_29938);
nor UO_1693 (O_1693,N_29810,N_29556);
nor UO_1694 (O_1694,N_29923,N_29931);
and UO_1695 (O_1695,N_29747,N_29560);
nand UO_1696 (O_1696,N_29843,N_29804);
or UO_1697 (O_1697,N_29599,N_29736);
or UO_1698 (O_1698,N_29951,N_29678);
xnor UO_1699 (O_1699,N_29535,N_29797);
and UO_1700 (O_1700,N_29586,N_29575);
xnor UO_1701 (O_1701,N_29521,N_29637);
and UO_1702 (O_1702,N_29737,N_29828);
nand UO_1703 (O_1703,N_29875,N_29937);
or UO_1704 (O_1704,N_29728,N_29917);
nor UO_1705 (O_1705,N_29616,N_29602);
and UO_1706 (O_1706,N_29647,N_29716);
nor UO_1707 (O_1707,N_29884,N_29704);
and UO_1708 (O_1708,N_29819,N_29855);
xor UO_1709 (O_1709,N_29806,N_29709);
xnor UO_1710 (O_1710,N_29759,N_29823);
or UO_1711 (O_1711,N_29894,N_29559);
xor UO_1712 (O_1712,N_29598,N_29850);
and UO_1713 (O_1713,N_29683,N_29640);
nor UO_1714 (O_1714,N_29503,N_29916);
and UO_1715 (O_1715,N_29515,N_29553);
nand UO_1716 (O_1716,N_29962,N_29539);
or UO_1717 (O_1717,N_29642,N_29745);
nand UO_1718 (O_1718,N_29535,N_29980);
or UO_1719 (O_1719,N_29881,N_29671);
nand UO_1720 (O_1720,N_29972,N_29617);
or UO_1721 (O_1721,N_29793,N_29733);
nor UO_1722 (O_1722,N_29892,N_29554);
and UO_1723 (O_1723,N_29996,N_29661);
xnor UO_1724 (O_1724,N_29793,N_29983);
xor UO_1725 (O_1725,N_29566,N_29794);
xor UO_1726 (O_1726,N_29765,N_29789);
nand UO_1727 (O_1727,N_29575,N_29595);
nand UO_1728 (O_1728,N_29566,N_29980);
xnor UO_1729 (O_1729,N_29659,N_29798);
or UO_1730 (O_1730,N_29832,N_29854);
or UO_1731 (O_1731,N_29724,N_29813);
nor UO_1732 (O_1732,N_29528,N_29508);
xnor UO_1733 (O_1733,N_29657,N_29877);
or UO_1734 (O_1734,N_29641,N_29984);
or UO_1735 (O_1735,N_29652,N_29807);
and UO_1736 (O_1736,N_29927,N_29969);
and UO_1737 (O_1737,N_29840,N_29537);
and UO_1738 (O_1738,N_29610,N_29673);
xnor UO_1739 (O_1739,N_29982,N_29508);
xor UO_1740 (O_1740,N_29501,N_29865);
nor UO_1741 (O_1741,N_29760,N_29592);
xnor UO_1742 (O_1742,N_29779,N_29876);
xor UO_1743 (O_1743,N_29528,N_29555);
and UO_1744 (O_1744,N_29729,N_29655);
or UO_1745 (O_1745,N_29556,N_29825);
and UO_1746 (O_1746,N_29522,N_29805);
nor UO_1747 (O_1747,N_29804,N_29514);
and UO_1748 (O_1748,N_29806,N_29710);
nand UO_1749 (O_1749,N_29848,N_29511);
xnor UO_1750 (O_1750,N_29862,N_29638);
or UO_1751 (O_1751,N_29542,N_29547);
or UO_1752 (O_1752,N_29568,N_29515);
and UO_1753 (O_1753,N_29614,N_29624);
nand UO_1754 (O_1754,N_29905,N_29752);
and UO_1755 (O_1755,N_29815,N_29576);
xor UO_1756 (O_1756,N_29870,N_29917);
xnor UO_1757 (O_1757,N_29945,N_29763);
nor UO_1758 (O_1758,N_29895,N_29935);
nor UO_1759 (O_1759,N_29994,N_29686);
or UO_1760 (O_1760,N_29761,N_29654);
or UO_1761 (O_1761,N_29841,N_29500);
or UO_1762 (O_1762,N_29582,N_29999);
and UO_1763 (O_1763,N_29531,N_29982);
or UO_1764 (O_1764,N_29877,N_29758);
or UO_1765 (O_1765,N_29553,N_29508);
or UO_1766 (O_1766,N_29858,N_29653);
nor UO_1767 (O_1767,N_29551,N_29714);
xnor UO_1768 (O_1768,N_29514,N_29925);
or UO_1769 (O_1769,N_29741,N_29573);
nand UO_1770 (O_1770,N_29688,N_29545);
or UO_1771 (O_1771,N_29611,N_29699);
or UO_1772 (O_1772,N_29611,N_29594);
and UO_1773 (O_1773,N_29984,N_29744);
nor UO_1774 (O_1774,N_29688,N_29813);
or UO_1775 (O_1775,N_29646,N_29500);
xnor UO_1776 (O_1776,N_29825,N_29963);
and UO_1777 (O_1777,N_29541,N_29547);
nand UO_1778 (O_1778,N_29768,N_29626);
or UO_1779 (O_1779,N_29687,N_29808);
xnor UO_1780 (O_1780,N_29919,N_29963);
nor UO_1781 (O_1781,N_29508,N_29664);
nand UO_1782 (O_1782,N_29832,N_29772);
and UO_1783 (O_1783,N_29571,N_29694);
or UO_1784 (O_1784,N_29773,N_29897);
nor UO_1785 (O_1785,N_29959,N_29619);
nor UO_1786 (O_1786,N_29670,N_29966);
nand UO_1787 (O_1787,N_29716,N_29673);
or UO_1788 (O_1788,N_29980,N_29955);
nor UO_1789 (O_1789,N_29758,N_29808);
or UO_1790 (O_1790,N_29929,N_29792);
and UO_1791 (O_1791,N_29659,N_29638);
nor UO_1792 (O_1792,N_29984,N_29858);
and UO_1793 (O_1793,N_29543,N_29794);
xnor UO_1794 (O_1794,N_29579,N_29667);
or UO_1795 (O_1795,N_29915,N_29994);
nor UO_1796 (O_1796,N_29632,N_29718);
nand UO_1797 (O_1797,N_29704,N_29702);
and UO_1798 (O_1798,N_29834,N_29723);
or UO_1799 (O_1799,N_29926,N_29749);
nand UO_1800 (O_1800,N_29726,N_29746);
and UO_1801 (O_1801,N_29866,N_29732);
or UO_1802 (O_1802,N_29562,N_29838);
and UO_1803 (O_1803,N_29532,N_29970);
nor UO_1804 (O_1804,N_29640,N_29820);
nand UO_1805 (O_1805,N_29921,N_29603);
and UO_1806 (O_1806,N_29817,N_29577);
xnor UO_1807 (O_1807,N_29884,N_29610);
nor UO_1808 (O_1808,N_29877,N_29606);
nand UO_1809 (O_1809,N_29560,N_29659);
nor UO_1810 (O_1810,N_29897,N_29747);
nand UO_1811 (O_1811,N_29765,N_29691);
xor UO_1812 (O_1812,N_29984,N_29813);
nor UO_1813 (O_1813,N_29678,N_29621);
nor UO_1814 (O_1814,N_29566,N_29903);
nand UO_1815 (O_1815,N_29602,N_29592);
xnor UO_1816 (O_1816,N_29512,N_29622);
nor UO_1817 (O_1817,N_29790,N_29743);
or UO_1818 (O_1818,N_29553,N_29853);
nor UO_1819 (O_1819,N_29815,N_29906);
and UO_1820 (O_1820,N_29954,N_29739);
nor UO_1821 (O_1821,N_29945,N_29778);
nand UO_1822 (O_1822,N_29665,N_29735);
or UO_1823 (O_1823,N_29700,N_29732);
and UO_1824 (O_1824,N_29709,N_29753);
nand UO_1825 (O_1825,N_29575,N_29652);
nor UO_1826 (O_1826,N_29775,N_29810);
nor UO_1827 (O_1827,N_29898,N_29746);
or UO_1828 (O_1828,N_29526,N_29664);
xor UO_1829 (O_1829,N_29858,N_29721);
or UO_1830 (O_1830,N_29889,N_29533);
nand UO_1831 (O_1831,N_29989,N_29701);
and UO_1832 (O_1832,N_29619,N_29504);
and UO_1833 (O_1833,N_29533,N_29541);
xor UO_1834 (O_1834,N_29973,N_29695);
xnor UO_1835 (O_1835,N_29789,N_29854);
nor UO_1836 (O_1836,N_29633,N_29749);
or UO_1837 (O_1837,N_29529,N_29580);
or UO_1838 (O_1838,N_29712,N_29848);
or UO_1839 (O_1839,N_29671,N_29751);
nand UO_1840 (O_1840,N_29708,N_29592);
xor UO_1841 (O_1841,N_29841,N_29981);
xnor UO_1842 (O_1842,N_29900,N_29922);
and UO_1843 (O_1843,N_29676,N_29558);
nand UO_1844 (O_1844,N_29517,N_29508);
or UO_1845 (O_1845,N_29845,N_29761);
or UO_1846 (O_1846,N_29588,N_29515);
and UO_1847 (O_1847,N_29523,N_29581);
xor UO_1848 (O_1848,N_29904,N_29806);
and UO_1849 (O_1849,N_29758,N_29666);
or UO_1850 (O_1850,N_29867,N_29817);
xnor UO_1851 (O_1851,N_29789,N_29882);
xnor UO_1852 (O_1852,N_29681,N_29605);
or UO_1853 (O_1853,N_29796,N_29831);
and UO_1854 (O_1854,N_29740,N_29889);
and UO_1855 (O_1855,N_29845,N_29548);
nor UO_1856 (O_1856,N_29993,N_29884);
and UO_1857 (O_1857,N_29842,N_29974);
and UO_1858 (O_1858,N_29610,N_29896);
and UO_1859 (O_1859,N_29642,N_29899);
or UO_1860 (O_1860,N_29556,N_29771);
or UO_1861 (O_1861,N_29696,N_29801);
or UO_1862 (O_1862,N_29847,N_29880);
and UO_1863 (O_1863,N_29596,N_29981);
or UO_1864 (O_1864,N_29655,N_29842);
or UO_1865 (O_1865,N_29879,N_29523);
and UO_1866 (O_1866,N_29737,N_29508);
or UO_1867 (O_1867,N_29952,N_29597);
or UO_1868 (O_1868,N_29638,N_29913);
xor UO_1869 (O_1869,N_29972,N_29708);
or UO_1870 (O_1870,N_29871,N_29757);
nor UO_1871 (O_1871,N_29713,N_29571);
and UO_1872 (O_1872,N_29886,N_29561);
xnor UO_1873 (O_1873,N_29821,N_29899);
nand UO_1874 (O_1874,N_29535,N_29955);
xor UO_1875 (O_1875,N_29897,N_29697);
xnor UO_1876 (O_1876,N_29922,N_29944);
nor UO_1877 (O_1877,N_29615,N_29922);
and UO_1878 (O_1878,N_29867,N_29772);
and UO_1879 (O_1879,N_29579,N_29836);
nor UO_1880 (O_1880,N_29621,N_29854);
nor UO_1881 (O_1881,N_29581,N_29658);
xor UO_1882 (O_1882,N_29691,N_29904);
and UO_1883 (O_1883,N_29974,N_29730);
nand UO_1884 (O_1884,N_29849,N_29553);
nand UO_1885 (O_1885,N_29784,N_29588);
nor UO_1886 (O_1886,N_29520,N_29518);
nor UO_1887 (O_1887,N_29775,N_29848);
xnor UO_1888 (O_1888,N_29928,N_29992);
nand UO_1889 (O_1889,N_29812,N_29555);
nor UO_1890 (O_1890,N_29801,N_29625);
nand UO_1891 (O_1891,N_29916,N_29580);
and UO_1892 (O_1892,N_29871,N_29819);
xnor UO_1893 (O_1893,N_29660,N_29817);
nand UO_1894 (O_1894,N_29608,N_29594);
and UO_1895 (O_1895,N_29996,N_29702);
nor UO_1896 (O_1896,N_29544,N_29619);
nand UO_1897 (O_1897,N_29680,N_29812);
nor UO_1898 (O_1898,N_29795,N_29774);
nor UO_1899 (O_1899,N_29753,N_29983);
nand UO_1900 (O_1900,N_29565,N_29778);
and UO_1901 (O_1901,N_29957,N_29637);
and UO_1902 (O_1902,N_29790,N_29504);
and UO_1903 (O_1903,N_29631,N_29694);
nand UO_1904 (O_1904,N_29725,N_29848);
xnor UO_1905 (O_1905,N_29694,N_29527);
nor UO_1906 (O_1906,N_29955,N_29748);
nand UO_1907 (O_1907,N_29847,N_29695);
and UO_1908 (O_1908,N_29500,N_29809);
nor UO_1909 (O_1909,N_29989,N_29660);
nand UO_1910 (O_1910,N_29587,N_29739);
nand UO_1911 (O_1911,N_29928,N_29966);
xnor UO_1912 (O_1912,N_29617,N_29942);
nor UO_1913 (O_1913,N_29548,N_29666);
and UO_1914 (O_1914,N_29803,N_29562);
nand UO_1915 (O_1915,N_29709,N_29841);
nor UO_1916 (O_1916,N_29918,N_29606);
nor UO_1917 (O_1917,N_29546,N_29850);
xnor UO_1918 (O_1918,N_29948,N_29530);
nor UO_1919 (O_1919,N_29711,N_29519);
nor UO_1920 (O_1920,N_29574,N_29867);
xor UO_1921 (O_1921,N_29968,N_29891);
xnor UO_1922 (O_1922,N_29746,N_29570);
or UO_1923 (O_1923,N_29637,N_29725);
and UO_1924 (O_1924,N_29717,N_29693);
or UO_1925 (O_1925,N_29838,N_29815);
nor UO_1926 (O_1926,N_29984,N_29712);
nor UO_1927 (O_1927,N_29703,N_29511);
nor UO_1928 (O_1928,N_29616,N_29514);
or UO_1929 (O_1929,N_29973,N_29877);
and UO_1930 (O_1930,N_29984,N_29620);
and UO_1931 (O_1931,N_29522,N_29665);
xor UO_1932 (O_1932,N_29952,N_29987);
nand UO_1933 (O_1933,N_29870,N_29591);
and UO_1934 (O_1934,N_29889,N_29511);
and UO_1935 (O_1935,N_29709,N_29963);
nand UO_1936 (O_1936,N_29797,N_29549);
or UO_1937 (O_1937,N_29935,N_29585);
nand UO_1938 (O_1938,N_29659,N_29756);
nand UO_1939 (O_1939,N_29502,N_29575);
and UO_1940 (O_1940,N_29766,N_29699);
and UO_1941 (O_1941,N_29551,N_29995);
nor UO_1942 (O_1942,N_29707,N_29695);
nor UO_1943 (O_1943,N_29954,N_29866);
or UO_1944 (O_1944,N_29840,N_29907);
and UO_1945 (O_1945,N_29954,N_29687);
nand UO_1946 (O_1946,N_29609,N_29599);
nand UO_1947 (O_1947,N_29936,N_29583);
and UO_1948 (O_1948,N_29744,N_29947);
nor UO_1949 (O_1949,N_29595,N_29849);
nand UO_1950 (O_1950,N_29695,N_29686);
and UO_1951 (O_1951,N_29749,N_29646);
and UO_1952 (O_1952,N_29613,N_29649);
or UO_1953 (O_1953,N_29745,N_29598);
xor UO_1954 (O_1954,N_29818,N_29530);
nor UO_1955 (O_1955,N_29718,N_29565);
xnor UO_1956 (O_1956,N_29533,N_29585);
nand UO_1957 (O_1957,N_29875,N_29609);
nor UO_1958 (O_1958,N_29950,N_29705);
nand UO_1959 (O_1959,N_29694,N_29518);
and UO_1960 (O_1960,N_29947,N_29747);
and UO_1961 (O_1961,N_29751,N_29588);
and UO_1962 (O_1962,N_29969,N_29964);
nor UO_1963 (O_1963,N_29910,N_29802);
and UO_1964 (O_1964,N_29687,N_29901);
or UO_1965 (O_1965,N_29832,N_29659);
nor UO_1966 (O_1966,N_29953,N_29547);
nor UO_1967 (O_1967,N_29978,N_29870);
nand UO_1968 (O_1968,N_29948,N_29536);
or UO_1969 (O_1969,N_29648,N_29839);
nor UO_1970 (O_1970,N_29947,N_29587);
or UO_1971 (O_1971,N_29993,N_29795);
nand UO_1972 (O_1972,N_29593,N_29850);
xor UO_1973 (O_1973,N_29526,N_29543);
nor UO_1974 (O_1974,N_29636,N_29721);
xor UO_1975 (O_1975,N_29685,N_29550);
and UO_1976 (O_1976,N_29616,N_29744);
nor UO_1977 (O_1977,N_29795,N_29706);
or UO_1978 (O_1978,N_29642,N_29891);
or UO_1979 (O_1979,N_29622,N_29680);
nor UO_1980 (O_1980,N_29512,N_29740);
or UO_1981 (O_1981,N_29826,N_29809);
or UO_1982 (O_1982,N_29540,N_29976);
and UO_1983 (O_1983,N_29887,N_29898);
nor UO_1984 (O_1984,N_29600,N_29797);
or UO_1985 (O_1985,N_29857,N_29751);
xor UO_1986 (O_1986,N_29753,N_29505);
nand UO_1987 (O_1987,N_29811,N_29759);
or UO_1988 (O_1988,N_29844,N_29595);
nor UO_1989 (O_1989,N_29667,N_29916);
xor UO_1990 (O_1990,N_29816,N_29537);
and UO_1991 (O_1991,N_29874,N_29966);
and UO_1992 (O_1992,N_29517,N_29770);
and UO_1993 (O_1993,N_29864,N_29952);
or UO_1994 (O_1994,N_29715,N_29542);
nand UO_1995 (O_1995,N_29962,N_29758);
or UO_1996 (O_1996,N_29760,N_29503);
xor UO_1997 (O_1997,N_29725,N_29549);
xnor UO_1998 (O_1998,N_29733,N_29664);
xnor UO_1999 (O_1999,N_29624,N_29868);
nand UO_2000 (O_2000,N_29758,N_29581);
or UO_2001 (O_2001,N_29851,N_29797);
xnor UO_2002 (O_2002,N_29946,N_29522);
or UO_2003 (O_2003,N_29791,N_29851);
or UO_2004 (O_2004,N_29823,N_29618);
nor UO_2005 (O_2005,N_29567,N_29902);
and UO_2006 (O_2006,N_29901,N_29821);
and UO_2007 (O_2007,N_29943,N_29717);
nand UO_2008 (O_2008,N_29814,N_29758);
and UO_2009 (O_2009,N_29929,N_29574);
xnor UO_2010 (O_2010,N_29661,N_29594);
or UO_2011 (O_2011,N_29836,N_29880);
nand UO_2012 (O_2012,N_29994,N_29510);
and UO_2013 (O_2013,N_29631,N_29714);
xor UO_2014 (O_2014,N_29814,N_29607);
xnor UO_2015 (O_2015,N_29892,N_29981);
nand UO_2016 (O_2016,N_29737,N_29929);
nor UO_2017 (O_2017,N_29552,N_29921);
nand UO_2018 (O_2018,N_29706,N_29842);
nor UO_2019 (O_2019,N_29875,N_29690);
xor UO_2020 (O_2020,N_29675,N_29593);
nor UO_2021 (O_2021,N_29593,N_29993);
nand UO_2022 (O_2022,N_29791,N_29637);
xor UO_2023 (O_2023,N_29634,N_29769);
nor UO_2024 (O_2024,N_29595,N_29989);
nand UO_2025 (O_2025,N_29737,N_29946);
and UO_2026 (O_2026,N_29656,N_29825);
xnor UO_2027 (O_2027,N_29617,N_29996);
or UO_2028 (O_2028,N_29767,N_29859);
or UO_2029 (O_2029,N_29806,N_29836);
and UO_2030 (O_2030,N_29539,N_29697);
and UO_2031 (O_2031,N_29655,N_29864);
or UO_2032 (O_2032,N_29509,N_29679);
or UO_2033 (O_2033,N_29808,N_29875);
xor UO_2034 (O_2034,N_29646,N_29681);
nand UO_2035 (O_2035,N_29721,N_29617);
nor UO_2036 (O_2036,N_29674,N_29858);
xnor UO_2037 (O_2037,N_29837,N_29594);
or UO_2038 (O_2038,N_29558,N_29628);
nand UO_2039 (O_2039,N_29649,N_29789);
xor UO_2040 (O_2040,N_29871,N_29728);
and UO_2041 (O_2041,N_29860,N_29934);
nand UO_2042 (O_2042,N_29733,N_29944);
and UO_2043 (O_2043,N_29869,N_29887);
and UO_2044 (O_2044,N_29689,N_29583);
or UO_2045 (O_2045,N_29622,N_29936);
xor UO_2046 (O_2046,N_29853,N_29504);
or UO_2047 (O_2047,N_29575,N_29625);
and UO_2048 (O_2048,N_29598,N_29812);
xor UO_2049 (O_2049,N_29542,N_29679);
and UO_2050 (O_2050,N_29578,N_29815);
nand UO_2051 (O_2051,N_29911,N_29834);
xnor UO_2052 (O_2052,N_29748,N_29510);
xor UO_2053 (O_2053,N_29815,N_29675);
nand UO_2054 (O_2054,N_29670,N_29982);
or UO_2055 (O_2055,N_29823,N_29943);
nor UO_2056 (O_2056,N_29873,N_29561);
nor UO_2057 (O_2057,N_29881,N_29771);
nor UO_2058 (O_2058,N_29959,N_29605);
xnor UO_2059 (O_2059,N_29879,N_29578);
nand UO_2060 (O_2060,N_29974,N_29834);
nand UO_2061 (O_2061,N_29571,N_29768);
nor UO_2062 (O_2062,N_29763,N_29719);
xor UO_2063 (O_2063,N_29635,N_29869);
and UO_2064 (O_2064,N_29860,N_29509);
nand UO_2065 (O_2065,N_29677,N_29690);
nand UO_2066 (O_2066,N_29583,N_29892);
nor UO_2067 (O_2067,N_29809,N_29537);
nand UO_2068 (O_2068,N_29501,N_29664);
nand UO_2069 (O_2069,N_29989,N_29916);
nand UO_2070 (O_2070,N_29835,N_29886);
nand UO_2071 (O_2071,N_29750,N_29588);
xor UO_2072 (O_2072,N_29543,N_29508);
or UO_2073 (O_2073,N_29548,N_29751);
and UO_2074 (O_2074,N_29605,N_29816);
nor UO_2075 (O_2075,N_29646,N_29610);
xor UO_2076 (O_2076,N_29762,N_29790);
or UO_2077 (O_2077,N_29956,N_29529);
and UO_2078 (O_2078,N_29901,N_29878);
xor UO_2079 (O_2079,N_29721,N_29841);
nor UO_2080 (O_2080,N_29948,N_29636);
and UO_2081 (O_2081,N_29870,N_29671);
or UO_2082 (O_2082,N_29806,N_29853);
nor UO_2083 (O_2083,N_29835,N_29663);
and UO_2084 (O_2084,N_29529,N_29818);
and UO_2085 (O_2085,N_29715,N_29682);
xor UO_2086 (O_2086,N_29726,N_29694);
xnor UO_2087 (O_2087,N_29685,N_29836);
or UO_2088 (O_2088,N_29948,N_29562);
or UO_2089 (O_2089,N_29605,N_29710);
and UO_2090 (O_2090,N_29849,N_29610);
and UO_2091 (O_2091,N_29705,N_29607);
and UO_2092 (O_2092,N_29605,N_29987);
xnor UO_2093 (O_2093,N_29540,N_29604);
nand UO_2094 (O_2094,N_29653,N_29756);
xor UO_2095 (O_2095,N_29954,N_29642);
xor UO_2096 (O_2096,N_29996,N_29887);
nand UO_2097 (O_2097,N_29705,N_29913);
nand UO_2098 (O_2098,N_29573,N_29982);
nor UO_2099 (O_2099,N_29582,N_29809);
xnor UO_2100 (O_2100,N_29717,N_29575);
nor UO_2101 (O_2101,N_29523,N_29768);
or UO_2102 (O_2102,N_29689,N_29898);
nor UO_2103 (O_2103,N_29711,N_29691);
or UO_2104 (O_2104,N_29505,N_29797);
and UO_2105 (O_2105,N_29674,N_29915);
and UO_2106 (O_2106,N_29591,N_29914);
nor UO_2107 (O_2107,N_29927,N_29724);
or UO_2108 (O_2108,N_29561,N_29894);
and UO_2109 (O_2109,N_29902,N_29972);
nor UO_2110 (O_2110,N_29926,N_29627);
nor UO_2111 (O_2111,N_29710,N_29854);
nor UO_2112 (O_2112,N_29730,N_29942);
nand UO_2113 (O_2113,N_29939,N_29756);
and UO_2114 (O_2114,N_29794,N_29883);
or UO_2115 (O_2115,N_29748,N_29706);
nor UO_2116 (O_2116,N_29637,N_29705);
nor UO_2117 (O_2117,N_29659,N_29584);
and UO_2118 (O_2118,N_29863,N_29974);
nand UO_2119 (O_2119,N_29912,N_29794);
xnor UO_2120 (O_2120,N_29511,N_29737);
and UO_2121 (O_2121,N_29571,N_29961);
xnor UO_2122 (O_2122,N_29514,N_29896);
nand UO_2123 (O_2123,N_29812,N_29911);
nand UO_2124 (O_2124,N_29778,N_29595);
or UO_2125 (O_2125,N_29775,N_29876);
or UO_2126 (O_2126,N_29514,N_29816);
or UO_2127 (O_2127,N_29680,N_29781);
nand UO_2128 (O_2128,N_29775,N_29817);
and UO_2129 (O_2129,N_29986,N_29700);
and UO_2130 (O_2130,N_29676,N_29783);
xnor UO_2131 (O_2131,N_29666,N_29914);
and UO_2132 (O_2132,N_29789,N_29539);
and UO_2133 (O_2133,N_29517,N_29795);
and UO_2134 (O_2134,N_29822,N_29782);
nand UO_2135 (O_2135,N_29501,N_29859);
xnor UO_2136 (O_2136,N_29689,N_29817);
nor UO_2137 (O_2137,N_29897,N_29862);
or UO_2138 (O_2138,N_29672,N_29606);
and UO_2139 (O_2139,N_29532,N_29774);
nor UO_2140 (O_2140,N_29661,N_29776);
nor UO_2141 (O_2141,N_29964,N_29814);
nand UO_2142 (O_2142,N_29865,N_29961);
nor UO_2143 (O_2143,N_29641,N_29826);
and UO_2144 (O_2144,N_29511,N_29808);
or UO_2145 (O_2145,N_29908,N_29856);
nand UO_2146 (O_2146,N_29540,N_29509);
nor UO_2147 (O_2147,N_29927,N_29835);
nor UO_2148 (O_2148,N_29503,N_29846);
nor UO_2149 (O_2149,N_29524,N_29924);
xnor UO_2150 (O_2150,N_29930,N_29926);
and UO_2151 (O_2151,N_29726,N_29892);
and UO_2152 (O_2152,N_29961,N_29669);
nor UO_2153 (O_2153,N_29628,N_29551);
and UO_2154 (O_2154,N_29779,N_29663);
nand UO_2155 (O_2155,N_29678,N_29521);
nand UO_2156 (O_2156,N_29584,N_29643);
nor UO_2157 (O_2157,N_29758,N_29507);
or UO_2158 (O_2158,N_29836,N_29588);
nand UO_2159 (O_2159,N_29999,N_29802);
xor UO_2160 (O_2160,N_29947,N_29641);
xor UO_2161 (O_2161,N_29668,N_29519);
xnor UO_2162 (O_2162,N_29624,N_29622);
or UO_2163 (O_2163,N_29928,N_29735);
nor UO_2164 (O_2164,N_29837,N_29693);
xor UO_2165 (O_2165,N_29834,N_29819);
or UO_2166 (O_2166,N_29790,N_29746);
or UO_2167 (O_2167,N_29568,N_29601);
and UO_2168 (O_2168,N_29852,N_29615);
xnor UO_2169 (O_2169,N_29883,N_29538);
and UO_2170 (O_2170,N_29822,N_29671);
and UO_2171 (O_2171,N_29536,N_29867);
nand UO_2172 (O_2172,N_29933,N_29557);
and UO_2173 (O_2173,N_29845,N_29565);
nand UO_2174 (O_2174,N_29993,N_29640);
nand UO_2175 (O_2175,N_29750,N_29791);
nor UO_2176 (O_2176,N_29591,N_29656);
and UO_2177 (O_2177,N_29796,N_29580);
nand UO_2178 (O_2178,N_29919,N_29678);
nor UO_2179 (O_2179,N_29785,N_29630);
xnor UO_2180 (O_2180,N_29636,N_29986);
or UO_2181 (O_2181,N_29759,N_29803);
nand UO_2182 (O_2182,N_29569,N_29515);
nand UO_2183 (O_2183,N_29977,N_29945);
xnor UO_2184 (O_2184,N_29980,N_29595);
nand UO_2185 (O_2185,N_29859,N_29634);
xor UO_2186 (O_2186,N_29849,N_29936);
nand UO_2187 (O_2187,N_29923,N_29983);
nand UO_2188 (O_2188,N_29522,N_29523);
and UO_2189 (O_2189,N_29540,N_29919);
nor UO_2190 (O_2190,N_29856,N_29719);
or UO_2191 (O_2191,N_29735,N_29985);
nor UO_2192 (O_2192,N_29956,N_29524);
or UO_2193 (O_2193,N_29592,N_29520);
xor UO_2194 (O_2194,N_29685,N_29914);
and UO_2195 (O_2195,N_29533,N_29995);
and UO_2196 (O_2196,N_29540,N_29517);
or UO_2197 (O_2197,N_29835,N_29538);
nand UO_2198 (O_2198,N_29774,N_29666);
nor UO_2199 (O_2199,N_29520,N_29958);
or UO_2200 (O_2200,N_29692,N_29957);
xnor UO_2201 (O_2201,N_29584,N_29744);
or UO_2202 (O_2202,N_29531,N_29657);
nor UO_2203 (O_2203,N_29739,N_29737);
nor UO_2204 (O_2204,N_29514,N_29868);
xor UO_2205 (O_2205,N_29806,N_29672);
xnor UO_2206 (O_2206,N_29965,N_29562);
nor UO_2207 (O_2207,N_29745,N_29877);
xnor UO_2208 (O_2208,N_29748,N_29765);
nand UO_2209 (O_2209,N_29624,N_29914);
or UO_2210 (O_2210,N_29696,N_29783);
and UO_2211 (O_2211,N_29945,N_29736);
and UO_2212 (O_2212,N_29547,N_29994);
nand UO_2213 (O_2213,N_29693,N_29901);
and UO_2214 (O_2214,N_29535,N_29851);
nor UO_2215 (O_2215,N_29608,N_29850);
or UO_2216 (O_2216,N_29698,N_29848);
and UO_2217 (O_2217,N_29622,N_29524);
and UO_2218 (O_2218,N_29648,N_29550);
nor UO_2219 (O_2219,N_29710,N_29909);
nand UO_2220 (O_2220,N_29906,N_29896);
nand UO_2221 (O_2221,N_29894,N_29837);
and UO_2222 (O_2222,N_29860,N_29879);
or UO_2223 (O_2223,N_29801,N_29597);
and UO_2224 (O_2224,N_29750,N_29902);
nor UO_2225 (O_2225,N_29551,N_29834);
xor UO_2226 (O_2226,N_29623,N_29890);
nor UO_2227 (O_2227,N_29927,N_29574);
and UO_2228 (O_2228,N_29810,N_29516);
nand UO_2229 (O_2229,N_29747,N_29506);
and UO_2230 (O_2230,N_29596,N_29989);
nand UO_2231 (O_2231,N_29737,N_29624);
and UO_2232 (O_2232,N_29505,N_29763);
nand UO_2233 (O_2233,N_29964,N_29945);
nor UO_2234 (O_2234,N_29775,N_29965);
or UO_2235 (O_2235,N_29595,N_29877);
and UO_2236 (O_2236,N_29527,N_29699);
or UO_2237 (O_2237,N_29579,N_29657);
or UO_2238 (O_2238,N_29705,N_29875);
nand UO_2239 (O_2239,N_29638,N_29631);
xor UO_2240 (O_2240,N_29511,N_29738);
and UO_2241 (O_2241,N_29762,N_29597);
xor UO_2242 (O_2242,N_29651,N_29753);
nand UO_2243 (O_2243,N_29840,N_29566);
and UO_2244 (O_2244,N_29540,N_29943);
xnor UO_2245 (O_2245,N_29515,N_29949);
nand UO_2246 (O_2246,N_29846,N_29917);
and UO_2247 (O_2247,N_29669,N_29742);
nand UO_2248 (O_2248,N_29578,N_29520);
and UO_2249 (O_2249,N_29933,N_29517);
nor UO_2250 (O_2250,N_29938,N_29716);
xor UO_2251 (O_2251,N_29953,N_29733);
nor UO_2252 (O_2252,N_29921,N_29869);
xor UO_2253 (O_2253,N_29672,N_29652);
or UO_2254 (O_2254,N_29793,N_29688);
xnor UO_2255 (O_2255,N_29572,N_29614);
and UO_2256 (O_2256,N_29839,N_29749);
nor UO_2257 (O_2257,N_29953,N_29976);
xnor UO_2258 (O_2258,N_29845,N_29559);
and UO_2259 (O_2259,N_29600,N_29745);
and UO_2260 (O_2260,N_29674,N_29574);
nand UO_2261 (O_2261,N_29827,N_29853);
xnor UO_2262 (O_2262,N_29635,N_29597);
or UO_2263 (O_2263,N_29809,N_29617);
nand UO_2264 (O_2264,N_29873,N_29815);
and UO_2265 (O_2265,N_29679,N_29647);
nor UO_2266 (O_2266,N_29531,N_29797);
nand UO_2267 (O_2267,N_29803,N_29700);
xor UO_2268 (O_2268,N_29875,N_29818);
nor UO_2269 (O_2269,N_29549,N_29561);
or UO_2270 (O_2270,N_29583,N_29802);
and UO_2271 (O_2271,N_29680,N_29519);
and UO_2272 (O_2272,N_29560,N_29842);
xor UO_2273 (O_2273,N_29501,N_29864);
xnor UO_2274 (O_2274,N_29932,N_29777);
nor UO_2275 (O_2275,N_29593,N_29686);
or UO_2276 (O_2276,N_29918,N_29501);
xnor UO_2277 (O_2277,N_29636,N_29609);
nor UO_2278 (O_2278,N_29907,N_29701);
nor UO_2279 (O_2279,N_29558,N_29909);
xor UO_2280 (O_2280,N_29970,N_29685);
and UO_2281 (O_2281,N_29505,N_29973);
nor UO_2282 (O_2282,N_29546,N_29555);
and UO_2283 (O_2283,N_29599,N_29929);
and UO_2284 (O_2284,N_29673,N_29650);
or UO_2285 (O_2285,N_29531,N_29952);
and UO_2286 (O_2286,N_29517,N_29677);
nor UO_2287 (O_2287,N_29564,N_29994);
or UO_2288 (O_2288,N_29996,N_29943);
and UO_2289 (O_2289,N_29514,N_29803);
nand UO_2290 (O_2290,N_29759,N_29842);
nor UO_2291 (O_2291,N_29906,N_29716);
or UO_2292 (O_2292,N_29533,N_29680);
and UO_2293 (O_2293,N_29929,N_29685);
nand UO_2294 (O_2294,N_29989,N_29956);
nor UO_2295 (O_2295,N_29993,N_29587);
nand UO_2296 (O_2296,N_29895,N_29616);
or UO_2297 (O_2297,N_29730,N_29831);
and UO_2298 (O_2298,N_29607,N_29748);
nand UO_2299 (O_2299,N_29784,N_29729);
and UO_2300 (O_2300,N_29805,N_29684);
nand UO_2301 (O_2301,N_29884,N_29823);
or UO_2302 (O_2302,N_29972,N_29532);
or UO_2303 (O_2303,N_29529,N_29504);
nand UO_2304 (O_2304,N_29638,N_29701);
nand UO_2305 (O_2305,N_29522,N_29514);
xor UO_2306 (O_2306,N_29968,N_29785);
and UO_2307 (O_2307,N_29913,N_29653);
or UO_2308 (O_2308,N_29916,N_29697);
nor UO_2309 (O_2309,N_29529,N_29671);
nand UO_2310 (O_2310,N_29628,N_29783);
nand UO_2311 (O_2311,N_29977,N_29888);
or UO_2312 (O_2312,N_29616,N_29527);
or UO_2313 (O_2313,N_29890,N_29884);
and UO_2314 (O_2314,N_29524,N_29858);
nor UO_2315 (O_2315,N_29986,N_29819);
xor UO_2316 (O_2316,N_29562,N_29693);
nor UO_2317 (O_2317,N_29986,N_29697);
xor UO_2318 (O_2318,N_29560,N_29535);
xor UO_2319 (O_2319,N_29747,N_29856);
nand UO_2320 (O_2320,N_29688,N_29808);
nor UO_2321 (O_2321,N_29601,N_29685);
nor UO_2322 (O_2322,N_29962,N_29762);
xnor UO_2323 (O_2323,N_29549,N_29719);
xnor UO_2324 (O_2324,N_29545,N_29787);
or UO_2325 (O_2325,N_29869,N_29724);
nand UO_2326 (O_2326,N_29501,N_29672);
and UO_2327 (O_2327,N_29797,N_29666);
nor UO_2328 (O_2328,N_29685,N_29916);
nor UO_2329 (O_2329,N_29664,N_29895);
xor UO_2330 (O_2330,N_29555,N_29817);
and UO_2331 (O_2331,N_29574,N_29871);
nand UO_2332 (O_2332,N_29909,N_29972);
nand UO_2333 (O_2333,N_29930,N_29998);
and UO_2334 (O_2334,N_29514,N_29768);
and UO_2335 (O_2335,N_29710,N_29936);
xnor UO_2336 (O_2336,N_29644,N_29506);
nor UO_2337 (O_2337,N_29803,N_29592);
xor UO_2338 (O_2338,N_29943,N_29662);
or UO_2339 (O_2339,N_29829,N_29986);
xor UO_2340 (O_2340,N_29649,N_29861);
or UO_2341 (O_2341,N_29865,N_29817);
xor UO_2342 (O_2342,N_29554,N_29875);
nor UO_2343 (O_2343,N_29726,N_29794);
xor UO_2344 (O_2344,N_29589,N_29795);
or UO_2345 (O_2345,N_29803,N_29634);
xor UO_2346 (O_2346,N_29706,N_29909);
xor UO_2347 (O_2347,N_29530,N_29709);
and UO_2348 (O_2348,N_29853,N_29963);
and UO_2349 (O_2349,N_29596,N_29647);
and UO_2350 (O_2350,N_29713,N_29763);
and UO_2351 (O_2351,N_29524,N_29512);
and UO_2352 (O_2352,N_29864,N_29867);
nand UO_2353 (O_2353,N_29703,N_29821);
nand UO_2354 (O_2354,N_29909,N_29634);
nand UO_2355 (O_2355,N_29922,N_29962);
xor UO_2356 (O_2356,N_29955,N_29809);
and UO_2357 (O_2357,N_29781,N_29636);
nand UO_2358 (O_2358,N_29518,N_29792);
nor UO_2359 (O_2359,N_29979,N_29760);
nor UO_2360 (O_2360,N_29794,N_29803);
xnor UO_2361 (O_2361,N_29905,N_29861);
nor UO_2362 (O_2362,N_29640,N_29803);
nand UO_2363 (O_2363,N_29662,N_29839);
xnor UO_2364 (O_2364,N_29951,N_29865);
or UO_2365 (O_2365,N_29814,N_29799);
nand UO_2366 (O_2366,N_29876,N_29837);
xnor UO_2367 (O_2367,N_29730,N_29858);
or UO_2368 (O_2368,N_29724,N_29876);
xor UO_2369 (O_2369,N_29912,N_29897);
nand UO_2370 (O_2370,N_29561,N_29950);
xnor UO_2371 (O_2371,N_29838,N_29515);
xnor UO_2372 (O_2372,N_29944,N_29948);
nor UO_2373 (O_2373,N_29507,N_29889);
and UO_2374 (O_2374,N_29687,N_29689);
nand UO_2375 (O_2375,N_29622,N_29995);
and UO_2376 (O_2376,N_29883,N_29889);
xnor UO_2377 (O_2377,N_29995,N_29891);
xnor UO_2378 (O_2378,N_29586,N_29559);
and UO_2379 (O_2379,N_29662,N_29753);
xnor UO_2380 (O_2380,N_29529,N_29904);
and UO_2381 (O_2381,N_29732,N_29994);
nor UO_2382 (O_2382,N_29550,N_29548);
xnor UO_2383 (O_2383,N_29564,N_29998);
and UO_2384 (O_2384,N_29674,N_29903);
nor UO_2385 (O_2385,N_29921,N_29835);
nor UO_2386 (O_2386,N_29540,N_29538);
and UO_2387 (O_2387,N_29979,N_29930);
nor UO_2388 (O_2388,N_29769,N_29963);
xnor UO_2389 (O_2389,N_29852,N_29944);
nor UO_2390 (O_2390,N_29637,N_29778);
nand UO_2391 (O_2391,N_29913,N_29656);
and UO_2392 (O_2392,N_29866,N_29642);
nor UO_2393 (O_2393,N_29757,N_29844);
and UO_2394 (O_2394,N_29883,N_29665);
nand UO_2395 (O_2395,N_29599,N_29712);
and UO_2396 (O_2396,N_29967,N_29782);
and UO_2397 (O_2397,N_29769,N_29797);
or UO_2398 (O_2398,N_29597,N_29832);
or UO_2399 (O_2399,N_29933,N_29916);
xnor UO_2400 (O_2400,N_29893,N_29555);
nor UO_2401 (O_2401,N_29674,N_29719);
xnor UO_2402 (O_2402,N_29730,N_29511);
or UO_2403 (O_2403,N_29636,N_29835);
and UO_2404 (O_2404,N_29768,N_29719);
and UO_2405 (O_2405,N_29896,N_29991);
and UO_2406 (O_2406,N_29623,N_29633);
nor UO_2407 (O_2407,N_29793,N_29920);
nor UO_2408 (O_2408,N_29511,N_29570);
nor UO_2409 (O_2409,N_29526,N_29924);
nor UO_2410 (O_2410,N_29932,N_29934);
or UO_2411 (O_2411,N_29664,N_29785);
or UO_2412 (O_2412,N_29614,N_29917);
nor UO_2413 (O_2413,N_29860,N_29989);
nand UO_2414 (O_2414,N_29513,N_29922);
xnor UO_2415 (O_2415,N_29606,N_29693);
and UO_2416 (O_2416,N_29669,N_29768);
and UO_2417 (O_2417,N_29931,N_29961);
and UO_2418 (O_2418,N_29689,N_29795);
xnor UO_2419 (O_2419,N_29701,N_29616);
or UO_2420 (O_2420,N_29719,N_29647);
and UO_2421 (O_2421,N_29851,N_29730);
nand UO_2422 (O_2422,N_29951,N_29800);
xnor UO_2423 (O_2423,N_29913,N_29832);
xor UO_2424 (O_2424,N_29580,N_29628);
nand UO_2425 (O_2425,N_29993,N_29513);
or UO_2426 (O_2426,N_29506,N_29978);
nor UO_2427 (O_2427,N_29876,N_29919);
xnor UO_2428 (O_2428,N_29871,N_29518);
nor UO_2429 (O_2429,N_29517,N_29777);
xnor UO_2430 (O_2430,N_29663,N_29970);
or UO_2431 (O_2431,N_29630,N_29958);
xor UO_2432 (O_2432,N_29953,N_29930);
and UO_2433 (O_2433,N_29870,N_29621);
xor UO_2434 (O_2434,N_29820,N_29873);
nor UO_2435 (O_2435,N_29531,N_29945);
or UO_2436 (O_2436,N_29981,N_29891);
nand UO_2437 (O_2437,N_29515,N_29780);
xnor UO_2438 (O_2438,N_29643,N_29997);
nor UO_2439 (O_2439,N_29909,N_29545);
nand UO_2440 (O_2440,N_29649,N_29637);
xor UO_2441 (O_2441,N_29880,N_29782);
and UO_2442 (O_2442,N_29633,N_29657);
xor UO_2443 (O_2443,N_29518,N_29509);
and UO_2444 (O_2444,N_29748,N_29611);
xor UO_2445 (O_2445,N_29846,N_29541);
nand UO_2446 (O_2446,N_29721,N_29904);
nor UO_2447 (O_2447,N_29978,N_29971);
xor UO_2448 (O_2448,N_29920,N_29515);
nand UO_2449 (O_2449,N_29697,N_29863);
or UO_2450 (O_2450,N_29979,N_29710);
or UO_2451 (O_2451,N_29812,N_29663);
xnor UO_2452 (O_2452,N_29555,N_29621);
nand UO_2453 (O_2453,N_29815,N_29741);
nor UO_2454 (O_2454,N_29977,N_29643);
and UO_2455 (O_2455,N_29506,N_29682);
xnor UO_2456 (O_2456,N_29607,N_29695);
xnor UO_2457 (O_2457,N_29790,N_29765);
nand UO_2458 (O_2458,N_29884,N_29651);
or UO_2459 (O_2459,N_29784,N_29576);
nand UO_2460 (O_2460,N_29654,N_29878);
or UO_2461 (O_2461,N_29744,N_29922);
and UO_2462 (O_2462,N_29995,N_29955);
nand UO_2463 (O_2463,N_29789,N_29547);
and UO_2464 (O_2464,N_29819,N_29612);
or UO_2465 (O_2465,N_29793,N_29933);
or UO_2466 (O_2466,N_29584,N_29801);
xor UO_2467 (O_2467,N_29883,N_29843);
nor UO_2468 (O_2468,N_29948,N_29557);
nor UO_2469 (O_2469,N_29710,N_29860);
nand UO_2470 (O_2470,N_29774,N_29967);
or UO_2471 (O_2471,N_29989,N_29725);
nand UO_2472 (O_2472,N_29824,N_29820);
and UO_2473 (O_2473,N_29509,N_29667);
xnor UO_2474 (O_2474,N_29790,N_29996);
nand UO_2475 (O_2475,N_29644,N_29745);
and UO_2476 (O_2476,N_29903,N_29539);
and UO_2477 (O_2477,N_29553,N_29624);
and UO_2478 (O_2478,N_29519,N_29887);
nand UO_2479 (O_2479,N_29543,N_29933);
nor UO_2480 (O_2480,N_29988,N_29619);
or UO_2481 (O_2481,N_29950,N_29778);
xnor UO_2482 (O_2482,N_29602,N_29773);
and UO_2483 (O_2483,N_29612,N_29914);
and UO_2484 (O_2484,N_29565,N_29562);
nand UO_2485 (O_2485,N_29848,N_29904);
or UO_2486 (O_2486,N_29816,N_29539);
or UO_2487 (O_2487,N_29955,N_29947);
or UO_2488 (O_2488,N_29872,N_29833);
or UO_2489 (O_2489,N_29645,N_29829);
or UO_2490 (O_2490,N_29627,N_29852);
or UO_2491 (O_2491,N_29824,N_29553);
nand UO_2492 (O_2492,N_29822,N_29705);
or UO_2493 (O_2493,N_29641,N_29975);
and UO_2494 (O_2494,N_29678,N_29606);
xor UO_2495 (O_2495,N_29517,N_29553);
and UO_2496 (O_2496,N_29708,N_29519);
xor UO_2497 (O_2497,N_29527,N_29951);
or UO_2498 (O_2498,N_29559,N_29769);
and UO_2499 (O_2499,N_29500,N_29664);
xor UO_2500 (O_2500,N_29800,N_29727);
xor UO_2501 (O_2501,N_29667,N_29552);
or UO_2502 (O_2502,N_29857,N_29599);
or UO_2503 (O_2503,N_29696,N_29966);
xor UO_2504 (O_2504,N_29904,N_29510);
or UO_2505 (O_2505,N_29887,N_29581);
and UO_2506 (O_2506,N_29595,N_29563);
and UO_2507 (O_2507,N_29850,N_29984);
and UO_2508 (O_2508,N_29861,N_29973);
and UO_2509 (O_2509,N_29854,N_29845);
and UO_2510 (O_2510,N_29698,N_29951);
or UO_2511 (O_2511,N_29648,N_29578);
nor UO_2512 (O_2512,N_29977,N_29842);
or UO_2513 (O_2513,N_29627,N_29919);
xor UO_2514 (O_2514,N_29970,N_29597);
nand UO_2515 (O_2515,N_29655,N_29848);
or UO_2516 (O_2516,N_29751,N_29655);
or UO_2517 (O_2517,N_29830,N_29671);
nand UO_2518 (O_2518,N_29607,N_29906);
and UO_2519 (O_2519,N_29832,N_29977);
or UO_2520 (O_2520,N_29583,N_29831);
xnor UO_2521 (O_2521,N_29925,N_29590);
nor UO_2522 (O_2522,N_29681,N_29808);
nand UO_2523 (O_2523,N_29965,N_29974);
and UO_2524 (O_2524,N_29676,N_29785);
nor UO_2525 (O_2525,N_29795,N_29695);
nand UO_2526 (O_2526,N_29842,N_29956);
nand UO_2527 (O_2527,N_29578,N_29631);
and UO_2528 (O_2528,N_29773,N_29605);
nand UO_2529 (O_2529,N_29897,N_29966);
or UO_2530 (O_2530,N_29770,N_29603);
or UO_2531 (O_2531,N_29521,N_29906);
and UO_2532 (O_2532,N_29942,N_29739);
xor UO_2533 (O_2533,N_29735,N_29518);
or UO_2534 (O_2534,N_29615,N_29926);
xnor UO_2535 (O_2535,N_29691,N_29893);
and UO_2536 (O_2536,N_29848,N_29987);
xnor UO_2537 (O_2537,N_29830,N_29500);
or UO_2538 (O_2538,N_29704,N_29826);
nand UO_2539 (O_2539,N_29891,N_29774);
and UO_2540 (O_2540,N_29518,N_29505);
and UO_2541 (O_2541,N_29741,N_29969);
xnor UO_2542 (O_2542,N_29519,N_29860);
nor UO_2543 (O_2543,N_29986,N_29803);
or UO_2544 (O_2544,N_29947,N_29637);
and UO_2545 (O_2545,N_29686,N_29823);
xnor UO_2546 (O_2546,N_29553,N_29876);
xor UO_2547 (O_2547,N_29784,N_29772);
nand UO_2548 (O_2548,N_29703,N_29761);
nand UO_2549 (O_2549,N_29703,N_29960);
or UO_2550 (O_2550,N_29976,N_29621);
nor UO_2551 (O_2551,N_29923,N_29686);
xnor UO_2552 (O_2552,N_29963,N_29921);
nand UO_2553 (O_2553,N_29975,N_29848);
nand UO_2554 (O_2554,N_29866,N_29882);
xor UO_2555 (O_2555,N_29698,N_29543);
or UO_2556 (O_2556,N_29637,N_29529);
nand UO_2557 (O_2557,N_29531,N_29766);
nor UO_2558 (O_2558,N_29782,N_29537);
or UO_2559 (O_2559,N_29975,N_29542);
xnor UO_2560 (O_2560,N_29679,N_29990);
nand UO_2561 (O_2561,N_29646,N_29981);
nand UO_2562 (O_2562,N_29999,N_29959);
xor UO_2563 (O_2563,N_29687,N_29957);
nand UO_2564 (O_2564,N_29615,N_29848);
or UO_2565 (O_2565,N_29925,N_29610);
nand UO_2566 (O_2566,N_29704,N_29554);
nand UO_2567 (O_2567,N_29505,N_29719);
nand UO_2568 (O_2568,N_29582,N_29629);
nor UO_2569 (O_2569,N_29519,N_29789);
nor UO_2570 (O_2570,N_29752,N_29935);
nor UO_2571 (O_2571,N_29918,N_29669);
xor UO_2572 (O_2572,N_29913,N_29657);
or UO_2573 (O_2573,N_29864,N_29933);
nor UO_2574 (O_2574,N_29841,N_29838);
nor UO_2575 (O_2575,N_29848,N_29880);
or UO_2576 (O_2576,N_29659,N_29698);
or UO_2577 (O_2577,N_29724,N_29972);
nand UO_2578 (O_2578,N_29999,N_29543);
xnor UO_2579 (O_2579,N_29976,N_29712);
xnor UO_2580 (O_2580,N_29754,N_29525);
and UO_2581 (O_2581,N_29792,N_29770);
nor UO_2582 (O_2582,N_29767,N_29564);
nor UO_2583 (O_2583,N_29540,N_29686);
xor UO_2584 (O_2584,N_29956,N_29875);
xor UO_2585 (O_2585,N_29699,N_29758);
nand UO_2586 (O_2586,N_29649,N_29528);
nor UO_2587 (O_2587,N_29996,N_29708);
nor UO_2588 (O_2588,N_29722,N_29625);
and UO_2589 (O_2589,N_29912,N_29662);
nand UO_2590 (O_2590,N_29709,N_29676);
nand UO_2591 (O_2591,N_29639,N_29748);
nand UO_2592 (O_2592,N_29810,N_29863);
nor UO_2593 (O_2593,N_29703,N_29914);
xor UO_2594 (O_2594,N_29909,N_29811);
xor UO_2595 (O_2595,N_29777,N_29572);
nand UO_2596 (O_2596,N_29711,N_29863);
and UO_2597 (O_2597,N_29583,N_29885);
or UO_2598 (O_2598,N_29971,N_29631);
or UO_2599 (O_2599,N_29962,N_29999);
nand UO_2600 (O_2600,N_29720,N_29901);
and UO_2601 (O_2601,N_29693,N_29949);
nand UO_2602 (O_2602,N_29850,N_29964);
nor UO_2603 (O_2603,N_29532,N_29716);
xnor UO_2604 (O_2604,N_29929,N_29818);
nand UO_2605 (O_2605,N_29952,N_29501);
nand UO_2606 (O_2606,N_29507,N_29618);
and UO_2607 (O_2607,N_29693,N_29841);
nand UO_2608 (O_2608,N_29942,N_29618);
or UO_2609 (O_2609,N_29557,N_29639);
and UO_2610 (O_2610,N_29832,N_29559);
or UO_2611 (O_2611,N_29919,N_29993);
xor UO_2612 (O_2612,N_29854,N_29616);
or UO_2613 (O_2613,N_29743,N_29782);
and UO_2614 (O_2614,N_29766,N_29737);
and UO_2615 (O_2615,N_29824,N_29881);
nand UO_2616 (O_2616,N_29506,N_29702);
or UO_2617 (O_2617,N_29614,N_29582);
nand UO_2618 (O_2618,N_29574,N_29580);
nand UO_2619 (O_2619,N_29938,N_29581);
and UO_2620 (O_2620,N_29788,N_29883);
nor UO_2621 (O_2621,N_29743,N_29745);
nand UO_2622 (O_2622,N_29684,N_29579);
xnor UO_2623 (O_2623,N_29839,N_29543);
or UO_2624 (O_2624,N_29510,N_29500);
xnor UO_2625 (O_2625,N_29884,N_29623);
nand UO_2626 (O_2626,N_29891,N_29776);
or UO_2627 (O_2627,N_29715,N_29570);
nand UO_2628 (O_2628,N_29609,N_29707);
and UO_2629 (O_2629,N_29631,N_29524);
xnor UO_2630 (O_2630,N_29935,N_29614);
and UO_2631 (O_2631,N_29835,N_29696);
nand UO_2632 (O_2632,N_29598,N_29844);
xnor UO_2633 (O_2633,N_29946,N_29765);
and UO_2634 (O_2634,N_29824,N_29520);
nand UO_2635 (O_2635,N_29596,N_29893);
nor UO_2636 (O_2636,N_29942,N_29789);
nand UO_2637 (O_2637,N_29698,N_29924);
and UO_2638 (O_2638,N_29773,N_29845);
or UO_2639 (O_2639,N_29995,N_29703);
nor UO_2640 (O_2640,N_29736,N_29567);
xor UO_2641 (O_2641,N_29913,N_29510);
and UO_2642 (O_2642,N_29555,N_29993);
nand UO_2643 (O_2643,N_29683,N_29998);
nand UO_2644 (O_2644,N_29724,N_29830);
nand UO_2645 (O_2645,N_29565,N_29945);
nor UO_2646 (O_2646,N_29519,N_29607);
or UO_2647 (O_2647,N_29844,N_29864);
or UO_2648 (O_2648,N_29699,N_29911);
or UO_2649 (O_2649,N_29543,N_29691);
nand UO_2650 (O_2650,N_29630,N_29611);
and UO_2651 (O_2651,N_29892,N_29524);
or UO_2652 (O_2652,N_29534,N_29759);
or UO_2653 (O_2653,N_29674,N_29979);
nand UO_2654 (O_2654,N_29672,N_29857);
or UO_2655 (O_2655,N_29697,N_29662);
xnor UO_2656 (O_2656,N_29817,N_29839);
xnor UO_2657 (O_2657,N_29953,N_29710);
or UO_2658 (O_2658,N_29611,N_29618);
nor UO_2659 (O_2659,N_29877,N_29520);
nand UO_2660 (O_2660,N_29869,N_29767);
and UO_2661 (O_2661,N_29715,N_29863);
or UO_2662 (O_2662,N_29592,N_29686);
xor UO_2663 (O_2663,N_29937,N_29893);
and UO_2664 (O_2664,N_29861,N_29995);
xnor UO_2665 (O_2665,N_29771,N_29610);
xnor UO_2666 (O_2666,N_29859,N_29969);
xnor UO_2667 (O_2667,N_29885,N_29717);
xor UO_2668 (O_2668,N_29828,N_29888);
and UO_2669 (O_2669,N_29678,N_29964);
or UO_2670 (O_2670,N_29659,N_29642);
xor UO_2671 (O_2671,N_29768,N_29628);
xnor UO_2672 (O_2672,N_29789,N_29627);
nand UO_2673 (O_2673,N_29545,N_29759);
or UO_2674 (O_2674,N_29573,N_29838);
or UO_2675 (O_2675,N_29642,N_29812);
or UO_2676 (O_2676,N_29674,N_29543);
xor UO_2677 (O_2677,N_29510,N_29940);
nor UO_2678 (O_2678,N_29901,N_29958);
and UO_2679 (O_2679,N_29677,N_29565);
or UO_2680 (O_2680,N_29676,N_29896);
or UO_2681 (O_2681,N_29956,N_29892);
or UO_2682 (O_2682,N_29600,N_29708);
nor UO_2683 (O_2683,N_29593,N_29748);
nor UO_2684 (O_2684,N_29971,N_29789);
nand UO_2685 (O_2685,N_29567,N_29846);
nor UO_2686 (O_2686,N_29665,N_29957);
nand UO_2687 (O_2687,N_29981,N_29884);
nor UO_2688 (O_2688,N_29763,N_29890);
nor UO_2689 (O_2689,N_29661,N_29824);
and UO_2690 (O_2690,N_29725,N_29926);
or UO_2691 (O_2691,N_29815,N_29948);
xor UO_2692 (O_2692,N_29888,N_29874);
or UO_2693 (O_2693,N_29665,N_29918);
nor UO_2694 (O_2694,N_29586,N_29626);
or UO_2695 (O_2695,N_29965,N_29923);
or UO_2696 (O_2696,N_29697,N_29909);
or UO_2697 (O_2697,N_29595,N_29678);
nand UO_2698 (O_2698,N_29517,N_29977);
xor UO_2699 (O_2699,N_29641,N_29905);
xnor UO_2700 (O_2700,N_29580,N_29870);
nor UO_2701 (O_2701,N_29542,N_29582);
nand UO_2702 (O_2702,N_29863,N_29709);
nand UO_2703 (O_2703,N_29873,N_29758);
or UO_2704 (O_2704,N_29542,N_29733);
and UO_2705 (O_2705,N_29600,N_29969);
nor UO_2706 (O_2706,N_29723,N_29735);
and UO_2707 (O_2707,N_29719,N_29968);
xor UO_2708 (O_2708,N_29922,N_29837);
nand UO_2709 (O_2709,N_29694,N_29900);
and UO_2710 (O_2710,N_29691,N_29698);
and UO_2711 (O_2711,N_29888,N_29565);
and UO_2712 (O_2712,N_29910,N_29767);
xnor UO_2713 (O_2713,N_29756,N_29769);
or UO_2714 (O_2714,N_29669,N_29973);
nand UO_2715 (O_2715,N_29565,N_29963);
or UO_2716 (O_2716,N_29950,N_29608);
xor UO_2717 (O_2717,N_29670,N_29919);
and UO_2718 (O_2718,N_29708,N_29765);
nand UO_2719 (O_2719,N_29769,N_29610);
xnor UO_2720 (O_2720,N_29954,N_29637);
xnor UO_2721 (O_2721,N_29868,N_29510);
nor UO_2722 (O_2722,N_29895,N_29693);
and UO_2723 (O_2723,N_29600,N_29519);
or UO_2724 (O_2724,N_29687,N_29609);
and UO_2725 (O_2725,N_29574,N_29560);
nor UO_2726 (O_2726,N_29621,N_29967);
nor UO_2727 (O_2727,N_29548,N_29527);
and UO_2728 (O_2728,N_29718,N_29521);
xnor UO_2729 (O_2729,N_29664,N_29769);
xnor UO_2730 (O_2730,N_29881,N_29694);
nor UO_2731 (O_2731,N_29880,N_29719);
and UO_2732 (O_2732,N_29741,N_29894);
nand UO_2733 (O_2733,N_29724,N_29857);
nor UO_2734 (O_2734,N_29901,N_29680);
xnor UO_2735 (O_2735,N_29690,N_29738);
xnor UO_2736 (O_2736,N_29730,N_29882);
xor UO_2737 (O_2737,N_29796,N_29721);
xor UO_2738 (O_2738,N_29742,N_29836);
nor UO_2739 (O_2739,N_29750,N_29929);
and UO_2740 (O_2740,N_29903,N_29728);
nand UO_2741 (O_2741,N_29649,N_29629);
or UO_2742 (O_2742,N_29904,N_29943);
or UO_2743 (O_2743,N_29616,N_29931);
nor UO_2744 (O_2744,N_29572,N_29697);
nand UO_2745 (O_2745,N_29792,N_29818);
or UO_2746 (O_2746,N_29868,N_29772);
nand UO_2747 (O_2747,N_29926,N_29800);
and UO_2748 (O_2748,N_29746,N_29682);
or UO_2749 (O_2749,N_29744,N_29680);
xnor UO_2750 (O_2750,N_29974,N_29544);
nor UO_2751 (O_2751,N_29527,N_29863);
nor UO_2752 (O_2752,N_29518,N_29620);
and UO_2753 (O_2753,N_29634,N_29843);
or UO_2754 (O_2754,N_29676,N_29957);
and UO_2755 (O_2755,N_29901,N_29791);
xnor UO_2756 (O_2756,N_29520,N_29972);
and UO_2757 (O_2757,N_29585,N_29863);
or UO_2758 (O_2758,N_29924,N_29855);
xnor UO_2759 (O_2759,N_29620,N_29797);
and UO_2760 (O_2760,N_29567,N_29854);
or UO_2761 (O_2761,N_29821,N_29898);
nand UO_2762 (O_2762,N_29615,N_29760);
and UO_2763 (O_2763,N_29688,N_29679);
or UO_2764 (O_2764,N_29516,N_29933);
xnor UO_2765 (O_2765,N_29638,N_29761);
xor UO_2766 (O_2766,N_29587,N_29823);
nand UO_2767 (O_2767,N_29766,N_29883);
xnor UO_2768 (O_2768,N_29844,N_29768);
or UO_2769 (O_2769,N_29591,N_29676);
nand UO_2770 (O_2770,N_29733,N_29921);
xnor UO_2771 (O_2771,N_29869,N_29611);
or UO_2772 (O_2772,N_29727,N_29963);
and UO_2773 (O_2773,N_29869,N_29693);
nor UO_2774 (O_2774,N_29715,N_29978);
xor UO_2775 (O_2775,N_29905,N_29675);
nor UO_2776 (O_2776,N_29824,N_29826);
or UO_2777 (O_2777,N_29559,N_29529);
nand UO_2778 (O_2778,N_29964,N_29642);
or UO_2779 (O_2779,N_29811,N_29961);
and UO_2780 (O_2780,N_29681,N_29584);
or UO_2781 (O_2781,N_29525,N_29538);
and UO_2782 (O_2782,N_29522,N_29648);
nand UO_2783 (O_2783,N_29644,N_29768);
and UO_2784 (O_2784,N_29796,N_29614);
xor UO_2785 (O_2785,N_29878,N_29634);
nand UO_2786 (O_2786,N_29941,N_29836);
xnor UO_2787 (O_2787,N_29569,N_29833);
xor UO_2788 (O_2788,N_29541,N_29536);
xnor UO_2789 (O_2789,N_29833,N_29790);
and UO_2790 (O_2790,N_29503,N_29926);
or UO_2791 (O_2791,N_29594,N_29898);
nor UO_2792 (O_2792,N_29934,N_29746);
xor UO_2793 (O_2793,N_29558,N_29720);
and UO_2794 (O_2794,N_29711,N_29646);
or UO_2795 (O_2795,N_29620,N_29527);
and UO_2796 (O_2796,N_29702,N_29969);
xor UO_2797 (O_2797,N_29859,N_29666);
and UO_2798 (O_2798,N_29531,N_29621);
or UO_2799 (O_2799,N_29959,N_29788);
xnor UO_2800 (O_2800,N_29863,N_29635);
and UO_2801 (O_2801,N_29764,N_29674);
or UO_2802 (O_2802,N_29960,N_29936);
or UO_2803 (O_2803,N_29803,N_29622);
xnor UO_2804 (O_2804,N_29805,N_29630);
or UO_2805 (O_2805,N_29845,N_29710);
nor UO_2806 (O_2806,N_29782,N_29841);
or UO_2807 (O_2807,N_29840,N_29794);
or UO_2808 (O_2808,N_29664,N_29780);
nand UO_2809 (O_2809,N_29879,N_29915);
nor UO_2810 (O_2810,N_29756,N_29958);
xor UO_2811 (O_2811,N_29668,N_29746);
or UO_2812 (O_2812,N_29970,N_29859);
nand UO_2813 (O_2813,N_29737,N_29675);
nand UO_2814 (O_2814,N_29983,N_29860);
and UO_2815 (O_2815,N_29768,N_29658);
and UO_2816 (O_2816,N_29560,N_29670);
and UO_2817 (O_2817,N_29695,N_29581);
or UO_2818 (O_2818,N_29628,N_29718);
or UO_2819 (O_2819,N_29983,N_29847);
nand UO_2820 (O_2820,N_29919,N_29565);
nor UO_2821 (O_2821,N_29508,N_29784);
and UO_2822 (O_2822,N_29833,N_29508);
and UO_2823 (O_2823,N_29513,N_29741);
or UO_2824 (O_2824,N_29564,N_29642);
xnor UO_2825 (O_2825,N_29545,N_29945);
nor UO_2826 (O_2826,N_29974,N_29503);
and UO_2827 (O_2827,N_29717,N_29680);
nand UO_2828 (O_2828,N_29857,N_29769);
or UO_2829 (O_2829,N_29649,N_29761);
xnor UO_2830 (O_2830,N_29894,N_29822);
nor UO_2831 (O_2831,N_29976,N_29928);
xnor UO_2832 (O_2832,N_29760,N_29995);
nand UO_2833 (O_2833,N_29886,N_29907);
xnor UO_2834 (O_2834,N_29960,N_29768);
nor UO_2835 (O_2835,N_29693,N_29667);
xor UO_2836 (O_2836,N_29626,N_29648);
and UO_2837 (O_2837,N_29726,N_29689);
nand UO_2838 (O_2838,N_29904,N_29554);
xor UO_2839 (O_2839,N_29888,N_29991);
or UO_2840 (O_2840,N_29837,N_29773);
nor UO_2841 (O_2841,N_29640,N_29501);
xnor UO_2842 (O_2842,N_29798,N_29609);
nand UO_2843 (O_2843,N_29549,N_29784);
nor UO_2844 (O_2844,N_29920,N_29608);
and UO_2845 (O_2845,N_29711,N_29884);
and UO_2846 (O_2846,N_29804,N_29529);
or UO_2847 (O_2847,N_29635,N_29533);
nor UO_2848 (O_2848,N_29892,N_29952);
nor UO_2849 (O_2849,N_29825,N_29644);
nand UO_2850 (O_2850,N_29813,N_29932);
xor UO_2851 (O_2851,N_29870,N_29937);
and UO_2852 (O_2852,N_29894,N_29928);
nand UO_2853 (O_2853,N_29900,N_29690);
nor UO_2854 (O_2854,N_29565,N_29500);
or UO_2855 (O_2855,N_29557,N_29553);
nand UO_2856 (O_2856,N_29873,N_29807);
and UO_2857 (O_2857,N_29657,N_29619);
or UO_2858 (O_2858,N_29772,N_29577);
xnor UO_2859 (O_2859,N_29923,N_29589);
nor UO_2860 (O_2860,N_29957,N_29699);
nand UO_2861 (O_2861,N_29933,N_29724);
and UO_2862 (O_2862,N_29737,N_29582);
and UO_2863 (O_2863,N_29838,N_29618);
nor UO_2864 (O_2864,N_29917,N_29760);
nor UO_2865 (O_2865,N_29989,N_29563);
nor UO_2866 (O_2866,N_29805,N_29701);
and UO_2867 (O_2867,N_29978,N_29939);
or UO_2868 (O_2868,N_29975,N_29684);
and UO_2869 (O_2869,N_29713,N_29703);
and UO_2870 (O_2870,N_29913,N_29933);
and UO_2871 (O_2871,N_29720,N_29749);
or UO_2872 (O_2872,N_29592,N_29999);
or UO_2873 (O_2873,N_29993,N_29779);
nand UO_2874 (O_2874,N_29522,N_29557);
and UO_2875 (O_2875,N_29502,N_29883);
and UO_2876 (O_2876,N_29994,N_29905);
or UO_2877 (O_2877,N_29888,N_29954);
and UO_2878 (O_2878,N_29716,N_29757);
and UO_2879 (O_2879,N_29740,N_29578);
nand UO_2880 (O_2880,N_29734,N_29861);
and UO_2881 (O_2881,N_29905,N_29626);
nor UO_2882 (O_2882,N_29891,N_29673);
and UO_2883 (O_2883,N_29893,N_29569);
or UO_2884 (O_2884,N_29526,N_29698);
nor UO_2885 (O_2885,N_29833,N_29931);
xor UO_2886 (O_2886,N_29813,N_29660);
nor UO_2887 (O_2887,N_29777,N_29864);
xnor UO_2888 (O_2888,N_29911,N_29632);
or UO_2889 (O_2889,N_29590,N_29879);
nor UO_2890 (O_2890,N_29905,N_29904);
and UO_2891 (O_2891,N_29868,N_29822);
nor UO_2892 (O_2892,N_29765,N_29994);
or UO_2893 (O_2893,N_29879,N_29584);
and UO_2894 (O_2894,N_29747,N_29687);
nand UO_2895 (O_2895,N_29946,N_29861);
nand UO_2896 (O_2896,N_29547,N_29992);
nor UO_2897 (O_2897,N_29684,N_29502);
nor UO_2898 (O_2898,N_29800,N_29628);
nor UO_2899 (O_2899,N_29700,N_29514);
and UO_2900 (O_2900,N_29898,N_29739);
and UO_2901 (O_2901,N_29681,N_29649);
nor UO_2902 (O_2902,N_29755,N_29547);
nor UO_2903 (O_2903,N_29695,N_29659);
nand UO_2904 (O_2904,N_29921,N_29936);
nand UO_2905 (O_2905,N_29924,N_29943);
and UO_2906 (O_2906,N_29880,N_29605);
and UO_2907 (O_2907,N_29553,N_29905);
nor UO_2908 (O_2908,N_29702,N_29765);
and UO_2909 (O_2909,N_29904,N_29507);
xnor UO_2910 (O_2910,N_29750,N_29637);
and UO_2911 (O_2911,N_29785,N_29717);
nor UO_2912 (O_2912,N_29698,N_29841);
and UO_2913 (O_2913,N_29582,N_29734);
or UO_2914 (O_2914,N_29606,N_29670);
nor UO_2915 (O_2915,N_29724,N_29619);
or UO_2916 (O_2916,N_29580,N_29969);
nand UO_2917 (O_2917,N_29960,N_29744);
and UO_2918 (O_2918,N_29894,N_29752);
and UO_2919 (O_2919,N_29573,N_29748);
xnor UO_2920 (O_2920,N_29811,N_29931);
xor UO_2921 (O_2921,N_29901,N_29970);
and UO_2922 (O_2922,N_29898,N_29872);
xor UO_2923 (O_2923,N_29534,N_29648);
or UO_2924 (O_2924,N_29786,N_29958);
nor UO_2925 (O_2925,N_29727,N_29784);
and UO_2926 (O_2926,N_29754,N_29534);
or UO_2927 (O_2927,N_29890,N_29918);
xnor UO_2928 (O_2928,N_29737,N_29897);
xnor UO_2929 (O_2929,N_29741,N_29798);
nor UO_2930 (O_2930,N_29555,N_29626);
and UO_2931 (O_2931,N_29547,N_29792);
xor UO_2932 (O_2932,N_29910,N_29934);
or UO_2933 (O_2933,N_29566,N_29750);
or UO_2934 (O_2934,N_29714,N_29683);
nor UO_2935 (O_2935,N_29954,N_29744);
xor UO_2936 (O_2936,N_29920,N_29886);
or UO_2937 (O_2937,N_29870,N_29982);
and UO_2938 (O_2938,N_29821,N_29829);
nand UO_2939 (O_2939,N_29642,N_29922);
xnor UO_2940 (O_2940,N_29533,N_29829);
nor UO_2941 (O_2941,N_29732,N_29947);
nor UO_2942 (O_2942,N_29975,N_29956);
nor UO_2943 (O_2943,N_29529,N_29599);
nand UO_2944 (O_2944,N_29686,N_29947);
nor UO_2945 (O_2945,N_29560,N_29511);
or UO_2946 (O_2946,N_29739,N_29909);
nor UO_2947 (O_2947,N_29760,N_29685);
and UO_2948 (O_2948,N_29633,N_29548);
nor UO_2949 (O_2949,N_29748,N_29731);
or UO_2950 (O_2950,N_29931,N_29905);
and UO_2951 (O_2951,N_29701,N_29579);
and UO_2952 (O_2952,N_29907,N_29585);
and UO_2953 (O_2953,N_29806,N_29777);
or UO_2954 (O_2954,N_29802,N_29990);
and UO_2955 (O_2955,N_29876,N_29688);
or UO_2956 (O_2956,N_29661,N_29669);
and UO_2957 (O_2957,N_29544,N_29683);
nor UO_2958 (O_2958,N_29725,N_29923);
xnor UO_2959 (O_2959,N_29669,N_29949);
or UO_2960 (O_2960,N_29597,N_29618);
nand UO_2961 (O_2961,N_29703,N_29855);
xnor UO_2962 (O_2962,N_29830,N_29624);
nand UO_2963 (O_2963,N_29854,N_29812);
nor UO_2964 (O_2964,N_29668,N_29612);
nand UO_2965 (O_2965,N_29752,N_29969);
or UO_2966 (O_2966,N_29904,N_29545);
or UO_2967 (O_2967,N_29581,N_29724);
nand UO_2968 (O_2968,N_29532,N_29677);
or UO_2969 (O_2969,N_29501,N_29746);
or UO_2970 (O_2970,N_29790,N_29987);
and UO_2971 (O_2971,N_29600,N_29842);
nor UO_2972 (O_2972,N_29719,N_29831);
nand UO_2973 (O_2973,N_29986,N_29809);
or UO_2974 (O_2974,N_29899,N_29686);
nand UO_2975 (O_2975,N_29515,N_29940);
nor UO_2976 (O_2976,N_29504,N_29940);
nand UO_2977 (O_2977,N_29945,N_29829);
or UO_2978 (O_2978,N_29606,N_29617);
xnor UO_2979 (O_2979,N_29650,N_29776);
nand UO_2980 (O_2980,N_29605,N_29512);
xor UO_2981 (O_2981,N_29978,N_29533);
nand UO_2982 (O_2982,N_29592,N_29512);
and UO_2983 (O_2983,N_29890,N_29719);
nor UO_2984 (O_2984,N_29643,N_29798);
or UO_2985 (O_2985,N_29577,N_29820);
xor UO_2986 (O_2986,N_29797,N_29838);
and UO_2987 (O_2987,N_29594,N_29586);
and UO_2988 (O_2988,N_29646,N_29573);
or UO_2989 (O_2989,N_29502,N_29941);
nand UO_2990 (O_2990,N_29612,N_29779);
and UO_2991 (O_2991,N_29822,N_29878);
xnor UO_2992 (O_2992,N_29792,N_29717);
nor UO_2993 (O_2993,N_29620,N_29541);
nor UO_2994 (O_2994,N_29969,N_29972);
or UO_2995 (O_2995,N_29589,N_29960);
and UO_2996 (O_2996,N_29621,N_29659);
nand UO_2997 (O_2997,N_29915,N_29849);
or UO_2998 (O_2998,N_29637,N_29732);
nand UO_2999 (O_2999,N_29638,N_29852);
or UO_3000 (O_3000,N_29737,N_29542);
nor UO_3001 (O_3001,N_29787,N_29753);
and UO_3002 (O_3002,N_29765,N_29639);
nand UO_3003 (O_3003,N_29631,N_29716);
nand UO_3004 (O_3004,N_29989,N_29751);
nor UO_3005 (O_3005,N_29578,N_29632);
nand UO_3006 (O_3006,N_29963,N_29581);
and UO_3007 (O_3007,N_29641,N_29775);
or UO_3008 (O_3008,N_29560,N_29579);
nand UO_3009 (O_3009,N_29879,N_29782);
nor UO_3010 (O_3010,N_29777,N_29845);
xor UO_3011 (O_3011,N_29994,N_29659);
nor UO_3012 (O_3012,N_29709,N_29535);
xor UO_3013 (O_3013,N_29744,N_29737);
xnor UO_3014 (O_3014,N_29664,N_29805);
xnor UO_3015 (O_3015,N_29739,N_29670);
nor UO_3016 (O_3016,N_29855,N_29541);
or UO_3017 (O_3017,N_29742,N_29821);
and UO_3018 (O_3018,N_29867,N_29534);
nor UO_3019 (O_3019,N_29721,N_29566);
xor UO_3020 (O_3020,N_29697,N_29514);
nand UO_3021 (O_3021,N_29661,N_29591);
xnor UO_3022 (O_3022,N_29930,N_29997);
or UO_3023 (O_3023,N_29571,N_29700);
and UO_3024 (O_3024,N_29855,N_29977);
nor UO_3025 (O_3025,N_29912,N_29645);
nor UO_3026 (O_3026,N_29795,N_29662);
or UO_3027 (O_3027,N_29884,N_29941);
and UO_3028 (O_3028,N_29539,N_29728);
xnor UO_3029 (O_3029,N_29769,N_29614);
nor UO_3030 (O_3030,N_29910,N_29870);
nand UO_3031 (O_3031,N_29820,N_29891);
nor UO_3032 (O_3032,N_29590,N_29839);
nand UO_3033 (O_3033,N_29675,N_29906);
and UO_3034 (O_3034,N_29752,N_29557);
xnor UO_3035 (O_3035,N_29905,N_29610);
nand UO_3036 (O_3036,N_29840,N_29898);
nand UO_3037 (O_3037,N_29692,N_29914);
xor UO_3038 (O_3038,N_29751,N_29901);
and UO_3039 (O_3039,N_29916,N_29894);
xnor UO_3040 (O_3040,N_29925,N_29723);
or UO_3041 (O_3041,N_29761,N_29928);
or UO_3042 (O_3042,N_29505,N_29768);
nand UO_3043 (O_3043,N_29978,N_29646);
xor UO_3044 (O_3044,N_29521,N_29566);
nand UO_3045 (O_3045,N_29555,N_29735);
nand UO_3046 (O_3046,N_29774,N_29552);
and UO_3047 (O_3047,N_29948,N_29912);
nor UO_3048 (O_3048,N_29951,N_29989);
nand UO_3049 (O_3049,N_29680,N_29662);
or UO_3050 (O_3050,N_29783,N_29564);
nand UO_3051 (O_3051,N_29948,N_29852);
and UO_3052 (O_3052,N_29748,N_29644);
or UO_3053 (O_3053,N_29613,N_29969);
xor UO_3054 (O_3054,N_29621,N_29685);
or UO_3055 (O_3055,N_29747,N_29757);
and UO_3056 (O_3056,N_29774,N_29946);
xnor UO_3057 (O_3057,N_29920,N_29679);
nand UO_3058 (O_3058,N_29633,N_29876);
nand UO_3059 (O_3059,N_29665,N_29803);
nor UO_3060 (O_3060,N_29666,N_29645);
and UO_3061 (O_3061,N_29931,N_29584);
and UO_3062 (O_3062,N_29977,N_29950);
and UO_3063 (O_3063,N_29710,N_29917);
or UO_3064 (O_3064,N_29811,N_29844);
or UO_3065 (O_3065,N_29956,N_29803);
xnor UO_3066 (O_3066,N_29975,N_29989);
nand UO_3067 (O_3067,N_29976,N_29680);
xor UO_3068 (O_3068,N_29678,N_29793);
and UO_3069 (O_3069,N_29929,N_29881);
xor UO_3070 (O_3070,N_29784,N_29973);
xor UO_3071 (O_3071,N_29756,N_29657);
or UO_3072 (O_3072,N_29762,N_29705);
nor UO_3073 (O_3073,N_29812,N_29913);
and UO_3074 (O_3074,N_29557,N_29644);
or UO_3075 (O_3075,N_29602,N_29835);
nand UO_3076 (O_3076,N_29858,N_29558);
and UO_3077 (O_3077,N_29660,N_29857);
xnor UO_3078 (O_3078,N_29625,N_29810);
or UO_3079 (O_3079,N_29688,N_29718);
and UO_3080 (O_3080,N_29777,N_29663);
nand UO_3081 (O_3081,N_29928,N_29910);
or UO_3082 (O_3082,N_29510,N_29512);
and UO_3083 (O_3083,N_29648,N_29553);
and UO_3084 (O_3084,N_29825,N_29796);
and UO_3085 (O_3085,N_29568,N_29925);
nand UO_3086 (O_3086,N_29983,N_29518);
nand UO_3087 (O_3087,N_29538,N_29861);
and UO_3088 (O_3088,N_29522,N_29543);
nor UO_3089 (O_3089,N_29567,N_29907);
or UO_3090 (O_3090,N_29589,N_29717);
xnor UO_3091 (O_3091,N_29534,N_29822);
nor UO_3092 (O_3092,N_29845,N_29970);
and UO_3093 (O_3093,N_29883,N_29936);
and UO_3094 (O_3094,N_29502,N_29999);
xor UO_3095 (O_3095,N_29725,N_29955);
nand UO_3096 (O_3096,N_29865,N_29984);
nand UO_3097 (O_3097,N_29792,N_29786);
and UO_3098 (O_3098,N_29707,N_29921);
xnor UO_3099 (O_3099,N_29675,N_29789);
nand UO_3100 (O_3100,N_29999,N_29971);
nand UO_3101 (O_3101,N_29604,N_29539);
nand UO_3102 (O_3102,N_29662,N_29564);
nand UO_3103 (O_3103,N_29779,N_29679);
nand UO_3104 (O_3104,N_29506,N_29636);
nand UO_3105 (O_3105,N_29605,N_29529);
or UO_3106 (O_3106,N_29847,N_29859);
or UO_3107 (O_3107,N_29744,N_29516);
nor UO_3108 (O_3108,N_29695,N_29611);
xor UO_3109 (O_3109,N_29608,N_29900);
nand UO_3110 (O_3110,N_29889,N_29990);
or UO_3111 (O_3111,N_29968,N_29904);
xor UO_3112 (O_3112,N_29517,N_29808);
and UO_3113 (O_3113,N_29628,N_29578);
or UO_3114 (O_3114,N_29850,N_29615);
and UO_3115 (O_3115,N_29799,N_29764);
nor UO_3116 (O_3116,N_29758,N_29846);
or UO_3117 (O_3117,N_29796,N_29654);
nor UO_3118 (O_3118,N_29929,N_29640);
or UO_3119 (O_3119,N_29708,N_29813);
and UO_3120 (O_3120,N_29782,N_29785);
nand UO_3121 (O_3121,N_29618,N_29577);
nor UO_3122 (O_3122,N_29530,N_29795);
xor UO_3123 (O_3123,N_29542,N_29786);
nand UO_3124 (O_3124,N_29512,N_29799);
nand UO_3125 (O_3125,N_29795,N_29800);
and UO_3126 (O_3126,N_29744,N_29842);
nor UO_3127 (O_3127,N_29753,N_29708);
nor UO_3128 (O_3128,N_29915,N_29606);
or UO_3129 (O_3129,N_29592,N_29633);
nand UO_3130 (O_3130,N_29802,N_29826);
and UO_3131 (O_3131,N_29977,N_29598);
and UO_3132 (O_3132,N_29570,N_29824);
or UO_3133 (O_3133,N_29930,N_29772);
and UO_3134 (O_3134,N_29730,N_29500);
xor UO_3135 (O_3135,N_29676,N_29669);
nand UO_3136 (O_3136,N_29838,N_29532);
xor UO_3137 (O_3137,N_29672,N_29908);
nand UO_3138 (O_3138,N_29699,N_29633);
xor UO_3139 (O_3139,N_29507,N_29601);
and UO_3140 (O_3140,N_29651,N_29678);
nand UO_3141 (O_3141,N_29542,N_29573);
nand UO_3142 (O_3142,N_29814,N_29896);
xnor UO_3143 (O_3143,N_29934,N_29904);
nand UO_3144 (O_3144,N_29806,N_29912);
nand UO_3145 (O_3145,N_29808,N_29932);
xor UO_3146 (O_3146,N_29603,N_29772);
and UO_3147 (O_3147,N_29538,N_29886);
nand UO_3148 (O_3148,N_29849,N_29902);
nand UO_3149 (O_3149,N_29567,N_29665);
nor UO_3150 (O_3150,N_29722,N_29860);
or UO_3151 (O_3151,N_29567,N_29642);
or UO_3152 (O_3152,N_29831,N_29577);
or UO_3153 (O_3153,N_29784,N_29716);
nand UO_3154 (O_3154,N_29784,N_29756);
xnor UO_3155 (O_3155,N_29956,N_29840);
or UO_3156 (O_3156,N_29612,N_29673);
or UO_3157 (O_3157,N_29558,N_29821);
nor UO_3158 (O_3158,N_29997,N_29619);
xnor UO_3159 (O_3159,N_29885,N_29568);
xor UO_3160 (O_3160,N_29886,N_29577);
nor UO_3161 (O_3161,N_29500,N_29680);
or UO_3162 (O_3162,N_29746,N_29760);
nand UO_3163 (O_3163,N_29531,N_29540);
nor UO_3164 (O_3164,N_29845,N_29823);
or UO_3165 (O_3165,N_29686,N_29565);
nand UO_3166 (O_3166,N_29722,N_29659);
nand UO_3167 (O_3167,N_29592,N_29634);
or UO_3168 (O_3168,N_29803,N_29855);
xnor UO_3169 (O_3169,N_29969,N_29512);
nor UO_3170 (O_3170,N_29770,N_29966);
xnor UO_3171 (O_3171,N_29562,N_29787);
nand UO_3172 (O_3172,N_29843,N_29933);
nand UO_3173 (O_3173,N_29907,N_29848);
or UO_3174 (O_3174,N_29967,N_29626);
and UO_3175 (O_3175,N_29564,N_29966);
xor UO_3176 (O_3176,N_29593,N_29886);
or UO_3177 (O_3177,N_29794,N_29538);
and UO_3178 (O_3178,N_29614,N_29800);
or UO_3179 (O_3179,N_29579,N_29883);
xor UO_3180 (O_3180,N_29844,N_29898);
xor UO_3181 (O_3181,N_29763,N_29655);
nand UO_3182 (O_3182,N_29742,N_29771);
nand UO_3183 (O_3183,N_29907,N_29690);
and UO_3184 (O_3184,N_29604,N_29645);
xor UO_3185 (O_3185,N_29735,N_29653);
or UO_3186 (O_3186,N_29944,N_29943);
and UO_3187 (O_3187,N_29972,N_29772);
or UO_3188 (O_3188,N_29999,N_29970);
xnor UO_3189 (O_3189,N_29512,N_29553);
and UO_3190 (O_3190,N_29760,N_29811);
nor UO_3191 (O_3191,N_29796,N_29644);
or UO_3192 (O_3192,N_29640,N_29907);
nor UO_3193 (O_3193,N_29703,N_29845);
and UO_3194 (O_3194,N_29581,N_29609);
nor UO_3195 (O_3195,N_29765,N_29931);
xnor UO_3196 (O_3196,N_29633,N_29718);
xnor UO_3197 (O_3197,N_29838,N_29678);
and UO_3198 (O_3198,N_29590,N_29862);
xnor UO_3199 (O_3199,N_29703,N_29735);
and UO_3200 (O_3200,N_29940,N_29740);
nand UO_3201 (O_3201,N_29643,N_29575);
or UO_3202 (O_3202,N_29814,N_29849);
nand UO_3203 (O_3203,N_29609,N_29652);
nand UO_3204 (O_3204,N_29615,N_29692);
nor UO_3205 (O_3205,N_29545,N_29636);
nand UO_3206 (O_3206,N_29827,N_29854);
xnor UO_3207 (O_3207,N_29526,N_29669);
nand UO_3208 (O_3208,N_29563,N_29583);
nor UO_3209 (O_3209,N_29919,N_29852);
nor UO_3210 (O_3210,N_29693,N_29722);
or UO_3211 (O_3211,N_29811,N_29791);
and UO_3212 (O_3212,N_29583,N_29544);
and UO_3213 (O_3213,N_29764,N_29543);
xnor UO_3214 (O_3214,N_29863,N_29818);
xnor UO_3215 (O_3215,N_29652,N_29798);
xor UO_3216 (O_3216,N_29647,N_29805);
nor UO_3217 (O_3217,N_29858,N_29750);
nand UO_3218 (O_3218,N_29609,N_29655);
xor UO_3219 (O_3219,N_29851,N_29821);
or UO_3220 (O_3220,N_29876,N_29550);
nand UO_3221 (O_3221,N_29652,N_29642);
or UO_3222 (O_3222,N_29733,N_29876);
xor UO_3223 (O_3223,N_29706,N_29629);
nand UO_3224 (O_3224,N_29621,N_29629);
nor UO_3225 (O_3225,N_29716,N_29738);
nand UO_3226 (O_3226,N_29951,N_29685);
and UO_3227 (O_3227,N_29759,N_29754);
xor UO_3228 (O_3228,N_29537,N_29629);
xor UO_3229 (O_3229,N_29560,N_29729);
and UO_3230 (O_3230,N_29946,N_29827);
or UO_3231 (O_3231,N_29547,N_29754);
or UO_3232 (O_3232,N_29715,N_29756);
nand UO_3233 (O_3233,N_29533,N_29590);
nand UO_3234 (O_3234,N_29754,N_29780);
nand UO_3235 (O_3235,N_29754,N_29969);
and UO_3236 (O_3236,N_29647,N_29793);
xor UO_3237 (O_3237,N_29685,N_29997);
and UO_3238 (O_3238,N_29520,N_29995);
nand UO_3239 (O_3239,N_29973,N_29763);
or UO_3240 (O_3240,N_29590,N_29987);
or UO_3241 (O_3241,N_29634,N_29943);
and UO_3242 (O_3242,N_29611,N_29741);
or UO_3243 (O_3243,N_29617,N_29600);
or UO_3244 (O_3244,N_29799,N_29876);
xnor UO_3245 (O_3245,N_29672,N_29555);
or UO_3246 (O_3246,N_29725,N_29877);
nor UO_3247 (O_3247,N_29888,N_29969);
xnor UO_3248 (O_3248,N_29501,N_29748);
or UO_3249 (O_3249,N_29624,N_29506);
xnor UO_3250 (O_3250,N_29541,N_29573);
xnor UO_3251 (O_3251,N_29836,N_29677);
xnor UO_3252 (O_3252,N_29516,N_29726);
or UO_3253 (O_3253,N_29832,N_29815);
xnor UO_3254 (O_3254,N_29506,N_29893);
nand UO_3255 (O_3255,N_29825,N_29827);
nor UO_3256 (O_3256,N_29674,N_29623);
and UO_3257 (O_3257,N_29740,N_29862);
nor UO_3258 (O_3258,N_29679,N_29557);
nor UO_3259 (O_3259,N_29729,N_29559);
or UO_3260 (O_3260,N_29860,N_29861);
or UO_3261 (O_3261,N_29776,N_29546);
nor UO_3262 (O_3262,N_29750,N_29695);
or UO_3263 (O_3263,N_29862,N_29951);
nand UO_3264 (O_3264,N_29613,N_29872);
or UO_3265 (O_3265,N_29719,N_29993);
xnor UO_3266 (O_3266,N_29670,N_29687);
or UO_3267 (O_3267,N_29584,N_29740);
nand UO_3268 (O_3268,N_29716,N_29545);
nor UO_3269 (O_3269,N_29582,N_29939);
or UO_3270 (O_3270,N_29589,N_29811);
and UO_3271 (O_3271,N_29978,N_29861);
nor UO_3272 (O_3272,N_29867,N_29807);
and UO_3273 (O_3273,N_29782,N_29679);
nand UO_3274 (O_3274,N_29656,N_29808);
nand UO_3275 (O_3275,N_29859,N_29675);
or UO_3276 (O_3276,N_29859,N_29822);
xnor UO_3277 (O_3277,N_29836,N_29839);
xor UO_3278 (O_3278,N_29819,N_29898);
and UO_3279 (O_3279,N_29885,N_29574);
nor UO_3280 (O_3280,N_29798,N_29815);
nor UO_3281 (O_3281,N_29827,N_29893);
nand UO_3282 (O_3282,N_29707,N_29944);
xor UO_3283 (O_3283,N_29870,N_29558);
and UO_3284 (O_3284,N_29692,N_29913);
or UO_3285 (O_3285,N_29702,N_29922);
or UO_3286 (O_3286,N_29926,N_29995);
or UO_3287 (O_3287,N_29939,N_29924);
xnor UO_3288 (O_3288,N_29601,N_29569);
nor UO_3289 (O_3289,N_29930,N_29887);
nor UO_3290 (O_3290,N_29815,N_29568);
nand UO_3291 (O_3291,N_29675,N_29505);
or UO_3292 (O_3292,N_29748,N_29826);
or UO_3293 (O_3293,N_29900,N_29500);
nand UO_3294 (O_3294,N_29628,N_29791);
or UO_3295 (O_3295,N_29843,N_29568);
or UO_3296 (O_3296,N_29574,N_29875);
nand UO_3297 (O_3297,N_29813,N_29525);
and UO_3298 (O_3298,N_29953,N_29509);
xnor UO_3299 (O_3299,N_29728,N_29885);
nand UO_3300 (O_3300,N_29523,N_29890);
nand UO_3301 (O_3301,N_29770,N_29771);
and UO_3302 (O_3302,N_29963,N_29549);
and UO_3303 (O_3303,N_29504,N_29924);
xor UO_3304 (O_3304,N_29648,N_29738);
nand UO_3305 (O_3305,N_29654,N_29528);
nand UO_3306 (O_3306,N_29802,N_29655);
or UO_3307 (O_3307,N_29845,N_29659);
nor UO_3308 (O_3308,N_29657,N_29713);
and UO_3309 (O_3309,N_29784,N_29935);
nand UO_3310 (O_3310,N_29661,N_29667);
nor UO_3311 (O_3311,N_29905,N_29753);
xnor UO_3312 (O_3312,N_29864,N_29631);
and UO_3313 (O_3313,N_29924,N_29680);
or UO_3314 (O_3314,N_29693,N_29736);
or UO_3315 (O_3315,N_29613,N_29918);
and UO_3316 (O_3316,N_29668,N_29503);
and UO_3317 (O_3317,N_29715,N_29855);
and UO_3318 (O_3318,N_29967,N_29554);
nor UO_3319 (O_3319,N_29557,N_29587);
nand UO_3320 (O_3320,N_29674,N_29893);
nand UO_3321 (O_3321,N_29655,N_29504);
nand UO_3322 (O_3322,N_29876,N_29545);
and UO_3323 (O_3323,N_29521,N_29782);
and UO_3324 (O_3324,N_29880,N_29623);
and UO_3325 (O_3325,N_29779,N_29865);
xor UO_3326 (O_3326,N_29866,N_29643);
nor UO_3327 (O_3327,N_29936,N_29536);
and UO_3328 (O_3328,N_29923,N_29732);
nand UO_3329 (O_3329,N_29849,N_29624);
nor UO_3330 (O_3330,N_29736,N_29562);
nor UO_3331 (O_3331,N_29749,N_29981);
nand UO_3332 (O_3332,N_29577,N_29592);
xnor UO_3333 (O_3333,N_29961,N_29920);
nor UO_3334 (O_3334,N_29612,N_29799);
nand UO_3335 (O_3335,N_29741,N_29593);
nand UO_3336 (O_3336,N_29533,N_29911);
nand UO_3337 (O_3337,N_29828,N_29790);
nor UO_3338 (O_3338,N_29691,N_29810);
and UO_3339 (O_3339,N_29680,N_29883);
nand UO_3340 (O_3340,N_29873,N_29591);
nor UO_3341 (O_3341,N_29874,N_29541);
nand UO_3342 (O_3342,N_29533,N_29900);
or UO_3343 (O_3343,N_29801,N_29715);
nand UO_3344 (O_3344,N_29899,N_29961);
nor UO_3345 (O_3345,N_29991,N_29940);
or UO_3346 (O_3346,N_29867,N_29835);
or UO_3347 (O_3347,N_29872,N_29735);
xor UO_3348 (O_3348,N_29932,N_29712);
xnor UO_3349 (O_3349,N_29874,N_29617);
or UO_3350 (O_3350,N_29523,N_29656);
and UO_3351 (O_3351,N_29820,N_29505);
nand UO_3352 (O_3352,N_29743,N_29817);
or UO_3353 (O_3353,N_29619,N_29650);
nand UO_3354 (O_3354,N_29517,N_29713);
or UO_3355 (O_3355,N_29588,N_29758);
or UO_3356 (O_3356,N_29979,N_29864);
and UO_3357 (O_3357,N_29972,N_29521);
and UO_3358 (O_3358,N_29952,N_29781);
and UO_3359 (O_3359,N_29621,N_29961);
and UO_3360 (O_3360,N_29811,N_29651);
and UO_3361 (O_3361,N_29664,N_29668);
nand UO_3362 (O_3362,N_29708,N_29723);
nand UO_3363 (O_3363,N_29857,N_29902);
nor UO_3364 (O_3364,N_29679,N_29729);
xnor UO_3365 (O_3365,N_29747,N_29733);
and UO_3366 (O_3366,N_29785,N_29928);
xnor UO_3367 (O_3367,N_29552,N_29743);
xnor UO_3368 (O_3368,N_29871,N_29741);
or UO_3369 (O_3369,N_29575,N_29532);
nand UO_3370 (O_3370,N_29964,N_29711);
or UO_3371 (O_3371,N_29966,N_29832);
or UO_3372 (O_3372,N_29679,N_29845);
nor UO_3373 (O_3373,N_29659,N_29928);
and UO_3374 (O_3374,N_29855,N_29740);
nand UO_3375 (O_3375,N_29508,N_29822);
nand UO_3376 (O_3376,N_29539,N_29995);
or UO_3377 (O_3377,N_29510,N_29971);
or UO_3378 (O_3378,N_29612,N_29705);
nor UO_3379 (O_3379,N_29771,N_29704);
nand UO_3380 (O_3380,N_29860,N_29757);
or UO_3381 (O_3381,N_29557,N_29783);
nor UO_3382 (O_3382,N_29766,N_29753);
xnor UO_3383 (O_3383,N_29851,N_29777);
nand UO_3384 (O_3384,N_29991,N_29988);
xor UO_3385 (O_3385,N_29513,N_29874);
nor UO_3386 (O_3386,N_29726,N_29874);
nand UO_3387 (O_3387,N_29662,N_29521);
and UO_3388 (O_3388,N_29590,N_29830);
nand UO_3389 (O_3389,N_29877,N_29803);
and UO_3390 (O_3390,N_29995,N_29987);
or UO_3391 (O_3391,N_29949,N_29789);
and UO_3392 (O_3392,N_29669,N_29647);
xnor UO_3393 (O_3393,N_29970,N_29631);
nand UO_3394 (O_3394,N_29895,N_29801);
and UO_3395 (O_3395,N_29582,N_29548);
and UO_3396 (O_3396,N_29580,N_29512);
xor UO_3397 (O_3397,N_29911,N_29945);
xnor UO_3398 (O_3398,N_29634,N_29625);
nor UO_3399 (O_3399,N_29758,N_29896);
nand UO_3400 (O_3400,N_29831,N_29726);
and UO_3401 (O_3401,N_29773,N_29891);
and UO_3402 (O_3402,N_29976,N_29800);
nand UO_3403 (O_3403,N_29519,N_29572);
nor UO_3404 (O_3404,N_29931,N_29541);
xor UO_3405 (O_3405,N_29874,N_29867);
or UO_3406 (O_3406,N_29733,N_29753);
or UO_3407 (O_3407,N_29639,N_29978);
or UO_3408 (O_3408,N_29502,N_29709);
or UO_3409 (O_3409,N_29964,N_29873);
nand UO_3410 (O_3410,N_29774,N_29947);
nand UO_3411 (O_3411,N_29871,N_29774);
nand UO_3412 (O_3412,N_29771,N_29725);
and UO_3413 (O_3413,N_29967,N_29736);
and UO_3414 (O_3414,N_29697,N_29728);
xnor UO_3415 (O_3415,N_29528,N_29530);
and UO_3416 (O_3416,N_29943,N_29686);
and UO_3417 (O_3417,N_29514,N_29790);
nor UO_3418 (O_3418,N_29536,N_29754);
nand UO_3419 (O_3419,N_29732,N_29725);
and UO_3420 (O_3420,N_29653,N_29727);
and UO_3421 (O_3421,N_29932,N_29698);
nand UO_3422 (O_3422,N_29917,N_29575);
xnor UO_3423 (O_3423,N_29979,N_29530);
or UO_3424 (O_3424,N_29906,N_29596);
and UO_3425 (O_3425,N_29570,N_29527);
nor UO_3426 (O_3426,N_29655,N_29639);
nand UO_3427 (O_3427,N_29828,N_29867);
and UO_3428 (O_3428,N_29633,N_29808);
xnor UO_3429 (O_3429,N_29614,N_29777);
nand UO_3430 (O_3430,N_29717,N_29722);
or UO_3431 (O_3431,N_29879,N_29651);
or UO_3432 (O_3432,N_29720,N_29961);
nand UO_3433 (O_3433,N_29964,N_29596);
nand UO_3434 (O_3434,N_29763,N_29884);
xor UO_3435 (O_3435,N_29577,N_29671);
or UO_3436 (O_3436,N_29976,N_29692);
and UO_3437 (O_3437,N_29597,N_29619);
nand UO_3438 (O_3438,N_29669,N_29734);
nand UO_3439 (O_3439,N_29969,N_29866);
or UO_3440 (O_3440,N_29805,N_29966);
or UO_3441 (O_3441,N_29824,N_29633);
or UO_3442 (O_3442,N_29610,N_29526);
nor UO_3443 (O_3443,N_29953,N_29937);
nor UO_3444 (O_3444,N_29765,N_29851);
nor UO_3445 (O_3445,N_29919,N_29693);
xnor UO_3446 (O_3446,N_29719,N_29635);
nand UO_3447 (O_3447,N_29766,N_29824);
nor UO_3448 (O_3448,N_29628,N_29567);
xor UO_3449 (O_3449,N_29732,N_29681);
nand UO_3450 (O_3450,N_29812,N_29879);
or UO_3451 (O_3451,N_29827,N_29614);
xnor UO_3452 (O_3452,N_29569,N_29603);
nand UO_3453 (O_3453,N_29657,N_29936);
nor UO_3454 (O_3454,N_29726,N_29925);
or UO_3455 (O_3455,N_29940,N_29816);
nand UO_3456 (O_3456,N_29791,N_29521);
nand UO_3457 (O_3457,N_29796,N_29860);
xnor UO_3458 (O_3458,N_29769,N_29570);
xnor UO_3459 (O_3459,N_29922,N_29994);
xnor UO_3460 (O_3460,N_29678,N_29557);
nor UO_3461 (O_3461,N_29635,N_29825);
or UO_3462 (O_3462,N_29934,N_29959);
nor UO_3463 (O_3463,N_29819,N_29893);
and UO_3464 (O_3464,N_29749,N_29825);
or UO_3465 (O_3465,N_29678,N_29815);
and UO_3466 (O_3466,N_29577,N_29546);
nand UO_3467 (O_3467,N_29983,N_29543);
and UO_3468 (O_3468,N_29814,N_29663);
nor UO_3469 (O_3469,N_29830,N_29980);
nor UO_3470 (O_3470,N_29586,N_29849);
nor UO_3471 (O_3471,N_29785,N_29979);
xor UO_3472 (O_3472,N_29987,N_29969);
or UO_3473 (O_3473,N_29602,N_29525);
nand UO_3474 (O_3474,N_29760,N_29821);
nor UO_3475 (O_3475,N_29962,N_29538);
nor UO_3476 (O_3476,N_29709,N_29810);
nand UO_3477 (O_3477,N_29523,N_29627);
and UO_3478 (O_3478,N_29916,N_29824);
or UO_3479 (O_3479,N_29662,N_29986);
nor UO_3480 (O_3480,N_29566,N_29856);
nor UO_3481 (O_3481,N_29746,N_29930);
or UO_3482 (O_3482,N_29999,N_29775);
and UO_3483 (O_3483,N_29888,N_29629);
nor UO_3484 (O_3484,N_29828,N_29994);
or UO_3485 (O_3485,N_29783,N_29754);
xnor UO_3486 (O_3486,N_29689,N_29823);
nor UO_3487 (O_3487,N_29527,N_29631);
and UO_3488 (O_3488,N_29953,N_29741);
or UO_3489 (O_3489,N_29851,N_29878);
nor UO_3490 (O_3490,N_29704,N_29808);
and UO_3491 (O_3491,N_29614,N_29876);
xor UO_3492 (O_3492,N_29672,N_29630);
nor UO_3493 (O_3493,N_29967,N_29622);
or UO_3494 (O_3494,N_29803,N_29785);
or UO_3495 (O_3495,N_29509,N_29740);
or UO_3496 (O_3496,N_29912,N_29604);
nor UO_3497 (O_3497,N_29892,N_29829);
or UO_3498 (O_3498,N_29556,N_29674);
nor UO_3499 (O_3499,N_29557,N_29860);
endmodule