module basic_5000_50000_5000_200_levels_10xor_9(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,In_3000,In_3001,In_3002,In_3003,In_3004,In_3005,In_3006,In_3007,In_3008,In_3009,In_3010,In_3011,In_3012,In_3013,In_3014,In_3015,In_3016,In_3017,In_3018,In_3019,In_3020,In_3021,In_3022,In_3023,In_3024,In_3025,In_3026,In_3027,In_3028,In_3029,In_3030,In_3031,In_3032,In_3033,In_3034,In_3035,In_3036,In_3037,In_3038,In_3039,In_3040,In_3041,In_3042,In_3043,In_3044,In_3045,In_3046,In_3047,In_3048,In_3049,In_3050,In_3051,In_3052,In_3053,In_3054,In_3055,In_3056,In_3057,In_3058,In_3059,In_3060,In_3061,In_3062,In_3063,In_3064,In_3065,In_3066,In_3067,In_3068,In_3069,In_3070,In_3071,In_3072,In_3073,In_3074,In_3075,In_3076,In_3077,In_3078,In_3079,In_3080,In_3081,In_3082,In_3083,In_3084,In_3085,In_3086,In_3087,In_3088,In_3089,In_3090,In_3091,In_3092,In_3093,In_3094,In_3095,In_3096,In_3097,In_3098,In_3099,In_3100,In_3101,In_3102,In_3103,In_3104,In_3105,In_3106,In_3107,In_3108,In_3109,In_3110,In_3111,In_3112,In_3113,In_3114,In_3115,In_3116,In_3117,In_3118,In_3119,In_3120,In_3121,In_3122,In_3123,In_3124,In_3125,In_3126,In_3127,In_3128,In_3129,In_3130,In_3131,In_3132,In_3133,In_3134,In_3135,In_3136,In_3137,In_3138,In_3139,In_3140,In_3141,In_3142,In_3143,In_3144,In_3145,In_3146,In_3147,In_3148,In_3149,In_3150,In_3151,In_3152,In_3153,In_3154,In_3155,In_3156,In_3157,In_3158,In_3159,In_3160,In_3161,In_3162,In_3163,In_3164,In_3165,In_3166,In_3167,In_3168,In_3169,In_3170,In_3171,In_3172,In_3173,In_3174,In_3175,In_3176,In_3177,In_3178,In_3179,In_3180,In_3181,In_3182,In_3183,In_3184,In_3185,In_3186,In_3187,In_3188,In_3189,In_3190,In_3191,In_3192,In_3193,In_3194,In_3195,In_3196,In_3197,In_3198,In_3199,In_3200,In_3201,In_3202,In_3203,In_3204,In_3205,In_3206,In_3207,In_3208,In_3209,In_3210,In_3211,In_3212,In_3213,In_3214,In_3215,In_3216,In_3217,In_3218,In_3219,In_3220,In_3221,In_3222,In_3223,In_3224,In_3225,In_3226,In_3227,In_3228,In_3229,In_3230,In_3231,In_3232,In_3233,In_3234,In_3235,In_3236,In_3237,In_3238,In_3239,In_3240,In_3241,In_3242,In_3243,In_3244,In_3245,In_3246,In_3247,In_3248,In_3249,In_3250,In_3251,In_3252,In_3253,In_3254,In_3255,In_3256,In_3257,In_3258,In_3259,In_3260,In_3261,In_3262,In_3263,In_3264,In_3265,In_3266,In_3267,In_3268,In_3269,In_3270,In_3271,In_3272,In_3273,In_3274,In_3275,In_3276,In_3277,In_3278,In_3279,In_3280,In_3281,In_3282,In_3283,In_3284,In_3285,In_3286,In_3287,In_3288,In_3289,In_3290,In_3291,In_3292,In_3293,In_3294,In_3295,In_3296,In_3297,In_3298,In_3299,In_3300,In_3301,In_3302,In_3303,In_3304,In_3305,In_3306,In_3307,In_3308,In_3309,In_3310,In_3311,In_3312,In_3313,In_3314,In_3315,In_3316,In_3317,In_3318,In_3319,In_3320,In_3321,In_3322,In_3323,In_3324,In_3325,In_3326,In_3327,In_3328,In_3329,In_3330,In_3331,In_3332,In_3333,In_3334,In_3335,In_3336,In_3337,In_3338,In_3339,In_3340,In_3341,In_3342,In_3343,In_3344,In_3345,In_3346,In_3347,In_3348,In_3349,In_3350,In_3351,In_3352,In_3353,In_3354,In_3355,In_3356,In_3357,In_3358,In_3359,In_3360,In_3361,In_3362,In_3363,In_3364,In_3365,In_3366,In_3367,In_3368,In_3369,In_3370,In_3371,In_3372,In_3373,In_3374,In_3375,In_3376,In_3377,In_3378,In_3379,In_3380,In_3381,In_3382,In_3383,In_3384,In_3385,In_3386,In_3387,In_3388,In_3389,In_3390,In_3391,In_3392,In_3393,In_3394,In_3395,In_3396,In_3397,In_3398,In_3399,In_3400,In_3401,In_3402,In_3403,In_3404,In_3405,In_3406,In_3407,In_3408,In_3409,In_3410,In_3411,In_3412,In_3413,In_3414,In_3415,In_3416,In_3417,In_3418,In_3419,In_3420,In_3421,In_3422,In_3423,In_3424,In_3425,In_3426,In_3427,In_3428,In_3429,In_3430,In_3431,In_3432,In_3433,In_3434,In_3435,In_3436,In_3437,In_3438,In_3439,In_3440,In_3441,In_3442,In_3443,In_3444,In_3445,In_3446,In_3447,In_3448,In_3449,In_3450,In_3451,In_3452,In_3453,In_3454,In_3455,In_3456,In_3457,In_3458,In_3459,In_3460,In_3461,In_3462,In_3463,In_3464,In_3465,In_3466,In_3467,In_3468,In_3469,In_3470,In_3471,In_3472,In_3473,In_3474,In_3475,In_3476,In_3477,In_3478,In_3479,In_3480,In_3481,In_3482,In_3483,In_3484,In_3485,In_3486,In_3487,In_3488,In_3489,In_3490,In_3491,In_3492,In_3493,In_3494,In_3495,In_3496,In_3497,In_3498,In_3499,In_3500,In_3501,In_3502,In_3503,In_3504,In_3505,In_3506,In_3507,In_3508,In_3509,In_3510,In_3511,In_3512,In_3513,In_3514,In_3515,In_3516,In_3517,In_3518,In_3519,In_3520,In_3521,In_3522,In_3523,In_3524,In_3525,In_3526,In_3527,In_3528,In_3529,In_3530,In_3531,In_3532,In_3533,In_3534,In_3535,In_3536,In_3537,In_3538,In_3539,In_3540,In_3541,In_3542,In_3543,In_3544,In_3545,In_3546,In_3547,In_3548,In_3549,In_3550,In_3551,In_3552,In_3553,In_3554,In_3555,In_3556,In_3557,In_3558,In_3559,In_3560,In_3561,In_3562,In_3563,In_3564,In_3565,In_3566,In_3567,In_3568,In_3569,In_3570,In_3571,In_3572,In_3573,In_3574,In_3575,In_3576,In_3577,In_3578,In_3579,In_3580,In_3581,In_3582,In_3583,In_3584,In_3585,In_3586,In_3587,In_3588,In_3589,In_3590,In_3591,In_3592,In_3593,In_3594,In_3595,In_3596,In_3597,In_3598,In_3599,In_3600,In_3601,In_3602,In_3603,In_3604,In_3605,In_3606,In_3607,In_3608,In_3609,In_3610,In_3611,In_3612,In_3613,In_3614,In_3615,In_3616,In_3617,In_3618,In_3619,In_3620,In_3621,In_3622,In_3623,In_3624,In_3625,In_3626,In_3627,In_3628,In_3629,In_3630,In_3631,In_3632,In_3633,In_3634,In_3635,In_3636,In_3637,In_3638,In_3639,In_3640,In_3641,In_3642,In_3643,In_3644,In_3645,In_3646,In_3647,In_3648,In_3649,In_3650,In_3651,In_3652,In_3653,In_3654,In_3655,In_3656,In_3657,In_3658,In_3659,In_3660,In_3661,In_3662,In_3663,In_3664,In_3665,In_3666,In_3667,In_3668,In_3669,In_3670,In_3671,In_3672,In_3673,In_3674,In_3675,In_3676,In_3677,In_3678,In_3679,In_3680,In_3681,In_3682,In_3683,In_3684,In_3685,In_3686,In_3687,In_3688,In_3689,In_3690,In_3691,In_3692,In_3693,In_3694,In_3695,In_3696,In_3697,In_3698,In_3699,In_3700,In_3701,In_3702,In_3703,In_3704,In_3705,In_3706,In_3707,In_3708,In_3709,In_3710,In_3711,In_3712,In_3713,In_3714,In_3715,In_3716,In_3717,In_3718,In_3719,In_3720,In_3721,In_3722,In_3723,In_3724,In_3725,In_3726,In_3727,In_3728,In_3729,In_3730,In_3731,In_3732,In_3733,In_3734,In_3735,In_3736,In_3737,In_3738,In_3739,In_3740,In_3741,In_3742,In_3743,In_3744,In_3745,In_3746,In_3747,In_3748,In_3749,In_3750,In_3751,In_3752,In_3753,In_3754,In_3755,In_3756,In_3757,In_3758,In_3759,In_3760,In_3761,In_3762,In_3763,In_3764,In_3765,In_3766,In_3767,In_3768,In_3769,In_3770,In_3771,In_3772,In_3773,In_3774,In_3775,In_3776,In_3777,In_3778,In_3779,In_3780,In_3781,In_3782,In_3783,In_3784,In_3785,In_3786,In_3787,In_3788,In_3789,In_3790,In_3791,In_3792,In_3793,In_3794,In_3795,In_3796,In_3797,In_3798,In_3799,In_3800,In_3801,In_3802,In_3803,In_3804,In_3805,In_3806,In_3807,In_3808,In_3809,In_3810,In_3811,In_3812,In_3813,In_3814,In_3815,In_3816,In_3817,In_3818,In_3819,In_3820,In_3821,In_3822,In_3823,In_3824,In_3825,In_3826,In_3827,In_3828,In_3829,In_3830,In_3831,In_3832,In_3833,In_3834,In_3835,In_3836,In_3837,In_3838,In_3839,In_3840,In_3841,In_3842,In_3843,In_3844,In_3845,In_3846,In_3847,In_3848,In_3849,In_3850,In_3851,In_3852,In_3853,In_3854,In_3855,In_3856,In_3857,In_3858,In_3859,In_3860,In_3861,In_3862,In_3863,In_3864,In_3865,In_3866,In_3867,In_3868,In_3869,In_3870,In_3871,In_3872,In_3873,In_3874,In_3875,In_3876,In_3877,In_3878,In_3879,In_3880,In_3881,In_3882,In_3883,In_3884,In_3885,In_3886,In_3887,In_3888,In_3889,In_3890,In_3891,In_3892,In_3893,In_3894,In_3895,In_3896,In_3897,In_3898,In_3899,In_3900,In_3901,In_3902,In_3903,In_3904,In_3905,In_3906,In_3907,In_3908,In_3909,In_3910,In_3911,In_3912,In_3913,In_3914,In_3915,In_3916,In_3917,In_3918,In_3919,In_3920,In_3921,In_3922,In_3923,In_3924,In_3925,In_3926,In_3927,In_3928,In_3929,In_3930,In_3931,In_3932,In_3933,In_3934,In_3935,In_3936,In_3937,In_3938,In_3939,In_3940,In_3941,In_3942,In_3943,In_3944,In_3945,In_3946,In_3947,In_3948,In_3949,In_3950,In_3951,In_3952,In_3953,In_3954,In_3955,In_3956,In_3957,In_3958,In_3959,In_3960,In_3961,In_3962,In_3963,In_3964,In_3965,In_3966,In_3967,In_3968,In_3969,In_3970,In_3971,In_3972,In_3973,In_3974,In_3975,In_3976,In_3977,In_3978,In_3979,In_3980,In_3981,In_3982,In_3983,In_3984,In_3985,In_3986,In_3987,In_3988,In_3989,In_3990,In_3991,In_3992,In_3993,In_3994,In_3995,In_3996,In_3997,In_3998,In_3999,In_4000,In_4001,In_4002,In_4003,In_4004,In_4005,In_4006,In_4007,In_4008,In_4009,In_4010,In_4011,In_4012,In_4013,In_4014,In_4015,In_4016,In_4017,In_4018,In_4019,In_4020,In_4021,In_4022,In_4023,In_4024,In_4025,In_4026,In_4027,In_4028,In_4029,In_4030,In_4031,In_4032,In_4033,In_4034,In_4035,In_4036,In_4037,In_4038,In_4039,In_4040,In_4041,In_4042,In_4043,In_4044,In_4045,In_4046,In_4047,In_4048,In_4049,In_4050,In_4051,In_4052,In_4053,In_4054,In_4055,In_4056,In_4057,In_4058,In_4059,In_4060,In_4061,In_4062,In_4063,In_4064,In_4065,In_4066,In_4067,In_4068,In_4069,In_4070,In_4071,In_4072,In_4073,In_4074,In_4075,In_4076,In_4077,In_4078,In_4079,In_4080,In_4081,In_4082,In_4083,In_4084,In_4085,In_4086,In_4087,In_4088,In_4089,In_4090,In_4091,In_4092,In_4093,In_4094,In_4095,In_4096,In_4097,In_4098,In_4099,In_4100,In_4101,In_4102,In_4103,In_4104,In_4105,In_4106,In_4107,In_4108,In_4109,In_4110,In_4111,In_4112,In_4113,In_4114,In_4115,In_4116,In_4117,In_4118,In_4119,In_4120,In_4121,In_4122,In_4123,In_4124,In_4125,In_4126,In_4127,In_4128,In_4129,In_4130,In_4131,In_4132,In_4133,In_4134,In_4135,In_4136,In_4137,In_4138,In_4139,In_4140,In_4141,In_4142,In_4143,In_4144,In_4145,In_4146,In_4147,In_4148,In_4149,In_4150,In_4151,In_4152,In_4153,In_4154,In_4155,In_4156,In_4157,In_4158,In_4159,In_4160,In_4161,In_4162,In_4163,In_4164,In_4165,In_4166,In_4167,In_4168,In_4169,In_4170,In_4171,In_4172,In_4173,In_4174,In_4175,In_4176,In_4177,In_4178,In_4179,In_4180,In_4181,In_4182,In_4183,In_4184,In_4185,In_4186,In_4187,In_4188,In_4189,In_4190,In_4191,In_4192,In_4193,In_4194,In_4195,In_4196,In_4197,In_4198,In_4199,In_4200,In_4201,In_4202,In_4203,In_4204,In_4205,In_4206,In_4207,In_4208,In_4209,In_4210,In_4211,In_4212,In_4213,In_4214,In_4215,In_4216,In_4217,In_4218,In_4219,In_4220,In_4221,In_4222,In_4223,In_4224,In_4225,In_4226,In_4227,In_4228,In_4229,In_4230,In_4231,In_4232,In_4233,In_4234,In_4235,In_4236,In_4237,In_4238,In_4239,In_4240,In_4241,In_4242,In_4243,In_4244,In_4245,In_4246,In_4247,In_4248,In_4249,In_4250,In_4251,In_4252,In_4253,In_4254,In_4255,In_4256,In_4257,In_4258,In_4259,In_4260,In_4261,In_4262,In_4263,In_4264,In_4265,In_4266,In_4267,In_4268,In_4269,In_4270,In_4271,In_4272,In_4273,In_4274,In_4275,In_4276,In_4277,In_4278,In_4279,In_4280,In_4281,In_4282,In_4283,In_4284,In_4285,In_4286,In_4287,In_4288,In_4289,In_4290,In_4291,In_4292,In_4293,In_4294,In_4295,In_4296,In_4297,In_4298,In_4299,In_4300,In_4301,In_4302,In_4303,In_4304,In_4305,In_4306,In_4307,In_4308,In_4309,In_4310,In_4311,In_4312,In_4313,In_4314,In_4315,In_4316,In_4317,In_4318,In_4319,In_4320,In_4321,In_4322,In_4323,In_4324,In_4325,In_4326,In_4327,In_4328,In_4329,In_4330,In_4331,In_4332,In_4333,In_4334,In_4335,In_4336,In_4337,In_4338,In_4339,In_4340,In_4341,In_4342,In_4343,In_4344,In_4345,In_4346,In_4347,In_4348,In_4349,In_4350,In_4351,In_4352,In_4353,In_4354,In_4355,In_4356,In_4357,In_4358,In_4359,In_4360,In_4361,In_4362,In_4363,In_4364,In_4365,In_4366,In_4367,In_4368,In_4369,In_4370,In_4371,In_4372,In_4373,In_4374,In_4375,In_4376,In_4377,In_4378,In_4379,In_4380,In_4381,In_4382,In_4383,In_4384,In_4385,In_4386,In_4387,In_4388,In_4389,In_4390,In_4391,In_4392,In_4393,In_4394,In_4395,In_4396,In_4397,In_4398,In_4399,In_4400,In_4401,In_4402,In_4403,In_4404,In_4405,In_4406,In_4407,In_4408,In_4409,In_4410,In_4411,In_4412,In_4413,In_4414,In_4415,In_4416,In_4417,In_4418,In_4419,In_4420,In_4421,In_4422,In_4423,In_4424,In_4425,In_4426,In_4427,In_4428,In_4429,In_4430,In_4431,In_4432,In_4433,In_4434,In_4435,In_4436,In_4437,In_4438,In_4439,In_4440,In_4441,In_4442,In_4443,In_4444,In_4445,In_4446,In_4447,In_4448,In_4449,In_4450,In_4451,In_4452,In_4453,In_4454,In_4455,In_4456,In_4457,In_4458,In_4459,In_4460,In_4461,In_4462,In_4463,In_4464,In_4465,In_4466,In_4467,In_4468,In_4469,In_4470,In_4471,In_4472,In_4473,In_4474,In_4475,In_4476,In_4477,In_4478,In_4479,In_4480,In_4481,In_4482,In_4483,In_4484,In_4485,In_4486,In_4487,In_4488,In_4489,In_4490,In_4491,In_4492,In_4493,In_4494,In_4495,In_4496,In_4497,In_4498,In_4499,In_4500,In_4501,In_4502,In_4503,In_4504,In_4505,In_4506,In_4507,In_4508,In_4509,In_4510,In_4511,In_4512,In_4513,In_4514,In_4515,In_4516,In_4517,In_4518,In_4519,In_4520,In_4521,In_4522,In_4523,In_4524,In_4525,In_4526,In_4527,In_4528,In_4529,In_4530,In_4531,In_4532,In_4533,In_4534,In_4535,In_4536,In_4537,In_4538,In_4539,In_4540,In_4541,In_4542,In_4543,In_4544,In_4545,In_4546,In_4547,In_4548,In_4549,In_4550,In_4551,In_4552,In_4553,In_4554,In_4555,In_4556,In_4557,In_4558,In_4559,In_4560,In_4561,In_4562,In_4563,In_4564,In_4565,In_4566,In_4567,In_4568,In_4569,In_4570,In_4571,In_4572,In_4573,In_4574,In_4575,In_4576,In_4577,In_4578,In_4579,In_4580,In_4581,In_4582,In_4583,In_4584,In_4585,In_4586,In_4587,In_4588,In_4589,In_4590,In_4591,In_4592,In_4593,In_4594,In_4595,In_4596,In_4597,In_4598,In_4599,In_4600,In_4601,In_4602,In_4603,In_4604,In_4605,In_4606,In_4607,In_4608,In_4609,In_4610,In_4611,In_4612,In_4613,In_4614,In_4615,In_4616,In_4617,In_4618,In_4619,In_4620,In_4621,In_4622,In_4623,In_4624,In_4625,In_4626,In_4627,In_4628,In_4629,In_4630,In_4631,In_4632,In_4633,In_4634,In_4635,In_4636,In_4637,In_4638,In_4639,In_4640,In_4641,In_4642,In_4643,In_4644,In_4645,In_4646,In_4647,In_4648,In_4649,In_4650,In_4651,In_4652,In_4653,In_4654,In_4655,In_4656,In_4657,In_4658,In_4659,In_4660,In_4661,In_4662,In_4663,In_4664,In_4665,In_4666,In_4667,In_4668,In_4669,In_4670,In_4671,In_4672,In_4673,In_4674,In_4675,In_4676,In_4677,In_4678,In_4679,In_4680,In_4681,In_4682,In_4683,In_4684,In_4685,In_4686,In_4687,In_4688,In_4689,In_4690,In_4691,In_4692,In_4693,In_4694,In_4695,In_4696,In_4697,In_4698,In_4699,In_4700,In_4701,In_4702,In_4703,In_4704,In_4705,In_4706,In_4707,In_4708,In_4709,In_4710,In_4711,In_4712,In_4713,In_4714,In_4715,In_4716,In_4717,In_4718,In_4719,In_4720,In_4721,In_4722,In_4723,In_4724,In_4725,In_4726,In_4727,In_4728,In_4729,In_4730,In_4731,In_4732,In_4733,In_4734,In_4735,In_4736,In_4737,In_4738,In_4739,In_4740,In_4741,In_4742,In_4743,In_4744,In_4745,In_4746,In_4747,In_4748,In_4749,In_4750,In_4751,In_4752,In_4753,In_4754,In_4755,In_4756,In_4757,In_4758,In_4759,In_4760,In_4761,In_4762,In_4763,In_4764,In_4765,In_4766,In_4767,In_4768,In_4769,In_4770,In_4771,In_4772,In_4773,In_4774,In_4775,In_4776,In_4777,In_4778,In_4779,In_4780,In_4781,In_4782,In_4783,In_4784,In_4785,In_4786,In_4787,In_4788,In_4789,In_4790,In_4791,In_4792,In_4793,In_4794,In_4795,In_4796,In_4797,In_4798,In_4799,In_4800,In_4801,In_4802,In_4803,In_4804,In_4805,In_4806,In_4807,In_4808,In_4809,In_4810,In_4811,In_4812,In_4813,In_4814,In_4815,In_4816,In_4817,In_4818,In_4819,In_4820,In_4821,In_4822,In_4823,In_4824,In_4825,In_4826,In_4827,In_4828,In_4829,In_4830,In_4831,In_4832,In_4833,In_4834,In_4835,In_4836,In_4837,In_4838,In_4839,In_4840,In_4841,In_4842,In_4843,In_4844,In_4845,In_4846,In_4847,In_4848,In_4849,In_4850,In_4851,In_4852,In_4853,In_4854,In_4855,In_4856,In_4857,In_4858,In_4859,In_4860,In_4861,In_4862,In_4863,In_4864,In_4865,In_4866,In_4867,In_4868,In_4869,In_4870,In_4871,In_4872,In_4873,In_4874,In_4875,In_4876,In_4877,In_4878,In_4879,In_4880,In_4881,In_4882,In_4883,In_4884,In_4885,In_4886,In_4887,In_4888,In_4889,In_4890,In_4891,In_4892,In_4893,In_4894,In_4895,In_4896,In_4897,In_4898,In_4899,In_4900,In_4901,In_4902,In_4903,In_4904,In_4905,In_4906,In_4907,In_4908,In_4909,In_4910,In_4911,In_4912,In_4913,In_4914,In_4915,In_4916,In_4917,In_4918,In_4919,In_4920,In_4921,In_4922,In_4923,In_4924,In_4925,In_4926,In_4927,In_4928,In_4929,In_4930,In_4931,In_4932,In_4933,In_4934,In_4935,In_4936,In_4937,In_4938,In_4939,In_4940,In_4941,In_4942,In_4943,In_4944,In_4945,In_4946,In_4947,In_4948,In_4949,In_4950,In_4951,In_4952,In_4953,In_4954,In_4955,In_4956,In_4957,In_4958,In_4959,In_4960,In_4961,In_4962,In_4963,In_4964,In_4965,In_4966,In_4967,In_4968,In_4969,In_4970,In_4971,In_4972,In_4973,In_4974,In_4975,In_4976,In_4977,In_4978,In_4979,In_4980,In_4981,In_4982,In_4983,In_4984,In_4985,In_4986,In_4987,In_4988,In_4989,In_4990,In_4991,In_4992,In_4993,In_4994,In_4995,In_4996,In_4997,In_4998,In_4999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499,O_3500,O_3501,O_3502,O_3503,O_3504,O_3505,O_3506,O_3507,O_3508,O_3509,O_3510,O_3511,O_3512,O_3513,O_3514,O_3515,O_3516,O_3517,O_3518,O_3519,O_3520,O_3521,O_3522,O_3523,O_3524,O_3525,O_3526,O_3527,O_3528,O_3529,O_3530,O_3531,O_3532,O_3533,O_3534,O_3535,O_3536,O_3537,O_3538,O_3539,O_3540,O_3541,O_3542,O_3543,O_3544,O_3545,O_3546,O_3547,O_3548,O_3549,O_3550,O_3551,O_3552,O_3553,O_3554,O_3555,O_3556,O_3557,O_3558,O_3559,O_3560,O_3561,O_3562,O_3563,O_3564,O_3565,O_3566,O_3567,O_3568,O_3569,O_3570,O_3571,O_3572,O_3573,O_3574,O_3575,O_3576,O_3577,O_3578,O_3579,O_3580,O_3581,O_3582,O_3583,O_3584,O_3585,O_3586,O_3587,O_3588,O_3589,O_3590,O_3591,O_3592,O_3593,O_3594,O_3595,O_3596,O_3597,O_3598,O_3599,O_3600,O_3601,O_3602,O_3603,O_3604,O_3605,O_3606,O_3607,O_3608,O_3609,O_3610,O_3611,O_3612,O_3613,O_3614,O_3615,O_3616,O_3617,O_3618,O_3619,O_3620,O_3621,O_3622,O_3623,O_3624,O_3625,O_3626,O_3627,O_3628,O_3629,O_3630,O_3631,O_3632,O_3633,O_3634,O_3635,O_3636,O_3637,O_3638,O_3639,O_3640,O_3641,O_3642,O_3643,O_3644,O_3645,O_3646,O_3647,O_3648,O_3649,O_3650,O_3651,O_3652,O_3653,O_3654,O_3655,O_3656,O_3657,O_3658,O_3659,O_3660,O_3661,O_3662,O_3663,O_3664,O_3665,O_3666,O_3667,O_3668,O_3669,O_3670,O_3671,O_3672,O_3673,O_3674,O_3675,O_3676,O_3677,O_3678,O_3679,O_3680,O_3681,O_3682,O_3683,O_3684,O_3685,O_3686,O_3687,O_3688,O_3689,O_3690,O_3691,O_3692,O_3693,O_3694,O_3695,O_3696,O_3697,O_3698,O_3699,O_3700,O_3701,O_3702,O_3703,O_3704,O_3705,O_3706,O_3707,O_3708,O_3709,O_3710,O_3711,O_3712,O_3713,O_3714,O_3715,O_3716,O_3717,O_3718,O_3719,O_3720,O_3721,O_3722,O_3723,O_3724,O_3725,O_3726,O_3727,O_3728,O_3729,O_3730,O_3731,O_3732,O_3733,O_3734,O_3735,O_3736,O_3737,O_3738,O_3739,O_3740,O_3741,O_3742,O_3743,O_3744,O_3745,O_3746,O_3747,O_3748,O_3749,O_3750,O_3751,O_3752,O_3753,O_3754,O_3755,O_3756,O_3757,O_3758,O_3759,O_3760,O_3761,O_3762,O_3763,O_3764,O_3765,O_3766,O_3767,O_3768,O_3769,O_3770,O_3771,O_3772,O_3773,O_3774,O_3775,O_3776,O_3777,O_3778,O_3779,O_3780,O_3781,O_3782,O_3783,O_3784,O_3785,O_3786,O_3787,O_3788,O_3789,O_3790,O_3791,O_3792,O_3793,O_3794,O_3795,O_3796,O_3797,O_3798,O_3799,O_3800,O_3801,O_3802,O_3803,O_3804,O_3805,O_3806,O_3807,O_3808,O_3809,O_3810,O_3811,O_3812,O_3813,O_3814,O_3815,O_3816,O_3817,O_3818,O_3819,O_3820,O_3821,O_3822,O_3823,O_3824,O_3825,O_3826,O_3827,O_3828,O_3829,O_3830,O_3831,O_3832,O_3833,O_3834,O_3835,O_3836,O_3837,O_3838,O_3839,O_3840,O_3841,O_3842,O_3843,O_3844,O_3845,O_3846,O_3847,O_3848,O_3849,O_3850,O_3851,O_3852,O_3853,O_3854,O_3855,O_3856,O_3857,O_3858,O_3859,O_3860,O_3861,O_3862,O_3863,O_3864,O_3865,O_3866,O_3867,O_3868,O_3869,O_3870,O_3871,O_3872,O_3873,O_3874,O_3875,O_3876,O_3877,O_3878,O_3879,O_3880,O_3881,O_3882,O_3883,O_3884,O_3885,O_3886,O_3887,O_3888,O_3889,O_3890,O_3891,O_3892,O_3893,O_3894,O_3895,O_3896,O_3897,O_3898,O_3899,O_3900,O_3901,O_3902,O_3903,O_3904,O_3905,O_3906,O_3907,O_3908,O_3909,O_3910,O_3911,O_3912,O_3913,O_3914,O_3915,O_3916,O_3917,O_3918,O_3919,O_3920,O_3921,O_3922,O_3923,O_3924,O_3925,O_3926,O_3927,O_3928,O_3929,O_3930,O_3931,O_3932,O_3933,O_3934,O_3935,O_3936,O_3937,O_3938,O_3939,O_3940,O_3941,O_3942,O_3943,O_3944,O_3945,O_3946,O_3947,O_3948,O_3949,O_3950,O_3951,O_3952,O_3953,O_3954,O_3955,O_3956,O_3957,O_3958,O_3959,O_3960,O_3961,O_3962,O_3963,O_3964,O_3965,O_3966,O_3967,O_3968,O_3969,O_3970,O_3971,O_3972,O_3973,O_3974,O_3975,O_3976,O_3977,O_3978,O_3979,O_3980,O_3981,O_3982,O_3983,O_3984,O_3985,O_3986,O_3987,O_3988,O_3989,O_3990,O_3991,O_3992,O_3993,O_3994,O_3995,O_3996,O_3997,O_3998,O_3999,O_4000,O_4001,O_4002,O_4003,O_4004,O_4005,O_4006,O_4007,O_4008,O_4009,O_4010,O_4011,O_4012,O_4013,O_4014,O_4015,O_4016,O_4017,O_4018,O_4019,O_4020,O_4021,O_4022,O_4023,O_4024,O_4025,O_4026,O_4027,O_4028,O_4029,O_4030,O_4031,O_4032,O_4033,O_4034,O_4035,O_4036,O_4037,O_4038,O_4039,O_4040,O_4041,O_4042,O_4043,O_4044,O_4045,O_4046,O_4047,O_4048,O_4049,O_4050,O_4051,O_4052,O_4053,O_4054,O_4055,O_4056,O_4057,O_4058,O_4059,O_4060,O_4061,O_4062,O_4063,O_4064,O_4065,O_4066,O_4067,O_4068,O_4069,O_4070,O_4071,O_4072,O_4073,O_4074,O_4075,O_4076,O_4077,O_4078,O_4079,O_4080,O_4081,O_4082,O_4083,O_4084,O_4085,O_4086,O_4087,O_4088,O_4089,O_4090,O_4091,O_4092,O_4093,O_4094,O_4095,O_4096,O_4097,O_4098,O_4099,O_4100,O_4101,O_4102,O_4103,O_4104,O_4105,O_4106,O_4107,O_4108,O_4109,O_4110,O_4111,O_4112,O_4113,O_4114,O_4115,O_4116,O_4117,O_4118,O_4119,O_4120,O_4121,O_4122,O_4123,O_4124,O_4125,O_4126,O_4127,O_4128,O_4129,O_4130,O_4131,O_4132,O_4133,O_4134,O_4135,O_4136,O_4137,O_4138,O_4139,O_4140,O_4141,O_4142,O_4143,O_4144,O_4145,O_4146,O_4147,O_4148,O_4149,O_4150,O_4151,O_4152,O_4153,O_4154,O_4155,O_4156,O_4157,O_4158,O_4159,O_4160,O_4161,O_4162,O_4163,O_4164,O_4165,O_4166,O_4167,O_4168,O_4169,O_4170,O_4171,O_4172,O_4173,O_4174,O_4175,O_4176,O_4177,O_4178,O_4179,O_4180,O_4181,O_4182,O_4183,O_4184,O_4185,O_4186,O_4187,O_4188,O_4189,O_4190,O_4191,O_4192,O_4193,O_4194,O_4195,O_4196,O_4197,O_4198,O_4199,O_4200,O_4201,O_4202,O_4203,O_4204,O_4205,O_4206,O_4207,O_4208,O_4209,O_4210,O_4211,O_4212,O_4213,O_4214,O_4215,O_4216,O_4217,O_4218,O_4219,O_4220,O_4221,O_4222,O_4223,O_4224,O_4225,O_4226,O_4227,O_4228,O_4229,O_4230,O_4231,O_4232,O_4233,O_4234,O_4235,O_4236,O_4237,O_4238,O_4239,O_4240,O_4241,O_4242,O_4243,O_4244,O_4245,O_4246,O_4247,O_4248,O_4249,O_4250,O_4251,O_4252,O_4253,O_4254,O_4255,O_4256,O_4257,O_4258,O_4259,O_4260,O_4261,O_4262,O_4263,O_4264,O_4265,O_4266,O_4267,O_4268,O_4269,O_4270,O_4271,O_4272,O_4273,O_4274,O_4275,O_4276,O_4277,O_4278,O_4279,O_4280,O_4281,O_4282,O_4283,O_4284,O_4285,O_4286,O_4287,O_4288,O_4289,O_4290,O_4291,O_4292,O_4293,O_4294,O_4295,O_4296,O_4297,O_4298,O_4299,O_4300,O_4301,O_4302,O_4303,O_4304,O_4305,O_4306,O_4307,O_4308,O_4309,O_4310,O_4311,O_4312,O_4313,O_4314,O_4315,O_4316,O_4317,O_4318,O_4319,O_4320,O_4321,O_4322,O_4323,O_4324,O_4325,O_4326,O_4327,O_4328,O_4329,O_4330,O_4331,O_4332,O_4333,O_4334,O_4335,O_4336,O_4337,O_4338,O_4339,O_4340,O_4341,O_4342,O_4343,O_4344,O_4345,O_4346,O_4347,O_4348,O_4349,O_4350,O_4351,O_4352,O_4353,O_4354,O_4355,O_4356,O_4357,O_4358,O_4359,O_4360,O_4361,O_4362,O_4363,O_4364,O_4365,O_4366,O_4367,O_4368,O_4369,O_4370,O_4371,O_4372,O_4373,O_4374,O_4375,O_4376,O_4377,O_4378,O_4379,O_4380,O_4381,O_4382,O_4383,O_4384,O_4385,O_4386,O_4387,O_4388,O_4389,O_4390,O_4391,O_4392,O_4393,O_4394,O_4395,O_4396,O_4397,O_4398,O_4399,O_4400,O_4401,O_4402,O_4403,O_4404,O_4405,O_4406,O_4407,O_4408,O_4409,O_4410,O_4411,O_4412,O_4413,O_4414,O_4415,O_4416,O_4417,O_4418,O_4419,O_4420,O_4421,O_4422,O_4423,O_4424,O_4425,O_4426,O_4427,O_4428,O_4429,O_4430,O_4431,O_4432,O_4433,O_4434,O_4435,O_4436,O_4437,O_4438,O_4439,O_4440,O_4441,O_4442,O_4443,O_4444,O_4445,O_4446,O_4447,O_4448,O_4449,O_4450,O_4451,O_4452,O_4453,O_4454,O_4455,O_4456,O_4457,O_4458,O_4459,O_4460,O_4461,O_4462,O_4463,O_4464,O_4465,O_4466,O_4467,O_4468,O_4469,O_4470,O_4471,O_4472,O_4473,O_4474,O_4475,O_4476,O_4477,O_4478,O_4479,O_4480,O_4481,O_4482,O_4483,O_4484,O_4485,O_4486,O_4487,O_4488,O_4489,O_4490,O_4491,O_4492,O_4493,O_4494,O_4495,O_4496,O_4497,O_4498,O_4499,O_4500,O_4501,O_4502,O_4503,O_4504,O_4505,O_4506,O_4507,O_4508,O_4509,O_4510,O_4511,O_4512,O_4513,O_4514,O_4515,O_4516,O_4517,O_4518,O_4519,O_4520,O_4521,O_4522,O_4523,O_4524,O_4525,O_4526,O_4527,O_4528,O_4529,O_4530,O_4531,O_4532,O_4533,O_4534,O_4535,O_4536,O_4537,O_4538,O_4539,O_4540,O_4541,O_4542,O_4543,O_4544,O_4545,O_4546,O_4547,O_4548,O_4549,O_4550,O_4551,O_4552,O_4553,O_4554,O_4555,O_4556,O_4557,O_4558,O_4559,O_4560,O_4561,O_4562,O_4563,O_4564,O_4565,O_4566,O_4567,O_4568,O_4569,O_4570,O_4571,O_4572,O_4573,O_4574,O_4575,O_4576,O_4577,O_4578,O_4579,O_4580,O_4581,O_4582,O_4583,O_4584,O_4585,O_4586,O_4587,O_4588,O_4589,O_4590,O_4591,O_4592,O_4593,O_4594,O_4595,O_4596,O_4597,O_4598,O_4599,O_4600,O_4601,O_4602,O_4603,O_4604,O_4605,O_4606,O_4607,O_4608,O_4609,O_4610,O_4611,O_4612,O_4613,O_4614,O_4615,O_4616,O_4617,O_4618,O_4619,O_4620,O_4621,O_4622,O_4623,O_4624,O_4625,O_4626,O_4627,O_4628,O_4629,O_4630,O_4631,O_4632,O_4633,O_4634,O_4635,O_4636,O_4637,O_4638,O_4639,O_4640,O_4641,O_4642,O_4643,O_4644,O_4645,O_4646,O_4647,O_4648,O_4649,O_4650,O_4651,O_4652,O_4653,O_4654,O_4655,O_4656,O_4657,O_4658,O_4659,O_4660,O_4661,O_4662,O_4663,O_4664,O_4665,O_4666,O_4667,O_4668,O_4669,O_4670,O_4671,O_4672,O_4673,O_4674,O_4675,O_4676,O_4677,O_4678,O_4679,O_4680,O_4681,O_4682,O_4683,O_4684,O_4685,O_4686,O_4687,O_4688,O_4689,O_4690,O_4691,O_4692,O_4693,O_4694,O_4695,O_4696,O_4697,O_4698,O_4699,O_4700,O_4701,O_4702,O_4703,O_4704,O_4705,O_4706,O_4707,O_4708,O_4709,O_4710,O_4711,O_4712,O_4713,O_4714,O_4715,O_4716,O_4717,O_4718,O_4719,O_4720,O_4721,O_4722,O_4723,O_4724,O_4725,O_4726,O_4727,O_4728,O_4729,O_4730,O_4731,O_4732,O_4733,O_4734,O_4735,O_4736,O_4737,O_4738,O_4739,O_4740,O_4741,O_4742,O_4743,O_4744,O_4745,O_4746,O_4747,O_4748,O_4749,O_4750,O_4751,O_4752,O_4753,O_4754,O_4755,O_4756,O_4757,O_4758,O_4759,O_4760,O_4761,O_4762,O_4763,O_4764,O_4765,O_4766,O_4767,O_4768,O_4769,O_4770,O_4771,O_4772,O_4773,O_4774,O_4775,O_4776,O_4777,O_4778,O_4779,O_4780,O_4781,O_4782,O_4783,O_4784,O_4785,O_4786,O_4787,O_4788,O_4789,O_4790,O_4791,O_4792,O_4793,O_4794,O_4795,O_4796,O_4797,O_4798,O_4799,O_4800,O_4801,O_4802,O_4803,O_4804,O_4805,O_4806,O_4807,O_4808,O_4809,O_4810,O_4811,O_4812,O_4813,O_4814,O_4815,O_4816,O_4817,O_4818,O_4819,O_4820,O_4821,O_4822,O_4823,O_4824,O_4825,O_4826,O_4827,O_4828,O_4829,O_4830,O_4831,O_4832,O_4833,O_4834,O_4835,O_4836,O_4837,O_4838,O_4839,O_4840,O_4841,O_4842,O_4843,O_4844,O_4845,O_4846,O_4847,O_4848,O_4849,O_4850,O_4851,O_4852,O_4853,O_4854,O_4855,O_4856,O_4857,O_4858,O_4859,O_4860,O_4861,O_4862,O_4863,O_4864,O_4865,O_4866,O_4867,O_4868,O_4869,O_4870,O_4871,O_4872,O_4873,O_4874,O_4875,O_4876,O_4877,O_4878,O_4879,O_4880,O_4881,O_4882,O_4883,O_4884,O_4885,O_4886,O_4887,O_4888,O_4889,O_4890,O_4891,O_4892,O_4893,O_4894,O_4895,O_4896,O_4897,O_4898,O_4899,O_4900,O_4901,O_4902,O_4903,O_4904,O_4905,O_4906,O_4907,O_4908,O_4909,O_4910,O_4911,O_4912,O_4913,O_4914,O_4915,O_4916,O_4917,O_4918,O_4919,O_4920,O_4921,O_4922,O_4923,O_4924,O_4925,O_4926,O_4927,O_4928,O_4929,O_4930,O_4931,O_4932,O_4933,O_4934,O_4935,O_4936,O_4937,O_4938,O_4939,O_4940,O_4941,O_4942,O_4943,O_4944,O_4945,O_4946,O_4947,O_4948,O_4949,O_4950,O_4951,O_4952,O_4953,O_4954,O_4955,O_4956,O_4957,O_4958,O_4959,O_4960,O_4961,O_4962,O_4963,O_4964,O_4965,O_4966,O_4967,O_4968,O_4969,O_4970,O_4971,O_4972,O_4973,O_4974,O_4975,O_4976,O_4977,O_4978,O_4979,O_4980,O_4981,O_4982,O_4983,O_4984,O_4985,O_4986,O_4987,O_4988,O_4989,O_4990,O_4991,O_4992,O_4993,O_4994,O_4995,O_4996,O_4997,O_4998,O_4999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,In_3000,In_3001,In_3002,In_3003,In_3004,In_3005,In_3006,In_3007,In_3008,In_3009,In_3010,In_3011,In_3012,In_3013,In_3014,In_3015,In_3016,In_3017,In_3018,In_3019,In_3020,In_3021,In_3022,In_3023,In_3024,In_3025,In_3026,In_3027,In_3028,In_3029,In_3030,In_3031,In_3032,In_3033,In_3034,In_3035,In_3036,In_3037,In_3038,In_3039,In_3040,In_3041,In_3042,In_3043,In_3044,In_3045,In_3046,In_3047,In_3048,In_3049,In_3050,In_3051,In_3052,In_3053,In_3054,In_3055,In_3056,In_3057,In_3058,In_3059,In_3060,In_3061,In_3062,In_3063,In_3064,In_3065,In_3066,In_3067,In_3068,In_3069,In_3070,In_3071,In_3072,In_3073,In_3074,In_3075,In_3076,In_3077,In_3078,In_3079,In_3080,In_3081,In_3082,In_3083,In_3084,In_3085,In_3086,In_3087,In_3088,In_3089,In_3090,In_3091,In_3092,In_3093,In_3094,In_3095,In_3096,In_3097,In_3098,In_3099,In_3100,In_3101,In_3102,In_3103,In_3104,In_3105,In_3106,In_3107,In_3108,In_3109,In_3110,In_3111,In_3112,In_3113,In_3114,In_3115,In_3116,In_3117,In_3118,In_3119,In_3120,In_3121,In_3122,In_3123,In_3124,In_3125,In_3126,In_3127,In_3128,In_3129,In_3130,In_3131,In_3132,In_3133,In_3134,In_3135,In_3136,In_3137,In_3138,In_3139,In_3140,In_3141,In_3142,In_3143,In_3144,In_3145,In_3146,In_3147,In_3148,In_3149,In_3150,In_3151,In_3152,In_3153,In_3154,In_3155,In_3156,In_3157,In_3158,In_3159,In_3160,In_3161,In_3162,In_3163,In_3164,In_3165,In_3166,In_3167,In_3168,In_3169,In_3170,In_3171,In_3172,In_3173,In_3174,In_3175,In_3176,In_3177,In_3178,In_3179,In_3180,In_3181,In_3182,In_3183,In_3184,In_3185,In_3186,In_3187,In_3188,In_3189,In_3190,In_3191,In_3192,In_3193,In_3194,In_3195,In_3196,In_3197,In_3198,In_3199,In_3200,In_3201,In_3202,In_3203,In_3204,In_3205,In_3206,In_3207,In_3208,In_3209,In_3210,In_3211,In_3212,In_3213,In_3214,In_3215,In_3216,In_3217,In_3218,In_3219,In_3220,In_3221,In_3222,In_3223,In_3224,In_3225,In_3226,In_3227,In_3228,In_3229,In_3230,In_3231,In_3232,In_3233,In_3234,In_3235,In_3236,In_3237,In_3238,In_3239,In_3240,In_3241,In_3242,In_3243,In_3244,In_3245,In_3246,In_3247,In_3248,In_3249,In_3250,In_3251,In_3252,In_3253,In_3254,In_3255,In_3256,In_3257,In_3258,In_3259,In_3260,In_3261,In_3262,In_3263,In_3264,In_3265,In_3266,In_3267,In_3268,In_3269,In_3270,In_3271,In_3272,In_3273,In_3274,In_3275,In_3276,In_3277,In_3278,In_3279,In_3280,In_3281,In_3282,In_3283,In_3284,In_3285,In_3286,In_3287,In_3288,In_3289,In_3290,In_3291,In_3292,In_3293,In_3294,In_3295,In_3296,In_3297,In_3298,In_3299,In_3300,In_3301,In_3302,In_3303,In_3304,In_3305,In_3306,In_3307,In_3308,In_3309,In_3310,In_3311,In_3312,In_3313,In_3314,In_3315,In_3316,In_3317,In_3318,In_3319,In_3320,In_3321,In_3322,In_3323,In_3324,In_3325,In_3326,In_3327,In_3328,In_3329,In_3330,In_3331,In_3332,In_3333,In_3334,In_3335,In_3336,In_3337,In_3338,In_3339,In_3340,In_3341,In_3342,In_3343,In_3344,In_3345,In_3346,In_3347,In_3348,In_3349,In_3350,In_3351,In_3352,In_3353,In_3354,In_3355,In_3356,In_3357,In_3358,In_3359,In_3360,In_3361,In_3362,In_3363,In_3364,In_3365,In_3366,In_3367,In_3368,In_3369,In_3370,In_3371,In_3372,In_3373,In_3374,In_3375,In_3376,In_3377,In_3378,In_3379,In_3380,In_3381,In_3382,In_3383,In_3384,In_3385,In_3386,In_3387,In_3388,In_3389,In_3390,In_3391,In_3392,In_3393,In_3394,In_3395,In_3396,In_3397,In_3398,In_3399,In_3400,In_3401,In_3402,In_3403,In_3404,In_3405,In_3406,In_3407,In_3408,In_3409,In_3410,In_3411,In_3412,In_3413,In_3414,In_3415,In_3416,In_3417,In_3418,In_3419,In_3420,In_3421,In_3422,In_3423,In_3424,In_3425,In_3426,In_3427,In_3428,In_3429,In_3430,In_3431,In_3432,In_3433,In_3434,In_3435,In_3436,In_3437,In_3438,In_3439,In_3440,In_3441,In_3442,In_3443,In_3444,In_3445,In_3446,In_3447,In_3448,In_3449,In_3450,In_3451,In_3452,In_3453,In_3454,In_3455,In_3456,In_3457,In_3458,In_3459,In_3460,In_3461,In_3462,In_3463,In_3464,In_3465,In_3466,In_3467,In_3468,In_3469,In_3470,In_3471,In_3472,In_3473,In_3474,In_3475,In_3476,In_3477,In_3478,In_3479,In_3480,In_3481,In_3482,In_3483,In_3484,In_3485,In_3486,In_3487,In_3488,In_3489,In_3490,In_3491,In_3492,In_3493,In_3494,In_3495,In_3496,In_3497,In_3498,In_3499,In_3500,In_3501,In_3502,In_3503,In_3504,In_3505,In_3506,In_3507,In_3508,In_3509,In_3510,In_3511,In_3512,In_3513,In_3514,In_3515,In_3516,In_3517,In_3518,In_3519,In_3520,In_3521,In_3522,In_3523,In_3524,In_3525,In_3526,In_3527,In_3528,In_3529,In_3530,In_3531,In_3532,In_3533,In_3534,In_3535,In_3536,In_3537,In_3538,In_3539,In_3540,In_3541,In_3542,In_3543,In_3544,In_3545,In_3546,In_3547,In_3548,In_3549,In_3550,In_3551,In_3552,In_3553,In_3554,In_3555,In_3556,In_3557,In_3558,In_3559,In_3560,In_3561,In_3562,In_3563,In_3564,In_3565,In_3566,In_3567,In_3568,In_3569,In_3570,In_3571,In_3572,In_3573,In_3574,In_3575,In_3576,In_3577,In_3578,In_3579,In_3580,In_3581,In_3582,In_3583,In_3584,In_3585,In_3586,In_3587,In_3588,In_3589,In_3590,In_3591,In_3592,In_3593,In_3594,In_3595,In_3596,In_3597,In_3598,In_3599,In_3600,In_3601,In_3602,In_3603,In_3604,In_3605,In_3606,In_3607,In_3608,In_3609,In_3610,In_3611,In_3612,In_3613,In_3614,In_3615,In_3616,In_3617,In_3618,In_3619,In_3620,In_3621,In_3622,In_3623,In_3624,In_3625,In_3626,In_3627,In_3628,In_3629,In_3630,In_3631,In_3632,In_3633,In_3634,In_3635,In_3636,In_3637,In_3638,In_3639,In_3640,In_3641,In_3642,In_3643,In_3644,In_3645,In_3646,In_3647,In_3648,In_3649,In_3650,In_3651,In_3652,In_3653,In_3654,In_3655,In_3656,In_3657,In_3658,In_3659,In_3660,In_3661,In_3662,In_3663,In_3664,In_3665,In_3666,In_3667,In_3668,In_3669,In_3670,In_3671,In_3672,In_3673,In_3674,In_3675,In_3676,In_3677,In_3678,In_3679,In_3680,In_3681,In_3682,In_3683,In_3684,In_3685,In_3686,In_3687,In_3688,In_3689,In_3690,In_3691,In_3692,In_3693,In_3694,In_3695,In_3696,In_3697,In_3698,In_3699,In_3700,In_3701,In_3702,In_3703,In_3704,In_3705,In_3706,In_3707,In_3708,In_3709,In_3710,In_3711,In_3712,In_3713,In_3714,In_3715,In_3716,In_3717,In_3718,In_3719,In_3720,In_3721,In_3722,In_3723,In_3724,In_3725,In_3726,In_3727,In_3728,In_3729,In_3730,In_3731,In_3732,In_3733,In_3734,In_3735,In_3736,In_3737,In_3738,In_3739,In_3740,In_3741,In_3742,In_3743,In_3744,In_3745,In_3746,In_3747,In_3748,In_3749,In_3750,In_3751,In_3752,In_3753,In_3754,In_3755,In_3756,In_3757,In_3758,In_3759,In_3760,In_3761,In_3762,In_3763,In_3764,In_3765,In_3766,In_3767,In_3768,In_3769,In_3770,In_3771,In_3772,In_3773,In_3774,In_3775,In_3776,In_3777,In_3778,In_3779,In_3780,In_3781,In_3782,In_3783,In_3784,In_3785,In_3786,In_3787,In_3788,In_3789,In_3790,In_3791,In_3792,In_3793,In_3794,In_3795,In_3796,In_3797,In_3798,In_3799,In_3800,In_3801,In_3802,In_3803,In_3804,In_3805,In_3806,In_3807,In_3808,In_3809,In_3810,In_3811,In_3812,In_3813,In_3814,In_3815,In_3816,In_3817,In_3818,In_3819,In_3820,In_3821,In_3822,In_3823,In_3824,In_3825,In_3826,In_3827,In_3828,In_3829,In_3830,In_3831,In_3832,In_3833,In_3834,In_3835,In_3836,In_3837,In_3838,In_3839,In_3840,In_3841,In_3842,In_3843,In_3844,In_3845,In_3846,In_3847,In_3848,In_3849,In_3850,In_3851,In_3852,In_3853,In_3854,In_3855,In_3856,In_3857,In_3858,In_3859,In_3860,In_3861,In_3862,In_3863,In_3864,In_3865,In_3866,In_3867,In_3868,In_3869,In_3870,In_3871,In_3872,In_3873,In_3874,In_3875,In_3876,In_3877,In_3878,In_3879,In_3880,In_3881,In_3882,In_3883,In_3884,In_3885,In_3886,In_3887,In_3888,In_3889,In_3890,In_3891,In_3892,In_3893,In_3894,In_3895,In_3896,In_3897,In_3898,In_3899,In_3900,In_3901,In_3902,In_3903,In_3904,In_3905,In_3906,In_3907,In_3908,In_3909,In_3910,In_3911,In_3912,In_3913,In_3914,In_3915,In_3916,In_3917,In_3918,In_3919,In_3920,In_3921,In_3922,In_3923,In_3924,In_3925,In_3926,In_3927,In_3928,In_3929,In_3930,In_3931,In_3932,In_3933,In_3934,In_3935,In_3936,In_3937,In_3938,In_3939,In_3940,In_3941,In_3942,In_3943,In_3944,In_3945,In_3946,In_3947,In_3948,In_3949,In_3950,In_3951,In_3952,In_3953,In_3954,In_3955,In_3956,In_3957,In_3958,In_3959,In_3960,In_3961,In_3962,In_3963,In_3964,In_3965,In_3966,In_3967,In_3968,In_3969,In_3970,In_3971,In_3972,In_3973,In_3974,In_3975,In_3976,In_3977,In_3978,In_3979,In_3980,In_3981,In_3982,In_3983,In_3984,In_3985,In_3986,In_3987,In_3988,In_3989,In_3990,In_3991,In_3992,In_3993,In_3994,In_3995,In_3996,In_3997,In_3998,In_3999,In_4000,In_4001,In_4002,In_4003,In_4004,In_4005,In_4006,In_4007,In_4008,In_4009,In_4010,In_4011,In_4012,In_4013,In_4014,In_4015,In_4016,In_4017,In_4018,In_4019,In_4020,In_4021,In_4022,In_4023,In_4024,In_4025,In_4026,In_4027,In_4028,In_4029,In_4030,In_4031,In_4032,In_4033,In_4034,In_4035,In_4036,In_4037,In_4038,In_4039,In_4040,In_4041,In_4042,In_4043,In_4044,In_4045,In_4046,In_4047,In_4048,In_4049,In_4050,In_4051,In_4052,In_4053,In_4054,In_4055,In_4056,In_4057,In_4058,In_4059,In_4060,In_4061,In_4062,In_4063,In_4064,In_4065,In_4066,In_4067,In_4068,In_4069,In_4070,In_4071,In_4072,In_4073,In_4074,In_4075,In_4076,In_4077,In_4078,In_4079,In_4080,In_4081,In_4082,In_4083,In_4084,In_4085,In_4086,In_4087,In_4088,In_4089,In_4090,In_4091,In_4092,In_4093,In_4094,In_4095,In_4096,In_4097,In_4098,In_4099,In_4100,In_4101,In_4102,In_4103,In_4104,In_4105,In_4106,In_4107,In_4108,In_4109,In_4110,In_4111,In_4112,In_4113,In_4114,In_4115,In_4116,In_4117,In_4118,In_4119,In_4120,In_4121,In_4122,In_4123,In_4124,In_4125,In_4126,In_4127,In_4128,In_4129,In_4130,In_4131,In_4132,In_4133,In_4134,In_4135,In_4136,In_4137,In_4138,In_4139,In_4140,In_4141,In_4142,In_4143,In_4144,In_4145,In_4146,In_4147,In_4148,In_4149,In_4150,In_4151,In_4152,In_4153,In_4154,In_4155,In_4156,In_4157,In_4158,In_4159,In_4160,In_4161,In_4162,In_4163,In_4164,In_4165,In_4166,In_4167,In_4168,In_4169,In_4170,In_4171,In_4172,In_4173,In_4174,In_4175,In_4176,In_4177,In_4178,In_4179,In_4180,In_4181,In_4182,In_4183,In_4184,In_4185,In_4186,In_4187,In_4188,In_4189,In_4190,In_4191,In_4192,In_4193,In_4194,In_4195,In_4196,In_4197,In_4198,In_4199,In_4200,In_4201,In_4202,In_4203,In_4204,In_4205,In_4206,In_4207,In_4208,In_4209,In_4210,In_4211,In_4212,In_4213,In_4214,In_4215,In_4216,In_4217,In_4218,In_4219,In_4220,In_4221,In_4222,In_4223,In_4224,In_4225,In_4226,In_4227,In_4228,In_4229,In_4230,In_4231,In_4232,In_4233,In_4234,In_4235,In_4236,In_4237,In_4238,In_4239,In_4240,In_4241,In_4242,In_4243,In_4244,In_4245,In_4246,In_4247,In_4248,In_4249,In_4250,In_4251,In_4252,In_4253,In_4254,In_4255,In_4256,In_4257,In_4258,In_4259,In_4260,In_4261,In_4262,In_4263,In_4264,In_4265,In_4266,In_4267,In_4268,In_4269,In_4270,In_4271,In_4272,In_4273,In_4274,In_4275,In_4276,In_4277,In_4278,In_4279,In_4280,In_4281,In_4282,In_4283,In_4284,In_4285,In_4286,In_4287,In_4288,In_4289,In_4290,In_4291,In_4292,In_4293,In_4294,In_4295,In_4296,In_4297,In_4298,In_4299,In_4300,In_4301,In_4302,In_4303,In_4304,In_4305,In_4306,In_4307,In_4308,In_4309,In_4310,In_4311,In_4312,In_4313,In_4314,In_4315,In_4316,In_4317,In_4318,In_4319,In_4320,In_4321,In_4322,In_4323,In_4324,In_4325,In_4326,In_4327,In_4328,In_4329,In_4330,In_4331,In_4332,In_4333,In_4334,In_4335,In_4336,In_4337,In_4338,In_4339,In_4340,In_4341,In_4342,In_4343,In_4344,In_4345,In_4346,In_4347,In_4348,In_4349,In_4350,In_4351,In_4352,In_4353,In_4354,In_4355,In_4356,In_4357,In_4358,In_4359,In_4360,In_4361,In_4362,In_4363,In_4364,In_4365,In_4366,In_4367,In_4368,In_4369,In_4370,In_4371,In_4372,In_4373,In_4374,In_4375,In_4376,In_4377,In_4378,In_4379,In_4380,In_4381,In_4382,In_4383,In_4384,In_4385,In_4386,In_4387,In_4388,In_4389,In_4390,In_4391,In_4392,In_4393,In_4394,In_4395,In_4396,In_4397,In_4398,In_4399,In_4400,In_4401,In_4402,In_4403,In_4404,In_4405,In_4406,In_4407,In_4408,In_4409,In_4410,In_4411,In_4412,In_4413,In_4414,In_4415,In_4416,In_4417,In_4418,In_4419,In_4420,In_4421,In_4422,In_4423,In_4424,In_4425,In_4426,In_4427,In_4428,In_4429,In_4430,In_4431,In_4432,In_4433,In_4434,In_4435,In_4436,In_4437,In_4438,In_4439,In_4440,In_4441,In_4442,In_4443,In_4444,In_4445,In_4446,In_4447,In_4448,In_4449,In_4450,In_4451,In_4452,In_4453,In_4454,In_4455,In_4456,In_4457,In_4458,In_4459,In_4460,In_4461,In_4462,In_4463,In_4464,In_4465,In_4466,In_4467,In_4468,In_4469,In_4470,In_4471,In_4472,In_4473,In_4474,In_4475,In_4476,In_4477,In_4478,In_4479,In_4480,In_4481,In_4482,In_4483,In_4484,In_4485,In_4486,In_4487,In_4488,In_4489,In_4490,In_4491,In_4492,In_4493,In_4494,In_4495,In_4496,In_4497,In_4498,In_4499,In_4500,In_4501,In_4502,In_4503,In_4504,In_4505,In_4506,In_4507,In_4508,In_4509,In_4510,In_4511,In_4512,In_4513,In_4514,In_4515,In_4516,In_4517,In_4518,In_4519,In_4520,In_4521,In_4522,In_4523,In_4524,In_4525,In_4526,In_4527,In_4528,In_4529,In_4530,In_4531,In_4532,In_4533,In_4534,In_4535,In_4536,In_4537,In_4538,In_4539,In_4540,In_4541,In_4542,In_4543,In_4544,In_4545,In_4546,In_4547,In_4548,In_4549,In_4550,In_4551,In_4552,In_4553,In_4554,In_4555,In_4556,In_4557,In_4558,In_4559,In_4560,In_4561,In_4562,In_4563,In_4564,In_4565,In_4566,In_4567,In_4568,In_4569,In_4570,In_4571,In_4572,In_4573,In_4574,In_4575,In_4576,In_4577,In_4578,In_4579,In_4580,In_4581,In_4582,In_4583,In_4584,In_4585,In_4586,In_4587,In_4588,In_4589,In_4590,In_4591,In_4592,In_4593,In_4594,In_4595,In_4596,In_4597,In_4598,In_4599,In_4600,In_4601,In_4602,In_4603,In_4604,In_4605,In_4606,In_4607,In_4608,In_4609,In_4610,In_4611,In_4612,In_4613,In_4614,In_4615,In_4616,In_4617,In_4618,In_4619,In_4620,In_4621,In_4622,In_4623,In_4624,In_4625,In_4626,In_4627,In_4628,In_4629,In_4630,In_4631,In_4632,In_4633,In_4634,In_4635,In_4636,In_4637,In_4638,In_4639,In_4640,In_4641,In_4642,In_4643,In_4644,In_4645,In_4646,In_4647,In_4648,In_4649,In_4650,In_4651,In_4652,In_4653,In_4654,In_4655,In_4656,In_4657,In_4658,In_4659,In_4660,In_4661,In_4662,In_4663,In_4664,In_4665,In_4666,In_4667,In_4668,In_4669,In_4670,In_4671,In_4672,In_4673,In_4674,In_4675,In_4676,In_4677,In_4678,In_4679,In_4680,In_4681,In_4682,In_4683,In_4684,In_4685,In_4686,In_4687,In_4688,In_4689,In_4690,In_4691,In_4692,In_4693,In_4694,In_4695,In_4696,In_4697,In_4698,In_4699,In_4700,In_4701,In_4702,In_4703,In_4704,In_4705,In_4706,In_4707,In_4708,In_4709,In_4710,In_4711,In_4712,In_4713,In_4714,In_4715,In_4716,In_4717,In_4718,In_4719,In_4720,In_4721,In_4722,In_4723,In_4724,In_4725,In_4726,In_4727,In_4728,In_4729,In_4730,In_4731,In_4732,In_4733,In_4734,In_4735,In_4736,In_4737,In_4738,In_4739,In_4740,In_4741,In_4742,In_4743,In_4744,In_4745,In_4746,In_4747,In_4748,In_4749,In_4750,In_4751,In_4752,In_4753,In_4754,In_4755,In_4756,In_4757,In_4758,In_4759,In_4760,In_4761,In_4762,In_4763,In_4764,In_4765,In_4766,In_4767,In_4768,In_4769,In_4770,In_4771,In_4772,In_4773,In_4774,In_4775,In_4776,In_4777,In_4778,In_4779,In_4780,In_4781,In_4782,In_4783,In_4784,In_4785,In_4786,In_4787,In_4788,In_4789,In_4790,In_4791,In_4792,In_4793,In_4794,In_4795,In_4796,In_4797,In_4798,In_4799,In_4800,In_4801,In_4802,In_4803,In_4804,In_4805,In_4806,In_4807,In_4808,In_4809,In_4810,In_4811,In_4812,In_4813,In_4814,In_4815,In_4816,In_4817,In_4818,In_4819,In_4820,In_4821,In_4822,In_4823,In_4824,In_4825,In_4826,In_4827,In_4828,In_4829,In_4830,In_4831,In_4832,In_4833,In_4834,In_4835,In_4836,In_4837,In_4838,In_4839,In_4840,In_4841,In_4842,In_4843,In_4844,In_4845,In_4846,In_4847,In_4848,In_4849,In_4850,In_4851,In_4852,In_4853,In_4854,In_4855,In_4856,In_4857,In_4858,In_4859,In_4860,In_4861,In_4862,In_4863,In_4864,In_4865,In_4866,In_4867,In_4868,In_4869,In_4870,In_4871,In_4872,In_4873,In_4874,In_4875,In_4876,In_4877,In_4878,In_4879,In_4880,In_4881,In_4882,In_4883,In_4884,In_4885,In_4886,In_4887,In_4888,In_4889,In_4890,In_4891,In_4892,In_4893,In_4894,In_4895,In_4896,In_4897,In_4898,In_4899,In_4900,In_4901,In_4902,In_4903,In_4904,In_4905,In_4906,In_4907,In_4908,In_4909,In_4910,In_4911,In_4912,In_4913,In_4914,In_4915,In_4916,In_4917,In_4918,In_4919,In_4920,In_4921,In_4922,In_4923,In_4924,In_4925,In_4926,In_4927,In_4928,In_4929,In_4930,In_4931,In_4932,In_4933,In_4934,In_4935,In_4936,In_4937,In_4938,In_4939,In_4940,In_4941,In_4942,In_4943,In_4944,In_4945,In_4946,In_4947,In_4948,In_4949,In_4950,In_4951,In_4952,In_4953,In_4954,In_4955,In_4956,In_4957,In_4958,In_4959,In_4960,In_4961,In_4962,In_4963,In_4964,In_4965,In_4966,In_4967,In_4968,In_4969,In_4970,In_4971,In_4972,In_4973,In_4974,In_4975,In_4976,In_4977,In_4978,In_4979,In_4980,In_4981,In_4982,In_4983,In_4984,In_4985,In_4986,In_4987,In_4988,In_4989,In_4990,In_4991,In_4992,In_4993,In_4994,In_4995,In_4996,In_4997,In_4998,In_4999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499,O_3500,O_3501,O_3502,O_3503,O_3504,O_3505,O_3506,O_3507,O_3508,O_3509,O_3510,O_3511,O_3512,O_3513,O_3514,O_3515,O_3516,O_3517,O_3518,O_3519,O_3520,O_3521,O_3522,O_3523,O_3524,O_3525,O_3526,O_3527,O_3528,O_3529,O_3530,O_3531,O_3532,O_3533,O_3534,O_3535,O_3536,O_3537,O_3538,O_3539,O_3540,O_3541,O_3542,O_3543,O_3544,O_3545,O_3546,O_3547,O_3548,O_3549,O_3550,O_3551,O_3552,O_3553,O_3554,O_3555,O_3556,O_3557,O_3558,O_3559,O_3560,O_3561,O_3562,O_3563,O_3564,O_3565,O_3566,O_3567,O_3568,O_3569,O_3570,O_3571,O_3572,O_3573,O_3574,O_3575,O_3576,O_3577,O_3578,O_3579,O_3580,O_3581,O_3582,O_3583,O_3584,O_3585,O_3586,O_3587,O_3588,O_3589,O_3590,O_3591,O_3592,O_3593,O_3594,O_3595,O_3596,O_3597,O_3598,O_3599,O_3600,O_3601,O_3602,O_3603,O_3604,O_3605,O_3606,O_3607,O_3608,O_3609,O_3610,O_3611,O_3612,O_3613,O_3614,O_3615,O_3616,O_3617,O_3618,O_3619,O_3620,O_3621,O_3622,O_3623,O_3624,O_3625,O_3626,O_3627,O_3628,O_3629,O_3630,O_3631,O_3632,O_3633,O_3634,O_3635,O_3636,O_3637,O_3638,O_3639,O_3640,O_3641,O_3642,O_3643,O_3644,O_3645,O_3646,O_3647,O_3648,O_3649,O_3650,O_3651,O_3652,O_3653,O_3654,O_3655,O_3656,O_3657,O_3658,O_3659,O_3660,O_3661,O_3662,O_3663,O_3664,O_3665,O_3666,O_3667,O_3668,O_3669,O_3670,O_3671,O_3672,O_3673,O_3674,O_3675,O_3676,O_3677,O_3678,O_3679,O_3680,O_3681,O_3682,O_3683,O_3684,O_3685,O_3686,O_3687,O_3688,O_3689,O_3690,O_3691,O_3692,O_3693,O_3694,O_3695,O_3696,O_3697,O_3698,O_3699,O_3700,O_3701,O_3702,O_3703,O_3704,O_3705,O_3706,O_3707,O_3708,O_3709,O_3710,O_3711,O_3712,O_3713,O_3714,O_3715,O_3716,O_3717,O_3718,O_3719,O_3720,O_3721,O_3722,O_3723,O_3724,O_3725,O_3726,O_3727,O_3728,O_3729,O_3730,O_3731,O_3732,O_3733,O_3734,O_3735,O_3736,O_3737,O_3738,O_3739,O_3740,O_3741,O_3742,O_3743,O_3744,O_3745,O_3746,O_3747,O_3748,O_3749,O_3750,O_3751,O_3752,O_3753,O_3754,O_3755,O_3756,O_3757,O_3758,O_3759,O_3760,O_3761,O_3762,O_3763,O_3764,O_3765,O_3766,O_3767,O_3768,O_3769,O_3770,O_3771,O_3772,O_3773,O_3774,O_3775,O_3776,O_3777,O_3778,O_3779,O_3780,O_3781,O_3782,O_3783,O_3784,O_3785,O_3786,O_3787,O_3788,O_3789,O_3790,O_3791,O_3792,O_3793,O_3794,O_3795,O_3796,O_3797,O_3798,O_3799,O_3800,O_3801,O_3802,O_3803,O_3804,O_3805,O_3806,O_3807,O_3808,O_3809,O_3810,O_3811,O_3812,O_3813,O_3814,O_3815,O_3816,O_3817,O_3818,O_3819,O_3820,O_3821,O_3822,O_3823,O_3824,O_3825,O_3826,O_3827,O_3828,O_3829,O_3830,O_3831,O_3832,O_3833,O_3834,O_3835,O_3836,O_3837,O_3838,O_3839,O_3840,O_3841,O_3842,O_3843,O_3844,O_3845,O_3846,O_3847,O_3848,O_3849,O_3850,O_3851,O_3852,O_3853,O_3854,O_3855,O_3856,O_3857,O_3858,O_3859,O_3860,O_3861,O_3862,O_3863,O_3864,O_3865,O_3866,O_3867,O_3868,O_3869,O_3870,O_3871,O_3872,O_3873,O_3874,O_3875,O_3876,O_3877,O_3878,O_3879,O_3880,O_3881,O_3882,O_3883,O_3884,O_3885,O_3886,O_3887,O_3888,O_3889,O_3890,O_3891,O_3892,O_3893,O_3894,O_3895,O_3896,O_3897,O_3898,O_3899,O_3900,O_3901,O_3902,O_3903,O_3904,O_3905,O_3906,O_3907,O_3908,O_3909,O_3910,O_3911,O_3912,O_3913,O_3914,O_3915,O_3916,O_3917,O_3918,O_3919,O_3920,O_3921,O_3922,O_3923,O_3924,O_3925,O_3926,O_3927,O_3928,O_3929,O_3930,O_3931,O_3932,O_3933,O_3934,O_3935,O_3936,O_3937,O_3938,O_3939,O_3940,O_3941,O_3942,O_3943,O_3944,O_3945,O_3946,O_3947,O_3948,O_3949,O_3950,O_3951,O_3952,O_3953,O_3954,O_3955,O_3956,O_3957,O_3958,O_3959,O_3960,O_3961,O_3962,O_3963,O_3964,O_3965,O_3966,O_3967,O_3968,O_3969,O_3970,O_3971,O_3972,O_3973,O_3974,O_3975,O_3976,O_3977,O_3978,O_3979,O_3980,O_3981,O_3982,O_3983,O_3984,O_3985,O_3986,O_3987,O_3988,O_3989,O_3990,O_3991,O_3992,O_3993,O_3994,O_3995,O_3996,O_3997,O_3998,O_3999,O_4000,O_4001,O_4002,O_4003,O_4004,O_4005,O_4006,O_4007,O_4008,O_4009,O_4010,O_4011,O_4012,O_4013,O_4014,O_4015,O_4016,O_4017,O_4018,O_4019,O_4020,O_4021,O_4022,O_4023,O_4024,O_4025,O_4026,O_4027,O_4028,O_4029,O_4030,O_4031,O_4032,O_4033,O_4034,O_4035,O_4036,O_4037,O_4038,O_4039,O_4040,O_4041,O_4042,O_4043,O_4044,O_4045,O_4046,O_4047,O_4048,O_4049,O_4050,O_4051,O_4052,O_4053,O_4054,O_4055,O_4056,O_4057,O_4058,O_4059,O_4060,O_4061,O_4062,O_4063,O_4064,O_4065,O_4066,O_4067,O_4068,O_4069,O_4070,O_4071,O_4072,O_4073,O_4074,O_4075,O_4076,O_4077,O_4078,O_4079,O_4080,O_4081,O_4082,O_4083,O_4084,O_4085,O_4086,O_4087,O_4088,O_4089,O_4090,O_4091,O_4092,O_4093,O_4094,O_4095,O_4096,O_4097,O_4098,O_4099,O_4100,O_4101,O_4102,O_4103,O_4104,O_4105,O_4106,O_4107,O_4108,O_4109,O_4110,O_4111,O_4112,O_4113,O_4114,O_4115,O_4116,O_4117,O_4118,O_4119,O_4120,O_4121,O_4122,O_4123,O_4124,O_4125,O_4126,O_4127,O_4128,O_4129,O_4130,O_4131,O_4132,O_4133,O_4134,O_4135,O_4136,O_4137,O_4138,O_4139,O_4140,O_4141,O_4142,O_4143,O_4144,O_4145,O_4146,O_4147,O_4148,O_4149,O_4150,O_4151,O_4152,O_4153,O_4154,O_4155,O_4156,O_4157,O_4158,O_4159,O_4160,O_4161,O_4162,O_4163,O_4164,O_4165,O_4166,O_4167,O_4168,O_4169,O_4170,O_4171,O_4172,O_4173,O_4174,O_4175,O_4176,O_4177,O_4178,O_4179,O_4180,O_4181,O_4182,O_4183,O_4184,O_4185,O_4186,O_4187,O_4188,O_4189,O_4190,O_4191,O_4192,O_4193,O_4194,O_4195,O_4196,O_4197,O_4198,O_4199,O_4200,O_4201,O_4202,O_4203,O_4204,O_4205,O_4206,O_4207,O_4208,O_4209,O_4210,O_4211,O_4212,O_4213,O_4214,O_4215,O_4216,O_4217,O_4218,O_4219,O_4220,O_4221,O_4222,O_4223,O_4224,O_4225,O_4226,O_4227,O_4228,O_4229,O_4230,O_4231,O_4232,O_4233,O_4234,O_4235,O_4236,O_4237,O_4238,O_4239,O_4240,O_4241,O_4242,O_4243,O_4244,O_4245,O_4246,O_4247,O_4248,O_4249,O_4250,O_4251,O_4252,O_4253,O_4254,O_4255,O_4256,O_4257,O_4258,O_4259,O_4260,O_4261,O_4262,O_4263,O_4264,O_4265,O_4266,O_4267,O_4268,O_4269,O_4270,O_4271,O_4272,O_4273,O_4274,O_4275,O_4276,O_4277,O_4278,O_4279,O_4280,O_4281,O_4282,O_4283,O_4284,O_4285,O_4286,O_4287,O_4288,O_4289,O_4290,O_4291,O_4292,O_4293,O_4294,O_4295,O_4296,O_4297,O_4298,O_4299,O_4300,O_4301,O_4302,O_4303,O_4304,O_4305,O_4306,O_4307,O_4308,O_4309,O_4310,O_4311,O_4312,O_4313,O_4314,O_4315,O_4316,O_4317,O_4318,O_4319,O_4320,O_4321,O_4322,O_4323,O_4324,O_4325,O_4326,O_4327,O_4328,O_4329,O_4330,O_4331,O_4332,O_4333,O_4334,O_4335,O_4336,O_4337,O_4338,O_4339,O_4340,O_4341,O_4342,O_4343,O_4344,O_4345,O_4346,O_4347,O_4348,O_4349,O_4350,O_4351,O_4352,O_4353,O_4354,O_4355,O_4356,O_4357,O_4358,O_4359,O_4360,O_4361,O_4362,O_4363,O_4364,O_4365,O_4366,O_4367,O_4368,O_4369,O_4370,O_4371,O_4372,O_4373,O_4374,O_4375,O_4376,O_4377,O_4378,O_4379,O_4380,O_4381,O_4382,O_4383,O_4384,O_4385,O_4386,O_4387,O_4388,O_4389,O_4390,O_4391,O_4392,O_4393,O_4394,O_4395,O_4396,O_4397,O_4398,O_4399,O_4400,O_4401,O_4402,O_4403,O_4404,O_4405,O_4406,O_4407,O_4408,O_4409,O_4410,O_4411,O_4412,O_4413,O_4414,O_4415,O_4416,O_4417,O_4418,O_4419,O_4420,O_4421,O_4422,O_4423,O_4424,O_4425,O_4426,O_4427,O_4428,O_4429,O_4430,O_4431,O_4432,O_4433,O_4434,O_4435,O_4436,O_4437,O_4438,O_4439,O_4440,O_4441,O_4442,O_4443,O_4444,O_4445,O_4446,O_4447,O_4448,O_4449,O_4450,O_4451,O_4452,O_4453,O_4454,O_4455,O_4456,O_4457,O_4458,O_4459,O_4460,O_4461,O_4462,O_4463,O_4464,O_4465,O_4466,O_4467,O_4468,O_4469,O_4470,O_4471,O_4472,O_4473,O_4474,O_4475,O_4476,O_4477,O_4478,O_4479,O_4480,O_4481,O_4482,O_4483,O_4484,O_4485,O_4486,O_4487,O_4488,O_4489,O_4490,O_4491,O_4492,O_4493,O_4494,O_4495,O_4496,O_4497,O_4498,O_4499,O_4500,O_4501,O_4502,O_4503,O_4504,O_4505,O_4506,O_4507,O_4508,O_4509,O_4510,O_4511,O_4512,O_4513,O_4514,O_4515,O_4516,O_4517,O_4518,O_4519,O_4520,O_4521,O_4522,O_4523,O_4524,O_4525,O_4526,O_4527,O_4528,O_4529,O_4530,O_4531,O_4532,O_4533,O_4534,O_4535,O_4536,O_4537,O_4538,O_4539,O_4540,O_4541,O_4542,O_4543,O_4544,O_4545,O_4546,O_4547,O_4548,O_4549,O_4550,O_4551,O_4552,O_4553,O_4554,O_4555,O_4556,O_4557,O_4558,O_4559,O_4560,O_4561,O_4562,O_4563,O_4564,O_4565,O_4566,O_4567,O_4568,O_4569,O_4570,O_4571,O_4572,O_4573,O_4574,O_4575,O_4576,O_4577,O_4578,O_4579,O_4580,O_4581,O_4582,O_4583,O_4584,O_4585,O_4586,O_4587,O_4588,O_4589,O_4590,O_4591,O_4592,O_4593,O_4594,O_4595,O_4596,O_4597,O_4598,O_4599,O_4600,O_4601,O_4602,O_4603,O_4604,O_4605,O_4606,O_4607,O_4608,O_4609,O_4610,O_4611,O_4612,O_4613,O_4614,O_4615,O_4616,O_4617,O_4618,O_4619,O_4620,O_4621,O_4622,O_4623,O_4624,O_4625,O_4626,O_4627,O_4628,O_4629,O_4630,O_4631,O_4632,O_4633,O_4634,O_4635,O_4636,O_4637,O_4638,O_4639,O_4640,O_4641,O_4642,O_4643,O_4644,O_4645,O_4646,O_4647,O_4648,O_4649,O_4650,O_4651,O_4652,O_4653,O_4654,O_4655,O_4656,O_4657,O_4658,O_4659,O_4660,O_4661,O_4662,O_4663,O_4664,O_4665,O_4666,O_4667,O_4668,O_4669,O_4670,O_4671,O_4672,O_4673,O_4674,O_4675,O_4676,O_4677,O_4678,O_4679,O_4680,O_4681,O_4682,O_4683,O_4684,O_4685,O_4686,O_4687,O_4688,O_4689,O_4690,O_4691,O_4692,O_4693,O_4694,O_4695,O_4696,O_4697,O_4698,O_4699,O_4700,O_4701,O_4702,O_4703,O_4704,O_4705,O_4706,O_4707,O_4708,O_4709,O_4710,O_4711,O_4712,O_4713,O_4714,O_4715,O_4716,O_4717,O_4718,O_4719,O_4720,O_4721,O_4722,O_4723,O_4724,O_4725,O_4726,O_4727,O_4728,O_4729,O_4730,O_4731,O_4732,O_4733,O_4734,O_4735,O_4736,O_4737,O_4738,O_4739,O_4740,O_4741,O_4742,O_4743,O_4744,O_4745,O_4746,O_4747,O_4748,O_4749,O_4750,O_4751,O_4752,O_4753,O_4754,O_4755,O_4756,O_4757,O_4758,O_4759,O_4760,O_4761,O_4762,O_4763,O_4764,O_4765,O_4766,O_4767,O_4768,O_4769,O_4770,O_4771,O_4772,O_4773,O_4774,O_4775,O_4776,O_4777,O_4778,O_4779,O_4780,O_4781,O_4782,O_4783,O_4784,O_4785,O_4786,O_4787,O_4788,O_4789,O_4790,O_4791,O_4792,O_4793,O_4794,O_4795,O_4796,O_4797,O_4798,O_4799,O_4800,O_4801,O_4802,O_4803,O_4804,O_4805,O_4806,O_4807,O_4808,O_4809,O_4810,O_4811,O_4812,O_4813,O_4814,O_4815,O_4816,O_4817,O_4818,O_4819,O_4820,O_4821,O_4822,O_4823,O_4824,O_4825,O_4826,O_4827,O_4828,O_4829,O_4830,O_4831,O_4832,O_4833,O_4834,O_4835,O_4836,O_4837,O_4838,O_4839,O_4840,O_4841,O_4842,O_4843,O_4844,O_4845,O_4846,O_4847,O_4848,O_4849,O_4850,O_4851,O_4852,O_4853,O_4854,O_4855,O_4856,O_4857,O_4858,O_4859,O_4860,O_4861,O_4862,O_4863,O_4864,O_4865,O_4866,O_4867,O_4868,O_4869,O_4870,O_4871,O_4872,O_4873,O_4874,O_4875,O_4876,O_4877,O_4878,O_4879,O_4880,O_4881,O_4882,O_4883,O_4884,O_4885,O_4886,O_4887,O_4888,O_4889,O_4890,O_4891,O_4892,O_4893,O_4894,O_4895,O_4896,O_4897,O_4898,O_4899,O_4900,O_4901,O_4902,O_4903,O_4904,O_4905,O_4906,O_4907,O_4908,O_4909,O_4910,O_4911,O_4912,O_4913,O_4914,O_4915,O_4916,O_4917,O_4918,O_4919,O_4920,O_4921,O_4922,O_4923,O_4924,O_4925,O_4926,O_4927,O_4928,O_4929,O_4930,O_4931,O_4932,O_4933,O_4934,O_4935,O_4936,O_4937,O_4938,O_4939,O_4940,O_4941,O_4942,O_4943,O_4944,O_4945,O_4946,O_4947,O_4948,O_4949,O_4950,O_4951,O_4952,O_4953,O_4954,O_4955,O_4956,O_4957,O_4958,O_4959,O_4960,O_4961,O_4962,O_4963,O_4964,O_4965,O_4966,O_4967,O_4968,O_4969,O_4970,O_4971,O_4972,O_4973,O_4974,O_4975,O_4976,O_4977,O_4978,O_4979,O_4980,O_4981,O_4982,O_4983,O_4984,O_4985,O_4986,O_4987,O_4988,O_4989,O_4990,O_4991,O_4992,O_4993,O_4994,O_4995,O_4996,O_4997,O_4998,O_4999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999,N_25000,N_25001,N_25002,N_25003,N_25004,N_25005,N_25006,N_25007,N_25008,N_25009,N_25010,N_25011,N_25012,N_25013,N_25014,N_25015,N_25016,N_25017,N_25018,N_25019,N_25020,N_25021,N_25022,N_25023,N_25024,N_25025,N_25026,N_25027,N_25028,N_25029,N_25030,N_25031,N_25032,N_25033,N_25034,N_25035,N_25036,N_25037,N_25038,N_25039,N_25040,N_25041,N_25042,N_25043,N_25044,N_25045,N_25046,N_25047,N_25048,N_25049,N_25050,N_25051,N_25052,N_25053,N_25054,N_25055,N_25056,N_25057,N_25058,N_25059,N_25060,N_25061,N_25062,N_25063,N_25064,N_25065,N_25066,N_25067,N_25068,N_25069,N_25070,N_25071,N_25072,N_25073,N_25074,N_25075,N_25076,N_25077,N_25078,N_25079,N_25080,N_25081,N_25082,N_25083,N_25084,N_25085,N_25086,N_25087,N_25088,N_25089,N_25090,N_25091,N_25092,N_25093,N_25094,N_25095,N_25096,N_25097,N_25098,N_25099,N_25100,N_25101,N_25102,N_25103,N_25104,N_25105,N_25106,N_25107,N_25108,N_25109,N_25110,N_25111,N_25112,N_25113,N_25114,N_25115,N_25116,N_25117,N_25118,N_25119,N_25120,N_25121,N_25122,N_25123,N_25124,N_25125,N_25126,N_25127,N_25128,N_25129,N_25130,N_25131,N_25132,N_25133,N_25134,N_25135,N_25136,N_25137,N_25138,N_25139,N_25140,N_25141,N_25142,N_25143,N_25144,N_25145,N_25146,N_25147,N_25148,N_25149,N_25150,N_25151,N_25152,N_25153,N_25154,N_25155,N_25156,N_25157,N_25158,N_25159,N_25160,N_25161,N_25162,N_25163,N_25164,N_25165,N_25166,N_25167,N_25168,N_25169,N_25170,N_25171,N_25172,N_25173,N_25174,N_25175,N_25176,N_25177,N_25178,N_25179,N_25180,N_25181,N_25182,N_25183,N_25184,N_25185,N_25186,N_25187,N_25188,N_25189,N_25190,N_25191,N_25192,N_25193,N_25194,N_25195,N_25196,N_25197,N_25198,N_25199,N_25200,N_25201,N_25202,N_25203,N_25204,N_25205,N_25206,N_25207,N_25208,N_25209,N_25210,N_25211,N_25212,N_25213,N_25214,N_25215,N_25216,N_25217,N_25218,N_25219,N_25220,N_25221,N_25222,N_25223,N_25224,N_25225,N_25226,N_25227,N_25228,N_25229,N_25230,N_25231,N_25232,N_25233,N_25234,N_25235,N_25236,N_25237,N_25238,N_25239,N_25240,N_25241,N_25242,N_25243,N_25244,N_25245,N_25246,N_25247,N_25248,N_25249,N_25250,N_25251,N_25252,N_25253,N_25254,N_25255,N_25256,N_25257,N_25258,N_25259,N_25260,N_25261,N_25262,N_25263,N_25264,N_25265,N_25266,N_25267,N_25268,N_25269,N_25270,N_25271,N_25272,N_25273,N_25274,N_25275,N_25276,N_25277,N_25278,N_25279,N_25280,N_25281,N_25282,N_25283,N_25284,N_25285,N_25286,N_25287,N_25288,N_25289,N_25290,N_25291,N_25292,N_25293,N_25294,N_25295,N_25296,N_25297,N_25298,N_25299,N_25300,N_25301,N_25302,N_25303,N_25304,N_25305,N_25306,N_25307,N_25308,N_25309,N_25310,N_25311,N_25312,N_25313,N_25314,N_25315,N_25316,N_25317,N_25318,N_25319,N_25320,N_25321,N_25322,N_25323,N_25324,N_25325,N_25326,N_25327,N_25328,N_25329,N_25330,N_25331,N_25332,N_25333,N_25334,N_25335,N_25336,N_25337,N_25338,N_25339,N_25340,N_25341,N_25342,N_25343,N_25344,N_25345,N_25346,N_25347,N_25348,N_25349,N_25350,N_25351,N_25352,N_25353,N_25354,N_25355,N_25356,N_25357,N_25358,N_25359,N_25360,N_25361,N_25362,N_25363,N_25364,N_25365,N_25366,N_25367,N_25368,N_25369,N_25370,N_25371,N_25372,N_25373,N_25374,N_25375,N_25376,N_25377,N_25378,N_25379,N_25380,N_25381,N_25382,N_25383,N_25384,N_25385,N_25386,N_25387,N_25388,N_25389,N_25390,N_25391,N_25392,N_25393,N_25394,N_25395,N_25396,N_25397,N_25398,N_25399,N_25400,N_25401,N_25402,N_25403,N_25404,N_25405,N_25406,N_25407,N_25408,N_25409,N_25410,N_25411,N_25412,N_25413,N_25414,N_25415,N_25416,N_25417,N_25418,N_25419,N_25420,N_25421,N_25422,N_25423,N_25424,N_25425,N_25426,N_25427,N_25428,N_25429,N_25430,N_25431,N_25432,N_25433,N_25434,N_25435,N_25436,N_25437,N_25438,N_25439,N_25440,N_25441,N_25442,N_25443,N_25444,N_25445,N_25446,N_25447,N_25448,N_25449,N_25450,N_25451,N_25452,N_25453,N_25454,N_25455,N_25456,N_25457,N_25458,N_25459,N_25460,N_25461,N_25462,N_25463,N_25464,N_25465,N_25466,N_25467,N_25468,N_25469,N_25470,N_25471,N_25472,N_25473,N_25474,N_25475,N_25476,N_25477,N_25478,N_25479,N_25480,N_25481,N_25482,N_25483,N_25484,N_25485,N_25486,N_25487,N_25488,N_25489,N_25490,N_25491,N_25492,N_25493,N_25494,N_25495,N_25496,N_25497,N_25498,N_25499,N_25500,N_25501,N_25502,N_25503,N_25504,N_25505,N_25506,N_25507,N_25508,N_25509,N_25510,N_25511,N_25512,N_25513,N_25514,N_25515,N_25516,N_25517,N_25518,N_25519,N_25520,N_25521,N_25522,N_25523,N_25524,N_25525,N_25526,N_25527,N_25528,N_25529,N_25530,N_25531,N_25532,N_25533,N_25534,N_25535,N_25536,N_25537,N_25538,N_25539,N_25540,N_25541,N_25542,N_25543,N_25544,N_25545,N_25546,N_25547,N_25548,N_25549,N_25550,N_25551,N_25552,N_25553,N_25554,N_25555,N_25556,N_25557,N_25558,N_25559,N_25560,N_25561,N_25562,N_25563,N_25564,N_25565,N_25566,N_25567,N_25568,N_25569,N_25570,N_25571,N_25572,N_25573,N_25574,N_25575,N_25576,N_25577,N_25578,N_25579,N_25580,N_25581,N_25582,N_25583,N_25584,N_25585,N_25586,N_25587,N_25588,N_25589,N_25590,N_25591,N_25592,N_25593,N_25594,N_25595,N_25596,N_25597,N_25598,N_25599,N_25600,N_25601,N_25602,N_25603,N_25604,N_25605,N_25606,N_25607,N_25608,N_25609,N_25610,N_25611,N_25612,N_25613,N_25614,N_25615,N_25616,N_25617,N_25618,N_25619,N_25620,N_25621,N_25622,N_25623,N_25624,N_25625,N_25626,N_25627,N_25628,N_25629,N_25630,N_25631,N_25632,N_25633,N_25634,N_25635,N_25636,N_25637,N_25638,N_25639,N_25640,N_25641,N_25642,N_25643,N_25644,N_25645,N_25646,N_25647,N_25648,N_25649,N_25650,N_25651,N_25652,N_25653,N_25654,N_25655,N_25656,N_25657,N_25658,N_25659,N_25660,N_25661,N_25662,N_25663,N_25664,N_25665,N_25666,N_25667,N_25668,N_25669,N_25670,N_25671,N_25672,N_25673,N_25674,N_25675,N_25676,N_25677,N_25678,N_25679,N_25680,N_25681,N_25682,N_25683,N_25684,N_25685,N_25686,N_25687,N_25688,N_25689,N_25690,N_25691,N_25692,N_25693,N_25694,N_25695,N_25696,N_25697,N_25698,N_25699,N_25700,N_25701,N_25702,N_25703,N_25704,N_25705,N_25706,N_25707,N_25708,N_25709,N_25710,N_25711,N_25712,N_25713,N_25714,N_25715,N_25716,N_25717,N_25718,N_25719,N_25720,N_25721,N_25722,N_25723,N_25724,N_25725,N_25726,N_25727,N_25728,N_25729,N_25730,N_25731,N_25732,N_25733,N_25734,N_25735,N_25736,N_25737,N_25738,N_25739,N_25740,N_25741,N_25742,N_25743,N_25744,N_25745,N_25746,N_25747,N_25748,N_25749,N_25750,N_25751,N_25752,N_25753,N_25754,N_25755,N_25756,N_25757,N_25758,N_25759,N_25760,N_25761,N_25762,N_25763,N_25764,N_25765,N_25766,N_25767,N_25768,N_25769,N_25770,N_25771,N_25772,N_25773,N_25774,N_25775,N_25776,N_25777,N_25778,N_25779,N_25780,N_25781,N_25782,N_25783,N_25784,N_25785,N_25786,N_25787,N_25788,N_25789,N_25790,N_25791,N_25792,N_25793,N_25794,N_25795,N_25796,N_25797,N_25798,N_25799,N_25800,N_25801,N_25802,N_25803,N_25804,N_25805,N_25806,N_25807,N_25808,N_25809,N_25810,N_25811,N_25812,N_25813,N_25814,N_25815,N_25816,N_25817,N_25818,N_25819,N_25820,N_25821,N_25822,N_25823,N_25824,N_25825,N_25826,N_25827,N_25828,N_25829,N_25830,N_25831,N_25832,N_25833,N_25834,N_25835,N_25836,N_25837,N_25838,N_25839,N_25840,N_25841,N_25842,N_25843,N_25844,N_25845,N_25846,N_25847,N_25848,N_25849,N_25850,N_25851,N_25852,N_25853,N_25854,N_25855,N_25856,N_25857,N_25858,N_25859,N_25860,N_25861,N_25862,N_25863,N_25864,N_25865,N_25866,N_25867,N_25868,N_25869,N_25870,N_25871,N_25872,N_25873,N_25874,N_25875,N_25876,N_25877,N_25878,N_25879,N_25880,N_25881,N_25882,N_25883,N_25884,N_25885,N_25886,N_25887,N_25888,N_25889,N_25890,N_25891,N_25892,N_25893,N_25894,N_25895,N_25896,N_25897,N_25898,N_25899,N_25900,N_25901,N_25902,N_25903,N_25904,N_25905,N_25906,N_25907,N_25908,N_25909,N_25910,N_25911,N_25912,N_25913,N_25914,N_25915,N_25916,N_25917,N_25918,N_25919,N_25920,N_25921,N_25922,N_25923,N_25924,N_25925,N_25926,N_25927,N_25928,N_25929,N_25930,N_25931,N_25932,N_25933,N_25934,N_25935,N_25936,N_25937,N_25938,N_25939,N_25940,N_25941,N_25942,N_25943,N_25944,N_25945,N_25946,N_25947,N_25948,N_25949,N_25950,N_25951,N_25952,N_25953,N_25954,N_25955,N_25956,N_25957,N_25958,N_25959,N_25960,N_25961,N_25962,N_25963,N_25964,N_25965,N_25966,N_25967,N_25968,N_25969,N_25970,N_25971,N_25972,N_25973,N_25974,N_25975,N_25976,N_25977,N_25978,N_25979,N_25980,N_25981,N_25982,N_25983,N_25984,N_25985,N_25986,N_25987,N_25988,N_25989,N_25990,N_25991,N_25992,N_25993,N_25994,N_25995,N_25996,N_25997,N_25998,N_25999,N_26000,N_26001,N_26002,N_26003,N_26004,N_26005,N_26006,N_26007,N_26008,N_26009,N_26010,N_26011,N_26012,N_26013,N_26014,N_26015,N_26016,N_26017,N_26018,N_26019,N_26020,N_26021,N_26022,N_26023,N_26024,N_26025,N_26026,N_26027,N_26028,N_26029,N_26030,N_26031,N_26032,N_26033,N_26034,N_26035,N_26036,N_26037,N_26038,N_26039,N_26040,N_26041,N_26042,N_26043,N_26044,N_26045,N_26046,N_26047,N_26048,N_26049,N_26050,N_26051,N_26052,N_26053,N_26054,N_26055,N_26056,N_26057,N_26058,N_26059,N_26060,N_26061,N_26062,N_26063,N_26064,N_26065,N_26066,N_26067,N_26068,N_26069,N_26070,N_26071,N_26072,N_26073,N_26074,N_26075,N_26076,N_26077,N_26078,N_26079,N_26080,N_26081,N_26082,N_26083,N_26084,N_26085,N_26086,N_26087,N_26088,N_26089,N_26090,N_26091,N_26092,N_26093,N_26094,N_26095,N_26096,N_26097,N_26098,N_26099,N_26100,N_26101,N_26102,N_26103,N_26104,N_26105,N_26106,N_26107,N_26108,N_26109,N_26110,N_26111,N_26112,N_26113,N_26114,N_26115,N_26116,N_26117,N_26118,N_26119,N_26120,N_26121,N_26122,N_26123,N_26124,N_26125,N_26126,N_26127,N_26128,N_26129,N_26130,N_26131,N_26132,N_26133,N_26134,N_26135,N_26136,N_26137,N_26138,N_26139,N_26140,N_26141,N_26142,N_26143,N_26144,N_26145,N_26146,N_26147,N_26148,N_26149,N_26150,N_26151,N_26152,N_26153,N_26154,N_26155,N_26156,N_26157,N_26158,N_26159,N_26160,N_26161,N_26162,N_26163,N_26164,N_26165,N_26166,N_26167,N_26168,N_26169,N_26170,N_26171,N_26172,N_26173,N_26174,N_26175,N_26176,N_26177,N_26178,N_26179,N_26180,N_26181,N_26182,N_26183,N_26184,N_26185,N_26186,N_26187,N_26188,N_26189,N_26190,N_26191,N_26192,N_26193,N_26194,N_26195,N_26196,N_26197,N_26198,N_26199,N_26200,N_26201,N_26202,N_26203,N_26204,N_26205,N_26206,N_26207,N_26208,N_26209,N_26210,N_26211,N_26212,N_26213,N_26214,N_26215,N_26216,N_26217,N_26218,N_26219,N_26220,N_26221,N_26222,N_26223,N_26224,N_26225,N_26226,N_26227,N_26228,N_26229,N_26230,N_26231,N_26232,N_26233,N_26234,N_26235,N_26236,N_26237,N_26238,N_26239,N_26240,N_26241,N_26242,N_26243,N_26244,N_26245,N_26246,N_26247,N_26248,N_26249,N_26250,N_26251,N_26252,N_26253,N_26254,N_26255,N_26256,N_26257,N_26258,N_26259,N_26260,N_26261,N_26262,N_26263,N_26264,N_26265,N_26266,N_26267,N_26268,N_26269,N_26270,N_26271,N_26272,N_26273,N_26274,N_26275,N_26276,N_26277,N_26278,N_26279,N_26280,N_26281,N_26282,N_26283,N_26284,N_26285,N_26286,N_26287,N_26288,N_26289,N_26290,N_26291,N_26292,N_26293,N_26294,N_26295,N_26296,N_26297,N_26298,N_26299,N_26300,N_26301,N_26302,N_26303,N_26304,N_26305,N_26306,N_26307,N_26308,N_26309,N_26310,N_26311,N_26312,N_26313,N_26314,N_26315,N_26316,N_26317,N_26318,N_26319,N_26320,N_26321,N_26322,N_26323,N_26324,N_26325,N_26326,N_26327,N_26328,N_26329,N_26330,N_26331,N_26332,N_26333,N_26334,N_26335,N_26336,N_26337,N_26338,N_26339,N_26340,N_26341,N_26342,N_26343,N_26344,N_26345,N_26346,N_26347,N_26348,N_26349,N_26350,N_26351,N_26352,N_26353,N_26354,N_26355,N_26356,N_26357,N_26358,N_26359,N_26360,N_26361,N_26362,N_26363,N_26364,N_26365,N_26366,N_26367,N_26368,N_26369,N_26370,N_26371,N_26372,N_26373,N_26374,N_26375,N_26376,N_26377,N_26378,N_26379,N_26380,N_26381,N_26382,N_26383,N_26384,N_26385,N_26386,N_26387,N_26388,N_26389,N_26390,N_26391,N_26392,N_26393,N_26394,N_26395,N_26396,N_26397,N_26398,N_26399,N_26400,N_26401,N_26402,N_26403,N_26404,N_26405,N_26406,N_26407,N_26408,N_26409,N_26410,N_26411,N_26412,N_26413,N_26414,N_26415,N_26416,N_26417,N_26418,N_26419,N_26420,N_26421,N_26422,N_26423,N_26424,N_26425,N_26426,N_26427,N_26428,N_26429,N_26430,N_26431,N_26432,N_26433,N_26434,N_26435,N_26436,N_26437,N_26438,N_26439,N_26440,N_26441,N_26442,N_26443,N_26444,N_26445,N_26446,N_26447,N_26448,N_26449,N_26450,N_26451,N_26452,N_26453,N_26454,N_26455,N_26456,N_26457,N_26458,N_26459,N_26460,N_26461,N_26462,N_26463,N_26464,N_26465,N_26466,N_26467,N_26468,N_26469,N_26470,N_26471,N_26472,N_26473,N_26474,N_26475,N_26476,N_26477,N_26478,N_26479,N_26480,N_26481,N_26482,N_26483,N_26484,N_26485,N_26486,N_26487,N_26488,N_26489,N_26490,N_26491,N_26492,N_26493,N_26494,N_26495,N_26496,N_26497,N_26498,N_26499,N_26500,N_26501,N_26502,N_26503,N_26504,N_26505,N_26506,N_26507,N_26508,N_26509,N_26510,N_26511,N_26512,N_26513,N_26514,N_26515,N_26516,N_26517,N_26518,N_26519,N_26520,N_26521,N_26522,N_26523,N_26524,N_26525,N_26526,N_26527,N_26528,N_26529,N_26530,N_26531,N_26532,N_26533,N_26534,N_26535,N_26536,N_26537,N_26538,N_26539,N_26540,N_26541,N_26542,N_26543,N_26544,N_26545,N_26546,N_26547,N_26548,N_26549,N_26550,N_26551,N_26552,N_26553,N_26554,N_26555,N_26556,N_26557,N_26558,N_26559,N_26560,N_26561,N_26562,N_26563,N_26564,N_26565,N_26566,N_26567,N_26568,N_26569,N_26570,N_26571,N_26572,N_26573,N_26574,N_26575,N_26576,N_26577,N_26578,N_26579,N_26580,N_26581,N_26582,N_26583,N_26584,N_26585,N_26586,N_26587,N_26588,N_26589,N_26590,N_26591,N_26592,N_26593,N_26594,N_26595,N_26596,N_26597,N_26598,N_26599,N_26600,N_26601,N_26602,N_26603,N_26604,N_26605,N_26606,N_26607,N_26608,N_26609,N_26610,N_26611,N_26612,N_26613,N_26614,N_26615,N_26616,N_26617,N_26618,N_26619,N_26620,N_26621,N_26622,N_26623,N_26624,N_26625,N_26626,N_26627,N_26628,N_26629,N_26630,N_26631,N_26632,N_26633,N_26634,N_26635,N_26636,N_26637,N_26638,N_26639,N_26640,N_26641,N_26642,N_26643,N_26644,N_26645,N_26646,N_26647,N_26648,N_26649,N_26650,N_26651,N_26652,N_26653,N_26654,N_26655,N_26656,N_26657,N_26658,N_26659,N_26660,N_26661,N_26662,N_26663,N_26664,N_26665,N_26666,N_26667,N_26668,N_26669,N_26670,N_26671,N_26672,N_26673,N_26674,N_26675,N_26676,N_26677,N_26678,N_26679,N_26680,N_26681,N_26682,N_26683,N_26684,N_26685,N_26686,N_26687,N_26688,N_26689,N_26690,N_26691,N_26692,N_26693,N_26694,N_26695,N_26696,N_26697,N_26698,N_26699,N_26700,N_26701,N_26702,N_26703,N_26704,N_26705,N_26706,N_26707,N_26708,N_26709,N_26710,N_26711,N_26712,N_26713,N_26714,N_26715,N_26716,N_26717,N_26718,N_26719,N_26720,N_26721,N_26722,N_26723,N_26724,N_26725,N_26726,N_26727,N_26728,N_26729,N_26730,N_26731,N_26732,N_26733,N_26734,N_26735,N_26736,N_26737,N_26738,N_26739,N_26740,N_26741,N_26742,N_26743,N_26744,N_26745,N_26746,N_26747,N_26748,N_26749,N_26750,N_26751,N_26752,N_26753,N_26754,N_26755,N_26756,N_26757,N_26758,N_26759,N_26760,N_26761,N_26762,N_26763,N_26764,N_26765,N_26766,N_26767,N_26768,N_26769,N_26770,N_26771,N_26772,N_26773,N_26774,N_26775,N_26776,N_26777,N_26778,N_26779,N_26780,N_26781,N_26782,N_26783,N_26784,N_26785,N_26786,N_26787,N_26788,N_26789,N_26790,N_26791,N_26792,N_26793,N_26794,N_26795,N_26796,N_26797,N_26798,N_26799,N_26800,N_26801,N_26802,N_26803,N_26804,N_26805,N_26806,N_26807,N_26808,N_26809,N_26810,N_26811,N_26812,N_26813,N_26814,N_26815,N_26816,N_26817,N_26818,N_26819,N_26820,N_26821,N_26822,N_26823,N_26824,N_26825,N_26826,N_26827,N_26828,N_26829,N_26830,N_26831,N_26832,N_26833,N_26834,N_26835,N_26836,N_26837,N_26838,N_26839,N_26840,N_26841,N_26842,N_26843,N_26844,N_26845,N_26846,N_26847,N_26848,N_26849,N_26850,N_26851,N_26852,N_26853,N_26854,N_26855,N_26856,N_26857,N_26858,N_26859,N_26860,N_26861,N_26862,N_26863,N_26864,N_26865,N_26866,N_26867,N_26868,N_26869,N_26870,N_26871,N_26872,N_26873,N_26874,N_26875,N_26876,N_26877,N_26878,N_26879,N_26880,N_26881,N_26882,N_26883,N_26884,N_26885,N_26886,N_26887,N_26888,N_26889,N_26890,N_26891,N_26892,N_26893,N_26894,N_26895,N_26896,N_26897,N_26898,N_26899,N_26900,N_26901,N_26902,N_26903,N_26904,N_26905,N_26906,N_26907,N_26908,N_26909,N_26910,N_26911,N_26912,N_26913,N_26914,N_26915,N_26916,N_26917,N_26918,N_26919,N_26920,N_26921,N_26922,N_26923,N_26924,N_26925,N_26926,N_26927,N_26928,N_26929,N_26930,N_26931,N_26932,N_26933,N_26934,N_26935,N_26936,N_26937,N_26938,N_26939,N_26940,N_26941,N_26942,N_26943,N_26944,N_26945,N_26946,N_26947,N_26948,N_26949,N_26950,N_26951,N_26952,N_26953,N_26954,N_26955,N_26956,N_26957,N_26958,N_26959,N_26960,N_26961,N_26962,N_26963,N_26964,N_26965,N_26966,N_26967,N_26968,N_26969,N_26970,N_26971,N_26972,N_26973,N_26974,N_26975,N_26976,N_26977,N_26978,N_26979,N_26980,N_26981,N_26982,N_26983,N_26984,N_26985,N_26986,N_26987,N_26988,N_26989,N_26990,N_26991,N_26992,N_26993,N_26994,N_26995,N_26996,N_26997,N_26998,N_26999,N_27000,N_27001,N_27002,N_27003,N_27004,N_27005,N_27006,N_27007,N_27008,N_27009,N_27010,N_27011,N_27012,N_27013,N_27014,N_27015,N_27016,N_27017,N_27018,N_27019,N_27020,N_27021,N_27022,N_27023,N_27024,N_27025,N_27026,N_27027,N_27028,N_27029,N_27030,N_27031,N_27032,N_27033,N_27034,N_27035,N_27036,N_27037,N_27038,N_27039,N_27040,N_27041,N_27042,N_27043,N_27044,N_27045,N_27046,N_27047,N_27048,N_27049,N_27050,N_27051,N_27052,N_27053,N_27054,N_27055,N_27056,N_27057,N_27058,N_27059,N_27060,N_27061,N_27062,N_27063,N_27064,N_27065,N_27066,N_27067,N_27068,N_27069,N_27070,N_27071,N_27072,N_27073,N_27074,N_27075,N_27076,N_27077,N_27078,N_27079,N_27080,N_27081,N_27082,N_27083,N_27084,N_27085,N_27086,N_27087,N_27088,N_27089,N_27090,N_27091,N_27092,N_27093,N_27094,N_27095,N_27096,N_27097,N_27098,N_27099,N_27100,N_27101,N_27102,N_27103,N_27104,N_27105,N_27106,N_27107,N_27108,N_27109,N_27110,N_27111,N_27112,N_27113,N_27114,N_27115,N_27116,N_27117,N_27118,N_27119,N_27120,N_27121,N_27122,N_27123,N_27124,N_27125,N_27126,N_27127,N_27128,N_27129,N_27130,N_27131,N_27132,N_27133,N_27134,N_27135,N_27136,N_27137,N_27138,N_27139,N_27140,N_27141,N_27142,N_27143,N_27144,N_27145,N_27146,N_27147,N_27148,N_27149,N_27150,N_27151,N_27152,N_27153,N_27154,N_27155,N_27156,N_27157,N_27158,N_27159,N_27160,N_27161,N_27162,N_27163,N_27164,N_27165,N_27166,N_27167,N_27168,N_27169,N_27170,N_27171,N_27172,N_27173,N_27174,N_27175,N_27176,N_27177,N_27178,N_27179,N_27180,N_27181,N_27182,N_27183,N_27184,N_27185,N_27186,N_27187,N_27188,N_27189,N_27190,N_27191,N_27192,N_27193,N_27194,N_27195,N_27196,N_27197,N_27198,N_27199,N_27200,N_27201,N_27202,N_27203,N_27204,N_27205,N_27206,N_27207,N_27208,N_27209,N_27210,N_27211,N_27212,N_27213,N_27214,N_27215,N_27216,N_27217,N_27218,N_27219,N_27220,N_27221,N_27222,N_27223,N_27224,N_27225,N_27226,N_27227,N_27228,N_27229,N_27230,N_27231,N_27232,N_27233,N_27234,N_27235,N_27236,N_27237,N_27238,N_27239,N_27240,N_27241,N_27242,N_27243,N_27244,N_27245,N_27246,N_27247,N_27248,N_27249,N_27250,N_27251,N_27252,N_27253,N_27254,N_27255,N_27256,N_27257,N_27258,N_27259,N_27260,N_27261,N_27262,N_27263,N_27264,N_27265,N_27266,N_27267,N_27268,N_27269,N_27270,N_27271,N_27272,N_27273,N_27274,N_27275,N_27276,N_27277,N_27278,N_27279,N_27280,N_27281,N_27282,N_27283,N_27284,N_27285,N_27286,N_27287,N_27288,N_27289,N_27290,N_27291,N_27292,N_27293,N_27294,N_27295,N_27296,N_27297,N_27298,N_27299,N_27300,N_27301,N_27302,N_27303,N_27304,N_27305,N_27306,N_27307,N_27308,N_27309,N_27310,N_27311,N_27312,N_27313,N_27314,N_27315,N_27316,N_27317,N_27318,N_27319,N_27320,N_27321,N_27322,N_27323,N_27324,N_27325,N_27326,N_27327,N_27328,N_27329,N_27330,N_27331,N_27332,N_27333,N_27334,N_27335,N_27336,N_27337,N_27338,N_27339,N_27340,N_27341,N_27342,N_27343,N_27344,N_27345,N_27346,N_27347,N_27348,N_27349,N_27350,N_27351,N_27352,N_27353,N_27354,N_27355,N_27356,N_27357,N_27358,N_27359,N_27360,N_27361,N_27362,N_27363,N_27364,N_27365,N_27366,N_27367,N_27368,N_27369,N_27370,N_27371,N_27372,N_27373,N_27374,N_27375,N_27376,N_27377,N_27378,N_27379,N_27380,N_27381,N_27382,N_27383,N_27384,N_27385,N_27386,N_27387,N_27388,N_27389,N_27390,N_27391,N_27392,N_27393,N_27394,N_27395,N_27396,N_27397,N_27398,N_27399,N_27400,N_27401,N_27402,N_27403,N_27404,N_27405,N_27406,N_27407,N_27408,N_27409,N_27410,N_27411,N_27412,N_27413,N_27414,N_27415,N_27416,N_27417,N_27418,N_27419,N_27420,N_27421,N_27422,N_27423,N_27424,N_27425,N_27426,N_27427,N_27428,N_27429,N_27430,N_27431,N_27432,N_27433,N_27434,N_27435,N_27436,N_27437,N_27438,N_27439,N_27440,N_27441,N_27442,N_27443,N_27444,N_27445,N_27446,N_27447,N_27448,N_27449,N_27450,N_27451,N_27452,N_27453,N_27454,N_27455,N_27456,N_27457,N_27458,N_27459,N_27460,N_27461,N_27462,N_27463,N_27464,N_27465,N_27466,N_27467,N_27468,N_27469,N_27470,N_27471,N_27472,N_27473,N_27474,N_27475,N_27476,N_27477,N_27478,N_27479,N_27480,N_27481,N_27482,N_27483,N_27484,N_27485,N_27486,N_27487,N_27488,N_27489,N_27490,N_27491,N_27492,N_27493,N_27494,N_27495,N_27496,N_27497,N_27498,N_27499,N_27500,N_27501,N_27502,N_27503,N_27504,N_27505,N_27506,N_27507,N_27508,N_27509,N_27510,N_27511,N_27512,N_27513,N_27514,N_27515,N_27516,N_27517,N_27518,N_27519,N_27520,N_27521,N_27522,N_27523,N_27524,N_27525,N_27526,N_27527,N_27528,N_27529,N_27530,N_27531,N_27532,N_27533,N_27534,N_27535,N_27536,N_27537,N_27538,N_27539,N_27540,N_27541,N_27542,N_27543,N_27544,N_27545,N_27546,N_27547,N_27548,N_27549,N_27550,N_27551,N_27552,N_27553,N_27554,N_27555,N_27556,N_27557,N_27558,N_27559,N_27560,N_27561,N_27562,N_27563,N_27564,N_27565,N_27566,N_27567,N_27568,N_27569,N_27570,N_27571,N_27572,N_27573,N_27574,N_27575,N_27576,N_27577,N_27578,N_27579,N_27580,N_27581,N_27582,N_27583,N_27584,N_27585,N_27586,N_27587,N_27588,N_27589,N_27590,N_27591,N_27592,N_27593,N_27594,N_27595,N_27596,N_27597,N_27598,N_27599,N_27600,N_27601,N_27602,N_27603,N_27604,N_27605,N_27606,N_27607,N_27608,N_27609,N_27610,N_27611,N_27612,N_27613,N_27614,N_27615,N_27616,N_27617,N_27618,N_27619,N_27620,N_27621,N_27622,N_27623,N_27624,N_27625,N_27626,N_27627,N_27628,N_27629,N_27630,N_27631,N_27632,N_27633,N_27634,N_27635,N_27636,N_27637,N_27638,N_27639,N_27640,N_27641,N_27642,N_27643,N_27644,N_27645,N_27646,N_27647,N_27648,N_27649,N_27650,N_27651,N_27652,N_27653,N_27654,N_27655,N_27656,N_27657,N_27658,N_27659,N_27660,N_27661,N_27662,N_27663,N_27664,N_27665,N_27666,N_27667,N_27668,N_27669,N_27670,N_27671,N_27672,N_27673,N_27674,N_27675,N_27676,N_27677,N_27678,N_27679,N_27680,N_27681,N_27682,N_27683,N_27684,N_27685,N_27686,N_27687,N_27688,N_27689,N_27690,N_27691,N_27692,N_27693,N_27694,N_27695,N_27696,N_27697,N_27698,N_27699,N_27700,N_27701,N_27702,N_27703,N_27704,N_27705,N_27706,N_27707,N_27708,N_27709,N_27710,N_27711,N_27712,N_27713,N_27714,N_27715,N_27716,N_27717,N_27718,N_27719,N_27720,N_27721,N_27722,N_27723,N_27724,N_27725,N_27726,N_27727,N_27728,N_27729,N_27730,N_27731,N_27732,N_27733,N_27734,N_27735,N_27736,N_27737,N_27738,N_27739,N_27740,N_27741,N_27742,N_27743,N_27744,N_27745,N_27746,N_27747,N_27748,N_27749,N_27750,N_27751,N_27752,N_27753,N_27754,N_27755,N_27756,N_27757,N_27758,N_27759,N_27760,N_27761,N_27762,N_27763,N_27764,N_27765,N_27766,N_27767,N_27768,N_27769,N_27770,N_27771,N_27772,N_27773,N_27774,N_27775,N_27776,N_27777,N_27778,N_27779,N_27780,N_27781,N_27782,N_27783,N_27784,N_27785,N_27786,N_27787,N_27788,N_27789,N_27790,N_27791,N_27792,N_27793,N_27794,N_27795,N_27796,N_27797,N_27798,N_27799,N_27800,N_27801,N_27802,N_27803,N_27804,N_27805,N_27806,N_27807,N_27808,N_27809,N_27810,N_27811,N_27812,N_27813,N_27814,N_27815,N_27816,N_27817,N_27818,N_27819,N_27820,N_27821,N_27822,N_27823,N_27824,N_27825,N_27826,N_27827,N_27828,N_27829,N_27830,N_27831,N_27832,N_27833,N_27834,N_27835,N_27836,N_27837,N_27838,N_27839,N_27840,N_27841,N_27842,N_27843,N_27844,N_27845,N_27846,N_27847,N_27848,N_27849,N_27850,N_27851,N_27852,N_27853,N_27854,N_27855,N_27856,N_27857,N_27858,N_27859,N_27860,N_27861,N_27862,N_27863,N_27864,N_27865,N_27866,N_27867,N_27868,N_27869,N_27870,N_27871,N_27872,N_27873,N_27874,N_27875,N_27876,N_27877,N_27878,N_27879,N_27880,N_27881,N_27882,N_27883,N_27884,N_27885,N_27886,N_27887,N_27888,N_27889,N_27890,N_27891,N_27892,N_27893,N_27894,N_27895,N_27896,N_27897,N_27898,N_27899,N_27900,N_27901,N_27902,N_27903,N_27904,N_27905,N_27906,N_27907,N_27908,N_27909,N_27910,N_27911,N_27912,N_27913,N_27914,N_27915,N_27916,N_27917,N_27918,N_27919,N_27920,N_27921,N_27922,N_27923,N_27924,N_27925,N_27926,N_27927,N_27928,N_27929,N_27930,N_27931,N_27932,N_27933,N_27934,N_27935,N_27936,N_27937,N_27938,N_27939,N_27940,N_27941,N_27942,N_27943,N_27944,N_27945,N_27946,N_27947,N_27948,N_27949,N_27950,N_27951,N_27952,N_27953,N_27954,N_27955,N_27956,N_27957,N_27958,N_27959,N_27960,N_27961,N_27962,N_27963,N_27964,N_27965,N_27966,N_27967,N_27968,N_27969,N_27970,N_27971,N_27972,N_27973,N_27974,N_27975,N_27976,N_27977,N_27978,N_27979,N_27980,N_27981,N_27982,N_27983,N_27984,N_27985,N_27986,N_27987,N_27988,N_27989,N_27990,N_27991,N_27992,N_27993,N_27994,N_27995,N_27996,N_27997,N_27998,N_27999,N_28000,N_28001,N_28002,N_28003,N_28004,N_28005,N_28006,N_28007,N_28008,N_28009,N_28010,N_28011,N_28012,N_28013,N_28014,N_28015,N_28016,N_28017,N_28018,N_28019,N_28020,N_28021,N_28022,N_28023,N_28024,N_28025,N_28026,N_28027,N_28028,N_28029,N_28030,N_28031,N_28032,N_28033,N_28034,N_28035,N_28036,N_28037,N_28038,N_28039,N_28040,N_28041,N_28042,N_28043,N_28044,N_28045,N_28046,N_28047,N_28048,N_28049,N_28050,N_28051,N_28052,N_28053,N_28054,N_28055,N_28056,N_28057,N_28058,N_28059,N_28060,N_28061,N_28062,N_28063,N_28064,N_28065,N_28066,N_28067,N_28068,N_28069,N_28070,N_28071,N_28072,N_28073,N_28074,N_28075,N_28076,N_28077,N_28078,N_28079,N_28080,N_28081,N_28082,N_28083,N_28084,N_28085,N_28086,N_28087,N_28088,N_28089,N_28090,N_28091,N_28092,N_28093,N_28094,N_28095,N_28096,N_28097,N_28098,N_28099,N_28100,N_28101,N_28102,N_28103,N_28104,N_28105,N_28106,N_28107,N_28108,N_28109,N_28110,N_28111,N_28112,N_28113,N_28114,N_28115,N_28116,N_28117,N_28118,N_28119,N_28120,N_28121,N_28122,N_28123,N_28124,N_28125,N_28126,N_28127,N_28128,N_28129,N_28130,N_28131,N_28132,N_28133,N_28134,N_28135,N_28136,N_28137,N_28138,N_28139,N_28140,N_28141,N_28142,N_28143,N_28144,N_28145,N_28146,N_28147,N_28148,N_28149,N_28150,N_28151,N_28152,N_28153,N_28154,N_28155,N_28156,N_28157,N_28158,N_28159,N_28160,N_28161,N_28162,N_28163,N_28164,N_28165,N_28166,N_28167,N_28168,N_28169,N_28170,N_28171,N_28172,N_28173,N_28174,N_28175,N_28176,N_28177,N_28178,N_28179,N_28180,N_28181,N_28182,N_28183,N_28184,N_28185,N_28186,N_28187,N_28188,N_28189,N_28190,N_28191,N_28192,N_28193,N_28194,N_28195,N_28196,N_28197,N_28198,N_28199,N_28200,N_28201,N_28202,N_28203,N_28204,N_28205,N_28206,N_28207,N_28208,N_28209,N_28210,N_28211,N_28212,N_28213,N_28214,N_28215,N_28216,N_28217,N_28218,N_28219,N_28220,N_28221,N_28222,N_28223,N_28224,N_28225,N_28226,N_28227,N_28228,N_28229,N_28230,N_28231,N_28232,N_28233,N_28234,N_28235,N_28236,N_28237,N_28238,N_28239,N_28240,N_28241,N_28242,N_28243,N_28244,N_28245,N_28246,N_28247,N_28248,N_28249,N_28250,N_28251,N_28252,N_28253,N_28254,N_28255,N_28256,N_28257,N_28258,N_28259,N_28260,N_28261,N_28262,N_28263,N_28264,N_28265,N_28266,N_28267,N_28268,N_28269,N_28270,N_28271,N_28272,N_28273,N_28274,N_28275,N_28276,N_28277,N_28278,N_28279,N_28280,N_28281,N_28282,N_28283,N_28284,N_28285,N_28286,N_28287,N_28288,N_28289,N_28290,N_28291,N_28292,N_28293,N_28294,N_28295,N_28296,N_28297,N_28298,N_28299,N_28300,N_28301,N_28302,N_28303,N_28304,N_28305,N_28306,N_28307,N_28308,N_28309,N_28310,N_28311,N_28312,N_28313,N_28314,N_28315,N_28316,N_28317,N_28318,N_28319,N_28320,N_28321,N_28322,N_28323,N_28324,N_28325,N_28326,N_28327,N_28328,N_28329,N_28330,N_28331,N_28332,N_28333,N_28334,N_28335,N_28336,N_28337,N_28338,N_28339,N_28340,N_28341,N_28342,N_28343,N_28344,N_28345,N_28346,N_28347,N_28348,N_28349,N_28350,N_28351,N_28352,N_28353,N_28354,N_28355,N_28356,N_28357,N_28358,N_28359,N_28360,N_28361,N_28362,N_28363,N_28364,N_28365,N_28366,N_28367,N_28368,N_28369,N_28370,N_28371,N_28372,N_28373,N_28374,N_28375,N_28376,N_28377,N_28378,N_28379,N_28380,N_28381,N_28382,N_28383,N_28384,N_28385,N_28386,N_28387,N_28388,N_28389,N_28390,N_28391,N_28392,N_28393,N_28394,N_28395,N_28396,N_28397,N_28398,N_28399,N_28400,N_28401,N_28402,N_28403,N_28404,N_28405,N_28406,N_28407,N_28408,N_28409,N_28410,N_28411,N_28412,N_28413,N_28414,N_28415,N_28416,N_28417,N_28418,N_28419,N_28420,N_28421,N_28422,N_28423,N_28424,N_28425,N_28426,N_28427,N_28428,N_28429,N_28430,N_28431,N_28432,N_28433,N_28434,N_28435,N_28436,N_28437,N_28438,N_28439,N_28440,N_28441,N_28442,N_28443,N_28444,N_28445,N_28446,N_28447,N_28448,N_28449,N_28450,N_28451,N_28452,N_28453,N_28454,N_28455,N_28456,N_28457,N_28458,N_28459,N_28460,N_28461,N_28462,N_28463,N_28464,N_28465,N_28466,N_28467,N_28468,N_28469,N_28470,N_28471,N_28472,N_28473,N_28474,N_28475,N_28476,N_28477,N_28478,N_28479,N_28480,N_28481,N_28482,N_28483,N_28484,N_28485,N_28486,N_28487,N_28488,N_28489,N_28490,N_28491,N_28492,N_28493,N_28494,N_28495,N_28496,N_28497,N_28498,N_28499,N_28500,N_28501,N_28502,N_28503,N_28504,N_28505,N_28506,N_28507,N_28508,N_28509,N_28510,N_28511,N_28512,N_28513,N_28514,N_28515,N_28516,N_28517,N_28518,N_28519,N_28520,N_28521,N_28522,N_28523,N_28524,N_28525,N_28526,N_28527,N_28528,N_28529,N_28530,N_28531,N_28532,N_28533,N_28534,N_28535,N_28536,N_28537,N_28538,N_28539,N_28540,N_28541,N_28542,N_28543,N_28544,N_28545,N_28546,N_28547,N_28548,N_28549,N_28550,N_28551,N_28552,N_28553,N_28554,N_28555,N_28556,N_28557,N_28558,N_28559,N_28560,N_28561,N_28562,N_28563,N_28564,N_28565,N_28566,N_28567,N_28568,N_28569,N_28570,N_28571,N_28572,N_28573,N_28574,N_28575,N_28576,N_28577,N_28578,N_28579,N_28580,N_28581,N_28582,N_28583,N_28584,N_28585,N_28586,N_28587,N_28588,N_28589,N_28590,N_28591,N_28592,N_28593,N_28594,N_28595,N_28596,N_28597,N_28598,N_28599,N_28600,N_28601,N_28602,N_28603,N_28604,N_28605,N_28606,N_28607,N_28608,N_28609,N_28610,N_28611,N_28612,N_28613,N_28614,N_28615,N_28616,N_28617,N_28618,N_28619,N_28620,N_28621,N_28622,N_28623,N_28624,N_28625,N_28626,N_28627,N_28628,N_28629,N_28630,N_28631,N_28632,N_28633,N_28634,N_28635,N_28636,N_28637,N_28638,N_28639,N_28640,N_28641,N_28642,N_28643,N_28644,N_28645,N_28646,N_28647,N_28648,N_28649,N_28650,N_28651,N_28652,N_28653,N_28654,N_28655,N_28656,N_28657,N_28658,N_28659,N_28660,N_28661,N_28662,N_28663,N_28664,N_28665,N_28666,N_28667,N_28668,N_28669,N_28670,N_28671,N_28672,N_28673,N_28674,N_28675,N_28676,N_28677,N_28678,N_28679,N_28680,N_28681,N_28682,N_28683,N_28684,N_28685,N_28686,N_28687,N_28688,N_28689,N_28690,N_28691,N_28692,N_28693,N_28694,N_28695,N_28696,N_28697,N_28698,N_28699,N_28700,N_28701,N_28702,N_28703,N_28704,N_28705,N_28706,N_28707,N_28708,N_28709,N_28710,N_28711,N_28712,N_28713,N_28714,N_28715,N_28716,N_28717,N_28718,N_28719,N_28720,N_28721,N_28722,N_28723,N_28724,N_28725,N_28726,N_28727,N_28728,N_28729,N_28730,N_28731,N_28732,N_28733,N_28734,N_28735,N_28736,N_28737,N_28738,N_28739,N_28740,N_28741,N_28742,N_28743,N_28744,N_28745,N_28746,N_28747,N_28748,N_28749,N_28750,N_28751,N_28752,N_28753,N_28754,N_28755,N_28756,N_28757,N_28758,N_28759,N_28760,N_28761,N_28762,N_28763,N_28764,N_28765,N_28766,N_28767,N_28768,N_28769,N_28770,N_28771,N_28772,N_28773,N_28774,N_28775,N_28776,N_28777,N_28778,N_28779,N_28780,N_28781,N_28782,N_28783,N_28784,N_28785,N_28786,N_28787,N_28788,N_28789,N_28790,N_28791,N_28792,N_28793,N_28794,N_28795,N_28796,N_28797,N_28798,N_28799,N_28800,N_28801,N_28802,N_28803,N_28804,N_28805,N_28806,N_28807,N_28808,N_28809,N_28810,N_28811,N_28812,N_28813,N_28814,N_28815,N_28816,N_28817,N_28818,N_28819,N_28820,N_28821,N_28822,N_28823,N_28824,N_28825,N_28826,N_28827,N_28828,N_28829,N_28830,N_28831,N_28832,N_28833,N_28834,N_28835,N_28836,N_28837,N_28838,N_28839,N_28840,N_28841,N_28842,N_28843,N_28844,N_28845,N_28846,N_28847,N_28848,N_28849,N_28850,N_28851,N_28852,N_28853,N_28854,N_28855,N_28856,N_28857,N_28858,N_28859,N_28860,N_28861,N_28862,N_28863,N_28864,N_28865,N_28866,N_28867,N_28868,N_28869,N_28870,N_28871,N_28872,N_28873,N_28874,N_28875,N_28876,N_28877,N_28878,N_28879,N_28880,N_28881,N_28882,N_28883,N_28884,N_28885,N_28886,N_28887,N_28888,N_28889,N_28890,N_28891,N_28892,N_28893,N_28894,N_28895,N_28896,N_28897,N_28898,N_28899,N_28900,N_28901,N_28902,N_28903,N_28904,N_28905,N_28906,N_28907,N_28908,N_28909,N_28910,N_28911,N_28912,N_28913,N_28914,N_28915,N_28916,N_28917,N_28918,N_28919,N_28920,N_28921,N_28922,N_28923,N_28924,N_28925,N_28926,N_28927,N_28928,N_28929,N_28930,N_28931,N_28932,N_28933,N_28934,N_28935,N_28936,N_28937,N_28938,N_28939,N_28940,N_28941,N_28942,N_28943,N_28944,N_28945,N_28946,N_28947,N_28948,N_28949,N_28950,N_28951,N_28952,N_28953,N_28954,N_28955,N_28956,N_28957,N_28958,N_28959,N_28960,N_28961,N_28962,N_28963,N_28964,N_28965,N_28966,N_28967,N_28968,N_28969,N_28970,N_28971,N_28972,N_28973,N_28974,N_28975,N_28976,N_28977,N_28978,N_28979,N_28980,N_28981,N_28982,N_28983,N_28984,N_28985,N_28986,N_28987,N_28988,N_28989,N_28990,N_28991,N_28992,N_28993,N_28994,N_28995,N_28996,N_28997,N_28998,N_28999,N_29000,N_29001,N_29002,N_29003,N_29004,N_29005,N_29006,N_29007,N_29008,N_29009,N_29010,N_29011,N_29012,N_29013,N_29014,N_29015,N_29016,N_29017,N_29018,N_29019,N_29020,N_29021,N_29022,N_29023,N_29024,N_29025,N_29026,N_29027,N_29028,N_29029,N_29030,N_29031,N_29032,N_29033,N_29034,N_29035,N_29036,N_29037,N_29038,N_29039,N_29040,N_29041,N_29042,N_29043,N_29044,N_29045,N_29046,N_29047,N_29048,N_29049,N_29050,N_29051,N_29052,N_29053,N_29054,N_29055,N_29056,N_29057,N_29058,N_29059,N_29060,N_29061,N_29062,N_29063,N_29064,N_29065,N_29066,N_29067,N_29068,N_29069,N_29070,N_29071,N_29072,N_29073,N_29074,N_29075,N_29076,N_29077,N_29078,N_29079,N_29080,N_29081,N_29082,N_29083,N_29084,N_29085,N_29086,N_29087,N_29088,N_29089,N_29090,N_29091,N_29092,N_29093,N_29094,N_29095,N_29096,N_29097,N_29098,N_29099,N_29100,N_29101,N_29102,N_29103,N_29104,N_29105,N_29106,N_29107,N_29108,N_29109,N_29110,N_29111,N_29112,N_29113,N_29114,N_29115,N_29116,N_29117,N_29118,N_29119,N_29120,N_29121,N_29122,N_29123,N_29124,N_29125,N_29126,N_29127,N_29128,N_29129,N_29130,N_29131,N_29132,N_29133,N_29134,N_29135,N_29136,N_29137,N_29138,N_29139,N_29140,N_29141,N_29142,N_29143,N_29144,N_29145,N_29146,N_29147,N_29148,N_29149,N_29150,N_29151,N_29152,N_29153,N_29154,N_29155,N_29156,N_29157,N_29158,N_29159,N_29160,N_29161,N_29162,N_29163,N_29164,N_29165,N_29166,N_29167,N_29168,N_29169,N_29170,N_29171,N_29172,N_29173,N_29174,N_29175,N_29176,N_29177,N_29178,N_29179,N_29180,N_29181,N_29182,N_29183,N_29184,N_29185,N_29186,N_29187,N_29188,N_29189,N_29190,N_29191,N_29192,N_29193,N_29194,N_29195,N_29196,N_29197,N_29198,N_29199,N_29200,N_29201,N_29202,N_29203,N_29204,N_29205,N_29206,N_29207,N_29208,N_29209,N_29210,N_29211,N_29212,N_29213,N_29214,N_29215,N_29216,N_29217,N_29218,N_29219,N_29220,N_29221,N_29222,N_29223,N_29224,N_29225,N_29226,N_29227,N_29228,N_29229,N_29230,N_29231,N_29232,N_29233,N_29234,N_29235,N_29236,N_29237,N_29238,N_29239,N_29240,N_29241,N_29242,N_29243,N_29244,N_29245,N_29246,N_29247,N_29248,N_29249,N_29250,N_29251,N_29252,N_29253,N_29254,N_29255,N_29256,N_29257,N_29258,N_29259,N_29260,N_29261,N_29262,N_29263,N_29264,N_29265,N_29266,N_29267,N_29268,N_29269,N_29270,N_29271,N_29272,N_29273,N_29274,N_29275,N_29276,N_29277,N_29278,N_29279,N_29280,N_29281,N_29282,N_29283,N_29284,N_29285,N_29286,N_29287,N_29288,N_29289,N_29290,N_29291,N_29292,N_29293,N_29294,N_29295,N_29296,N_29297,N_29298,N_29299,N_29300,N_29301,N_29302,N_29303,N_29304,N_29305,N_29306,N_29307,N_29308,N_29309,N_29310,N_29311,N_29312,N_29313,N_29314,N_29315,N_29316,N_29317,N_29318,N_29319,N_29320,N_29321,N_29322,N_29323,N_29324,N_29325,N_29326,N_29327,N_29328,N_29329,N_29330,N_29331,N_29332,N_29333,N_29334,N_29335,N_29336,N_29337,N_29338,N_29339,N_29340,N_29341,N_29342,N_29343,N_29344,N_29345,N_29346,N_29347,N_29348,N_29349,N_29350,N_29351,N_29352,N_29353,N_29354,N_29355,N_29356,N_29357,N_29358,N_29359,N_29360,N_29361,N_29362,N_29363,N_29364,N_29365,N_29366,N_29367,N_29368,N_29369,N_29370,N_29371,N_29372,N_29373,N_29374,N_29375,N_29376,N_29377,N_29378,N_29379,N_29380,N_29381,N_29382,N_29383,N_29384,N_29385,N_29386,N_29387,N_29388,N_29389,N_29390,N_29391,N_29392,N_29393,N_29394,N_29395,N_29396,N_29397,N_29398,N_29399,N_29400,N_29401,N_29402,N_29403,N_29404,N_29405,N_29406,N_29407,N_29408,N_29409,N_29410,N_29411,N_29412,N_29413,N_29414,N_29415,N_29416,N_29417,N_29418,N_29419,N_29420,N_29421,N_29422,N_29423,N_29424,N_29425,N_29426,N_29427,N_29428,N_29429,N_29430,N_29431,N_29432,N_29433,N_29434,N_29435,N_29436,N_29437,N_29438,N_29439,N_29440,N_29441,N_29442,N_29443,N_29444,N_29445,N_29446,N_29447,N_29448,N_29449,N_29450,N_29451,N_29452,N_29453,N_29454,N_29455,N_29456,N_29457,N_29458,N_29459,N_29460,N_29461,N_29462,N_29463,N_29464,N_29465,N_29466,N_29467,N_29468,N_29469,N_29470,N_29471,N_29472,N_29473,N_29474,N_29475,N_29476,N_29477,N_29478,N_29479,N_29480,N_29481,N_29482,N_29483,N_29484,N_29485,N_29486,N_29487,N_29488,N_29489,N_29490,N_29491,N_29492,N_29493,N_29494,N_29495,N_29496,N_29497,N_29498,N_29499,N_29500,N_29501,N_29502,N_29503,N_29504,N_29505,N_29506,N_29507,N_29508,N_29509,N_29510,N_29511,N_29512,N_29513,N_29514,N_29515,N_29516,N_29517,N_29518,N_29519,N_29520,N_29521,N_29522,N_29523,N_29524,N_29525,N_29526,N_29527,N_29528,N_29529,N_29530,N_29531,N_29532,N_29533,N_29534,N_29535,N_29536,N_29537,N_29538,N_29539,N_29540,N_29541,N_29542,N_29543,N_29544,N_29545,N_29546,N_29547,N_29548,N_29549,N_29550,N_29551,N_29552,N_29553,N_29554,N_29555,N_29556,N_29557,N_29558,N_29559,N_29560,N_29561,N_29562,N_29563,N_29564,N_29565,N_29566,N_29567,N_29568,N_29569,N_29570,N_29571,N_29572,N_29573,N_29574,N_29575,N_29576,N_29577,N_29578,N_29579,N_29580,N_29581,N_29582,N_29583,N_29584,N_29585,N_29586,N_29587,N_29588,N_29589,N_29590,N_29591,N_29592,N_29593,N_29594,N_29595,N_29596,N_29597,N_29598,N_29599,N_29600,N_29601,N_29602,N_29603,N_29604,N_29605,N_29606,N_29607,N_29608,N_29609,N_29610,N_29611,N_29612,N_29613,N_29614,N_29615,N_29616,N_29617,N_29618,N_29619,N_29620,N_29621,N_29622,N_29623,N_29624,N_29625,N_29626,N_29627,N_29628,N_29629,N_29630,N_29631,N_29632,N_29633,N_29634,N_29635,N_29636,N_29637,N_29638,N_29639,N_29640,N_29641,N_29642,N_29643,N_29644,N_29645,N_29646,N_29647,N_29648,N_29649,N_29650,N_29651,N_29652,N_29653,N_29654,N_29655,N_29656,N_29657,N_29658,N_29659,N_29660,N_29661,N_29662,N_29663,N_29664,N_29665,N_29666,N_29667,N_29668,N_29669,N_29670,N_29671,N_29672,N_29673,N_29674,N_29675,N_29676,N_29677,N_29678,N_29679,N_29680,N_29681,N_29682,N_29683,N_29684,N_29685,N_29686,N_29687,N_29688,N_29689,N_29690,N_29691,N_29692,N_29693,N_29694,N_29695,N_29696,N_29697,N_29698,N_29699,N_29700,N_29701,N_29702,N_29703,N_29704,N_29705,N_29706,N_29707,N_29708,N_29709,N_29710,N_29711,N_29712,N_29713,N_29714,N_29715,N_29716,N_29717,N_29718,N_29719,N_29720,N_29721,N_29722,N_29723,N_29724,N_29725,N_29726,N_29727,N_29728,N_29729,N_29730,N_29731,N_29732,N_29733,N_29734,N_29735,N_29736,N_29737,N_29738,N_29739,N_29740,N_29741,N_29742,N_29743,N_29744,N_29745,N_29746,N_29747,N_29748,N_29749,N_29750,N_29751,N_29752,N_29753,N_29754,N_29755,N_29756,N_29757,N_29758,N_29759,N_29760,N_29761,N_29762,N_29763,N_29764,N_29765,N_29766,N_29767,N_29768,N_29769,N_29770,N_29771,N_29772,N_29773,N_29774,N_29775,N_29776,N_29777,N_29778,N_29779,N_29780,N_29781,N_29782,N_29783,N_29784,N_29785,N_29786,N_29787,N_29788,N_29789,N_29790,N_29791,N_29792,N_29793,N_29794,N_29795,N_29796,N_29797,N_29798,N_29799,N_29800,N_29801,N_29802,N_29803,N_29804,N_29805,N_29806,N_29807,N_29808,N_29809,N_29810,N_29811,N_29812,N_29813,N_29814,N_29815,N_29816,N_29817,N_29818,N_29819,N_29820,N_29821,N_29822,N_29823,N_29824,N_29825,N_29826,N_29827,N_29828,N_29829,N_29830,N_29831,N_29832,N_29833,N_29834,N_29835,N_29836,N_29837,N_29838,N_29839,N_29840,N_29841,N_29842,N_29843,N_29844,N_29845,N_29846,N_29847,N_29848,N_29849,N_29850,N_29851,N_29852,N_29853,N_29854,N_29855,N_29856,N_29857,N_29858,N_29859,N_29860,N_29861,N_29862,N_29863,N_29864,N_29865,N_29866,N_29867,N_29868,N_29869,N_29870,N_29871,N_29872,N_29873,N_29874,N_29875,N_29876,N_29877,N_29878,N_29879,N_29880,N_29881,N_29882,N_29883,N_29884,N_29885,N_29886,N_29887,N_29888,N_29889,N_29890,N_29891,N_29892,N_29893,N_29894,N_29895,N_29896,N_29897,N_29898,N_29899,N_29900,N_29901,N_29902,N_29903,N_29904,N_29905,N_29906,N_29907,N_29908,N_29909,N_29910,N_29911,N_29912,N_29913,N_29914,N_29915,N_29916,N_29917,N_29918,N_29919,N_29920,N_29921,N_29922,N_29923,N_29924,N_29925,N_29926,N_29927,N_29928,N_29929,N_29930,N_29931,N_29932,N_29933,N_29934,N_29935,N_29936,N_29937,N_29938,N_29939,N_29940,N_29941,N_29942,N_29943,N_29944,N_29945,N_29946,N_29947,N_29948,N_29949,N_29950,N_29951,N_29952,N_29953,N_29954,N_29955,N_29956,N_29957,N_29958,N_29959,N_29960,N_29961,N_29962,N_29963,N_29964,N_29965,N_29966,N_29967,N_29968,N_29969,N_29970,N_29971,N_29972,N_29973,N_29974,N_29975,N_29976,N_29977,N_29978,N_29979,N_29980,N_29981,N_29982,N_29983,N_29984,N_29985,N_29986,N_29987,N_29988,N_29989,N_29990,N_29991,N_29992,N_29993,N_29994,N_29995,N_29996,N_29997,N_29998,N_29999,N_30000,N_30001,N_30002,N_30003,N_30004,N_30005,N_30006,N_30007,N_30008,N_30009,N_30010,N_30011,N_30012,N_30013,N_30014,N_30015,N_30016,N_30017,N_30018,N_30019,N_30020,N_30021,N_30022,N_30023,N_30024,N_30025,N_30026,N_30027,N_30028,N_30029,N_30030,N_30031,N_30032,N_30033,N_30034,N_30035,N_30036,N_30037,N_30038,N_30039,N_30040,N_30041,N_30042,N_30043,N_30044,N_30045,N_30046,N_30047,N_30048,N_30049,N_30050,N_30051,N_30052,N_30053,N_30054,N_30055,N_30056,N_30057,N_30058,N_30059,N_30060,N_30061,N_30062,N_30063,N_30064,N_30065,N_30066,N_30067,N_30068,N_30069,N_30070,N_30071,N_30072,N_30073,N_30074,N_30075,N_30076,N_30077,N_30078,N_30079,N_30080,N_30081,N_30082,N_30083,N_30084,N_30085,N_30086,N_30087,N_30088,N_30089,N_30090,N_30091,N_30092,N_30093,N_30094,N_30095,N_30096,N_30097,N_30098,N_30099,N_30100,N_30101,N_30102,N_30103,N_30104,N_30105,N_30106,N_30107,N_30108,N_30109,N_30110,N_30111,N_30112,N_30113,N_30114,N_30115,N_30116,N_30117,N_30118,N_30119,N_30120,N_30121,N_30122,N_30123,N_30124,N_30125,N_30126,N_30127,N_30128,N_30129,N_30130,N_30131,N_30132,N_30133,N_30134,N_30135,N_30136,N_30137,N_30138,N_30139,N_30140,N_30141,N_30142,N_30143,N_30144,N_30145,N_30146,N_30147,N_30148,N_30149,N_30150,N_30151,N_30152,N_30153,N_30154,N_30155,N_30156,N_30157,N_30158,N_30159,N_30160,N_30161,N_30162,N_30163,N_30164,N_30165,N_30166,N_30167,N_30168,N_30169,N_30170,N_30171,N_30172,N_30173,N_30174,N_30175,N_30176,N_30177,N_30178,N_30179,N_30180,N_30181,N_30182,N_30183,N_30184,N_30185,N_30186,N_30187,N_30188,N_30189,N_30190,N_30191,N_30192,N_30193,N_30194,N_30195,N_30196,N_30197,N_30198,N_30199,N_30200,N_30201,N_30202,N_30203,N_30204,N_30205,N_30206,N_30207,N_30208,N_30209,N_30210,N_30211,N_30212,N_30213,N_30214,N_30215,N_30216,N_30217,N_30218,N_30219,N_30220,N_30221,N_30222,N_30223,N_30224,N_30225,N_30226,N_30227,N_30228,N_30229,N_30230,N_30231,N_30232,N_30233,N_30234,N_30235,N_30236,N_30237,N_30238,N_30239,N_30240,N_30241,N_30242,N_30243,N_30244,N_30245,N_30246,N_30247,N_30248,N_30249,N_30250,N_30251,N_30252,N_30253,N_30254,N_30255,N_30256,N_30257,N_30258,N_30259,N_30260,N_30261,N_30262,N_30263,N_30264,N_30265,N_30266,N_30267,N_30268,N_30269,N_30270,N_30271,N_30272,N_30273,N_30274,N_30275,N_30276,N_30277,N_30278,N_30279,N_30280,N_30281,N_30282,N_30283,N_30284,N_30285,N_30286,N_30287,N_30288,N_30289,N_30290,N_30291,N_30292,N_30293,N_30294,N_30295,N_30296,N_30297,N_30298,N_30299,N_30300,N_30301,N_30302,N_30303,N_30304,N_30305,N_30306,N_30307,N_30308,N_30309,N_30310,N_30311,N_30312,N_30313,N_30314,N_30315,N_30316,N_30317,N_30318,N_30319,N_30320,N_30321,N_30322,N_30323,N_30324,N_30325,N_30326,N_30327,N_30328,N_30329,N_30330,N_30331,N_30332,N_30333,N_30334,N_30335,N_30336,N_30337,N_30338,N_30339,N_30340,N_30341,N_30342,N_30343,N_30344,N_30345,N_30346,N_30347,N_30348,N_30349,N_30350,N_30351,N_30352,N_30353,N_30354,N_30355,N_30356,N_30357,N_30358,N_30359,N_30360,N_30361,N_30362,N_30363,N_30364,N_30365,N_30366,N_30367,N_30368,N_30369,N_30370,N_30371,N_30372,N_30373,N_30374,N_30375,N_30376,N_30377,N_30378,N_30379,N_30380,N_30381,N_30382,N_30383,N_30384,N_30385,N_30386,N_30387,N_30388,N_30389,N_30390,N_30391,N_30392,N_30393,N_30394,N_30395,N_30396,N_30397,N_30398,N_30399,N_30400,N_30401,N_30402,N_30403,N_30404,N_30405,N_30406,N_30407,N_30408,N_30409,N_30410,N_30411,N_30412,N_30413,N_30414,N_30415,N_30416,N_30417,N_30418,N_30419,N_30420,N_30421,N_30422,N_30423,N_30424,N_30425,N_30426,N_30427,N_30428,N_30429,N_30430,N_30431,N_30432,N_30433,N_30434,N_30435,N_30436,N_30437,N_30438,N_30439,N_30440,N_30441,N_30442,N_30443,N_30444,N_30445,N_30446,N_30447,N_30448,N_30449,N_30450,N_30451,N_30452,N_30453,N_30454,N_30455,N_30456,N_30457,N_30458,N_30459,N_30460,N_30461,N_30462,N_30463,N_30464,N_30465,N_30466,N_30467,N_30468,N_30469,N_30470,N_30471,N_30472,N_30473,N_30474,N_30475,N_30476,N_30477,N_30478,N_30479,N_30480,N_30481,N_30482,N_30483,N_30484,N_30485,N_30486,N_30487,N_30488,N_30489,N_30490,N_30491,N_30492,N_30493,N_30494,N_30495,N_30496,N_30497,N_30498,N_30499,N_30500,N_30501,N_30502,N_30503,N_30504,N_30505,N_30506,N_30507,N_30508,N_30509,N_30510,N_30511,N_30512,N_30513,N_30514,N_30515,N_30516,N_30517,N_30518,N_30519,N_30520,N_30521,N_30522,N_30523,N_30524,N_30525,N_30526,N_30527,N_30528,N_30529,N_30530,N_30531,N_30532,N_30533,N_30534,N_30535,N_30536,N_30537,N_30538,N_30539,N_30540,N_30541,N_30542,N_30543,N_30544,N_30545,N_30546,N_30547,N_30548,N_30549,N_30550,N_30551,N_30552,N_30553,N_30554,N_30555,N_30556,N_30557,N_30558,N_30559,N_30560,N_30561,N_30562,N_30563,N_30564,N_30565,N_30566,N_30567,N_30568,N_30569,N_30570,N_30571,N_30572,N_30573,N_30574,N_30575,N_30576,N_30577,N_30578,N_30579,N_30580,N_30581,N_30582,N_30583,N_30584,N_30585,N_30586,N_30587,N_30588,N_30589,N_30590,N_30591,N_30592,N_30593,N_30594,N_30595,N_30596,N_30597,N_30598,N_30599,N_30600,N_30601,N_30602,N_30603,N_30604,N_30605,N_30606,N_30607,N_30608,N_30609,N_30610,N_30611,N_30612,N_30613,N_30614,N_30615,N_30616,N_30617,N_30618,N_30619,N_30620,N_30621,N_30622,N_30623,N_30624,N_30625,N_30626,N_30627,N_30628,N_30629,N_30630,N_30631,N_30632,N_30633,N_30634,N_30635,N_30636,N_30637,N_30638,N_30639,N_30640,N_30641,N_30642,N_30643,N_30644,N_30645,N_30646,N_30647,N_30648,N_30649,N_30650,N_30651,N_30652,N_30653,N_30654,N_30655,N_30656,N_30657,N_30658,N_30659,N_30660,N_30661,N_30662,N_30663,N_30664,N_30665,N_30666,N_30667,N_30668,N_30669,N_30670,N_30671,N_30672,N_30673,N_30674,N_30675,N_30676,N_30677,N_30678,N_30679,N_30680,N_30681,N_30682,N_30683,N_30684,N_30685,N_30686,N_30687,N_30688,N_30689,N_30690,N_30691,N_30692,N_30693,N_30694,N_30695,N_30696,N_30697,N_30698,N_30699,N_30700,N_30701,N_30702,N_30703,N_30704,N_30705,N_30706,N_30707,N_30708,N_30709,N_30710,N_30711,N_30712,N_30713,N_30714,N_30715,N_30716,N_30717,N_30718,N_30719,N_30720,N_30721,N_30722,N_30723,N_30724,N_30725,N_30726,N_30727,N_30728,N_30729,N_30730,N_30731,N_30732,N_30733,N_30734,N_30735,N_30736,N_30737,N_30738,N_30739,N_30740,N_30741,N_30742,N_30743,N_30744,N_30745,N_30746,N_30747,N_30748,N_30749,N_30750,N_30751,N_30752,N_30753,N_30754,N_30755,N_30756,N_30757,N_30758,N_30759,N_30760,N_30761,N_30762,N_30763,N_30764,N_30765,N_30766,N_30767,N_30768,N_30769,N_30770,N_30771,N_30772,N_30773,N_30774,N_30775,N_30776,N_30777,N_30778,N_30779,N_30780,N_30781,N_30782,N_30783,N_30784,N_30785,N_30786,N_30787,N_30788,N_30789,N_30790,N_30791,N_30792,N_30793,N_30794,N_30795,N_30796,N_30797,N_30798,N_30799,N_30800,N_30801,N_30802,N_30803,N_30804,N_30805,N_30806,N_30807,N_30808,N_30809,N_30810,N_30811,N_30812,N_30813,N_30814,N_30815,N_30816,N_30817,N_30818,N_30819,N_30820,N_30821,N_30822,N_30823,N_30824,N_30825,N_30826,N_30827,N_30828,N_30829,N_30830,N_30831,N_30832,N_30833,N_30834,N_30835,N_30836,N_30837,N_30838,N_30839,N_30840,N_30841,N_30842,N_30843,N_30844,N_30845,N_30846,N_30847,N_30848,N_30849,N_30850,N_30851,N_30852,N_30853,N_30854,N_30855,N_30856,N_30857,N_30858,N_30859,N_30860,N_30861,N_30862,N_30863,N_30864,N_30865,N_30866,N_30867,N_30868,N_30869,N_30870,N_30871,N_30872,N_30873,N_30874,N_30875,N_30876,N_30877,N_30878,N_30879,N_30880,N_30881,N_30882,N_30883,N_30884,N_30885,N_30886,N_30887,N_30888,N_30889,N_30890,N_30891,N_30892,N_30893,N_30894,N_30895,N_30896,N_30897,N_30898,N_30899,N_30900,N_30901,N_30902,N_30903,N_30904,N_30905,N_30906,N_30907,N_30908,N_30909,N_30910,N_30911,N_30912,N_30913,N_30914,N_30915,N_30916,N_30917,N_30918,N_30919,N_30920,N_30921,N_30922,N_30923,N_30924,N_30925,N_30926,N_30927,N_30928,N_30929,N_30930,N_30931,N_30932,N_30933,N_30934,N_30935,N_30936,N_30937,N_30938,N_30939,N_30940,N_30941,N_30942,N_30943,N_30944,N_30945,N_30946,N_30947,N_30948,N_30949,N_30950,N_30951,N_30952,N_30953,N_30954,N_30955,N_30956,N_30957,N_30958,N_30959,N_30960,N_30961,N_30962,N_30963,N_30964,N_30965,N_30966,N_30967,N_30968,N_30969,N_30970,N_30971,N_30972,N_30973,N_30974,N_30975,N_30976,N_30977,N_30978,N_30979,N_30980,N_30981,N_30982,N_30983,N_30984,N_30985,N_30986,N_30987,N_30988,N_30989,N_30990,N_30991,N_30992,N_30993,N_30994,N_30995,N_30996,N_30997,N_30998,N_30999,N_31000,N_31001,N_31002,N_31003,N_31004,N_31005,N_31006,N_31007,N_31008,N_31009,N_31010,N_31011,N_31012,N_31013,N_31014,N_31015,N_31016,N_31017,N_31018,N_31019,N_31020,N_31021,N_31022,N_31023,N_31024,N_31025,N_31026,N_31027,N_31028,N_31029,N_31030,N_31031,N_31032,N_31033,N_31034,N_31035,N_31036,N_31037,N_31038,N_31039,N_31040,N_31041,N_31042,N_31043,N_31044,N_31045,N_31046,N_31047,N_31048,N_31049,N_31050,N_31051,N_31052,N_31053,N_31054,N_31055,N_31056,N_31057,N_31058,N_31059,N_31060,N_31061,N_31062,N_31063,N_31064,N_31065,N_31066,N_31067,N_31068,N_31069,N_31070,N_31071,N_31072,N_31073,N_31074,N_31075,N_31076,N_31077,N_31078,N_31079,N_31080,N_31081,N_31082,N_31083,N_31084,N_31085,N_31086,N_31087,N_31088,N_31089,N_31090,N_31091,N_31092,N_31093,N_31094,N_31095,N_31096,N_31097,N_31098,N_31099,N_31100,N_31101,N_31102,N_31103,N_31104,N_31105,N_31106,N_31107,N_31108,N_31109,N_31110,N_31111,N_31112,N_31113,N_31114,N_31115,N_31116,N_31117,N_31118,N_31119,N_31120,N_31121,N_31122,N_31123,N_31124,N_31125,N_31126,N_31127,N_31128,N_31129,N_31130,N_31131,N_31132,N_31133,N_31134,N_31135,N_31136,N_31137,N_31138,N_31139,N_31140,N_31141,N_31142,N_31143,N_31144,N_31145,N_31146,N_31147,N_31148,N_31149,N_31150,N_31151,N_31152,N_31153,N_31154,N_31155,N_31156,N_31157,N_31158,N_31159,N_31160,N_31161,N_31162,N_31163,N_31164,N_31165,N_31166,N_31167,N_31168,N_31169,N_31170,N_31171,N_31172,N_31173,N_31174,N_31175,N_31176,N_31177,N_31178,N_31179,N_31180,N_31181,N_31182,N_31183,N_31184,N_31185,N_31186,N_31187,N_31188,N_31189,N_31190,N_31191,N_31192,N_31193,N_31194,N_31195,N_31196,N_31197,N_31198,N_31199,N_31200,N_31201,N_31202,N_31203,N_31204,N_31205,N_31206,N_31207,N_31208,N_31209,N_31210,N_31211,N_31212,N_31213,N_31214,N_31215,N_31216,N_31217,N_31218,N_31219,N_31220,N_31221,N_31222,N_31223,N_31224,N_31225,N_31226,N_31227,N_31228,N_31229,N_31230,N_31231,N_31232,N_31233,N_31234,N_31235,N_31236,N_31237,N_31238,N_31239,N_31240,N_31241,N_31242,N_31243,N_31244,N_31245,N_31246,N_31247,N_31248,N_31249,N_31250,N_31251,N_31252,N_31253,N_31254,N_31255,N_31256,N_31257,N_31258,N_31259,N_31260,N_31261,N_31262,N_31263,N_31264,N_31265,N_31266,N_31267,N_31268,N_31269,N_31270,N_31271,N_31272,N_31273,N_31274,N_31275,N_31276,N_31277,N_31278,N_31279,N_31280,N_31281,N_31282,N_31283,N_31284,N_31285,N_31286,N_31287,N_31288,N_31289,N_31290,N_31291,N_31292,N_31293,N_31294,N_31295,N_31296,N_31297,N_31298,N_31299,N_31300,N_31301,N_31302,N_31303,N_31304,N_31305,N_31306,N_31307,N_31308,N_31309,N_31310,N_31311,N_31312,N_31313,N_31314,N_31315,N_31316,N_31317,N_31318,N_31319,N_31320,N_31321,N_31322,N_31323,N_31324,N_31325,N_31326,N_31327,N_31328,N_31329,N_31330,N_31331,N_31332,N_31333,N_31334,N_31335,N_31336,N_31337,N_31338,N_31339,N_31340,N_31341,N_31342,N_31343,N_31344,N_31345,N_31346,N_31347,N_31348,N_31349,N_31350,N_31351,N_31352,N_31353,N_31354,N_31355,N_31356,N_31357,N_31358,N_31359,N_31360,N_31361,N_31362,N_31363,N_31364,N_31365,N_31366,N_31367,N_31368,N_31369,N_31370,N_31371,N_31372,N_31373,N_31374,N_31375,N_31376,N_31377,N_31378,N_31379,N_31380,N_31381,N_31382,N_31383,N_31384,N_31385,N_31386,N_31387,N_31388,N_31389,N_31390,N_31391,N_31392,N_31393,N_31394,N_31395,N_31396,N_31397,N_31398,N_31399,N_31400,N_31401,N_31402,N_31403,N_31404,N_31405,N_31406,N_31407,N_31408,N_31409,N_31410,N_31411,N_31412,N_31413,N_31414,N_31415,N_31416,N_31417,N_31418,N_31419,N_31420,N_31421,N_31422,N_31423,N_31424,N_31425,N_31426,N_31427,N_31428,N_31429,N_31430,N_31431,N_31432,N_31433,N_31434,N_31435,N_31436,N_31437,N_31438,N_31439,N_31440,N_31441,N_31442,N_31443,N_31444,N_31445,N_31446,N_31447,N_31448,N_31449,N_31450,N_31451,N_31452,N_31453,N_31454,N_31455,N_31456,N_31457,N_31458,N_31459,N_31460,N_31461,N_31462,N_31463,N_31464,N_31465,N_31466,N_31467,N_31468,N_31469,N_31470,N_31471,N_31472,N_31473,N_31474,N_31475,N_31476,N_31477,N_31478,N_31479,N_31480,N_31481,N_31482,N_31483,N_31484,N_31485,N_31486,N_31487,N_31488,N_31489,N_31490,N_31491,N_31492,N_31493,N_31494,N_31495,N_31496,N_31497,N_31498,N_31499,N_31500,N_31501,N_31502,N_31503,N_31504,N_31505,N_31506,N_31507,N_31508,N_31509,N_31510,N_31511,N_31512,N_31513,N_31514,N_31515,N_31516,N_31517,N_31518,N_31519,N_31520,N_31521,N_31522,N_31523,N_31524,N_31525,N_31526,N_31527,N_31528,N_31529,N_31530,N_31531,N_31532,N_31533,N_31534,N_31535,N_31536,N_31537,N_31538,N_31539,N_31540,N_31541,N_31542,N_31543,N_31544,N_31545,N_31546,N_31547,N_31548,N_31549,N_31550,N_31551,N_31552,N_31553,N_31554,N_31555,N_31556,N_31557,N_31558,N_31559,N_31560,N_31561,N_31562,N_31563,N_31564,N_31565,N_31566,N_31567,N_31568,N_31569,N_31570,N_31571,N_31572,N_31573,N_31574,N_31575,N_31576,N_31577,N_31578,N_31579,N_31580,N_31581,N_31582,N_31583,N_31584,N_31585,N_31586,N_31587,N_31588,N_31589,N_31590,N_31591,N_31592,N_31593,N_31594,N_31595,N_31596,N_31597,N_31598,N_31599,N_31600,N_31601,N_31602,N_31603,N_31604,N_31605,N_31606,N_31607,N_31608,N_31609,N_31610,N_31611,N_31612,N_31613,N_31614,N_31615,N_31616,N_31617,N_31618,N_31619,N_31620,N_31621,N_31622,N_31623,N_31624,N_31625,N_31626,N_31627,N_31628,N_31629,N_31630,N_31631,N_31632,N_31633,N_31634,N_31635,N_31636,N_31637,N_31638,N_31639,N_31640,N_31641,N_31642,N_31643,N_31644,N_31645,N_31646,N_31647,N_31648,N_31649,N_31650,N_31651,N_31652,N_31653,N_31654,N_31655,N_31656,N_31657,N_31658,N_31659,N_31660,N_31661,N_31662,N_31663,N_31664,N_31665,N_31666,N_31667,N_31668,N_31669,N_31670,N_31671,N_31672,N_31673,N_31674,N_31675,N_31676,N_31677,N_31678,N_31679,N_31680,N_31681,N_31682,N_31683,N_31684,N_31685,N_31686,N_31687,N_31688,N_31689,N_31690,N_31691,N_31692,N_31693,N_31694,N_31695,N_31696,N_31697,N_31698,N_31699,N_31700,N_31701,N_31702,N_31703,N_31704,N_31705,N_31706,N_31707,N_31708,N_31709,N_31710,N_31711,N_31712,N_31713,N_31714,N_31715,N_31716,N_31717,N_31718,N_31719,N_31720,N_31721,N_31722,N_31723,N_31724,N_31725,N_31726,N_31727,N_31728,N_31729,N_31730,N_31731,N_31732,N_31733,N_31734,N_31735,N_31736,N_31737,N_31738,N_31739,N_31740,N_31741,N_31742,N_31743,N_31744,N_31745,N_31746,N_31747,N_31748,N_31749,N_31750,N_31751,N_31752,N_31753,N_31754,N_31755,N_31756,N_31757,N_31758,N_31759,N_31760,N_31761,N_31762,N_31763,N_31764,N_31765,N_31766,N_31767,N_31768,N_31769,N_31770,N_31771,N_31772,N_31773,N_31774,N_31775,N_31776,N_31777,N_31778,N_31779,N_31780,N_31781,N_31782,N_31783,N_31784,N_31785,N_31786,N_31787,N_31788,N_31789,N_31790,N_31791,N_31792,N_31793,N_31794,N_31795,N_31796,N_31797,N_31798,N_31799,N_31800,N_31801,N_31802,N_31803,N_31804,N_31805,N_31806,N_31807,N_31808,N_31809,N_31810,N_31811,N_31812,N_31813,N_31814,N_31815,N_31816,N_31817,N_31818,N_31819,N_31820,N_31821,N_31822,N_31823,N_31824,N_31825,N_31826,N_31827,N_31828,N_31829,N_31830,N_31831,N_31832,N_31833,N_31834,N_31835,N_31836,N_31837,N_31838,N_31839,N_31840,N_31841,N_31842,N_31843,N_31844,N_31845,N_31846,N_31847,N_31848,N_31849,N_31850,N_31851,N_31852,N_31853,N_31854,N_31855,N_31856,N_31857,N_31858,N_31859,N_31860,N_31861,N_31862,N_31863,N_31864,N_31865,N_31866,N_31867,N_31868,N_31869,N_31870,N_31871,N_31872,N_31873,N_31874,N_31875,N_31876,N_31877,N_31878,N_31879,N_31880,N_31881,N_31882,N_31883,N_31884,N_31885,N_31886,N_31887,N_31888,N_31889,N_31890,N_31891,N_31892,N_31893,N_31894,N_31895,N_31896,N_31897,N_31898,N_31899,N_31900,N_31901,N_31902,N_31903,N_31904,N_31905,N_31906,N_31907,N_31908,N_31909,N_31910,N_31911,N_31912,N_31913,N_31914,N_31915,N_31916,N_31917,N_31918,N_31919,N_31920,N_31921,N_31922,N_31923,N_31924,N_31925,N_31926,N_31927,N_31928,N_31929,N_31930,N_31931,N_31932,N_31933,N_31934,N_31935,N_31936,N_31937,N_31938,N_31939,N_31940,N_31941,N_31942,N_31943,N_31944,N_31945,N_31946,N_31947,N_31948,N_31949,N_31950,N_31951,N_31952,N_31953,N_31954,N_31955,N_31956,N_31957,N_31958,N_31959,N_31960,N_31961,N_31962,N_31963,N_31964,N_31965,N_31966,N_31967,N_31968,N_31969,N_31970,N_31971,N_31972,N_31973,N_31974,N_31975,N_31976,N_31977,N_31978,N_31979,N_31980,N_31981,N_31982,N_31983,N_31984,N_31985,N_31986,N_31987,N_31988,N_31989,N_31990,N_31991,N_31992,N_31993,N_31994,N_31995,N_31996,N_31997,N_31998,N_31999,N_32000,N_32001,N_32002,N_32003,N_32004,N_32005,N_32006,N_32007,N_32008,N_32009,N_32010,N_32011,N_32012,N_32013,N_32014,N_32015,N_32016,N_32017,N_32018,N_32019,N_32020,N_32021,N_32022,N_32023,N_32024,N_32025,N_32026,N_32027,N_32028,N_32029,N_32030,N_32031,N_32032,N_32033,N_32034,N_32035,N_32036,N_32037,N_32038,N_32039,N_32040,N_32041,N_32042,N_32043,N_32044,N_32045,N_32046,N_32047,N_32048,N_32049,N_32050,N_32051,N_32052,N_32053,N_32054,N_32055,N_32056,N_32057,N_32058,N_32059,N_32060,N_32061,N_32062,N_32063,N_32064,N_32065,N_32066,N_32067,N_32068,N_32069,N_32070,N_32071,N_32072,N_32073,N_32074,N_32075,N_32076,N_32077,N_32078,N_32079,N_32080,N_32081,N_32082,N_32083,N_32084,N_32085,N_32086,N_32087,N_32088,N_32089,N_32090,N_32091,N_32092,N_32093,N_32094,N_32095,N_32096,N_32097,N_32098,N_32099,N_32100,N_32101,N_32102,N_32103,N_32104,N_32105,N_32106,N_32107,N_32108,N_32109,N_32110,N_32111,N_32112,N_32113,N_32114,N_32115,N_32116,N_32117,N_32118,N_32119,N_32120,N_32121,N_32122,N_32123,N_32124,N_32125,N_32126,N_32127,N_32128,N_32129,N_32130,N_32131,N_32132,N_32133,N_32134,N_32135,N_32136,N_32137,N_32138,N_32139,N_32140,N_32141,N_32142,N_32143,N_32144,N_32145,N_32146,N_32147,N_32148,N_32149,N_32150,N_32151,N_32152,N_32153,N_32154,N_32155,N_32156,N_32157,N_32158,N_32159,N_32160,N_32161,N_32162,N_32163,N_32164,N_32165,N_32166,N_32167,N_32168,N_32169,N_32170,N_32171,N_32172,N_32173,N_32174,N_32175,N_32176,N_32177,N_32178,N_32179,N_32180,N_32181,N_32182,N_32183,N_32184,N_32185,N_32186,N_32187,N_32188,N_32189,N_32190,N_32191,N_32192,N_32193,N_32194,N_32195,N_32196,N_32197,N_32198,N_32199,N_32200,N_32201,N_32202,N_32203,N_32204,N_32205,N_32206,N_32207,N_32208,N_32209,N_32210,N_32211,N_32212,N_32213,N_32214,N_32215,N_32216,N_32217,N_32218,N_32219,N_32220,N_32221,N_32222,N_32223,N_32224,N_32225,N_32226,N_32227,N_32228,N_32229,N_32230,N_32231,N_32232,N_32233,N_32234,N_32235,N_32236,N_32237,N_32238,N_32239,N_32240,N_32241,N_32242,N_32243,N_32244,N_32245,N_32246,N_32247,N_32248,N_32249,N_32250,N_32251,N_32252,N_32253,N_32254,N_32255,N_32256,N_32257,N_32258,N_32259,N_32260,N_32261,N_32262,N_32263,N_32264,N_32265,N_32266,N_32267,N_32268,N_32269,N_32270,N_32271,N_32272,N_32273,N_32274,N_32275,N_32276,N_32277,N_32278,N_32279,N_32280,N_32281,N_32282,N_32283,N_32284,N_32285,N_32286,N_32287,N_32288,N_32289,N_32290,N_32291,N_32292,N_32293,N_32294,N_32295,N_32296,N_32297,N_32298,N_32299,N_32300,N_32301,N_32302,N_32303,N_32304,N_32305,N_32306,N_32307,N_32308,N_32309,N_32310,N_32311,N_32312,N_32313,N_32314,N_32315,N_32316,N_32317,N_32318,N_32319,N_32320,N_32321,N_32322,N_32323,N_32324,N_32325,N_32326,N_32327,N_32328,N_32329,N_32330,N_32331,N_32332,N_32333,N_32334,N_32335,N_32336,N_32337,N_32338,N_32339,N_32340,N_32341,N_32342,N_32343,N_32344,N_32345,N_32346,N_32347,N_32348,N_32349,N_32350,N_32351,N_32352,N_32353,N_32354,N_32355,N_32356,N_32357,N_32358,N_32359,N_32360,N_32361,N_32362,N_32363,N_32364,N_32365,N_32366,N_32367,N_32368,N_32369,N_32370,N_32371,N_32372,N_32373,N_32374,N_32375,N_32376,N_32377,N_32378,N_32379,N_32380,N_32381,N_32382,N_32383,N_32384,N_32385,N_32386,N_32387,N_32388,N_32389,N_32390,N_32391,N_32392,N_32393,N_32394,N_32395,N_32396,N_32397,N_32398,N_32399,N_32400,N_32401,N_32402,N_32403,N_32404,N_32405,N_32406,N_32407,N_32408,N_32409,N_32410,N_32411,N_32412,N_32413,N_32414,N_32415,N_32416,N_32417,N_32418,N_32419,N_32420,N_32421,N_32422,N_32423,N_32424,N_32425,N_32426,N_32427,N_32428,N_32429,N_32430,N_32431,N_32432,N_32433,N_32434,N_32435,N_32436,N_32437,N_32438,N_32439,N_32440,N_32441,N_32442,N_32443,N_32444,N_32445,N_32446,N_32447,N_32448,N_32449,N_32450,N_32451,N_32452,N_32453,N_32454,N_32455,N_32456,N_32457,N_32458,N_32459,N_32460,N_32461,N_32462,N_32463,N_32464,N_32465,N_32466,N_32467,N_32468,N_32469,N_32470,N_32471,N_32472,N_32473,N_32474,N_32475,N_32476,N_32477,N_32478,N_32479,N_32480,N_32481,N_32482,N_32483,N_32484,N_32485,N_32486,N_32487,N_32488,N_32489,N_32490,N_32491,N_32492,N_32493,N_32494,N_32495,N_32496,N_32497,N_32498,N_32499,N_32500,N_32501,N_32502,N_32503,N_32504,N_32505,N_32506,N_32507,N_32508,N_32509,N_32510,N_32511,N_32512,N_32513,N_32514,N_32515,N_32516,N_32517,N_32518,N_32519,N_32520,N_32521,N_32522,N_32523,N_32524,N_32525,N_32526,N_32527,N_32528,N_32529,N_32530,N_32531,N_32532,N_32533,N_32534,N_32535,N_32536,N_32537,N_32538,N_32539,N_32540,N_32541,N_32542,N_32543,N_32544,N_32545,N_32546,N_32547,N_32548,N_32549,N_32550,N_32551,N_32552,N_32553,N_32554,N_32555,N_32556,N_32557,N_32558,N_32559,N_32560,N_32561,N_32562,N_32563,N_32564,N_32565,N_32566,N_32567,N_32568,N_32569,N_32570,N_32571,N_32572,N_32573,N_32574,N_32575,N_32576,N_32577,N_32578,N_32579,N_32580,N_32581,N_32582,N_32583,N_32584,N_32585,N_32586,N_32587,N_32588,N_32589,N_32590,N_32591,N_32592,N_32593,N_32594,N_32595,N_32596,N_32597,N_32598,N_32599,N_32600,N_32601,N_32602,N_32603,N_32604,N_32605,N_32606,N_32607,N_32608,N_32609,N_32610,N_32611,N_32612,N_32613,N_32614,N_32615,N_32616,N_32617,N_32618,N_32619,N_32620,N_32621,N_32622,N_32623,N_32624,N_32625,N_32626,N_32627,N_32628,N_32629,N_32630,N_32631,N_32632,N_32633,N_32634,N_32635,N_32636,N_32637,N_32638,N_32639,N_32640,N_32641,N_32642,N_32643,N_32644,N_32645,N_32646,N_32647,N_32648,N_32649,N_32650,N_32651,N_32652,N_32653,N_32654,N_32655,N_32656,N_32657,N_32658,N_32659,N_32660,N_32661,N_32662,N_32663,N_32664,N_32665,N_32666,N_32667,N_32668,N_32669,N_32670,N_32671,N_32672,N_32673,N_32674,N_32675,N_32676,N_32677,N_32678,N_32679,N_32680,N_32681,N_32682,N_32683,N_32684,N_32685,N_32686,N_32687,N_32688,N_32689,N_32690,N_32691,N_32692,N_32693,N_32694,N_32695,N_32696,N_32697,N_32698,N_32699,N_32700,N_32701,N_32702,N_32703,N_32704,N_32705,N_32706,N_32707,N_32708,N_32709,N_32710,N_32711,N_32712,N_32713,N_32714,N_32715,N_32716,N_32717,N_32718,N_32719,N_32720,N_32721,N_32722,N_32723,N_32724,N_32725,N_32726,N_32727,N_32728,N_32729,N_32730,N_32731,N_32732,N_32733,N_32734,N_32735,N_32736,N_32737,N_32738,N_32739,N_32740,N_32741,N_32742,N_32743,N_32744,N_32745,N_32746,N_32747,N_32748,N_32749,N_32750,N_32751,N_32752,N_32753,N_32754,N_32755,N_32756,N_32757,N_32758,N_32759,N_32760,N_32761,N_32762,N_32763,N_32764,N_32765,N_32766,N_32767,N_32768,N_32769,N_32770,N_32771,N_32772,N_32773,N_32774,N_32775,N_32776,N_32777,N_32778,N_32779,N_32780,N_32781,N_32782,N_32783,N_32784,N_32785,N_32786,N_32787,N_32788,N_32789,N_32790,N_32791,N_32792,N_32793,N_32794,N_32795,N_32796,N_32797,N_32798,N_32799,N_32800,N_32801,N_32802,N_32803,N_32804,N_32805,N_32806,N_32807,N_32808,N_32809,N_32810,N_32811,N_32812,N_32813,N_32814,N_32815,N_32816,N_32817,N_32818,N_32819,N_32820,N_32821,N_32822,N_32823,N_32824,N_32825,N_32826,N_32827,N_32828,N_32829,N_32830,N_32831,N_32832,N_32833,N_32834,N_32835,N_32836,N_32837,N_32838,N_32839,N_32840,N_32841,N_32842,N_32843,N_32844,N_32845,N_32846,N_32847,N_32848,N_32849,N_32850,N_32851,N_32852,N_32853,N_32854,N_32855,N_32856,N_32857,N_32858,N_32859,N_32860,N_32861,N_32862,N_32863,N_32864,N_32865,N_32866,N_32867,N_32868,N_32869,N_32870,N_32871,N_32872,N_32873,N_32874,N_32875,N_32876,N_32877,N_32878,N_32879,N_32880,N_32881,N_32882,N_32883,N_32884,N_32885,N_32886,N_32887,N_32888,N_32889,N_32890,N_32891,N_32892,N_32893,N_32894,N_32895,N_32896,N_32897,N_32898,N_32899,N_32900,N_32901,N_32902,N_32903,N_32904,N_32905,N_32906,N_32907,N_32908,N_32909,N_32910,N_32911,N_32912,N_32913,N_32914,N_32915,N_32916,N_32917,N_32918,N_32919,N_32920,N_32921,N_32922,N_32923,N_32924,N_32925,N_32926,N_32927,N_32928,N_32929,N_32930,N_32931,N_32932,N_32933,N_32934,N_32935,N_32936,N_32937,N_32938,N_32939,N_32940,N_32941,N_32942,N_32943,N_32944,N_32945,N_32946,N_32947,N_32948,N_32949,N_32950,N_32951,N_32952,N_32953,N_32954,N_32955,N_32956,N_32957,N_32958,N_32959,N_32960,N_32961,N_32962,N_32963,N_32964,N_32965,N_32966,N_32967,N_32968,N_32969,N_32970,N_32971,N_32972,N_32973,N_32974,N_32975,N_32976,N_32977,N_32978,N_32979,N_32980,N_32981,N_32982,N_32983,N_32984,N_32985,N_32986,N_32987,N_32988,N_32989,N_32990,N_32991,N_32992,N_32993,N_32994,N_32995,N_32996,N_32997,N_32998,N_32999,N_33000,N_33001,N_33002,N_33003,N_33004,N_33005,N_33006,N_33007,N_33008,N_33009,N_33010,N_33011,N_33012,N_33013,N_33014,N_33015,N_33016,N_33017,N_33018,N_33019,N_33020,N_33021,N_33022,N_33023,N_33024,N_33025,N_33026,N_33027,N_33028,N_33029,N_33030,N_33031,N_33032,N_33033,N_33034,N_33035,N_33036,N_33037,N_33038,N_33039,N_33040,N_33041,N_33042,N_33043,N_33044,N_33045,N_33046,N_33047,N_33048,N_33049,N_33050,N_33051,N_33052,N_33053,N_33054,N_33055,N_33056,N_33057,N_33058,N_33059,N_33060,N_33061,N_33062,N_33063,N_33064,N_33065,N_33066,N_33067,N_33068,N_33069,N_33070,N_33071,N_33072,N_33073,N_33074,N_33075,N_33076,N_33077,N_33078,N_33079,N_33080,N_33081,N_33082,N_33083,N_33084,N_33085,N_33086,N_33087,N_33088,N_33089,N_33090,N_33091,N_33092,N_33093,N_33094,N_33095,N_33096,N_33097,N_33098,N_33099,N_33100,N_33101,N_33102,N_33103,N_33104,N_33105,N_33106,N_33107,N_33108,N_33109,N_33110,N_33111,N_33112,N_33113,N_33114,N_33115,N_33116,N_33117,N_33118,N_33119,N_33120,N_33121,N_33122,N_33123,N_33124,N_33125,N_33126,N_33127,N_33128,N_33129,N_33130,N_33131,N_33132,N_33133,N_33134,N_33135,N_33136,N_33137,N_33138,N_33139,N_33140,N_33141,N_33142,N_33143,N_33144,N_33145,N_33146,N_33147,N_33148,N_33149,N_33150,N_33151,N_33152,N_33153,N_33154,N_33155,N_33156,N_33157,N_33158,N_33159,N_33160,N_33161,N_33162,N_33163,N_33164,N_33165,N_33166,N_33167,N_33168,N_33169,N_33170,N_33171,N_33172,N_33173,N_33174,N_33175,N_33176,N_33177,N_33178,N_33179,N_33180,N_33181,N_33182,N_33183,N_33184,N_33185,N_33186,N_33187,N_33188,N_33189,N_33190,N_33191,N_33192,N_33193,N_33194,N_33195,N_33196,N_33197,N_33198,N_33199,N_33200,N_33201,N_33202,N_33203,N_33204,N_33205,N_33206,N_33207,N_33208,N_33209,N_33210,N_33211,N_33212,N_33213,N_33214,N_33215,N_33216,N_33217,N_33218,N_33219,N_33220,N_33221,N_33222,N_33223,N_33224,N_33225,N_33226,N_33227,N_33228,N_33229,N_33230,N_33231,N_33232,N_33233,N_33234,N_33235,N_33236,N_33237,N_33238,N_33239,N_33240,N_33241,N_33242,N_33243,N_33244,N_33245,N_33246,N_33247,N_33248,N_33249,N_33250,N_33251,N_33252,N_33253,N_33254,N_33255,N_33256,N_33257,N_33258,N_33259,N_33260,N_33261,N_33262,N_33263,N_33264,N_33265,N_33266,N_33267,N_33268,N_33269,N_33270,N_33271,N_33272,N_33273,N_33274,N_33275,N_33276,N_33277,N_33278,N_33279,N_33280,N_33281,N_33282,N_33283,N_33284,N_33285,N_33286,N_33287,N_33288,N_33289,N_33290,N_33291,N_33292,N_33293,N_33294,N_33295,N_33296,N_33297,N_33298,N_33299,N_33300,N_33301,N_33302,N_33303,N_33304,N_33305,N_33306,N_33307,N_33308,N_33309,N_33310,N_33311,N_33312,N_33313,N_33314,N_33315,N_33316,N_33317,N_33318,N_33319,N_33320,N_33321,N_33322,N_33323,N_33324,N_33325,N_33326,N_33327,N_33328,N_33329,N_33330,N_33331,N_33332,N_33333,N_33334,N_33335,N_33336,N_33337,N_33338,N_33339,N_33340,N_33341,N_33342,N_33343,N_33344,N_33345,N_33346,N_33347,N_33348,N_33349,N_33350,N_33351,N_33352,N_33353,N_33354,N_33355,N_33356,N_33357,N_33358,N_33359,N_33360,N_33361,N_33362,N_33363,N_33364,N_33365,N_33366,N_33367,N_33368,N_33369,N_33370,N_33371,N_33372,N_33373,N_33374,N_33375,N_33376,N_33377,N_33378,N_33379,N_33380,N_33381,N_33382,N_33383,N_33384,N_33385,N_33386,N_33387,N_33388,N_33389,N_33390,N_33391,N_33392,N_33393,N_33394,N_33395,N_33396,N_33397,N_33398,N_33399,N_33400,N_33401,N_33402,N_33403,N_33404,N_33405,N_33406,N_33407,N_33408,N_33409,N_33410,N_33411,N_33412,N_33413,N_33414,N_33415,N_33416,N_33417,N_33418,N_33419,N_33420,N_33421,N_33422,N_33423,N_33424,N_33425,N_33426,N_33427,N_33428,N_33429,N_33430,N_33431,N_33432,N_33433,N_33434,N_33435,N_33436,N_33437,N_33438,N_33439,N_33440,N_33441,N_33442,N_33443,N_33444,N_33445,N_33446,N_33447,N_33448,N_33449,N_33450,N_33451,N_33452,N_33453,N_33454,N_33455,N_33456,N_33457,N_33458,N_33459,N_33460,N_33461,N_33462,N_33463,N_33464,N_33465,N_33466,N_33467,N_33468,N_33469,N_33470,N_33471,N_33472,N_33473,N_33474,N_33475,N_33476,N_33477,N_33478,N_33479,N_33480,N_33481,N_33482,N_33483,N_33484,N_33485,N_33486,N_33487,N_33488,N_33489,N_33490,N_33491,N_33492,N_33493,N_33494,N_33495,N_33496,N_33497,N_33498,N_33499,N_33500,N_33501,N_33502,N_33503,N_33504,N_33505,N_33506,N_33507,N_33508,N_33509,N_33510,N_33511,N_33512,N_33513,N_33514,N_33515,N_33516,N_33517,N_33518,N_33519,N_33520,N_33521,N_33522,N_33523,N_33524,N_33525,N_33526,N_33527,N_33528,N_33529,N_33530,N_33531,N_33532,N_33533,N_33534,N_33535,N_33536,N_33537,N_33538,N_33539,N_33540,N_33541,N_33542,N_33543,N_33544,N_33545,N_33546,N_33547,N_33548,N_33549,N_33550,N_33551,N_33552,N_33553,N_33554,N_33555,N_33556,N_33557,N_33558,N_33559,N_33560,N_33561,N_33562,N_33563,N_33564,N_33565,N_33566,N_33567,N_33568,N_33569,N_33570,N_33571,N_33572,N_33573,N_33574,N_33575,N_33576,N_33577,N_33578,N_33579,N_33580,N_33581,N_33582,N_33583,N_33584,N_33585,N_33586,N_33587,N_33588,N_33589,N_33590,N_33591,N_33592,N_33593,N_33594,N_33595,N_33596,N_33597,N_33598,N_33599,N_33600,N_33601,N_33602,N_33603,N_33604,N_33605,N_33606,N_33607,N_33608,N_33609,N_33610,N_33611,N_33612,N_33613,N_33614,N_33615,N_33616,N_33617,N_33618,N_33619,N_33620,N_33621,N_33622,N_33623,N_33624,N_33625,N_33626,N_33627,N_33628,N_33629,N_33630,N_33631,N_33632,N_33633,N_33634,N_33635,N_33636,N_33637,N_33638,N_33639,N_33640,N_33641,N_33642,N_33643,N_33644,N_33645,N_33646,N_33647,N_33648,N_33649,N_33650,N_33651,N_33652,N_33653,N_33654,N_33655,N_33656,N_33657,N_33658,N_33659,N_33660,N_33661,N_33662,N_33663,N_33664,N_33665,N_33666,N_33667,N_33668,N_33669,N_33670,N_33671,N_33672,N_33673,N_33674,N_33675,N_33676,N_33677,N_33678,N_33679,N_33680,N_33681,N_33682,N_33683,N_33684,N_33685,N_33686,N_33687,N_33688,N_33689,N_33690,N_33691,N_33692,N_33693,N_33694,N_33695,N_33696,N_33697,N_33698,N_33699,N_33700,N_33701,N_33702,N_33703,N_33704,N_33705,N_33706,N_33707,N_33708,N_33709,N_33710,N_33711,N_33712,N_33713,N_33714,N_33715,N_33716,N_33717,N_33718,N_33719,N_33720,N_33721,N_33722,N_33723,N_33724,N_33725,N_33726,N_33727,N_33728,N_33729,N_33730,N_33731,N_33732,N_33733,N_33734,N_33735,N_33736,N_33737,N_33738,N_33739,N_33740,N_33741,N_33742,N_33743,N_33744,N_33745,N_33746,N_33747,N_33748,N_33749,N_33750,N_33751,N_33752,N_33753,N_33754,N_33755,N_33756,N_33757,N_33758,N_33759,N_33760,N_33761,N_33762,N_33763,N_33764,N_33765,N_33766,N_33767,N_33768,N_33769,N_33770,N_33771,N_33772,N_33773,N_33774,N_33775,N_33776,N_33777,N_33778,N_33779,N_33780,N_33781,N_33782,N_33783,N_33784,N_33785,N_33786,N_33787,N_33788,N_33789,N_33790,N_33791,N_33792,N_33793,N_33794,N_33795,N_33796,N_33797,N_33798,N_33799,N_33800,N_33801,N_33802,N_33803,N_33804,N_33805,N_33806,N_33807,N_33808,N_33809,N_33810,N_33811,N_33812,N_33813,N_33814,N_33815,N_33816,N_33817,N_33818,N_33819,N_33820,N_33821,N_33822,N_33823,N_33824,N_33825,N_33826,N_33827,N_33828,N_33829,N_33830,N_33831,N_33832,N_33833,N_33834,N_33835,N_33836,N_33837,N_33838,N_33839,N_33840,N_33841,N_33842,N_33843,N_33844,N_33845,N_33846,N_33847,N_33848,N_33849,N_33850,N_33851,N_33852,N_33853,N_33854,N_33855,N_33856,N_33857,N_33858,N_33859,N_33860,N_33861,N_33862,N_33863,N_33864,N_33865,N_33866,N_33867,N_33868,N_33869,N_33870,N_33871,N_33872,N_33873,N_33874,N_33875,N_33876,N_33877,N_33878,N_33879,N_33880,N_33881,N_33882,N_33883,N_33884,N_33885,N_33886,N_33887,N_33888,N_33889,N_33890,N_33891,N_33892,N_33893,N_33894,N_33895,N_33896,N_33897,N_33898,N_33899,N_33900,N_33901,N_33902,N_33903,N_33904,N_33905,N_33906,N_33907,N_33908,N_33909,N_33910,N_33911,N_33912,N_33913,N_33914,N_33915,N_33916,N_33917,N_33918,N_33919,N_33920,N_33921,N_33922,N_33923,N_33924,N_33925,N_33926,N_33927,N_33928,N_33929,N_33930,N_33931,N_33932,N_33933,N_33934,N_33935,N_33936,N_33937,N_33938,N_33939,N_33940,N_33941,N_33942,N_33943,N_33944,N_33945,N_33946,N_33947,N_33948,N_33949,N_33950,N_33951,N_33952,N_33953,N_33954,N_33955,N_33956,N_33957,N_33958,N_33959,N_33960,N_33961,N_33962,N_33963,N_33964,N_33965,N_33966,N_33967,N_33968,N_33969,N_33970,N_33971,N_33972,N_33973,N_33974,N_33975,N_33976,N_33977,N_33978,N_33979,N_33980,N_33981,N_33982,N_33983,N_33984,N_33985,N_33986,N_33987,N_33988,N_33989,N_33990,N_33991,N_33992,N_33993,N_33994,N_33995,N_33996,N_33997,N_33998,N_33999,N_34000,N_34001,N_34002,N_34003,N_34004,N_34005,N_34006,N_34007,N_34008,N_34009,N_34010,N_34011,N_34012,N_34013,N_34014,N_34015,N_34016,N_34017,N_34018,N_34019,N_34020,N_34021,N_34022,N_34023,N_34024,N_34025,N_34026,N_34027,N_34028,N_34029,N_34030,N_34031,N_34032,N_34033,N_34034,N_34035,N_34036,N_34037,N_34038,N_34039,N_34040,N_34041,N_34042,N_34043,N_34044,N_34045,N_34046,N_34047,N_34048,N_34049,N_34050,N_34051,N_34052,N_34053,N_34054,N_34055,N_34056,N_34057,N_34058,N_34059,N_34060,N_34061,N_34062,N_34063,N_34064,N_34065,N_34066,N_34067,N_34068,N_34069,N_34070,N_34071,N_34072,N_34073,N_34074,N_34075,N_34076,N_34077,N_34078,N_34079,N_34080,N_34081,N_34082,N_34083,N_34084,N_34085,N_34086,N_34087,N_34088,N_34089,N_34090,N_34091,N_34092,N_34093,N_34094,N_34095,N_34096,N_34097,N_34098,N_34099,N_34100,N_34101,N_34102,N_34103,N_34104,N_34105,N_34106,N_34107,N_34108,N_34109,N_34110,N_34111,N_34112,N_34113,N_34114,N_34115,N_34116,N_34117,N_34118,N_34119,N_34120,N_34121,N_34122,N_34123,N_34124,N_34125,N_34126,N_34127,N_34128,N_34129,N_34130,N_34131,N_34132,N_34133,N_34134,N_34135,N_34136,N_34137,N_34138,N_34139,N_34140,N_34141,N_34142,N_34143,N_34144,N_34145,N_34146,N_34147,N_34148,N_34149,N_34150,N_34151,N_34152,N_34153,N_34154,N_34155,N_34156,N_34157,N_34158,N_34159,N_34160,N_34161,N_34162,N_34163,N_34164,N_34165,N_34166,N_34167,N_34168,N_34169,N_34170,N_34171,N_34172,N_34173,N_34174,N_34175,N_34176,N_34177,N_34178,N_34179,N_34180,N_34181,N_34182,N_34183,N_34184,N_34185,N_34186,N_34187,N_34188,N_34189,N_34190,N_34191,N_34192,N_34193,N_34194,N_34195,N_34196,N_34197,N_34198,N_34199,N_34200,N_34201,N_34202,N_34203,N_34204,N_34205,N_34206,N_34207,N_34208,N_34209,N_34210,N_34211,N_34212,N_34213,N_34214,N_34215,N_34216,N_34217,N_34218,N_34219,N_34220,N_34221,N_34222,N_34223,N_34224,N_34225,N_34226,N_34227,N_34228,N_34229,N_34230,N_34231,N_34232,N_34233,N_34234,N_34235,N_34236,N_34237,N_34238,N_34239,N_34240,N_34241,N_34242,N_34243,N_34244,N_34245,N_34246,N_34247,N_34248,N_34249,N_34250,N_34251,N_34252,N_34253,N_34254,N_34255,N_34256,N_34257,N_34258,N_34259,N_34260,N_34261,N_34262,N_34263,N_34264,N_34265,N_34266,N_34267,N_34268,N_34269,N_34270,N_34271,N_34272,N_34273,N_34274,N_34275,N_34276,N_34277,N_34278,N_34279,N_34280,N_34281,N_34282,N_34283,N_34284,N_34285,N_34286,N_34287,N_34288,N_34289,N_34290,N_34291,N_34292,N_34293,N_34294,N_34295,N_34296,N_34297,N_34298,N_34299,N_34300,N_34301,N_34302,N_34303,N_34304,N_34305,N_34306,N_34307,N_34308,N_34309,N_34310,N_34311,N_34312,N_34313,N_34314,N_34315,N_34316,N_34317,N_34318,N_34319,N_34320,N_34321,N_34322,N_34323,N_34324,N_34325,N_34326,N_34327,N_34328,N_34329,N_34330,N_34331,N_34332,N_34333,N_34334,N_34335,N_34336,N_34337,N_34338,N_34339,N_34340,N_34341,N_34342,N_34343,N_34344,N_34345,N_34346,N_34347,N_34348,N_34349,N_34350,N_34351,N_34352,N_34353,N_34354,N_34355,N_34356,N_34357,N_34358,N_34359,N_34360,N_34361,N_34362,N_34363,N_34364,N_34365,N_34366,N_34367,N_34368,N_34369,N_34370,N_34371,N_34372,N_34373,N_34374,N_34375,N_34376,N_34377,N_34378,N_34379,N_34380,N_34381,N_34382,N_34383,N_34384,N_34385,N_34386,N_34387,N_34388,N_34389,N_34390,N_34391,N_34392,N_34393,N_34394,N_34395,N_34396,N_34397,N_34398,N_34399,N_34400,N_34401,N_34402,N_34403,N_34404,N_34405,N_34406,N_34407,N_34408,N_34409,N_34410,N_34411,N_34412,N_34413,N_34414,N_34415,N_34416,N_34417,N_34418,N_34419,N_34420,N_34421,N_34422,N_34423,N_34424,N_34425,N_34426,N_34427,N_34428,N_34429,N_34430,N_34431,N_34432,N_34433,N_34434,N_34435,N_34436,N_34437,N_34438,N_34439,N_34440,N_34441,N_34442,N_34443,N_34444,N_34445,N_34446,N_34447,N_34448,N_34449,N_34450,N_34451,N_34452,N_34453,N_34454,N_34455,N_34456,N_34457,N_34458,N_34459,N_34460,N_34461,N_34462,N_34463,N_34464,N_34465,N_34466,N_34467,N_34468,N_34469,N_34470,N_34471,N_34472,N_34473,N_34474,N_34475,N_34476,N_34477,N_34478,N_34479,N_34480,N_34481,N_34482,N_34483,N_34484,N_34485,N_34486,N_34487,N_34488,N_34489,N_34490,N_34491,N_34492,N_34493,N_34494,N_34495,N_34496,N_34497,N_34498,N_34499,N_34500,N_34501,N_34502,N_34503,N_34504,N_34505,N_34506,N_34507,N_34508,N_34509,N_34510,N_34511,N_34512,N_34513,N_34514,N_34515,N_34516,N_34517,N_34518,N_34519,N_34520,N_34521,N_34522,N_34523,N_34524,N_34525,N_34526,N_34527,N_34528,N_34529,N_34530,N_34531,N_34532,N_34533,N_34534,N_34535,N_34536,N_34537,N_34538,N_34539,N_34540,N_34541,N_34542,N_34543,N_34544,N_34545,N_34546,N_34547,N_34548,N_34549,N_34550,N_34551,N_34552,N_34553,N_34554,N_34555,N_34556,N_34557,N_34558,N_34559,N_34560,N_34561,N_34562,N_34563,N_34564,N_34565,N_34566,N_34567,N_34568,N_34569,N_34570,N_34571,N_34572,N_34573,N_34574,N_34575,N_34576,N_34577,N_34578,N_34579,N_34580,N_34581,N_34582,N_34583,N_34584,N_34585,N_34586,N_34587,N_34588,N_34589,N_34590,N_34591,N_34592,N_34593,N_34594,N_34595,N_34596,N_34597,N_34598,N_34599,N_34600,N_34601,N_34602,N_34603,N_34604,N_34605,N_34606,N_34607,N_34608,N_34609,N_34610,N_34611,N_34612,N_34613,N_34614,N_34615,N_34616,N_34617,N_34618,N_34619,N_34620,N_34621,N_34622,N_34623,N_34624,N_34625,N_34626,N_34627,N_34628,N_34629,N_34630,N_34631,N_34632,N_34633,N_34634,N_34635,N_34636,N_34637,N_34638,N_34639,N_34640,N_34641,N_34642,N_34643,N_34644,N_34645,N_34646,N_34647,N_34648,N_34649,N_34650,N_34651,N_34652,N_34653,N_34654,N_34655,N_34656,N_34657,N_34658,N_34659,N_34660,N_34661,N_34662,N_34663,N_34664,N_34665,N_34666,N_34667,N_34668,N_34669,N_34670,N_34671,N_34672,N_34673,N_34674,N_34675,N_34676,N_34677,N_34678,N_34679,N_34680,N_34681,N_34682,N_34683,N_34684,N_34685,N_34686,N_34687,N_34688,N_34689,N_34690,N_34691,N_34692,N_34693,N_34694,N_34695,N_34696,N_34697,N_34698,N_34699,N_34700,N_34701,N_34702,N_34703,N_34704,N_34705,N_34706,N_34707,N_34708,N_34709,N_34710,N_34711,N_34712,N_34713,N_34714,N_34715,N_34716,N_34717,N_34718,N_34719,N_34720,N_34721,N_34722,N_34723,N_34724,N_34725,N_34726,N_34727,N_34728,N_34729,N_34730,N_34731,N_34732,N_34733,N_34734,N_34735,N_34736,N_34737,N_34738,N_34739,N_34740,N_34741,N_34742,N_34743,N_34744,N_34745,N_34746,N_34747,N_34748,N_34749,N_34750,N_34751,N_34752,N_34753,N_34754,N_34755,N_34756,N_34757,N_34758,N_34759,N_34760,N_34761,N_34762,N_34763,N_34764,N_34765,N_34766,N_34767,N_34768,N_34769,N_34770,N_34771,N_34772,N_34773,N_34774,N_34775,N_34776,N_34777,N_34778,N_34779,N_34780,N_34781,N_34782,N_34783,N_34784,N_34785,N_34786,N_34787,N_34788,N_34789,N_34790,N_34791,N_34792,N_34793,N_34794,N_34795,N_34796,N_34797,N_34798,N_34799,N_34800,N_34801,N_34802,N_34803,N_34804,N_34805,N_34806,N_34807,N_34808,N_34809,N_34810,N_34811,N_34812,N_34813,N_34814,N_34815,N_34816,N_34817,N_34818,N_34819,N_34820,N_34821,N_34822,N_34823,N_34824,N_34825,N_34826,N_34827,N_34828,N_34829,N_34830,N_34831,N_34832,N_34833,N_34834,N_34835,N_34836,N_34837,N_34838,N_34839,N_34840,N_34841,N_34842,N_34843,N_34844,N_34845,N_34846,N_34847,N_34848,N_34849,N_34850,N_34851,N_34852,N_34853,N_34854,N_34855,N_34856,N_34857,N_34858,N_34859,N_34860,N_34861,N_34862,N_34863,N_34864,N_34865,N_34866,N_34867,N_34868,N_34869,N_34870,N_34871,N_34872,N_34873,N_34874,N_34875,N_34876,N_34877,N_34878,N_34879,N_34880,N_34881,N_34882,N_34883,N_34884,N_34885,N_34886,N_34887,N_34888,N_34889,N_34890,N_34891,N_34892,N_34893,N_34894,N_34895,N_34896,N_34897,N_34898,N_34899,N_34900,N_34901,N_34902,N_34903,N_34904,N_34905,N_34906,N_34907,N_34908,N_34909,N_34910,N_34911,N_34912,N_34913,N_34914,N_34915,N_34916,N_34917,N_34918,N_34919,N_34920,N_34921,N_34922,N_34923,N_34924,N_34925,N_34926,N_34927,N_34928,N_34929,N_34930,N_34931,N_34932,N_34933,N_34934,N_34935,N_34936,N_34937,N_34938,N_34939,N_34940,N_34941,N_34942,N_34943,N_34944,N_34945,N_34946,N_34947,N_34948,N_34949,N_34950,N_34951,N_34952,N_34953,N_34954,N_34955,N_34956,N_34957,N_34958,N_34959,N_34960,N_34961,N_34962,N_34963,N_34964,N_34965,N_34966,N_34967,N_34968,N_34969,N_34970,N_34971,N_34972,N_34973,N_34974,N_34975,N_34976,N_34977,N_34978,N_34979,N_34980,N_34981,N_34982,N_34983,N_34984,N_34985,N_34986,N_34987,N_34988,N_34989,N_34990,N_34991,N_34992,N_34993,N_34994,N_34995,N_34996,N_34997,N_34998,N_34999,N_35000,N_35001,N_35002,N_35003,N_35004,N_35005,N_35006,N_35007,N_35008,N_35009,N_35010,N_35011,N_35012,N_35013,N_35014,N_35015,N_35016,N_35017,N_35018,N_35019,N_35020,N_35021,N_35022,N_35023,N_35024,N_35025,N_35026,N_35027,N_35028,N_35029,N_35030,N_35031,N_35032,N_35033,N_35034,N_35035,N_35036,N_35037,N_35038,N_35039,N_35040,N_35041,N_35042,N_35043,N_35044,N_35045,N_35046,N_35047,N_35048,N_35049,N_35050,N_35051,N_35052,N_35053,N_35054,N_35055,N_35056,N_35057,N_35058,N_35059,N_35060,N_35061,N_35062,N_35063,N_35064,N_35065,N_35066,N_35067,N_35068,N_35069,N_35070,N_35071,N_35072,N_35073,N_35074,N_35075,N_35076,N_35077,N_35078,N_35079,N_35080,N_35081,N_35082,N_35083,N_35084,N_35085,N_35086,N_35087,N_35088,N_35089,N_35090,N_35091,N_35092,N_35093,N_35094,N_35095,N_35096,N_35097,N_35098,N_35099,N_35100,N_35101,N_35102,N_35103,N_35104,N_35105,N_35106,N_35107,N_35108,N_35109,N_35110,N_35111,N_35112,N_35113,N_35114,N_35115,N_35116,N_35117,N_35118,N_35119,N_35120,N_35121,N_35122,N_35123,N_35124,N_35125,N_35126,N_35127,N_35128,N_35129,N_35130,N_35131,N_35132,N_35133,N_35134,N_35135,N_35136,N_35137,N_35138,N_35139,N_35140,N_35141,N_35142,N_35143,N_35144,N_35145,N_35146,N_35147,N_35148,N_35149,N_35150,N_35151,N_35152,N_35153,N_35154,N_35155,N_35156,N_35157,N_35158,N_35159,N_35160,N_35161,N_35162,N_35163,N_35164,N_35165,N_35166,N_35167,N_35168,N_35169,N_35170,N_35171,N_35172,N_35173,N_35174,N_35175,N_35176,N_35177,N_35178,N_35179,N_35180,N_35181,N_35182,N_35183,N_35184,N_35185,N_35186,N_35187,N_35188,N_35189,N_35190,N_35191,N_35192,N_35193,N_35194,N_35195,N_35196,N_35197,N_35198,N_35199,N_35200,N_35201,N_35202,N_35203,N_35204,N_35205,N_35206,N_35207,N_35208,N_35209,N_35210,N_35211,N_35212,N_35213,N_35214,N_35215,N_35216,N_35217,N_35218,N_35219,N_35220,N_35221,N_35222,N_35223,N_35224,N_35225,N_35226,N_35227,N_35228,N_35229,N_35230,N_35231,N_35232,N_35233,N_35234,N_35235,N_35236,N_35237,N_35238,N_35239,N_35240,N_35241,N_35242,N_35243,N_35244,N_35245,N_35246,N_35247,N_35248,N_35249,N_35250,N_35251,N_35252,N_35253,N_35254,N_35255,N_35256,N_35257,N_35258,N_35259,N_35260,N_35261,N_35262,N_35263,N_35264,N_35265,N_35266,N_35267,N_35268,N_35269,N_35270,N_35271,N_35272,N_35273,N_35274,N_35275,N_35276,N_35277,N_35278,N_35279,N_35280,N_35281,N_35282,N_35283,N_35284,N_35285,N_35286,N_35287,N_35288,N_35289,N_35290,N_35291,N_35292,N_35293,N_35294,N_35295,N_35296,N_35297,N_35298,N_35299,N_35300,N_35301,N_35302,N_35303,N_35304,N_35305,N_35306,N_35307,N_35308,N_35309,N_35310,N_35311,N_35312,N_35313,N_35314,N_35315,N_35316,N_35317,N_35318,N_35319,N_35320,N_35321,N_35322,N_35323,N_35324,N_35325,N_35326,N_35327,N_35328,N_35329,N_35330,N_35331,N_35332,N_35333,N_35334,N_35335,N_35336,N_35337,N_35338,N_35339,N_35340,N_35341,N_35342,N_35343,N_35344,N_35345,N_35346,N_35347,N_35348,N_35349,N_35350,N_35351,N_35352,N_35353,N_35354,N_35355,N_35356,N_35357,N_35358,N_35359,N_35360,N_35361,N_35362,N_35363,N_35364,N_35365,N_35366,N_35367,N_35368,N_35369,N_35370,N_35371,N_35372,N_35373,N_35374,N_35375,N_35376,N_35377,N_35378,N_35379,N_35380,N_35381,N_35382,N_35383,N_35384,N_35385,N_35386,N_35387,N_35388,N_35389,N_35390,N_35391,N_35392,N_35393,N_35394,N_35395,N_35396,N_35397,N_35398,N_35399,N_35400,N_35401,N_35402,N_35403,N_35404,N_35405,N_35406,N_35407,N_35408,N_35409,N_35410,N_35411,N_35412,N_35413,N_35414,N_35415,N_35416,N_35417,N_35418,N_35419,N_35420,N_35421,N_35422,N_35423,N_35424,N_35425,N_35426,N_35427,N_35428,N_35429,N_35430,N_35431,N_35432,N_35433,N_35434,N_35435,N_35436,N_35437,N_35438,N_35439,N_35440,N_35441,N_35442,N_35443,N_35444,N_35445,N_35446,N_35447,N_35448,N_35449,N_35450,N_35451,N_35452,N_35453,N_35454,N_35455,N_35456,N_35457,N_35458,N_35459,N_35460,N_35461,N_35462,N_35463,N_35464,N_35465,N_35466,N_35467,N_35468,N_35469,N_35470,N_35471,N_35472,N_35473,N_35474,N_35475,N_35476,N_35477,N_35478,N_35479,N_35480,N_35481,N_35482,N_35483,N_35484,N_35485,N_35486,N_35487,N_35488,N_35489,N_35490,N_35491,N_35492,N_35493,N_35494,N_35495,N_35496,N_35497,N_35498,N_35499,N_35500,N_35501,N_35502,N_35503,N_35504,N_35505,N_35506,N_35507,N_35508,N_35509,N_35510,N_35511,N_35512,N_35513,N_35514,N_35515,N_35516,N_35517,N_35518,N_35519,N_35520,N_35521,N_35522,N_35523,N_35524,N_35525,N_35526,N_35527,N_35528,N_35529,N_35530,N_35531,N_35532,N_35533,N_35534,N_35535,N_35536,N_35537,N_35538,N_35539,N_35540,N_35541,N_35542,N_35543,N_35544,N_35545,N_35546,N_35547,N_35548,N_35549,N_35550,N_35551,N_35552,N_35553,N_35554,N_35555,N_35556,N_35557,N_35558,N_35559,N_35560,N_35561,N_35562,N_35563,N_35564,N_35565,N_35566,N_35567,N_35568,N_35569,N_35570,N_35571,N_35572,N_35573,N_35574,N_35575,N_35576,N_35577,N_35578,N_35579,N_35580,N_35581,N_35582,N_35583,N_35584,N_35585,N_35586,N_35587,N_35588,N_35589,N_35590,N_35591,N_35592,N_35593,N_35594,N_35595,N_35596,N_35597,N_35598,N_35599,N_35600,N_35601,N_35602,N_35603,N_35604,N_35605,N_35606,N_35607,N_35608,N_35609,N_35610,N_35611,N_35612,N_35613,N_35614,N_35615,N_35616,N_35617,N_35618,N_35619,N_35620,N_35621,N_35622,N_35623,N_35624,N_35625,N_35626,N_35627,N_35628,N_35629,N_35630,N_35631,N_35632,N_35633,N_35634,N_35635,N_35636,N_35637,N_35638,N_35639,N_35640,N_35641,N_35642,N_35643,N_35644,N_35645,N_35646,N_35647,N_35648,N_35649,N_35650,N_35651,N_35652,N_35653,N_35654,N_35655,N_35656,N_35657,N_35658,N_35659,N_35660,N_35661,N_35662,N_35663,N_35664,N_35665,N_35666,N_35667,N_35668,N_35669,N_35670,N_35671,N_35672,N_35673,N_35674,N_35675,N_35676,N_35677,N_35678,N_35679,N_35680,N_35681,N_35682,N_35683,N_35684,N_35685,N_35686,N_35687,N_35688,N_35689,N_35690,N_35691,N_35692,N_35693,N_35694,N_35695,N_35696,N_35697,N_35698,N_35699,N_35700,N_35701,N_35702,N_35703,N_35704,N_35705,N_35706,N_35707,N_35708,N_35709,N_35710,N_35711,N_35712,N_35713,N_35714,N_35715,N_35716,N_35717,N_35718,N_35719,N_35720,N_35721,N_35722,N_35723,N_35724,N_35725,N_35726,N_35727,N_35728,N_35729,N_35730,N_35731,N_35732,N_35733,N_35734,N_35735,N_35736,N_35737,N_35738,N_35739,N_35740,N_35741,N_35742,N_35743,N_35744,N_35745,N_35746,N_35747,N_35748,N_35749,N_35750,N_35751,N_35752,N_35753,N_35754,N_35755,N_35756,N_35757,N_35758,N_35759,N_35760,N_35761,N_35762,N_35763,N_35764,N_35765,N_35766,N_35767,N_35768,N_35769,N_35770,N_35771,N_35772,N_35773,N_35774,N_35775,N_35776,N_35777,N_35778,N_35779,N_35780,N_35781,N_35782,N_35783,N_35784,N_35785,N_35786,N_35787,N_35788,N_35789,N_35790,N_35791,N_35792,N_35793,N_35794,N_35795,N_35796,N_35797,N_35798,N_35799,N_35800,N_35801,N_35802,N_35803,N_35804,N_35805,N_35806,N_35807,N_35808,N_35809,N_35810,N_35811,N_35812,N_35813,N_35814,N_35815,N_35816,N_35817,N_35818,N_35819,N_35820,N_35821,N_35822,N_35823,N_35824,N_35825,N_35826,N_35827,N_35828,N_35829,N_35830,N_35831,N_35832,N_35833,N_35834,N_35835,N_35836,N_35837,N_35838,N_35839,N_35840,N_35841,N_35842,N_35843,N_35844,N_35845,N_35846,N_35847,N_35848,N_35849,N_35850,N_35851,N_35852,N_35853,N_35854,N_35855,N_35856,N_35857,N_35858,N_35859,N_35860,N_35861,N_35862,N_35863,N_35864,N_35865,N_35866,N_35867,N_35868,N_35869,N_35870,N_35871,N_35872,N_35873,N_35874,N_35875,N_35876,N_35877,N_35878,N_35879,N_35880,N_35881,N_35882,N_35883,N_35884,N_35885,N_35886,N_35887,N_35888,N_35889,N_35890,N_35891,N_35892,N_35893,N_35894,N_35895,N_35896,N_35897,N_35898,N_35899,N_35900,N_35901,N_35902,N_35903,N_35904,N_35905,N_35906,N_35907,N_35908,N_35909,N_35910,N_35911,N_35912,N_35913,N_35914,N_35915,N_35916,N_35917,N_35918,N_35919,N_35920,N_35921,N_35922,N_35923,N_35924,N_35925,N_35926,N_35927,N_35928,N_35929,N_35930,N_35931,N_35932,N_35933,N_35934,N_35935,N_35936,N_35937,N_35938,N_35939,N_35940,N_35941,N_35942,N_35943,N_35944,N_35945,N_35946,N_35947,N_35948,N_35949,N_35950,N_35951,N_35952,N_35953,N_35954,N_35955,N_35956,N_35957,N_35958,N_35959,N_35960,N_35961,N_35962,N_35963,N_35964,N_35965,N_35966,N_35967,N_35968,N_35969,N_35970,N_35971,N_35972,N_35973,N_35974,N_35975,N_35976,N_35977,N_35978,N_35979,N_35980,N_35981,N_35982,N_35983,N_35984,N_35985,N_35986,N_35987,N_35988,N_35989,N_35990,N_35991,N_35992,N_35993,N_35994,N_35995,N_35996,N_35997,N_35998,N_35999,N_36000,N_36001,N_36002,N_36003,N_36004,N_36005,N_36006,N_36007,N_36008,N_36009,N_36010,N_36011,N_36012,N_36013,N_36014,N_36015,N_36016,N_36017,N_36018,N_36019,N_36020,N_36021,N_36022,N_36023,N_36024,N_36025,N_36026,N_36027,N_36028,N_36029,N_36030,N_36031,N_36032,N_36033,N_36034,N_36035,N_36036,N_36037,N_36038,N_36039,N_36040,N_36041,N_36042,N_36043,N_36044,N_36045,N_36046,N_36047,N_36048,N_36049,N_36050,N_36051,N_36052,N_36053,N_36054,N_36055,N_36056,N_36057,N_36058,N_36059,N_36060,N_36061,N_36062,N_36063,N_36064,N_36065,N_36066,N_36067,N_36068,N_36069,N_36070,N_36071,N_36072,N_36073,N_36074,N_36075,N_36076,N_36077,N_36078,N_36079,N_36080,N_36081,N_36082,N_36083,N_36084,N_36085,N_36086,N_36087,N_36088,N_36089,N_36090,N_36091,N_36092,N_36093,N_36094,N_36095,N_36096,N_36097,N_36098,N_36099,N_36100,N_36101,N_36102,N_36103,N_36104,N_36105,N_36106,N_36107,N_36108,N_36109,N_36110,N_36111,N_36112,N_36113,N_36114,N_36115,N_36116,N_36117,N_36118,N_36119,N_36120,N_36121,N_36122,N_36123,N_36124,N_36125,N_36126,N_36127,N_36128,N_36129,N_36130,N_36131,N_36132,N_36133,N_36134,N_36135,N_36136,N_36137,N_36138,N_36139,N_36140,N_36141,N_36142,N_36143,N_36144,N_36145,N_36146,N_36147,N_36148,N_36149,N_36150,N_36151,N_36152,N_36153,N_36154,N_36155,N_36156,N_36157,N_36158,N_36159,N_36160,N_36161,N_36162,N_36163,N_36164,N_36165,N_36166,N_36167,N_36168,N_36169,N_36170,N_36171,N_36172,N_36173,N_36174,N_36175,N_36176,N_36177,N_36178,N_36179,N_36180,N_36181,N_36182,N_36183,N_36184,N_36185,N_36186,N_36187,N_36188,N_36189,N_36190,N_36191,N_36192,N_36193,N_36194,N_36195,N_36196,N_36197,N_36198,N_36199,N_36200,N_36201,N_36202,N_36203,N_36204,N_36205,N_36206,N_36207,N_36208,N_36209,N_36210,N_36211,N_36212,N_36213,N_36214,N_36215,N_36216,N_36217,N_36218,N_36219,N_36220,N_36221,N_36222,N_36223,N_36224,N_36225,N_36226,N_36227,N_36228,N_36229,N_36230,N_36231,N_36232,N_36233,N_36234,N_36235,N_36236,N_36237,N_36238,N_36239,N_36240,N_36241,N_36242,N_36243,N_36244,N_36245,N_36246,N_36247,N_36248,N_36249,N_36250,N_36251,N_36252,N_36253,N_36254,N_36255,N_36256,N_36257,N_36258,N_36259,N_36260,N_36261,N_36262,N_36263,N_36264,N_36265,N_36266,N_36267,N_36268,N_36269,N_36270,N_36271,N_36272,N_36273,N_36274,N_36275,N_36276,N_36277,N_36278,N_36279,N_36280,N_36281,N_36282,N_36283,N_36284,N_36285,N_36286,N_36287,N_36288,N_36289,N_36290,N_36291,N_36292,N_36293,N_36294,N_36295,N_36296,N_36297,N_36298,N_36299,N_36300,N_36301,N_36302,N_36303,N_36304,N_36305,N_36306,N_36307,N_36308,N_36309,N_36310,N_36311,N_36312,N_36313,N_36314,N_36315,N_36316,N_36317,N_36318,N_36319,N_36320,N_36321,N_36322,N_36323,N_36324,N_36325,N_36326,N_36327,N_36328,N_36329,N_36330,N_36331,N_36332,N_36333,N_36334,N_36335,N_36336,N_36337,N_36338,N_36339,N_36340,N_36341,N_36342,N_36343,N_36344,N_36345,N_36346,N_36347,N_36348,N_36349,N_36350,N_36351,N_36352,N_36353,N_36354,N_36355,N_36356,N_36357,N_36358,N_36359,N_36360,N_36361,N_36362,N_36363,N_36364,N_36365,N_36366,N_36367,N_36368,N_36369,N_36370,N_36371,N_36372,N_36373,N_36374,N_36375,N_36376,N_36377,N_36378,N_36379,N_36380,N_36381,N_36382,N_36383,N_36384,N_36385,N_36386,N_36387,N_36388,N_36389,N_36390,N_36391,N_36392,N_36393,N_36394,N_36395,N_36396,N_36397,N_36398,N_36399,N_36400,N_36401,N_36402,N_36403,N_36404,N_36405,N_36406,N_36407,N_36408,N_36409,N_36410,N_36411,N_36412,N_36413,N_36414,N_36415,N_36416,N_36417,N_36418,N_36419,N_36420,N_36421,N_36422,N_36423,N_36424,N_36425,N_36426,N_36427,N_36428,N_36429,N_36430,N_36431,N_36432,N_36433,N_36434,N_36435,N_36436,N_36437,N_36438,N_36439,N_36440,N_36441,N_36442,N_36443,N_36444,N_36445,N_36446,N_36447,N_36448,N_36449,N_36450,N_36451,N_36452,N_36453,N_36454,N_36455,N_36456,N_36457,N_36458,N_36459,N_36460,N_36461,N_36462,N_36463,N_36464,N_36465,N_36466,N_36467,N_36468,N_36469,N_36470,N_36471,N_36472,N_36473,N_36474,N_36475,N_36476,N_36477,N_36478,N_36479,N_36480,N_36481,N_36482,N_36483,N_36484,N_36485,N_36486,N_36487,N_36488,N_36489,N_36490,N_36491,N_36492,N_36493,N_36494,N_36495,N_36496,N_36497,N_36498,N_36499,N_36500,N_36501,N_36502,N_36503,N_36504,N_36505,N_36506,N_36507,N_36508,N_36509,N_36510,N_36511,N_36512,N_36513,N_36514,N_36515,N_36516,N_36517,N_36518,N_36519,N_36520,N_36521,N_36522,N_36523,N_36524,N_36525,N_36526,N_36527,N_36528,N_36529,N_36530,N_36531,N_36532,N_36533,N_36534,N_36535,N_36536,N_36537,N_36538,N_36539,N_36540,N_36541,N_36542,N_36543,N_36544,N_36545,N_36546,N_36547,N_36548,N_36549,N_36550,N_36551,N_36552,N_36553,N_36554,N_36555,N_36556,N_36557,N_36558,N_36559,N_36560,N_36561,N_36562,N_36563,N_36564,N_36565,N_36566,N_36567,N_36568,N_36569,N_36570,N_36571,N_36572,N_36573,N_36574,N_36575,N_36576,N_36577,N_36578,N_36579,N_36580,N_36581,N_36582,N_36583,N_36584,N_36585,N_36586,N_36587,N_36588,N_36589,N_36590,N_36591,N_36592,N_36593,N_36594,N_36595,N_36596,N_36597,N_36598,N_36599,N_36600,N_36601,N_36602,N_36603,N_36604,N_36605,N_36606,N_36607,N_36608,N_36609,N_36610,N_36611,N_36612,N_36613,N_36614,N_36615,N_36616,N_36617,N_36618,N_36619,N_36620,N_36621,N_36622,N_36623,N_36624,N_36625,N_36626,N_36627,N_36628,N_36629,N_36630,N_36631,N_36632,N_36633,N_36634,N_36635,N_36636,N_36637,N_36638,N_36639,N_36640,N_36641,N_36642,N_36643,N_36644,N_36645,N_36646,N_36647,N_36648,N_36649,N_36650,N_36651,N_36652,N_36653,N_36654,N_36655,N_36656,N_36657,N_36658,N_36659,N_36660,N_36661,N_36662,N_36663,N_36664,N_36665,N_36666,N_36667,N_36668,N_36669,N_36670,N_36671,N_36672,N_36673,N_36674,N_36675,N_36676,N_36677,N_36678,N_36679,N_36680,N_36681,N_36682,N_36683,N_36684,N_36685,N_36686,N_36687,N_36688,N_36689,N_36690,N_36691,N_36692,N_36693,N_36694,N_36695,N_36696,N_36697,N_36698,N_36699,N_36700,N_36701,N_36702,N_36703,N_36704,N_36705,N_36706,N_36707,N_36708,N_36709,N_36710,N_36711,N_36712,N_36713,N_36714,N_36715,N_36716,N_36717,N_36718,N_36719,N_36720,N_36721,N_36722,N_36723,N_36724,N_36725,N_36726,N_36727,N_36728,N_36729,N_36730,N_36731,N_36732,N_36733,N_36734,N_36735,N_36736,N_36737,N_36738,N_36739,N_36740,N_36741,N_36742,N_36743,N_36744,N_36745,N_36746,N_36747,N_36748,N_36749,N_36750,N_36751,N_36752,N_36753,N_36754,N_36755,N_36756,N_36757,N_36758,N_36759,N_36760,N_36761,N_36762,N_36763,N_36764,N_36765,N_36766,N_36767,N_36768,N_36769,N_36770,N_36771,N_36772,N_36773,N_36774,N_36775,N_36776,N_36777,N_36778,N_36779,N_36780,N_36781,N_36782,N_36783,N_36784,N_36785,N_36786,N_36787,N_36788,N_36789,N_36790,N_36791,N_36792,N_36793,N_36794,N_36795,N_36796,N_36797,N_36798,N_36799,N_36800,N_36801,N_36802,N_36803,N_36804,N_36805,N_36806,N_36807,N_36808,N_36809,N_36810,N_36811,N_36812,N_36813,N_36814,N_36815,N_36816,N_36817,N_36818,N_36819,N_36820,N_36821,N_36822,N_36823,N_36824,N_36825,N_36826,N_36827,N_36828,N_36829,N_36830,N_36831,N_36832,N_36833,N_36834,N_36835,N_36836,N_36837,N_36838,N_36839,N_36840,N_36841,N_36842,N_36843,N_36844,N_36845,N_36846,N_36847,N_36848,N_36849,N_36850,N_36851,N_36852,N_36853,N_36854,N_36855,N_36856,N_36857,N_36858,N_36859,N_36860,N_36861,N_36862,N_36863,N_36864,N_36865,N_36866,N_36867,N_36868,N_36869,N_36870,N_36871,N_36872,N_36873,N_36874,N_36875,N_36876,N_36877,N_36878,N_36879,N_36880,N_36881,N_36882,N_36883,N_36884,N_36885,N_36886,N_36887,N_36888,N_36889,N_36890,N_36891,N_36892,N_36893,N_36894,N_36895,N_36896,N_36897,N_36898,N_36899,N_36900,N_36901,N_36902,N_36903,N_36904,N_36905,N_36906,N_36907,N_36908,N_36909,N_36910,N_36911,N_36912,N_36913,N_36914,N_36915,N_36916,N_36917,N_36918,N_36919,N_36920,N_36921,N_36922,N_36923,N_36924,N_36925,N_36926,N_36927,N_36928,N_36929,N_36930,N_36931,N_36932,N_36933,N_36934,N_36935,N_36936,N_36937,N_36938,N_36939,N_36940,N_36941,N_36942,N_36943,N_36944,N_36945,N_36946,N_36947,N_36948,N_36949,N_36950,N_36951,N_36952,N_36953,N_36954,N_36955,N_36956,N_36957,N_36958,N_36959,N_36960,N_36961,N_36962,N_36963,N_36964,N_36965,N_36966,N_36967,N_36968,N_36969,N_36970,N_36971,N_36972,N_36973,N_36974,N_36975,N_36976,N_36977,N_36978,N_36979,N_36980,N_36981,N_36982,N_36983,N_36984,N_36985,N_36986,N_36987,N_36988,N_36989,N_36990,N_36991,N_36992,N_36993,N_36994,N_36995,N_36996,N_36997,N_36998,N_36999,N_37000,N_37001,N_37002,N_37003,N_37004,N_37005,N_37006,N_37007,N_37008,N_37009,N_37010,N_37011,N_37012,N_37013,N_37014,N_37015,N_37016,N_37017,N_37018,N_37019,N_37020,N_37021,N_37022,N_37023,N_37024,N_37025,N_37026,N_37027,N_37028,N_37029,N_37030,N_37031,N_37032,N_37033,N_37034,N_37035,N_37036,N_37037,N_37038,N_37039,N_37040,N_37041,N_37042,N_37043,N_37044,N_37045,N_37046,N_37047,N_37048,N_37049,N_37050,N_37051,N_37052,N_37053,N_37054,N_37055,N_37056,N_37057,N_37058,N_37059,N_37060,N_37061,N_37062,N_37063,N_37064,N_37065,N_37066,N_37067,N_37068,N_37069,N_37070,N_37071,N_37072,N_37073,N_37074,N_37075,N_37076,N_37077,N_37078,N_37079,N_37080,N_37081,N_37082,N_37083,N_37084,N_37085,N_37086,N_37087,N_37088,N_37089,N_37090,N_37091,N_37092,N_37093,N_37094,N_37095,N_37096,N_37097,N_37098,N_37099,N_37100,N_37101,N_37102,N_37103,N_37104,N_37105,N_37106,N_37107,N_37108,N_37109,N_37110,N_37111,N_37112,N_37113,N_37114,N_37115,N_37116,N_37117,N_37118,N_37119,N_37120,N_37121,N_37122,N_37123,N_37124,N_37125,N_37126,N_37127,N_37128,N_37129,N_37130,N_37131,N_37132,N_37133,N_37134,N_37135,N_37136,N_37137,N_37138,N_37139,N_37140,N_37141,N_37142,N_37143,N_37144,N_37145,N_37146,N_37147,N_37148,N_37149,N_37150,N_37151,N_37152,N_37153,N_37154,N_37155,N_37156,N_37157,N_37158,N_37159,N_37160,N_37161,N_37162,N_37163,N_37164,N_37165,N_37166,N_37167,N_37168,N_37169,N_37170,N_37171,N_37172,N_37173,N_37174,N_37175,N_37176,N_37177,N_37178,N_37179,N_37180,N_37181,N_37182,N_37183,N_37184,N_37185,N_37186,N_37187,N_37188,N_37189,N_37190,N_37191,N_37192,N_37193,N_37194,N_37195,N_37196,N_37197,N_37198,N_37199,N_37200,N_37201,N_37202,N_37203,N_37204,N_37205,N_37206,N_37207,N_37208,N_37209,N_37210,N_37211,N_37212,N_37213,N_37214,N_37215,N_37216,N_37217,N_37218,N_37219,N_37220,N_37221,N_37222,N_37223,N_37224,N_37225,N_37226,N_37227,N_37228,N_37229,N_37230,N_37231,N_37232,N_37233,N_37234,N_37235,N_37236,N_37237,N_37238,N_37239,N_37240,N_37241,N_37242,N_37243,N_37244,N_37245,N_37246,N_37247,N_37248,N_37249,N_37250,N_37251,N_37252,N_37253,N_37254,N_37255,N_37256,N_37257,N_37258,N_37259,N_37260,N_37261,N_37262,N_37263,N_37264,N_37265,N_37266,N_37267,N_37268,N_37269,N_37270,N_37271,N_37272,N_37273,N_37274,N_37275,N_37276,N_37277,N_37278,N_37279,N_37280,N_37281,N_37282,N_37283,N_37284,N_37285,N_37286,N_37287,N_37288,N_37289,N_37290,N_37291,N_37292,N_37293,N_37294,N_37295,N_37296,N_37297,N_37298,N_37299,N_37300,N_37301,N_37302,N_37303,N_37304,N_37305,N_37306,N_37307,N_37308,N_37309,N_37310,N_37311,N_37312,N_37313,N_37314,N_37315,N_37316,N_37317,N_37318,N_37319,N_37320,N_37321,N_37322,N_37323,N_37324,N_37325,N_37326,N_37327,N_37328,N_37329,N_37330,N_37331,N_37332,N_37333,N_37334,N_37335,N_37336,N_37337,N_37338,N_37339,N_37340,N_37341,N_37342,N_37343,N_37344,N_37345,N_37346,N_37347,N_37348,N_37349,N_37350,N_37351,N_37352,N_37353,N_37354,N_37355,N_37356,N_37357,N_37358,N_37359,N_37360,N_37361,N_37362,N_37363,N_37364,N_37365,N_37366,N_37367,N_37368,N_37369,N_37370,N_37371,N_37372,N_37373,N_37374,N_37375,N_37376,N_37377,N_37378,N_37379,N_37380,N_37381,N_37382,N_37383,N_37384,N_37385,N_37386,N_37387,N_37388,N_37389,N_37390,N_37391,N_37392,N_37393,N_37394,N_37395,N_37396,N_37397,N_37398,N_37399,N_37400,N_37401,N_37402,N_37403,N_37404,N_37405,N_37406,N_37407,N_37408,N_37409,N_37410,N_37411,N_37412,N_37413,N_37414,N_37415,N_37416,N_37417,N_37418,N_37419,N_37420,N_37421,N_37422,N_37423,N_37424,N_37425,N_37426,N_37427,N_37428,N_37429,N_37430,N_37431,N_37432,N_37433,N_37434,N_37435,N_37436,N_37437,N_37438,N_37439,N_37440,N_37441,N_37442,N_37443,N_37444,N_37445,N_37446,N_37447,N_37448,N_37449,N_37450,N_37451,N_37452,N_37453,N_37454,N_37455,N_37456,N_37457,N_37458,N_37459,N_37460,N_37461,N_37462,N_37463,N_37464,N_37465,N_37466,N_37467,N_37468,N_37469,N_37470,N_37471,N_37472,N_37473,N_37474,N_37475,N_37476,N_37477,N_37478,N_37479,N_37480,N_37481,N_37482,N_37483,N_37484,N_37485,N_37486,N_37487,N_37488,N_37489,N_37490,N_37491,N_37492,N_37493,N_37494,N_37495,N_37496,N_37497,N_37498,N_37499,N_37500,N_37501,N_37502,N_37503,N_37504,N_37505,N_37506,N_37507,N_37508,N_37509,N_37510,N_37511,N_37512,N_37513,N_37514,N_37515,N_37516,N_37517,N_37518,N_37519,N_37520,N_37521,N_37522,N_37523,N_37524,N_37525,N_37526,N_37527,N_37528,N_37529,N_37530,N_37531,N_37532,N_37533,N_37534,N_37535,N_37536,N_37537,N_37538,N_37539,N_37540,N_37541,N_37542,N_37543,N_37544,N_37545,N_37546,N_37547,N_37548,N_37549,N_37550,N_37551,N_37552,N_37553,N_37554,N_37555,N_37556,N_37557,N_37558,N_37559,N_37560,N_37561,N_37562,N_37563,N_37564,N_37565,N_37566,N_37567,N_37568,N_37569,N_37570,N_37571,N_37572,N_37573,N_37574,N_37575,N_37576,N_37577,N_37578,N_37579,N_37580,N_37581,N_37582,N_37583,N_37584,N_37585,N_37586,N_37587,N_37588,N_37589,N_37590,N_37591,N_37592,N_37593,N_37594,N_37595,N_37596,N_37597,N_37598,N_37599,N_37600,N_37601,N_37602,N_37603,N_37604,N_37605,N_37606,N_37607,N_37608,N_37609,N_37610,N_37611,N_37612,N_37613,N_37614,N_37615,N_37616,N_37617,N_37618,N_37619,N_37620,N_37621,N_37622,N_37623,N_37624,N_37625,N_37626,N_37627,N_37628,N_37629,N_37630,N_37631,N_37632,N_37633,N_37634,N_37635,N_37636,N_37637,N_37638,N_37639,N_37640,N_37641,N_37642,N_37643,N_37644,N_37645,N_37646,N_37647,N_37648,N_37649,N_37650,N_37651,N_37652,N_37653,N_37654,N_37655,N_37656,N_37657,N_37658,N_37659,N_37660,N_37661,N_37662,N_37663,N_37664,N_37665,N_37666,N_37667,N_37668,N_37669,N_37670,N_37671,N_37672,N_37673,N_37674,N_37675,N_37676,N_37677,N_37678,N_37679,N_37680,N_37681,N_37682,N_37683,N_37684,N_37685,N_37686,N_37687,N_37688,N_37689,N_37690,N_37691,N_37692,N_37693,N_37694,N_37695,N_37696,N_37697,N_37698,N_37699,N_37700,N_37701,N_37702,N_37703,N_37704,N_37705,N_37706,N_37707,N_37708,N_37709,N_37710,N_37711,N_37712,N_37713,N_37714,N_37715,N_37716,N_37717,N_37718,N_37719,N_37720,N_37721,N_37722,N_37723,N_37724,N_37725,N_37726,N_37727,N_37728,N_37729,N_37730,N_37731,N_37732,N_37733,N_37734,N_37735,N_37736,N_37737,N_37738,N_37739,N_37740,N_37741,N_37742,N_37743,N_37744,N_37745,N_37746,N_37747,N_37748,N_37749,N_37750,N_37751,N_37752,N_37753,N_37754,N_37755,N_37756,N_37757,N_37758,N_37759,N_37760,N_37761,N_37762,N_37763,N_37764,N_37765,N_37766,N_37767,N_37768,N_37769,N_37770,N_37771,N_37772,N_37773,N_37774,N_37775,N_37776,N_37777,N_37778,N_37779,N_37780,N_37781,N_37782,N_37783,N_37784,N_37785,N_37786,N_37787,N_37788,N_37789,N_37790,N_37791,N_37792,N_37793,N_37794,N_37795,N_37796,N_37797,N_37798,N_37799,N_37800,N_37801,N_37802,N_37803,N_37804,N_37805,N_37806,N_37807,N_37808,N_37809,N_37810,N_37811,N_37812,N_37813,N_37814,N_37815,N_37816,N_37817,N_37818,N_37819,N_37820,N_37821,N_37822,N_37823,N_37824,N_37825,N_37826,N_37827,N_37828,N_37829,N_37830,N_37831,N_37832,N_37833,N_37834,N_37835,N_37836,N_37837,N_37838,N_37839,N_37840,N_37841,N_37842,N_37843,N_37844,N_37845,N_37846,N_37847,N_37848,N_37849,N_37850,N_37851,N_37852,N_37853,N_37854,N_37855,N_37856,N_37857,N_37858,N_37859,N_37860,N_37861,N_37862,N_37863,N_37864,N_37865,N_37866,N_37867,N_37868,N_37869,N_37870,N_37871,N_37872,N_37873,N_37874,N_37875,N_37876,N_37877,N_37878,N_37879,N_37880,N_37881,N_37882,N_37883,N_37884,N_37885,N_37886,N_37887,N_37888,N_37889,N_37890,N_37891,N_37892,N_37893,N_37894,N_37895,N_37896,N_37897,N_37898,N_37899,N_37900,N_37901,N_37902,N_37903,N_37904,N_37905,N_37906,N_37907,N_37908,N_37909,N_37910,N_37911,N_37912,N_37913,N_37914,N_37915,N_37916,N_37917,N_37918,N_37919,N_37920,N_37921,N_37922,N_37923,N_37924,N_37925,N_37926,N_37927,N_37928,N_37929,N_37930,N_37931,N_37932,N_37933,N_37934,N_37935,N_37936,N_37937,N_37938,N_37939,N_37940,N_37941,N_37942,N_37943,N_37944,N_37945,N_37946,N_37947,N_37948,N_37949,N_37950,N_37951,N_37952,N_37953,N_37954,N_37955,N_37956,N_37957,N_37958,N_37959,N_37960,N_37961,N_37962,N_37963,N_37964,N_37965,N_37966,N_37967,N_37968,N_37969,N_37970,N_37971,N_37972,N_37973,N_37974,N_37975,N_37976,N_37977,N_37978,N_37979,N_37980,N_37981,N_37982,N_37983,N_37984,N_37985,N_37986,N_37987,N_37988,N_37989,N_37990,N_37991,N_37992,N_37993,N_37994,N_37995,N_37996,N_37997,N_37998,N_37999,N_38000,N_38001,N_38002,N_38003,N_38004,N_38005,N_38006,N_38007,N_38008,N_38009,N_38010,N_38011,N_38012,N_38013,N_38014,N_38015,N_38016,N_38017,N_38018,N_38019,N_38020,N_38021,N_38022,N_38023,N_38024,N_38025,N_38026,N_38027,N_38028,N_38029,N_38030,N_38031,N_38032,N_38033,N_38034,N_38035,N_38036,N_38037,N_38038,N_38039,N_38040,N_38041,N_38042,N_38043,N_38044,N_38045,N_38046,N_38047,N_38048,N_38049,N_38050,N_38051,N_38052,N_38053,N_38054,N_38055,N_38056,N_38057,N_38058,N_38059,N_38060,N_38061,N_38062,N_38063,N_38064,N_38065,N_38066,N_38067,N_38068,N_38069,N_38070,N_38071,N_38072,N_38073,N_38074,N_38075,N_38076,N_38077,N_38078,N_38079,N_38080,N_38081,N_38082,N_38083,N_38084,N_38085,N_38086,N_38087,N_38088,N_38089,N_38090,N_38091,N_38092,N_38093,N_38094,N_38095,N_38096,N_38097,N_38098,N_38099,N_38100,N_38101,N_38102,N_38103,N_38104,N_38105,N_38106,N_38107,N_38108,N_38109,N_38110,N_38111,N_38112,N_38113,N_38114,N_38115,N_38116,N_38117,N_38118,N_38119,N_38120,N_38121,N_38122,N_38123,N_38124,N_38125,N_38126,N_38127,N_38128,N_38129,N_38130,N_38131,N_38132,N_38133,N_38134,N_38135,N_38136,N_38137,N_38138,N_38139,N_38140,N_38141,N_38142,N_38143,N_38144,N_38145,N_38146,N_38147,N_38148,N_38149,N_38150,N_38151,N_38152,N_38153,N_38154,N_38155,N_38156,N_38157,N_38158,N_38159,N_38160,N_38161,N_38162,N_38163,N_38164,N_38165,N_38166,N_38167,N_38168,N_38169,N_38170,N_38171,N_38172,N_38173,N_38174,N_38175,N_38176,N_38177,N_38178,N_38179,N_38180,N_38181,N_38182,N_38183,N_38184,N_38185,N_38186,N_38187,N_38188,N_38189,N_38190,N_38191,N_38192,N_38193,N_38194,N_38195,N_38196,N_38197,N_38198,N_38199,N_38200,N_38201,N_38202,N_38203,N_38204,N_38205,N_38206,N_38207,N_38208,N_38209,N_38210,N_38211,N_38212,N_38213,N_38214,N_38215,N_38216,N_38217,N_38218,N_38219,N_38220,N_38221,N_38222,N_38223,N_38224,N_38225,N_38226,N_38227,N_38228,N_38229,N_38230,N_38231,N_38232,N_38233,N_38234,N_38235,N_38236,N_38237,N_38238,N_38239,N_38240,N_38241,N_38242,N_38243,N_38244,N_38245,N_38246,N_38247,N_38248,N_38249,N_38250,N_38251,N_38252,N_38253,N_38254,N_38255,N_38256,N_38257,N_38258,N_38259,N_38260,N_38261,N_38262,N_38263,N_38264,N_38265,N_38266,N_38267,N_38268,N_38269,N_38270,N_38271,N_38272,N_38273,N_38274,N_38275,N_38276,N_38277,N_38278,N_38279,N_38280,N_38281,N_38282,N_38283,N_38284,N_38285,N_38286,N_38287,N_38288,N_38289,N_38290,N_38291,N_38292,N_38293,N_38294,N_38295,N_38296,N_38297,N_38298,N_38299,N_38300,N_38301,N_38302,N_38303,N_38304,N_38305,N_38306,N_38307,N_38308,N_38309,N_38310,N_38311,N_38312,N_38313,N_38314,N_38315,N_38316,N_38317,N_38318,N_38319,N_38320,N_38321,N_38322,N_38323,N_38324,N_38325,N_38326,N_38327,N_38328,N_38329,N_38330,N_38331,N_38332,N_38333,N_38334,N_38335,N_38336,N_38337,N_38338,N_38339,N_38340,N_38341,N_38342,N_38343,N_38344,N_38345,N_38346,N_38347,N_38348,N_38349,N_38350,N_38351,N_38352,N_38353,N_38354,N_38355,N_38356,N_38357,N_38358,N_38359,N_38360,N_38361,N_38362,N_38363,N_38364,N_38365,N_38366,N_38367,N_38368,N_38369,N_38370,N_38371,N_38372,N_38373,N_38374,N_38375,N_38376,N_38377,N_38378,N_38379,N_38380,N_38381,N_38382,N_38383,N_38384,N_38385,N_38386,N_38387,N_38388,N_38389,N_38390,N_38391,N_38392,N_38393,N_38394,N_38395,N_38396,N_38397,N_38398,N_38399,N_38400,N_38401,N_38402,N_38403,N_38404,N_38405,N_38406,N_38407,N_38408,N_38409,N_38410,N_38411,N_38412,N_38413,N_38414,N_38415,N_38416,N_38417,N_38418,N_38419,N_38420,N_38421,N_38422,N_38423,N_38424,N_38425,N_38426,N_38427,N_38428,N_38429,N_38430,N_38431,N_38432,N_38433,N_38434,N_38435,N_38436,N_38437,N_38438,N_38439,N_38440,N_38441,N_38442,N_38443,N_38444,N_38445,N_38446,N_38447,N_38448,N_38449,N_38450,N_38451,N_38452,N_38453,N_38454,N_38455,N_38456,N_38457,N_38458,N_38459,N_38460,N_38461,N_38462,N_38463,N_38464,N_38465,N_38466,N_38467,N_38468,N_38469,N_38470,N_38471,N_38472,N_38473,N_38474,N_38475,N_38476,N_38477,N_38478,N_38479,N_38480,N_38481,N_38482,N_38483,N_38484,N_38485,N_38486,N_38487,N_38488,N_38489,N_38490,N_38491,N_38492,N_38493,N_38494,N_38495,N_38496,N_38497,N_38498,N_38499,N_38500,N_38501,N_38502,N_38503,N_38504,N_38505,N_38506,N_38507,N_38508,N_38509,N_38510,N_38511,N_38512,N_38513,N_38514,N_38515,N_38516,N_38517,N_38518,N_38519,N_38520,N_38521,N_38522,N_38523,N_38524,N_38525,N_38526,N_38527,N_38528,N_38529,N_38530,N_38531,N_38532,N_38533,N_38534,N_38535,N_38536,N_38537,N_38538,N_38539,N_38540,N_38541,N_38542,N_38543,N_38544,N_38545,N_38546,N_38547,N_38548,N_38549,N_38550,N_38551,N_38552,N_38553,N_38554,N_38555,N_38556,N_38557,N_38558,N_38559,N_38560,N_38561,N_38562,N_38563,N_38564,N_38565,N_38566,N_38567,N_38568,N_38569,N_38570,N_38571,N_38572,N_38573,N_38574,N_38575,N_38576,N_38577,N_38578,N_38579,N_38580,N_38581,N_38582,N_38583,N_38584,N_38585,N_38586,N_38587,N_38588,N_38589,N_38590,N_38591,N_38592,N_38593,N_38594,N_38595,N_38596,N_38597,N_38598,N_38599,N_38600,N_38601,N_38602,N_38603,N_38604,N_38605,N_38606,N_38607,N_38608,N_38609,N_38610,N_38611,N_38612,N_38613,N_38614,N_38615,N_38616,N_38617,N_38618,N_38619,N_38620,N_38621,N_38622,N_38623,N_38624,N_38625,N_38626,N_38627,N_38628,N_38629,N_38630,N_38631,N_38632,N_38633,N_38634,N_38635,N_38636,N_38637,N_38638,N_38639,N_38640,N_38641,N_38642,N_38643,N_38644,N_38645,N_38646,N_38647,N_38648,N_38649,N_38650,N_38651,N_38652,N_38653,N_38654,N_38655,N_38656,N_38657,N_38658,N_38659,N_38660,N_38661,N_38662,N_38663,N_38664,N_38665,N_38666,N_38667,N_38668,N_38669,N_38670,N_38671,N_38672,N_38673,N_38674,N_38675,N_38676,N_38677,N_38678,N_38679,N_38680,N_38681,N_38682,N_38683,N_38684,N_38685,N_38686,N_38687,N_38688,N_38689,N_38690,N_38691,N_38692,N_38693,N_38694,N_38695,N_38696,N_38697,N_38698,N_38699,N_38700,N_38701,N_38702,N_38703,N_38704,N_38705,N_38706,N_38707,N_38708,N_38709,N_38710,N_38711,N_38712,N_38713,N_38714,N_38715,N_38716,N_38717,N_38718,N_38719,N_38720,N_38721,N_38722,N_38723,N_38724,N_38725,N_38726,N_38727,N_38728,N_38729,N_38730,N_38731,N_38732,N_38733,N_38734,N_38735,N_38736,N_38737,N_38738,N_38739,N_38740,N_38741,N_38742,N_38743,N_38744,N_38745,N_38746,N_38747,N_38748,N_38749,N_38750,N_38751,N_38752,N_38753,N_38754,N_38755,N_38756,N_38757,N_38758,N_38759,N_38760,N_38761,N_38762,N_38763,N_38764,N_38765,N_38766,N_38767,N_38768,N_38769,N_38770,N_38771,N_38772,N_38773,N_38774,N_38775,N_38776,N_38777,N_38778,N_38779,N_38780,N_38781,N_38782,N_38783,N_38784,N_38785,N_38786,N_38787,N_38788,N_38789,N_38790,N_38791,N_38792,N_38793,N_38794,N_38795,N_38796,N_38797,N_38798,N_38799,N_38800,N_38801,N_38802,N_38803,N_38804,N_38805,N_38806,N_38807,N_38808,N_38809,N_38810,N_38811,N_38812,N_38813,N_38814,N_38815,N_38816,N_38817,N_38818,N_38819,N_38820,N_38821,N_38822,N_38823,N_38824,N_38825,N_38826,N_38827,N_38828,N_38829,N_38830,N_38831,N_38832,N_38833,N_38834,N_38835,N_38836,N_38837,N_38838,N_38839,N_38840,N_38841,N_38842,N_38843,N_38844,N_38845,N_38846,N_38847,N_38848,N_38849,N_38850,N_38851,N_38852,N_38853,N_38854,N_38855,N_38856,N_38857,N_38858,N_38859,N_38860,N_38861,N_38862,N_38863,N_38864,N_38865,N_38866,N_38867,N_38868,N_38869,N_38870,N_38871,N_38872,N_38873,N_38874,N_38875,N_38876,N_38877,N_38878,N_38879,N_38880,N_38881,N_38882,N_38883,N_38884,N_38885,N_38886,N_38887,N_38888,N_38889,N_38890,N_38891,N_38892,N_38893,N_38894,N_38895,N_38896,N_38897,N_38898,N_38899,N_38900,N_38901,N_38902,N_38903,N_38904,N_38905,N_38906,N_38907,N_38908,N_38909,N_38910,N_38911,N_38912,N_38913,N_38914,N_38915,N_38916,N_38917,N_38918,N_38919,N_38920,N_38921,N_38922,N_38923,N_38924,N_38925,N_38926,N_38927,N_38928,N_38929,N_38930,N_38931,N_38932,N_38933,N_38934,N_38935,N_38936,N_38937,N_38938,N_38939,N_38940,N_38941,N_38942,N_38943,N_38944,N_38945,N_38946,N_38947,N_38948,N_38949,N_38950,N_38951,N_38952,N_38953,N_38954,N_38955,N_38956,N_38957,N_38958,N_38959,N_38960,N_38961,N_38962,N_38963,N_38964,N_38965,N_38966,N_38967,N_38968,N_38969,N_38970,N_38971,N_38972,N_38973,N_38974,N_38975,N_38976,N_38977,N_38978,N_38979,N_38980,N_38981,N_38982,N_38983,N_38984,N_38985,N_38986,N_38987,N_38988,N_38989,N_38990,N_38991,N_38992,N_38993,N_38994,N_38995,N_38996,N_38997,N_38998,N_38999,N_39000,N_39001,N_39002,N_39003,N_39004,N_39005,N_39006,N_39007,N_39008,N_39009,N_39010,N_39011,N_39012,N_39013,N_39014,N_39015,N_39016,N_39017,N_39018,N_39019,N_39020,N_39021,N_39022,N_39023,N_39024,N_39025,N_39026,N_39027,N_39028,N_39029,N_39030,N_39031,N_39032,N_39033,N_39034,N_39035,N_39036,N_39037,N_39038,N_39039,N_39040,N_39041,N_39042,N_39043,N_39044,N_39045,N_39046,N_39047,N_39048,N_39049,N_39050,N_39051,N_39052,N_39053,N_39054,N_39055,N_39056,N_39057,N_39058,N_39059,N_39060,N_39061,N_39062,N_39063,N_39064,N_39065,N_39066,N_39067,N_39068,N_39069,N_39070,N_39071,N_39072,N_39073,N_39074,N_39075,N_39076,N_39077,N_39078,N_39079,N_39080,N_39081,N_39082,N_39083,N_39084,N_39085,N_39086,N_39087,N_39088,N_39089,N_39090,N_39091,N_39092,N_39093,N_39094,N_39095,N_39096,N_39097,N_39098,N_39099,N_39100,N_39101,N_39102,N_39103,N_39104,N_39105,N_39106,N_39107,N_39108,N_39109,N_39110,N_39111,N_39112,N_39113,N_39114,N_39115,N_39116,N_39117,N_39118,N_39119,N_39120,N_39121,N_39122,N_39123,N_39124,N_39125,N_39126,N_39127,N_39128,N_39129,N_39130,N_39131,N_39132,N_39133,N_39134,N_39135,N_39136,N_39137,N_39138,N_39139,N_39140,N_39141,N_39142,N_39143,N_39144,N_39145,N_39146,N_39147,N_39148,N_39149,N_39150,N_39151,N_39152,N_39153,N_39154,N_39155,N_39156,N_39157,N_39158,N_39159,N_39160,N_39161,N_39162,N_39163,N_39164,N_39165,N_39166,N_39167,N_39168,N_39169,N_39170,N_39171,N_39172,N_39173,N_39174,N_39175,N_39176,N_39177,N_39178,N_39179,N_39180,N_39181,N_39182,N_39183,N_39184,N_39185,N_39186,N_39187,N_39188,N_39189,N_39190,N_39191,N_39192,N_39193,N_39194,N_39195,N_39196,N_39197,N_39198,N_39199,N_39200,N_39201,N_39202,N_39203,N_39204,N_39205,N_39206,N_39207,N_39208,N_39209,N_39210,N_39211,N_39212,N_39213,N_39214,N_39215,N_39216,N_39217,N_39218,N_39219,N_39220,N_39221,N_39222,N_39223,N_39224,N_39225,N_39226,N_39227,N_39228,N_39229,N_39230,N_39231,N_39232,N_39233,N_39234,N_39235,N_39236,N_39237,N_39238,N_39239,N_39240,N_39241,N_39242,N_39243,N_39244,N_39245,N_39246,N_39247,N_39248,N_39249,N_39250,N_39251,N_39252,N_39253,N_39254,N_39255,N_39256,N_39257,N_39258,N_39259,N_39260,N_39261,N_39262,N_39263,N_39264,N_39265,N_39266,N_39267,N_39268,N_39269,N_39270,N_39271,N_39272,N_39273,N_39274,N_39275,N_39276,N_39277,N_39278,N_39279,N_39280,N_39281,N_39282,N_39283,N_39284,N_39285,N_39286,N_39287,N_39288,N_39289,N_39290,N_39291,N_39292,N_39293,N_39294,N_39295,N_39296,N_39297,N_39298,N_39299,N_39300,N_39301,N_39302,N_39303,N_39304,N_39305,N_39306,N_39307,N_39308,N_39309,N_39310,N_39311,N_39312,N_39313,N_39314,N_39315,N_39316,N_39317,N_39318,N_39319,N_39320,N_39321,N_39322,N_39323,N_39324,N_39325,N_39326,N_39327,N_39328,N_39329,N_39330,N_39331,N_39332,N_39333,N_39334,N_39335,N_39336,N_39337,N_39338,N_39339,N_39340,N_39341,N_39342,N_39343,N_39344,N_39345,N_39346,N_39347,N_39348,N_39349,N_39350,N_39351,N_39352,N_39353,N_39354,N_39355,N_39356,N_39357,N_39358,N_39359,N_39360,N_39361,N_39362,N_39363,N_39364,N_39365,N_39366,N_39367,N_39368,N_39369,N_39370,N_39371,N_39372,N_39373,N_39374,N_39375,N_39376,N_39377,N_39378,N_39379,N_39380,N_39381,N_39382,N_39383,N_39384,N_39385,N_39386,N_39387,N_39388,N_39389,N_39390,N_39391,N_39392,N_39393,N_39394,N_39395,N_39396,N_39397,N_39398,N_39399,N_39400,N_39401,N_39402,N_39403,N_39404,N_39405,N_39406,N_39407,N_39408,N_39409,N_39410,N_39411,N_39412,N_39413,N_39414,N_39415,N_39416,N_39417,N_39418,N_39419,N_39420,N_39421,N_39422,N_39423,N_39424,N_39425,N_39426,N_39427,N_39428,N_39429,N_39430,N_39431,N_39432,N_39433,N_39434,N_39435,N_39436,N_39437,N_39438,N_39439,N_39440,N_39441,N_39442,N_39443,N_39444,N_39445,N_39446,N_39447,N_39448,N_39449,N_39450,N_39451,N_39452,N_39453,N_39454,N_39455,N_39456,N_39457,N_39458,N_39459,N_39460,N_39461,N_39462,N_39463,N_39464,N_39465,N_39466,N_39467,N_39468,N_39469,N_39470,N_39471,N_39472,N_39473,N_39474,N_39475,N_39476,N_39477,N_39478,N_39479,N_39480,N_39481,N_39482,N_39483,N_39484,N_39485,N_39486,N_39487,N_39488,N_39489,N_39490,N_39491,N_39492,N_39493,N_39494,N_39495,N_39496,N_39497,N_39498,N_39499,N_39500,N_39501,N_39502,N_39503,N_39504,N_39505,N_39506,N_39507,N_39508,N_39509,N_39510,N_39511,N_39512,N_39513,N_39514,N_39515,N_39516,N_39517,N_39518,N_39519,N_39520,N_39521,N_39522,N_39523,N_39524,N_39525,N_39526,N_39527,N_39528,N_39529,N_39530,N_39531,N_39532,N_39533,N_39534,N_39535,N_39536,N_39537,N_39538,N_39539,N_39540,N_39541,N_39542,N_39543,N_39544,N_39545,N_39546,N_39547,N_39548,N_39549,N_39550,N_39551,N_39552,N_39553,N_39554,N_39555,N_39556,N_39557,N_39558,N_39559,N_39560,N_39561,N_39562,N_39563,N_39564,N_39565,N_39566,N_39567,N_39568,N_39569,N_39570,N_39571,N_39572,N_39573,N_39574,N_39575,N_39576,N_39577,N_39578,N_39579,N_39580,N_39581,N_39582,N_39583,N_39584,N_39585,N_39586,N_39587,N_39588,N_39589,N_39590,N_39591,N_39592,N_39593,N_39594,N_39595,N_39596,N_39597,N_39598,N_39599,N_39600,N_39601,N_39602,N_39603,N_39604,N_39605,N_39606,N_39607,N_39608,N_39609,N_39610,N_39611,N_39612,N_39613,N_39614,N_39615,N_39616,N_39617,N_39618,N_39619,N_39620,N_39621,N_39622,N_39623,N_39624,N_39625,N_39626,N_39627,N_39628,N_39629,N_39630,N_39631,N_39632,N_39633,N_39634,N_39635,N_39636,N_39637,N_39638,N_39639,N_39640,N_39641,N_39642,N_39643,N_39644,N_39645,N_39646,N_39647,N_39648,N_39649,N_39650,N_39651,N_39652,N_39653,N_39654,N_39655,N_39656,N_39657,N_39658,N_39659,N_39660,N_39661,N_39662,N_39663,N_39664,N_39665,N_39666,N_39667,N_39668,N_39669,N_39670,N_39671,N_39672,N_39673,N_39674,N_39675,N_39676,N_39677,N_39678,N_39679,N_39680,N_39681,N_39682,N_39683,N_39684,N_39685,N_39686,N_39687,N_39688,N_39689,N_39690,N_39691,N_39692,N_39693,N_39694,N_39695,N_39696,N_39697,N_39698,N_39699,N_39700,N_39701,N_39702,N_39703,N_39704,N_39705,N_39706,N_39707,N_39708,N_39709,N_39710,N_39711,N_39712,N_39713,N_39714,N_39715,N_39716,N_39717,N_39718,N_39719,N_39720,N_39721,N_39722,N_39723,N_39724,N_39725,N_39726,N_39727,N_39728,N_39729,N_39730,N_39731,N_39732,N_39733,N_39734,N_39735,N_39736,N_39737,N_39738,N_39739,N_39740,N_39741,N_39742,N_39743,N_39744,N_39745,N_39746,N_39747,N_39748,N_39749,N_39750,N_39751,N_39752,N_39753,N_39754,N_39755,N_39756,N_39757,N_39758,N_39759,N_39760,N_39761,N_39762,N_39763,N_39764,N_39765,N_39766,N_39767,N_39768,N_39769,N_39770,N_39771,N_39772,N_39773,N_39774,N_39775,N_39776,N_39777,N_39778,N_39779,N_39780,N_39781,N_39782,N_39783,N_39784,N_39785,N_39786,N_39787,N_39788,N_39789,N_39790,N_39791,N_39792,N_39793,N_39794,N_39795,N_39796,N_39797,N_39798,N_39799,N_39800,N_39801,N_39802,N_39803,N_39804,N_39805,N_39806,N_39807,N_39808,N_39809,N_39810,N_39811,N_39812,N_39813,N_39814,N_39815,N_39816,N_39817,N_39818,N_39819,N_39820,N_39821,N_39822,N_39823,N_39824,N_39825,N_39826,N_39827,N_39828,N_39829,N_39830,N_39831,N_39832,N_39833,N_39834,N_39835,N_39836,N_39837,N_39838,N_39839,N_39840,N_39841,N_39842,N_39843,N_39844,N_39845,N_39846,N_39847,N_39848,N_39849,N_39850,N_39851,N_39852,N_39853,N_39854,N_39855,N_39856,N_39857,N_39858,N_39859,N_39860,N_39861,N_39862,N_39863,N_39864,N_39865,N_39866,N_39867,N_39868,N_39869,N_39870,N_39871,N_39872,N_39873,N_39874,N_39875,N_39876,N_39877,N_39878,N_39879,N_39880,N_39881,N_39882,N_39883,N_39884,N_39885,N_39886,N_39887,N_39888,N_39889,N_39890,N_39891,N_39892,N_39893,N_39894,N_39895,N_39896,N_39897,N_39898,N_39899,N_39900,N_39901,N_39902,N_39903,N_39904,N_39905,N_39906,N_39907,N_39908,N_39909,N_39910,N_39911,N_39912,N_39913,N_39914,N_39915,N_39916,N_39917,N_39918,N_39919,N_39920,N_39921,N_39922,N_39923,N_39924,N_39925,N_39926,N_39927,N_39928,N_39929,N_39930,N_39931,N_39932,N_39933,N_39934,N_39935,N_39936,N_39937,N_39938,N_39939,N_39940,N_39941,N_39942,N_39943,N_39944,N_39945,N_39946,N_39947,N_39948,N_39949,N_39950,N_39951,N_39952,N_39953,N_39954,N_39955,N_39956,N_39957,N_39958,N_39959,N_39960,N_39961,N_39962,N_39963,N_39964,N_39965,N_39966,N_39967,N_39968,N_39969,N_39970,N_39971,N_39972,N_39973,N_39974,N_39975,N_39976,N_39977,N_39978,N_39979,N_39980,N_39981,N_39982,N_39983,N_39984,N_39985,N_39986,N_39987,N_39988,N_39989,N_39990,N_39991,N_39992,N_39993,N_39994,N_39995,N_39996,N_39997,N_39998,N_39999,N_40000,N_40001,N_40002,N_40003,N_40004,N_40005,N_40006,N_40007,N_40008,N_40009,N_40010,N_40011,N_40012,N_40013,N_40014,N_40015,N_40016,N_40017,N_40018,N_40019,N_40020,N_40021,N_40022,N_40023,N_40024,N_40025,N_40026,N_40027,N_40028,N_40029,N_40030,N_40031,N_40032,N_40033,N_40034,N_40035,N_40036,N_40037,N_40038,N_40039,N_40040,N_40041,N_40042,N_40043,N_40044,N_40045,N_40046,N_40047,N_40048,N_40049,N_40050,N_40051,N_40052,N_40053,N_40054,N_40055,N_40056,N_40057,N_40058,N_40059,N_40060,N_40061,N_40062,N_40063,N_40064,N_40065,N_40066,N_40067,N_40068,N_40069,N_40070,N_40071,N_40072,N_40073,N_40074,N_40075,N_40076,N_40077,N_40078,N_40079,N_40080,N_40081,N_40082,N_40083,N_40084,N_40085,N_40086,N_40087,N_40088,N_40089,N_40090,N_40091,N_40092,N_40093,N_40094,N_40095,N_40096,N_40097,N_40098,N_40099,N_40100,N_40101,N_40102,N_40103,N_40104,N_40105,N_40106,N_40107,N_40108,N_40109,N_40110,N_40111,N_40112,N_40113,N_40114,N_40115,N_40116,N_40117,N_40118,N_40119,N_40120,N_40121,N_40122,N_40123,N_40124,N_40125,N_40126,N_40127,N_40128,N_40129,N_40130,N_40131,N_40132,N_40133,N_40134,N_40135,N_40136,N_40137,N_40138,N_40139,N_40140,N_40141,N_40142,N_40143,N_40144,N_40145,N_40146,N_40147,N_40148,N_40149,N_40150,N_40151,N_40152,N_40153,N_40154,N_40155,N_40156,N_40157,N_40158,N_40159,N_40160,N_40161,N_40162,N_40163,N_40164,N_40165,N_40166,N_40167,N_40168,N_40169,N_40170,N_40171,N_40172,N_40173,N_40174,N_40175,N_40176,N_40177,N_40178,N_40179,N_40180,N_40181,N_40182,N_40183,N_40184,N_40185,N_40186,N_40187,N_40188,N_40189,N_40190,N_40191,N_40192,N_40193,N_40194,N_40195,N_40196,N_40197,N_40198,N_40199,N_40200,N_40201,N_40202,N_40203,N_40204,N_40205,N_40206,N_40207,N_40208,N_40209,N_40210,N_40211,N_40212,N_40213,N_40214,N_40215,N_40216,N_40217,N_40218,N_40219,N_40220,N_40221,N_40222,N_40223,N_40224,N_40225,N_40226,N_40227,N_40228,N_40229,N_40230,N_40231,N_40232,N_40233,N_40234,N_40235,N_40236,N_40237,N_40238,N_40239,N_40240,N_40241,N_40242,N_40243,N_40244,N_40245,N_40246,N_40247,N_40248,N_40249,N_40250,N_40251,N_40252,N_40253,N_40254,N_40255,N_40256,N_40257,N_40258,N_40259,N_40260,N_40261,N_40262,N_40263,N_40264,N_40265,N_40266,N_40267,N_40268,N_40269,N_40270,N_40271,N_40272,N_40273,N_40274,N_40275,N_40276,N_40277,N_40278,N_40279,N_40280,N_40281,N_40282,N_40283,N_40284,N_40285,N_40286,N_40287,N_40288,N_40289,N_40290,N_40291,N_40292,N_40293,N_40294,N_40295,N_40296,N_40297,N_40298,N_40299,N_40300,N_40301,N_40302,N_40303,N_40304,N_40305,N_40306,N_40307,N_40308,N_40309,N_40310,N_40311,N_40312,N_40313,N_40314,N_40315,N_40316,N_40317,N_40318,N_40319,N_40320,N_40321,N_40322,N_40323,N_40324,N_40325,N_40326,N_40327,N_40328,N_40329,N_40330,N_40331,N_40332,N_40333,N_40334,N_40335,N_40336,N_40337,N_40338,N_40339,N_40340,N_40341,N_40342,N_40343,N_40344,N_40345,N_40346,N_40347,N_40348,N_40349,N_40350,N_40351,N_40352,N_40353,N_40354,N_40355,N_40356,N_40357,N_40358,N_40359,N_40360,N_40361,N_40362,N_40363,N_40364,N_40365,N_40366,N_40367,N_40368,N_40369,N_40370,N_40371,N_40372,N_40373,N_40374,N_40375,N_40376,N_40377,N_40378,N_40379,N_40380,N_40381,N_40382,N_40383,N_40384,N_40385,N_40386,N_40387,N_40388,N_40389,N_40390,N_40391,N_40392,N_40393,N_40394,N_40395,N_40396,N_40397,N_40398,N_40399,N_40400,N_40401,N_40402,N_40403,N_40404,N_40405,N_40406,N_40407,N_40408,N_40409,N_40410,N_40411,N_40412,N_40413,N_40414,N_40415,N_40416,N_40417,N_40418,N_40419,N_40420,N_40421,N_40422,N_40423,N_40424,N_40425,N_40426,N_40427,N_40428,N_40429,N_40430,N_40431,N_40432,N_40433,N_40434,N_40435,N_40436,N_40437,N_40438,N_40439,N_40440,N_40441,N_40442,N_40443,N_40444,N_40445,N_40446,N_40447,N_40448,N_40449,N_40450,N_40451,N_40452,N_40453,N_40454,N_40455,N_40456,N_40457,N_40458,N_40459,N_40460,N_40461,N_40462,N_40463,N_40464,N_40465,N_40466,N_40467,N_40468,N_40469,N_40470,N_40471,N_40472,N_40473,N_40474,N_40475,N_40476,N_40477,N_40478,N_40479,N_40480,N_40481,N_40482,N_40483,N_40484,N_40485,N_40486,N_40487,N_40488,N_40489,N_40490,N_40491,N_40492,N_40493,N_40494,N_40495,N_40496,N_40497,N_40498,N_40499,N_40500,N_40501,N_40502,N_40503,N_40504,N_40505,N_40506,N_40507,N_40508,N_40509,N_40510,N_40511,N_40512,N_40513,N_40514,N_40515,N_40516,N_40517,N_40518,N_40519,N_40520,N_40521,N_40522,N_40523,N_40524,N_40525,N_40526,N_40527,N_40528,N_40529,N_40530,N_40531,N_40532,N_40533,N_40534,N_40535,N_40536,N_40537,N_40538,N_40539,N_40540,N_40541,N_40542,N_40543,N_40544,N_40545,N_40546,N_40547,N_40548,N_40549,N_40550,N_40551,N_40552,N_40553,N_40554,N_40555,N_40556,N_40557,N_40558,N_40559,N_40560,N_40561,N_40562,N_40563,N_40564,N_40565,N_40566,N_40567,N_40568,N_40569,N_40570,N_40571,N_40572,N_40573,N_40574,N_40575,N_40576,N_40577,N_40578,N_40579,N_40580,N_40581,N_40582,N_40583,N_40584,N_40585,N_40586,N_40587,N_40588,N_40589,N_40590,N_40591,N_40592,N_40593,N_40594,N_40595,N_40596,N_40597,N_40598,N_40599,N_40600,N_40601,N_40602,N_40603,N_40604,N_40605,N_40606,N_40607,N_40608,N_40609,N_40610,N_40611,N_40612,N_40613,N_40614,N_40615,N_40616,N_40617,N_40618,N_40619,N_40620,N_40621,N_40622,N_40623,N_40624,N_40625,N_40626,N_40627,N_40628,N_40629,N_40630,N_40631,N_40632,N_40633,N_40634,N_40635,N_40636,N_40637,N_40638,N_40639,N_40640,N_40641,N_40642,N_40643,N_40644,N_40645,N_40646,N_40647,N_40648,N_40649,N_40650,N_40651,N_40652,N_40653,N_40654,N_40655,N_40656,N_40657,N_40658,N_40659,N_40660,N_40661,N_40662,N_40663,N_40664,N_40665,N_40666,N_40667,N_40668,N_40669,N_40670,N_40671,N_40672,N_40673,N_40674,N_40675,N_40676,N_40677,N_40678,N_40679,N_40680,N_40681,N_40682,N_40683,N_40684,N_40685,N_40686,N_40687,N_40688,N_40689,N_40690,N_40691,N_40692,N_40693,N_40694,N_40695,N_40696,N_40697,N_40698,N_40699,N_40700,N_40701,N_40702,N_40703,N_40704,N_40705,N_40706,N_40707,N_40708,N_40709,N_40710,N_40711,N_40712,N_40713,N_40714,N_40715,N_40716,N_40717,N_40718,N_40719,N_40720,N_40721,N_40722,N_40723,N_40724,N_40725,N_40726,N_40727,N_40728,N_40729,N_40730,N_40731,N_40732,N_40733,N_40734,N_40735,N_40736,N_40737,N_40738,N_40739,N_40740,N_40741,N_40742,N_40743,N_40744,N_40745,N_40746,N_40747,N_40748,N_40749,N_40750,N_40751,N_40752,N_40753,N_40754,N_40755,N_40756,N_40757,N_40758,N_40759,N_40760,N_40761,N_40762,N_40763,N_40764,N_40765,N_40766,N_40767,N_40768,N_40769,N_40770,N_40771,N_40772,N_40773,N_40774,N_40775,N_40776,N_40777,N_40778,N_40779,N_40780,N_40781,N_40782,N_40783,N_40784,N_40785,N_40786,N_40787,N_40788,N_40789,N_40790,N_40791,N_40792,N_40793,N_40794,N_40795,N_40796,N_40797,N_40798,N_40799,N_40800,N_40801,N_40802,N_40803,N_40804,N_40805,N_40806,N_40807,N_40808,N_40809,N_40810,N_40811,N_40812,N_40813,N_40814,N_40815,N_40816,N_40817,N_40818,N_40819,N_40820,N_40821,N_40822,N_40823,N_40824,N_40825,N_40826,N_40827,N_40828,N_40829,N_40830,N_40831,N_40832,N_40833,N_40834,N_40835,N_40836,N_40837,N_40838,N_40839,N_40840,N_40841,N_40842,N_40843,N_40844,N_40845,N_40846,N_40847,N_40848,N_40849,N_40850,N_40851,N_40852,N_40853,N_40854,N_40855,N_40856,N_40857,N_40858,N_40859,N_40860,N_40861,N_40862,N_40863,N_40864,N_40865,N_40866,N_40867,N_40868,N_40869,N_40870,N_40871,N_40872,N_40873,N_40874,N_40875,N_40876,N_40877,N_40878,N_40879,N_40880,N_40881,N_40882,N_40883,N_40884,N_40885,N_40886,N_40887,N_40888,N_40889,N_40890,N_40891,N_40892,N_40893,N_40894,N_40895,N_40896,N_40897,N_40898,N_40899,N_40900,N_40901,N_40902,N_40903,N_40904,N_40905,N_40906,N_40907,N_40908,N_40909,N_40910,N_40911,N_40912,N_40913,N_40914,N_40915,N_40916,N_40917,N_40918,N_40919,N_40920,N_40921,N_40922,N_40923,N_40924,N_40925,N_40926,N_40927,N_40928,N_40929,N_40930,N_40931,N_40932,N_40933,N_40934,N_40935,N_40936,N_40937,N_40938,N_40939,N_40940,N_40941,N_40942,N_40943,N_40944,N_40945,N_40946,N_40947,N_40948,N_40949,N_40950,N_40951,N_40952,N_40953,N_40954,N_40955,N_40956,N_40957,N_40958,N_40959,N_40960,N_40961,N_40962,N_40963,N_40964,N_40965,N_40966,N_40967,N_40968,N_40969,N_40970,N_40971,N_40972,N_40973,N_40974,N_40975,N_40976,N_40977,N_40978,N_40979,N_40980,N_40981,N_40982,N_40983,N_40984,N_40985,N_40986,N_40987,N_40988,N_40989,N_40990,N_40991,N_40992,N_40993,N_40994,N_40995,N_40996,N_40997,N_40998,N_40999,N_41000,N_41001,N_41002,N_41003,N_41004,N_41005,N_41006,N_41007,N_41008,N_41009,N_41010,N_41011,N_41012,N_41013,N_41014,N_41015,N_41016,N_41017,N_41018,N_41019,N_41020,N_41021,N_41022,N_41023,N_41024,N_41025,N_41026,N_41027,N_41028,N_41029,N_41030,N_41031,N_41032,N_41033,N_41034,N_41035,N_41036,N_41037,N_41038,N_41039,N_41040,N_41041,N_41042,N_41043,N_41044,N_41045,N_41046,N_41047,N_41048,N_41049,N_41050,N_41051,N_41052,N_41053,N_41054,N_41055,N_41056,N_41057,N_41058,N_41059,N_41060,N_41061,N_41062,N_41063,N_41064,N_41065,N_41066,N_41067,N_41068,N_41069,N_41070,N_41071,N_41072,N_41073,N_41074,N_41075,N_41076,N_41077,N_41078,N_41079,N_41080,N_41081,N_41082,N_41083,N_41084,N_41085,N_41086,N_41087,N_41088,N_41089,N_41090,N_41091,N_41092,N_41093,N_41094,N_41095,N_41096,N_41097,N_41098,N_41099,N_41100,N_41101,N_41102,N_41103,N_41104,N_41105,N_41106,N_41107,N_41108,N_41109,N_41110,N_41111,N_41112,N_41113,N_41114,N_41115,N_41116,N_41117,N_41118,N_41119,N_41120,N_41121,N_41122,N_41123,N_41124,N_41125,N_41126,N_41127,N_41128,N_41129,N_41130,N_41131,N_41132,N_41133,N_41134,N_41135,N_41136,N_41137,N_41138,N_41139,N_41140,N_41141,N_41142,N_41143,N_41144,N_41145,N_41146,N_41147,N_41148,N_41149,N_41150,N_41151,N_41152,N_41153,N_41154,N_41155,N_41156,N_41157,N_41158,N_41159,N_41160,N_41161,N_41162,N_41163,N_41164,N_41165,N_41166,N_41167,N_41168,N_41169,N_41170,N_41171,N_41172,N_41173,N_41174,N_41175,N_41176,N_41177,N_41178,N_41179,N_41180,N_41181,N_41182,N_41183,N_41184,N_41185,N_41186,N_41187,N_41188,N_41189,N_41190,N_41191,N_41192,N_41193,N_41194,N_41195,N_41196,N_41197,N_41198,N_41199,N_41200,N_41201,N_41202,N_41203,N_41204,N_41205,N_41206,N_41207,N_41208,N_41209,N_41210,N_41211,N_41212,N_41213,N_41214,N_41215,N_41216,N_41217,N_41218,N_41219,N_41220,N_41221,N_41222,N_41223,N_41224,N_41225,N_41226,N_41227,N_41228,N_41229,N_41230,N_41231,N_41232,N_41233,N_41234,N_41235,N_41236,N_41237,N_41238,N_41239,N_41240,N_41241,N_41242,N_41243,N_41244,N_41245,N_41246,N_41247,N_41248,N_41249,N_41250,N_41251,N_41252,N_41253,N_41254,N_41255,N_41256,N_41257,N_41258,N_41259,N_41260,N_41261,N_41262,N_41263,N_41264,N_41265,N_41266,N_41267,N_41268,N_41269,N_41270,N_41271,N_41272,N_41273,N_41274,N_41275,N_41276,N_41277,N_41278,N_41279,N_41280,N_41281,N_41282,N_41283,N_41284,N_41285,N_41286,N_41287,N_41288,N_41289,N_41290,N_41291,N_41292,N_41293,N_41294,N_41295,N_41296,N_41297,N_41298,N_41299,N_41300,N_41301,N_41302,N_41303,N_41304,N_41305,N_41306,N_41307,N_41308,N_41309,N_41310,N_41311,N_41312,N_41313,N_41314,N_41315,N_41316,N_41317,N_41318,N_41319,N_41320,N_41321,N_41322,N_41323,N_41324,N_41325,N_41326,N_41327,N_41328,N_41329,N_41330,N_41331,N_41332,N_41333,N_41334,N_41335,N_41336,N_41337,N_41338,N_41339,N_41340,N_41341,N_41342,N_41343,N_41344,N_41345,N_41346,N_41347,N_41348,N_41349,N_41350,N_41351,N_41352,N_41353,N_41354,N_41355,N_41356,N_41357,N_41358,N_41359,N_41360,N_41361,N_41362,N_41363,N_41364,N_41365,N_41366,N_41367,N_41368,N_41369,N_41370,N_41371,N_41372,N_41373,N_41374,N_41375,N_41376,N_41377,N_41378,N_41379,N_41380,N_41381,N_41382,N_41383,N_41384,N_41385,N_41386,N_41387,N_41388,N_41389,N_41390,N_41391,N_41392,N_41393,N_41394,N_41395,N_41396,N_41397,N_41398,N_41399,N_41400,N_41401,N_41402,N_41403,N_41404,N_41405,N_41406,N_41407,N_41408,N_41409,N_41410,N_41411,N_41412,N_41413,N_41414,N_41415,N_41416,N_41417,N_41418,N_41419,N_41420,N_41421,N_41422,N_41423,N_41424,N_41425,N_41426,N_41427,N_41428,N_41429,N_41430,N_41431,N_41432,N_41433,N_41434,N_41435,N_41436,N_41437,N_41438,N_41439,N_41440,N_41441,N_41442,N_41443,N_41444,N_41445,N_41446,N_41447,N_41448,N_41449,N_41450,N_41451,N_41452,N_41453,N_41454,N_41455,N_41456,N_41457,N_41458,N_41459,N_41460,N_41461,N_41462,N_41463,N_41464,N_41465,N_41466,N_41467,N_41468,N_41469,N_41470,N_41471,N_41472,N_41473,N_41474,N_41475,N_41476,N_41477,N_41478,N_41479,N_41480,N_41481,N_41482,N_41483,N_41484,N_41485,N_41486,N_41487,N_41488,N_41489,N_41490,N_41491,N_41492,N_41493,N_41494,N_41495,N_41496,N_41497,N_41498,N_41499,N_41500,N_41501,N_41502,N_41503,N_41504,N_41505,N_41506,N_41507,N_41508,N_41509,N_41510,N_41511,N_41512,N_41513,N_41514,N_41515,N_41516,N_41517,N_41518,N_41519,N_41520,N_41521,N_41522,N_41523,N_41524,N_41525,N_41526,N_41527,N_41528,N_41529,N_41530,N_41531,N_41532,N_41533,N_41534,N_41535,N_41536,N_41537,N_41538,N_41539,N_41540,N_41541,N_41542,N_41543,N_41544,N_41545,N_41546,N_41547,N_41548,N_41549,N_41550,N_41551,N_41552,N_41553,N_41554,N_41555,N_41556,N_41557,N_41558,N_41559,N_41560,N_41561,N_41562,N_41563,N_41564,N_41565,N_41566,N_41567,N_41568,N_41569,N_41570,N_41571,N_41572,N_41573,N_41574,N_41575,N_41576,N_41577,N_41578,N_41579,N_41580,N_41581,N_41582,N_41583,N_41584,N_41585,N_41586,N_41587,N_41588,N_41589,N_41590,N_41591,N_41592,N_41593,N_41594,N_41595,N_41596,N_41597,N_41598,N_41599,N_41600,N_41601,N_41602,N_41603,N_41604,N_41605,N_41606,N_41607,N_41608,N_41609,N_41610,N_41611,N_41612,N_41613,N_41614,N_41615,N_41616,N_41617,N_41618,N_41619,N_41620,N_41621,N_41622,N_41623,N_41624,N_41625,N_41626,N_41627,N_41628,N_41629,N_41630,N_41631,N_41632,N_41633,N_41634,N_41635,N_41636,N_41637,N_41638,N_41639,N_41640,N_41641,N_41642,N_41643,N_41644,N_41645,N_41646,N_41647,N_41648,N_41649,N_41650,N_41651,N_41652,N_41653,N_41654,N_41655,N_41656,N_41657,N_41658,N_41659,N_41660,N_41661,N_41662,N_41663,N_41664,N_41665,N_41666,N_41667,N_41668,N_41669,N_41670,N_41671,N_41672,N_41673,N_41674,N_41675,N_41676,N_41677,N_41678,N_41679,N_41680,N_41681,N_41682,N_41683,N_41684,N_41685,N_41686,N_41687,N_41688,N_41689,N_41690,N_41691,N_41692,N_41693,N_41694,N_41695,N_41696,N_41697,N_41698,N_41699,N_41700,N_41701,N_41702,N_41703,N_41704,N_41705,N_41706,N_41707,N_41708,N_41709,N_41710,N_41711,N_41712,N_41713,N_41714,N_41715,N_41716,N_41717,N_41718,N_41719,N_41720,N_41721,N_41722,N_41723,N_41724,N_41725,N_41726,N_41727,N_41728,N_41729,N_41730,N_41731,N_41732,N_41733,N_41734,N_41735,N_41736,N_41737,N_41738,N_41739,N_41740,N_41741,N_41742,N_41743,N_41744,N_41745,N_41746,N_41747,N_41748,N_41749,N_41750,N_41751,N_41752,N_41753,N_41754,N_41755,N_41756,N_41757,N_41758,N_41759,N_41760,N_41761,N_41762,N_41763,N_41764,N_41765,N_41766,N_41767,N_41768,N_41769,N_41770,N_41771,N_41772,N_41773,N_41774,N_41775,N_41776,N_41777,N_41778,N_41779,N_41780,N_41781,N_41782,N_41783,N_41784,N_41785,N_41786,N_41787,N_41788,N_41789,N_41790,N_41791,N_41792,N_41793,N_41794,N_41795,N_41796,N_41797,N_41798,N_41799,N_41800,N_41801,N_41802,N_41803,N_41804,N_41805,N_41806,N_41807,N_41808,N_41809,N_41810,N_41811,N_41812,N_41813,N_41814,N_41815,N_41816,N_41817,N_41818,N_41819,N_41820,N_41821,N_41822,N_41823,N_41824,N_41825,N_41826,N_41827,N_41828,N_41829,N_41830,N_41831,N_41832,N_41833,N_41834,N_41835,N_41836,N_41837,N_41838,N_41839,N_41840,N_41841,N_41842,N_41843,N_41844,N_41845,N_41846,N_41847,N_41848,N_41849,N_41850,N_41851,N_41852,N_41853,N_41854,N_41855,N_41856,N_41857,N_41858,N_41859,N_41860,N_41861,N_41862,N_41863,N_41864,N_41865,N_41866,N_41867,N_41868,N_41869,N_41870,N_41871,N_41872,N_41873,N_41874,N_41875,N_41876,N_41877,N_41878,N_41879,N_41880,N_41881,N_41882,N_41883,N_41884,N_41885,N_41886,N_41887,N_41888,N_41889,N_41890,N_41891,N_41892,N_41893,N_41894,N_41895,N_41896,N_41897,N_41898,N_41899,N_41900,N_41901,N_41902,N_41903,N_41904,N_41905,N_41906,N_41907,N_41908,N_41909,N_41910,N_41911,N_41912,N_41913,N_41914,N_41915,N_41916,N_41917,N_41918,N_41919,N_41920,N_41921,N_41922,N_41923,N_41924,N_41925,N_41926,N_41927,N_41928,N_41929,N_41930,N_41931,N_41932,N_41933,N_41934,N_41935,N_41936,N_41937,N_41938,N_41939,N_41940,N_41941,N_41942,N_41943,N_41944,N_41945,N_41946,N_41947,N_41948,N_41949,N_41950,N_41951,N_41952,N_41953,N_41954,N_41955,N_41956,N_41957,N_41958,N_41959,N_41960,N_41961,N_41962,N_41963,N_41964,N_41965,N_41966,N_41967,N_41968,N_41969,N_41970,N_41971,N_41972,N_41973,N_41974,N_41975,N_41976,N_41977,N_41978,N_41979,N_41980,N_41981,N_41982,N_41983,N_41984,N_41985,N_41986,N_41987,N_41988,N_41989,N_41990,N_41991,N_41992,N_41993,N_41994,N_41995,N_41996,N_41997,N_41998,N_41999,N_42000,N_42001,N_42002,N_42003,N_42004,N_42005,N_42006,N_42007,N_42008,N_42009,N_42010,N_42011,N_42012,N_42013,N_42014,N_42015,N_42016,N_42017,N_42018,N_42019,N_42020,N_42021,N_42022,N_42023,N_42024,N_42025,N_42026,N_42027,N_42028,N_42029,N_42030,N_42031,N_42032,N_42033,N_42034,N_42035,N_42036,N_42037,N_42038,N_42039,N_42040,N_42041,N_42042,N_42043,N_42044,N_42045,N_42046,N_42047,N_42048,N_42049,N_42050,N_42051,N_42052,N_42053,N_42054,N_42055,N_42056,N_42057,N_42058,N_42059,N_42060,N_42061,N_42062,N_42063,N_42064,N_42065,N_42066,N_42067,N_42068,N_42069,N_42070,N_42071,N_42072,N_42073,N_42074,N_42075,N_42076,N_42077,N_42078,N_42079,N_42080,N_42081,N_42082,N_42083,N_42084,N_42085,N_42086,N_42087,N_42088,N_42089,N_42090,N_42091,N_42092,N_42093,N_42094,N_42095,N_42096,N_42097,N_42098,N_42099,N_42100,N_42101,N_42102,N_42103,N_42104,N_42105,N_42106,N_42107,N_42108,N_42109,N_42110,N_42111,N_42112,N_42113,N_42114,N_42115,N_42116,N_42117,N_42118,N_42119,N_42120,N_42121,N_42122,N_42123,N_42124,N_42125,N_42126,N_42127,N_42128,N_42129,N_42130,N_42131,N_42132,N_42133,N_42134,N_42135,N_42136,N_42137,N_42138,N_42139,N_42140,N_42141,N_42142,N_42143,N_42144,N_42145,N_42146,N_42147,N_42148,N_42149,N_42150,N_42151,N_42152,N_42153,N_42154,N_42155,N_42156,N_42157,N_42158,N_42159,N_42160,N_42161,N_42162,N_42163,N_42164,N_42165,N_42166,N_42167,N_42168,N_42169,N_42170,N_42171,N_42172,N_42173,N_42174,N_42175,N_42176,N_42177,N_42178,N_42179,N_42180,N_42181,N_42182,N_42183,N_42184,N_42185,N_42186,N_42187,N_42188,N_42189,N_42190,N_42191,N_42192,N_42193,N_42194,N_42195,N_42196,N_42197,N_42198,N_42199,N_42200,N_42201,N_42202,N_42203,N_42204,N_42205,N_42206,N_42207,N_42208,N_42209,N_42210,N_42211,N_42212,N_42213,N_42214,N_42215,N_42216,N_42217,N_42218,N_42219,N_42220,N_42221,N_42222,N_42223,N_42224,N_42225,N_42226,N_42227,N_42228,N_42229,N_42230,N_42231,N_42232,N_42233,N_42234,N_42235,N_42236,N_42237,N_42238,N_42239,N_42240,N_42241,N_42242,N_42243,N_42244,N_42245,N_42246,N_42247,N_42248,N_42249,N_42250,N_42251,N_42252,N_42253,N_42254,N_42255,N_42256,N_42257,N_42258,N_42259,N_42260,N_42261,N_42262,N_42263,N_42264,N_42265,N_42266,N_42267,N_42268,N_42269,N_42270,N_42271,N_42272,N_42273,N_42274,N_42275,N_42276,N_42277,N_42278,N_42279,N_42280,N_42281,N_42282,N_42283,N_42284,N_42285,N_42286,N_42287,N_42288,N_42289,N_42290,N_42291,N_42292,N_42293,N_42294,N_42295,N_42296,N_42297,N_42298,N_42299,N_42300,N_42301,N_42302,N_42303,N_42304,N_42305,N_42306,N_42307,N_42308,N_42309,N_42310,N_42311,N_42312,N_42313,N_42314,N_42315,N_42316,N_42317,N_42318,N_42319,N_42320,N_42321,N_42322,N_42323,N_42324,N_42325,N_42326,N_42327,N_42328,N_42329,N_42330,N_42331,N_42332,N_42333,N_42334,N_42335,N_42336,N_42337,N_42338,N_42339,N_42340,N_42341,N_42342,N_42343,N_42344,N_42345,N_42346,N_42347,N_42348,N_42349,N_42350,N_42351,N_42352,N_42353,N_42354,N_42355,N_42356,N_42357,N_42358,N_42359,N_42360,N_42361,N_42362,N_42363,N_42364,N_42365,N_42366,N_42367,N_42368,N_42369,N_42370,N_42371,N_42372,N_42373,N_42374,N_42375,N_42376,N_42377,N_42378,N_42379,N_42380,N_42381,N_42382,N_42383,N_42384,N_42385,N_42386,N_42387,N_42388,N_42389,N_42390,N_42391,N_42392,N_42393,N_42394,N_42395,N_42396,N_42397,N_42398,N_42399,N_42400,N_42401,N_42402,N_42403,N_42404,N_42405,N_42406,N_42407,N_42408,N_42409,N_42410,N_42411,N_42412,N_42413,N_42414,N_42415,N_42416,N_42417,N_42418,N_42419,N_42420,N_42421,N_42422,N_42423,N_42424,N_42425,N_42426,N_42427,N_42428,N_42429,N_42430,N_42431,N_42432,N_42433,N_42434,N_42435,N_42436,N_42437,N_42438,N_42439,N_42440,N_42441,N_42442,N_42443,N_42444,N_42445,N_42446,N_42447,N_42448,N_42449,N_42450,N_42451,N_42452,N_42453,N_42454,N_42455,N_42456,N_42457,N_42458,N_42459,N_42460,N_42461,N_42462,N_42463,N_42464,N_42465,N_42466,N_42467,N_42468,N_42469,N_42470,N_42471,N_42472,N_42473,N_42474,N_42475,N_42476,N_42477,N_42478,N_42479,N_42480,N_42481,N_42482,N_42483,N_42484,N_42485,N_42486,N_42487,N_42488,N_42489,N_42490,N_42491,N_42492,N_42493,N_42494,N_42495,N_42496,N_42497,N_42498,N_42499,N_42500,N_42501,N_42502,N_42503,N_42504,N_42505,N_42506,N_42507,N_42508,N_42509,N_42510,N_42511,N_42512,N_42513,N_42514,N_42515,N_42516,N_42517,N_42518,N_42519,N_42520,N_42521,N_42522,N_42523,N_42524,N_42525,N_42526,N_42527,N_42528,N_42529,N_42530,N_42531,N_42532,N_42533,N_42534,N_42535,N_42536,N_42537,N_42538,N_42539,N_42540,N_42541,N_42542,N_42543,N_42544,N_42545,N_42546,N_42547,N_42548,N_42549,N_42550,N_42551,N_42552,N_42553,N_42554,N_42555,N_42556,N_42557,N_42558,N_42559,N_42560,N_42561,N_42562,N_42563,N_42564,N_42565,N_42566,N_42567,N_42568,N_42569,N_42570,N_42571,N_42572,N_42573,N_42574,N_42575,N_42576,N_42577,N_42578,N_42579,N_42580,N_42581,N_42582,N_42583,N_42584,N_42585,N_42586,N_42587,N_42588,N_42589,N_42590,N_42591,N_42592,N_42593,N_42594,N_42595,N_42596,N_42597,N_42598,N_42599,N_42600,N_42601,N_42602,N_42603,N_42604,N_42605,N_42606,N_42607,N_42608,N_42609,N_42610,N_42611,N_42612,N_42613,N_42614,N_42615,N_42616,N_42617,N_42618,N_42619,N_42620,N_42621,N_42622,N_42623,N_42624,N_42625,N_42626,N_42627,N_42628,N_42629,N_42630,N_42631,N_42632,N_42633,N_42634,N_42635,N_42636,N_42637,N_42638,N_42639,N_42640,N_42641,N_42642,N_42643,N_42644,N_42645,N_42646,N_42647,N_42648,N_42649,N_42650,N_42651,N_42652,N_42653,N_42654,N_42655,N_42656,N_42657,N_42658,N_42659,N_42660,N_42661,N_42662,N_42663,N_42664,N_42665,N_42666,N_42667,N_42668,N_42669,N_42670,N_42671,N_42672,N_42673,N_42674,N_42675,N_42676,N_42677,N_42678,N_42679,N_42680,N_42681,N_42682,N_42683,N_42684,N_42685,N_42686,N_42687,N_42688,N_42689,N_42690,N_42691,N_42692,N_42693,N_42694,N_42695,N_42696,N_42697,N_42698,N_42699,N_42700,N_42701,N_42702,N_42703,N_42704,N_42705,N_42706,N_42707,N_42708,N_42709,N_42710,N_42711,N_42712,N_42713,N_42714,N_42715,N_42716,N_42717,N_42718,N_42719,N_42720,N_42721,N_42722,N_42723,N_42724,N_42725,N_42726,N_42727,N_42728,N_42729,N_42730,N_42731,N_42732,N_42733,N_42734,N_42735,N_42736,N_42737,N_42738,N_42739,N_42740,N_42741,N_42742,N_42743,N_42744,N_42745,N_42746,N_42747,N_42748,N_42749,N_42750,N_42751,N_42752,N_42753,N_42754,N_42755,N_42756,N_42757,N_42758,N_42759,N_42760,N_42761,N_42762,N_42763,N_42764,N_42765,N_42766,N_42767,N_42768,N_42769,N_42770,N_42771,N_42772,N_42773,N_42774,N_42775,N_42776,N_42777,N_42778,N_42779,N_42780,N_42781,N_42782,N_42783,N_42784,N_42785,N_42786,N_42787,N_42788,N_42789,N_42790,N_42791,N_42792,N_42793,N_42794,N_42795,N_42796,N_42797,N_42798,N_42799,N_42800,N_42801,N_42802,N_42803,N_42804,N_42805,N_42806,N_42807,N_42808,N_42809,N_42810,N_42811,N_42812,N_42813,N_42814,N_42815,N_42816,N_42817,N_42818,N_42819,N_42820,N_42821,N_42822,N_42823,N_42824,N_42825,N_42826,N_42827,N_42828,N_42829,N_42830,N_42831,N_42832,N_42833,N_42834,N_42835,N_42836,N_42837,N_42838,N_42839,N_42840,N_42841,N_42842,N_42843,N_42844,N_42845,N_42846,N_42847,N_42848,N_42849,N_42850,N_42851,N_42852,N_42853,N_42854,N_42855,N_42856,N_42857,N_42858,N_42859,N_42860,N_42861,N_42862,N_42863,N_42864,N_42865,N_42866,N_42867,N_42868,N_42869,N_42870,N_42871,N_42872,N_42873,N_42874,N_42875,N_42876,N_42877,N_42878,N_42879,N_42880,N_42881,N_42882,N_42883,N_42884,N_42885,N_42886,N_42887,N_42888,N_42889,N_42890,N_42891,N_42892,N_42893,N_42894,N_42895,N_42896,N_42897,N_42898,N_42899,N_42900,N_42901,N_42902,N_42903,N_42904,N_42905,N_42906,N_42907,N_42908,N_42909,N_42910,N_42911,N_42912,N_42913,N_42914,N_42915,N_42916,N_42917,N_42918,N_42919,N_42920,N_42921,N_42922,N_42923,N_42924,N_42925,N_42926,N_42927,N_42928,N_42929,N_42930,N_42931,N_42932,N_42933,N_42934,N_42935,N_42936,N_42937,N_42938,N_42939,N_42940,N_42941,N_42942,N_42943,N_42944,N_42945,N_42946,N_42947,N_42948,N_42949,N_42950,N_42951,N_42952,N_42953,N_42954,N_42955,N_42956,N_42957,N_42958,N_42959,N_42960,N_42961,N_42962,N_42963,N_42964,N_42965,N_42966,N_42967,N_42968,N_42969,N_42970,N_42971,N_42972,N_42973,N_42974,N_42975,N_42976,N_42977,N_42978,N_42979,N_42980,N_42981,N_42982,N_42983,N_42984,N_42985,N_42986,N_42987,N_42988,N_42989,N_42990,N_42991,N_42992,N_42993,N_42994,N_42995,N_42996,N_42997,N_42998,N_42999,N_43000,N_43001,N_43002,N_43003,N_43004,N_43005,N_43006,N_43007,N_43008,N_43009,N_43010,N_43011,N_43012,N_43013,N_43014,N_43015,N_43016,N_43017,N_43018,N_43019,N_43020,N_43021,N_43022,N_43023,N_43024,N_43025,N_43026,N_43027,N_43028,N_43029,N_43030,N_43031,N_43032,N_43033,N_43034,N_43035,N_43036,N_43037,N_43038,N_43039,N_43040,N_43041,N_43042,N_43043,N_43044,N_43045,N_43046,N_43047,N_43048,N_43049,N_43050,N_43051,N_43052,N_43053,N_43054,N_43055,N_43056,N_43057,N_43058,N_43059,N_43060,N_43061,N_43062,N_43063,N_43064,N_43065,N_43066,N_43067,N_43068,N_43069,N_43070,N_43071,N_43072,N_43073,N_43074,N_43075,N_43076,N_43077,N_43078,N_43079,N_43080,N_43081,N_43082,N_43083,N_43084,N_43085,N_43086,N_43087,N_43088,N_43089,N_43090,N_43091,N_43092,N_43093,N_43094,N_43095,N_43096,N_43097,N_43098,N_43099,N_43100,N_43101,N_43102,N_43103,N_43104,N_43105,N_43106,N_43107,N_43108,N_43109,N_43110,N_43111,N_43112,N_43113,N_43114,N_43115,N_43116,N_43117,N_43118,N_43119,N_43120,N_43121,N_43122,N_43123,N_43124,N_43125,N_43126,N_43127,N_43128,N_43129,N_43130,N_43131,N_43132,N_43133,N_43134,N_43135,N_43136,N_43137,N_43138,N_43139,N_43140,N_43141,N_43142,N_43143,N_43144,N_43145,N_43146,N_43147,N_43148,N_43149,N_43150,N_43151,N_43152,N_43153,N_43154,N_43155,N_43156,N_43157,N_43158,N_43159,N_43160,N_43161,N_43162,N_43163,N_43164,N_43165,N_43166,N_43167,N_43168,N_43169,N_43170,N_43171,N_43172,N_43173,N_43174,N_43175,N_43176,N_43177,N_43178,N_43179,N_43180,N_43181,N_43182,N_43183,N_43184,N_43185,N_43186,N_43187,N_43188,N_43189,N_43190,N_43191,N_43192,N_43193,N_43194,N_43195,N_43196,N_43197,N_43198,N_43199,N_43200,N_43201,N_43202,N_43203,N_43204,N_43205,N_43206,N_43207,N_43208,N_43209,N_43210,N_43211,N_43212,N_43213,N_43214,N_43215,N_43216,N_43217,N_43218,N_43219,N_43220,N_43221,N_43222,N_43223,N_43224,N_43225,N_43226,N_43227,N_43228,N_43229,N_43230,N_43231,N_43232,N_43233,N_43234,N_43235,N_43236,N_43237,N_43238,N_43239,N_43240,N_43241,N_43242,N_43243,N_43244,N_43245,N_43246,N_43247,N_43248,N_43249,N_43250,N_43251,N_43252,N_43253,N_43254,N_43255,N_43256,N_43257,N_43258,N_43259,N_43260,N_43261,N_43262,N_43263,N_43264,N_43265,N_43266,N_43267,N_43268,N_43269,N_43270,N_43271,N_43272,N_43273,N_43274,N_43275,N_43276,N_43277,N_43278,N_43279,N_43280,N_43281,N_43282,N_43283,N_43284,N_43285,N_43286,N_43287,N_43288,N_43289,N_43290,N_43291,N_43292,N_43293,N_43294,N_43295,N_43296,N_43297,N_43298,N_43299,N_43300,N_43301,N_43302,N_43303,N_43304,N_43305,N_43306,N_43307,N_43308,N_43309,N_43310,N_43311,N_43312,N_43313,N_43314,N_43315,N_43316,N_43317,N_43318,N_43319,N_43320,N_43321,N_43322,N_43323,N_43324,N_43325,N_43326,N_43327,N_43328,N_43329,N_43330,N_43331,N_43332,N_43333,N_43334,N_43335,N_43336,N_43337,N_43338,N_43339,N_43340,N_43341,N_43342,N_43343,N_43344,N_43345,N_43346,N_43347,N_43348,N_43349,N_43350,N_43351,N_43352,N_43353,N_43354,N_43355,N_43356,N_43357,N_43358,N_43359,N_43360,N_43361,N_43362,N_43363,N_43364,N_43365,N_43366,N_43367,N_43368,N_43369,N_43370,N_43371,N_43372,N_43373,N_43374,N_43375,N_43376,N_43377,N_43378,N_43379,N_43380,N_43381,N_43382,N_43383,N_43384,N_43385,N_43386,N_43387,N_43388,N_43389,N_43390,N_43391,N_43392,N_43393,N_43394,N_43395,N_43396,N_43397,N_43398,N_43399,N_43400,N_43401,N_43402,N_43403,N_43404,N_43405,N_43406,N_43407,N_43408,N_43409,N_43410,N_43411,N_43412,N_43413,N_43414,N_43415,N_43416,N_43417,N_43418,N_43419,N_43420,N_43421,N_43422,N_43423,N_43424,N_43425,N_43426,N_43427,N_43428,N_43429,N_43430,N_43431,N_43432,N_43433,N_43434,N_43435,N_43436,N_43437,N_43438,N_43439,N_43440,N_43441,N_43442,N_43443,N_43444,N_43445,N_43446,N_43447,N_43448,N_43449,N_43450,N_43451,N_43452,N_43453,N_43454,N_43455,N_43456,N_43457,N_43458,N_43459,N_43460,N_43461,N_43462,N_43463,N_43464,N_43465,N_43466,N_43467,N_43468,N_43469,N_43470,N_43471,N_43472,N_43473,N_43474,N_43475,N_43476,N_43477,N_43478,N_43479,N_43480,N_43481,N_43482,N_43483,N_43484,N_43485,N_43486,N_43487,N_43488,N_43489,N_43490,N_43491,N_43492,N_43493,N_43494,N_43495,N_43496,N_43497,N_43498,N_43499,N_43500,N_43501,N_43502,N_43503,N_43504,N_43505,N_43506,N_43507,N_43508,N_43509,N_43510,N_43511,N_43512,N_43513,N_43514,N_43515,N_43516,N_43517,N_43518,N_43519,N_43520,N_43521,N_43522,N_43523,N_43524,N_43525,N_43526,N_43527,N_43528,N_43529,N_43530,N_43531,N_43532,N_43533,N_43534,N_43535,N_43536,N_43537,N_43538,N_43539,N_43540,N_43541,N_43542,N_43543,N_43544,N_43545,N_43546,N_43547,N_43548,N_43549,N_43550,N_43551,N_43552,N_43553,N_43554,N_43555,N_43556,N_43557,N_43558,N_43559,N_43560,N_43561,N_43562,N_43563,N_43564,N_43565,N_43566,N_43567,N_43568,N_43569,N_43570,N_43571,N_43572,N_43573,N_43574,N_43575,N_43576,N_43577,N_43578,N_43579,N_43580,N_43581,N_43582,N_43583,N_43584,N_43585,N_43586,N_43587,N_43588,N_43589,N_43590,N_43591,N_43592,N_43593,N_43594,N_43595,N_43596,N_43597,N_43598,N_43599,N_43600,N_43601,N_43602,N_43603,N_43604,N_43605,N_43606,N_43607,N_43608,N_43609,N_43610,N_43611,N_43612,N_43613,N_43614,N_43615,N_43616,N_43617,N_43618,N_43619,N_43620,N_43621,N_43622,N_43623,N_43624,N_43625,N_43626,N_43627,N_43628,N_43629,N_43630,N_43631,N_43632,N_43633,N_43634,N_43635,N_43636,N_43637,N_43638,N_43639,N_43640,N_43641,N_43642,N_43643,N_43644,N_43645,N_43646,N_43647,N_43648,N_43649,N_43650,N_43651,N_43652,N_43653,N_43654,N_43655,N_43656,N_43657,N_43658,N_43659,N_43660,N_43661,N_43662,N_43663,N_43664,N_43665,N_43666,N_43667,N_43668,N_43669,N_43670,N_43671,N_43672,N_43673,N_43674,N_43675,N_43676,N_43677,N_43678,N_43679,N_43680,N_43681,N_43682,N_43683,N_43684,N_43685,N_43686,N_43687,N_43688,N_43689,N_43690,N_43691,N_43692,N_43693,N_43694,N_43695,N_43696,N_43697,N_43698,N_43699,N_43700,N_43701,N_43702,N_43703,N_43704,N_43705,N_43706,N_43707,N_43708,N_43709,N_43710,N_43711,N_43712,N_43713,N_43714,N_43715,N_43716,N_43717,N_43718,N_43719,N_43720,N_43721,N_43722,N_43723,N_43724,N_43725,N_43726,N_43727,N_43728,N_43729,N_43730,N_43731,N_43732,N_43733,N_43734,N_43735,N_43736,N_43737,N_43738,N_43739,N_43740,N_43741,N_43742,N_43743,N_43744,N_43745,N_43746,N_43747,N_43748,N_43749,N_43750,N_43751,N_43752,N_43753,N_43754,N_43755,N_43756,N_43757,N_43758,N_43759,N_43760,N_43761,N_43762,N_43763,N_43764,N_43765,N_43766,N_43767,N_43768,N_43769,N_43770,N_43771,N_43772,N_43773,N_43774,N_43775,N_43776,N_43777,N_43778,N_43779,N_43780,N_43781,N_43782,N_43783,N_43784,N_43785,N_43786,N_43787,N_43788,N_43789,N_43790,N_43791,N_43792,N_43793,N_43794,N_43795,N_43796,N_43797,N_43798,N_43799,N_43800,N_43801,N_43802,N_43803,N_43804,N_43805,N_43806,N_43807,N_43808,N_43809,N_43810,N_43811,N_43812,N_43813,N_43814,N_43815,N_43816,N_43817,N_43818,N_43819,N_43820,N_43821,N_43822,N_43823,N_43824,N_43825,N_43826,N_43827,N_43828,N_43829,N_43830,N_43831,N_43832,N_43833,N_43834,N_43835,N_43836,N_43837,N_43838,N_43839,N_43840,N_43841,N_43842,N_43843,N_43844,N_43845,N_43846,N_43847,N_43848,N_43849,N_43850,N_43851,N_43852,N_43853,N_43854,N_43855,N_43856,N_43857,N_43858,N_43859,N_43860,N_43861,N_43862,N_43863,N_43864,N_43865,N_43866,N_43867,N_43868,N_43869,N_43870,N_43871,N_43872,N_43873,N_43874,N_43875,N_43876,N_43877,N_43878,N_43879,N_43880,N_43881,N_43882,N_43883,N_43884,N_43885,N_43886,N_43887,N_43888,N_43889,N_43890,N_43891,N_43892,N_43893,N_43894,N_43895,N_43896,N_43897,N_43898,N_43899,N_43900,N_43901,N_43902,N_43903,N_43904,N_43905,N_43906,N_43907,N_43908,N_43909,N_43910,N_43911,N_43912,N_43913,N_43914,N_43915,N_43916,N_43917,N_43918,N_43919,N_43920,N_43921,N_43922,N_43923,N_43924,N_43925,N_43926,N_43927,N_43928,N_43929,N_43930,N_43931,N_43932,N_43933,N_43934,N_43935,N_43936,N_43937,N_43938,N_43939,N_43940,N_43941,N_43942,N_43943,N_43944,N_43945,N_43946,N_43947,N_43948,N_43949,N_43950,N_43951,N_43952,N_43953,N_43954,N_43955,N_43956,N_43957,N_43958,N_43959,N_43960,N_43961,N_43962,N_43963,N_43964,N_43965,N_43966,N_43967,N_43968,N_43969,N_43970,N_43971,N_43972,N_43973,N_43974,N_43975,N_43976,N_43977,N_43978,N_43979,N_43980,N_43981,N_43982,N_43983,N_43984,N_43985,N_43986,N_43987,N_43988,N_43989,N_43990,N_43991,N_43992,N_43993,N_43994,N_43995,N_43996,N_43997,N_43998,N_43999,N_44000,N_44001,N_44002,N_44003,N_44004,N_44005,N_44006,N_44007,N_44008,N_44009,N_44010,N_44011,N_44012,N_44013,N_44014,N_44015,N_44016,N_44017,N_44018,N_44019,N_44020,N_44021,N_44022,N_44023,N_44024,N_44025,N_44026,N_44027,N_44028,N_44029,N_44030,N_44031,N_44032,N_44033,N_44034,N_44035,N_44036,N_44037,N_44038,N_44039,N_44040,N_44041,N_44042,N_44043,N_44044,N_44045,N_44046,N_44047,N_44048,N_44049,N_44050,N_44051,N_44052,N_44053,N_44054,N_44055,N_44056,N_44057,N_44058,N_44059,N_44060,N_44061,N_44062,N_44063,N_44064,N_44065,N_44066,N_44067,N_44068,N_44069,N_44070,N_44071,N_44072,N_44073,N_44074,N_44075,N_44076,N_44077,N_44078,N_44079,N_44080,N_44081,N_44082,N_44083,N_44084,N_44085,N_44086,N_44087,N_44088,N_44089,N_44090,N_44091,N_44092,N_44093,N_44094,N_44095,N_44096,N_44097,N_44098,N_44099,N_44100,N_44101,N_44102,N_44103,N_44104,N_44105,N_44106,N_44107,N_44108,N_44109,N_44110,N_44111,N_44112,N_44113,N_44114,N_44115,N_44116,N_44117,N_44118,N_44119,N_44120,N_44121,N_44122,N_44123,N_44124,N_44125,N_44126,N_44127,N_44128,N_44129,N_44130,N_44131,N_44132,N_44133,N_44134,N_44135,N_44136,N_44137,N_44138,N_44139,N_44140,N_44141,N_44142,N_44143,N_44144,N_44145,N_44146,N_44147,N_44148,N_44149,N_44150,N_44151,N_44152,N_44153,N_44154,N_44155,N_44156,N_44157,N_44158,N_44159,N_44160,N_44161,N_44162,N_44163,N_44164,N_44165,N_44166,N_44167,N_44168,N_44169,N_44170,N_44171,N_44172,N_44173,N_44174,N_44175,N_44176,N_44177,N_44178,N_44179,N_44180,N_44181,N_44182,N_44183,N_44184,N_44185,N_44186,N_44187,N_44188,N_44189,N_44190,N_44191,N_44192,N_44193,N_44194,N_44195,N_44196,N_44197,N_44198,N_44199,N_44200,N_44201,N_44202,N_44203,N_44204,N_44205,N_44206,N_44207,N_44208,N_44209,N_44210,N_44211,N_44212,N_44213,N_44214,N_44215,N_44216,N_44217,N_44218,N_44219,N_44220,N_44221,N_44222,N_44223,N_44224,N_44225,N_44226,N_44227,N_44228,N_44229,N_44230,N_44231,N_44232,N_44233,N_44234,N_44235,N_44236,N_44237,N_44238,N_44239,N_44240,N_44241,N_44242,N_44243,N_44244,N_44245,N_44246,N_44247,N_44248,N_44249,N_44250,N_44251,N_44252,N_44253,N_44254,N_44255,N_44256,N_44257,N_44258,N_44259,N_44260,N_44261,N_44262,N_44263,N_44264,N_44265,N_44266,N_44267,N_44268,N_44269,N_44270,N_44271,N_44272,N_44273,N_44274,N_44275,N_44276,N_44277,N_44278,N_44279,N_44280,N_44281,N_44282,N_44283,N_44284,N_44285,N_44286,N_44287,N_44288,N_44289,N_44290,N_44291,N_44292,N_44293,N_44294,N_44295,N_44296,N_44297,N_44298,N_44299,N_44300,N_44301,N_44302,N_44303,N_44304,N_44305,N_44306,N_44307,N_44308,N_44309,N_44310,N_44311,N_44312,N_44313,N_44314,N_44315,N_44316,N_44317,N_44318,N_44319,N_44320,N_44321,N_44322,N_44323,N_44324,N_44325,N_44326,N_44327,N_44328,N_44329,N_44330,N_44331,N_44332,N_44333,N_44334,N_44335,N_44336,N_44337,N_44338,N_44339,N_44340,N_44341,N_44342,N_44343,N_44344,N_44345,N_44346,N_44347,N_44348,N_44349,N_44350,N_44351,N_44352,N_44353,N_44354,N_44355,N_44356,N_44357,N_44358,N_44359,N_44360,N_44361,N_44362,N_44363,N_44364,N_44365,N_44366,N_44367,N_44368,N_44369,N_44370,N_44371,N_44372,N_44373,N_44374,N_44375,N_44376,N_44377,N_44378,N_44379,N_44380,N_44381,N_44382,N_44383,N_44384,N_44385,N_44386,N_44387,N_44388,N_44389,N_44390,N_44391,N_44392,N_44393,N_44394,N_44395,N_44396,N_44397,N_44398,N_44399,N_44400,N_44401,N_44402,N_44403,N_44404,N_44405,N_44406,N_44407,N_44408,N_44409,N_44410,N_44411,N_44412,N_44413,N_44414,N_44415,N_44416,N_44417,N_44418,N_44419,N_44420,N_44421,N_44422,N_44423,N_44424,N_44425,N_44426,N_44427,N_44428,N_44429,N_44430,N_44431,N_44432,N_44433,N_44434,N_44435,N_44436,N_44437,N_44438,N_44439,N_44440,N_44441,N_44442,N_44443,N_44444,N_44445,N_44446,N_44447,N_44448,N_44449,N_44450,N_44451,N_44452,N_44453,N_44454,N_44455,N_44456,N_44457,N_44458,N_44459,N_44460,N_44461,N_44462,N_44463,N_44464,N_44465,N_44466,N_44467,N_44468,N_44469,N_44470,N_44471,N_44472,N_44473,N_44474,N_44475,N_44476,N_44477,N_44478,N_44479,N_44480,N_44481,N_44482,N_44483,N_44484,N_44485,N_44486,N_44487,N_44488,N_44489,N_44490,N_44491,N_44492,N_44493,N_44494,N_44495,N_44496,N_44497,N_44498,N_44499,N_44500,N_44501,N_44502,N_44503,N_44504,N_44505,N_44506,N_44507,N_44508,N_44509,N_44510,N_44511,N_44512,N_44513,N_44514,N_44515,N_44516,N_44517,N_44518,N_44519,N_44520,N_44521,N_44522,N_44523,N_44524,N_44525,N_44526,N_44527,N_44528,N_44529,N_44530,N_44531,N_44532,N_44533,N_44534,N_44535,N_44536,N_44537,N_44538,N_44539,N_44540,N_44541,N_44542,N_44543,N_44544,N_44545,N_44546,N_44547,N_44548,N_44549,N_44550,N_44551,N_44552,N_44553,N_44554,N_44555,N_44556,N_44557,N_44558,N_44559,N_44560,N_44561,N_44562,N_44563,N_44564,N_44565,N_44566,N_44567,N_44568,N_44569,N_44570,N_44571,N_44572,N_44573,N_44574,N_44575,N_44576,N_44577,N_44578,N_44579,N_44580,N_44581,N_44582,N_44583,N_44584,N_44585,N_44586,N_44587,N_44588,N_44589,N_44590,N_44591,N_44592,N_44593,N_44594,N_44595,N_44596,N_44597,N_44598,N_44599,N_44600,N_44601,N_44602,N_44603,N_44604,N_44605,N_44606,N_44607,N_44608,N_44609,N_44610,N_44611,N_44612,N_44613,N_44614,N_44615,N_44616,N_44617,N_44618,N_44619,N_44620,N_44621,N_44622,N_44623,N_44624,N_44625,N_44626,N_44627,N_44628,N_44629,N_44630,N_44631,N_44632,N_44633,N_44634,N_44635,N_44636,N_44637,N_44638,N_44639,N_44640,N_44641,N_44642,N_44643,N_44644,N_44645,N_44646,N_44647,N_44648,N_44649,N_44650,N_44651,N_44652,N_44653,N_44654,N_44655,N_44656,N_44657,N_44658,N_44659,N_44660,N_44661,N_44662,N_44663,N_44664,N_44665,N_44666,N_44667,N_44668,N_44669,N_44670,N_44671,N_44672,N_44673,N_44674,N_44675,N_44676,N_44677,N_44678,N_44679,N_44680,N_44681,N_44682,N_44683,N_44684,N_44685,N_44686,N_44687,N_44688,N_44689,N_44690,N_44691,N_44692,N_44693,N_44694,N_44695,N_44696,N_44697,N_44698,N_44699,N_44700,N_44701,N_44702,N_44703,N_44704,N_44705,N_44706,N_44707,N_44708,N_44709,N_44710,N_44711,N_44712,N_44713,N_44714,N_44715,N_44716,N_44717,N_44718,N_44719,N_44720,N_44721,N_44722,N_44723,N_44724,N_44725,N_44726,N_44727,N_44728,N_44729,N_44730,N_44731,N_44732,N_44733,N_44734,N_44735,N_44736,N_44737,N_44738,N_44739,N_44740,N_44741,N_44742,N_44743,N_44744,N_44745,N_44746,N_44747,N_44748,N_44749,N_44750,N_44751,N_44752,N_44753,N_44754,N_44755,N_44756,N_44757,N_44758,N_44759,N_44760,N_44761,N_44762,N_44763,N_44764,N_44765,N_44766,N_44767,N_44768,N_44769,N_44770,N_44771,N_44772,N_44773,N_44774,N_44775,N_44776,N_44777,N_44778,N_44779,N_44780,N_44781,N_44782,N_44783,N_44784,N_44785,N_44786,N_44787,N_44788,N_44789,N_44790,N_44791,N_44792,N_44793,N_44794,N_44795,N_44796,N_44797,N_44798,N_44799,N_44800,N_44801,N_44802,N_44803,N_44804,N_44805,N_44806,N_44807,N_44808,N_44809,N_44810,N_44811,N_44812,N_44813,N_44814,N_44815,N_44816,N_44817,N_44818,N_44819,N_44820,N_44821,N_44822,N_44823,N_44824,N_44825,N_44826,N_44827,N_44828,N_44829,N_44830,N_44831,N_44832,N_44833,N_44834,N_44835,N_44836,N_44837,N_44838,N_44839,N_44840,N_44841,N_44842,N_44843,N_44844,N_44845,N_44846,N_44847,N_44848,N_44849,N_44850,N_44851,N_44852,N_44853,N_44854,N_44855,N_44856,N_44857,N_44858,N_44859,N_44860,N_44861,N_44862,N_44863,N_44864,N_44865,N_44866,N_44867,N_44868,N_44869,N_44870,N_44871,N_44872,N_44873,N_44874,N_44875,N_44876,N_44877,N_44878,N_44879,N_44880,N_44881,N_44882,N_44883,N_44884,N_44885,N_44886,N_44887,N_44888,N_44889,N_44890,N_44891,N_44892,N_44893,N_44894,N_44895,N_44896,N_44897,N_44898,N_44899,N_44900,N_44901,N_44902,N_44903,N_44904,N_44905,N_44906,N_44907,N_44908,N_44909,N_44910,N_44911,N_44912,N_44913,N_44914,N_44915,N_44916,N_44917,N_44918,N_44919,N_44920,N_44921,N_44922,N_44923,N_44924,N_44925,N_44926,N_44927,N_44928,N_44929,N_44930,N_44931,N_44932,N_44933,N_44934,N_44935,N_44936,N_44937,N_44938,N_44939,N_44940,N_44941,N_44942,N_44943,N_44944,N_44945,N_44946,N_44947,N_44948,N_44949,N_44950,N_44951,N_44952,N_44953,N_44954,N_44955,N_44956,N_44957,N_44958,N_44959,N_44960,N_44961,N_44962,N_44963,N_44964,N_44965,N_44966,N_44967,N_44968,N_44969,N_44970,N_44971,N_44972,N_44973,N_44974,N_44975,N_44976,N_44977,N_44978,N_44979,N_44980,N_44981,N_44982,N_44983,N_44984,N_44985,N_44986,N_44987,N_44988,N_44989,N_44990,N_44991,N_44992,N_44993,N_44994,N_44995,N_44996,N_44997,N_44998,N_44999,N_45000,N_45001,N_45002,N_45003,N_45004,N_45005,N_45006,N_45007,N_45008,N_45009,N_45010,N_45011,N_45012,N_45013,N_45014,N_45015,N_45016,N_45017,N_45018,N_45019,N_45020,N_45021,N_45022,N_45023,N_45024,N_45025,N_45026,N_45027,N_45028,N_45029,N_45030,N_45031,N_45032,N_45033,N_45034,N_45035,N_45036,N_45037,N_45038,N_45039,N_45040,N_45041,N_45042,N_45043,N_45044,N_45045,N_45046,N_45047,N_45048,N_45049,N_45050,N_45051,N_45052,N_45053,N_45054,N_45055,N_45056,N_45057,N_45058,N_45059,N_45060,N_45061,N_45062,N_45063,N_45064,N_45065,N_45066,N_45067,N_45068,N_45069,N_45070,N_45071,N_45072,N_45073,N_45074,N_45075,N_45076,N_45077,N_45078,N_45079,N_45080,N_45081,N_45082,N_45083,N_45084,N_45085,N_45086,N_45087,N_45088,N_45089,N_45090,N_45091,N_45092,N_45093,N_45094,N_45095,N_45096,N_45097,N_45098,N_45099,N_45100,N_45101,N_45102,N_45103,N_45104,N_45105,N_45106,N_45107,N_45108,N_45109,N_45110,N_45111,N_45112,N_45113,N_45114,N_45115,N_45116,N_45117,N_45118,N_45119,N_45120,N_45121,N_45122,N_45123,N_45124,N_45125,N_45126,N_45127,N_45128,N_45129,N_45130,N_45131,N_45132,N_45133,N_45134,N_45135,N_45136,N_45137,N_45138,N_45139,N_45140,N_45141,N_45142,N_45143,N_45144,N_45145,N_45146,N_45147,N_45148,N_45149,N_45150,N_45151,N_45152,N_45153,N_45154,N_45155,N_45156,N_45157,N_45158,N_45159,N_45160,N_45161,N_45162,N_45163,N_45164,N_45165,N_45166,N_45167,N_45168,N_45169,N_45170,N_45171,N_45172,N_45173,N_45174,N_45175,N_45176,N_45177,N_45178,N_45179,N_45180,N_45181,N_45182,N_45183,N_45184,N_45185,N_45186,N_45187,N_45188,N_45189,N_45190,N_45191,N_45192,N_45193,N_45194,N_45195,N_45196,N_45197,N_45198,N_45199,N_45200,N_45201,N_45202,N_45203,N_45204,N_45205,N_45206,N_45207,N_45208,N_45209,N_45210,N_45211,N_45212,N_45213,N_45214,N_45215,N_45216,N_45217,N_45218,N_45219,N_45220,N_45221,N_45222,N_45223,N_45224,N_45225,N_45226,N_45227,N_45228,N_45229,N_45230,N_45231,N_45232,N_45233,N_45234,N_45235,N_45236,N_45237,N_45238,N_45239,N_45240,N_45241,N_45242,N_45243,N_45244,N_45245,N_45246,N_45247,N_45248,N_45249,N_45250,N_45251,N_45252,N_45253,N_45254,N_45255,N_45256,N_45257,N_45258,N_45259,N_45260,N_45261,N_45262,N_45263,N_45264,N_45265,N_45266,N_45267,N_45268,N_45269,N_45270,N_45271,N_45272,N_45273,N_45274,N_45275,N_45276,N_45277,N_45278,N_45279,N_45280,N_45281,N_45282,N_45283,N_45284,N_45285,N_45286,N_45287,N_45288,N_45289,N_45290,N_45291,N_45292,N_45293,N_45294,N_45295,N_45296,N_45297,N_45298,N_45299,N_45300,N_45301,N_45302,N_45303,N_45304,N_45305,N_45306,N_45307,N_45308,N_45309,N_45310,N_45311,N_45312,N_45313,N_45314,N_45315,N_45316,N_45317,N_45318,N_45319,N_45320,N_45321,N_45322,N_45323,N_45324,N_45325,N_45326,N_45327,N_45328,N_45329,N_45330,N_45331,N_45332,N_45333,N_45334,N_45335,N_45336,N_45337,N_45338,N_45339,N_45340,N_45341,N_45342,N_45343,N_45344,N_45345,N_45346,N_45347,N_45348,N_45349,N_45350,N_45351,N_45352,N_45353,N_45354,N_45355,N_45356,N_45357,N_45358,N_45359,N_45360,N_45361,N_45362,N_45363,N_45364,N_45365,N_45366,N_45367,N_45368,N_45369,N_45370,N_45371,N_45372,N_45373,N_45374,N_45375,N_45376,N_45377,N_45378,N_45379,N_45380,N_45381,N_45382,N_45383,N_45384,N_45385,N_45386,N_45387,N_45388,N_45389,N_45390,N_45391,N_45392,N_45393,N_45394,N_45395,N_45396,N_45397,N_45398,N_45399,N_45400,N_45401,N_45402,N_45403,N_45404,N_45405,N_45406,N_45407,N_45408,N_45409,N_45410,N_45411,N_45412,N_45413,N_45414,N_45415,N_45416,N_45417,N_45418,N_45419,N_45420,N_45421,N_45422,N_45423,N_45424,N_45425,N_45426,N_45427,N_45428,N_45429,N_45430,N_45431,N_45432,N_45433,N_45434,N_45435,N_45436,N_45437,N_45438,N_45439,N_45440,N_45441,N_45442,N_45443,N_45444,N_45445,N_45446,N_45447,N_45448,N_45449,N_45450,N_45451,N_45452,N_45453,N_45454,N_45455,N_45456,N_45457,N_45458,N_45459,N_45460,N_45461,N_45462,N_45463,N_45464,N_45465,N_45466,N_45467,N_45468,N_45469,N_45470,N_45471,N_45472,N_45473,N_45474,N_45475,N_45476,N_45477,N_45478,N_45479,N_45480,N_45481,N_45482,N_45483,N_45484,N_45485,N_45486,N_45487,N_45488,N_45489,N_45490,N_45491,N_45492,N_45493,N_45494,N_45495,N_45496,N_45497,N_45498,N_45499,N_45500,N_45501,N_45502,N_45503,N_45504,N_45505,N_45506,N_45507,N_45508,N_45509,N_45510,N_45511,N_45512,N_45513,N_45514,N_45515,N_45516,N_45517,N_45518,N_45519,N_45520,N_45521,N_45522,N_45523,N_45524,N_45525,N_45526,N_45527,N_45528,N_45529,N_45530,N_45531,N_45532,N_45533,N_45534,N_45535,N_45536,N_45537,N_45538,N_45539,N_45540,N_45541,N_45542,N_45543,N_45544,N_45545,N_45546,N_45547,N_45548,N_45549,N_45550,N_45551,N_45552,N_45553,N_45554,N_45555,N_45556,N_45557,N_45558,N_45559,N_45560,N_45561,N_45562,N_45563,N_45564,N_45565,N_45566,N_45567,N_45568,N_45569,N_45570,N_45571,N_45572,N_45573,N_45574,N_45575,N_45576,N_45577,N_45578,N_45579,N_45580,N_45581,N_45582,N_45583,N_45584,N_45585,N_45586,N_45587,N_45588,N_45589,N_45590,N_45591,N_45592,N_45593,N_45594,N_45595,N_45596,N_45597,N_45598,N_45599,N_45600,N_45601,N_45602,N_45603,N_45604,N_45605,N_45606,N_45607,N_45608,N_45609,N_45610,N_45611,N_45612,N_45613,N_45614,N_45615,N_45616,N_45617,N_45618,N_45619,N_45620,N_45621,N_45622,N_45623,N_45624,N_45625,N_45626,N_45627,N_45628,N_45629,N_45630,N_45631,N_45632,N_45633,N_45634,N_45635,N_45636,N_45637,N_45638,N_45639,N_45640,N_45641,N_45642,N_45643,N_45644,N_45645,N_45646,N_45647,N_45648,N_45649,N_45650,N_45651,N_45652,N_45653,N_45654,N_45655,N_45656,N_45657,N_45658,N_45659,N_45660,N_45661,N_45662,N_45663,N_45664,N_45665,N_45666,N_45667,N_45668,N_45669,N_45670,N_45671,N_45672,N_45673,N_45674,N_45675,N_45676,N_45677,N_45678,N_45679,N_45680,N_45681,N_45682,N_45683,N_45684,N_45685,N_45686,N_45687,N_45688,N_45689,N_45690,N_45691,N_45692,N_45693,N_45694,N_45695,N_45696,N_45697,N_45698,N_45699,N_45700,N_45701,N_45702,N_45703,N_45704,N_45705,N_45706,N_45707,N_45708,N_45709,N_45710,N_45711,N_45712,N_45713,N_45714,N_45715,N_45716,N_45717,N_45718,N_45719,N_45720,N_45721,N_45722,N_45723,N_45724,N_45725,N_45726,N_45727,N_45728,N_45729,N_45730,N_45731,N_45732,N_45733,N_45734,N_45735,N_45736,N_45737,N_45738,N_45739,N_45740,N_45741,N_45742,N_45743,N_45744,N_45745,N_45746,N_45747,N_45748,N_45749,N_45750,N_45751,N_45752,N_45753,N_45754,N_45755,N_45756,N_45757,N_45758,N_45759,N_45760,N_45761,N_45762,N_45763,N_45764,N_45765,N_45766,N_45767,N_45768,N_45769,N_45770,N_45771,N_45772,N_45773,N_45774,N_45775,N_45776,N_45777,N_45778,N_45779,N_45780,N_45781,N_45782,N_45783,N_45784,N_45785,N_45786,N_45787,N_45788,N_45789,N_45790,N_45791,N_45792,N_45793,N_45794,N_45795,N_45796,N_45797,N_45798,N_45799,N_45800,N_45801,N_45802,N_45803,N_45804,N_45805,N_45806,N_45807,N_45808,N_45809,N_45810,N_45811,N_45812,N_45813,N_45814,N_45815,N_45816,N_45817,N_45818,N_45819,N_45820,N_45821,N_45822,N_45823,N_45824,N_45825,N_45826,N_45827,N_45828,N_45829,N_45830,N_45831,N_45832,N_45833,N_45834,N_45835,N_45836,N_45837,N_45838,N_45839,N_45840,N_45841,N_45842,N_45843,N_45844,N_45845,N_45846,N_45847,N_45848,N_45849,N_45850,N_45851,N_45852,N_45853,N_45854,N_45855,N_45856,N_45857,N_45858,N_45859,N_45860,N_45861,N_45862,N_45863,N_45864,N_45865,N_45866,N_45867,N_45868,N_45869,N_45870,N_45871,N_45872,N_45873,N_45874,N_45875,N_45876,N_45877,N_45878,N_45879,N_45880,N_45881,N_45882,N_45883,N_45884,N_45885,N_45886,N_45887,N_45888,N_45889,N_45890,N_45891,N_45892,N_45893,N_45894,N_45895,N_45896,N_45897,N_45898,N_45899,N_45900,N_45901,N_45902,N_45903,N_45904,N_45905,N_45906,N_45907,N_45908,N_45909,N_45910,N_45911,N_45912,N_45913,N_45914,N_45915,N_45916,N_45917,N_45918,N_45919,N_45920,N_45921,N_45922,N_45923,N_45924,N_45925,N_45926,N_45927,N_45928,N_45929,N_45930,N_45931,N_45932,N_45933,N_45934,N_45935,N_45936,N_45937,N_45938,N_45939,N_45940,N_45941,N_45942,N_45943,N_45944,N_45945,N_45946,N_45947,N_45948,N_45949,N_45950,N_45951,N_45952,N_45953,N_45954,N_45955,N_45956,N_45957,N_45958,N_45959,N_45960,N_45961,N_45962,N_45963,N_45964,N_45965,N_45966,N_45967,N_45968,N_45969,N_45970,N_45971,N_45972,N_45973,N_45974,N_45975,N_45976,N_45977,N_45978,N_45979,N_45980,N_45981,N_45982,N_45983,N_45984,N_45985,N_45986,N_45987,N_45988,N_45989,N_45990,N_45991,N_45992,N_45993,N_45994,N_45995,N_45996,N_45997,N_45998,N_45999,N_46000,N_46001,N_46002,N_46003,N_46004,N_46005,N_46006,N_46007,N_46008,N_46009,N_46010,N_46011,N_46012,N_46013,N_46014,N_46015,N_46016,N_46017,N_46018,N_46019,N_46020,N_46021,N_46022,N_46023,N_46024,N_46025,N_46026,N_46027,N_46028,N_46029,N_46030,N_46031,N_46032,N_46033,N_46034,N_46035,N_46036,N_46037,N_46038,N_46039,N_46040,N_46041,N_46042,N_46043,N_46044,N_46045,N_46046,N_46047,N_46048,N_46049,N_46050,N_46051,N_46052,N_46053,N_46054,N_46055,N_46056,N_46057,N_46058,N_46059,N_46060,N_46061,N_46062,N_46063,N_46064,N_46065,N_46066,N_46067,N_46068,N_46069,N_46070,N_46071,N_46072,N_46073,N_46074,N_46075,N_46076,N_46077,N_46078,N_46079,N_46080,N_46081,N_46082,N_46083,N_46084,N_46085,N_46086,N_46087,N_46088,N_46089,N_46090,N_46091,N_46092,N_46093,N_46094,N_46095,N_46096,N_46097,N_46098,N_46099,N_46100,N_46101,N_46102,N_46103,N_46104,N_46105,N_46106,N_46107,N_46108,N_46109,N_46110,N_46111,N_46112,N_46113,N_46114,N_46115,N_46116,N_46117,N_46118,N_46119,N_46120,N_46121,N_46122,N_46123,N_46124,N_46125,N_46126,N_46127,N_46128,N_46129,N_46130,N_46131,N_46132,N_46133,N_46134,N_46135,N_46136,N_46137,N_46138,N_46139,N_46140,N_46141,N_46142,N_46143,N_46144,N_46145,N_46146,N_46147,N_46148,N_46149,N_46150,N_46151,N_46152,N_46153,N_46154,N_46155,N_46156,N_46157,N_46158,N_46159,N_46160,N_46161,N_46162,N_46163,N_46164,N_46165,N_46166,N_46167,N_46168,N_46169,N_46170,N_46171,N_46172,N_46173,N_46174,N_46175,N_46176,N_46177,N_46178,N_46179,N_46180,N_46181,N_46182,N_46183,N_46184,N_46185,N_46186,N_46187,N_46188,N_46189,N_46190,N_46191,N_46192,N_46193,N_46194,N_46195,N_46196,N_46197,N_46198,N_46199,N_46200,N_46201,N_46202,N_46203,N_46204,N_46205,N_46206,N_46207,N_46208,N_46209,N_46210,N_46211,N_46212,N_46213,N_46214,N_46215,N_46216,N_46217,N_46218,N_46219,N_46220,N_46221,N_46222,N_46223,N_46224,N_46225,N_46226,N_46227,N_46228,N_46229,N_46230,N_46231,N_46232,N_46233,N_46234,N_46235,N_46236,N_46237,N_46238,N_46239,N_46240,N_46241,N_46242,N_46243,N_46244,N_46245,N_46246,N_46247,N_46248,N_46249,N_46250,N_46251,N_46252,N_46253,N_46254,N_46255,N_46256,N_46257,N_46258,N_46259,N_46260,N_46261,N_46262,N_46263,N_46264,N_46265,N_46266,N_46267,N_46268,N_46269,N_46270,N_46271,N_46272,N_46273,N_46274,N_46275,N_46276,N_46277,N_46278,N_46279,N_46280,N_46281,N_46282,N_46283,N_46284,N_46285,N_46286,N_46287,N_46288,N_46289,N_46290,N_46291,N_46292,N_46293,N_46294,N_46295,N_46296,N_46297,N_46298,N_46299,N_46300,N_46301,N_46302,N_46303,N_46304,N_46305,N_46306,N_46307,N_46308,N_46309,N_46310,N_46311,N_46312,N_46313,N_46314,N_46315,N_46316,N_46317,N_46318,N_46319,N_46320,N_46321,N_46322,N_46323,N_46324,N_46325,N_46326,N_46327,N_46328,N_46329,N_46330,N_46331,N_46332,N_46333,N_46334,N_46335,N_46336,N_46337,N_46338,N_46339,N_46340,N_46341,N_46342,N_46343,N_46344,N_46345,N_46346,N_46347,N_46348,N_46349,N_46350,N_46351,N_46352,N_46353,N_46354,N_46355,N_46356,N_46357,N_46358,N_46359,N_46360,N_46361,N_46362,N_46363,N_46364,N_46365,N_46366,N_46367,N_46368,N_46369,N_46370,N_46371,N_46372,N_46373,N_46374,N_46375,N_46376,N_46377,N_46378,N_46379,N_46380,N_46381,N_46382,N_46383,N_46384,N_46385,N_46386,N_46387,N_46388,N_46389,N_46390,N_46391,N_46392,N_46393,N_46394,N_46395,N_46396,N_46397,N_46398,N_46399,N_46400,N_46401,N_46402,N_46403,N_46404,N_46405,N_46406,N_46407,N_46408,N_46409,N_46410,N_46411,N_46412,N_46413,N_46414,N_46415,N_46416,N_46417,N_46418,N_46419,N_46420,N_46421,N_46422,N_46423,N_46424,N_46425,N_46426,N_46427,N_46428,N_46429,N_46430,N_46431,N_46432,N_46433,N_46434,N_46435,N_46436,N_46437,N_46438,N_46439,N_46440,N_46441,N_46442,N_46443,N_46444,N_46445,N_46446,N_46447,N_46448,N_46449,N_46450,N_46451,N_46452,N_46453,N_46454,N_46455,N_46456,N_46457,N_46458,N_46459,N_46460,N_46461,N_46462,N_46463,N_46464,N_46465,N_46466,N_46467,N_46468,N_46469,N_46470,N_46471,N_46472,N_46473,N_46474,N_46475,N_46476,N_46477,N_46478,N_46479,N_46480,N_46481,N_46482,N_46483,N_46484,N_46485,N_46486,N_46487,N_46488,N_46489,N_46490,N_46491,N_46492,N_46493,N_46494,N_46495,N_46496,N_46497,N_46498,N_46499,N_46500,N_46501,N_46502,N_46503,N_46504,N_46505,N_46506,N_46507,N_46508,N_46509,N_46510,N_46511,N_46512,N_46513,N_46514,N_46515,N_46516,N_46517,N_46518,N_46519,N_46520,N_46521,N_46522,N_46523,N_46524,N_46525,N_46526,N_46527,N_46528,N_46529,N_46530,N_46531,N_46532,N_46533,N_46534,N_46535,N_46536,N_46537,N_46538,N_46539,N_46540,N_46541,N_46542,N_46543,N_46544,N_46545,N_46546,N_46547,N_46548,N_46549,N_46550,N_46551,N_46552,N_46553,N_46554,N_46555,N_46556,N_46557,N_46558,N_46559,N_46560,N_46561,N_46562,N_46563,N_46564,N_46565,N_46566,N_46567,N_46568,N_46569,N_46570,N_46571,N_46572,N_46573,N_46574,N_46575,N_46576,N_46577,N_46578,N_46579,N_46580,N_46581,N_46582,N_46583,N_46584,N_46585,N_46586,N_46587,N_46588,N_46589,N_46590,N_46591,N_46592,N_46593,N_46594,N_46595,N_46596,N_46597,N_46598,N_46599,N_46600,N_46601,N_46602,N_46603,N_46604,N_46605,N_46606,N_46607,N_46608,N_46609,N_46610,N_46611,N_46612,N_46613,N_46614,N_46615,N_46616,N_46617,N_46618,N_46619,N_46620,N_46621,N_46622,N_46623,N_46624,N_46625,N_46626,N_46627,N_46628,N_46629,N_46630,N_46631,N_46632,N_46633,N_46634,N_46635,N_46636,N_46637,N_46638,N_46639,N_46640,N_46641,N_46642,N_46643,N_46644,N_46645,N_46646,N_46647,N_46648,N_46649,N_46650,N_46651,N_46652,N_46653,N_46654,N_46655,N_46656,N_46657,N_46658,N_46659,N_46660,N_46661,N_46662,N_46663,N_46664,N_46665,N_46666,N_46667,N_46668,N_46669,N_46670,N_46671,N_46672,N_46673,N_46674,N_46675,N_46676,N_46677,N_46678,N_46679,N_46680,N_46681,N_46682,N_46683,N_46684,N_46685,N_46686,N_46687,N_46688,N_46689,N_46690,N_46691,N_46692,N_46693,N_46694,N_46695,N_46696,N_46697,N_46698,N_46699,N_46700,N_46701,N_46702,N_46703,N_46704,N_46705,N_46706,N_46707,N_46708,N_46709,N_46710,N_46711,N_46712,N_46713,N_46714,N_46715,N_46716,N_46717,N_46718,N_46719,N_46720,N_46721,N_46722,N_46723,N_46724,N_46725,N_46726,N_46727,N_46728,N_46729,N_46730,N_46731,N_46732,N_46733,N_46734,N_46735,N_46736,N_46737,N_46738,N_46739,N_46740,N_46741,N_46742,N_46743,N_46744,N_46745,N_46746,N_46747,N_46748,N_46749,N_46750,N_46751,N_46752,N_46753,N_46754,N_46755,N_46756,N_46757,N_46758,N_46759,N_46760,N_46761,N_46762,N_46763,N_46764,N_46765,N_46766,N_46767,N_46768,N_46769,N_46770,N_46771,N_46772,N_46773,N_46774,N_46775,N_46776,N_46777,N_46778,N_46779,N_46780,N_46781,N_46782,N_46783,N_46784,N_46785,N_46786,N_46787,N_46788,N_46789,N_46790,N_46791,N_46792,N_46793,N_46794,N_46795,N_46796,N_46797,N_46798,N_46799,N_46800,N_46801,N_46802,N_46803,N_46804,N_46805,N_46806,N_46807,N_46808,N_46809,N_46810,N_46811,N_46812,N_46813,N_46814,N_46815,N_46816,N_46817,N_46818,N_46819,N_46820,N_46821,N_46822,N_46823,N_46824,N_46825,N_46826,N_46827,N_46828,N_46829,N_46830,N_46831,N_46832,N_46833,N_46834,N_46835,N_46836,N_46837,N_46838,N_46839,N_46840,N_46841,N_46842,N_46843,N_46844,N_46845,N_46846,N_46847,N_46848,N_46849,N_46850,N_46851,N_46852,N_46853,N_46854,N_46855,N_46856,N_46857,N_46858,N_46859,N_46860,N_46861,N_46862,N_46863,N_46864,N_46865,N_46866,N_46867,N_46868,N_46869,N_46870,N_46871,N_46872,N_46873,N_46874,N_46875,N_46876,N_46877,N_46878,N_46879,N_46880,N_46881,N_46882,N_46883,N_46884,N_46885,N_46886,N_46887,N_46888,N_46889,N_46890,N_46891,N_46892,N_46893,N_46894,N_46895,N_46896,N_46897,N_46898,N_46899,N_46900,N_46901,N_46902,N_46903,N_46904,N_46905,N_46906,N_46907,N_46908,N_46909,N_46910,N_46911,N_46912,N_46913,N_46914,N_46915,N_46916,N_46917,N_46918,N_46919,N_46920,N_46921,N_46922,N_46923,N_46924,N_46925,N_46926,N_46927,N_46928,N_46929,N_46930,N_46931,N_46932,N_46933,N_46934,N_46935,N_46936,N_46937,N_46938,N_46939,N_46940,N_46941,N_46942,N_46943,N_46944,N_46945,N_46946,N_46947,N_46948,N_46949,N_46950,N_46951,N_46952,N_46953,N_46954,N_46955,N_46956,N_46957,N_46958,N_46959,N_46960,N_46961,N_46962,N_46963,N_46964,N_46965,N_46966,N_46967,N_46968,N_46969,N_46970,N_46971,N_46972,N_46973,N_46974,N_46975,N_46976,N_46977,N_46978,N_46979,N_46980,N_46981,N_46982,N_46983,N_46984,N_46985,N_46986,N_46987,N_46988,N_46989,N_46990,N_46991,N_46992,N_46993,N_46994,N_46995,N_46996,N_46997,N_46998,N_46999,N_47000,N_47001,N_47002,N_47003,N_47004,N_47005,N_47006,N_47007,N_47008,N_47009,N_47010,N_47011,N_47012,N_47013,N_47014,N_47015,N_47016,N_47017,N_47018,N_47019,N_47020,N_47021,N_47022,N_47023,N_47024,N_47025,N_47026,N_47027,N_47028,N_47029,N_47030,N_47031,N_47032,N_47033,N_47034,N_47035,N_47036,N_47037,N_47038,N_47039,N_47040,N_47041,N_47042,N_47043,N_47044,N_47045,N_47046,N_47047,N_47048,N_47049,N_47050,N_47051,N_47052,N_47053,N_47054,N_47055,N_47056,N_47057,N_47058,N_47059,N_47060,N_47061,N_47062,N_47063,N_47064,N_47065,N_47066,N_47067,N_47068,N_47069,N_47070,N_47071,N_47072,N_47073,N_47074,N_47075,N_47076,N_47077,N_47078,N_47079,N_47080,N_47081,N_47082,N_47083,N_47084,N_47085,N_47086,N_47087,N_47088,N_47089,N_47090,N_47091,N_47092,N_47093,N_47094,N_47095,N_47096,N_47097,N_47098,N_47099,N_47100,N_47101,N_47102,N_47103,N_47104,N_47105,N_47106,N_47107,N_47108,N_47109,N_47110,N_47111,N_47112,N_47113,N_47114,N_47115,N_47116,N_47117,N_47118,N_47119,N_47120,N_47121,N_47122,N_47123,N_47124,N_47125,N_47126,N_47127,N_47128,N_47129,N_47130,N_47131,N_47132,N_47133,N_47134,N_47135,N_47136,N_47137,N_47138,N_47139,N_47140,N_47141,N_47142,N_47143,N_47144,N_47145,N_47146,N_47147,N_47148,N_47149,N_47150,N_47151,N_47152,N_47153,N_47154,N_47155,N_47156,N_47157,N_47158,N_47159,N_47160,N_47161,N_47162,N_47163,N_47164,N_47165,N_47166,N_47167,N_47168,N_47169,N_47170,N_47171,N_47172,N_47173,N_47174,N_47175,N_47176,N_47177,N_47178,N_47179,N_47180,N_47181,N_47182,N_47183,N_47184,N_47185,N_47186,N_47187,N_47188,N_47189,N_47190,N_47191,N_47192,N_47193,N_47194,N_47195,N_47196,N_47197,N_47198,N_47199,N_47200,N_47201,N_47202,N_47203,N_47204,N_47205,N_47206,N_47207,N_47208,N_47209,N_47210,N_47211,N_47212,N_47213,N_47214,N_47215,N_47216,N_47217,N_47218,N_47219,N_47220,N_47221,N_47222,N_47223,N_47224,N_47225,N_47226,N_47227,N_47228,N_47229,N_47230,N_47231,N_47232,N_47233,N_47234,N_47235,N_47236,N_47237,N_47238,N_47239,N_47240,N_47241,N_47242,N_47243,N_47244,N_47245,N_47246,N_47247,N_47248,N_47249,N_47250,N_47251,N_47252,N_47253,N_47254,N_47255,N_47256,N_47257,N_47258,N_47259,N_47260,N_47261,N_47262,N_47263,N_47264,N_47265,N_47266,N_47267,N_47268,N_47269,N_47270,N_47271,N_47272,N_47273,N_47274,N_47275,N_47276,N_47277,N_47278,N_47279,N_47280,N_47281,N_47282,N_47283,N_47284,N_47285,N_47286,N_47287,N_47288,N_47289,N_47290,N_47291,N_47292,N_47293,N_47294,N_47295,N_47296,N_47297,N_47298,N_47299,N_47300,N_47301,N_47302,N_47303,N_47304,N_47305,N_47306,N_47307,N_47308,N_47309,N_47310,N_47311,N_47312,N_47313,N_47314,N_47315,N_47316,N_47317,N_47318,N_47319,N_47320,N_47321,N_47322,N_47323,N_47324,N_47325,N_47326,N_47327,N_47328,N_47329,N_47330,N_47331,N_47332,N_47333,N_47334,N_47335,N_47336,N_47337,N_47338,N_47339,N_47340,N_47341,N_47342,N_47343,N_47344,N_47345,N_47346,N_47347,N_47348,N_47349,N_47350,N_47351,N_47352,N_47353,N_47354,N_47355,N_47356,N_47357,N_47358,N_47359,N_47360,N_47361,N_47362,N_47363,N_47364,N_47365,N_47366,N_47367,N_47368,N_47369,N_47370,N_47371,N_47372,N_47373,N_47374,N_47375,N_47376,N_47377,N_47378,N_47379,N_47380,N_47381,N_47382,N_47383,N_47384,N_47385,N_47386,N_47387,N_47388,N_47389,N_47390,N_47391,N_47392,N_47393,N_47394,N_47395,N_47396,N_47397,N_47398,N_47399,N_47400,N_47401,N_47402,N_47403,N_47404,N_47405,N_47406,N_47407,N_47408,N_47409,N_47410,N_47411,N_47412,N_47413,N_47414,N_47415,N_47416,N_47417,N_47418,N_47419,N_47420,N_47421,N_47422,N_47423,N_47424,N_47425,N_47426,N_47427,N_47428,N_47429,N_47430,N_47431,N_47432,N_47433,N_47434,N_47435,N_47436,N_47437,N_47438,N_47439,N_47440,N_47441,N_47442,N_47443,N_47444,N_47445,N_47446,N_47447,N_47448,N_47449,N_47450,N_47451,N_47452,N_47453,N_47454,N_47455,N_47456,N_47457,N_47458,N_47459,N_47460,N_47461,N_47462,N_47463,N_47464,N_47465,N_47466,N_47467,N_47468,N_47469,N_47470,N_47471,N_47472,N_47473,N_47474,N_47475,N_47476,N_47477,N_47478,N_47479,N_47480,N_47481,N_47482,N_47483,N_47484,N_47485,N_47486,N_47487,N_47488,N_47489,N_47490,N_47491,N_47492,N_47493,N_47494,N_47495,N_47496,N_47497,N_47498,N_47499,N_47500,N_47501,N_47502,N_47503,N_47504,N_47505,N_47506,N_47507,N_47508,N_47509,N_47510,N_47511,N_47512,N_47513,N_47514,N_47515,N_47516,N_47517,N_47518,N_47519,N_47520,N_47521,N_47522,N_47523,N_47524,N_47525,N_47526,N_47527,N_47528,N_47529,N_47530,N_47531,N_47532,N_47533,N_47534,N_47535,N_47536,N_47537,N_47538,N_47539,N_47540,N_47541,N_47542,N_47543,N_47544,N_47545,N_47546,N_47547,N_47548,N_47549,N_47550,N_47551,N_47552,N_47553,N_47554,N_47555,N_47556,N_47557,N_47558,N_47559,N_47560,N_47561,N_47562,N_47563,N_47564,N_47565,N_47566,N_47567,N_47568,N_47569,N_47570,N_47571,N_47572,N_47573,N_47574,N_47575,N_47576,N_47577,N_47578,N_47579,N_47580,N_47581,N_47582,N_47583,N_47584,N_47585,N_47586,N_47587,N_47588,N_47589,N_47590,N_47591,N_47592,N_47593,N_47594,N_47595,N_47596,N_47597,N_47598,N_47599,N_47600,N_47601,N_47602,N_47603,N_47604,N_47605,N_47606,N_47607,N_47608,N_47609,N_47610,N_47611,N_47612,N_47613,N_47614,N_47615,N_47616,N_47617,N_47618,N_47619,N_47620,N_47621,N_47622,N_47623,N_47624,N_47625,N_47626,N_47627,N_47628,N_47629,N_47630,N_47631,N_47632,N_47633,N_47634,N_47635,N_47636,N_47637,N_47638,N_47639,N_47640,N_47641,N_47642,N_47643,N_47644,N_47645,N_47646,N_47647,N_47648,N_47649,N_47650,N_47651,N_47652,N_47653,N_47654,N_47655,N_47656,N_47657,N_47658,N_47659,N_47660,N_47661,N_47662,N_47663,N_47664,N_47665,N_47666,N_47667,N_47668,N_47669,N_47670,N_47671,N_47672,N_47673,N_47674,N_47675,N_47676,N_47677,N_47678,N_47679,N_47680,N_47681,N_47682,N_47683,N_47684,N_47685,N_47686,N_47687,N_47688,N_47689,N_47690,N_47691,N_47692,N_47693,N_47694,N_47695,N_47696,N_47697,N_47698,N_47699,N_47700,N_47701,N_47702,N_47703,N_47704,N_47705,N_47706,N_47707,N_47708,N_47709,N_47710,N_47711,N_47712,N_47713,N_47714,N_47715,N_47716,N_47717,N_47718,N_47719,N_47720,N_47721,N_47722,N_47723,N_47724,N_47725,N_47726,N_47727,N_47728,N_47729,N_47730,N_47731,N_47732,N_47733,N_47734,N_47735,N_47736,N_47737,N_47738,N_47739,N_47740,N_47741,N_47742,N_47743,N_47744,N_47745,N_47746,N_47747,N_47748,N_47749,N_47750,N_47751,N_47752,N_47753,N_47754,N_47755,N_47756,N_47757,N_47758,N_47759,N_47760,N_47761,N_47762,N_47763,N_47764,N_47765,N_47766,N_47767,N_47768,N_47769,N_47770,N_47771,N_47772,N_47773,N_47774,N_47775,N_47776,N_47777,N_47778,N_47779,N_47780,N_47781,N_47782,N_47783,N_47784,N_47785,N_47786,N_47787,N_47788,N_47789,N_47790,N_47791,N_47792,N_47793,N_47794,N_47795,N_47796,N_47797,N_47798,N_47799,N_47800,N_47801,N_47802,N_47803,N_47804,N_47805,N_47806,N_47807,N_47808,N_47809,N_47810,N_47811,N_47812,N_47813,N_47814,N_47815,N_47816,N_47817,N_47818,N_47819,N_47820,N_47821,N_47822,N_47823,N_47824,N_47825,N_47826,N_47827,N_47828,N_47829,N_47830,N_47831,N_47832,N_47833,N_47834,N_47835,N_47836,N_47837,N_47838,N_47839,N_47840,N_47841,N_47842,N_47843,N_47844,N_47845,N_47846,N_47847,N_47848,N_47849,N_47850,N_47851,N_47852,N_47853,N_47854,N_47855,N_47856,N_47857,N_47858,N_47859,N_47860,N_47861,N_47862,N_47863,N_47864,N_47865,N_47866,N_47867,N_47868,N_47869,N_47870,N_47871,N_47872,N_47873,N_47874,N_47875,N_47876,N_47877,N_47878,N_47879,N_47880,N_47881,N_47882,N_47883,N_47884,N_47885,N_47886,N_47887,N_47888,N_47889,N_47890,N_47891,N_47892,N_47893,N_47894,N_47895,N_47896,N_47897,N_47898,N_47899,N_47900,N_47901,N_47902,N_47903,N_47904,N_47905,N_47906,N_47907,N_47908,N_47909,N_47910,N_47911,N_47912,N_47913,N_47914,N_47915,N_47916,N_47917,N_47918,N_47919,N_47920,N_47921,N_47922,N_47923,N_47924,N_47925,N_47926,N_47927,N_47928,N_47929,N_47930,N_47931,N_47932,N_47933,N_47934,N_47935,N_47936,N_47937,N_47938,N_47939,N_47940,N_47941,N_47942,N_47943,N_47944,N_47945,N_47946,N_47947,N_47948,N_47949,N_47950,N_47951,N_47952,N_47953,N_47954,N_47955,N_47956,N_47957,N_47958,N_47959,N_47960,N_47961,N_47962,N_47963,N_47964,N_47965,N_47966,N_47967,N_47968,N_47969,N_47970,N_47971,N_47972,N_47973,N_47974,N_47975,N_47976,N_47977,N_47978,N_47979,N_47980,N_47981,N_47982,N_47983,N_47984,N_47985,N_47986,N_47987,N_47988,N_47989,N_47990,N_47991,N_47992,N_47993,N_47994,N_47995,N_47996,N_47997,N_47998,N_47999,N_48000,N_48001,N_48002,N_48003,N_48004,N_48005,N_48006,N_48007,N_48008,N_48009,N_48010,N_48011,N_48012,N_48013,N_48014,N_48015,N_48016,N_48017,N_48018,N_48019,N_48020,N_48021,N_48022,N_48023,N_48024,N_48025,N_48026,N_48027,N_48028,N_48029,N_48030,N_48031,N_48032,N_48033,N_48034,N_48035,N_48036,N_48037,N_48038,N_48039,N_48040,N_48041,N_48042,N_48043,N_48044,N_48045,N_48046,N_48047,N_48048,N_48049,N_48050,N_48051,N_48052,N_48053,N_48054,N_48055,N_48056,N_48057,N_48058,N_48059,N_48060,N_48061,N_48062,N_48063,N_48064,N_48065,N_48066,N_48067,N_48068,N_48069,N_48070,N_48071,N_48072,N_48073,N_48074,N_48075,N_48076,N_48077,N_48078,N_48079,N_48080,N_48081,N_48082,N_48083,N_48084,N_48085,N_48086,N_48087,N_48088,N_48089,N_48090,N_48091,N_48092,N_48093,N_48094,N_48095,N_48096,N_48097,N_48098,N_48099,N_48100,N_48101,N_48102,N_48103,N_48104,N_48105,N_48106,N_48107,N_48108,N_48109,N_48110,N_48111,N_48112,N_48113,N_48114,N_48115,N_48116,N_48117,N_48118,N_48119,N_48120,N_48121,N_48122,N_48123,N_48124,N_48125,N_48126,N_48127,N_48128,N_48129,N_48130,N_48131,N_48132,N_48133,N_48134,N_48135,N_48136,N_48137,N_48138,N_48139,N_48140,N_48141,N_48142,N_48143,N_48144,N_48145,N_48146,N_48147,N_48148,N_48149,N_48150,N_48151,N_48152,N_48153,N_48154,N_48155,N_48156,N_48157,N_48158,N_48159,N_48160,N_48161,N_48162,N_48163,N_48164,N_48165,N_48166,N_48167,N_48168,N_48169,N_48170,N_48171,N_48172,N_48173,N_48174,N_48175,N_48176,N_48177,N_48178,N_48179,N_48180,N_48181,N_48182,N_48183,N_48184,N_48185,N_48186,N_48187,N_48188,N_48189,N_48190,N_48191,N_48192,N_48193,N_48194,N_48195,N_48196,N_48197,N_48198,N_48199,N_48200,N_48201,N_48202,N_48203,N_48204,N_48205,N_48206,N_48207,N_48208,N_48209,N_48210,N_48211,N_48212,N_48213,N_48214,N_48215,N_48216,N_48217,N_48218,N_48219,N_48220,N_48221,N_48222,N_48223,N_48224,N_48225,N_48226,N_48227,N_48228,N_48229,N_48230,N_48231,N_48232,N_48233,N_48234,N_48235,N_48236,N_48237,N_48238,N_48239,N_48240,N_48241,N_48242,N_48243,N_48244,N_48245,N_48246,N_48247,N_48248,N_48249,N_48250,N_48251,N_48252,N_48253,N_48254,N_48255,N_48256,N_48257,N_48258,N_48259,N_48260,N_48261,N_48262,N_48263,N_48264,N_48265,N_48266,N_48267,N_48268,N_48269,N_48270,N_48271,N_48272,N_48273,N_48274,N_48275,N_48276,N_48277,N_48278,N_48279,N_48280,N_48281,N_48282,N_48283,N_48284,N_48285,N_48286,N_48287,N_48288,N_48289,N_48290,N_48291,N_48292,N_48293,N_48294,N_48295,N_48296,N_48297,N_48298,N_48299,N_48300,N_48301,N_48302,N_48303,N_48304,N_48305,N_48306,N_48307,N_48308,N_48309,N_48310,N_48311,N_48312,N_48313,N_48314,N_48315,N_48316,N_48317,N_48318,N_48319,N_48320,N_48321,N_48322,N_48323,N_48324,N_48325,N_48326,N_48327,N_48328,N_48329,N_48330,N_48331,N_48332,N_48333,N_48334,N_48335,N_48336,N_48337,N_48338,N_48339,N_48340,N_48341,N_48342,N_48343,N_48344,N_48345,N_48346,N_48347,N_48348,N_48349,N_48350,N_48351,N_48352,N_48353,N_48354,N_48355,N_48356,N_48357,N_48358,N_48359,N_48360,N_48361,N_48362,N_48363,N_48364,N_48365,N_48366,N_48367,N_48368,N_48369,N_48370,N_48371,N_48372,N_48373,N_48374,N_48375,N_48376,N_48377,N_48378,N_48379,N_48380,N_48381,N_48382,N_48383,N_48384,N_48385,N_48386,N_48387,N_48388,N_48389,N_48390,N_48391,N_48392,N_48393,N_48394,N_48395,N_48396,N_48397,N_48398,N_48399,N_48400,N_48401,N_48402,N_48403,N_48404,N_48405,N_48406,N_48407,N_48408,N_48409,N_48410,N_48411,N_48412,N_48413,N_48414,N_48415,N_48416,N_48417,N_48418,N_48419,N_48420,N_48421,N_48422,N_48423,N_48424,N_48425,N_48426,N_48427,N_48428,N_48429,N_48430,N_48431,N_48432,N_48433,N_48434,N_48435,N_48436,N_48437,N_48438,N_48439,N_48440,N_48441,N_48442,N_48443,N_48444,N_48445,N_48446,N_48447,N_48448,N_48449,N_48450,N_48451,N_48452,N_48453,N_48454,N_48455,N_48456,N_48457,N_48458,N_48459,N_48460,N_48461,N_48462,N_48463,N_48464,N_48465,N_48466,N_48467,N_48468,N_48469,N_48470,N_48471,N_48472,N_48473,N_48474,N_48475,N_48476,N_48477,N_48478,N_48479,N_48480,N_48481,N_48482,N_48483,N_48484,N_48485,N_48486,N_48487,N_48488,N_48489,N_48490,N_48491,N_48492,N_48493,N_48494,N_48495,N_48496,N_48497,N_48498,N_48499,N_48500,N_48501,N_48502,N_48503,N_48504,N_48505,N_48506,N_48507,N_48508,N_48509,N_48510,N_48511,N_48512,N_48513,N_48514,N_48515,N_48516,N_48517,N_48518,N_48519,N_48520,N_48521,N_48522,N_48523,N_48524,N_48525,N_48526,N_48527,N_48528,N_48529,N_48530,N_48531,N_48532,N_48533,N_48534,N_48535,N_48536,N_48537,N_48538,N_48539,N_48540,N_48541,N_48542,N_48543,N_48544,N_48545,N_48546,N_48547,N_48548,N_48549,N_48550,N_48551,N_48552,N_48553,N_48554,N_48555,N_48556,N_48557,N_48558,N_48559,N_48560,N_48561,N_48562,N_48563,N_48564,N_48565,N_48566,N_48567,N_48568,N_48569,N_48570,N_48571,N_48572,N_48573,N_48574,N_48575,N_48576,N_48577,N_48578,N_48579,N_48580,N_48581,N_48582,N_48583,N_48584,N_48585,N_48586,N_48587,N_48588,N_48589,N_48590,N_48591,N_48592,N_48593,N_48594,N_48595,N_48596,N_48597,N_48598,N_48599,N_48600,N_48601,N_48602,N_48603,N_48604,N_48605,N_48606,N_48607,N_48608,N_48609,N_48610,N_48611,N_48612,N_48613,N_48614,N_48615,N_48616,N_48617,N_48618,N_48619,N_48620,N_48621,N_48622,N_48623,N_48624,N_48625,N_48626,N_48627,N_48628,N_48629,N_48630,N_48631,N_48632,N_48633,N_48634,N_48635,N_48636,N_48637,N_48638,N_48639,N_48640,N_48641,N_48642,N_48643,N_48644,N_48645,N_48646,N_48647,N_48648,N_48649,N_48650,N_48651,N_48652,N_48653,N_48654,N_48655,N_48656,N_48657,N_48658,N_48659,N_48660,N_48661,N_48662,N_48663,N_48664,N_48665,N_48666,N_48667,N_48668,N_48669,N_48670,N_48671,N_48672,N_48673,N_48674,N_48675,N_48676,N_48677,N_48678,N_48679,N_48680,N_48681,N_48682,N_48683,N_48684,N_48685,N_48686,N_48687,N_48688,N_48689,N_48690,N_48691,N_48692,N_48693,N_48694,N_48695,N_48696,N_48697,N_48698,N_48699,N_48700,N_48701,N_48702,N_48703,N_48704,N_48705,N_48706,N_48707,N_48708,N_48709,N_48710,N_48711,N_48712,N_48713,N_48714,N_48715,N_48716,N_48717,N_48718,N_48719,N_48720,N_48721,N_48722,N_48723,N_48724,N_48725,N_48726,N_48727,N_48728,N_48729,N_48730,N_48731,N_48732,N_48733,N_48734,N_48735,N_48736,N_48737,N_48738,N_48739,N_48740,N_48741,N_48742,N_48743,N_48744,N_48745,N_48746,N_48747,N_48748,N_48749,N_48750,N_48751,N_48752,N_48753,N_48754,N_48755,N_48756,N_48757,N_48758,N_48759,N_48760,N_48761,N_48762,N_48763,N_48764,N_48765,N_48766,N_48767,N_48768,N_48769,N_48770,N_48771,N_48772,N_48773,N_48774,N_48775,N_48776,N_48777,N_48778,N_48779,N_48780,N_48781,N_48782,N_48783,N_48784,N_48785,N_48786,N_48787,N_48788,N_48789,N_48790,N_48791,N_48792,N_48793,N_48794,N_48795,N_48796,N_48797,N_48798,N_48799,N_48800,N_48801,N_48802,N_48803,N_48804,N_48805,N_48806,N_48807,N_48808,N_48809,N_48810,N_48811,N_48812,N_48813,N_48814,N_48815,N_48816,N_48817,N_48818,N_48819,N_48820,N_48821,N_48822,N_48823,N_48824,N_48825,N_48826,N_48827,N_48828,N_48829,N_48830,N_48831,N_48832,N_48833,N_48834,N_48835,N_48836,N_48837,N_48838,N_48839,N_48840,N_48841,N_48842,N_48843,N_48844,N_48845,N_48846,N_48847,N_48848,N_48849,N_48850,N_48851,N_48852,N_48853,N_48854,N_48855,N_48856,N_48857,N_48858,N_48859,N_48860,N_48861,N_48862,N_48863,N_48864,N_48865,N_48866,N_48867,N_48868,N_48869,N_48870,N_48871,N_48872,N_48873,N_48874,N_48875,N_48876,N_48877,N_48878,N_48879,N_48880,N_48881,N_48882,N_48883,N_48884,N_48885,N_48886,N_48887,N_48888,N_48889,N_48890,N_48891,N_48892,N_48893,N_48894,N_48895,N_48896,N_48897,N_48898,N_48899,N_48900,N_48901,N_48902,N_48903,N_48904,N_48905,N_48906,N_48907,N_48908,N_48909,N_48910,N_48911,N_48912,N_48913,N_48914,N_48915,N_48916,N_48917,N_48918,N_48919,N_48920,N_48921,N_48922,N_48923,N_48924,N_48925,N_48926,N_48927,N_48928,N_48929,N_48930,N_48931,N_48932,N_48933,N_48934,N_48935,N_48936,N_48937,N_48938,N_48939,N_48940,N_48941,N_48942,N_48943,N_48944,N_48945,N_48946,N_48947,N_48948,N_48949,N_48950,N_48951,N_48952,N_48953,N_48954,N_48955,N_48956,N_48957,N_48958,N_48959,N_48960,N_48961,N_48962,N_48963,N_48964,N_48965,N_48966,N_48967,N_48968,N_48969,N_48970,N_48971,N_48972,N_48973,N_48974,N_48975,N_48976,N_48977,N_48978,N_48979,N_48980,N_48981,N_48982,N_48983,N_48984,N_48985,N_48986,N_48987,N_48988,N_48989,N_48990,N_48991,N_48992,N_48993,N_48994,N_48995,N_48996,N_48997,N_48998,N_48999,N_49000,N_49001,N_49002,N_49003,N_49004,N_49005,N_49006,N_49007,N_49008,N_49009,N_49010,N_49011,N_49012,N_49013,N_49014,N_49015,N_49016,N_49017,N_49018,N_49019,N_49020,N_49021,N_49022,N_49023,N_49024,N_49025,N_49026,N_49027,N_49028,N_49029,N_49030,N_49031,N_49032,N_49033,N_49034,N_49035,N_49036,N_49037,N_49038,N_49039,N_49040,N_49041,N_49042,N_49043,N_49044,N_49045,N_49046,N_49047,N_49048,N_49049,N_49050,N_49051,N_49052,N_49053,N_49054,N_49055,N_49056,N_49057,N_49058,N_49059,N_49060,N_49061,N_49062,N_49063,N_49064,N_49065,N_49066,N_49067,N_49068,N_49069,N_49070,N_49071,N_49072,N_49073,N_49074,N_49075,N_49076,N_49077,N_49078,N_49079,N_49080,N_49081,N_49082,N_49083,N_49084,N_49085,N_49086,N_49087,N_49088,N_49089,N_49090,N_49091,N_49092,N_49093,N_49094,N_49095,N_49096,N_49097,N_49098,N_49099,N_49100,N_49101,N_49102,N_49103,N_49104,N_49105,N_49106,N_49107,N_49108,N_49109,N_49110,N_49111,N_49112,N_49113,N_49114,N_49115,N_49116,N_49117,N_49118,N_49119,N_49120,N_49121,N_49122,N_49123,N_49124,N_49125,N_49126,N_49127,N_49128,N_49129,N_49130,N_49131,N_49132,N_49133,N_49134,N_49135,N_49136,N_49137,N_49138,N_49139,N_49140,N_49141,N_49142,N_49143,N_49144,N_49145,N_49146,N_49147,N_49148,N_49149,N_49150,N_49151,N_49152,N_49153,N_49154,N_49155,N_49156,N_49157,N_49158,N_49159,N_49160,N_49161,N_49162,N_49163,N_49164,N_49165,N_49166,N_49167,N_49168,N_49169,N_49170,N_49171,N_49172,N_49173,N_49174,N_49175,N_49176,N_49177,N_49178,N_49179,N_49180,N_49181,N_49182,N_49183,N_49184,N_49185,N_49186,N_49187,N_49188,N_49189,N_49190,N_49191,N_49192,N_49193,N_49194,N_49195,N_49196,N_49197,N_49198,N_49199,N_49200,N_49201,N_49202,N_49203,N_49204,N_49205,N_49206,N_49207,N_49208,N_49209,N_49210,N_49211,N_49212,N_49213,N_49214,N_49215,N_49216,N_49217,N_49218,N_49219,N_49220,N_49221,N_49222,N_49223,N_49224,N_49225,N_49226,N_49227,N_49228,N_49229,N_49230,N_49231,N_49232,N_49233,N_49234,N_49235,N_49236,N_49237,N_49238,N_49239,N_49240,N_49241,N_49242,N_49243,N_49244,N_49245,N_49246,N_49247,N_49248,N_49249,N_49250,N_49251,N_49252,N_49253,N_49254,N_49255,N_49256,N_49257,N_49258,N_49259,N_49260,N_49261,N_49262,N_49263,N_49264,N_49265,N_49266,N_49267,N_49268,N_49269,N_49270,N_49271,N_49272,N_49273,N_49274,N_49275,N_49276,N_49277,N_49278,N_49279,N_49280,N_49281,N_49282,N_49283,N_49284,N_49285,N_49286,N_49287,N_49288,N_49289,N_49290,N_49291,N_49292,N_49293,N_49294,N_49295,N_49296,N_49297,N_49298,N_49299,N_49300,N_49301,N_49302,N_49303,N_49304,N_49305,N_49306,N_49307,N_49308,N_49309,N_49310,N_49311,N_49312,N_49313,N_49314,N_49315,N_49316,N_49317,N_49318,N_49319,N_49320,N_49321,N_49322,N_49323,N_49324,N_49325,N_49326,N_49327,N_49328,N_49329,N_49330,N_49331,N_49332,N_49333,N_49334,N_49335,N_49336,N_49337,N_49338,N_49339,N_49340,N_49341,N_49342,N_49343,N_49344,N_49345,N_49346,N_49347,N_49348,N_49349,N_49350,N_49351,N_49352,N_49353,N_49354,N_49355,N_49356,N_49357,N_49358,N_49359,N_49360,N_49361,N_49362,N_49363,N_49364,N_49365,N_49366,N_49367,N_49368,N_49369,N_49370,N_49371,N_49372,N_49373,N_49374,N_49375,N_49376,N_49377,N_49378,N_49379,N_49380,N_49381,N_49382,N_49383,N_49384,N_49385,N_49386,N_49387,N_49388,N_49389,N_49390,N_49391,N_49392,N_49393,N_49394,N_49395,N_49396,N_49397,N_49398,N_49399,N_49400,N_49401,N_49402,N_49403,N_49404,N_49405,N_49406,N_49407,N_49408,N_49409,N_49410,N_49411,N_49412,N_49413,N_49414,N_49415,N_49416,N_49417,N_49418,N_49419,N_49420,N_49421,N_49422,N_49423,N_49424,N_49425,N_49426,N_49427,N_49428,N_49429,N_49430,N_49431,N_49432,N_49433,N_49434,N_49435,N_49436,N_49437,N_49438,N_49439,N_49440,N_49441,N_49442,N_49443,N_49444,N_49445,N_49446,N_49447,N_49448,N_49449,N_49450,N_49451,N_49452,N_49453,N_49454,N_49455,N_49456,N_49457,N_49458,N_49459,N_49460,N_49461,N_49462,N_49463,N_49464,N_49465,N_49466,N_49467,N_49468,N_49469,N_49470,N_49471,N_49472,N_49473,N_49474,N_49475,N_49476,N_49477,N_49478,N_49479,N_49480,N_49481,N_49482,N_49483,N_49484,N_49485,N_49486,N_49487,N_49488,N_49489,N_49490,N_49491,N_49492,N_49493,N_49494,N_49495,N_49496,N_49497,N_49498,N_49499,N_49500,N_49501,N_49502,N_49503,N_49504,N_49505,N_49506,N_49507,N_49508,N_49509,N_49510,N_49511,N_49512,N_49513,N_49514,N_49515,N_49516,N_49517,N_49518,N_49519,N_49520,N_49521,N_49522,N_49523,N_49524,N_49525,N_49526,N_49527,N_49528,N_49529,N_49530,N_49531,N_49532,N_49533,N_49534,N_49535,N_49536,N_49537,N_49538,N_49539,N_49540,N_49541,N_49542,N_49543,N_49544,N_49545,N_49546,N_49547,N_49548,N_49549,N_49550,N_49551,N_49552,N_49553,N_49554,N_49555,N_49556,N_49557,N_49558,N_49559,N_49560,N_49561,N_49562,N_49563,N_49564,N_49565,N_49566,N_49567,N_49568,N_49569,N_49570,N_49571,N_49572,N_49573,N_49574,N_49575,N_49576,N_49577,N_49578,N_49579,N_49580,N_49581,N_49582,N_49583,N_49584,N_49585,N_49586,N_49587,N_49588,N_49589,N_49590,N_49591,N_49592,N_49593,N_49594,N_49595,N_49596,N_49597,N_49598,N_49599,N_49600,N_49601,N_49602,N_49603,N_49604,N_49605,N_49606,N_49607,N_49608,N_49609,N_49610,N_49611,N_49612,N_49613,N_49614,N_49615,N_49616,N_49617,N_49618,N_49619,N_49620,N_49621,N_49622,N_49623,N_49624,N_49625,N_49626,N_49627,N_49628,N_49629,N_49630,N_49631,N_49632,N_49633,N_49634,N_49635,N_49636,N_49637,N_49638,N_49639,N_49640,N_49641,N_49642,N_49643,N_49644,N_49645,N_49646,N_49647,N_49648,N_49649,N_49650,N_49651,N_49652,N_49653,N_49654,N_49655,N_49656,N_49657,N_49658,N_49659,N_49660,N_49661,N_49662,N_49663,N_49664,N_49665,N_49666,N_49667,N_49668,N_49669,N_49670,N_49671,N_49672,N_49673,N_49674,N_49675,N_49676,N_49677,N_49678,N_49679,N_49680,N_49681,N_49682,N_49683,N_49684,N_49685,N_49686,N_49687,N_49688,N_49689,N_49690,N_49691,N_49692,N_49693,N_49694,N_49695,N_49696,N_49697,N_49698,N_49699,N_49700,N_49701,N_49702,N_49703,N_49704,N_49705,N_49706,N_49707,N_49708,N_49709,N_49710,N_49711,N_49712,N_49713,N_49714,N_49715,N_49716,N_49717,N_49718,N_49719,N_49720,N_49721,N_49722,N_49723,N_49724,N_49725,N_49726,N_49727,N_49728,N_49729,N_49730,N_49731,N_49732,N_49733,N_49734,N_49735,N_49736,N_49737,N_49738,N_49739,N_49740,N_49741,N_49742,N_49743,N_49744,N_49745,N_49746,N_49747,N_49748,N_49749,N_49750,N_49751,N_49752,N_49753,N_49754,N_49755,N_49756,N_49757,N_49758,N_49759,N_49760,N_49761,N_49762,N_49763,N_49764,N_49765,N_49766,N_49767,N_49768,N_49769,N_49770,N_49771,N_49772,N_49773,N_49774,N_49775,N_49776,N_49777,N_49778,N_49779,N_49780,N_49781,N_49782,N_49783,N_49784,N_49785,N_49786,N_49787,N_49788,N_49789,N_49790,N_49791,N_49792,N_49793,N_49794,N_49795,N_49796,N_49797,N_49798,N_49799,N_49800,N_49801,N_49802,N_49803,N_49804,N_49805,N_49806,N_49807,N_49808,N_49809,N_49810,N_49811,N_49812,N_49813,N_49814,N_49815,N_49816,N_49817,N_49818,N_49819,N_49820,N_49821,N_49822,N_49823,N_49824,N_49825,N_49826,N_49827,N_49828,N_49829,N_49830,N_49831,N_49832,N_49833,N_49834,N_49835,N_49836,N_49837,N_49838,N_49839,N_49840,N_49841,N_49842,N_49843,N_49844,N_49845,N_49846,N_49847,N_49848,N_49849,N_49850,N_49851,N_49852,N_49853,N_49854,N_49855,N_49856,N_49857,N_49858,N_49859,N_49860,N_49861,N_49862,N_49863,N_49864,N_49865,N_49866,N_49867,N_49868,N_49869,N_49870,N_49871,N_49872,N_49873,N_49874,N_49875,N_49876,N_49877,N_49878,N_49879,N_49880,N_49881,N_49882,N_49883,N_49884,N_49885,N_49886,N_49887,N_49888,N_49889,N_49890,N_49891,N_49892,N_49893,N_49894,N_49895,N_49896,N_49897,N_49898,N_49899,N_49900,N_49901,N_49902,N_49903,N_49904,N_49905,N_49906,N_49907,N_49908,N_49909,N_49910,N_49911,N_49912,N_49913,N_49914,N_49915,N_49916,N_49917,N_49918,N_49919,N_49920,N_49921,N_49922,N_49923,N_49924,N_49925,N_49926,N_49927,N_49928,N_49929,N_49930,N_49931,N_49932,N_49933,N_49934,N_49935,N_49936,N_49937,N_49938,N_49939,N_49940,N_49941,N_49942,N_49943,N_49944,N_49945,N_49946,N_49947,N_49948,N_49949,N_49950,N_49951,N_49952,N_49953,N_49954,N_49955,N_49956,N_49957,N_49958,N_49959,N_49960,N_49961,N_49962,N_49963,N_49964,N_49965,N_49966,N_49967,N_49968,N_49969,N_49970,N_49971,N_49972,N_49973,N_49974,N_49975,N_49976,N_49977,N_49978,N_49979,N_49980,N_49981,N_49982,N_49983,N_49984,N_49985,N_49986,N_49987,N_49988,N_49989,N_49990,N_49991,N_49992,N_49993,N_49994,N_49995,N_49996,N_49997,N_49998,N_49999;
nor U0 (N_0,In_3520,In_961);
or U1 (N_1,In_4661,In_3662);
and U2 (N_2,In_2220,In_3333);
nand U3 (N_3,In_4673,In_1914);
and U4 (N_4,In_3618,In_1180);
nor U5 (N_5,In_3714,In_3381);
or U6 (N_6,In_1931,In_1772);
nand U7 (N_7,In_2112,In_2120);
nand U8 (N_8,In_4739,In_792);
xor U9 (N_9,In_2796,In_3179);
xnor U10 (N_10,In_625,In_3152);
or U11 (N_11,In_2318,In_3776);
nand U12 (N_12,In_1576,In_271);
or U13 (N_13,In_3752,In_1184);
nor U14 (N_14,In_2821,In_2744);
nand U15 (N_15,In_3822,In_3149);
nor U16 (N_16,In_859,In_1498);
xnor U17 (N_17,In_2986,In_4019);
nor U18 (N_18,In_1535,In_1913);
and U19 (N_19,In_919,In_483);
nand U20 (N_20,In_198,In_4885);
nand U21 (N_21,In_3316,In_4964);
nand U22 (N_22,In_2185,In_1432);
xnor U23 (N_23,In_2941,In_3873);
or U24 (N_24,In_2763,In_1816);
nor U25 (N_25,In_1136,In_1400);
xnor U26 (N_26,In_2865,In_1072);
xnor U27 (N_27,In_1274,In_1522);
nor U28 (N_28,In_2543,In_2514);
xor U29 (N_29,In_2042,In_1443);
xnor U30 (N_30,In_851,In_690);
nor U31 (N_31,In_2663,In_1842);
nor U32 (N_32,In_1450,In_3175);
and U33 (N_33,In_3246,In_1199);
nor U34 (N_34,In_2657,In_2231);
nor U35 (N_35,In_127,In_2127);
and U36 (N_36,In_4333,In_2939);
or U37 (N_37,In_292,In_2554);
xor U38 (N_38,In_1241,In_2907);
xor U39 (N_39,In_2882,In_4513);
nor U40 (N_40,In_3590,In_1797);
nor U41 (N_41,In_4801,In_4980);
nor U42 (N_42,In_1336,In_440);
or U43 (N_43,In_313,In_241);
and U44 (N_44,In_1925,In_2337);
and U45 (N_45,In_3047,In_144);
and U46 (N_46,In_1082,In_1561);
or U47 (N_47,In_1848,In_2178);
nand U48 (N_48,In_4957,In_3664);
nor U49 (N_49,In_1837,In_2974);
nor U50 (N_50,In_3761,In_1203);
or U51 (N_51,In_2587,In_2955);
xnor U52 (N_52,In_53,In_1322);
xor U53 (N_53,In_881,In_935);
nand U54 (N_54,In_4071,In_2733);
xnor U55 (N_55,In_1048,In_2038);
nand U56 (N_56,In_2141,In_4698);
or U57 (N_57,In_1442,In_3842);
and U58 (N_58,In_335,In_837);
nor U59 (N_59,In_4669,In_3362);
xnor U60 (N_60,In_2515,In_4566);
xnor U61 (N_61,In_3661,In_944);
nor U62 (N_62,In_1373,In_4114);
and U63 (N_63,In_126,In_2299);
nand U64 (N_64,In_2945,In_2064);
nand U65 (N_65,In_2177,In_2491);
or U66 (N_66,In_3021,In_2192);
and U67 (N_67,In_2791,In_1210);
nor U68 (N_68,In_1883,In_2146);
and U69 (N_69,In_1889,In_2991);
xnor U70 (N_70,In_1305,In_3588);
and U71 (N_71,In_3726,In_4671);
xor U72 (N_72,In_4568,In_3566);
nor U73 (N_73,In_4914,In_3305);
xnor U74 (N_74,In_1100,In_3787);
or U75 (N_75,In_1891,In_1167);
nor U76 (N_76,In_3373,In_820);
xnor U77 (N_77,In_1987,In_906);
nor U78 (N_78,In_2467,In_2397);
nand U79 (N_79,In_988,In_3355);
and U80 (N_80,In_4195,In_3608);
or U81 (N_81,In_3137,In_4381);
nor U82 (N_82,In_3370,In_392);
nor U83 (N_83,In_4633,In_1585);
or U84 (N_84,In_4391,In_3285);
and U85 (N_85,In_4982,In_2903);
and U86 (N_86,In_2808,In_4276);
and U87 (N_87,In_3414,In_265);
xnor U88 (N_88,In_3976,In_3670);
nand U89 (N_89,In_4696,In_3484);
and U90 (N_90,In_2875,In_1852);
nand U91 (N_91,In_336,In_1938);
or U92 (N_92,In_1412,In_4238);
nor U93 (N_93,In_2540,In_3867);
or U94 (N_94,In_2445,In_1557);
xnor U95 (N_95,In_3091,In_1032);
nor U96 (N_96,In_3014,In_226);
nand U97 (N_97,In_1052,In_2693);
nand U98 (N_98,In_1533,In_773);
nor U99 (N_99,In_1586,In_393);
or U100 (N_100,In_700,In_4394);
nor U101 (N_101,In_542,In_1517);
and U102 (N_102,In_3613,In_1558);
xnor U103 (N_103,In_2207,In_3206);
xor U104 (N_104,In_3811,In_4003);
or U105 (N_105,In_2929,In_4967);
xnor U106 (N_106,In_4679,In_2608);
nand U107 (N_107,In_4053,In_1009);
xnor U108 (N_108,In_2825,In_3708);
nor U109 (N_109,In_2876,In_2473);
xor U110 (N_110,In_4354,In_1768);
and U111 (N_111,In_887,In_959);
xor U112 (N_112,In_1428,In_808);
nand U113 (N_113,In_4854,In_1666);
nand U114 (N_114,In_4951,In_2970);
and U115 (N_115,In_3509,In_4931);
nor U116 (N_116,In_4873,In_3090);
or U117 (N_117,In_1829,In_1968);
or U118 (N_118,In_4628,In_4449);
nand U119 (N_119,In_4152,In_2131);
and U120 (N_120,In_4653,In_1149);
nand U121 (N_121,In_369,In_531);
nand U122 (N_122,In_3512,In_499);
and U123 (N_123,In_2352,In_839);
or U124 (N_124,In_2123,In_3095);
and U125 (N_125,In_1355,In_3154);
or U126 (N_126,In_105,In_1446);
nand U127 (N_127,In_3301,In_3382);
or U128 (N_128,In_1876,In_4553);
xor U129 (N_129,In_234,In_4907);
xor U130 (N_130,In_4487,In_3092);
nor U131 (N_131,In_2928,In_2132);
or U132 (N_132,In_1537,In_39);
nand U133 (N_133,In_728,In_4488);
xor U134 (N_134,In_3022,In_842);
xnor U135 (N_135,In_1740,In_2534);
nand U136 (N_136,In_2464,In_357);
and U137 (N_137,In_4091,In_4672);
xor U138 (N_138,In_3671,In_976);
nand U139 (N_139,In_498,In_2920);
and U140 (N_140,In_1865,In_178);
nor U141 (N_141,In_3232,In_449);
nand U142 (N_142,In_4561,In_966);
nor U143 (N_143,In_4693,In_2469);
or U144 (N_144,In_2351,In_3839);
or U145 (N_145,In_3797,In_4230);
xor U146 (N_146,In_493,In_2148);
nor U147 (N_147,In_2408,In_4100);
nand U148 (N_148,In_3307,In_2427);
nor U149 (N_149,In_4159,In_4384);
nand U150 (N_150,In_2443,In_1980);
or U151 (N_151,In_140,In_2359);
or U152 (N_152,In_2930,In_1097);
xnor U153 (N_153,In_953,In_1732);
nand U154 (N_154,In_1062,In_3527);
nand U155 (N_155,In_1946,In_2829);
nor U156 (N_156,In_3383,In_4532);
nand U157 (N_157,In_1050,In_1109);
and U158 (N_158,In_2577,In_4969);
nand U159 (N_159,In_3279,In_4606);
nor U160 (N_160,In_2936,In_1781);
xnor U161 (N_161,In_2694,In_1658);
or U162 (N_162,In_379,In_2827);
and U163 (N_163,In_4917,In_3689);
nand U164 (N_164,In_4796,In_3835);
nor U165 (N_165,In_218,In_322);
nand U166 (N_166,In_2350,In_2251);
nand U167 (N_167,In_1362,In_4906);
xnor U168 (N_168,In_4389,In_3485);
xor U169 (N_169,In_642,In_4594);
xor U170 (N_170,In_2539,In_4301);
and U171 (N_171,In_1279,In_1008);
and U172 (N_172,In_2788,In_56);
nand U173 (N_173,In_1552,In_4234);
xnor U174 (N_174,In_309,In_1312);
nand U175 (N_175,In_3412,In_3293);
xor U176 (N_176,In_4239,In_1381);
xor U177 (N_177,In_239,In_2755);
and U178 (N_178,In_3200,In_1299);
or U179 (N_179,In_4625,In_529);
nor U180 (N_180,In_1012,In_3390);
nor U181 (N_181,In_4259,In_356);
nand U182 (N_182,In_3648,In_48);
and U183 (N_183,In_1483,In_1663);
and U184 (N_184,In_2592,In_1458);
or U185 (N_185,In_1773,In_1832);
and U186 (N_186,In_402,In_4039);
xnor U187 (N_187,In_478,In_515);
xnor U188 (N_188,In_4421,In_785);
nor U189 (N_189,In_2306,In_689);
and U190 (N_190,In_654,In_4962);
nand U191 (N_191,In_3789,In_2668);
nand U192 (N_192,In_1361,In_4450);
or U193 (N_193,In_1118,In_3304);
nand U194 (N_194,In_3473,In_2360);
nand U195 (N_195,In_2302,In_2949);
nor U196 (N_196,In_4476,In_4134);
and U197 (N_197,In_1667,In_1472);
nand U198 (N_198,In_806,In_4406);
and U199 (N_199,In_3430,In_1744);
or U200 (N_200,In_1023,In_4210);
and U201 (N_201,In_4346,In_3134);
xnor U202 (N_202,In_2396,In_1391);
nor U203 (N_203,In_852,In_213);
nor U204 (N_204,In_4383,In_2583);
xnor U205 (N_205,In_2642,In_1642);
and U206 (N_206,In_4156,In_3616);
nor U207 (N_207,In_1749,In_103);
nand U208 (N_208,In_3562,In_1467);
and U209 (N_209,In_420,In_399);
nand U210 (N_210,In_1031,In_921);
and U211 (N_211,In_2794,In_1250);
and U212 (N_212,In_1792,In_3564);
nor U213 (N_213,In_1952,In_2600);
nand U214 (N_214,In_4556,In_151);
nor U215 (N_215,In_1195,In_3108);
xor U216 (N_216,In_4541,In_90);
or U217 (N_217,In_1359,In_25);
nand U218 (N_218,In_518,In_4014);
nor U219 (N_219,In_3039,In_1831);
xnor U220 (N_220,In_693,In_3238);
and U221 (N_221,In_4533,In_805);
xor U222 (N_222,In_3457,In_854);
nand U223 (N_223,In_3173,In_27);
and U224 (N_224,In_1699,In_2115);
nand U225 (N_225,In_1090,In_4648);
xor U226 (N_226,In_962,In_1810);
nand U227 (N_227,In_2206,In_4147);
nand U228 (N_228,In_4143,In_4680);
nand U229 (N_229,In_1027,In_3208);
and U230 (N_230,In_391,In_681);
nand U231 (N_231,In_4438,In_2954);
xnor U232 (N_232,In_3893,In_4252);
nand U233 (N_233,In_3494,In_4932);
nor U234 (N_234,In_3303,In_4930);
nor U235 (N_235,In_2226,In_4960);
or U236 (N_236,In_3313,In_1588);
nor U237 (N_237,In_1545,In_1329);
or U238 (N_238,In_3821,In_445);
xor U239 (N_239,In_337,In_992);
xnor U240 (N_240,In_4954,In_555);
and U241 (N_241,In_2578,In_1890);
xor U242 (N_242,In_2637,In_3848);
and U243 (N_243,In_4246,In_2559);
or U244 (N_244,In_904,In_2003);
nor U245 (N_245,In_658,In_4756);
and U246 (N_246,In_4049,In_1998);
xor U247 (N_247,In_3254,In_3031);
nor U248 (N_248,In_3621,In_1054);
nand U249 (N_249,In_2338,In_4617);
nand U250 (N_250,In_164,In_2304);
nor U251 (N_251,In_2701,In_118);
or U252 (N_252,In_1775,In_2997);
xor U253 (N_253,In_960,In_2118);
and U254 (N_254,In_3034,N_11);
nand U255 (N_255,In_2274,In_2116);
nand U256 (N_256,In_3569,In_2398);
or U257 (N_257,In_2676,In_1431);
or U258 (N_258,In_3968,In_4206);
or U259 (N_259,In_2447,In_4085);
xor U260 (N_260,In_4111,In_3701);
nand U261 (N_261,In_3944,In_4292);
and U262 (N_262,In_3500,In_1785);
nand U263 (N_263,In_3683,N_97);
or U264 (N_264,In_1334,In_1904);
nor U265 (N_265,In_568,In_2728);
xnor U266 (N_266,N_52,In_2914);
or U267 (N_267,In_4794,In_4697);
nand U268 (N_268,In_3183,In_4463);
xnor U269 (N_269,In_2312,In_3429);
and U270 (N_270,In_11,In_3191);
and U271 (N_271,In_3543,In_249);
or U272 (N_272,In_2376,In_4274);
or U273 (N_273,In_1673,In_2414);
and U274 (N_274,In_2653,In_4121);
or U275 (N_275,In_2004,In_1709);
and U276 (N_276,In_4642,In_422);
nand U277 (N_277,In_1736,In_4538);
xor U278 (N_278,In_2591,In_4067);
and U279 (N_279,In_4754,In_2493);
xnor U280 (N_280,In_632,In_129);
and U281 (N_281,In_2697,In_964);
nand U282 (N_282,In_4789,In_169);
xor U283 (N_283,In_1132,In_3239);
nand U284 (N_284,In_4768,In_1901);
xnor U285 (N_285,In_7,In_4379);
and U286 (N_286,In_1360,In_344);
nor U287 (N_287,In_2501,In_3326);
and U288 (N_288,In_3946,N_116);
xnor U289 (N_289,In_1873,In_2859);
and U290 (N_290,In_4593,In_931);
or U291 (N_291,In_3369,In_908);
nor U292 (N_292,In_1248,N_30);
and U293 (N_293,In_2237,In_1249);
and U294 (N_294,In_3779,N_106);
and U295 (N_295,In_4780,In_4430);
and U296 (N_296,In_4809,In_1000);
or U297 (N_297,In_3529,In_77);
nor U298 (N_298,In_827,In_2969);
nor U299 (N_299,In_2606,In_3446);
and U300 (N_300,In_3748,In_3918);
or U301 (N_301,In_4686,In_710);
and U302 (N_302,N_125,In_1930);
nor U303 (N_303,In_4665,In_1011);
and U304 (N_304,In_4992,In_3450);
and U305 (N_305,In_3989,N_220);
xor U306 (N_306,In_3231,In_2331);
nand U307 (N_307,In_3780,In_2593);
or U308 (N_308,In_2589,In_4824);
xnor U309 (N_309,In_831,In_2441);
nand U310 (N_310,In_4848,In_1003);
nand U311 (N_311,In_3653,In_4150);
xnor U312 (N_312,In_4355,In_1553);
xnor U313 (N_313,In_1317,In_4734);
and U314 (N_314,In_2734,In_3458);
xor U315 (N_315,In_2387,In_1941);
or U316 (N_316,In_210,In_2561);
and U317 (N_317,In_3974,In_4802);
nand U318 (N_318,In_2552,In_4763);
and U319 (N_319,In_2639,In_1337);
or U320 (N_320,In_41,In_4138);
nor U321 (N_321,In_4903,In_1710);
xor U322 (N_322,In_1018,In_3120);
nand U323 (N_323,In_4280,In_4572);
nand U324 (N_324,In_2266,In_1019);
nor U325 (N_325,In_2328,In_567);
xnor U326 (N_326,In_3029,In_4339);
nor U327 (N_327,In_54,In_1654);
or U328 (N_328,In_2544,In_2332);
xnor U329 (N_329,In_2363,In_4546);
and U330 (N_330,In_4144,In_4877);
or U331 (N_331,In_4523,In_116);
and U332 (N_332,In_3991,In_4161);
nor U333 (N_333,In_2841,In_65);
or U334 (N_334,In_3539,In_1225);
or U335 (N_335,N_72,In_1789);
nand U336 (N_336,In_171,In_640);
nand U337 (N_337,In_125,In_3573);
nor U338 (N_338,In_1200,In_4843);
nor U339 (N_339,In_4001,In_3812);
xor U340 (N_340,In_1911,In_3234);
and U341 (N_341,N_154,In_366);
nor U342 (N_342,In_1310,In_1327);
and U343 (N_343,In_2495,In_3363);
and U344 (N_344,In_1242,In_3150);
xor U345 (N_345,In_2671,In_1193);
nor U346 (N_346,In_1067,In_4677);
nand U347 (N_347,In_2373,In_3749);
xnor U348 (N_348,In_2486,In_4704);
xnor U349 (N_349,In_3262,In_1518);
nor U350 (N_350,In_3640,In_3853);
and U351 (N_351,In_4823,In_2981);
and U352 (N_352,In_521,N_62);
and U353 (N_353,In_2310,In_29);
nand U354 (N_354,In_2984,In_2095);
or U355 (N_355,In_3549,In_3256);
nand U356 (N_356,In_1176,In_3441);
nor U357 (N_357,In_2035,In_4022);
xor U358 (N_358,In_346,In_2611);
nor U359 (N_359,In_787,In_136);
and U360 (N_360,In_1997,In_922);
nand U361 (N_361,In_3139,In_4821);
nand U362 (N_362,In_1079,In_1655);
nor U363 (N_363,In_4602,In_2910);
nand U364 (N_364,N_138,In_1961);
or U365 (N_365,In_3583,In_2630);
nor U366 (N_366,In_184,In_3763);
xor U367 (N_367,In_1323,In_1041);
nor U368 (N_368,In_4128,In_1216);
nor U369 (N_369,In_768,In_4583);
and U370 (N_370,In_3734,In_4424);
xor U371 (N_371,In_2636,In_603);
and U372 (N_372,In_2564,In_3985);
or U373 (N_373,In_3386,In_629);
nor U374 (N_374,In_2287,In_3829);
nor U375 (N_375,In_2169,In_4835);
xnor U376 (N_376,In_2111,In_3766);
nor U377 (N_377,In_2366,In_3535);
or U378 (N_378,In_713,In_3937);
and U379 (N_379,In_2725,In_2348);
or U380 (N_380,In_3243,In_2656);
and U381 (N_381,In_3907,In_2635);
and U382 (N_382,In_4284,In_2647);
xor U383 (N_383,In_3586,In_464);
and U384 (N_384,In_2390,In_388);
xor U385 (N_385,In_3795,In_2176);
nand U386 (N_386,In_3168,In_1053);
and U387 (N_387,In_3508,In_2194);
nand U388 (N_388,In_2891,In_186);
and U389 (N_389,In_3060,In_3207);
and U390 (N_390,In_443,In_3693);
xnor U391 (N_391,In_4330,In_3275);
or U392 (N_392,In_120,In_682);
nor U393 (N_393,N_126,In_2382);
nand U394 (N_394,In_4678,In_91);
and U395 (N_395,In_4211,In_3028);
nor U396 (N_396,In_3808,In_3665);
nor U397 (N_397,In_352,N_183);
xnor U398 (N_398,In_832,In_349);
and U399 (N_399,In_256,In_733);
and U400 (N_400,In_1659,In_101);
xor U401 (N_401,In_4242,In_3128);
or U402 (N_402,In_2124,In_162);
nor U403 (N_403,In_3916,In_2844);
xnor U404 (N_404,In_3525,In_311);
nor U405 (N_405,In_3841,In_1021);
or U406 (N_406,In_3467,In_3404);
nor U407 (N_407,In_4760,In_2279);
or U408 (N_408,In_2105,In_1798);
xor U409 (N_409,In_511,In_2025);
or U410 (N_410,In_1653,In_1543);
and U411 (N_411,In_3147,In_638);
xnor U412 (N_412,In_2677,In_1212);
or U413 (N_413,In_1218,In_4485);
and U414 (N_414,In_4770,In_1183);
xor U415 (N_415,In_2460,N_48);
and U416 (N_416,In_390,N_142);
xor U417 (N_417,In_3744,N_56);
and U418 (N_418,In_3133,In_537);
nor U419 (N_419,In_4431,In_220);
nor U420 (N_420,In_982,In_589);
nand U421 (N_421,N_171,In_141);
xor U422 (N_422,In_3926,In_751);
and U423 (N_423,In_4462,In_43);
nor U424 (N_424,In_4325,In_2524);
nor U425 (N_425,In_4953,In_2235);
xnor U426 (N_426,In_1614,In_2670);
xnor U427 (N_427,In_679,In_2159);
nor U428 (N_428,In_4816,In_2339);
xor U429 (N_429,In_3559,In_3614);
nand U430 (N_430,In_2193,In_4889);
nand U431 (N_431,In_2977,In_3610);
nor U432 (N_432,In_2150,In_2904);
and U433 (N_433,In_1959,N_15);
nand U434 (N_434,In_4574,In_4664);
nor U435 (N_435,In_419,In_1888);
xnor U436 (N_436,In_4190,In_691);
xnor U437 (N_437,In_4622,In_1129);
or U438 (N_438,In_4882,In_4318);
nor U439 (N_439,In_1524,In_1578);
or U440 (N_440,In_1903,In_4486);
nand U441 (N_441,In_2980,In_2823);
nor U442 (N_442,In_519,N_96);
xnor U443 (N_443,In_1684,In_3016);
or U444 (N_444,In_152,In_3423);
nor U445 (N_445,In_3792,In_639);
nor U446 (N_446,In_4308,In_4392);
xor U447 (N_447,In_745,In_4737);
nor U448 (N_448,In_1825,In_2164);
or U449 (N_449,In_2240,In_3477);
or U450 (N_450,In_3984,In_1962);
and U451 (N_451,In_3377,In_585);
xnor U452 (N_452,In_4342,In_766);
nand U453 (N_453,In_2502,In_4312);
xnor U454 (N_454,In_4051,In_4724);
nand U455 (N_455,In_4390,N_225);
or U456 (N_456,In_410,In_2288);
and U457 (N_457,In_2284,In_3089);
or U458 (N_458,In_2817,In_1396);
nand U459 (N_459,In_1237,In_1429);
nor U460 (N_460,In_4510,In_4576);
nor U461 (N_461,In_3129,In_2950);
or U462 (N_462,In_4235,In_759);
nor U463 (N_463,In_3594,In_5);
nor U464 (N_464,In_3690,In_2405);
nor U465 (N_465,In_3105,In_3691);
xor U466 (N_466,In_3315,In_3901);
nor U467 (N_467,In_572,In_2076);
nand U468 (N_468,In_1301,In_4459);
or U469 (N_469,In_2742,In_3958);
xor U470 (N_470,N_35,In_4560);
or U471 (N_471,In_888,In_930);
and U472 (N_472,In_4637,In_958);
xor U473 (N_473,In_4413,In_4109);
and U474 (N_474,In_3177,In_2293);
or U475 (N_475,In_3519,In_1680);
xnor U476 (N_476,In_374,In_3558);
nand U477 (N_477,In_1628,In_4225);
xor U478 (N_478,In_2110,In_462);
nor U479 (N_479,In_1868,In_2581);
and U480 (N_480,In_4611,In_2411);
and U481 (N_481,In_2437,In_4047);
and U482 (N_482,In_1126,In_3913);
and U483 (N_483,In_747,In_406);
and U484 (N_484,In_2901,In_4006);
xnor U485 (N_485,In_2511,In_1110);
nand U486 (N_486,In_45,In_1624);
nand U487 (N_487,N_179,In_199);
nor U488 (N_488,In_50,In_4295);
and U489 (N_489,In_1939,In_3263);
xnor U490 (N_490,In_4831,N_43);
nand U491 (N_491,In_783,In_1729);
or U492 (N_492,In_2819,In_873);
xnor U493 (N_493,In_3654,In_3827);
and U494 (N_494,In_2919,N_94);
nor U495 (N_495,In_1609,In_3327);
xor U496 (N_496,In_2440,N_23);
xnor U497 (N_497,In_3522,In_1820);
or U498 (N_498,In_4160,In_2199);
or U499 (N_499,In_4057,In_2049);
and U500 (N_500,N_120,In_3190);
nand U501 (N_501,In_4101,In_4554);
nand U502 (N_502,In_243,In_2391);
nand U503 (N_503,In_4790,In_361);
nand U504 (N_504,In_878,In_615);
xnor U505 (N_505,In_1945,In_28);
xnor U506 (N_506,In_4779,In_1229);
nand U507 (N_507,In_253,In_4371);
nand U508 (N_508,In_4961,In_4856);
nor U509 (N_509,In_951,In_2031);
xnor U510 (N_510,In_3557,In_3528);
or U511 (N_511,In_4456,In_1783);
xnor U512 (N_512,In_2263,In_1185);
xnor U513 (N_513,In_1627,N_343);
and U514 (N_514,In_4551,In_216);
nand U515 (N_515,In_646,In_749);
nand U516 (N_516,In_1881,N_166);
nor U517 (N_517,In_2669,In_3140);
and U518 (N_518,N_332,In_4812);
xor U519 (N_519,In_3943,In_1763);
xnor U520 (N_520,In_861,In_350);
nor U521 (N_521,In_2354,In_4194);
nor U522 (N_522,In_3425,In_3894);
and U523 (N_523,N_438,In_1920);
nor U524 (N_524,In_2080,In_1051);
and U525 (N_525,In_3637,In_2720);
and U526 (N_526,In_3281,In_671);
nor U527 (N_527,In_3837,N_204);
nor U528 (N_528,In_4249,In_2062);
nor U529 (N_529,In_696,In_2685);
and U530 (N_530,In_2995,In_3550);
or U531 (N_531,In_2261,In_3006);
or U532 (N_532,In_879,In_1374);
nand U533 (N_533,N_460,In_3591);
xor U534 (N_534,In_4189,In_2547);
xor U535 (N_535,In_1343,In_1917);
or U536 (N_536,In_1092,In_2758);
nor U537 (N_537,In_2322,In_994);
or U538 (N_538,In_1625,In_2043);
xnor U539 (N_539,N_363,N_435);
nor U540 (N_540,In_4199,In_3925);
nor U541 (N_541,In_1502,In_4614);
nor U542 (N_542,In_2071,In_305);
or U543 (N_543,In_1127,In_3574);
nor U544 (N_544,In_4328,N_347);
and U545 (N_545,In_772,In_3202);
or U546 (N_546,In_586,In_2662);
xor U547 (N_547,In_4294,In_3674);
nand U548 (N_548,In_4626,In_4287);
nand U549 (N_549,N_447,In_2798);
xnor U550 (N_550,In_1434,In_2174);
and U551 (N_551,In_2078,N_387);
and U552 (N_552,N_370,In_4971);
nand U553 (N_553,In_1144,In_4863);
nand U554 (N_554,N_246,In_208);
nor U555 (N_555,N_362,N_151);
nor U556 (N_556,In_546,In_1022);
nor U557 (N_557,In_3554,In_3542);
nor U558 (N_558,In_4500,In_2333);
and U559 (N_559,In_817,In_2384);
xor U560 (N_560,In_1368,In_1905);
or U561 (N_561,In_2257,In_897);
and U562 (N_562,In_4915,In_4277);
nor U563 (N_563,In_486,N_104);
xor U564 (N_564,In_3334,In_3824);
xor U565 (N_565,In_360,In_993);
and U566 (N_566,In_2278,In_1158);
nand U567 (N_567,In_3681,In_3953);
nor U568 (N_568,In_2861,In_1761);
nand U569 (N_569,In_341,In_554);
or U570 (N_570,In_3831,In_989);
xnor U571 (N_571,In_4155,In_4986);
nor U572 (N_572,In_3879,In_2171);
nand U573 (N_573,In_4514,N_77);
nor U574 (N_574,In_1423,In_3949);
xnor U575 (N_575,In_252,In_3284);
nand U576 (N_576,In_1143,N_0);
nand U577 (N_577,In_2476,In_4097);
and U578 (N_578,In_3858,In_3132);
or U579 (N_579,In_266,In_675);
nor U580 (N_580,In_4911,In_3682);
xnor U581 (N_581,In_2654,N_314);
and U582 (N_582,In_4110,In_1015);
xor U583 (N_583,In_308,In_1696);
xnor U584 (N_584,In_812,In_4520);
nand U585 (N_585,In_1120,In_929);
and U586 (N_586,In_1966,In_952);
and U587 (N_587,N_492,N_87);
nor U588 (N_588,In_1856,In_0);
nand U589 (N_589,In_2029,In_807);
xnor U590 (N_590,In_3395,In_3196);
xor U591 (N_591,In_4562,In_2336);
or U592 (N_592,In_4204,In_2831);
and U593 (N_593,N_315,In_4118);
nand U594 (N_594,In_2922,In_4434);
or U595 (N_595,In_3306,In_1101);
nor U596 (N_596,In_619,In_4929);
and U597 (N_597,In_3124,In_4007);
nand U598 (N_598,In_1424,In_2168);
nand U599 (N_599,In_3052,In_4184);
and U600 (N_600,In_4426,In_2957);
and U601 (N_601,In_4508,In_4529);
and U602 (N_602,N_205,In_4869);
xnor U603 (N_603,In_2113,In_189);
or U604 (N_604,In_4319,In_161);
nor U605 (N_605,In_2528,In_36);
nor U606 (N_606,In_1847,In_4829);
or U607 (N_607,N_209,In_1860);
or U608 (N_608,In_3438,N_161);
nor U609 (N_609,In_620,In_4094);
xnor U610 (N_610,N_122,N_413);
and U611 (N_611,In_3631,In_2747);
nand U612 (N_612,In_3253,N_137);
nor U613 (N_613,In_4621,In_4183);
nor U614 (N_614,In_3950,In_3420);
or U615 (N_615,In_3264,N_1);
or U616 (N_616,In_3939,In_948);
xnor U617 (N_617,In_1232,In_4151);
and U618 (N_618,N_444,In_466);
nand U619 (N_619,In_3875,In_2752);
nor U620 (N_620,In_2316,In_4273);
nand U621 (N_621,In_4644,In_1045);
nand U622 (N_622,In_2937,In_1252);
or U623 (N_623,In_1778,In_2992);
nand U624 (N_624,In_533,In_2353);
and U625 (N_625,In_520,In_4709);
nand U626 (N_626,In_1076,In_1350);
nand U627 (N_627,In_4429,N_481);
xnor U628 (N_628,In_1995,In_617);
or U629 (N_629,In_1715,In_4985);
xnor U630 (N_630,In_4857,N_421);
nand U631 (N_631,In_2573,In_2424);
or U632 (N_632,In_1958,N_378);
and U633 (N_633,In_3040,In_1767);
and U634 (N_634,N_365,In_592);
nand U635 (N_635,N_46,In_522);
and U636 (N_636,In_3010,In_1004);
and U637 (N_637,In_439,In_995);
xor U638 (N_638,In_798,In_3389);
or U639 (N_639,In_963,In_351);
xor U640 (N_640,N_337,In_4125);
or U641 (N_641,In_3405,In_2215);
nor U642 (N_642,In_3580,In_3453);
nor U643 (N_643,In_4304,In_1949);
nand U644 (N_644,In_2622,In_3288);
xnor U645 (N_645,In_2155,In_2335);
and U646 (N_646,In_2628,In_2369);
and U647 (N_647,In_4077,In_4193);
or U648 (N_648,In_145,In_4684);
and U649 (N_649,In_1664,In_1957);
nand U650 (N_650,In_4933,In_3607);
and U651 (N_651,In_1448,In_1181);
nand U652 (N_652,N_464,In_121);
nand U653 (N_653,In_676,In_3340);
and U654 (N_654,In_469,In_2000);
nor U655 (N_655,In_2433,In_1977);
xor U656 (N_656,In_3240,In_4886);
or U657 (N_657,In_2401,In_2218);
or U658 (N_658,In_3595,N_422);
xor U659 (N_659,In_1268,In_2667);
nor U660 (N_660,In_801,In_4944);
nor U661 (N_661,In_3765,N_13);
xnor U662 (N_662,N_78,In_1927);
nor U663 (N_663,In_784,In_3647);
and U664 (N_664,In_3068,In_2840);
nand U665 (N_665,In_3345,In_2145);
xor U666 (N_666,In_4008,In_480);
xor U667 (N_667,N_71,In_2731);
and U668 (N_668,In_637,In_4437);
nor U669 (N_669,N_200,In_652);
xnor U670 (N_670,In_4176,In_3758);
nand U671 (N_671,In_4928,In_3220);
and U672 (N_672,In_877,In_4956);
or U673 (N_673,In_1178,In_3760);
nand U674 (N_674,In_261,N_448);
and U675 (N_675,In_2065,N_274);
and U676 (N_676,In_4070,N_251);
and U677 (N_677,In_576,In_4341);
xor U678 (N_678,In_3617,In_3959);
or U679 (N_679,In_3267,In_3773);
nand U680 (N_680,In_1202,In_3265);
and U681 (N_681,In_3130,In_2165);
or U682 (N_682,In_4826,In_3273);
nor U683 (N_683,In_3324,N_419);
xnor U684 (N_684,In_2687,In_814);
nand U685 (N_685,In_4396,In_4332);
nand U686 (N_686,In_1146,In_1765);
or U687 (N_687,In_1964,In_299);
nand U688 (N_688,In_1536,In_1975);
nor U689 (N_689,In_2283,In_3909);
and U690 (N_690,In_3515,In_1811);
nand U691 (N_691,In_762,In_2045);
xnor U692 (N_692,In_3990,In_1984);
and U693 (N_693,In_914,In_2403);
and U694 (N_694,In_3464,In_3437);
nand U695 (N_695,In_2484,N_95);
and U696 (N_696,In_1430,In_290);
or U697 (N_697,In_2456,In_130);
xor U698 (N_698,In_324,In_3881);
nand U699 (N_699,In_3531,N_415);
xnor U700 (N_700,In_4069,In_3365);
nor U701 (N_701,In_735,In_849);
xnor U702 (N_702,In_4226,In_3312);
or U703 (N_703,In_739,In_2979);
nor U704 (N_704,In_1963,In_3071);
xnor U705 (N_705,In_3655,In_4375);
nand U706 (N_706,In_1,N_226);
nor U707 (N_707,In_2597,N_461);
xor U708 (N_708,In_1214,In_514);
or U709 (N_709,In_2565,In_4721);
nand U710 (N_710,In_3398,In_1437);
or U711 (N_711,In_1660,N_373);
and U712 (N_712,In_2329,N_384);
or U713 (N_713,In_47,In_44);
xor U714 (N_714,In_4866,In_3767);
and U715 (N_715,In_1674,In_37);
xor U716 (N_716,In_3002,In_2345);
and U717 (N_717,In_4781,In_2399);
nand U718 (N_718,In_3735,In_137);
xnor U719 (N_719,In_3628,In_686);
and U720 (N_720,In_3249,In_2889);
and U721 (N_721,In_212,In_2782);
nor U722 (N_722,In_3245,In_3552);
nor U723 (N_723,In_221,In_501);
or U724 (N_724,In_3189,N_287);
nor U725 (N_725,In_3560,In_4918);
nor U726 (N_726,In_3545,In_1897);
nor U727 (N_727,In_598,In_332);
or U728 (N_728,In_3532,In_2344);
and U729 (N_729,In_3495,N_342);
nand U730 (N_730,N_252,In_895);
nand U731 (N_731,In_2802,In_211);
xnor U732 (N_732,In_385,In_228);
and U733 (N_733,In_3709,In_838);
and U734 (N_734,In_1565,In_204);
nand U735 (N_735,In_4592,In_1534);
nor U736 (N_736,In_3460,In_315);
xor U737 (N_737,In_3897,In_3440);
xnor U738 (N_738,In_4478,In_794);
or U739 (N_739,In_1065,In_1573);
and U740 (N_740,In_3857,In_2535);
and U741 (N_741,In_132,In_3013);
nand U742 (N_742,In_525,In_2142);
xnor U743 (N_743,N_452,In_326);
nor U744 (N_744,In_3287,In_3042);
nor U745 (N_745,In_1731,In_4037);
nor U746 (N_746,In_1967,N_453);
xor U747 (N_747,In_564,In_1728);
or U748 (N_748,In_3170,In_1113);
nor U749 (N_749,In_1509,In_3660);
nand U750 (N_750,In_485,In_1926);
nand U751 (N_751,In_1591,In_2682);
nand U752 (N_752,N_279,In_491);
nor U753 (N_753,In_4516,In_2426);
nor U754 (N_754,In_3004,N_394);
nand U755 (N_755,In_4852,In_3225);
or U756 (N_756,In_1639,In_3250);
nand U757 (N_757,In_1189,In_3826);
nor U758 (N_758,In_4528,In_4405);
xor U759 (N_759,In_1117,In_4140);
nand U760 (N_760,In_100,In_1646);
nand U761 (N_761,In_1220,In_4605);
xnor U762 (N_762,In_3018,In_594);
xnor U763 (N_763,In_1929,In_1404);
nor U764 (N_764,In_578,N_257);
and U765 (N_765,In_3818,N_515);
or U766 (N_766,In_1339,In_3435);
nand U767 (N_767,In_1239,N_7);
nand U768 (N_768,In_277,In_4367);
and U769 (N_769,In_4167,N_398);
xnor U770 (N_770,In_4464,In_4649);
nor U771 (N_771,In_1809,In_4557);
and U772 (N_772,In_4972,In_3971);
and U773 (N_773,In_2208,In_883);
and U774 (N_774,In_4454,In_3998);
xnor U775 (N_775,N_475,N_653);
and U776 (N_776,In_1338,In_4447);
and U777 (N_777,In_2298,In_2272);
nand U778 (N_778,In_3300,In_1206);
and U779 (N_779,In_2358,In_4901);
or U780 (N_780,In_2277,In_955);
or U781 (N_781,In_2976,In_4044);
xor U782 (N_782,In_3629,In_687);
nor U783 (N_783,In_1874,In_131);
xnor U784 (N_784,In_2870,In_285);
or U785 (N_785,In_111,In_2553);
xnor U786 (N_786,In_1754,N_583);
nand U787 (N_787,In_4772,N_269);
xor U788 (N_788,In_2740,In_3910);
xor U789 (N_789,N_51,In_2027);
xor U790 (N_790,In_1457,In_438);
xnor U791 (N_791,In_3427,In_1307);
nand U792 (N_792,N_410,In_3242);
nand U793 (N_793,In_2911,In_2550);
nand U794 (N_794,In_1084,N_493);
nor U795 (N_795,In_1033,In_1923);
or U796 (N_796,In_377,In_1034);
nand U797 (N_797,In_1649,In_2805);
nand U798 (N_798,In_936,In_4031);
nor U799 (N_799,In_404,In_702);
nor U800 (N_800,In_3782,In_1152);
nor U801 (N_801,In_3367,In_1858);
xor U802 (N_802,In_4804,In_3882);
nor U803 (N_803,In_4511,In_1515);
xor U804 (N_804,N_584,In_4503);
nand U805 (N_805,In_3713,N_434);
and U806 (N_806,In_282,N_480);
and U807 (N_807,In_3886,N_428);
or U808 (N_808,In_306,N_532);
or U809 (N_809,In_2993,In_4257);
or U810 (N_810,In_4616,In_1879);
or U811 (N_811,In_2204,In_584);
or U812 (N_812,In_405,In_3411);
nand U813 (N_813,In_4248,In_927);
or U814 (N_814,In_46,In_1992);
nand U815 (N_815,In_2830,In_1918);
or U816 (N_816,In_1141,In_524);
and U817 (N_817,N_353,In_1413);
and U818 (N_818,In_574,In_365);
nand U819 (N_819,In_3899,In_4567);
xor U820 (N_820,In_874,In_4136);
and U821 (N_821,In_2769,In_453);
nor U822 (N_822,In_2269,In_3584);
or U823 (N_823,In_4518,In_990);
nand U824 (N_824,In_1933,In_858);
or U825 (N_825,N_443,In_3790);
or U826 (N_826,In_765,N_284);
xnor U827 (N_827,In_853,N_417);
nor U828 (N_828,In_236,N_108);
or U829 (N_829,In_2037,In_4810);
xor U830 (N_830,In_2879,In_4207);
nand U831 (N_831,In_2030,In_1640);
and U832 (N_832,In_4731,In_3252);
or U833 (N_833,In_1880,N_683);
nand U834 (N_834,In_3278,In_3724);
nor U835 (N_835,In_4105,In_506);
or U836 (N_836,In_722,In_3399);
xor U837 (N_837,In_232,In_67);
nand U838 (N_838,In_1013,In_744);
xnor U839 (N_839,In_726,In_4416);
nor U840 (N_840,In_4496,In_2570);
xor U841 (N_841,N_712,In_4943);
and U842 (N_842,N_354,N_677);
or U843 (N_843,In_3210,In_3538);
nor U844 (N_844,In_1956,In_2856);
nand U845 (N_845,In_441,In_2483);
or U846 (N_846,In_4530,In_4834);
or U847 (N_847,In_4934,In_716);
nand U848 (N_848,In_2761,In_651);
or U849 (N_849,In_217,In_2104);
or U850 (N_850,In_3698,In_2575);
nand U851 (N_851,In_1570,In_1056);
nor U852 (N_852,In_3431,N_50);
xor U853 (N_853,In_3741,In_4475);
xor U854 (N_854,In_3221,In_259);
nand U855 (N_855,In_4937,In_3657);
nor U856 (N_856,In_4650,N_150);
xor U857 (N_857,In_3570,In_3280);
nor U858 (N_858,In_2784,In_3820);
xnor U859 (N_859,In_4278,In_58);
or U860 (N_860,In_4820,In_3504);
and U861 (N_861,In_2355,N_357);
and U862 (N_862,In_1372,In_3094);
nand U863 (N_863,In_683,In_1098);
nand U864 (N_864,In_761,In_394);
or U865 (N_865,N_404,In_1638);
or U866 (N_866,In_2324,N_153);
xnor U867 (N_867,In_4545,In_3292);
or U868 (N_868,In_1505,In_4620);
or U869 (N_869,In_42,In_2481);
nor U870 (N_870,In_4359,In_1603);
or U871 (N_871,In_4412,In_3076);
and U872 (N_872,In_389,In_730);
or U873 (N_873,N_65,In_1460);
nand U874 (N_874,N_392,In_3198);
xnor U875 (N_875,In_3546,In_1621);
and U876 (N_876,In_1251,In_3144);
xnor U877 (N_877,In_1147,In_1716);
nand U878 (N_878,In_1346,N_336);
nand U879 (N_879,In_300,In_206);
nand U880 (N_880,In_2908,N_676);
nand U881 (N_881,N_21,In_4490);
and U882 (N_882,In_1358,In_201);
nand U883 (N_883,In_1102,In_2144);
nand U884 (N_884,In_2392,In_500);
nor U885 (N_885,In_4262,In_2014);
nand U886 (N_886,In_63,In_31);
nand U887 (N_887,In_1730,N_259);
or U888 (N_888,In_4060,In_2946);
or U889 (N_889,In_4595,N_262);
or U890 (N_890,In_421,In_1342);
nor U891 (N_891,In_4850,In_2743);
and U892 (N_892,N_577,In_570);
nor U893 (N_893,In_4846,In_386);
nor U894 (N_894,N_335,In_3890);
nor U895 (N_895,In_4635,In_3219);
xor U896 (N_896,In_163,In_2947);
xor U897 (N_897,In_1213,In_1993);
xor U898 (N_898,In_2948,N_566);
nand U899 (N_899,In_811,In_4229);
or U900 (N_900,In_1161,In_753);
nor U901 (N_901,N_724,In_325);
and U902 (N_902,In_3401,In_923);
xor U903 (N_903,N_189,In_4149);
or U904 (N_904,In_1983,In_2518);
nor U905 (N_905,In_200,N_330);
nand U906 (N_906,In_2210,In_296);
nor U907 (N_907,In_3915,In_4058);
nand U908 (N_908,In_2541,In_1262);
nor U909 (N_909,In_4788,N_184);
xor U910 (N_910,In_1618,In_3117);
xnor U911 (N_911,In_1538,In_4115);
xnor U912 (N_912,In_4350,In_4963);
nand U913 (N_913,In_4723,In_3502);
nand U914 (N_914,In_636,In_2776);
xnor U915 (N_915,In_545,In_3349);
xor U916 (N_916,In_1451,In_1759);
nand U917 (N_917,In_4504,In_3409);
xnor U918 (N_918,In_2166,N_28);
nand U919 (N_919,In_3337,In_4663);
nand U920 (N_920,In_3496,In_1629);
xor U921 (N_921,In_4895,In_1854);
xor U922 (N_922,In_2809,In_1494);
nor U923 (N_923,N_124,In_4491);
nor U924 (N_924,In_2072,In_2890);
xor U925 (N_925,In_1283,In_2075);
xnor U926 (N_926,In_1676,N_309);
and U927 (N_927,In_3917,In_2780);
xor U928 (N_928,In_1574,In_3999);
xnor U929 (N_929,In_1815,In_12);
or U930 (N_930,In_415,N_497);
and U931 (N_931,In_886,In_1756);
nor U932 (N_932,In_2086,In_3107);
and U933 (N_933,In_3145,In_1454);
nor U934 (N_934,N_316,In_4517);
nor U935 (N_935,N_479,In_94);
nand U936 (N_936,In_4286,In_3181);
nor U937 (N_937,In_1791,In_23);
nor U938 (N_938,In_2163,N_738);
or U939 (N_939,In_1752,In_2666);
nor U940 (N_940,In_170,N_426);
nand U941 (N_941,In_2470,In_138);
nor U942 (N_942,In_1982,In_2417);
nand U943 (N_943,In_3571,In_1402);
or U944 (N_944,In_2107,In_4188);
nor U945 (N_945,In_1258,N_615);
or U946 (N_946,In_2866,In_4388);
or U947 (N_947,In_2201,In_4634);
and U948 (N_948,In_721,In_970);
or U949 (N_949,N_534,In_3443);
or U950 (N_950,In_1416,In_1064);
and U951 (N_951,In_734,In_1717);
and U952 (N_952,In_4191,In_4601);
and U953 (N_953,In_237,In_2551);
and U954 (N_954,In_396,N_260);
nand U955 (N_955,In_1814,In_3339);
nand U956 (N_956,In_3193,In_2343);
or U957 (N_957,In_1275,In_4708);
or U958 (N_958,In_4407,In_3578);
and U959 (N_959,In_2222,In_1397);
and U960 (N_960,In_3033,In_1315);
and U961 (N_961,In_4657,In_4442);
nand U962 (N_962,In_1297,In_1162);
nand U963 (N_963,In_3729,In_767);
nand U964 (N_964,In_3146,In_3211);
xor U965 (N_965,In_3186,In_4201);
nor U966 (N_966,In_1261,In_1077);
nand U967 (N_967,In_3491,N_61);
and U968 (N_968,In_4771,In_1972);
nand U969 (N_969,In_1843,In_2280);
nand U970 (N_970,N_14,In_4910);
xor U971 (N_971,In_2601,In_3856);
nand U972 (N_972,In_4888,N_650);
xor U973 (N_973,In_3226,In_455);
nor U974 (N_974,In_3994,In_2710);
nand U975 (N_975,N_211,In_1073);
nand U976 (N_976,In_669,In_3075);
nor U977 (N_977,In_3385,In_2393);
and U978 (N_978,In_4828,N_689);
or U979 (N_979,In_3563,In_4305);
or U980 (N_980,N_619,In_616);
nand U981 (N_981,In_4298,In_911);
nor U982 (N_982,In_1895,In_3104);
nand U983 (N_983,In_294,In_3832);
and U984 (N_984,In_3816,In_4299);
or U985 (N_985,In_1937,In_4913);
nand U986 (N_986,In_1550,In_1344);
xor U987 (N_987,N_745,In_2212);
xor U988 (N_988,In_3771,In_61);
or U989 (N_989,In_3627,In_1726);
nor U990 (N_990,N_562,In_2994);
xnor U991 (N_991,In_2327,In_3669);
and U992 (N_992,N_512,In_3379);
xor U993 (N_993,In_1779,In_3544);
xor U994 (N_994,N_367,In_2094);
nor U995 (N_995,In_3687,N_552);
xnor U996 (N_996,In_4894,N_320);
nand U997 (N_997,In_1971,In_937);
and U998 (N_998,In_2522,In_482);
or U999 (N_999,In_3479,In_3805);
nand U1000 (N_1000,In_3676,In_2878);
xor U1001 (N_1001,N_788,In_4417);
xor U1002 (N_1002,N_143,In_4582);
xnor U1003 (N_1003,In_1745,In_896);
nand U1004 (N_1004,In_998,In_92);
xnor U1005 (N_1005,In_3742,N_103);
or U1006 (N_1006,In_3017,In_2307);
nor U1007 (N_1007,N_974,N_70);
or U1008 (N_1008,N_799,In_3672);
nor U1009 (N_1009,In_3298,In_2843);
or U1010 (N_1010,In_1508,In_2932);
xnor U1011 (N_1011,In_2139,N_899);
and U1012 (N_1012,N_75,In_1341);
and U1013 (N_1013,N_668,In_436);
nand U1014 (N_1014,N_945,N_272);
and U1015 (N_1015,N_731,In_4775);
xnor U1016 (N_1016,In_4218,In_2513);
or U1017 (N_1017,In_4942,In_2059);
nor U1018 (N_1018,In_3957,In_3673);
nor U1019 (N_1019,In_2634,In_569);
nor U1020 (N_1020,In_2341,In_1406);
xnor U1021 (N_1021,In_3121,In_1747);
and U1022 (N_1022,N_952,N_655);
or U1023 (N_1023,In_1107,In_3228);
or U1024 (N_1024,In_3695,In_1155);
nor U1025 (N_1025,In_2998,In_3770);
nor U1026 (N_1026,In_606,In_2183);
nand U1027 (N_1027,In_4537,In_3077);
nor U1028 (N_1028,In_1039,In_3073);
and U1029 (N_1029,In_1115,In_2096);
or U1030 (N_1030,In_3456,In_219);
or U1031 (N_1031,In_2643,N_406);
nand U1032 (N_1032,In_1857,N_304);
and U1033 (N_1033,In_954,In_2698);
nor U1034 (N_1034,In_69,In_4726);
and U1035 (N_1035,In_1698,In_3056);
or U1036 (N_1036,In_2783,In_4168);
and U1037 (N_1037,In_866,In_235);
nand U1038 (N_1038,N_407,In_4400);
and U1039 (N_1039,In_3235,In_1735);
and U1040 (N_1040,In_2054,In_891);
nor U1041 (N_1041,In_1198,In_4870);
nor U1042 (N_1042,In_3895,In_3992);
nor U1043 (N_1043,In_1803,In_3151);
nand U1044 (N_1044,In_1234,In_2252);
or U1045 (N_1045,In_1990,In_1285);
or U1046 (N_1046,In_1112,In_4337);
or U1047 (N_1047,In_224,N_486);
or U1048 (N_1048,N_323,In_2872);
or U1049 (N_1049,In_321,In_2494);
nor U1050 (N_1050,In_4550,In_4336);
xnor U1051 (N_1051,N_462,In_1688);
nor U1052 (N_1052,In_2244,N_900);
and U1053 (N_1053,In_2549,In_4531);
nand U1054 (N_1054,In_4536,In_4187);
nand U1055 (N_1055,N_765,In_1643);
nor U1056 (N_1056,In_775,In_503);
or U1057 (N_1057,In_867,In_1380);
or U1058 (N_1058,In_1295,In_4973);
nor U1059 (N_1059,N_895,In_3813);
xnor U1060 (N_1060,N_485,In_78);
or U1061 (N_1061,In_4749,In_2289);
nor U1062 (N_1062,In_4512,In_2400);
nor U1063 (N_1063,In_2531,In_4880);
xnor U1064 (N_1064,In_3475,N_196);
nand U1065 (N_1065,In_4192,In_2044);
nand U1066 (N_1066,In_1255,In_2326);
or U1067 (N_1067,In_4148,In_1762);
nand U1068 (N_1068,In_3675,In_2726);
xor U1069 (N_1069,In_4883,In_2665);
or U1070 (N_1070,In_2746,In_4643);
nand U1071 (N_1071,In_4107,In_4351);
xor U1072 (N_1072,In_1540,N_793);
or U1073 (N_1073,N_167,In_4099);
nor U1074 (N_1074,In_4166,N_69);
and U1075 (N_1075,In_247,In_3928);
xnor U1076 (N_1076,In_370,In_3169);
or U1077 (N_1077,In_763,In_2081);
nand U1078 (N_1078,In_1567,In_4040);
and U1079 (N_1079,In_621,In_3876);
or U1080 (N_1080,In_1083,In_4844);
and U1081 (N_1081,N_820,In_712);
xor U1082 (N_1082,In_1441,In_3274);
nor U1083 (N_1083,In_4769,In_3996);
nor U1084 (N_1084,In_2015,In_3840);
and U1085 (N_1085,In_3498,In_4428);
or U1086 (N_1086,In_4623,In_2621);
or U1087 (N_1087,In_4921,In_665);
nor U1088 (N_1088,In_641,In_437);
nor U1089 (N_1089,In_2229,In_2446);
nor U1090 (N_1090,N_176,In_1108);
nor U1091 (N_1091,N_688,In_1622);
nand U1092 (N_1092,N_923,In_508);
and U1093 (N_1093,N_914,In_2197);
nand U1094 (N_1094,In_4435,N_666);
nor U1095 (N_1095,In_3103,In_3600);
and U1096 (N_1096,In_4433,N_665);
nand U1097 (N_1097,In_1131,In_3069);
and U1098 (N_1098,In_2723,In_2778);
and U1099 (N_1099,In_2051,In_934);
xor U1100 (N_1100,In_714,N_382);
nor U1101 (N_1101,In_1304,In_645);
and U1102 (N_1102,In_1392,N_381);
nand U1103 (N_1103,N_947,In_3777);
and U1104 (N_1104,In_504,In_3388);
xor U1105 (N_1105,In_2745,In_4076);
or U1106 (N_1106,In_358,N_467);
nor U1107 (N_1107,In_4372,In_1139);
nand U1108 (N_1108,In_1823,In_3164);
xnor U1109 (N_1109,N_446,In_4761);
xnor U1110 (N_1110,In_2286,In_3174);
nor U1111 (N_1111,In_3898,N_33);
or U1112 (N_1112,In_4088,In_648);
nand U1113 (N_1113,N_705,In_1318);
xnor U1114 (N_1114,In_1104,In_3592);
xor U1115 (N_1115,In_2971,In_4145);
nor U1116 (N_1116,In_3050,In_924);
nand U1117 (N_1117,In_1153,N_710);
nand U1118 (N_1118,In_4524,In_3934);
nand U1119 (N_1119,In_4055,In_3970);
xnor U1120 (N_1120,N_789,N_580);
and U1121 (N_1121,In_1804,In_2357);
nor U1122 (N_1122,In_4261,In_2063);
xnor U1123 (N_1123,In_1179,In_4178);
or U1124 (N_1124,In_1493,N_682);
and U1125 (N_1125,N_815,N_736);
nor U1126 (N_1126,N_216,N_313);
or U1127 (N_1127,In_1123,In_3666);
nand U1128 (N_1128,N_684,In_3011);
nand U1129 (N_1129,In_2455,In_1116);
xnor U1130 (N_1130,In_2005,In_2962);
nand U1131 (N_1131,In_2952,In_2787);
and U1132 (N_1132,In_3526,In_1606);
or U1133 (N_1133,In_1613,In_97);
or U1134 (N_1134,In_3116,In_2273);
nand U1135 (N_1135,In_2321,In_2036);
and U1136 (N_1136,In_2311,In_968);
nor U1137 (N_1137,In_2248,In_1645);
and U1138 (N_1138,N_960,In_362);
and U1139 (N_1139,N_38,N_996);
and U1140 (N_1140,In_2982,N_445);
nand U1141 (N_1141,In_986,In_628);
xor U1142 (N_1142,In_1291,N_891);
and U1143 (N_1143,N_291,In_1345);
xnor U1144 (N_1144,N_904,In_487);
nand U1145 (N_1145,In_432,N_889);
or U1146 (N_1146,In_3977,In_3419);
or U1147 (N_1147,In_3986,N_338);
nor U1148 (N_1148,In_950,N_159);
nor U1149 (N_1149,N_995,N_757);
or U1150 (N_1150,In_1174,In_4871);
nor U1151 (N_1151,N_100,In_4640);
or U1152 (N_1152,In_857,In_2395);
and U1153 (N_1153,In_3295,N_341);
and U1154 (N_1154,In_4005,N_199);
and U1155 (N_1155,N_412,In_3630);
or U1156 (N_1156,In_4699,N_58);
nor U1157 (N_1157,N_693,N_308);
nor U1158 (N_1158,In_1375,In_4116);
nand U1159 (N_1159,In_4687,In_4586);
and U1160 (N_1160,N_640,In_461);
xor U1161 (N_1161,In_3723,In_2610);
nor U1162 (N_1162,In_3732,In_1288);
xor U1163 (N_1163,In_4746,N_160);
or U1164 (N_1164,N_519,In_2846);
nor U1165 (N_1165,In_4169,In_4352);
or U1166 (N_1166,In_3930,N_540);
or U1167 (N_1167,N_518,N_647);
or U1168 (N_1168,In_717,N_310);
nand U1169 (N_1169,In_1581,In_3987);
and U1170 (N_1170,In_2002,In_1165);
and U1171 (N_1171,In_4066,In_4399);
and U1172 (N_1172,In_2314,N_609);
and U1173 (N_1173,In_1170,N_841);
or U1174 (N_1174,In_2349,In_4119);
and U1175 (N_1175,In_1347,In_4327);
nor U1176 (N_1176,N_661,In_4297);
xor U1177 (N_1177,In_2582,In_979);
nor U1178 (N_1178,In_2021,In_1787);
and U1179 (N_1179,In_2699,In_4890);
or U1180 (N_1180,In_2268,In_2507);
nand U1181 (N_1181,In_2842,In_4717);
nor U1182 (N_1182,N_720,In_1029);
nand U1183 (N_1183,In_269,N_823);
and U1184 (N_1184,In_3924,N_560);
xor U1185 (N_1185,In_3093,In_2368);
nand U1186 (N_1186,In_3061,N_117);
nor U1187 (N_1187,In_1328,In_926);
nand U1188 (N_1188,In_2330,In_3474);
xnor U1189 (N_1189,N_255,N_856);
nand U1190 (N_1190,In_833,In_4272);
and U1191 (N_1191,In_1046,In_1544);
and U1192 (N_1192,In_1040,In_3948);
nand U1193 (N_1193,In_663,In_2295);
xnor U1194 (N_1194,In_270,In_631);
nand U1195 (N_1195,In_1838,In_4493);
xnor U1196 (N_1196,N_824,In_1974);
or U1197 (N_1197,In_1217,In_1370);
nand U1198 (N_1198,In_2563,In_1002);
or U1199 (N_1199,In_2795,In_1559);
or U1200 (N_1200,In_1947,N_80);
nor U1201 (N_1201,In_188,In_2965);
nor U1202 (N_1202,N_520,In_3344);
and U1203 (N_1203,In_2828,In_3463);
nand U1204 (N_1204,In_139,In_1806);
or U1205 (N_1205,N_739,In_57);
nand U1206 (N_1206,In_2627,In_4842);
or U1207 (N_1207,In_1449,In_1171);
nand U1208 (N_1208,In_2546,In_2616);
and U1209 (N_1209,In_2586,In_2951);
nor U1210 (N_1210,In_2474,In_4893);
nand U1211 (N_1211,In_1861,In_1024);
nor U1212 (N_1212,In_2276,In_607);
and U1213 (N_1213,In_2864,In_2254);
nor U1214 (N_1214,In_3863,In_1592);
or U1215 (N_1215,In_2607,In_2722);
and U1216 (N_1216,In_2431,In_855);
nor U1217 (N_1217,N_698,In_4764);
xor U1218 (N_1218,In_4578,N_174);
and U1219 (N_1219,In_507,In_2519);
and U1220 (N_1220,In_435,In_4279);
nand U1221 (N_1221,N_190,In_3100);
nor U1222 (N_1222,In_3318,In_4241);
nand U1223 (N_1223,N_212,In_4197);
or U1224 (N_1224,In_488,In_264);
and U1225 (N_1225,N_482,In_3967);
xor U1226 (N_1226,N_586,In_4315);
or U1227 (N_1227,In_3668,In_1626);
nand U1228 (N_1228,In_2785,In_695);
and U1229 (N_1229,In_2706,In_4753);
or U1230 (N_1230,N_525,In_2845);
nand U1231 (N_1231,In_3492,N_644);
and U1232 (N_1232,In_1333,N_935);
nor U1233 (N_1233,In_1532,In_2759);
nand U1234 (N_1234,In_1049,In_1546);
xor U1235 (N_1235,In_1490,In_1324);
or U1236 (N_1236,N_221,In_819);
and U1237 (N_1237,N_790,N_326);
xnor U1238 (N_1238,In_268,In_1353);
xor U1239 (N_1239,In_2942,In_4380);
xor U1240 (N_1240,In_4522,In_17);
or U1241 (N_1241,In_1572,In_1043);
xnor U1242 (N_1242,In_3320,N_408);
nor U1243 (N_1243,N_545,N_981);
xor U1244 (N_1244,In_1936,In_4712);
and U1245 (N_1245,In_2249,In_2093);
nand U1246 (N_1246,N_155,In_3127);
or U1247 (N_1247,In_4947,In_2836);
and U1248 (N_1248,N_833,In_4715);
nand U1249 (N_1249,N_872,In_62);
xor U1250 (N_1250,In_35,In_3599);
and U1251 (N_1251,N_838,In_4126);
xor U1252 (N_1252,In_4819,In_4683);
and U1253 (N_1253,In_4415,In_917);
xnor U1254 (N_1254,N_1111,In_623);
xnor U1255 (N_1255,N_403,In_1114);
nand U1256 (N_1256,In_2631,In_1440);
xnor U1257 (N_1257,N_839,In_2537);
nor U1258 (N_1258,In_452,In_2377);
and U1259 (N_1259,In_580,In_2466);
or U1260 (N_1260,In_2058,In_1026);
or U1261 (N_1261,In_149,N_986);
and U1262 (N_1262,N_961,In_2504);
xnor U1263 (N_1263,In_3651,In_112);
and U1264 (N_1264,In_3330,In_894);
or U1265 (N_1265,In_2964,N_12);
or U1266 (N_1266,N_709,In_596);
or U1267 (N_1267,In_4232,In_3375);
xor U1268 (N_1268,N_66,In_327);
nor U1269 (N_1269,N_1150,In_2057);
xnor U1270 (N_1270,In_4647,In_841);
or U1271 (N_1271,In_363,In_4408);
or U1272 (N_1272,In_1612,In_942);
xor U1273 (N_1273,In_813,In_2749);
nand U1274 (N_1274,In_4747,N_599);
or U1275 (N_1275,In_2371,In_579);
nor U1276 (N_1276,In_2119,In_3111);
nand U1277 (N_1277,In_3936,In_2217);
and U1278 (N_1278,In_2214,In_2082);
or U1279 (N_1279,In_1091,In_3785);
nor U1280 (N_1280,N_181,N_185);
xnor U1281 (N_1281,In_4373,In_1748);
and U1282 (N_1282,In_1793,In_229);
xnor U1283 (N_1283,In_3125,N_454);
xor U1284 (N_1284,In_4542,In_1569);
nor U1285 (N_1285,N_785,In_3023);
and U1286 (N_1286,N_198,In_424);
nor U1287 (N_1287,In_999,In_2533);
xnor U1288 (N_1288,In_2270,In_3317);
xnor U1289 (N_1289,In_3880,In_458);
nor U1290 (N_1290,In_2603,N_16);
xnor U1291 (N_1291,In_3846,In_1827);
and U1292 (N_1292,In_2380,In_4676);
nor U1293 (N_1293,N_1012,N_1136);
and U1294 (N_1294,In_2800,In_2958);
xnor U1295 (N_1295,N_1207,In_1970);
nand U1296 (N_1296,In_1632,In_1824);
or U1297 (N_1297,In_2989,In_2604);
or U1298 (N_1298,In_1794,In_3932);
and U1299 (N_1299,In_1969,In_724);
and U1300 (N_1300,In_444,N_873);
nand U1301 (N_1301,N_749,In_3085);
nor U1302 (N_1302,N_477,In_3255);
xor U1303 (N_1303,In_2739,N_913);
nand U1304 (N_1304,N_1026,In_1934);
nand U1305 (N_1305,N_791,In_1677);
nand U1306 (N_1306,In_540,In_2230);
xnor U1307 (N_1307,In_1284,In_2147);
nor U1308 (N_1308,In_939,In_2375);
and U1309 (N_1309,In_2334,In_154);
or U1310 (N_1310,N_1004,In_2751);
nor U1311 (N_1311,In_20,In_3003);
nor U1312 (N_1312,In_1555,In_1186);
and U1313 (N_1313,In_4084,In_973);
and U1314 (N_1314,In_1447,In_2877);
nor U1315 (N_1315,N_192,In_657);
nand U1316 (N_1316,In_4588,In_3442);
nand U1317 (N_1317,In_1421,N_182);
xor U1318 (N_1318,In_799,In_1420);
and U1319 (N_1319,In_4173,In_2585);
and U1320 (N_1320,In_4171,In_1871);
nor U1321 (N_1321,N_994,In_407);
or U1322 (N_1322,N_451,N_925);
nor U1323 (N_1323,In_1795,In_3062);
and U1324 (N_1324,In_4865,In_1025);
xor U1325 (N_1325,In_1834,In_60);
nand U1326 (N_1326,N_9,In_175);
xor U1327 (N_1327,In_4662,In_2187);
xnor U1328 (N_1328,In_4365,N_253);
xor U1329 (N_1329,In_4996,In_1743);
or U1330 (N_1330,In_612,N_850);
or U1331 (N_1331,In_1910,N_706);
nor U1332 (N_1332,In_3609,In_3507);
or U1333 (N_1333,In_477,In_3960);
and U1334 (N_1334,N_1074,In_489);
or U1335 (N_1335,In_1681,In_1037);
nor U1336 (N_1336,In_2182,In_3374);
nand U1337 (N_1337,In_378,In_659);
nor U1338 (N_1338,In_3323,In_556);
nor U1339 (N_1339,In_1201,In_1257);
nand U1340 (N_1340,In_22,In_692);
and U1341 (N_1341,In_1271,In_433);
and U1342 (N_1342,N_1152,N_431);
or U1343 (N_1343,In_2618,In_183);
nor U1344 (N_1344,N_1133,In_4909);
xor U1345 (N_1345,In_3258,In_411);
xnor U1346 (N_1346,In_3598,In_2181);
or U1347 (N_1347,In_3759,N_496);
and U1348 (N_1348,In_4317,In_3236);
or U1349 (N_1349,In_4102,In_2019);
nor U1350 (N_1350,In_1529,In_1590);
or U1351 (N_1351,In_4803,In_2775);
xor U1352 (N_1352,N_680,In_2851);
xor U1353 (N_1353,In_3784,N_617);
xnor U1354 (N_1354,N_848,N_470);
and U1355 (N_1355,In_4024,N_222);
or U1356 (N_1356,In_3099,N_639);
and U1357 (N_1357,In_4867,N_537);
nand U1358 (N_1358,N_557,In_4581);
and U1359 (N_1359,N_331,In_3555);
nand U1360 (N_1360,In_3266,In_423);
nor U1361 (N_1361,In_3634,In_4938);
nor U1362 (N_1362,In_2490,N_905);
or U1363 (N_1363,In_1399,In_3448);
and U1364 (N_1364,In_4497,N_821);
and U1365 (N_1365,In_4469,N_127);
nor U1366 (N_1366,In_3001,In_3868);
xor U1367 (N_1367,In_4922,In_1369);
xnor U1368 (N_1368,N_1092,In_2806);
xnor U1369 (N_1369,In_2818,In_2084);
xor U1370 (N_1370,In_2512,In_287);
xor U1371 (N_1371,N_970,In_3537);
xor U1372 (N_1372,In_1630,N_690);
or U1373 (N_1373,In_4484,In_85);
and U1374 (N_1374,In_442,N_1245);
xor U1375 (N_1375,In_84,In_4185);
or U1376 (N_1376,In_4264,In_3110);
nor U1377 (N_1377,In_1864,N_761);
nand U1378 (N_1378,In_4131,In_2125);
and U1379 (N_1379,N_567,N_836);
and U1380 (N_1380,In_2323,N_1230);
and U1381 (N_1381,In_4896,In_3044);
nand U1382 (N_1382,N_1043,N_748);
nand U1383 (N_1383,In_3490,N_614);
xor U1384 (N_1384,N_1044,In_3413);
xor U1385 (N_1385,In_3706,In_13);
or U1386 (N_1386,N_299,In_4994);
or U1387 (N_1387,In_2862,In_4927);
and U1388 (N_1388,In_3045,N_173);
nor U1389 (N_1389,In_750,In_4692);
xnor U1390 (N_1390,N_114,In_4215);
and U1391 (N_1391,In_274,N_507);
or U1392 (N_1392,In_3244,In_345);
or U1393 (N_1393,In_1671,N_587);
nor U1394 (N_1394,In_4778,In_2926);
or U1395 (N_1395,In_3194,In_426);
xor U1396 (N_1396,In_1245,N_869);
nand U1397 (N_1397,In_4563,In_1499);
nand U1398 (N_1398,In_1138,In_2708);
nand U1399 (N_1399,In_1985,In_4275);
or U1400 (N_1400,N_374,In_737);
and U1401 (N_1401,In_4624,In_4231);
and U1402 (N_1402,In_2378,In_1148);
or U1403 (N_1403,In_2990,N_311);
nor U1404 (N_1404,In_2886,In_677);
xnor U1405 (N_1405,In_2083,N_685);
xnor U1406 (N_1406,In_719,In_4059);
xor U1407 (N_1407,In_4021,In_2801);
nand U1408 (N_1408,In_2153,N_669);
nor U1409 (N_1409,In_409,In_4323);
nand U1410 (N_1410,In_3364,In_2506);
nand U1411 (N_1411,N_809,In_2291);
or U1412 (N_1412,In_182,In_1953);
nor U1413 (N_1413,In_457,In_1652);
and U1414 (N_1414,N_933,In_3951);
xor U1415 (N_1415,In_2978,In_601);
xnor U1416 (N_1416,In_4766,In_826);
or U1417 (N_1417,In_575,N_1076);
and U1418 (N_1418,In_3954,In_558);
nand U1419 (N_1419,In_2294,In_3793);
or U1420 (N_1420,N_1161,In_114);
xor U1421 (N_1421,N_468,In_368);
nor U1422 (N_1422,In_1686,In_3000);
or U1423 (N_1423,In_383,N_429);
and U1424 (N_1424,In_1331,In_4307);
or U1425 (N_1425,In_1157,N_144);
xor U1426 (N_1426,In_408,In_3860);
nand U1427 (N_1427,In_2434,N_957);
nand U1428 (N_1428,In_3904,In_4868);
xnor U1429 (N_1429,In_2140,In_4123);
nor U1430 (N_1430,N_758,In_757);
or U1431 (N_1431,In_684,N_1100);
and U1432 (N_1432,N_1138,N_966);
nand U1433 (N_1433,In_334,N_574);
nand U1434 (N_1434,N_1112,In_387);
xnor U1435 (N_1435,In_2023,In_75);
xnor U1436 (N_1436,N_535,In_4499);
nor U1437 (N_1437,N_1014,In_2319);
xor U1438 (N_1438,N_390,N_1030);
or U1439 (N_1439,In_3180,In_1095);
or U1440 (N_1440,N_664,N_1046);
xor U1441 (N_1441,In_4494,In_3739);
nor U1442 (N_1442,N_589,In_2915);
nor U1443 (N_1443,In_3384,N_551);
and U1444 (N_1444,In_2313,N_951);
xnor U1445 (N_1445,In_3900,N_906);
and U1446 (N_1446,In_4936,In_2451);
and U1447 (N_1447,In_1321,N_1184);
and U1448 (N_1448,In_4758,N_263);
and U1449 (N_1449,N_1090,In_3844);
and U1450 (N_1450,In_289,In_1637);
and U1451 (N_1451,N_210,In_3309);
or U1452 (N_1452,In_1724,In_902);
and U1453 (N_1453,In_342,N_1190);
nor U1454 (N_1454,In_4376,In_1469);
and U1455 (N_1455,In_4681,N_604);
xnor U1456 (N_1456,In_2418,In_2143);
and U1457 (N_1457,N_265,In_1137);
nor U1458 (N_1458,In_3612,N_1168);
nor U1459 (N_1459,In_348,In_882);
nor U1460 (N_1460,In_1899,In_4872);
nand U1461 (N_1461,In_3214,In_2361);
nand U1462 (N_1462,In_4254,In_1260);
nor U1463 (N_1463,In_2202,In_1514);
xnor U1464 (N_1464,N_541,N_140);
xnor U1465 (N_1465,N_950,In_1647);
and U1466 (N_1466,In_3862,In_4154);
or U1467 (N_1467,N_630,In_3799);
xnor U1468 (N_1468,In_3497,N_707);
xor U1469 (N_1469,In_2241,In_4549);
xnor U1470 (N_1470,N_383,In_2661);
nor U1471 (N_1471,In_3743,In_3102);
nor U1472 (N_1472,In_2250,In_4711);
and U1473 (N_1473,In_528,N_837);
nand U1474 (N_1474,N_105,In_222);
xnor U1475 (N_1475,In_4607,In_1487);
xor U1476 (N_1476,N_409,In_2032);
xnor U1477 (N_1477,In_89,In_2479);
or U1478 (N_1478,In_3623,In_3774);
or U1479 (N_1479,N_998,In_3493);
nand U1480 (N_1480,N_621,In_401);
or U1481 (N_1481,In_343,N_471);
or U1482 (N_1482,In_803,In_3470);
or U1483 (N_1483,In_3636,N_825);
xnor U1484 (N_1484,In_1511,N_623);
nor U1485 (N_1485,N_1149,In_4338);
xnor U1486 (N_1486,In_723,N_955);
xor U1487 (N_1487,N_509,In_2975);
and U1488 (N_1488,In_2154,N_546);
xnor U1489 (N_1489,In_2509,In_1751);
nand U1490 (N_1490,In_1403,In_660);
nand U1491 (N_1491,In_4175,N_550);
nor U1492 (N_1492,N_767,In_991);
nor U1493 (N_1493,In_463,In_510);
or U1494 (N_1494,In_1898,N_708);
and U1495 (N_1495,In_2771,N_1163);
xor U1496 (N_1496,In_3417,N_340);
xnor U1497 (N_1497,In_1481,In_3715);
and U1498 (N_1498,In_4135,In_583);
xor U1499 (N_1499,N_548,N_3);
and U1500 (N_1500,In_650,In_2198);
nand U1501 (N_1501,In_3596,N_1274);
nand U1502 (N_1502,In_3717,In_3756);
and U1503 (N_1503,N_830,In_2953);
nand U1504 (N_1504,N_271,In_1135);
xnor U1505 (N_1505,In_941,In_1096);
and U1506 (N_1506,In_3171,In_1253);
nand U1507 (N_1507,In_1452,In_4291);
nor U1508 (N_1508,In_3074,In_2100);
or U1509 (N_1509,N_884,In_2203);
and U1510 (N_1510,N_449,In_3769);
nand U1511 (N_1511,In_4468,In_2770);
and U1512 (N_1512,In_4004,N_822);
nand U1513 (N_1513,In_3394,In_3038);
xnor U1514 (N_1514,In_776,In_1721);
and U1515 (N_1515,In_4587,In_4987);
or U1516 (N_1516,In_2523,In_2888);
or U1517 (N_1517,N_1307,In_3663);
xnor U1518 (N_1518,In_2101,In_3869);
and U1519 (N_1519,N_719,In_2686);
nand U1520 (N_1520,In_34,In_4492);
and U1521 (N_1521,N_1415,N_1122);
or U1522 (N_1522,In_4013,In_429);
and U1523 (N_1523,N_503,N_1419);
and U1524 (N_1524,In_4061,In_655);
and U1525 (N_1525,In_2897,N_1318);
or U1526 (N_1526,In_3622,N_699);
and U1527 (N_1527,In_3877,In_2394);
xor U1528 (N_1528,In_4833,In_2223);
nand U1529 (N_1529,In_2620,N_474);
xor U1530 (N_1530,In_653,In_4422);
xnor U1531 (N_1531,In_3065,In_4141);
xor U1532 (N_1532,N_232,N_1414);
nor U1533 (N_1533,In_3679,In_4570);
nor U1534 (N_1534,N_439,In_3524);
or U1535 (N_1535,In_4946,In_214);
xor U1536 (N_1536,In_2454,N_1449);
or U1537 (N_1537,In_4580,In_128);
nor U1538 (N_1538,In_3290,In_4598);
nand U1539 (N_1539,N_910,In_4420);
xor U1540 (N_1540,N_490,N_63);
nor U1541 (N_1541,In_3587,N_555);
and U1542 (N_1542,In_1228,N_938);
or U1543 (N_1543,In_3088,In_3711);
and U1544 (N_1544,In_1996,In_2562);
and U1545 (N_1545,In_3980,N_854);
and U1546 (N_1546,N_667,N_1164);
xnor U1547 (N_1547,In_4705,In_2264);
xnor U1548 (N_1548,N_1080,In_758);
nor U1549 (N_1549,In_1679,In_1474);
or U1550 (N_1550,In_4106,N_1096);
or U1551 (N_1551,In_1757,N_1317);
and U1552 (N_1552,In_4033,N_1120);
nand U1553 (N_1553,In_72,In_4740);
xnor U1554 (N_1554,In_4900,In_3489);
xor U1555 (N_1555,In_932,In_4293);
xor U1556 (N_1556,In_532,N_68);
and U1557 (N_1557,N_1219,In_4316);
and U1558 (N_1558,In_1919,In_2017);
and U1559 (N_1559,In_1028,In_1313);
nand U1560 (N_1560,In_4773,N_1248);
nand U1561 (N_1561,In_2066,N_687);
nor U1562 (N_1562,In_2675,N_553);
or U1563 (N_1563,In_2255,In_3677);
or U1564 (N_1564,N_652,In_3396);
nor U1565 (N_1565,In_1712,In_2482);
nand U1566 (N_1566,N_1359,N_244);
and U1567 (N_1567,N_115,N_642);
xnor U1568 (N_1568,In_4898,In_2730);
xor U1569 (N_1569,In_4793,In_3008);
and U1570 (N_1570,N_673,In_4251);
nor U1571 (N_1571,In_4063,In_3115);
nand U1572 (N_1572,In_1289,In_4281);
xor U1573 (N_1573,In_122,In_4694);
or U1574 (N_1574,In_1786,In_3332);
nor U1575 (N_1575,N_959,In_4030);
nand U1576 (N_1576,In_3392,In_3471);
nor U1577 (N_1577,In_4879,N_695);
and U1578 (N_1578,In_562,In_375);
nand U1579 (N_1579,N_1225,N_98);
nor U1580 (N_1580,In_3938,In_2406);
nand U1581 (N_1581,In_1547,In_1683);
xor U1582 (N_1582,In_3325,In_549);
nor U1583 (N_1583,In_2505,In_2503);
or U1584 (N_1584,In_82,N_1347);
and U1585 (N_1585,In_3424,In_1168);
nor U1586 (N_1586,In_4966,N_965);
nor U1587 (N_1587,In_4090,In_1159);
and U1588 (N_1588,In_3054,In_3185);
nand U1589 (N_1589,N_107,In_4977);
nor U1590 (N_1590,In_3892,In_4056);
and U1591 (N_1591,In_339,In_1296);
nand U1592 (N_1592,In_196,In_317);
xor U1593 (N_1593,In_133,In_1086);
and U1594 (N_1594,In_2545,In_4345);
or U1595 (N_1595,In_4130,In_1259);
and U1596 (N_1596,N_777,In_4792);
nor U1597 (N_1597,In_2034,In_4409);
nor U1598 (N_1598,N_1470,In_4050);
xnor U1599 (N_1599,In_3329,In_2458);
nor U1600 (N_1600,In_928,In_4668);
and U1601 (N_1601,In_250,In_1465);
and U1602 (N_1602,In_49,In_490);
nor U1603 (N_1603,N_1197,In_2114);
and U1604 (N_1604,In_2179,N_178);
and U1605 (N_1605,In_4618,N_230);
nand U1606 (N_1606,In_2099,In_413);
nand U1607 (N_1607,In_3533,In_4505);
or U1608 (N_1608,N_1068,In_534);
and U1609 (N_1609,In_3030,In_4213);
xnor U1610 (N_1610,In_3796,In_1697);
xor U1611 (N_1611,In_2873,In_3466);
xnor U1612 (N_1612,N_808,N_921);
or U1613 (N_1613,In_376,N_294);
xnor U1614 (N_1614,N_876,In_1693);
and U1615 (N_1615,N_1457,In_1209);
xnor U1616 (N_1616,In_2516,N_1202);
nor U1617 (N_1617,In_146,In_618);
nand U1618 (N_1618,In_4356,In_3024);
nand U1619 (N_1619,In_4222,In_3834);
xor U1620 (N_1620,N_1135,In_1846);
and U1621 (N_1621,N_730,In_4028);
nor U1622 (N_1622,In_2122,In_187);
nand U1623 (N_1623,In_781,In_3270);
nand U1624 (N_1624,N_1312,N_524);
nor U1625 (N_1625,In_3357,In_1063);
xor U1626 (N_1626,In_3969,In_157);
nor U1627 (N_1627,In_2472,In_3057);
and U1628 (N_1628,N_975,In_4599);
nor U1629 (N_1629,In_945,In_3911);
xor U1630 (N_1630,In_1853,In_3866);
nor U1631 (N_1631,In_4129,In_770);
nor U1632 (N_1632,In_1177,N_844);
nand U1633 (N_1633,N_1006,In_4912);
or U1634 (N_1634,In_2128,In_177);
or U1635 (N_1635,In_3487,N_882);
nor U1636 (N_1636,In_1700,In_4172);
or U1637 (N_1637,In_969,In_756);
nor U1638 (N_1638,In_2717,N_926);
nand U1639 (N_1639,In_3736,N_722);
nand U1640 (N_1640,N_19,In_1500);
or U1641 (N_1641,In_1802,In_3036);
nor U1642 (N_1642,In_1492,In_4797);
and U1643 (N_1643,In_3920,N_1461);
or U1644 (N_1644,In_1818,In_1226);
nand U1645 (N_1645,In_318,In_1273);
nand U1646 (N_1646,N_1251,In_4266);
and U1647 (N_1647,In_3161,In_3603);
nor U1648 (N_1648,N_268,In_1839);
nor U1649 (N_1649,In_1169,In_2633);
and U1650 (N_1650,In_2736,N_893);
nor U1651 (N_1651,In_547,In_1635);
or U1652 (N_1652,In_4544,N_1280);
or U1653 (N_1653,In_10,In_2008);
nor U1654 (N_1654,In_4427,N_249);
nand U1655 (N_1655,N_568,In_4645);
nand U1656 (N_1656,N_1383,In_380);
nand U1657 (N_1657,In_1081,N_113);
and U1658 (N_1658,In_3727,In_3883);
or U1659 (N_1659,In_4691,In_2715);
or U1660 (N_1660,N_1388,N_727);
nand U1661 (N_1661,In_4082,N_1475);
and U1662 (N_1662,In_2599,In_2536);
and U1663 (N_1663,In_1290,N_733);
nor U1664 (N_1664,N_1087,In_2612);
nand U1665 (N_1665,In_1885,In_1542);
nor U1666 (N_1666,In_4443,In_1600);
or U1667 (N_1667,In_258,In_2732);
nor U1668 (N_1668,In_4489,N_608);
or U1669 (N_1669,N_894,N_747);
or U1670 (N_1670,N_547,In_2020);
xor U1671 (N_1671,In_1470,In_1718);
nor U1672 (N_1672,N_1261,In_3241);
nor U1673 (N_1673,In_1657,In_4117);
xor U1674 (N_1674,In_2615,In_1900);
xnor U1675 (N_1675,In_4579,In_2705);
nor U1676 (N_1676,N_1303,In_769);
nand U1677 (N_1677,N_1060,In_1932);
nand U1678 (N_1678,In_4916,In_2260);
xor U1679 (N_1679,In_123,N_686);
nor U1680 (N_1680,In_295,N_1294);
or U1681 (N_1681,In_2275,In_2895);
nor U1682 (N_1682,N_827,In_3572);
nand U1683 (N_1683,In_1651,In_3585);
and U1684 (N_1684,N_197,In_4685);
xor U1685 (N_1685,In_302,In_1187);
xnor U1686 (N_1686,N_267,In_3302);
and U1687 (N_1687,N_1395,In_4703);
nand U1688 (N_1688,In_4410,In_3403);
and U1689 (N_1689,N_1067,In_1014);
or U1690 (N_1690,In_4177,In_2623);
nand U1691 (N_1691,In_3025,In_2130);
or U1692 (N_1692,In_561,N_702);
and U1693 (N_1693,In_3517,In_1769);
xnor U1694 (N_1694,N_1436,In_3855);
or U1695 (N_1695,In_977,N_1485);
nand U1696 (N_1696,N_1393,In_3510);
xnor U1697 (N_1697,N_1002,In_3680);
and U1698 (N_1698,N_1416,In_3747);
nand U1699 (N_1699,N_1275,In_2247);
nor U1700 (N_1700,N_8,In_2457);
nor U1701 (N_1701,In_384,In_2881);
or U1702 (N_1702,N_1233,In_872);
nand U1703 (N_1703,In_68,In_4112);
or U1704 (N_1704,In_71,N_375);
and U1705 (N_1705,In_3964,In_889);
nor U1706 (N_1706,In_1692,In_1006);
nand U1707 (N_1707,N_1229,In_3109);
xnor U1708 (N_1708,N_1192,In_1057);
nand U1709 (N_1709,N_752,In_1616);
xnor U1710 (N_1710,N_302,In_2558);
and U1711 (N_1711,In_3269,N_1095);
or U1712 (N_1712,In_1564,In_246);
and U1713 (N_1713,In_2849,N_1341);
xnor U1714 (N_1714,In_4482,In_3086);
or U1715 (N_1715,N_753,In_3775);
or U1716 (N_1716,In_2238,In_3801);
or U1717 (N_1717,In_2822,In_1988);
nor U1718 (N_1718,In_4303,In_2768);
and U1719 (N_1719,N_180,In_3605);
nor U1720 (N_1720,In_3703,In_4603);
nor U1721 (N_1721,N_1139,N_506);
xor U1722 (N_1722,In_2061,In_2655);
nand U1723 (N_1723,N_881,In_3387);
or U1724 (N_1724,In_2500,In_3923);
and U1725 (N_1725,N_380,N_57);
and U1726 (N_1726,In_913,In_4658);
and U1727 (N_1727,In_818,In_2556);
and U1728 (N_1728,In_3118,In_4777);
and U1729 (N_1729,In_4081,In_1478);
nand U1730 (N_1730,N_1005,In_2764);
xnor U1731 (N_1731,N_1211,In_2108);
xor U1732 (N_1732,In_1894,In_26);
nand U1733 (N_1733,In_3836,In_4441);
or U1734 (N_1734,In_1256,In_1916);
xnor U1735 (N_1735,In_3872,In_793);
or U1736 (N_1736,In_3141,N_755);
nand U1737 (N_1737,N_1191,In_3019);
and U1738 (N_1738,N_866,In_3754);
and U1739 (N_1739,In_3975,In_1280);
and U1740 (N_1740,N_843,In_3786);
xnor U1741 (N_1741,In_1124,N_863);
xor U1742 (N_1742,In_3597,N_37);
and U1743 (N_1743,N_303,N_1375);
nor U1744 (N_1744,In_1706,N_201);
or U1745 (N_1745,In_2983,In_3854);
or U1746 (N_1746,N_53,N_60);
or U1747 (N_1747,In_280,In_4706);
xnor U1748 (N_1748,In_3368,N_1253);
xnor U1749 (N_1749,In_1036,N_648);
nor U1750 (N_1750,N_564,In_1579);
or U1751 (N_1751,In_1293,In_153);
or U1752 (N_1752,N_600,N_1397);
nand U1753 (N_1753,In_2816,N_1327);
or U1754 (N_1754,In_3257,In_705);
xor U1755 (N_1755,In_4808,N_1629);
nand U1756 (N_1756,In_1909,N_1456);
and U1757 (N_1757,In_3020,N_1520);
and U1758 (N_1758,In_2852,N_828);
xor U1759 (N_1759,N_1086,In_3452);
nor U1760 (N_1760,N_1035,N_704);
nand U1761 (N_1761,N_1580,In_3046);
nor U1762 (N_1762,In_3346,In_903);
nor U1763 (N_1763,In_4688,N_1705);
xor U1764 (N_1764,N_849,In_4358);
and U1765 (N_1765,N_1662,In_548);
nor U1766 (N_1766,In_4527,In_4089);
or U1767 (N_1767,N_1377,In_2421);
nand U1768 (N_1768,N_1737,N_847);
nand U1769 (N_1769,In_4202,In_1263);
nor U1770 (N_1770,In_2850,In_2912);
or U1771 (N_1771,N_266,N_1648);
nor U1772 (N_1772,In_2542,N_880);
and U1773 (N_1773,In_1238,N_1151);
and U1774 (N_1774,In_467,N_601);
xor U1775 (N_1775,N_1684,In_4787);
nand U1776 (N_1776,In_2422,N_607);
nand U1777 (N_1777,In_2383,N_1003);
xnor U1778 (N_1778,In_1734,In_2022);
nor U1779 (N_1779,N_531,N_1306);
nor U1780 (N_1780,N_1235,N_1380);
nor U1781 (N_1781,N_1309,In_4357);
or U1782 (N_1782,N_49,N_22);
xor U1783 (N_1783,In_279,N_1365);
nor U1784 (N_1784,In_2672,In_946);
nand U1785 (N_1785,N_1669,N_1301);
nor U1786 (N_1786,N_1728,N_769);
or U1787 (N_1787,In_3037,In_4958);
nor U1788 (N_1788,In_1575,N_111);
xnor U1789 (N_1789,N_875,N_344);
nand U1790 (N_1790,In_1738,N_1539);
nor U1791 (N_1791,N_766,In_1986);
xor U1792 (N_1792,In_2572,In_4480);
or U1793 (N_1793,In_509,In_1150);
xnor U1794 (N_1794,N_83,In_209);
or U1795 (N_1795,N_1215,In_1833);
nand U1796 (N_1796,In_4613,In_2103);
and U1797 (N_1797,In_1796,In_2485);
nor U1798 (N_1798,N_888,N_517);
or U1799 (N_1799,In_2356,N_472);
xor U1800 (N_1800,In_2156,N_1497);
nand U1801 (N_1801,In_1604,In_1921);
xnor U1802 (N_1802,N_188,In_786);
and U1803 (N_1803,In_3961,In_4198);
xnor U1804 (N_1804,In_4660,N_1692);
xor U1805 (N_1805,In_2874,N_213);
and U1806 (N_1806,In_2258,In_1140);
or U1807 (N_1807,In_2050,In_395);
or U1808 (N_1808,N_1278,N_206);
or U1809 (N_1809,N_1496,In_2475);
or U1810 (N_1810,N_1231,N_1355);
nand U1811 (N_1811,In_3282,In_530);
and U1812 (N_1812,In_4016,In_4539);
or U1813 (N_1813,In_1456,In_3271);
nand U1814 (N_1814,In_3084,In_551);
nand U1815 (N_1815,N_1600,In_4874);
or U1816 (N_1816,N_1308,N_280);
or U1817 (N_1817,In_2463,In_4627);
nand U1818 (N_1818,In_2180,N_118);
nand U1819 (N_1819,In_1035,In_2638);
or U1820 (N_1820,In_2262,In_2815);
or U1821 (N_1821,N_67,In_1598);
xor U1822 (N_1822,N_781,N_1450);
and U1823 (N_1823,In_1316,N_852);
and U1824 (N_1824,N_463,In_4104);
xnor U1825 (N_1825,In_1872,N_1260);
or U1826 (N_1826,In_3781,In_3080);
nand U1827 (N_1827,N_1503,N_1606);
nor U1828 (N_1828,In_456,N_324);
nor U1829 (N_1829,In_2943,In_2216);
nand U1830 (N_1830,In_2737,N_1256);
nor U1831 (N_1831,N_1656,In_3982);
nand U1832 (N_1832,N_1382,N_591);
and U1833 (N_1833,In_79,In_3063);
or U1834 (N_1834,In_4310,In_197);
nand U1835 (N_1835,In_96,In_4048);
and U1836 (N_1836,N_554,In_3940);
or U1837 (N_1837,N_10,N_1593);
or U1838 (N_1838,In_3350,In_3223);
xor U1839 (N_1839,In_87,N_1627);
xnor U1840 (N_1840,In_1531,In_1608);
nor U1841 (N_1841,In_4370,In_752);
or U1842 (N_1842,In_644,N_846);
nor U1843 (N_1843,N_1266,In_1340);
xor U1844 (N_1844,N_922,In_99);
nand U1845 (N_1845,N_549,N_1102);
xnor U1846 (N_1846,In_4837,In_985);
or U1847 (N_1847,N_293,In_1924);
or U1848 (N_1848,In_3310,N_1063);
nor U1849 (N_1849,In_791,In_2430);
or U1850 (N_1850,In_1488,In_4905);
xnor U1851 (N_1851,In_1468,N_1495);
xor U1852 (N_1852,N_1289,In_460);
nand U1853 (N_1853,N_1165,N_779);
nand U1854 (N_1854,In_3733,N_1367);
nor U1855 (N_1855,In_1070,N_1667);
nand U1856 (N_1856,N_1170,In_3436);
xor U1857 (N_1857,In_2415,N_917);
nand U1858 (N_1858,N_247,N_396);
xor U1859 (N_1859,In_3372,N_1130);
and U1860 (N_1860,N_1302,N_742);
or U1861 (N_1861,N_1586,In_4968);
xnor U1862 (N_1862,N_513,N_578);
nand U1863 (N_1863,N_1736,In_4838);
nor U1864 (N_1864,In_2548,In_2157);
nand U1865 (N_1865,N_1244,In_4255);
and U1866 (N_1866,N_1446,In_3852);
nand U1867 (N_1867,In_1845,N_1597);
nand U1868 (N_1868,In_885,In_310);
and U1869 (N_1869,In_3850,In_2407);
nand U1870 (N_1870,In_3963,N_1482);
and U1871 (N_1871,In_2727,In_2056);
nand U1872 (N_1872,In_1495,N_1709);
nor U1873 (N_1873,In_577,N_976);
xnor U1874 (N_1874,In_3331,In_978);
xor U1875 (N_1875,In_3153,In_3819);
nand U1876 (N_1876,In_3988,In_949);
nand U1877 (N_1877,In_263,In_4120);
or U1878 (N_1878,In_3722,N_1045);
nor U1879 (N_1879,In_1685,In_240);
nand U1880 (N_1880,In_2285,N_1494);
and U1881 (N_1881,In_517,In_1254);
nand U1882 (N_1882,In_333,In_4604);
or U1883 (N_1883,In_3087,In_278);
nand U1884 (N_1884,N_1543,In_319);
and U1885 (N_1885,In_3755,N_227);
or U1886 (N_1886,In_732,In_3380);
nor U1887 (N_1887,In_3126,In_1005);
nand U1888 (N_1888,N_1646,N_1371);
or U1889 (N_1889,N_1440,In_231);
or U1890 (N_1890,N_1735,In_2602);
xnor U1891 (N_1891,In_2184,In_4046);
nand U1892 (N_1892,In_2158,In_1882);
nand U1893 (N_1893,In_2301,In_495);
nand U1894 (N_1894,N_1321,N_973);
nor U1895 (N_1895,In_93,N_1048);
or U1896 (N_1896,In_4439,In_3503);
nor U1897 (N_1897,In_1466,N_45);
or U1898 (N_1898,N_1581,N_217);
and U1899 (N_1899,In_1599,In_4402);
xnor U1900 (N_1900,In_3576,N_1406);
and U1901 (N_1901,N_1226,In_2010);
or U1902 (N_1902,In_3947,In_1497);
and U1903 (N_1903,N_817,In_1723);
or U1904 (N_1904,N_1297,In_3215);
nand U1905 (N_1905,In_3772,In_2305);
or U1906 (N_1906,N_1530,In_3289);
or U1907 (N_1907,N_322,N_1304);
or U1908 (N_1908,In_3342,N_1361);
or U1909 (N_1909,In_74,In_2233);
nor U1910 (N_1910,In_876,In_1038);
nand U1911 (N_1911,In_314,In_1093);
and U1912 (N_1912,In_4340,In_667);
and U1913 (N_1913,N_778,In_4805);
xor U1914 (N_1914,N_1689,In_291);
or U1915 (N_1915,In_459,In_4414);
xor U1916 (N_1916,N_1059,In_4009);
and U1917 (N_1917,N_1350,In_2315);
or U1918 (N_1918,In_1641,In_502);
and U1919 (N_1919,In_4075,N_1389);
xor U1920 (N_1920,In_4035,N_1634);
xor U1921 (N_1921,In_1648,N_258);
xnor U1922 (N_1922,In_3712,N_1010);
and U1923 (N_1923,N_1270,In_4822);
nor U1924 (N_1924,In_150,N_281);
or U1925 (N_1925,N_1423,In_451);
nand U1926 (N_1926,In_1620,In_40);
or U1927 (N_1927,N_1137,In_3005);
or U1928 (N_1928,N_1699,N_865);
or U1929 (N_1929,In_4385,N_1607);
xnor U1930 (N_1930,In_1512,In_4092);
xor U1931 (N_1931,N_501,N_1657);
xor U1932 (N_1932,In_2521,N_963);
xor U1933 (N_1933,In_1080,In_4757);
and U1934 (N_1934,In_1484,In_610);
xnor U1935 (N_1935,N_511,In_4466);
xnor U1936 (N_1936,In_1780,In_862);
xnor U1937 (N_1937,N_42,In_1394);
nor U1938 (N_1938,N_1481,In_4990);
and U1939 (N_1939,In_109,In_3201);
and U1940 (N_1940,In_4923,N_1490);
nand U1941 (N_1941,In_3635,N_883);
xor U1942 (N_1942,In_4432,In_2718);
or U1943 (N_1943,N_832,N_1366);
and U1944 (N_1944,In_4334,In_4364);
nand U1945 (N_1945,In_4289,In_4534);
xor U1946 (N_1946,N_860,In_2047);
and U1947 (N_1947,In_614,N_1566);
nand U1948 (N_1948,In_472,In_4765);
nor U1949 (N_1949,In_4314,In_1395);
and U1950 (N_1950,In_412,N_526);
and U1951 (N_1951,N_1117,In_2738);
or U1952 (N_1952,N_240,N_1647);
or U1953 (N_1953,In_168,In_3874);
and U1954 (N_1954,N_711,In_2097);
or U1955 (N_1955,In_3009,In_179);
nor U1956 (N_1956,N_1198,N_813);
nand U1957 (N_1957,In_3536,In_3802);
nor U1958 (N_1958,N_405,In_3667);
xnor U1959 (N_1959,In_1739,In_4884);
or U1960 (N_1960,N_498,In_2530);
nand U1961 (N_1961,In_1078,In_1704);
nand U1962 (N_1962,In_24,In_2259);
or U1963 (N_1963,In_4403,In_3351);
nand U1964 (N_1964,In_2596,N_1549);
nor U1965 (N_1965,N_641,N_1480);
or U1966 (N_1966,In_535,N_1670);
and U1967 (N_1967,N_1655,In_2477);
nor U1968 (N_1968,In_2325,In_142);
nor U1969 (N_1969,In_496,N_1509);
and U1970 (N_1970,In_4659,N_325);
nand U1971 (N_1971,In_3051,N_620);
nand U1972 (N_1972,N_937,N_214);
and U1973 (N_1973,N_1065,In_4165);
or U1974 (N_1974,In_4875,In_1541);
or U1975 (N_1975,In_3807,N_675);
xor U1976 (N_1976,In_2073,N_194);
nor U1977 (N_1977,In_2200,In_1836);
nor U1978 (N_1978,N_1079,In_4086);
nor U1979 (N_1979,In_3530,In_1999);
nor U1980 (N_1980,N_1338,N_780);
and U1981 (N_1981,In_4807,In_4999);
nor U1982 (N_1982,In_1855,N_1590);
nand U1983 (N_1983,N_646,In_1154);
xnor U1984 (N_1984,N_301,In_972);
or U1985 (N_1985,N_1115,In_4965);
nand U1986 (N_1986,In_2006,In_2425);
nand U1987 (N_1987,In_4860,N_93);
and U1988 (N_1988,N_1326,In_1589);
nand U1989 (N_1989,In_4555,In_2707);
nand U1990 (N_1990,In_3625,In_3632);
and U1991 (N_1991,In_694,N_1316);
xnor U1992 (N_1992,N_1159,N_593);
nor U1993 (N_1993,N_295,N_31);
or U1994 (N_1994,N_254,In_2959);
nor U1995 (N_1995,In_4453,In_4851);
and U1996 (N_1996,In_2221,N_376);
nor U1997 (N_1997,N_1473,N_892);
and U1998 (N_1998,In_1094,In_3407);
nand U1999 (N_1999,In_1377,In_697);
or U2000 (N_2000,In_2088,In_3488);
xor U2001 (N_2001,In_1527,N_1695);
nand U2002 (N_2002,In_825,N_476);
or U2003 (N_2003,In_316,In_1548);
and U2004 (N_2004,N_442,In_821);
nor U2005 (N_2005,N_297,In_38);
xnor U2006 (N_2006,N_1519,N_1865);
or U2007 (N_2007,N_1971,In_4670);
nor U2008 (N_2008,In_1935,In_2900);
nand U2009 (N_2009,N_110,N_1803);
xor U2010 (N_2010,In_1577,N_1967);
xor U2011 (N_2011,N_1426,In_4919);
or U2012 (N_2012,In_1303,In_3421);
or U2013 (N_2013,N_505,In_1503);
and U2014 (N_2014,In_1835,N_47);
xor U2015 (N_2015,In_2789,N_1852);
nand U2016 (N_2016,In_3426,In_2389);
xor U2017 (N_2017,N_1688,N_1943);
nor U2018 (N_2018,In_4465,In_3887);
nor U2019 (N_2019,In_1215,In_3343);
xnor U2020 (N_2020,N_1162,N_800);
or U2021 (N_2021,N_1585,N_603);
and U2022 (N_2022,In_796,In_703);
and U2023 (N_2023,In_1172,N_1323);
or U2024 (N_2024,In_3172,In_4597);
nand U2025 (N_2025,In_3462,In_1300);
xnor U2026 (N_2026,In_4236,N_318);
and U2027 (N_2027,In_4521,N_276);
or U2028 (N_2028,N_224,N_241);
xor U2029 (N_2029,In_3973,In_2449);
nand U2030 (N_2030,In_1156,In_2190);
nand U2031 (N_2031,In_1436,In_2242);
nor U2032 (N_2032,In_3393,N_1373);
nand U2033 (N_2033,In_4564,N_1125);
nand U2034 (N_2034,In_1507,N_721);
nor U2035 (N_2035,In_3314,N_1756);
nand U2036 (N_2036,In_4743,In_4064);
nor U2037 (N_2037,N_1979,In_364);
xnor U2038 (N_2038,N_1474,In_283);
nor U2039 (N_2039,N_1927,In_656);
or U2040 (N_2040,In_847,N_121);
xnor U2041 (N_2041,N_734,N_1262);
nor U2042 (N_2042,N_1433,N_1712);
and U2043 (N_2043,N_897,N_528);
nor U2044 (N_2044,N_1913,In_1702);
and U2045 (N_2045,N_1675,N_1123);
nor U2046 (N_2046,N_1546,In_844);
xnor U2047 (N_2047,In_3849,In_635);
nor U2048 (N_2048,N_1224,N_616);
xor U2049 (N_2049,N_1602,In_1272);
and U2050 (N_2050,N_679,N_1058);
and U2051 (N_2051,In_331,In_2658);
or U2052 (N_2052,In_3079,N_1477);
and U2053 (N_2053,N_741,N_416);
nor U2054 (N_2054,In_338,In_4083);
nand U2055 (N_2055,In_892,N_1091);
and U2056 (N_2056,N_1764,N_1733);
and U2057 (N_2057,N_930,In_624);
xor U2058 (N_2058,N_1757,In_4736);
or U2059 (N_2059,N_1890,N_1937);
or U2060 (N_2060,In_605,In_943);
nand U2061 (N_2061,N_356,N_1486);
nand U2062 (N_2062,In_1650,In_2317);
and U2063 (N_2063,In_4483,In_1302);
and U2064 (N_2064,N_1642,In_1979);
xnor U2065 (N_2065,In_4783,In_1830);
and U2066 (N_2066,N_1276,In_4839);
nand U2067 (N_2067,N_1998,In_1244);
nand U2068 (N_2068,In_2569,In_2574);
nand U2069 (N_2069,N_715,N_1742);
and U2070 (N_2070,In_2256,N_953);
xnor U2071 (N_2071,N_1912,In_4639);
nor U2072 (N_2072,In_4446,In_3187);
nor U2073 (N_2073,In_938,In_3308);
nor U2074 (N_2074,In_1850,N_696);
nand U2075 (N_2075,In_729,In_1122);
nand U2076 (N_2076,N_1369,N_1362);
or U2077 (N_2077,In_3919,In_4710);
xor U2078 (N_2078,In_4904,N_1932);
nor U2079 (N_2079,In_3912,N_1707);
nand U2080 (N_2080,In_559,In_573);
nor U2081 (N_2081,In_4214,In_4719);
and U2082 (N_2082,N_364,N_149);
nor U2083 (N_2083,In_3972,In_293);
nor U2084 (N_2084,In_3035,In_4260);
nand U2085 (N_2085,N_596,In_1243);
and U2086 (N_2086,In_1633,In_1892);
and U2087 (N_2087,N_1089,N_1220);
nor U2088 (N_2088,In_1733,N_1545);
and U2089 (N_2089,In_3859,N_1432);
nand U2090 (N_2090,N_1652,In_3541);
nor U2091 (N_2091,In_809,N_402);
nor U2092 (N_2092,In_1405,In_1777);
or U2093 (N_2093,In_1675,In_2868);
or U2094 (N_2094,In_2896,In_1960);
nand U2095 (N_2095,In_3929,In_3476);
nand U2096 (N_2096,In_1822,N_611);
xor U2097 (N_2097,N_991,In_868);
nand U2098 (N_2098,N_1801,In_4795);
xor U2099 (N_2099,N_1021,In_2517);
nand U2100 (N_2100,N_1899,In_1444);
or U2101 (N_2101,N_1811,In_2213);
xor U2102 (N_2102,N_1093,In_1973);
nor U2103 (N_2103,In_3058,In_2487);
and U2104 (N_2104,N_229,In_2659);
nand U2105 (N_2105,N_1381,In_2966);
and U2106 (N_2106,In_3845,In_742);
or U2107 (N_2107,In_18,In_3371);
nand U2108 (N_2108,N_504,In_3209);
nor U2109 (N_2109,N_992,In_1596);
nor U2110 (N_2110,In_1766,N_243);
and U2111 (N_2111,N_1841,In_1501);
or U2112 (N_2112,N_565,In_207);
and U2113 (N_2113,N_1623,In_4738);
xnor U2114 (N_2114,In_3347,N_692);
nor U2115 (N_2115,In_3798,In_3810);
nand U2116 (N_2116,In_2079,N_1287);
or U2117 (N_2117,In_430,In_1711);
and U2118 (N_2118,N_1077,In_1583);
xnor U2119 (N_2119,In_4012,N_1833);
nand U2120 (N_2120,N_1948,N_1834);
or U2121 (N_2121,N_1379,N_1257);
and U2122 (N_2122,N_1107,In_3360);
or U2123 (N_2123,In_4612,In_1504);
nor U2124 (N_2124,N_441,N_1716);
xor U2125 (N_2125,N_1109,In_3582);
and U2126 (N_2126,N_502,In_1593);
and U2127 (N_2127,In_3865,In_3012);
nor U2128 (N_2128,N_237,N_1336);
nor U2129 (N_2129,In_3658,In_4718);
nand U2130 (N_2130,N_1263,In_668);
nand U2131 (N_2131,N_1041,In_1513);
and U2132 (N_2132,In_2838,N_1854);
nand U2133 (N_2133,In_588,N_979);
and U2134 (N_2134,In_32,In_3026);
or U2135 (N_2135,N_1182,In_1602);
nor U2136 (N_2136,In_3788,In_4042);
and U2137 (N_2137,N_1510,In_1383);
or U2138 (N_2138,In_3156,In_1419);
or U2139 (N_2139,N_1281,N_1315);
nand U2140 (N_2140,In_3568,In_587);
nor U2141 (N_2141,N_1420,In_1978);
and U2142 (N_2142,In_3433,N_1871);
nand U2143 (N_2143,N_1945,N_1410);
nand U2144 (N_2144,In_2760,In_4498);
or U2145 (N_2145,N_1761,N_878);
and U2146 (N_2146,In_3378,In_2855);
and U2147 (N_2147,N_420,N_1980);
nor U2148 (N_2148,In_2126,In_4784);
and U2149 (N_2149,In_1163,In_4224);
nor U2150 (N_2150,In_1519,N_1608);
nand U2151 (N_2151,N_1587,In_4629);
xor U2152 (N_2152,In_119,N_1823);
nand U2153 (N_2153,In_815,In_2931);
or U2154 (N_2154,N_759,N_1442);
and U2155 (N_2155,In_1455,In_666);
nand U2156 (N_2156,In_1103,In_2917);
and U2157 (N_2157,In_4526,N_1240);
nand U2158 (N_2158,N_1951,In_3136);
nor U2159 (N_2159,In_4845,N_756);
nor U2160 (N_2160,N_1343,In_1678);
or U2161 (N_2161,N_1997,N_984);
and U2162 (N_2162,In_4477,In_3794);
or U2163 (N_2163,In_1714,In_3995);
or U2164 (N_2164,N_371,In_143);
and U2165 (N_2165,N_339,N_857);
nor U2166 (N_2166,N_1836,In_4610);
or U2167 (N_2167,In_2935,N_466);
nand U2168 (N_2168,In_2916,In_2571);
or U2169 (N_2169,N_1011,In_4774);
nand U2170 (N_2170,N_1413,In_4899);
or U2171 (N_2171,In_2812,In_446);
and U2172 (N_2172,In_2684,In_4329);
or U2173 (N_2173,In_1411,In_3406);
and U2174 (N_2174,In_447,In_2138);
and U2175 (N_2175,In_3721,In_846);
nand U2176 (N_2176,N_102,N_1935);
or U2177 (N_2177,In_983,N_1838);
nor U2178 (N_2178,In_1130,In_2729);
or U2179 (N_2179,In_593,N_1807);
xnor U2180 (N_2180,In_933,N_148);
and U2181 (N_2181,N_1888,In_4714);
nand U2182 (N_2182,N_1332,In_4481);
xor U2183 (N_2183,In_802,In_1750);
and U2184 (N_2184,In_2089,In_1915);
nor U2185 (N_2185,In_2300,In_1902);
nand U2186 (N_2186,In_3072,In_774);
nand U2187 (N_2187,N_1931,In_899);
nand U2188 (N_2188,In_3828,N_1141);
xnor U2189 (N_2189,In_3870,In_233);
and U2190 (N_2190,N_1715,N_1015);
and U2191 (N_2191,N_1357,In_3815);
xnor U2192 (N_2192,N_1084,In_354);
or U2193 (N_2193,In_4153,N_851);
nand U2194 (N_2194,N_1588,In_4023);
nand U2195 (N_2195,N_909,In_2756);
nor U2196 (N_2196,N_1119,In_104);
xnor U2197 (N_2197,In_4000,In_330);
nand U2198 (N_2198,N_1008,N_663);
and U2199 (N_2199,In_1320,N_1903);
or U2200 (N_2200,In_4752,In_3518);
nand U2201 (N_2201,In_2681,In_2683);
nand U2202 (N_2202,In_4170,In_901);
xor U2203 (N_2203,In_2779,In_1955);
or U2204 (N_2204,In_1737,In_2985);
xor U2205 (N_2205,In_4455,N_1725);
nor U2206 (N_2206,N_1827,N_489);
and U2207 (N_2207,In_1278,N_530);
xor U2208 (N_2208,In_3746,N_1977);
nand U2209 (N_2209,In_3993,N_1018);
nand U2210 (N_2210,In_1207,In_2053);
xnor U2211 (N_2211,In_3778,In_746);
and U2212 (N_2212,In_1281,N_743);
xor U2213 (N_2213,In_816,N_1028);
xnor U2214 (N_2214,In_4108,N_1180);
and U2215 (N_2215,In_1286,N_1893);
nor U2216 (N_2216,N_1353,N_1847);
nor U2217 (N_2217,In_4320,In_4020);
xor U2218 (N_2218,N_579,In_4174);
nor U2219 (N_2219,In_3188,In_347);
xnor U2220 (N_2220,In_2880,In_3);
nor U2221 (N_2221,In_1125,N_1007);
and U2222 (N_2222,N_1145,In_2781);
and U2223 (N_2223,In_2972,In_4265);
or U2224 (N_2224,N_1268,In_4113);
nand U2225 (N_2225,N_275,N_1218);
or U2226 (N_2226,N_156,N_870);
nand U2227 (N_2227,In_760,In_2386);
xnor U2228 (N_2228,N_1605,N_1690);
nor U2229 (N_2229,In_672,N_1466);
xor U2230 (N_2230,In_1314,N_533);
nor U2231 (N_2231,N_202,In_3851);
and U2232 (N_2232,N_1778,In_602);
and U2233 (N_2233,N_1555,In_4589);
nor U2234 (N_2234,N_1500,N_1788);
nor U2235 (N_2235,In_3725,In_3861);
nor U2236 (N_2236,N_627,N_542);
and U2237 (N_2237,N_714,In_4847);
nor U2238 (N_2238,In_3444,In_2290);
xnor U2239 (N_2239,N_1583,In_3335);
and U2240 (N_2240,N_1507,In_4347);
nor U2241 (N_2241,In_1190,In_1869);
xor U2242 (N_2242,N_1908,N_581);
and U2243 (N_2243,N_812,In_1151);
and U2244 (N_2244,N_34,N_1038);
and U2245 (N_2245,In_3806,N_41);
or U2246 (N_2246,In_3652,N_1907);
nor U2247 (N_2247,In_680,In_835);
nand U2248 (N_2248,In_2786,N_1247);
and U2249 (N_2249,N_1926,In_1510);
and U2250 (N_2250,In_3067,In_622);
and U2251 (N_2251,N_1575,N_2074);
nor U2252 (N_2252,In_591,In_1491);
xnor U2253 (N_2253,In_1142,In_1211);
xor U2254 (N_2254,In_736,In_3415);
and U2255 (N_2255,N_130,N_2177);
xnor U2256 (N_2256,N_807,In_4452);
and U2257 (N_2257,N_797,In_1523);
nand U2258 (N_2258,In_4054,N_1938);
nor U2259 (N_2259,In_160,In_4864);
or U2260 (N_2260,N_654,In_1701);
and U2261 (N_2261,N_1522,N_556);
nand U2262 (N_2262,In_1991,N_2136);
xnor U2263 (N_2263,In_2525,In_3540);
or U2264 (N_2264,N_2217,N_2001);
nor U2265 (N_2265,N_927,In_1587);
nand U2266 (N_2266,N_1524,N_1430);
and U2267 (N_2267,N_726,In_3157);
nand U2268 (N_2268,In_1182,N_662);
nor U2269 (N_2269,N_1738,N_1447);
nor U2270 (N_2270,N_538,N_874);
nor U2271 (N_2271,In_3352,In_2646);
xor U2272 (N_2272,N_391,N_1239);
nor U2273 (N_2273,In_2584,N_1849);
xnor U2274 (N_2274,In_2385,In_3158);
nor U2275 (N_2275,N_1960,N_1901);
nand U2276 (N_2276,N_2085,N_2191);
xor U2277 (N_2277,In_1563,N_529);
nor U2278 (N_2278,N_2189,In_3768);
or U2279 (N_2279,N_1488,In_3283);
or U2280 (N_2280,N_2205,N_1134);
nor U2281 (N_2281,In_397,In_1705);
xor U2282 (N_2282,N_427,N_2105);
and U2283 (N_2283,N_1174,In_1134);
nor U2284 (N_2284,In_3942,In_4565);
nor U2285 (N_2285,N_2117,N_1518);
xor U2286 (N_2286,In_4137,In_1319);
nand U2287 (N_2287,In_3328,N_2130);
nand U2288 (N_2288,In_2033,In_3361);
nand U2289 (N_2289,In_4348,N_1837);
or U2290 (N_2290,N_1421,In_4950);
xnor U2291 (N_2291,In_3402,N_39);
xnor U2292 (N_2292,In_2018,N_1264);
and U2293 (N_2293,In_275,In_3962);
and U2294 (N_2294,N_1813,N_1800);
nor U2295 (N_2295,N_1394,N_81);
and U2296 (N_2296,In_1227,In_1145);
or U2297 (N_2297,N_1673,N_1056);
nor U2298 (N_2298,N_1506,In_1105);
and U2299 (N_2299,In_3499,N_1292);
nor U2300 (N_2300,N_1552,In_1461);
xor U2301 (N_2301,N_1428,N_1437);
nand U2302 (N_2302,N_1644,In_1689);
nor U2303 (N_2303,N_1700,N_473);
or U2304 (N_2304,N_1636,In_1691);
xor U2305 (N_2305,N_867,In_4631);
or U2306 (N_2306,N_2185,In_417);
or U2307 (N_2307,N_2183,In_3131);
nor U2308 (N_2308,In_3142,In_764);
xor U2309 (N_2309,N_2099,N_1774);
xor U2310 (N_2310,In_980,N_2152);
or U2311 (N_2311,In_245,In_3751);
xnor U2312 (N_2312,N_510,N_2089);
or U2313 (N_2313,In_1760,In_4311);
or U2314 (N_2314,In_2814,In_4393);
or U2315 (N_2315,In_2716,In_2303);
xor U2316 (N_2316,N_170,N_988);
xnor U2317 (N_2317,In_3114,N_1744);
nand U2318 (N_2318,In_2625,In_1776);
xor U2319 (N_2319,N_1062,N_1396);
nand U2320 (N_2320,N_1934,In_202);
nor U2321 (N_2321,N_2014,In_173);
and U2322 (N_2322,In_1875,N_147);
nor U2323 (N_2323,In_1453,N_414);
nand U2324 (N_2324,In_2648,In_1267);
nor U2325 (N_2325,In_4052,N_1835);
xor U2326 (N_2326,In_4748,N_2199);
nand U2327 (N_2327,N_346,N_2013);
nor U2328 (N_2328,In_1525,In_1634);
nand U2329 (N_2329,In_1601,N_1472);
nand U2330 (N_2330,N_1324,In_479);
nand U2331 (N_2331,N_985,In_4615);
nand U2332 (N_2332,In_3896,N_1958);
nor U2333 (N_2333,In_1486,N_1228);
xor U2334 (N_2334,N_385,N_2035);
nand U2335 (N_2335,N_948,N_1540);
and U2336 (N_2336,N_2087,N_2135);
xor U2337 (N_2337,In_450,In_1231);
nor U2338 (N_2338,In_3624,N_2248);
or U2339 (N_2339,N_1734,In_3454);
xnor U2340 (N_2340,In_2614,N_1252);
and U2341 (N_2341,N_2129,N_1201);
or U2342 (N_2342,N_543,N_1614);
or U2343 (N_2343,In_4569,N_2194);
xnor U2344 (N_2344,N_1390,N_1897);
xnor U2345 (N_2345,N_1185,N_1241);
xnor U2346 (N_2346,In_3581,N_1805);
xnor U2347 (N_2347,In_704,In_3952);
nand U2348 (N_2348,In_3113,N_829);
and U2349 (N_2349,N_1895,In_3641);
or U2350 (N_2350,N_625,In_4799);
or U2351 (N_2351,In_4479,In_353);
and U2352 (N_2352,In_4559,In_1906);
nand U2353 (N_2353,N_1645,In_3353);
nand U2354 (N_2354,In_55,N_907);
xnor U2355 (N_2355,N_1721,N_305);
and U2356 (N_2356,In_3321,In_4474);
nand U2357 (N_2357,In_4655,N_1403);
nor U2358 (N_2358,In_2068,N_2180);
xnor U2359 (N_2359,In_4785,In_242);
and U2360 (N_2360,In_2098,In_3864);
nand U2361 (N_2361,N_527,N_1189);
and U2362 (N_2362,In_3237,N_135);
and U2363 (N_2363,N_349,In_21);
xor U2364 (N_2364,In_4547,N_1952);
nor U2365 (N_2365,N_2204,N_2000);
nor U2366 (N_2366,In_1668,N_2081);
or U2367 (N_2367,N_228,N_559);
nand U2368 (N_2368,N_2019,In_2664);
nand U2369 (N_2369,In_4296,N_1169);
and U2370 (N_2370,In_975,In_4425);
nor U2371 (N_2371,In_4813,In_267);
xor U2372 (N_2372,N_2114,In_2404);
nand U2373 (N_2373,N_2095,N_2169);
xor U2374 (N_2374,N_1194,N_2032);
nor U2375 (N_2375,N_1066,N_941);
and U2376 (N_2376,In_797,In_2413);
xnor U2377 (N_2377,N_1680,In_4306);
nand U2378 (N_2378,N_649,In_4223);
or U2379 (N_2379,N_2025,In_4237);
nand U2380 (N_2380,N_1525,In_795);
nor U2381 (N_2381,In_3750,N_1753);
or U2382 (N_2382,N_1033,N_92);
nand U2383 (N_2383,N_1814,In_2012);
nor U2384 (N_2384,N_1929,N_1946);
or U2385 (N_2385,In_117,N_321);
nor U2386 (N_2386,In_1119,N_1772);
xor U2387 (N_2387,N_1820,In_2807);
xnor U2388 (N_2388,In_884,N_2140);
xnor U2389 (N_2389,N_1016,In_4471);
nand U2390 (N_2390,N_890,In_1562);
xnor U2391 (N_2391,In_543,In_698);
nand U2392 (N_2392,N_1493,N_1822);
nor U2393 (N_2393,N_1630,N_134);
nand U2394 (N_2394,N_1491,N_2149);
and U2395 (N_2395,In_633,In_4948);
xnor U2396 (N_2396,In_4811,N_1328);
nor U2397 (N_2397,N_571,In_4378);
xor U2398 (N_2398,N_1334,In_355);
nand U2399 (N_2399,In_3906,N_1311);
xor U2400 (N_2400,In_865,N_670);
and U2401 (N_2401,In_4997,N_2064);
nand U2402 (N_2402,N_1770,In_2757);
or U2403 (N_2403,In_2134,In_1665);
xnor U2404 (N_2404,In_1219,In_147);
nor U2405 (N_2405,In_1235,In_1335);
nor U2406 (N_2406,N_784,N_1179);
xor U2407 (N_2407,N_163,In_599);
nor U2408 (N_2408,N_678,N_632);
nand U2409 (N_2409,In_2465,In_4419);
nor U2410 (N_2410,N_1553,In_465);
or U2411 (N_2411,In_1594,N_18);
nand U2412 (N_2412,In_2750,In_1819);
or U2413 (N_2413,N_1592,N_59);
nand U2414 (N_2414,N_1363,N_2009);
xor U2415 (N_2415,In_4157,N_2123);
and U2416 (N_2416,In_1030,In_2412);
nand U2417 (N_2417,In_3804,N_1676);
nand U2418 (N_2418,In_1042,N_2226);
and U2419 (N_2419,N_694,In_1840);
or U2420 (N_2420,N_1333,In_1221);
nand U2421 (N_2421,In_3645,In_1644);
nand U2422 (N_2422,In_4395,In_1866);
nand U2423 (N_2423,N_1408,N_1283);
xor U2424 (N_2424,In_4989,In_4377);
nor U2425 (N_2425,N_2178,In_2598);
and U2426 (N_2426,In_2428,In_1942);
or U2427 (N_2427,In_3032,In_4361);
xor U2428 (N_2428,In_1390,N_2084);
or U2429 (N_2429,N_1708,N_1855);
nor U2430 (N_2430,N_1411,In_4288);
and U2431 (N_2431,N_1156,In_4386);
nand U2432 (N_2432,N_1984,In_3178);
or U2433 (N_2433,In_4509,N_1463);
nand U2434 (N_2434,In_1893,In_4205);
nor U2435 (N_2435,In_2060,N_2246);
and U2436 (N_2436,N_450,In_1425);
nor U2437 (N_2437,In_1066,In_73);
xor U2438 (N_2438,In_1387,N_2125);
and U2439 (N_2439,N_1848,In_4285);
and U2440 (N_2440,In_3348,In_670);
nor U2441 (N_2441,N_2154,N_352);
nor U2442 (N_2442,N_215,In_3311);
and U2443 (N_2443,In_2246,In_2792);
nand U2444 (N_2444,N_424,N_1113);
or U2445 (N_2445,In_4200,N_1976);
nor U2446 (N_2446,In_3478,In_3213);
and U2447 (N_2447,In_3921,N_2156);
xor U2448 (N_2448,N_1039,In_2568);
nor U2449 (N_2449,In_1298,In_2209);
or U2450 (N_2450,In_3979,In_2410);
and U2451 (N_2451,In_4212,N_290);
xnor U2452 (N_2452,N_2029,In_2011);
xnor U2453 (N_2453,N_2175,In_3098);
nor U2454 (N_2454,In_4742,N_1142);
nor U2455 (N_2455,In_1384,In_2824);
and U2456 (N_2456,In_4654,In_468);
and U2457 (N_2457,In_165,N_234);
or U2458 (N_2458,N_1740,N_1265);
nand U2459 (N_2459,In_870,In_3644);
xor U2460 (N_2460,In_2673,In_3445);
and U2461 (N_2461,N_859,In_6);
and U2462 (N_2462,In_156,N_1961);
and U2463 (N_2463,N_203,In_1867);
and U2464 (N_2464,N_1758,In_2167);
xnor U2465 (N_2465,In_3408,In_3204);
nand U2466 (N_2466,In_3547,In_4018);
xnor U2467 (N_2467,In_918,N_1501);
or U2468 (N_2468,In_720,N_1534);
or U2469 (N_2469,In_1863,N_573);
nand U2470 (N_2470,In_1426,N_2003);
nor U2471 (N_2471,N_2102,N_1221);
or U2472 (N_2472,N_2060,In_4840);
nand U2473 (N_2473,In_3465,In_755);
xor U2474 (N_2474,In_1364,N_1628);
or U2475 (N_2475,In_2453,In_381);
nand U2476 (N_2476,In_2899,N_1081);
nor U2477 (N_2477,In_1133,In_4897);
xnor U2478 (N_2478,N_487,N_1521);
xor U2479 (N_2479,In_2892,N_1384);
nor U2480 (N_2480,N_1991,In_3843);
nor U2481 (N_2481,In_1489,In_3184);
nor U2482 (N_2482,In_4501,In_3908);
or U2483 (N_2483,In_1240,In_2191);
xor U2484 (N_2484,N_139,In_2052);
and U2485 (N_2485,N_288,In_4072);
nor U2486 (N_2486,In_1859,N_1078);
or U2487 (N_2487,In_3376,N_1259);
nor U2488 (N_2488,In_4636,N_1242);
nor U2489 (N_2489,N_1978,In_2496);
nand U2490 (N_2490,In_627,In_2074);
xnor U2491 (N_2491,In_3710,N_1269);
nand U2492 (N_2492,In_789,N_1232);
nor U2493 (N_2493,In_4032,N_598);
and U2494 (N_2494,In_2374,N_1613);
and U2495 (N_2495,In_1782,N_1143);
or U2496 (N_2496,In_1770,N_29);
nand U2497 (N_2497,In_1828,N_1128);
and U2498 (N_2498,N_1370,N_236);
or U2499 (N_2499,In_536,N_1124);
nor U2500 (N_2500,N_2356,N_1794);
nand U2501 (N_2501,In_2867,N_2453);
nand U2502 (N_2502,In_2712,N_2491);
xor U2503 (N_2503,N_2015,In_782);
or U2504 (N_2504,In_2347,N_1968);
or U2505 (N_2505,N_2450,In_3481);
nor U2506 (N_2506,N_436,N_1458);
and U2507 (N_2507,N_987,In_1106);
nand U2508 (N_2508,N_1036,N_2227);
nand U2509 (N_2509,In_1417,N_2238);
xor U2510 (N_2510,N_1659,N_298);
xnor U2511 (N_2511,N_1559,N_2466);
nand U2512 (N_2512,In_4411,N_2258);
nor U2513 (N_2513,In_2799,In_2423);
nor U2514 (N_2514,N_2254,N_886);
and U2515 (N_2515,In_1479,N_432);
nand U2516 (N_2516,In_2297,N_771);
or U2517 (N_2517,N_2002,In_3482);
nand U2518 (N_2518,In_3299,In_1784);
nor U2519 (N_2519,N_2239,In_4827);
or U2520 (N_2520,In_1951,N_1027);
nor U2521 (N_2521,In_4036,N_388);
nand U2522 (N_2522,In_2651,N_2173);
nand U2523 (N_2523,In_2409,In_1418);
and U2524 (N_2524,N_1515,N_1930);
nand U2525 (N_2525,N_2285,In_2754);
xor U2526 (N_2526,N_2352,In_4095);
nand U2527 (N_2527,N_1994,N_1498);
nor U2528 (N_2528,N_1293,N_1565);
or U2529 (N_2529,N_1925,In_2527);
and U2530 (N_2530,N_2324,N_440);
nand U2531 (N_2531,In_2869,In_4445);
nand U2532 (N_2532,N_725,N_1508);
nor U2533 (N_2533,In_2652,N_2030);
and U2534 (N_2534,N_2122,In_3551);
nor U2535 (N_2535,In_4725,N_329);
or U2536 (N_2536,N_898,In_553);
and U2537 (N_2537,N_1872,In_997);
and U2538 (N_2538,In_276,In_4716);
xor U2539 (N_2539,N_2245,In_2137);
nor U2540 (N_2540,N_1860,N_88);
xor U2541 (N_2541,In_3160,N_942);
xor U2542 (N_2542,In_4353,N_2444);
nor U2543 (N_2543,In_565,N_25);
nor U2544 (N_2544,In_1059,N_2400);
or U2545 (N_2545,In_1309,N_1859);
or U2546 (N_2546,N_1789,N_2415);
and U2547 (N_2547,N_826,N_1919);
and U2548 (N_2548,N_1320,N_1812);
nand U2549 (N_2549,N_842,N_2265);
xor U2550 (N_2550,In_4397,N_1999);
and U2551 (N_2551,In_1352,N_2335);
nor U2552 (N_2552,N_796,N_1917);
xnor U2553 (N_2553,In_836,In_2232);
and U2554 (N_2554,N_908,In_3097);
and U2555 (N_2555,N_2157,N_1325);
xor U2556 (N_2556,N_569,In_1306);
or U2557 (N_2557,In_699,N_1618);
nand U2558 (N_2558,In_1463,N_1691);
and U2559 (N_2559,N_1199,N_1391);
nand U2560 (N_2560,In_2624,In_2704);
and U2561 (N_2561,In_1055,In_3162);
and U2562 (N_2562,N_250,N_2004);
nor U2563 (N_2563,N_861,N_1776);
or U2564 (N_2564,N_1748,N_2027);
nand U2565 (N_2565,In_1047,In_1205);
or U2566 (N_2566,In_957,In_2724);
xor U2567 (N_2567,In_4219,In_643);
or U2568 (N_2568,N_2100,N_637);
xor U2569 (N_2569,N_261,In_1571);
and U2570 (N_2570,In_2162,In_4025);
or U2571 (N_2571,In_340,In_223);
nor U2572 (N_2572,N_2341,In_4735);
nor U2573 (N_2573,N_1729,N_1955);
nand U2574 (N_2574,In_4103,N_2369);
or U2575 (N_2575,In_4892,In_1713);
and U2576 (N_2576,N_1722,In_4240);
nand U2577 (N_2577,In_1584,In_167);
nor U2578 (N_2578,N_2336,In_320);
or U2579 (N_2579,In_875,In_257);
xnor U2580 (N_2580,In_1741,N_2346);
nand U2581 (N_2581,N_718,In_3685);
nand U2582 (N_2582,In_2499,N_1879);
xor U2583 (N_2583,N_1863,N_145);
nor U2584 (N_2584,In_2613,N_967);
or U2585 (N_2585,In_3945,In_1817);
nor U2586 (N_2586,In_3083,In_3643);
nand U2587 (N_2587,In_4776,In_4571);
and U2588 (N_2588,In_947,In_4440);
nor U2589 (N_2589,In_1907,In_2721);
xnor U2590 (N_2590,N_2124,N_1153);
or U2591 (N_2591,In_974,N_740);
nand U2592 (N_2592,In_1774,N_334);
and U2593 (N_2593,N_672,N_700);
xnor U2594 (N_2594,N_2387,N_2448);
nand U2595 (N_2595,In_2234,N_939);
and U2596 (N_2596,In_3356,N_1887);
nor U2597 (N_2597,N_626,N_920);
nand U2598 (N_2598,In_1223,In_174);
and U2599 (N_2599,In_3871,N_2273);
xnor U2600 (N_2600,N_86,In_425);
or U2601 (N_2601,N_2291,N_296);
xor U2602 (N_2602,N_2390,N_1532);
nor U2603 (N_2603,In_3101,N_1448);
and U2604 (N_2604,N_1471,In_4941);
xnor U2605 (N_2605,N_2306,In_1433);
nand U2606 (N_2606,N_1718,In_3941);
nand U2607 (N_2607,In_4762,In_2689);
and U2608 (N_2608,In_740,N_2458);
nand U2609 (N_2609,In_4720,In_3015);
or U2610 (N_2610,In_1197,In_2767);
or U2611 (N_2611,N_1650,In_1687);
nor U2612 (N_2612,N_2398,N_810);
nand U2613 (N_2613,N_2112,In_2644);
xnor U2614 (N_2614,In_3809,N_2385);
xnor U2615 (N_2615,N_1760,In_1690);
and U2616 (N_2616,In_1408,N_219);
or U2617 (N_2617,In_829,N_2311);
nand U2618 (N_2618,In_1746,In_3043);
nand U2619 (N_2619,In_1194,N_2063);
nand U2620 (N_2620,N_728,In_3884);
and U2621 (N_2621,N_1889,In_1708);
nand U2622 (N_2622,In_1075,In_2858);
nand U2623 (N_2623,In_159,N_1051);
xor U2624 (N_2624,N_2126,N_1797);
xnor U2625 (N_2625,N_2277,In_4270);
nor U2626 (N_2626,N_2022,N_1121);
and U2627 (N_2627,N_2388,N_1828);
or U2628 (N_2628,N_1484,In_2046);
or U2629 (N_2629,In_15,N_792);
xor U2630 (N_2630,In_4878,N_2434);
nand U2631 (N_2631,N_2452,In_2609);
xor U2632 (N_2632,N_1285,N_1237);
or U2633 (N_2633,In_3268,N_2193);
xor U2634 (N_2634,In_4849,N_2427);
xor U2635 (N_2635,N_2481,N_1617);
nand U2636 (N_2636,In_609,N_1658);
or U2637 (N_2637,N_1661,In_4374);
or U2638 (N_2638,N_1564,N_1465);
nand U2639 (N_2639,In_2364,N_2429);
and U2640 (N_2640,N_1861,N_1407);
or U2641 (N_2641,N_350,N_2143);
nand U2642 (N_2642,N_1795,In_678);
xor U2643 (N_2643,N_2413,N_2323);
and U2644 (N_2644,N_2109,N_1631);
or U2645 (N_2645,In_3981,In_1887);
or U2646 (N_2646,N_1910,N_2409);
xor U2647 (N_2647,N_1042,N_1025);
or U2648 (N_2648,In_4133,N_2068);
nor U2649 (N_2649,In_4268,In_359);
nand U2650 (N_2650,N_2280,N_2276);
and U2651 (N_2651,N_2184,N_1874);
nor U2652 (N_2652,In_4730,In_244);
and U2653 (N_2653,N_2467,In_4674);
and U2654 (N_2654,N_1906,In_3626);
nor U2655 (N_2655,In_1943,In_1976);
or U2656 (N_2656,N_2282,In_4026);
nor U2657 (N_2657,In_1526,In_685);
and U2658 (N_2658,In_3825,In_1401);
or U2659 (N_2659,N_1401,N_2475);
nand U2660 (N_2660,In_981,N_1344);
or U2661 (N_2661,N_1576,In_3927);
nand U2662 (N_2662,In_2968,In_4646);
nor U2663 (N_2663,In_707,N_576);
and U2664 (N_2664,N_2377,In_987);
nor U2665 (N_2665,N_1452,N_962);
or U2666 (N_2666,In_2973,In_1269);
nand U2667 (N_2667,N_2331,In_3762);
nand U2668 (N_2668,N_2329,N_1271);
xnor U2669 (N_2669,N_2138,In_1017);
or U2670 (N_2670,N_2462,In_780);
or U2671 (N_2671,In_190,In_106);
or U2672 (N_2672,N_1857,In_1367);
nand U2673 (N_2673,In_3459,In_371);
or U2674 (N_2674,N_2382,In_3933);
and U2675 (N_2675,In_2151,N_1400);
xnor U2676 (N_2676,In_3227,In_3646);
or U2677 (N_2677,N_1773,In_1597);
or U2678 (N_2678,N_2086,N_6);
or U2679 (N_2679,N_1816,In_1376);
nand U2680 (N_2680,N_2098,N_1331);
or U2681 (N_2681,In_3259,In_4244);
and U2682 (N_2682,N_1747,In_3575);
or U2683 (N_2683,In_1074,In_3720);
nor U2684 (N_2684,In_709,In_2420);
or U2685 (N_2685,N_1453,In_476);
xnor U2686 (N_2686,In_3914,N_2288);
xnor U2687 (N_2687,In_3410,N_929);
xor U2688 (N_2688,N_1178,In_822);
xor U2689 (N_2689,N_1595,In_3611);
nand U2690 (N_2690,In_2013,In_3830);
xor U2691 (N_2691,N_2174,N_2250);
and U2692 (N_2692,N_2223,In_3366);
or U2693 (N_2693,In_4322,N_2110);
nor U2694 (N_2694,N_868,In_516);
xnor U2695 (N_2695,N_2165,In_2239);
xor U2696 (N_2696,N_597,N_2459);
or U2697 (N_2697,In_4074,N_2023);
nor U2698 (N_2698,N_1743,N_2113);
or U2699 (N_2699,N_1533,In_4369);
nor U2700 (N_2700,In_3700,N_1724);
and U2701 (N_2701,In_1464,N_1845);
or U2702 (N_2702,N_2411,N_2101);
xnor U2703 (N_2703,N_2431,N_90);
and U2704 (N_2704,N_2182,N_2375);
xnor U2705 (N_2705,In_2885,In_4818);
or U2706 (N_2706,In_2367,N_1203);
or U2707 (N_2707,In_86,In_3516);
nand U2708 (N_2708,N_2225,In_4);
or U2709 (N_2709,In_3070,In_1896);
nor U2710 (N_2710,In_83,N_2202);
or U2711 (N_2711,In_230,N_2386);
nor U2712 (N_2712,N_1941,In_2526);
nand U2713 (N_2713,In_2679,N_1677);
or U2714 (N_2714,N_1864,N_2186);
and U2715 (N_2715,In_298,N_2269);
or U2716 (N_2716,In_2967,N_656);
nor U2717 (N_2717,In_1111,In_2629);
nand U2718 (N_2718,In_3432,N_2111);
nor U2719 (N_2719,N_2487,In_4467);
and U2720 (N_2720,N_2456,In_611);
nand U2721 (N_2721,N_1714,N_2091);
xor U2722 (N_2722,N_2039,N_1582);
nand U2723 (N_2723,N_2044,N_133);
nand U2724 (N_2724,N_2404,In_51);
nor U2725 (N_2725,In_3224,In_2839);
or U2726 (N_2726,In_4062,In_2372);
or U2727 (N_2727,N_1654,N_2082);
nand U2728 (N_2728,N_2144,In_2448);
xor U2729 (N_2729,In_4707,N_1250);
xnor U2730 (N_2730,In_2342,In_2362);
nand U2731 (N_2731,In_3699,In_494);
nor U2732 (N_2732,In_195,In_3656);
nand U2733 (N_2733,N_1052,N_2399);
nor U2734 (N_2734,In_454,In_1247);
nor U2735 (N_2735,N_1986,N_2120);
xnor U2736 (N_2736,In_4949,N_729);
and U2737 (N_2737,N_1070,In_2811);
nor U2738 (N_2738,In_3642,In_3451);
nand U2739 (N_2739,In_2442,In_1821);
nor U2740 (N_2740,In_1060,N_2041);
xnor U2741 (N_2741,N_1548,N_1529);
nor U2742 (N_2742,N_1023,N_1790);
or U2743 (N_2743,N_2275,In_4182);
xnor U2744 (N_2744,In_3165,N_1829);
nand U2745 (N_2745,In_484,In_2660);
and U2746 (N_2746,N_2121,In_649);
nand U2747 (N_2747,In_3192,N_1815);
xnor U2748 (N_2748,N_2485,In_2265);
nor U2749 (N_2749,N_1418,N_27);
nand U2750 (N_2750,In_708,In_76);
or U2751 (N_2751,In_4309,N_2441);
nor U2752 (N_2752,N_993,N_1878);
or U2753 (N_2753,In_3730,In_1378);
and U2754 (N_2754,In_3556,N_2058);
nand U2755 (N_2755,In_3511,In_4858);
or U2756 (N_2756,N_2052,In_2690);
or U2757 (N_2757,In_2195,In_2854);
and U2758 (N_2758,N_2158,In_108);
xnor U2759 (N_2759,In_4908,In_3885);
nand U2760 (N_2760,N_956,In_1191);
and U2761 (N_2761,N_1358,N_2484);
or U2762 (N_2762,In_1682,N_657);
nand U2763 (N_2763,N_1563,In_4689);
xnor U2764 (N_2764,In_474,In_2432);
nand U2765 (N_2765,N_1710,In_3686);
nor U2766 (N_2766,N_972,N_91);
xor U2767 (N_2767,N_2694,N_2590);
and U2768 (N_2768,N_2264,N_2407);
or U2769 (N_2769,N_1288,N_128);
and U2770 (N_2770,N_2428,N_1513);
nand U2771 (N_2771,In_4782,N_459);
nor U2772 (N_2772,In_2996,In_4585);
xnor U2773 (N_2773,In_1121,N_1616);
nand U2774 (N_2774,N_1208,In_2680);
nor U2775 (N_2775,In_497,In_2172);
nor U2776 (N_2776,N_307,In_3449);
nor U2777 (N_2777,In_1480,In_255);
xor U2778 (N_2778,In_3143,In_2645);
xnor U2779 (N_2779,In_626,In_2444);
and U2780 (N_2780,In_727,In_4127);
nor U2781 (N_2781,N_2359,In_1389);
and U2782 (N_2782,N_2502,In_2069);
nand U2783 (N_2783,N_2176,In_2803);
nand U2784 (N_2784,In_909,N_425);
or U2785 (N_2785,In_1061,N_264);
nor U2786 (N_2786,In_3251,N_2435);
nor U2787 (N_2787,In_248,N_1193);
nand U2788 (N_2788,In_4460,N_2195);
or U2789 (N_2789,In_1069,N_2392);
or U2790 (N_2790,In_70,N_1176);
xnor U2791 (N_2791,N_2721,In_2253);
or U2792 (N_2792,In_4461,N_1840);
nor U2793 (N_2793,N_2119,N_2270);
and U2794 (N_2794,In_661,In_3472);
and U2795 (N_2795,In_4902,In_4515);
xor U2796 (N_2796,N_746,N_1920);
or U2797 (N_2797,In_1349,In_2243);
and U2798 (N_2798,In_3791,N_703);
xnor U2799 (N_2799,N_433,N_2639);
nor U2800 (N_2800,N_2445,N_1686);
or U2801 (N_2801,N_1996,N_1354);
or U2802 (N_2802,In_1922,N_2408);
nand U2803 (N_2803,N_2524,N_2543);
or U2804 (N_2804,In_2189,In_3716);
xor U2805 (N_2805,N_2433,In_403);
nand U2806 (N_2806,N_195,N_369);
xnor U2807 (N_2807,N_368,In_1160);
or U2808 (N_2808,In_1173,N_1187);
nor U2809 (N_2809,In_3286,In_4247);
or U2810 (N_2810,N_602,N_1558);
nand U2811 (N_2811,In_1619,N_1098);
and U2812 (N_2812,N_2351,N_1322);
and U2813 (N_2813,In_571,N_1438);
nor U2814 (N_2814,N_1364,N_1246);
or U2815 (N_2815,N_2598,N_2034);
nor U2816 (N_2816,N_1637,In_448);
nand U2817 (N_2817,N_2279,N_1387);
xor U2818 (N_2818,In_4859,N_1615);
nor U2819 (N_2819,N_418,In_2271);
nand U2820 (N_2820,N_1731,In_2863);
nor U2821 (N_2821,N_2446,N_1993);
and U2822 (N_2822,In_1727,N_2330);
nor U2823 (N_2823,In_4507,N_1001);
or U2824 (N_2824,In_3966,In_3601);
nor U2825 (N_2825,N_1061,In_4073);
and U2826 (N_2826,N_782,In_1410);
xnor U2827 (N_2827,N_2738,In_4132);
nor U2828 (N_2828,In_2186,N_2662);
nand U2829 (N_2829,N_924,N_2493);
nor U2830 (N_2830,In_871,In_828);
xnor U2831 (N_2831,N_2163,N_2710);
and U2832 (N_2832,N_1766,In_674);
and U2833 (N_2833,N_2142,N_818);
or U2834 (N_2834,N_2730,N_990);
or U2835 (N_2835,N_1866,N_1210);
or U2836 (N_2836,N_2078,In_3922);
or U2837 (N_2837,In_527,N_701);
nand U2838 (N_2838,N_2215,N_2332);
nor U2839 (N_2839,In_434,N_2553);
nor U2840 (N_2840,N_2641,In_4181);
nand U2841 (N_2841,N_2302,N_1017);
xnor U2842 (N_2842,In_523,In_2921);
xnor U2843 (N_2843,N_2558,N_1172);
and U2844 (N_2844,N_1940,N_186);
nor U2845 (N_2845,In_2320,In_4124);
or U2846 (N_2846,In_777,N_2286);
xor U2847 (N_2847,N_2213,N_764);
nand U2848 (N_2848,In_2365,N_2252);
xor U2849 (N_2849,N_2161,N_1277);
xor U2850 (N_2850,In_3455,N_1514);
or U2851 (N_2851,N_1939,N_2692);
nor U2852 (N_2852,N_1755,N_2010);
nor U2853 (N_2853,In_4220,N_2066);
xor U2854 (N_2854,In_4029,In_810);
and U2855 (N_2855,N_1399,N_2501);
and U2856 (N_2856,N_1964,In_4245);
and U2857 (N_2857,N_2372,In_4217);
nand U2858 (N_2858,In_4015,N_2537);
nand U2859 (N_2859,N_2097,In_3359);
and U2860 (N_2860,In_4815,N_2317);
nor U2861 (N_2861,In_3692,In_303);
xnor U2862 (N_2862,N_1116,N_911);
xor U2863 (N_2863,In_1001,In_1566);
xnor U2864 (N_2864,N_2056,In_915);
nor U2865 (N_2865,N_1883,In_984);
and U2866 (N_2866,In_4027,N_610);
nand U2867 (N_2867,N_1013,N_248);
nor U2868 (N_2868,N_1693,N_1412);
or U2869 (N_2869,In_1636,N_2495);
or U2870 (N_2870,N_879,In_64);
nand U2871 (N_2871,In_1311,In_3217);
nand U2872 (N_2872,In_1276,In_741);
and U2873 (N_2873,In_1325,N_2652);
xor U2874 (N_2874,N_1641,N_1745);
nor U2875 (N_2875,N_2560,In_59);
and U2876 (N_2876,N_2634,In_4401);
nand U2877 (N_2877,N_2043,In_1965);
nand U2878 (N_2878,In_2576,N_2251);
xor U2879 (N_2879,N_716,In_2695);
or U2880 (N_2880,N_1598,In_3081);
nor U2881 (N_2881,In_3577,In_3066);
nor U2882 (N_2882,N_2218,N_2548);
xnor U2883 (N_2883,N_1601,In_172);
and U2884 (N_2884,N_1664,N_1911);
xnor U2885 (N_2885,In_1393,N_902);
or U2886 (N_2886,In_3096,N_2221);
and U2887 (N_2887,N_1329,N_1768);
nand U2888 (N_2888,In_4179,N_1499);
nand U2889 (N_2889,N_278,N_2241);
and U2890 (N_2890,In_4952,In_754);
nor U2891 (N_2891,In_1366,N_772);
xor U2892 (N_2892,N_1300,In_4751);
nor U2893 (N_2893,N_172,In_4163);
or U2894 (N_2894,N_2625,In_2835);
or U2895 (N_2895,In_1805,In_281);
nor U2896 (N_2896,N_2532,In_824);
and U2897 (N_2897,N_2072,In_1801);
or U2898 (N_2898,In_2346,In_4324);
or U2899 (N_2899,N_896,In_1595);
and U2900 (N_2900,N_786,N_2608);
and U2901 (N_2901,N_377,In_2804);
or U2902 (N_2902,N_109,In_1224);
nor U2903 (N_2903,N_1902,N_345);
xnor U2904 (N_2904,In_180,In_3276);
nand U2905 (N_2905,In_890,In_2492);
and U2906 (N_2906,N_2305,In_4368);
nand U2907 (N_2907,N_2322,In_2160);
and U2908 (N_2908,In_2498,N_1435);
or U2909 (N_2909,In_2837,N_2059);
xor U2910 (N_2910,In_916,N_1254);
nor U2911 (N_2911,N_1290,N_2539);
nand U2912 (N_2912,N_1517,In_238);
and U2913 (N_2913,N_1983,In_2580);
xnor U2914 (N_2914,N_2362,N_2172);
nor U2915 (N_2915,N_2705,N_1780);
and U2916 (N_2916,N_2345,N_1249);
xnor U2917 (N_2917,N_1726,In_1388);
or U2918 (N_2918,In_1422,N_2300);
nand U2919 (N_2919,In_414,In_3565);
xnor U2920 (N_2920,In_1807,N_157);
xor U2921 (N_2921,N_191,N_328);
or U2922 (N_2922,N_2747,N_1653);
nand U2923 (N_2923,In_2566,In_134);
nand U2924 (N_2924,N_1985,In_1071);
and U2925 (N_2925,N_2545,In_2236);
and U2926 (N_2926,N_2519,In_3553);
nand U2927 (N_2927,In_1356,N_2374);
nand U2928 (N_2928,N_1427,N_2201);
and U2929 (N_2929,N_2531,In_3486);
xor U2930 (N_2930,N_2164,In_1016);
nor U2931 (N_2931,In_1196,N_635);
and U2932 (N_2932,In_2640,In_4891);
nand U2933 (N_2933,N_2723,N_1335);
nor U2934 (N_2934,In_2927,N_770);
xor U2935 (N_2935,In_30,In_600);
xnor U2936 (N_2936,In_3322,In_550);
xnor U2937 (N_2937,N_806,N_814);
nor U2938 (N_2938,N_193,N_1767);
or U2939 (N_2939,N_1088,N_2370);
or U2940 (N_2940,In_2832,N_2621);
xnor U2941 (N_2941,N_2197,N_2360);
and U2942 (N_2942,In_2913,N_2686);
nor U2943 (N_2943,In_4444,In_1841);
xor U2944 (N_2944,N_2512,In_2906);
and U2945 (N_2945,In_2459,In_4041);
or U2946 (N_2946,In_4577,In_1755);
nor U2947 (N_2947,N_697,N_2570);
nand U2948 (N_2948,In_2766,N_2660);
nor U2949 (N_2949,N_1922,N_499);
xnor U2950 (N_2950,In_4519,N_2339);
nor U2951 (N_2951,N_582,N_2671);
nor U2952 (N_2952,N_2083,N_1392);
or U2953 (N_2953,N_2650,N_2526);
nand U2954 (N_2954,N_2148,In_4695);
and U2955 (N_2955,In_2588,In_4228);
nor U2956 (N_2956,In_2009,N_1746);
xnor U2957 (N_2957,N_2170,N_2343);
or U2958 (N_2958,In_2961,N_622);
and U2959 (N_2959,N_2420,In_2091);
or U2960 (N_2960,N_2573,In_2793);
and U2961 (N_2961,N_940,N_1468);
xnor U2962 (N_2962,N_2257,N_2595);
nor U2963 (N_2963,In_1615,In_2820);
nor U2964 (N_2964,In_1617,N_794);
nand U2965 (N_2965,N_2716,N_1704);
nand U2966 (N_2966,In_590,N_2293);
or U2967 (N_2967,N_2555,In_3997);
or U2968 (N_2968,N_1072,N_1603);
nand U2969 (N_2969,N_317,In_4608);
nand U2970 (N_2970,In_1385,In_1742);
nand U2971 (N_2971,In_3277,N_2150);
xnor U2972 (N_2972,In_2489,In_3480);
nor U2973 (N_2973,N_1779,N_2676);
and U2974 (N_2974,In_2567,N_1858);
xor U2975 (N_2975,In_2281,In_2529);
and U2976 (N_2976,N_89,N_24);
nand U2977 (N_2977,In_2853,N_2337);
nor U2978 (N_2978,N_1802,N_1981);
and U2979 (N_2979,In_1365,N_292);
and U2980 (N_2980,N_658,In_3296);
nand U2981 (N_2981,N_932,N_2490);
or U2982 (N_2982,In_779,In_4387);
xnor U2983 (N_2983,N_2520,In_4002);
or U2984 (N_2984,In_967,N_2620);
and U2985 (N_2985,N_2659,In_3272);
and U2986 (N_2986,N_1966,N_2243);
or U2987 (N_2987,In_4573,In_1944);
and U2988 (N_2988,In_4495,In_2438);
nand U2989 (N_2989,N_55,In_4472);
nor U2990 (N_2990,N_1604,In_1790);
nor U2991 (N_2991,N_2368,N_1868);
nor U2992 (N_2992,N_1898,In_1438);
nand U2993 (N_2993,N_735,N_355);
and U2994 (N_2994,N_2695,N_233);
xor U2995 (N_2995,In_566,In_2092);
xnor U2996 (N_2996,N_2463,N_2295);
xor U2997 (N_2997,N_2414,N_2615);
xnor U2998 (N_2998,In_9,In_3416);
nor U2999 (N_2999,N_1537,N_1963);
nand U3000 (N_3000,In_2938,In_647);
nor U3001 (N_3001,N_2663,In_3155);
or U3002 (N_3002,N_238,In_3702);
xnor U3003 (N_3003,In_4817,In_2370);
and U3004 (N_3004,N_946,N_2073);
or U3005 (N_3005,N_146,N_1904);
xor U3006 (N_3006,In_284,In_1560);
and U3007 (N_3007,In_539,In_1287);
or U3008 (N_3008,In_2619,N_1957);
and U3009 (N_3009,N_2912,N_1620);
nor U3010 (N_3010,N_2770,N_1154);
nand U3011 (N_3011,In_2925,N_2540);
nor U3012 (N_3012,In_135,In_1208);
nand U3013 (N_3013,N_2829,N_2889);
and U3014 (N_3014,In_3291,N_2267);
or U3015 (N_3015,N_570,N_2479);
and U3016 (N_3016,N_2926,In_4253);
and U3017 (N_3017,N_2393,N_2775);
nor U3018 (N_3018,In_3633,N_2994);
or U3019 (N_3019,N_2292,In_4034);
and U3020 (N_3020,N_2606,N_2296);
and U3021 (N_3021,In_2956,In_2175);
nand U3022 (N_3022,N_1129,In_3891);
xnor U3023 (N_3023,N_916,N_1238);
and U3024 (N_3024,N_2883,In_2028);
nor U3025 (N_3025,N_971,In_4366);
and U3026 (N_3026,In_2719,In_3203);
nor U3027 (N_3027,N_2672,In_3222);
or U3028 (N_3028,N_2932,N_1894);
and U3029 (N_3029,N_2963,In_1188);
and U3030 (N_3030,N_1973,N_2037);
or U3031 (N_3031,In_4078,N_2326);
nand U3032 (N_3032,N_2821,N_2698);
or U3033 (N_3033,In_1485,N_2697);
or U3034 (N_3034,N_1195,N_2900);
xor U3035 (N_3035,In_2461,N_123);
nand U3036 (N_3036,N_2997,N_411);
nand U3037 (N_3037,In_3469,N_2993);
nor U3038 (N_3038,N_1751,N_2925);
nand U3039 (N_3039,N_2405,In_3197);
xnor U3040 (N_3040,N_2905,N_2929);
nor U3041 (N_3041,N_2559,N_2364);
nand U3042 (N_3042,N_2054,N_2389);
and U3043 (N_3043,N_1668,N_1749);
nand U3044 (N_3044,In_4079,In_898);
nor U3045 (N_3045,N_2461,N_2874);
nand U3046 (N_3046,In_907,N_1019);
nand U3047 (N_3047,N_1720,N_1784);
nand U3048 (N_3048,In_850,In_1788);
or U3049 (N_3049,In_4146,In_2292);
xnor U3050 (N_3050,N_2506,N_2645);
nand U3051 (N_3051,In_2632,N_2941);
nand U3052 (N_3052,N_2209,N_372);
nor U3053 (N_3053,In_1332,N_1799);
or U3054 (N_3054,N_1785,In_1568);
nand U3055 (N_3055,In_4043,In_205);
nand U3056 (N_3056,N_1050,In_1164);
xnor U3057 (N_3057,In_2039,In_1844);
nor U3058 (N_3058,N_207,N_2069);
nand U3059 (N_3059,N_1826,N_969);
and U3060 (N_3060,N_2316,In_4502);
nor U3061 (N_3061,In_1631,N_643);
and U3062 (N_3062,In_1085,In_2077);
and U3063 (N_3063,N_2394,N_2612);
xnor U3064 (N_3064,N_2893,In_3354);
nand U3065 (N_3065,N_2688,N_2436);
and U3066 (N_3066,In_3135,N_1487);
xor U3067 (N_3067,N_1216,In_2205);
nand U3068 (N_3068,N_1022,N_674);
and U3069 (N_3069,N_283,N_1069);
and U3070 (N_3070,N_1923,N_1610);
or U3071 (N_3071,N_169,In_4945);
and U3072 (N_3072,N_1299,N_1451);
or U3073 (N_3073,N_613,N_2733);
and U3074 (N_3074,N_787,In_2129);
and U3075 (N_3075,In_3731,N_903);
nor U3076 (N_3076,In_4830,In_2267);
nor U3077 (N_3077,N_2640,In_1549);
and U3078 (N_3078,N_218,N_1970);
xnor U3079 (N_3079,In_2497,N_2825);
nand U3080 (N_3080,In_2898,N_2160);
nand U3081 (N_3081,In_2678,In_3707);
nor U3082 (N_3082,N_2596,In_3823);
nor U3083 (N_3083,N_2996,N_2278);
nor U3084 (N_3084,N_2594,N_26);
and U3085 (N_3085,In_4186,In_1427);
nand U3086 (N_3086,In_1669,N_1572);
or U3087 (N_3087,N_399,In_2918);
nand U3088 (N_3088,In_823,N_2839);
nor U3089 (N_3089,N_2833,N_2704);
nand U3090 (N_3090,In_4591,N_2406);
nor U3091 (N_3091,N_1649,N_2882);
or U3092 (N_3092,N_651,In_3163);
or U3093 (N_3093,N_2864,In_3230);
or U3094 (N_3094,N_2070,In_1884);
and U3095 (N_3095,In_400,N_713);
and U3096 (N_3096,N_2700,N_2959);
and U3097 (N_3097,In_4256,N_2719);
and U3098 (N_3098,In_367,In_3753);
nand U3099 (N_3099,In_3983,In_925);
nor U3100 (N_3100,In_1270,N_2563);
xnor U3101 (N_3101,In_2848,N_1905);
nand U3102 (N_3102,In_194,In_304);
and U3103 (N_3103,N_2624,N_2793);
nor U3104 (N_3104,In_900,N_1155);
and U3105 (N_3105,N_2486,N_2918);
or U3106 (N_3106,In_2452,N_2867);
or U3107 (N_3107,N_1571,In_4995);
nand U3108 (N_3108,In_192,N_488);
nor U3109 (N_3109,N_1422,N_1651);
and U3110 (N_3110,In_4087,N_2290);
and U3111 (N_3111,In_4700,In_1813);
xor U3112 (N_3112,N_853,N_1204);
and U3113 (N_3113,N_1057,N_1953);
nor U3114 (N_3114,N_1101,In_2987);
and U3115 (N_3115,N_2910,N_2574);
nor U3116 (N_3116,In_2026,N_1830);
xor U3117 (N_3117,N_2464,N_2609);
and U3118 (N_3118,N_2785,N_2886);
or U3119 (N_3119,In_1799,In_2813);
nand U3120 (N_3120,In_4732,N_2586);
and U3121 (N_3121,In_4926,N_2380);
nand U3122 (N_3122,N_1114,In_595);
and U3123 (N_3123,In_1294,In_3650);
nand U3124 (N_3124,In_869,N_2903);
and U3125 (N_3125,N_516,N_2159);
and U3126 (N_3126,N_1305,N_2106);
nand U3127 (N_3127,In_1439,N_2313);
and U3128 (N_3128,In_4552,N_2971);
nand U3129 (N_3129,N_1158,N_2872);
or U3130 (N_3130,N_1900,N_1037);
xor U3131 (N_3131,N_1279,N_2836);
xor U3132 (N_3132,In_2702,N_2214);
xnor U3133 (N_3133,In_1266,In_1476);
nand U3134 (N_3134,N_2827,In_3336);
and U3135 (N_3135,N_2530,N_2950);
and U3136 (N_3136,In_203,N_605);
xor U3137 (N_3137,N_805,N_2658);
nor U3138 (N_3138,In_4701,N_1825);
nor U3139 (N_3139,N_2551,N_2863);
xor U3140 (N_3140,In_3461,N_2538);
or U3141 (N_3141,In_4998,In_2924);
nand U3142 (N_3142,In_2923,N_1173);
or U3143 (N_3143,N_1082,N_1884);
and U3144 (N_3144,N_2107,In_52);
or U3145 (N_3145,In_4733,In_1623);
xnor U3146 (N_3146,N_2500,In_2135);
xnor U3147 (N_3147,In_552,N_2153);
nor U3148 (N_3148,N_119,N_1639);
nor U3149 (N_3149,N_2788,N_2514);
or U3150 (N_3150,In_4690,N_455);
and U3151 (N_3151,In_3659,N_1804);
and U3152 (N_3152,N_1579,N_2957);
or U3153 (N_3153,N_2196,N_2944);
xnor U3154 (N_3154,N_1990,In_181);
xor U3155 (N_3155,In_4836,N_2812);
or U3156 (N_3156,In_800,N_270);
and U3157 (N_3157,In_2227,N_2381);
or U3158 (N_3158,N_2678,N_2939);
xnor U3159 (N_3159,N_1516,In_3294);
xor U3160 (N_3160,N_1348,In_4326);
xor U3161 (N_3161,N_1454,In_4853);
nand U3162 (N_3162,In_1656,N_1047);
nor U3163 (N_3163,N_2965,N_2077);
xor U3164 (N_3164,N_2047,N_887);
nand U3165 (N_3165,N_2504,N_2954);
xor U3166 (N_3166,N_1284,N_2807);
xnor U3167 (N_3167,N_2549,In_2902);
nor U3168 (N_3168,In_297,N_2792);
xor U3169 (N_3169,N_1094,In_3684);
nand U3170 (N_3170,In_860,N_1886);
xnor U3171 (N_3171,N_1752,N_2643);
nand U3172 (N_3172,In_2772,N_2811);
nand U3173 (N_3173,N_2986,N_1223);
or U3174 (N_3174,N_136,N_2284);
nand U3175 (N_3175,In_4959,N_1460);
nor U3176 (N_3176,N_2516,N_2534);
xnor U3177 (N_3177,In_3738,In_14);
xor U3178 (N_3178,N_2344,In_4162);
nand U3179 (N_3179,N_2133,N_2357);
and U3180 (N_3180,N_2774,In_3397);
or U3181 (N_3181,In_2388,N_2442);
or U3182 (N_3182,N_2093,N_2656);
and U3183 (N_3183,In_4632,N_2421);
or U3184 (N_3184,In_1554,N_1132);
nor U3185 (N_3185,N_2046,In_2379);
xnor U3186 (N_3186,N_2146,N_2137);
and U3187 (N_3187,N_1739,N_2437);
xnor U3188 (N_3188,In_3182,N_1577);
or U3189 (N_3189,N_1817,In_4313);
nand U3190 (N_3190,In_4250,N_2834);
or U3191 (N_3191,N_1148,N_2679);
nand U3192 (N_3192,In_4158,N_1443);
or U3193 (N_3193,In_971,N_491);
nor U3194 (N_3194,N_2861,N_469);
or U3195 (N_3195,In_2070,N_2691);
nor U3196 (N_3196,N_2447,N_1118);
and U3197 (N_3197,In_4436,N_495);
or U3198 (N_3198,N_85,N_2945);
nand U3199 (N_3199,N_2220,N_1568);
and U3200 (N_3200,In_743,N_1398);
nor U3201 (N_3201,In_4979,N_2860);
xor U3202 (N_3202,N_2820,N_2936);
xnor U3203 (N_3203,N_1727,N_999);
nand U3204 (N_3204,N_2342,In_2595);
nand U3205 (N_3205,N_2619,In_4991);
xor U3206 (N_3206,In_538,N_2048);
nand U3207 (N_3207,N_2667,N_2340);
or U3208 (N_3208,In_3218,N_1694);
nor U3209 (N_3209,N_2911,N_2477);
nor U3210 (N_3210,N_2919,N_2554);
or U3211 (N_3211,N_2281,N_2921);
nand U3212 (N_3212,N_2,N_1762);
xor U3213 (N_3213,N_1083,In_1277);
nand U3214 (N_3214,N_2557,N_2879);
xor U3215 (N_3215,N_2492,N_2852);
nand U3216 (N_3216,N_2894,In_286);
nand U3217 (N_3217,N_2365,In_2381);
nand U3218 (N_3218,In_4271,In_3123);
nand U3219 (N_3219,N_1697,N_2521);
and U3220 (N_3220,N_1536,N_521);
nor U3221 (N_3221,In_4525,N_816);
or U3222 (N_3222,N_1167,In_323);
xor U3223 (N_3223,N_2168,N_2503);
xnor U3224 (N_3224,N_2752,In_863);
nor U3225 (N_3225,In_1044,In_3697);
and U3226 (N_3226,N_2256,N_949);
or U3227 (N_3227,In_4862,In_3338);
nor U3228 (N_3228,N_1402,In_3728);
nand U3229 (N_3229,N_2617,N_2507);
or U3230 (N_3230,N_775,In_3838);
xor U3231 (N_3231,In_1607,N_2933);
or U3232 (N_3232,N_2703,In_1192);
or U3233 (N_3233,N_1918,In_3604);
and U3234 (N_3234,N_885,In_3468);
and U3235 (N_3235,N_2851,N_2767);
and U3236 (N_3236,In_4418,N_2657);
or U3237 (N_3237,N_2962,In_4786);
or U3238 (N_3238,N_1295,In_3696);
xnor U3239 (N_3239,N_1425,N_2628);
or U3240 (N_3240,N_2784,In_4010);
xor U3241 (N_3241,N_2020,In_1236);
or U3242 (N_3242,N_1511,N_2830);
nand U3243 (N_3243,N_2805,In_2797);
and U3244 (N_3244,N_2301,In_4993);
nand U3245 (N_3245,In_4543,N_223);
or U3246 (N_3246,N_162,N_2067);
nor U3247 (N_3247,N_2729,N_2556);
and U3248 (N_3248,N_795,N_361);
xor U3249 (N_3249,N_2778,N_2402);
nand U3250 (N_3250,N_2465,N_1431);
xnor U3251 (N_3251,N_2471,In_3567);
nor U3252 (N_3252,N_44,N_2017);
or U3253 (N_3253,N_2735,N_1965);
nor U3254 (N_3254,N_1346,In_4243);
nor U3255 (N_3255,N_3183,N_2949);
or U3256 (N_3256,In_581,N_1108);
nand U3257 (N_3257,N_2134,N_2208);
nand U3258 (N_3258,N_3049,In_1010);
or U3259 (N_3259,In_2462,In_4269);
nand U3260 (N_3260,N_2132,N_2607);
and U3261 (N_3261,N_3052,In_2617);
nand U3262 (N_3262,In_3501,N_2610);
nand U3263 (N_3263,N_2424,N_3242);
xor U3264 (N_3264,N_3092,N_2815);
xor U3265 (N_3265,N_2234,N_2315);
and U3266 (N_3266,N_1439,In_3055);
nand U3267 (N_3267,N_2042,N_1573);
nor U3268 (N_3268,N_2536,In_956);
xnor U3269 (N_3269,N_2992,N_2585);
and U3270 (N_3270,N_1638,In_418);
and U3271 (N_3271,N_1349,N_1962);
or U3272 (N_3272,N_2266,In_4767);
and U3273 (N_3273,In_4208,N_2489);
xor U3274 (N_3274,N_3083,N_3028);
or U3275 (N_3275,In_2224,N_2999);
or U3276 (N_3276,In_2579,N_3202);
nand U3277 (N_3277,N_1987,N_3058);
nand U3278 (N_3278,In_563,In_1661);
nor U3279 (N_3279,N_751,N_300);
xnor U3280 (N_3280,In_1954,N_2631);
or U3281 (N_3281,N_2440,N_3079);
nor U3282 (N_3282,N_327,N_1103);
and U3283 (N_3283,In_4984,N_3055);
nand U3284 (N_3284,N_1741,N_478);
or U3285 (N_3285,In_2109,N_3122);
and U3286 (N_3286,N_2983,In_191);
xnor U3287 (N_3287,In_2711,N_1053);
or U3288 (N_3288,N_3249,In_905);
or U3289 (N_3289,N_2780,N_2720);
or U3290 (N_3290,In_4638,In_4940);
and U3291 (N_3291,N_2263,N_1569);
xnor U3292 (N_3292,N_3001,In_4806);
or U3293 (N_3293,N_20,N_2547);
nor U3294 (N_3294,In_3602,In_3593);
nor U3295 (N_3295,N_3102,In_1611);
or U3296 (N_3296,N_2513,In_2228);
or U3297 (N_3297,N_3170,N_1337);
and U3298 (N_3298,In_2508,N_2673);
nor U3299 (N_3299,N_2970,N_2094);
xnor U3300 (N_3300,N_1345,N_3222);
or U3301 (N_3301,In_840,N_351);
nor U3302 (N_3302,In_473,N_1914);
and U3303 (N_3303,N_2826,N_458);
or U3304 (N_3304,N_2871,In_664);
xnor U3305 (N_3305,N_3248,N_3045);
and U3306 (N_3306,N_5,N_3132);
or U3307 (N_3307,In_4988,N_2236);
xnor U3308 (N_3308,N_2589,N_2746);
nor U3309 (N_3309,N_2216,N_2396);
or U3310 (N_3310,In_1379,N_1706);
xnor U3311 (N_3311,N_1444,N_2951);
or U3312 (N_3312,N_2571,N_54);
nand U3313 (N_3313,N_360,In_4981);
nor U3314 (N_3314,In_3833,N_2701);
xnor U3315 (N_3315,N_2990,In_262);
and U3316 (N_3316,N_3149,N_386);
or U3317 (N_3317,N_2953,In_95);
and U3318 (N_3318,N_1146,In_1230);
nor U3319 (N_3319,N_1313,N_3158);
nand U3320 (N_3320,N_2722,N_3209);
or U3321 (N_3321,N_306,N_3030);
xor U3322 (N_3322,In_3606,N_1523);
and U3323 (N_3323,In_2161,N_3023);
or U3324 (N_3324,N_208,In_893);
xnor U3325 (N_3325,N_2769,In_1414);
xor U3326 (N_3326,N_1040,In_88);
xnor U3327 (N_3327,N_2443,N_2798);
nor U3328 (N_3328,N_1551,N_3175);
and U3329 (N_3329,N_2881,N_3133);
and U3330 (N_3330,N_1846,N_798);
or U3331 (N_3331,N_1928,N_2505);
nor U3332 (N_3332,N_2240,N_1200);
and U3333 (N_3333,N_2976,N_3226);
xnor U3334 (N_3334,N_1798,In_4535);
or U3335 (N_3335,N_2862,N_2763);
and U3336 (N_3336,In_3757,In_4196);
nand U3337 (N_3337,N_2509,N_2611);
xor U3338 (N_3338,N_3186,N_2597);
and U3339 (N_3339,N_1969,N_2588);
nand U3340 (N_3340,N_1282,In_4203);
and U3341 (N_3341,N_855,In_3007);
or U3342 (N_3342,In_3506,N_954);
xnor U3343 (N_3343,N_3038,N_2287);
or U3344 (N_3344,N_1542,N_3181);
or U3345 (N_3345,N_1921,In_4975);
nor U3346 (N_3346,N_2835,N_2299);
xor U3347 (N_3347,N_3012,N_737);
nor U3348 (N_3348,N_2828,In_2934);
and U3349 (N_3349,N_982,N_2891);
nor U3350 (N_3350,N_2564,N_1528);
xnor U3351 (N_3351,In_4983,In_3027);
nor U3352 (N_3352,N_1853,N_1554);
xor U3353 (N_3353,N_3179,N_2425);
and U3354 (N_3354,In_1610,N_2754);
or U3355 (N_3355,In_4935,N_3223);
xnor U3356 (N_3356,N_456,N_2664);
xor U3357 (N_3357,N_3208,N_2975);
nor U3358 (N_3358,N_2751,In_513);
xnor U3359 (N_3359,N_158,N_3192);
nor U3360 (N_3360,N_2600,N_1372);
xor U3361 (N_3361,N_2682,N_3232);
and U3362 (N_3362,In_560,N_2987);
and U3363 (N_3363,In_3589,N_2304);
nand U3364 (N_3364,N_1769,In_4473);
or U3365 (N_3365,N_2814,N_2230);
nand U3366 (N_3366,N_2934,In_1204);
or U3367 (N_3367,N_2809,In_2649);
xor U3368 (N_3368,In_3483,N_2748);
or U3369 (N_3369,N_1687,In_227);
nor U3370 (N_3370,N_2294,In_1582);
xnor U3371 (N_3371,N_2255,N_636);
xnor U3372 (N_3372,In_4702,N_1462);
nor U3373 (N_3373,N_2542,N_3190);
and U3374 (N_3374,In_1886,N_3067);
xor U3375 (N_3375,In_2087,N_717);
xor U3376 (N_3376,N_2522,In_4596);
xor U3377 (N_3377,In_158,N_2708);
xnor U3378 (N_3378,In_1308,In_3199);
nor U3379 (N_3379,N_3167,N_3095);
or U3380 (N_3380,N_2090,N_2989);
nor U3381 (N_3381,In_4590,N_1949);
or U3382 (N_3382,In_3694,N_3206);
or U3383 (N_3383,N_3180,N_2451);
xnor U3384 (N_3384,N_1954,N_348);
or U3385 (N_3385,N_1679,N_3054);
and U3386 (N_3386,In_193,N_245);
nand U3387 (N_3387,N_1550,N_3184);
or U3388 (N_3388,In_4258,N_2850);
nand U3389 (N_3389,N_3059,N_2940);
and U3390 (N_3390,N_1924,In_3579);
or U3391 (N_3391,N_2712,N_36);
nor U3392 (N_3392,In_80,N_2483);
xnor U3393 (N_3393,N_333,In_3229);
xor U3394 (N_3394,N_2469,N_1227);
xnor U3395 (N_3395,N_1989,N_1291);
xnor U3396 (N_3396,N_2984,In_4360);
nor U3397 (N_3397,In_541,N_3005);
nor U3398 (N_3398,N_1319,N_1469);
nor U3399 (N_3399,In_4122,In_1851);
or U3400 (N_3400,N_286,N_3101);
nor U3401 (N_3401,N_3009,N_1459);
or U3402 (N_3402,In_3965,N_2991);
and U3403 (N_3403,In_3122,N_2499);
nand U3404 (N_3404,N_2790,N_3146);
and U3405 (N_3405,N_2920,N_2028);
xor U3406 (N_3406,N_484,N_2403);
nor U3407 (N_3407,N_3032,N_978);
and U3408 (N_3408,N_1567,N_3156);
nand U3409 (N_3409,N_3178,In_475);
or U3410 (N_3410,N_3159,In_4727);
xor U3411 (N_3411,In_4667,N_2838);
xor U3412 (N_3412,N_2670,In_3705);
nor U3413 (N_3413,N_3064,N_1624);
or U3414 (N_3414,N_3057,In_2674);
or U3415 (N_3415,N_2745,N_803);
nor U3416 (N_3416,In_4263,N_1992);
nor U3417 (N_3417,N_732,N_2426);
xnor U3418 (N_3418,N_1791,N_2397);
or U3419 (N_3419,N_1183,N_1360);
xnor U3420 (N_3420,In_4300,N_2283);
xnor U3421 (N_3421,N_2079,N_1703);
nor U3422 (N_3422,N_2938,N_508);
nand U3423 (N_3423,In_4540,In_2007);
nand U3424 (N_3424,N_2036,N_1097);
xor U3425 (N_3425,N_400,In_1386);
xor U3426 (N_3426,N_1754,N_2873);
xnor U3427 (N_3427,In_215,In_2894);
or U3428 (N_3428,In_4925,N_2756);
and U3429 (N_3429,N_1844,N_3075);
nor U3430 (N_3430,N_1055,N_3000);
or U3431 (N_3431,N_2808,In_1351);
xnor U3432 (N_3432,N_1196,N_2057);
or U3433 (N_3433,N_3161,N_3042);
and U3434 (N_3434,N_1479,In_4970);
and U3435 (N_3435,N_3123,In_1928);
or U3436 (N_3436,In_2340,N_1711);
or U3437 (N_3437,N_3110,N_1892);
and U3438 (N_3438,In_1363,N_2973);
and U3439 (N_3439,N_2736,N_1594);
nand U3440 (N_3440,N_2801,In_2085);
and U3441 (N_3441,In_2106,N_3017);
or U3442 (N_3442,In_4976,In_1877);
and U3443 (N_3443,In_834,In_738);
nand U3444 (N_3444,N_2007,N_3125);
nor U3445 (N_3445,In_4209,N_2599);
nor U3446 (N_3446,In_3195,N_1944);
nand U3447 (N_3447,N_3217,In_4448);
or U3448 (N_3448,In_4458,N_256);
xnor U3449 (N_3449,In_2713,In_2471);
and U3450 (N_3450,N_2779,N_2802);
and U3451 (N_3451,N_3109,In_3434);
nand U3452 (N_3452,N_3241,N_2819);
and U3453 (N_3453,N_2630,In_3718);
or U3454 (N_3454,In_251,N_840);
and U3455 (N_3455,N_834,N_3063);
nand U3456 (N_3456,N_3195,N_2115);
nand U3457 (N_3457,N_3014,N_575);
nand U3458 (N_3458,N_3056,N_1085);
nand U3459 (N_3459,In_1908,N_3129);
xor U3460 (N_3460,In_2468,N_968);
nor U3461 (N_3461,In_1265,In_3391);
xnor U3462 (N_3462,N_2049,N_1342);
nand U3463 (N_3463,In_3112,N_2837);
and U3464 (N_3464,N_2904,In_1007);
or U3465 (N_3465,N_1950,In_1808);
nand U3466 (N_3466,N_2371,In_1950);
nor U3467 (N_3467,N_312,N_1640);
and U3468 (N_3468,N_2334,In_1695);
xnor U3469 (N_3469,N_2759,N_2909);
and U3470 (N_3470,N_2636,N_3207);
and U3471 (N_3471,N_101,N_3084);
nand U3472 (N_3472,N_1236,In_512);
nand U3473 (N_3473,In_715,N_2449);
nand U3474 (N_3474,N_1808,N_84);
or U3475 (N_3475,N_3150,N_3210);
xnor U3476 (N_3476,N_3213,In_2136);
nand U3477 (N_3477,N_437,N_3233);
nand U3478 (N_3478,N_3165,N_2842);
nand U3479 (N_3479,In_771,N_1527);
xnor U3480 (N_3480,N_2026,N_3137);
nor U3481 (N_3481,N_2272,N_3085);
nor U3482 (N_3482,N_1578,N_750);
nor U3483 (N_3483,N_273,N_915);
nor U3484 (N_3484,N_2312,In_3166);
nand U3485 (N_3485,In_597,N_3246);
nand U3486 (N_3486,N_3188,N_3006);
nand U3487 (N_3487,N_2966,N_2454);
xnor U3488 (N_3488,N_2859,In_102);
xnor U3489 (N_3489,N_2783,In_2102);
and U3490 (N_3490,N_2219,N_1701);
nor U3491 (N_3491,N_3088,N_2567);
xor U3492 (N_3492,N_901,N_500);
xnor U3493 (N_3493,In_4398,In_3638);
or U3494 (N_3494,N_235,In_3931);
nand U3495 (N_3495,In_1530,N_2613);
nand U3496 (N_3496,N_2709,N_2637);
xnor U3497 (N_3497,N_2853,N_2128);
xor U3498 (N_3498,N_2376,In_4558);
nor U3499 (N_3499,N_2416,In_2402);
and U3500 (N_3500,N_3087,N_544);
or U3501 (N_3501,In_4290,N_2318);
nand U3502 (N_3502,N_2061,In_3719);
and U3503 (N_3503,N_3182,In_630);
and U3504 (N_3504,In_2152,N_2699);
nand U3505 (N_3505,N_2869,N_2865);
and U3506 (N_3506,In_3737,N_2457);
and U3507 (N_3507,In_1089,N_3419);
nand U3508 (N_3508,N_3314,N_3153);
nand U3509 (N_3509,N_164,N_3376);
xor U3510 (N_3510,In_2905,In_2055);
nor U3511 (N_3511,In_3978,N_1612);
xnor U3512 (N_3512,N_2181,In_1812);
or U3513 (N_3513,N_2367,N_2076);
nand U3514 (N_3514,N_2843,N_3351);
xnor U3515 (N_3515,N_2075,In_4609);
nand U3516 (N_3516,N_3078,In_2735);
xnor U3517 (N_3517,N_2192,N_2913);
and U3518 (N_3518,N_389,In_2188);
xnor U3519 (N_3519,N_1810,N_3359);
and U3520 (N_3520,N_1777,N_1974);
xnor U3521 (N_3521,N_1531,N_2744);
xor U3522 (N_3522,N_3345,N_3388);
and U3523 (N_3523,In_1371,N_2053);
xor U3524 (N_3524,In_3935,N_2806);
and U3525 (N_3525,In_166,N_1127);
nand U3526 (N_3526,N_3478,N_2895);
xnor U3527 (N_3527,N_3363,N_3236);
xnor U3528 (N_3528,N_1982,N_3198);
nand U3529 (N_3529,In_4011,N_588);
nor U3530 (N_3530,N_3406,N_3367);
nor U3531 (N_3531,In_1435,In_3905);
xor U3532 (N_3532,N_3229,N_2092);
or U3533 (N_3533,N_1054,N_3234);
xnor U3534 (N_3534,In_1222,In_2833);
xor U3535 (N_3535,N_912,N_3237);
nor U3536 (N_3536,In_3903,N_3162);
nor U3537 (N_3537,In_1722,N_2917);
nor U3538 (N_3538,N_1818,N_2482);
or U3539 (N_3539,N_3261,N_3120);
or U3540 (N_3540,N_762,N_2569);
and U3541 (N_3541,N_2525,In_2133);
xnor U3542 (N_3542,N_612,N_3257);
nor U3543 (N_3543,In_2860,In_398);
nor U3544 (N_3544,In_4955,N_2740);
and U3545 (N_3545,In_845,N_2654);
nand U3546 (N_3546,In_4741,In_996);
or U3547 (N_3547,N_3456,N_3046);
xnor U3548 (N_3548,N_3301,In_725);
nand U3549 (N_3549,N_629,N_2787);
xor U3550 (N_3550,In_2225,N_1339);
and U3551 (N_3551,In_4656,N_1781);
or U3552 (N_3552,N_2496,In_4093);
nand U3553 (N_3553,In_778,N_1909);
xor U3554 (N_3554,In_2001,N_2680);
and U3555 (N_3555,N_3362,N_3131);
nor U3556 (N_3556,N_3285,N_3041);
xor U3557 (N_3557,In_557,In_416);
xor U3558 (N_3558,N_2760,N_1626);
xnor U3559 (N_3559,N_3453,In_427);
nor U3560 (N_3560,In_613,In_3513);
xnor U3561 (N_3561,N_2998,N_3004);
nor U3562 (N_3562,N_1356,N_3293);
or U3563 (N_3563,In_431,In_3447);
and U3564 (N_3564,In_526,N_2714);
nor U3565 (N_3565,N_141,N_2016);
xor U3566 (N_3566,In_1720,In_2016);
nand U3567 (N_3567,N_3027,N_2854);
xor U3568 (N_3568,N_1258,N_2050);
and U3569 (N_3569,N_2822,N_2139);
or U3570 (N_3570,N_1188,N_2978);
nor U3571 (N_3571,N_3225,N_1429);
nor U3572 (N_3572,N_1561,N_2006);
nor U3573 (N_3573,N_3139,N_2528);
nor U3574 (N_3574,N_1870,N_3338);
nand U3575 (N_3575,N_74,N_1404);
xor U3576 (N_3576,N_1157,N_1541);
nor U3577 (N_3577,N_3157,N_1663);
or U3578 (N_3578,N_3379,N_2718);
or U3579 (N_3579,N_2947,N_1255);
xor U3580 (N_3580,N_2901,N_2766);
xnor U3581 (N_3581,N_592,N_862);
or U3582 (N_3582,N_3108,In_1800);
nor U3583 (N_3583,N_3218,N_522);
nor U3584 (N_3584,In_1445,N_379);
xnor U3585 (N_3585,N_3047,N_3071);
nand U3586 (N_3586,N_3228,In_4457);
or U3587 (N_3587,N_3276,N_2541);
nand U3588 (N_3588,N_1678,In_3955);
and U3589 (N_3589,N_801,In_3167);
and U3590 (N_3590,N_2685,N_3317);
or U3591 (N_3591,N_1665,N_3355);
nand U3592 (N_3592,N_1947,N_1793);
or U3593 (N_3593,N_3215,N_1144);
nand U3594 (N_3594,N_3034,N_3196);
nand U3595 (N_3595,N_1024,In_1516);
xor U3596 (N_3596,In_4728,N_1713);
or U3597 (N_3597,In_2688,N_1099);
nor U3598 (N_3598,N_1478,In_1719);
and U3599 (N_3599,N_1611,In_3148);
nand U3600 (N_3600,N_2795,In_3817);
nor U3601 (N_3601,N_3097,N_3077);
nand U3602 (N_3602,N_2732,N_3168);
nor U3603 (N_3603,N_1869,N_2896);
nor U3604 (N_3604,In_4349,N_1839);
xnor U3605 (N_3605,N_2179,In_2555);
or U3606 (N_3606,In_3248,In_1670);
and U3607 (N_3607,N_1106,N_1682);
nand U3608 (N_3608,In_1473,In_1528);
and U3609 (N_3609,N_3340,N_3262);
xor U3610 (N_3610,In_2560,N_3243);
or U3611 (N_3611,In_2282,In_1233);
xnor U3612 (N_3612,N_3466,N_1821);
or U3613 (N_3613,In_920,In_3297);
nor U3614 (N_3614,N_3320,In_3548);
nand U3615 (N_3615,N_1314,In_1870);
and U3616 (N_3616,N_819,N_1843);
nand U3617 (N_3617,N_3312,N_1205);
xor U3618 (N_3618,In_544,In_940);
and U3619 (N_3619,In_1471,N_1126);
and U3620 (N_3620,N_3366,In_4404);
nor U3621 (N_3621,N_3348,In_1758);
xor U3622 (N_3622,N_3141,N_1916);
and U3623 (N_3623,In_1088,N_358);
or U3624 (N_3624,N_3060,In_225);
nor U3625 (N_3625,N_1073,In_4974);
and U3626 (N_3626,In_1128,N_3499);
and U3627 (N_3627,In_4920,In_98);
nand U3628 (N_3628,N_2561,N_2237);
xnor U3629 (N_3629,N_2715,N_152);
and U3630 (N_3630,N_3472,N_2162);
xnor U3631 (N_3631,N_2480,N_1071);
xnor U3632 (N_3632,In_1764,N_2943);
or U3633 (N_3633,N_2131,N_3310);
and U3634 (N_3634,N_2668,In_4652);
or U3635 (N_3635,N_2488,N_2088);
or U3636 (N_3636,N_3124,N_2206);
and U3637 (N_3637,N_3344,In_4045);
nand U3638 (N_3638,In_4744,N_3307);
nor U3639 (N_3639,In_4800,In_2435);
xnor U3640 (N_3640,N_681,In_748);
and U3641 (N_3641,N_1915,N_1891);
and U3642 (N_3642,N_1544,In_2532);
xor U3643 (N_3643,N_3417,In_312);
and U3644 (N_3644,N_3490,N_3392);
xnor U3645 (N_3645,In_2488,N_2644);
or U3646 (N_3646,N_3013,N_2960);
or U3647 (N_3647,N_1502,In_1354);
nor U3648 (N_3648,In_3053,N_3201);
and U3649 (N_3649,In_3619,N_3138);
nor U3650 (N_3650,N_2618,N_3400);
nor U3651 (N_3651,N_1417,N_3203);
nor U3652 (N_3652,In_16,N_2166);
nor U3653 (N_3653,N_395,N_3076);
xor U3654 (N_3654,N_132,N_2578);
nor U3655 (N_3655,N_1995,N_2515);
or U3656 (N_3656,N_1340,N_3306);
nor U3657 (N_3657,N_1492,N_1222);
xor U3658 (N_3658,N_3263,In_2933);
xnor U3659 (N_3659,N_3384,N_3291);
xor U3660 (N_3660,N_1557,In_3159);
xor U3661 (N_3661,N_2190,N_3302);
and U3662 (N_3662,N_2410,N_2980);
nand U3663 (N_3663,In_1662,N_2616);
nor U3664 (N_3664,N_3394,N_3418);
xnor U3665 (N_3665,N_2967,N_3134);
or U3666 (N_3666,N_3245,N_2391);
xnor U3667 (N_3667,N_1885,N_3140);
nand U3668 (N_3668,N_3255,In_1940);
nor U3669 (N_3669,N_3062,N_401);
or U3670 (N_3670,N_3360,In_2999);
or U3671 (N_3671,In_662,N_3189);
nand U3672 (N_3672,N_2517,N_3114);
nand U3673 (N_3673,In_3119,N_1625);
nand U3674 (N_3674,N_99,N_3116);
nand U3675 (N_3675,N_3477,N_3311);
xor U3676 (N_3676,N_1856,N_723);
nand U3677 (N_3677,In_2696,In_1475);
and U3678 (N_3678,N_2622,N_3482);
nor U3679 (N_3679,In_1246,N_3100);
and U3680 (N_3680,N_2803,N_3160);
or U3681 (N_3681,N_2593,N_2581);
xnor U3682 (N_3682,N_2728,In_1878);
xnor U3683 (N_3683,N_1942,In_254);
xor U3684 (N_3684,In_3439,N_2858);
xor U3685 (N_3685,N_774,N_3354);
or U3686 (N_3686,In_4227,In_1725);
or U3687 (N_3687,N_3391,N_3377);
nor U3688 (N_3688,In_2429,N_3264);
xnor U3689 (N_3689,In_1398,N_2310);
nor U3690 (N_3690,In_4233,In_2748);
nor U3691 (N_3691,In_1292,In_4382);
nor U3692 (N_3692,N_1862,N_3274);
or U3693 (N_3693,N_3048,In_2245);
or U3694 (N_3694,N_2568,N_2232);
nand U3695 (N_3695,N_3434,N_3147);
nand U3696 (N_3696,In_4096,In_706);
nor U3697 (N_3697,N_1455,In_4887);
nor U3698 (N_3698,N_2948,N_1526);
and U3699 (N_3699,N_2627,In_2041);
nor U3700 (N_3700,N_2888,In_2641);
and U3701 (N_3701,N_2690,N_2878);
and U3702 (N_3702,N_3026,In_3740);
xor U3703 (N_3703,In_148,N_1213);
and U3704 (N_3704,In_804,N_3211);
nor U3705 (N_3705,In_124,N_595);
or U3706 (N_3706,N_2632,N_3287);
xor U3707 (N_3707,N_3308,In_1520);
or U3708 (N_3708,In_3260,N_563);
and U3709 (N_3709,In_4825,N_3475);
nor U3710 (N_3710,N_3409,N_1842);
nand U3711 (N_3711,N_3381,N_177);
nand U3712 (N_3712,In_4283,N_3416);
or U3713 (N_3713,N_2535,N_2347);
nor U3714 (N_3714,N_3096,N_864);
and U3715 (N_3715,N_2188,N_3002);
or U3716 (N_3716,N_2727,In_3078);
nor U3717 (N_3717,In_4939,N_3173);
and U3718 (N_3718,In_2884,N_1666);
and U3719 (N_3719,N_1424,N_2804);
xnor U3720 (N_3720,N_1298,N_3284);
nor U3721 (N_3721,N_3117,N_3396);
or U3722 (N_3722,In_718,In_1282);
nand U3723 (N_3723,N_2849,In_4363);
and U3724 (N_3724,In_1539,N_2439);
nand U3725 (N_3725,N_2033,In_185);
nor U3726 (N_3726,N_1806,In_1672);
xor U3727 (N_3727,N_3003,N_2432);
or U3728 (N_3728,N_3430,In_3341);
nand U3729 (N_3729,N_2724,N_1851);
nor U3730 (N_3730,In_4876,In_4180);
and U3731 (N_3731,N_2935,N_2915);
nor U3732 (N_3732,N_2823,N_831);
xnor U3733 (N_3733,In_4798,N_3050);
xnor U3734 (N_3734,N_3336,N_3011);
xnor U3735 (N_3735,N_2687,N_2648);
or U3736 (N_3736,N_2211,N_2274);
nand U3737 (N_3737,N_3281,N_2955);
and U3738 (N_3738,N_2742,N_2601);
or U3739 (N_3739,N_3169,N_73);
and U3740 (N_3740,In_4861,In_2510);
nor U3741 (N_3741,N_2633,N_3343);
nand U3742 (N_3742,N_2661,N_871);
nor U3743 (N_3743,N_2021,N_585);
xor U3744 (N_3744,N_3428,N_3313);
or U3745 (N_3745,In_3639,N_1330);
or U3746 (N_3746,N_2261,N_3385);
nor U3747 (N_3747,N_2824,In_372);
nand U3748 (N_3748,In_1496,N_1609);
and U3749 (N_3749,N_2693,N_1685);
nor U3750 (N_3750,N_3703,In_382);
nand U3751 (N_3751,N_168,In_1753);
xnor U3752 (N_3752,In_4216,N_2579);
nand U3753 (N_3753,N_3719,N_3205);
nor U3754 (N_3754,N_3152,N_2321);
xor U3755 (N_3755,N_1765,N_2651);
and U3756 (N_3756,N_2927,N_3035);
or U3757 (N_3757,N_1310,N_3269);
or U3758 (N_3758,N_2583,N_2665);
nand U3759 (N_3759,N_2898,N_3099);
nand U3760 (N_3760,N_2438,N_3177);
nor U3761 (N_3761,N_2899,In_604);
nand U3762 (N_3762,N_2071,N_2314);
nand U3763 (N_3763,N_3070,In_701);
nand U3764 (N_3764,N_2604,In_3247);
nand U3765 (N_3765,N_2497,N_3305);
and U3766 (N_3766,N_2813,N_3500);
nor U3767 (N_3767,In_3847,In_2871);
or U3768 (N_3768,N_397,N_2412);
nor U3769 (N_3769,N_2031,N_2580);
and U3770 (N_3770,In_113,N_3128);
xnor U3771 (N_3771,N_2529,In_3428);
and U3772 (N_3772,N_3671,In_4267);
and U3773 (N_3773,N_2379,N_1075);
nand U3774 (N_3774,N_3352,N_3491);
and U3775 (N_3775,N_3699,N_3552);
or U3776 (N_3776,N_3669,N_1378);
xnor U3777 (N_3777,N_845,N_3069);
xnor U3778 (N_3778,N_2880,N_1621);
and U3779 (N_3779,In_1058,N_3044);
and U3780 (N_3780,N_2062,N_3675);
nand U3781 (N_3781,N_1376,In_2887);
and U3782 (N_3782,N_3627,N_2666);
nand U3783 (N_3783,N_3670,N_1792);
xor U3784 (N_3784,N_3642,N_239);
xnor U3785 (N_3785,N_977,N_3705);
or U3786 (N_3786,N_2055,In_2211);
nor U3787 (N_3787,N_3709,In_3764);
xor U3788 (N_3788,N_919,In_1348);
and U3789 (N_3789,N_2647,In_3814);
and U3790 (N_3790,N_2533,N_3688);
nand U3791 (N_3791,N_2419,N_1296);
xor U3792 (N_3792,N_3235,N_2523);
xnor U3793 (N_3793,N_3332,N_3503);
nor U3794 (N_3794,In_66,N_3717);
xor U3795 (N_3795,N_3460,N_2946);
nand U3796 (N_3796,In_471,In_2826);
or U3797 (N_3797,N_2870,N_3441);
xor U3798 (N_3798,N_1787,N_3008);
xor U3799 (N_3799,N_3335,N_2474);
and U3800 (N_3800,N_1160,N_3533);
or U3801 (N_3801,In_1087,N_3437);
nor U3802 (N_3802,N_958,N_1599);
xor U3803 (N_3803,N_3504,In_4584);
nor U3804 (N_3804,In_1556,N_2167);
nand U3805 (N_3805,N_3036,N_964);
xor U3806 (N_3806,N_1177,In_4832);
and U3807 (N_3807,In_4068,N_3510);
nor U3808 (N_3808,N_1702,N_2931);
nor U3809 (N_3809,N_2603,N_2866);
and U3810 (N_3810,In_608,N_1875);
nand U3811 (N_3811,In_864,N_3403);
and U3812 (N_3812,N_3272,N_3534);
xor U3813 (N_3813,In_2765,N_3524);
nor U3814 (N_3814,N_3292,N_2739);
xor U3815 (N_3815,N_1763,N_1049);
nand U3816 (N_3816,N_3435,N_1512);
and U3817 (N_3817,N_1732,N_2271);
xnor U3818 (N_3818,N_2713,N_3333);
nand U3819 (N_3819,N_3424,N_3072);
and U3820 (N_3820,N_3692,N_2566);
nand U3821 (N_3821,N_3509,N_2470);
xnor U3822 (N_3822,N_3724,In_2024);
xnor U3823 (N_3823,N_2207,In_272);
xnor U3824 (N_3824,In_3678,In_4619);
and U3825 (N_3825,In_4451,N_1880);
nor U3826 (N_3826,In_4282,N_2773);
nor U3827 (N_3827,In_3422,N_3297);
xnor U3828 (N_3828,N_1975,N_514);
xnor U3829 (N_3829,N_3445,N_2198);
and U3830 (N_3830,N_2384,In_4017);
nor U3831 (N_3831,N_3025,In_1771);
xnor U3832 (N_3832,N_2818,N_2892);
and U3833 (N_3833,N_2473,N_82);
nand U3834 (N_3834,N_3741,N_3682);
nor U3835 (N_3835,N_1181,N_2964);
or U3836 (N_3836,N_3322,N_2831);
and U3837 (N_3837,N_3663,N_2200);
nand U3838 (N_3838,N_1750,In_4038);
or U3839 (N_3839,N_1635,N_3677);
or U3840 (N_3840,N_1535,N_2765);
xnor U3841 (N_3841,N_3318,N_3695);
xnor U3842 (N_3842,N_3696,N_3747);
nand U3843 (N_3843,N_1368,N_1476);
nor U3844 (N_3844,In_107,N_1351);
xnor U3845 (N_3845,N_1556,In_3514);
nor U3846 (N_3846,N_3112,N_3398);
xnor U3847 (N_3847,In_1415,N_3626);
or U3848 (N_3848,N_980,N_2309);
nand U3849 (N_3849,In_1551,N_2675);
nor U3850 (N_3850,N_3375,In_3205);
and U3851 (N_3851,N_3593,N_3039);
or U3852 (N_3852,In_2847,N_3623);
or U3853 (N_3853,N_1441,In_3561);
and U3854 (N_3854,N_2799,N_2800);
nand U3855 (N_3855,In_4729,N_3549);
xnor U3856 (N_3856,N_1140,N_1850);
xor U3857 (N_3857,N_3572,N_2231);
or U3858 (N_3858,N_2562,In_2834);
or U3859 (N_3859,N_3421,N_1445);
nor U3860 (N_3860,N_1972,N_3545);
or U3861 (N_3861,N_1660,N_2510);
xnor U3862 (N_3862,N_1873,In_3902);
nor U3863 (N_3863,N_3163,N_2726);
or U3864 (N_3864,N_3300,N_3619);
and U3865 (N_3865,N_1464,N_660);
xor U3866 (N_3866,N_2855,N_590);
nor U3867 (N_3867,N_131,N_3227);
or U3868 (N_3868,N_2848,In_1407);
nor U3869 (N_3869,N_3143,In_3138);
xnor U3870 (N_3870,N_2772,N_2141);
nor U3871 (N_3871,In_1264,In_4080);
nor U3872 (N_3872,N_2741,N_2749);
nand U3873 (N_3873,N_3516,N_3415);
xor U3874 (N_3874,In_2703,N_3600);
nand U3875 (N_3875,In_1862,In_3041);
or U3876 (N_3876,N_3399,N_3588);
xnor U3877 (N_3877,N_3294,N_989);
and U3878 (N_3878,In_1912,N_3364);
and U3879 (N_3879,N_2468,N_3587);
and U3880 (N_3880,N_2320,In_4221);
xnor U3881 (N_3881,N_2979,N_3412);
nor U3882 (N_3882,N_3483,N_3187);
xor U3883 (N_3883,In_2121,N_2930);
nand U3884 (N_3884,N_3748,N_2681);
and U3885 (N_3885,N_2734,In_2741);
or U3886 (N_3886,N_2591,In_3212);
xnor U3887 (N_3887,In_2067,N_2974);
and U3888 (N_3888,N_1696,In_273);
nor U3889 (N_3889,In_2810,In_1068);
and U3890 (N_3890,In_3620,In_731);
xnor U3891 (N_3891,N_2847,In_2308);
xor U3892 (N_3892,In_2590,N_3607);
nand U3893 (N_3893,N_2928,N_3254);
nor U3894 (N_3894,N_618,N_3265);
nand U3895 (N_3895,N_3590,N_2478);
nor U3896 (N_3896,N_2797,In_3745);
or U3897 (N_3897,N_3361,N_3273);
xnor U3898 (N_3898,N_64,N_3484);
and U3899 (N_3899,In_2520,N_776);
xor U3900 (N_3900,N_2552,N_3474);
nor U3901 (N_3901,N_1683,N_1622);
or U3902 (N_3902,N_3742,N_3327);
xnor U3903 (N_3903,N_3569,N_3105);
and U3904 (N_3904,N_943,In_2);
nor U3905 (N_3905,N_3485,N_1881);
and U3906 (N_3906,N_430,N_3260);
nor U3907 (N_3907,In_4331,In_3059);
nand U3908 (N_3908,N_2902,N_3672);
xnor U3909 (N_3909,N_3020,N_3583);
or U3910 (N_3910,N_3689,N_3447);
and U3911 (N_3911,N_2924,In_1099);
and U3912 (N_3912,N_277,N_3635);
nand U3913 (N_3913,N_3382,N_2702);
xor U3914 (N_3914,In_2450,N_2981);
nand U3915 (N_3915,N_3638,N_2875);
xor U3916 (N_3916,N_3728,In_1506);
nor U3917 (N_3917,N_1131,N_1171);
or U3918 (N_3918,N_3444,N_2985);
or U3919 (N_3919,N_3136,In_2480);
nor U3920 (N_3920,In_1166,In_115);
nand U3921 (N_3921,N_2856,N_2592);
or U3922 (N_3922,N_2796,N_2642);
or U3923 (N_3923,N_3514,N_3629);
or U3924 (N_3924,N_3621,N_2155);
and U3925 (N_3925,N_3631,In_307);
xnor U3926 (N_3926,N_3174,N_3154);
and U3927 (N_3927,N_3446,N_3315);
or U3928 (N_3928,N_2575,N_3684);
nor U3929 (N_3929,N_3562,In_2762);
xnor U3930 (N_3930,N_3135,N_3508);
and U3931 (N_3931,In_3064,N_2969);
nand U3932 (N_3932,In_2090,N_3480);
and U3933 (N_3933,N_3522,N_2383);
xor U3934 (N_3934,N_3530,N_3666);
nor U3935 (N_3935,N_1538,N_2212);
xnor U3936 (N_3936,N_3636,In_1707);
xnor U3937 (N_3937,N_3468,N_2988);
or U3938 (N_3938,N_3473,N_3015);
xnor U3939 (N_3939,N_3093,N_2755);
nand U3940 (N_3940,N_3668,N_3220);
nand U3941 (N_3941,N_3618,N_3707);
xnor U3942 (N_3942,In_3176,N_1434);
and U3943 (N_3943,N_3649,N_3650);
nand U3944 (N_3944,N_2717,N_3632);
nor U3945 (N_3945,N_2363,N_3687);
nand U3946 (N_3946,N_2103,N_2840);
and U3947 (N_3947,N_2885,N_3519);
and U3948 (N_3948,N_3658,In_4600);
nor U3949 (N_3949,N_2810,N_3452);
nor U3950 (N_3950,N_1589,N_3591);
nor U3951 (N_3951,In_2149,N_2096);
or U3952 (N_3952,N_2430,N_3598);
and U3953 (N_3953,N_289,N_2743);
nand U3954 (N_3954,N_2303,N_3496);
nand U3955 (N_3955,N_3288,N_2565);
nand U3956 (N_3956,N_760,N_3405);
or U3957 (N_3957,N_3090,In_965);
nand U3958 (N_3958,N_3716,N_3710);
xnor U3959 (N_3959,N_3573,N_3740);
xor U3960 (N_3960,N_594,N_3303);
xor U3961 (N_3961,In_3783,N_3489);
xor U3962 (N_3962,N_3221,N_3712);
and U3963 (N_3963,N_3609,N_3451);
or U3964 (N_3964,N_3290,N_2635);
nor U3965 (N_3965,N_3550,N_1483);
nand U3966 (N_3966,N_3694,N_3280);
and U3967 (N_3967,N_3596,N_3511);
and U3968 (N_3968,N_2104,N_2576);
xnor U3969 (N_3969,N_2857,In_3878);
or U3970 (N_3970,N_3553,In_3534);
nand U3971 (N_3971,N_936,N_1596);
and U3972 (N_3972,N_2242,In_110);
or U3973 (N_3973,N_3732,N_3531);
nor U3974 (N_3974,In_1694,In_1175);
nand U3975 (N_3975,N_3461,N_3200);
and U3976 (N_3976,N_539,In_2040);
nand U3977 (N_3977,N_877,N_3347);
and U3978 (N_3978,N_3330,N_2725);
and U3979 (N_3979,N_2649,N_3664);
and U3980 (N_3980,N_3380,N_3469);
nor U3981 (N_3981,N_3082,N_3479);
nand U3982 (N_3982,N_3701,N_2018);
nand U3983 (N_3983,N_175,N_1374);
nand U3984 (N_3984,N_3224,N_3449);
or U3985 (N_3985,N_2080,N_3559);
or U3986 (N_3986,N_3592,N_3620);
or U3987 (N_3987,N_3458,N_3350);
nor U3988 (N_3988,N_3356,N_918);
nand U3989 (N_3989,N_3674,In_711);
or U3990 (N_3990,N_1671,N_2711);
or U3991 (N_3991,N_1730,N_3540);
or U3992 (N_3992,N_3711,N_2626);
xnor U3993 (N_3993,N_3373,N_3086);
nand U3994 (N_3994,N_1584,N_1771);
xor U3995 (N_3995,N_3155,N_2460);
nand U3996 (N_3996,N_523,N_3113);
nor U3997 (N_3997,N_2977,N_2498);
or U3998 (N_3998,In_505,In_3800);
nor U3999 (N_3999,N_3686,N_3749);
nor U4000 (N_4000,N_3283,N_2353);
or U4001 (N_4001,In_4791,N_3106);
xnor U4002 (N_4002,N_3556,N_2012);
and U4003 (N_4003,N_3778,N_3230);
nand U4004 (N_4004,N_457,In_3956);
and U4005 (N_4005,N_3564,N_3467);
nor U4006 (N_4006,N_3440,N_3898);
or U4007 (N_4007,N_3993,N_3397);
and U4008 (N_4008,N_3585,N_3040);
nand U4009 (N_4009,N_3582,N_2890);
nor U4010 (N_4010,N_3402,In_4362);
or U4011 (N_4011,N_1267,N_3966);
nand U4012 (N_4012,N_3943,N_3680);
nor U4013 (N_4013,N_3080,N_2696);
and U4014 (N_4014,N_3932,N_3746);
nor U4015 (N_4015,N_3144,N_2707);
nor U4016 (N_4016,N_3907,In_3521);
nor U4017 (N_4017,N_3247,N_3949);
xor U4018 (N_4018,N_3130,N_2876);
or U4019 (N_4019,N_624,N_3810);
or U4020 (N_4020,N_3497,N_2422);
nor U4021 (N_4021,N_3611,N_3872);
nand U4022 (N_4022,N_3625,In_3688);
xnor U4023 (N_4023,N_3830,N_3643);
and U4024 (N_4024,N_483,N_3925);
or U4025 (N_4025,N_3782,N_3547);
nand U4026 (N_4026,N_2646,N_2907);
nand U4027 (N_4027,N_3339,N_2366);
nand U4028 (N_4028,N_3698,N_3800);
nand U4029 (N_4029,In_4841,N_3765);
nand U4030 (N_4030,N_3568,N_3852);
and U4031 (N_4031,In_155,N_3867);
nor U4032 (N_4032,N_2328,In_2940);
xnor U4033 (N_4033,N_3506,N_3945);
nor U4034 (N_4034,N_3690,N_2297);
xnor U4035 (N_4035,N_2171,N_3544);
xor U4036 (N_4036,N_3455,N_1104);
nor U4037 (N_4037,N_3216,N_3507);
or U4038 (N_4038,N_2244,N_2841);
nor U4039 (N_4039,N_3481,N_3752);
and U4040 (N_4040,N_3803,N_3194);
xnor U4041 (N_4041,In_2691,N_1877);
xnor U4042 (N_4042,In_4065,N_3879);
or U4043 (N_4043,N_3575,N_3868);
xor U4044 (N_4044,N_3574,N_3798);
nor U4045 (N_4045,N_3439,N_3845);
xor U4046 (N_4046,N_3697,N_3848);
nand U4047 (N_4047,N_768,N_631);
xnor U4048 (N_4048,N_2040,N_3476);
xnor U4049 (N_4049,N_744,N_3959);
xor U4050 (N_4050,N_3927,N_3148);
and U4051 (N_4051,N_3683,N_3608);
and U4052 (N_4052,N_3801,N_3018);
and U4053 (N_4053,N_2455,N_2706);
or U4054 (N_4054,N_112,N_3834);
or U4055 (N_4055,N_3119,N_2249);
xor U4056 (N_4056,N_3425,N_3442);
nand U4057 (N_4057,N_2753,N_3817);
or U4058 (N_4058,N_3994,N_3457);
and U4059 (N_4059,N_3827,N_2262);
or U4060 (N_4060,In_373,N_983);
and U4061 (N_4061,N_3081,N_3995);
nand U4062 (N_4062,N_3915,N_3358);
nand U4063 (N_4063,N_3877,N_3443);
and U4064 (N_4064,N_3614,N_2737);
nand U4065 (N_4065,In_2714,N_3630);
and U4066 (N_4066,N_1681,N_2677);
and U4067 (N_4067,N_4,N_3610);
xnor U4068 (N_4068,N_2816,N_3515);
or U4069 (N_4069,In_1948,N_3776);
nand U4070 (N_4070,N_3856,N_3902);
nand U4071 (N_4071,N_3414,N_3761);
or U4072 (N_4072,N_3423,N_835);
and U4073 (N_4073,N_3316,N_997);
and U4074 (N_4074,In_1482,N_3252);
nand U4075 (N_4075,N_1988,In_2117);
or U4076 (N_4076,N_3968,N_3910);
xor U4077 (N_4077,N_3804,In_3615);
nand U4078 (N_4078,N_763,N_1896);
or U4079 (N_4079,N_2260,N_2228);
xor U4080 (N_4080,N_3185,N_3859);
nor U4081 (N_4081,N_2782,N_2147);
nand U4082 (N_4082,In_1605,N_3652);
xnor U4083 (N_4083,N_3999,In_4675);
nand U4084 (N_4084,N_3802,N_3924);
xnor U4085 (N_4085,N_3870,N_3431);
or U4086 (N_4086,In_3233,N_3557);
or U4087 (N_4087,N_3826,N_1547);
xnor U4088 (N_4088,N_2358,N_1209);
nor U4089 (N_4089,N_2527,N_242);
nor U4090 (N_4090,N_2629,N_3849);
and U4091 (N_4091,N_3667,N_3796);
or U4092 (N_4092,N_3616,N_3997);
nor U4093 (N_4093,N_2373,N_3334);
xor U4094 (N_4094,N_3462,N_1214);
xnor U4095 (N_4095,N_3861,N_3678);
nand U4096 (N_4096,N_3759,N_3604);
xor U4097 (N_4097,N_3962,N_3754);
xor U4098 (N_4098,In_4423,N_3794);
xor U4099 (N_4099,N_3912,N_3895);
xnor U4100 (N_4100,N_3882,N_3745);
nor U4101 (N_4101,In_1459,N_3875);
or U4102 (N_4102,N_3987,N_2045);
or U4103 (N_4103,N_3107,N_3634);
nand U4104 (N_4104,N_3454,N_3864);
nand U4105 (N_4105,N_3843,N_3401);
and U4106 (N_4106,In_4978,N_1956);
nand U4107 (N_4107,N_1352,N_2884);
nand U4108 (N_4108,N_3068,N_3744);
xnor U4109 (N_4109,In_1989,N_3603);
nor U4110 (N_4110,N_3777,N_3679);
nand U4111 (N_4111,In_2626,N_2605);
or U4112 (N_4112,N_1105,N_3985);
and U4113 (N_4113,In_3505,In_1357);
and U4114 (N_4114,N_3259,N_2762);
xnor U4115 (N_4115,N_3411,N_3323);
and U4116 (N_4116,N_3881,N_2653);
or U4117 (N_4117,N_3577,N_3874);
nand U4118 (N_4118,N_3021,N_1759);
xnor U4119 (N_4119,In_2196,N_3639);
nand U4120 (N_4120,N_3073,N_3580);
nand U4121 (N_4121,N_2952,N_1212);
nand U4122 (N_4122,N_2877,N_3386);
xor U4123 (N_4123,N_3521,N_3967);
xor U4124 (N_4124,N_1560,N_3888);
xnor U4125 (N_4125,N_3896,N_3094);
or U4126 (N_4126,N_3726,N_3647);
and U4127 (N_4127,In_788,N_659);
or U4128 (N_4128,N_3858,N_3277);
or U4129 (N_4129,N_3219,N_3653);
nand U4130 (N_4130,N_3470,N_671);
nor U4131 (N_4131,N_3337,N_3739);
or U4132 (N_4132,N_2325,N_3369);
nor U4133 (N_4133,N_3756,N_3904);
or U4134 (N_4134,N_3757,N_3911);
nor U4135 (N_4135,N_3427,N_3863);
nor U4136 (N_4136,In_3704,N_1619);
nand U4137 (N_4137,N_858,In_260);
or U4138 (N_4138,N_2602,N_3151);
xor U4139 (N_4139,N_3751,N_3127);
and U4140 (N_4140,N_3942,N_3790);
or U4141 (N_4141,N_1234,N_3065);
xor U4142 (N_4142,N_3926,N_3525);
xnor U4143 (N_4143,N_3488,N_3542);
nor U4144 (N_4144,N_3899,N_3597);
nand U4145 (N_4145,N_3991,N_3561);
and U4146 (N_4146,N_773,N_3498);
nor U4147 (N_4147,N_3729,In_176);
or U4148 (N_4148,N_231,N_2145);
nor U4149 (N_4149,N_3492,N_3700);
or U4150 (N_4150,N_2333,N_3432);
nand U4151 (N_4151,N_2844,N_1698);
nand U4152 (N_4152,N_3880,N_1020);
xor U4153 (N_4153,In_1382,In_2296);
and U4154 (N_4154,N_2908,N_3111);
or U4155 (N_4155,N_2897,N_3816);
nor U4156 (N_4156,N_3887,N_3061);
and U4157 (N_4157,N_3860,In_4506);
and U4158 (N_4158,In_1981,N_2781);
nor U4159 (N_4159,N_3066,N_3383);
nand U4160 (N_4160,N_3972,N_2319);
nand U4161 (N_4161,N_3917,N_2572);
nor U4162 (N_4162,N_3785,N_3622);
xor U4163 (N_4163,N_3906,N_2511);
nand U4164 (N_4164,N_3964,N_465);
xor U4165 (N_4165,N_3873,N_3037);
nand U4166 (N_4166,N_3371,N_3957);
nor U4167 (N_4167,N_3532,N_3822);
nor U4168 (N_4168,N_3231,N_3022);
nor U4169 (N_4169,N_3971,N_2937);
nand U4170 (N_4170,In_2753,N_3718);
nand U4171 (N_4171,N_3946,N_3876);
nor U4172 (N_4172,N_2307,N_3787);
nor U4173 (N_4173,In_1477,N_3857);
nor U4174 (N_4174,N_2674,In_2700);
and U4175 (N_4175,N_811,In_2988);
nand U4176 (N_4176,N_3494,N_3797);
xor U4177 (N_4177,N_1206,In_3649);
xor U4178 (N_4178,N_1882,N_3951);
and U4179 (N_4179,N_3091,N_3842);
and U4180 (N_4180,N_931,N_3727);
nand U4181 (N_4181,In_830,N_3121);
xnor U4182 (N_4182,N_3702,N_3779);
or U4183 (N_4183,N_3520,N_1876);
nor U4184 (N_4184,N_2776,In_2909);
nor U4185 (N_4185,N_3372,N_3570);
nor U4186 (N_4186,In_3261,N_2972);
and U4187 (N_4187,N_3436,N_3685);
nor U4188 (N_4188,In_1703,N_3433);
and U4189 (N_4189,N_3963,N_3998);
nor U4190 (N_4190,N_1719,N_2247);
xor U4191 (N_4191,N_1574,N_3862);
and U4192 (N_4192,N_1147,N_3824);
xnor U4193 (N_4193,N_3929,N_3253);
or U4194 (N_4194,N_3633,In_4814);
xor U4195 (N_4195,N_2355,N_3813);
and U4196 (N_4196,N_3829,N_3973);
and U4197 (N_4197,N_3464,N_3837);
nand U4198 (N_4198,N_3517,N_17);
and U4199 (N_4199,N_2757,N_3450);
or U4200 (N_4200,N_1775,N_3589);
or U4201 (N_4201,In_2048,N_3342);
and U4202 (N_4202,N_3762,N_3933);
nor U4203 (N_4203,N_3846,N_2210);
or U4204 (N_4204,N_3548,In_3048);
xnor U4205 (N_4205,N_3996,In_3523);
nand U4206 (N_4206,In_3358,N_1409);
nor U4207 (N_4207,N_3546,N_3126);
and U4208 (N_4208,N_3976,N_3555);
nor U4209 (N_4209,N_3878,N_1831);
nand U4210 (N_4210,In_4924,N_1936);
and U4211 (N_4211,N_1796,N_3526);
nand U4212 (N_4212,In_2893,N_3275);
nor U4213 (N_4213,N_3387,N_3357);
and U4214 (N_4214,N_3145,N_3940);
nor U4215 (N_4215,N_3640,N_1959);
nor U4216 (N_4216,N_3518,N_3818);
and U4217 (N_4217,N_3814,N_3965);
and U4218 (N_4218,N_1591,N_572);
xor U4219 (N_4219,N_3605,N_3566);
xnor U4220 (N_4220,N_3390,N_2224);
and U4221 (N_4221,N_633,N_3908);
xnor U4222 (N_4222,N_1782,N_3983);
or U4223 (N_4223,In_1849,N_3730);
or U4224 (N_4224,N_3743,N_3919);
or U4225 (N_4225,N_1000,N_3952);
nand U4226 (N_4226,N_2731,In_4575);
nand U4227 (N_4227,N_3900,N_1217);
nand U4228 (N_4228,N_3897,N_3581);
nand U4229 (N_4229,N_3918,N_561);
nor U4230 (N_4230,N_1570,In_2416);
nand U4231 (N_4231,N_3660,N_3786);
xnor U4232 (N_4232,N_3955,N_3282);
xor U4233 (N_4233,N_3948,N_3007);
nand U4234 (N_4234,N_558,N_3502);
nand U4235 (N_4235,N_3708,N_3586);
or U4236 (N_4236,N_3990,N_3901);
or U4237 (N_4237,N_3770,N_3733);
nor U4238 (N_4238,N_3774,N_3978);
nand U4239 (N_4239,N_3602,N_2338);
xnor U4240 (N_4240,In_4713,In_582);
nor U4241 (N_4241,N_3031,N_3471);
xnor U4242 (N_4242,N_1029,In_2419);
and U4243 (N_4243,N_3753,N_3851);
nor U4244 (N_4244,In_329,N_3854);
nand U4245 (N_4245,N_3920,N_3270);
nor U4246 (N_4246,In_2170,N_2922);
nor U4247 (N_4247,In_2478,N_3975);
nor U4248 (N_4248,N_3289,N_3956);
nand U4249 (N_4249,N_804,N_2832);
nor U4250 (N_4250,N_3953,N_4016);
nor U4251 (N_4251,N_4027,N_3326);
or U4252 (N_4252,N_3676,N_4224);
or U4253 (N_4253,N_2233,N_3463);
or U4254 (N_4254,N_638,N_4155);
nand U4255 (N_4255,N_3871,N_4165);
and U4256 (N_4256,N_3961,N_4103);
xnor U4257 (N_4257,N_4189,N_1110);
xor U4258 (N_4258,N_4195,N_359);
or U4259 (N_4259,N_3341,N_3935);
nand U4260 (N_4260,N_4007,N_4194);
and U4261 (N_4261,N_4003,N_3268);
and U4262 (N_4262,N_4096,N_4204);
or U4263 (N_4263,N_4166,N_4218);
and U4264 (N_4264,N_2289,N_2108);
or U4265 (N_4265,N_3853,N_3768);
and U4266 (N_4266,N_3267,N_4219);
nand U4267 (N_4267,N_2127,N_4221);
or U4268 (N_4268,N_4029,In_2857);
and U4269 (N_4269,In_4855,N_3389);
nand U4270 (N_4270,N_4118,N_2914);
nor U4271 (N_4271,N_2011,N_4009);
or U4272 (N_4272,N_3560,N_4156);
nand U4273 (N_4273,N_3244,N_3370);
nor U4274 (N_4274,N_165,N_3805);
or U4275 (N_4275,N_1272,N_4105);
nand U4276 (N_4276,N_2203,N_4191);
or U4277 (N_4277,N_3536,N_3795);
xor U4278 (N_4278,In_790,N_3554);
or U4279 (N_4279,In_1521,N_2982);
and U4280 (N_4280,N_3374,N_4159);
xnor U4281 (N_4281,N_934,N_3922);
nor U4282 (N_4282,N_3847,N_3089);
and U4283 (N_4283,N_2923,N_2906);
xnor U4284 (N_4284,N_3395,In_428);
nor U4285 (N_4285,N_2229,N_3537);
nor U4286 (N_4286,In_4755,N_4059);
or U4287 (N_4287,N_4223,N_4053);
xnor U4288 (N_4288,In_2774,N_1674);
nor U4289 (N_4289,N_3841,N_3673);
nor U4290 (N_4290,N_3766,N_3019);
xnor U4291 (N_4291,N_1009,N_1031);
xor U4292 (N_4292,N_2476,N_3986);
nand U4293 (N_4293,N_4117,N_4070);
or U4294 (N_4294,N_3721,In_2773);
or U4295 (N_4295,In_3082,N_1933);
xnor U4296 (N_4296,N_4177,N_3735);
and U4297 (N_4297,N_3296,N_3764);
xnor U4298 (N_4298,N_1175,N_2268);
xor U4299 (N_4299,N_3806,N_4044);
nor U4300 (N_4300,N_4182,N_3763);
and U4301 (N_4301,N_3958,N_3850);
nand U4302 (N_4302,N_3913,N_3771);
and U4303 (N_4303,N_628,N_4169);
nor U4304 (N_4304,N_4056,N_3164);
nor U4305 (N_4305,N_2638,N_3723);
xnor U4306 (N_4306,In_4164,N_4081);
and U4307 (N_4307,N_634,In_3889);
or U4308 (N_4308,N_4222,N_3637);
and U4309 (N_4309,N_4023,In_856);
xor U4310 (N_4310,N_3487,N_2868);
and U4311 (N_4311,N_423,N_802);
or U4312 (N_4312,In_4682,N_4104);
nor U4313 (N_4313,In_19,N_187);
xnor U4314 (N_4314,N_4122,N_4208);
xor U4315 (N_4315,N_3171,N_4026);
or U4316 (N_4316,N_4022,N_3807);
and U4317 (N_4317,N_3256,N_3212);
xor U4318 (N_4318,N_2546,N_4030);
nand U4319 (N_4319,N_3923,N_4077);
nor U4320 (N_4320,N_40,N_3578);
nand U4321 (N_4321,N_3819,N_4212);
and U4322 (N_4322,N_4123,N_3459);
nand U4323 (N_4323,N_2348,N_2354);
nor U4324 (N_4324,N_3977,N_393);
nor U4325 (N_4325,N_3844,N_3429);
or U4326 (N_4326,N_3954,N_1032);
nor U4327 (N_4327,N_4227,N_4019);
nand U4328 (N_4328,N_3214,In_4335);
or U4329 (N_4329,N_2008,N_3098);
nand U4330 (N_4330,N_3947,N_3755);
nor U4331 (N_4331,N_3823,N_1243);
nand U4332 (N_4332,N_645,N_4137);
nor U4333 (N_4333,N_4057,N_3644);
nor U4334 (N_4334,N_754,N_1504);
nand U4335 (N_4335,N_3825,N_3974);
xor U4336 (N_4336,N_4141,N_4079);
nor U4337 (N_4337,N_3565,N_2222);
nand U4338 (N_4338,N_4179,N_4125);
xnor U4339 (N_4339,N_3980,N_3793);
xnor U4340 (N_4340,N_4184,In_4750);
xnor U4341 (N_4341,N_2786,N_4099);
or U4342 (N_4342,N_2544,N_3529);
nand U4343 (N_4343,N_4225,N_3513);
or U4344 (N_4344,N_4151,N_3176);
xnor U4345 (N_4345,N_2845,N_4051);
or U4346 (N_4346,N_3641,N_536);
and U4347 (N_4347,In_673,N_4013);
nor U4348 (N_4348,In_2944,N_282);
and U4349 (N_4349,N_4201,N_4094);
nor U4350 (N_4350,N_4163,N_4046);
nor U4351 (N_4351,N_1786,N_2750);
and U4352 (N_4352,N_1867,N_4097);
nor U4353 (N_4353,In_1462,In_2594);
nor U4354 (N_4354,N_3505,N_3328);
or U4355 (N_4355,N_4092,N_2395);
nor U4356 (N_4356,N_3982,N_4045);
nor U4357 (N_4357,N_3979,N_3240);
or U4358 (N_4358,In_33,N_3937);
and U4359 (N_4359,N_2401,N_4236);
nand U4360 (N_4360,N_4229,N_4232);
and U4361 (N_4361,N_3567,N_3349);
and U4362 (N_4362,N_4231,N_1633);
and U4363 (N_4363,N_3199,In_301);
xnor U4364 (N_4364,N_4149,N_3894);
nand U4365 (N_4365,In_4722,N_3936);
or U4366 (N_4366,N_2614,N_3831);
nor U4367 (N_4367,N_3760,N_4139);
nor U4368 (N_4368,N_3251,N_3969);
or U4369 (N_4369,N_3921,N_4213);
and U4370 (N_4370,N_4135,In_843);
xnor U4371 (N_4371,N_3309,N_4158);
or U4372 (N_4372,N_4124,N_494);
nand U4373 (N_4373,N_3775,In_4470);
xor U4374 (N_4374,N_4028,N_4199);
nor U4375 (N_4375,N_4090,N_2817);
and U4376 (N_4376,N_3799,N_4185);
nor U4377 (N_4377,N_3438,N_4072);
nand U4378 (N_4378,N_3909,N_3809);
nor U4379 (N_4379,N_4084,N_4054);
nand U4380 (N_4380,N_4032,N_1723);
and U4381 (N_4381,N_3734,N_4043);
nor U4382 (N_4382,N_4120,N_3914);
or U4383 (N_4383,N_3266,N_3033);
and U4384 (N_4384,N_4112,In_288);
and U4385 (N_4385,N_4113,N_1286);
and U4386 (N_4386,N_1643,N_4095);
nand U4387 (N_4387,N_3319,N_3886);
nand U4388 (N_4388,N_3885,In_2309);
nand U4389 (N_4389,N_4068,In_2960);
or U4390 (N_4390,N_3258,In_4666);
or U4391 (N_4391,N_3615,N_3928);
or U4392 (N_4392,N_4196,N_3543);
nor U4393 (N_4393,N_3836,N_4187);
nand U4394 (N_4394,N_3905,N_3197);
and U4395 (N_4395,N_3501,N_4154);
nand U4396 (N_4396,N_4237,N_3324);
or U4397 (N_4397,In_2692,N_2494);
or U4398 (N_4398,N_4065,N_1467);
xnor U4399 (N_4399,N_3791,N_3838);
or U4400 (N_4400,N_4146,N_3346);
nand U4401 (N_4401,In_3106,N_4198);
nor U4402 (N_4402,N_4167,N_4015);
or U4403 (N_4403,In_3888,N_4183);
nand U4404 (N_4404,N_1632,N_3884);
and U4405 (N_4405,N_4245,N_3193);
nor U4406 (N_4406,N_2846,N_2995);
and U4407 (N_4407,N_3731,N_2235);
nand U4408 (N_4408,N_3780,N_3448);
and U4409 (N_4409,N_3665,In_1580);
nand U4410 (N_4410,N_3365,N_3903);
xor U4411 (N_4411,N_2418,In_2557);
nand U4412 (N_4412,N_319,N_3528);
or U4413 (N_4413,N_4186,N_3408);
or U4414 (N_4414,N_4025,N_4173);
or U4415 (N_4415,N_4150,N_3422);
and U4416 (N_4416,N_3238,N_4210);
or U4417 (N_4417,N_4064,N_3722);
and U4418 (N_4418,N_4002,N_3645);
nor U4419 (N_4419,N_3828,N_3893);
nand U4420 (N_4420,N_2005,N_32);
nand U4421 (N_4421,In_4142,N_3992);
and U4422 (N_4422,N_3191,N_4087);
xor U4423 (N_4423,N_3892,N_2961);
nand U4424 (N_4424,N_4109,N_3250);
and U4425 (N_4425,N_2655,N_1809);
or U4426 (N_4426,In_1020,N_928);
nor U4427 (N_4427,N_4055,In_4344);
nand U4428 (N_4428,N_4101,N_4164);
or U4429 (N_4429,N_3720,N_1405);
or U4430 (N_4430,N_3839,N_4241);
xnor U4431 (N_4431,N_3407,N_4001);
nor U4432 (N_4432,N_79,In_2538);
and U4433 (N_4433,N_4134,N_1386);
xnor U4434 (N_4434,N_4133,N_3393);
nand U4435 (N_4435,N_4038,N_2253);
nor U4436 (N_4436,N_4217,N_4121);
nand U4437 (N_4437,N_4233,N_3656);
nand U4438 (N_4438,N_2942,N_3889);
nor U4439 (N_4439,N_3713,N_4178);
and U4440 (N_4440,N_3539,N_2417);
and U4441 (N_4441,N_4126,N_3426);
nor U4442 (N_4442,N_3551,N_3118);
and U4443 (N_4443,N_4153,N_3812);
nand U4444 (N_4444,N_4011,N_2350);
or U4445 (N_4445,N_4102,N_4136);
or U4446 (N_4446,N_4008,N_3527);
xor U4447 (N_4447,N_2349,N_4172);
xnor U4448 (N_4448,N_3655,N_1273);
xor U4449 (N_4449,N_2051,N_4010);
nor U4450 (N_4450,N_4106,In_688);
and U4451 (N_4451,N_3654,N_3612);
and U4452 (N_4452,N_3989,N_4215);
and U4453 (N_4453,N_3166,N_4000);
nor U4454 (N_4454,N_3773,In_4548);
or U4455 (N_4455,N_4176,In_4745);
or U4456 (N_4456,N_2958,N_3624);
nor U4457 (N_4457,N_4246,N_4180);
or U4458 (N_4458,N_3821,N_4047);
and U4459 (N_4459,N_4234,N_2956);
or U4460 (N_4460,N_4160,N_3891);
xnor U4461 (N_4461,N_1385,N_1166);
nand U4462 (N_4462,N_4004,N_4205);
or U4463 (N_4463,In_2173,N_3988);
nand U4464 (N_4464,N_3938,N_4203);
or U4465 (N_4465,N_3579,In_880);
nand U4466 (N_4466,N_3736,N_2761);
and U4467 (N_4467,N_2582,N_4220);
xor U4468 (N_4468,N_3538,N_3304);
or U4469 (N_4469,N_4131,N_4049);
and U4470 (N_4470,N_4076,N_2518);
nand U4471 (N_4471,N_2887,N_4039);
nor U4472 (N_4472,N_3681,N_4243);
or U4473 (N_4473,N_4089,N_3662);
xnor U4474 (N_4474,N_3495,N_3486);
xor U4475 (N_4475,N_3691,N_4129);
or U4476 (N_4476,N_1832,N_3725);
nand U4477 (N_4477,N_285,N_3278);
nand U4478 (N_4478,N_2298,N_4193);
or U4479 (N_4479,N_4140,In_2605);
and U4480 (N_4480,N_3043,N_3541);
and U4481 (N_4481,N_3029,N_4078);
or U4482 (N_4482,N_4037,N_4066);
xor U4483 (N_4483,N_2764,N_2187);
and U4484 (N_4484,N_4042,N_4052);
or U4485 (N_4485,In_4321,N_4247);
and U4486 (N_4486,In_3049,N_4181);
and U4487 (N_4487,N_4152,N_4238);
xor U4488 (N_4488,In_910,N_3325);
nand U4489 (N_4489,In_2219,N_1824);
nand U4490 (N_4490,N_4127,In_634);
nand U4491 (N_4491,In_4630,N_4216);
nor U4492 (N_4492,N_1186,N_3706);
xor U4493 (N_4493,N_4209,N_3767);
and U4494 (N_4494,In_2436,N_3628);
nor U4495 (N_4495,N_4075,N_944);
and U4496 (N_4496,N_3869,N_4188);
xnor U4497 (N_4497,N_3693,N_3104);
nor U4498 (N_4498,N_4200,N_4130);
nand U4499 (N_4499,N_4145,N_4114);
xnor U4500 (N_4500,N_2623,N_2259);
nor U4501 (N_4501,N_2472,N_4410);
nand U4502 (N_4502,N_4175,N_4297);
nand U4503 (N_4503,N_3239,N_4091);
nand U4504 (N_4504,N_4399,N_4372);
xor U4505 (N_4505,N_4487,N_4274);
xnor U4506 (N_4506,N_4479,N_4235);
nor U4507 (N_4507,N_4085,N_4414);
xnor U4508 (N_4508,N_4386,N_4481);
nor U4509 (N_4509,In_2777,N_4086);
nand U4510 (N_4510,N_4486,N_4317);
xor U4511 (N_4511,N_4431,N_4422);
nor U4512 (N_4512,N_4398,N_4263);
xor U4513 (N_4513,N_2771,N_4393);
xnor U4514 (N_4514,N_4282,N_2508);
nand U4515 (N_4515,N_4380,N_3051);
nor U4516 (N_4516,N_4285,N_4415);
and U4517 (N_4517,N_3840,In_4881);
nand U4518 (N_4518,N_4293,N_2669);
and U4519 (N_4519,N_4484,N_2684);
nand U4520 (N_4520,N_4465,N_4460);
nor U4521 (N_4521,In_328,N_4368);
nand U4522 (N_4522,N_4337,N_3142);
nor U4523 (N_4523,N_3970,N_3404);
or U4524 (N_4524,N_4424,N_3024);
nand U4525 (N_4525,N_4300,N_1672);
or U4526 (N_4526,N_3410,N_4192);
xnor U4527 (N_4527,N_3563,N_3420);
or U4528 (N_4528,N_2038,N_4271);
or U4529 (N_4529,N_4335,N_4423);
nor U4530 (N_4530,N_4311,N_4041);
nor U4531 (N_4531,N_4254,N_3074);
or U4532 (N_4532,N_3571,N_3883);
nor U4533 (N_4533,N_4275,N_2065);
and U4534 (N_4534,N_4017,N_4062);
or U4535 (N_4535,N_4093,N_4457);
nand U4536 (N_4536,N_4347,N_3331);
and U4537 (N_4537,N_4286,N_4403);
or U4538 (N_4538,N_4143,N_4338);
xnor U4539 (N_4539,N_3594,N_4387);
nand U4540 (N_4540,N_3329,In_2650);
and U4541 (N_4541,N_4379,N_4291);
nand U4542 (N_4542,N_2151,N_4144);
xor U4543 (N_4543,In_1826,N_4350);
xor U4544 (N_4544,N_4436,N_3950);
nor U4545 (N_4545,N_3595,N_4492);
or U4546 (N_4546,N_3811,In_4343);
or U4547 (N_4547,N_4331,N_4390);
xnor U4548 (N_4548,N_3815,N_4228);
nor U4549 (N_4549,N_3648,N_4313);
xor U4550 (N_4550,N_4268,N_4384);
xor U4551 (N_4551,N_4463,N_4314);
xnor U4552 (N_4552,N_4407,N_4248);
nand U4553 (N_4553,N_4394,N_129);
or U4554 (N_4554,N_4128,N_4269);
nor U4555 (N_4555,N_4466,N_1717);
nor U4556 (N_4556,N_4478,N_3535);
or U4557 (N_4557,N_4239,N_2587);
and U4558 (N_4558,N_3599,N_4467);
or U4559 (N_4559,N_4475,N_4437);
nand U4560 (N_4560,N_4207,N_3368);
and U4561 (N_4561,N_4294,N_3792);
nand U4562 (N_4562,N_4206,N_3783);
nor U4563 (N_4563,N_4342,N_4302);
nand U4564 (N_4564,N_4280,N_4388);
or U4565 (N_4565,N_4382,N_4443);
nor U4566 (N_4566,N_4288,In_481);
or U4567 (N_4567,N_3789,N_4434);
or U4568 (N_4568,N_4111,N_691);
xor U4569 (N_4569,N_4346,N_4345);
nor U4570 (N_4570,N_4284,N_3321);
nor U4571 (N_4571,N_4495,N_4416);
and U4572 (N_4572,N_4061,In_4139);
and U4573 (N_4573,N_4279,N_2327);
or U4574 (N_4574,N_4035,N_3512);
xnor U4575 (N_4575,N_4100,N_4489);
or U4576 (N_4576,N_3758,N_4276);
xor U4577 (N_4577,N_4267,N_4021);
nor U4578 (N_4578,N_4270,N_4354);
or U4579 (N_4579,N_3378,N_4340);
xnor U4580 (N_4580,N_4329,In_4098);
nor U4581 (N_4581,N_4107,N_3715);
nand U4582 (N_4582,In_8,N_3053);
nand U4583 (N_4583,N_3172,N_4355);
or U4584 (N_4584,N_4067,N_4447);
and U4585 (N_4585,N_4402,N_4454);
and U4586 (N_4586,N_4377,N_1562);
nand U4587 (N_4587,N_4411,N_4006);
or U4588 (N_4588,N_4162,N_4256);
nor U4589 (N_4589,N_4352,N_4366);
xnor U4590 (N_4590,N_4050,N_4080);
and U4591 (N_4591,N_3941,N_3781);
nor U4592 (N_4592,N_4308,In_3216);
nor U4593 (N_4593,N_4033,N_4365);
and U4594 (N_4594,N_4468,N_4230);
nor U4595 (N_4595,N_4496,N_4458);
nand U4596 (N_4596,N_4073,In_4302);
nand U4597 (N_4597,N_3659,N_4364);
nor U4598 (N_4598,N_3738,N_2794);
or U4599 (N_4599,N_4283,N_4473);
nand U4600 (N_4600,N_4483,N_3584);
or U4601 (N_4601,N_2118,In_2709);
xor U4602 (N_4602,N_4482,N_3661);
xor U4603 (N_4603,N_3016,N_4389);
nor U4604 (N_4604,N_4339,N_4452);
nor U4605 (N_4605,N_4369,N_4412);
or U4606 (N_4606,N_4119,N_4349);
nor U4607 (N_4607,In_492,N_4497);
nor U4608 (N_4608,N_4132,N_4353);
nor U4609 (N_4609,N_4252,N_3704);
nor U4610 (N_4610,N_3493,N_4014);
or U4611 (N_4611,N_4408,N_4323);
or U4612 (N_4612,N_4455,N_3558);
nand U4613 (N_4613,In_1994,N_4240);
and U4614 (N_4614,N_2024,N_4296);
nand U4615 (N_4615,N_3784,N_4448);
nand U4616 (N_4616,N_4295,N_76);
and U4617 (N_4617,N_3298,N_4383);
or U4618 (N_4618,N_4292,N_4110);
and U4619 (N_4619,N_4202,N_4381);
xor U4620 (N_4620,N_4453,N_4433);
nor U4621 (N_4621,N_4356,N_4397);
or U4622 (N_4622,N_2791,N_4494);
nand U4623 (N_4623,N_3890,N_2378);
xnor U4624 (N_4624,N_4357,N_4378);
or U4625 (N_4625,N_4305,N_3413);
nand U4626 (N_4626,N_4298,N_4083);
and U4627 (N_4627,N_1819,N_3353);
nand U4628 (N_4628,N_4063,N_3279);
xnor U4629 (N_4629,N_4316,N_4242);
xor U4630 (N_4630,N_4161,N_1505);
xnor U4631 (N_4631,N_4417,N_4405);
nor U4632 (N_4632,N_4438,In_1330);
nand U4633 (N_4633,In_2439,N_4088);
nor U4634 (N_4634,N_4024,N_4343);
nand U4635 (N_4635,N_366,In_4759);
or U4636 (N_4636,N_4020,N_4315);
nand U4637 (N_4637,N_2916,N_4264);
nand U4638 (N_4638,N_3601,N_4250);
xor U4639 (N_4639,N_3576,N_2308);
nor U4640 (N_4640,In_81,N_4012);
and U4641 (N_4641,N_4273,In_3319);
and U4642 (N_4642,N_4036,N_4082);
nand U4643 (N_4643,N_4429,N_3808);
and U4644 (N_4644,N_2361,N_4168);
nand U4645 (N_4645,In_848,N_3960);
nor U4646 (N_4646,N_3465,N_4450);
nand U4647 (N_4647,N_4476,N_2550);
xor U4648 (N_4648,In_3803,N_3606);
xnor U4649 (N_4649,N_4304,N_4490);
nor U4650 (N_4650,N_1783,N_4147);
or U4651 (N_4651,In_2790,N_4071);
nand U4652 (N_4652,N_1064,N_4048);
or U4653 (N_4653,N_4171,N_4174);
nor U4654 (N_4654,N_3934,N_3835);
nor U4655 (N_4655,N_4320,N_4058);
xnor U4656 (N_4656,N_4312,N_4018);
nor U4657 (N_4657,N_4303,N_4287);
and U4658 (N_4658,In_2963,N_3204);
xnor U4659 (N_4659,N_4318,N_4373);
or U4660 (N_4660,N_4170,In_3418);
or U4661 (N_4661,N_4469,N_1034);
xor U4662 (N_4662,N_3617,N_3866);
nand U4663 (N_4663,N_4306,N_4301);
nor U4664 (N_4664,N_3271,N_4461);
xor U4665 (N_4665,N_4261,N_783);
and U4666 (N_4666,N_3984,N_3944);
and U4667 (N_4667,N_4142,N_4251);
or U4668 (N_4668,N_4074,N_4328);
xnor U4669 (N_4669,N_4040,N_4257);
xor U4670 (N_4670,N_3651,N_4418);
nand U4671 (N_4671,N_4258,N_4148);
and U4672 (N_4672,N_4367,N_4472);
xnor U4673 (N_4673,N_4474,N_4098);
and U4674 (N_4674,N_4299,N_3613);
nand U4675 (N_4675,N_3737,N_3115);
and U4676 (N_4676,N_2758,N_4375);
or U4677 (N_4677,N_4442,N_4249);
nand U4678 (N_4678,N_3772,N_4259);
xor U4679 (N_4679,N_4360,N_4326);
xor U4680 (N_4680,N_2116,N_4435);
nand U4681 (N_4681,N_4499,N_4451);
or U4682 (N_4682,N_3855,N_4197);
and U4683 (N_4683,In_470,N_4376);
xor U4684 (N_4684,N_4395,N_4477);
xor U4685 (N_4685,N_2777,N_4464);
xor U4686 (N_4686,N_4255,In_4651);
or U4687 (N_4687,N_4060,N_4430);
nand U4688 (N_4688,N_4272,N_4440);
nor U4689 (N_4689,N_4444,N_4370);
or U4690 (N_4690,N_1489,N_4281);
and U4691 (N_4691,N_4488,N_4449);
nand U4692 (N_4692,N_3788,N_4266);
xnor U4693 (N_4693,N_3820,N_4470);
nand U4694 (N_4694,N_2423,N_4322);
nand U4695 (N_4695,N_4361,N_4363);
nand U4696 (N_4696,N_4498,N_4277);
nor U4697 (N_4697,N_3295,N_3939);
or U4698 (N_4698,In_1409,N_4348);
nor U4699 (N_4699,N_3299,N_4462);
or U4700 (N_4700,N_4432,N_4362);
or U4701 (N_4701,N_4359,N_4005);
or U4702 (N_4702,N_4392,N_4321);
xor U4703 (N_4703,N_4480,In_2883);
nor U4704 (N_4704,N_4253,N_4409);
xor U4705 (N_4705,N_3750,N_4324);
and U4706 (N_4706,N_4138,N_3286);
nand U4707 (N_4707,N_4351,N_4471);
nand U4708 (N_4708,N_4226,N_4336);
nand U4709 (N_4709,N_4401,N_606);
nand U4710 (N_4710,N_4265,N_4115);
or U4711 (N_4711,N_4446,N_4385);
nor U4712 (N_4712,N_4439,N_4244);
nand U4713 (N_4713,N_4413,N_2768);
nor U4714 (N_4714,N_3930,N_4325);
and U4715 (N_4715,N_4420,N_4491);
nand U4716 (N_4716,N_4419,N_4374);
xor U4717 (N_4717,N_4327,N_4358);
or U4718 (N_4718,N_4459,N_2577);
xnor U4719 (N_4719,N_4341,N_4214);
nor U4720 (N_4720,N_4108,N_4391);
nand U4721 (N_4721,N_4262,N_4034);
and U4722 (N_4722,N_4333,N_2689);
nor U4723 (N_4723,N_4427,N_3646);
or U4724 (N_4724,N_3769,N_4493);
nand U4725 (N_4725,N_4310,N_4445);
nand U4726 (N_4726,N_4031,N_2968);
xnor U4727 (N_4727,N_3657,In_912);
or U4728 (N_4728,N_3010,N_4441);
xor U4729 (N_4729,N_4309,N_4319);
nor U4730 (N_4730,N_4307,N_2789);
xnor U4731 (N_4731,N_4396,N_4456);
xnor U4732 (N_4732,N_4400,N_4290);
nand U4733 (N_4733,N_4289,N_4332);
or U4734 (N_4734,N_4116,N_4404);
xor U4735 (N_4735,N_3931,N_4485);
and U4736 (N_4736,N_4428,N_2584);
or U4737 (N_4737,In_1326,N_3832);
and U4738 (N_4738,N_3714,N_4190);
and U4739 (N_4739,In_4641,N_4157);
xnor U4740 (N_4740,N_3916,N_3523);
nand U4741 (N_4741,N_4260,N_4406);
xnor U4742 (N_4742,N_4330,N_4426);
or U4743 (N_4743,N_4344,In_3400);
nand U4744 (N_4744,N_4069,N_3833);
xor U4745 (N_4745,N_3981,N_4371);
or U4746 (N_4746,N_4278,N_4211);
nand U4747 (N_4747,N_2683,N_4425);
nand U4748 (N_4748,N_4421,N_4334);
nand U4749 (N_4749,N_3103,N_3865);
nor U4750 (N_4750,N_4652,N_4640);
nand U4751 (N_4751,N_4663,N_4621);
and U4752 (N_4752,N_4741,N_4556);
xnor U4753 (N_4753,N_4605,N_4705);
nand U4754 (N_4754,N_4505,N_4544);
or U4755 (N_4755,N_4537,N_4571);
nor U4756 (N_4756,N_4699,N_4515);
xor U4757 (N_4757,N_4600,N_4655);
nand U4758 (N_4758,N_4536,N_4518);
and U4759 (N_4759,N_4582,N_4688);
and U4760 (N_4760,N_4619,N_4674);
xnor U4761 (N_4761,N_4524,N_4501);
xnor U4762 (N_4762,N_4506,N_4716);
and U4763 (N_4763,N_4546,N_4570);
nor U4764 (N_4764,N_4586,N_4659);
or U4765 (N_4765,N_4539,N_4647);
nor U4766 (N_4766,N_4661,N_4511);
and U4767 (N_4767,N_4625,N_4743);
or U4768 (N_4768,N_4673,N_4660);
and U4769 (N_4769,N_4563,N_4599);
or U4770 (N_4770,N_4503,N_4612);
or U4771 (N_4771,N_4637,N_4709);
xor U4772 (N_4772,N_4560,N_4670);
nand U4773 (N_4773,N_4739,N_4692);
nor U4774 (N_4774,N_4644,N_4642);
or U4775 (N_4775,N_4729,N_4650);
nand U4776 (N_4776,N_4620,N_4579);
and U4777 (N_4777,N_4554,N_4545);
and U4778 (N_4778,N_4710,N_4725);
nor U4779 (N_4779,N_4575,N_4726);
nand U4780 (N_4780,N_4551,N_4658);
and U4781 (N_4781,N_4531,N_4684);
nor U4782 (N_4782,N_4541,N_4527);
nand U4783 (N_4783,N_4730,N_4580);
nor U4784 (N_4784,N_4578,N_4685);
nor U4785 (N_4785,N_4606,N_4689);
or U4786 (N_4786,N_4628,N_4549);
xor U4787 (N_4787,N_4649,N_4616);
xor U4788 (N_4788,N_4508,N_4698);
or U4789 (N_4789,N_4717,N_4576);
or U4790 (N_4790,N_4588,N_4744);
or U4791 (N_4791,N_4559,N_4585);
or U4792 (N_4792,N_4636,N_4617);
nand U4793 (N_4793,N_4533,N_4596);
nand U4794 (N_4794,N_4645,N_4747);
xnor U4795 (N_4795,N_4614,N_4706);
nand U4796 (N_4796,N_4548,N_4566);
nor U4797 (N_4797,N_4603,N_4514);
nor U4798 (N_4798,N_4662,N_4654);
and U4799 (N_4799,N_4629,N_4722);
xor U4800 (N_4800,N_4607,N_4540);
and U4801 (N_4801,N_4587,N_4610);
or U4802 (N_4802,N_4723,N_4589);
nor U4803 (N_4803,N_4719,N_4641);
xor U4804 (N_4804,N_4535,N_4569);
and U4805 (N_4805,N_4721,N_4510);
nand U4806 (N_4806,N_4639,N_4746);
and U4807 (N_4807,N_4622,N_4601);
xor U4808 (N_4808,N_4704,N_4609);
and U4809 (N_4809,N_4665,N_4550);
and U4810 (N_4810,N_4532,N_4517);
and U4811 (N_4811,N_4718,N_4568);
nand U4812 (N_4812,N_4565,N_4555);
nor U4813 (N_4813,N_4552,N_4562);
xor U4814 (N_4814,N_4664,N_4584);
nand U4815 (N_4815,N_4651,N_4693);
xor U4816 (N_4816,N_4543,N_4690);
or U4817 (N_4817,N_4516,N_4736);
nand U4818 (N_4818,N_4525,N_4681);
xnor U4819 (N_4819,N_4509,N_4627);
nand U4820 (N_4820,N_4683,N_4731);
nand U4821 (N_4821,N_4737,N_4695);
xor U4822 (N_4822,N_4679,N_4686);
or U4823 (N_4823,N_4748,N_4523);
nor U4824 (N_4824,N_4703,N_4595);
or U4825 (N_4825,N_4635,N_4590);
nand U4826 (N_4826,N_4672,N_4745);
nand U4827 (N_4827,N_4526,N_4694);
nor U4828 (N_4828,N_4522,N_4631);
nor U4829 (N_4829,N_4656,N_4702);
nand U4830 (N_4830,N_4538,N_4643);
xnor U4831 (N_4831,N_4696,N_4597);
and U4832 (N_4832,N_4675,N_4502);
nor U4833 (N_4833,N_4734,N_4712);
xnor U4834 (N_4834,N_4504,N_4500);
nor U4835 (N_4835,N_4707,N_4604);
and U4836 (N_4836,N_4715,N_4733);
nor U4837 (N_4837,N_4700,N_4680);
nand U4838 (N_4838,N_4667,N_4732);
and U4839 (N_4839,N_4713,N_4691);
and U4840 (N_4840,N_4611,N_4735);
or U4841 (N_4841,N_4558,N_4534);
and U4842 (N_4842,N_4564,N_4615);
xor U4843 (N_4843,N_4697,N_4520);
nand U4844 (N_4844,N_4714,N_4711);
nand U4845 (N_4845,N_4676,N_4653);
or U4846 (N_4846,N_4521,N_4646);
and U4847 (N_4847,N_4574,N_4687);
xnor U4848 (N_4848,N_4630,N_4572);
nand U4849 (N_4849,N_4677,N_4530);
nor U4850 (N_4850,N_4618,N_4528);
nor U4851 (N_4851,N_4624,N_4593);
or U4852 (N_4852,N_4720,N_4547);
nand U4853 (N_4853,N_4613,N_4633);
xnor U4854 (N_4854,N_4632,N_4738);
and U4855 (N_4855,N_4634,N_4671);
and U4856 (N_4856,N_4657,N_4742);
or U4857 (N_4857,N_4749,N_4567);
and U4858 (N_4858,N_4701,N_4727);
nand U4859 (N_4859,N_4638,N_4592);
and U4860 (N_4860,N_4561,N_4594);
nand U4861 (N_4861,N_4581,N_4728);
nand U4862 (N_4862,N_4668,N_4708);
nor U4863 (N_4863,N_4623,N_4666);
or U4864 (N_4864,N_4583,N_4682);
or U4865 (N_4865,N_4591,N_4529);
and U4866 (N_4866,N_4513,N_4573);
nand U4867 (N_4867,N_4678,N_4648);
or U4868 (N_4868,N_4724,N_4557);
or U4869 (N_4869,N_4512,N_4740);
and U4870 (N_4870,N_4542,N_4602);
and U4871 (N_4871,N_4598,N_4608);
nor U4872 (N_4872,N_4507,N_4669);
xnor U4873 (N_4873,N_4577,N_4553);
nand U4874 (N_4874,N_4519,N_4626);
or U4875 (N_4875,N_4626,N_4740);
nand U4876 (N_4876,N_4501,N_4690);
nand U4877 (N_4877,N_4604,N_4685);
xor U4878 (N_4878,N_4629,N_4532);
or U4879 (N_4879,N_4563,N_4639);
nand U4880 (N_4880,N_4625,N_4667);
nand U4881 (N_4881,N_4679,N_4510);
xnor U4882 (N_4882,N_4589,N_4630);
and U4883 (N_4883,N_4549,N_4576);
or U4884 (N_4884,N_4674,N_4524);
and U4885 (N_4885,N_4500,N_4545);
nand U4886 (N_4886,N_4611,N_4602);
nor U4887 (N_4887,N_4556,N_4581);
xor U4888 (N_4888,N_4520,N_4502);
or U4889 (N_4889,N_4677,N_4578);
and U4890 (N_4890,N_4711,N_4550);
nand U4891 (N_4891,N_4650,N_4514);
or U4892 (N_4892,N_4514,N_4609);
and U4893 (N_4893,N_4602,N_4704);
xnor U4894 (N_4894,N_4558,N_4693);
xor U4895 (N_4895,N_4507,N_4663);
and U4896 (N_4896,N_4647,N_4553);
nand U4897 (N_4897,N_4542,N_4726);
nand U4898 (N_4898,N_4564,N_4654);
nand U4899 (N_4899,N_4526,N_4529);
nand U4900 (N_4900,N_4657,N_4557);
and U4901 (N_4901,N_4630,N_4547);
and U4902 (N_4902,N_4573,N_4516);
nor U4903 (N_4903,N_4517,N_4653);
xnor U4904 (N_4904,N_4634,N_4648);
xnor U4905 (N_4905,N_4733,N_4577);
nor U4906 (N_4906,N_4629,N_4598);
or U4907 (N_4907,N_4522,N_4617);
nor U4908 (N_4908,N_4569,N_4743);
xor U4909 (N_4909,N_4663,N_4696);
nand U4910 (N_4910,N_4746,N_4675);
nand U4911 (N_4911,N_4708,N_4717);
nor U4912 (N_4912,N_4513,N_4586);
xor U4913 (N_4913,N_4591,N_4560);
nand U4914 (N_4914,N_4683,N_4740);
nor U4915 (N_4915,N_4657,N_4733);
nand U4916 (N_4916,N_4638,N_4712);
xor U4917 (N_4917,N_4612,N_4502);
xnor U4918 (N_4918,N_4746,N_4622);
xor U4919 (N_4919,N_4575,N_4694);
nand U4920 (N_4920,N_4684,N_4665);
or U4921 (N_4921,N_4607,N_4567);
xor U4922 (N_4922,N_4707,N_4745);
nand U4923 (N_4923,N_4690,N_4507);
nand U4924 (N_4924,N_4503,N_4630);
nor U4925 (N_4925,N_4673,N_4656);
nand U4926 (N_4926,N_4568,N_4529);
nor U4927 (N_4927,N_4552,N_4697);
or U4928 (N_4928,N_4712,N_4627);
and U4929 (N_4929,N_4556,N_4689);
or U4930 (N_4930,N_4638,N_4736);
nor U4931 (N_4931,N_4645,N_4521);
nand U4932 (N_4932,N_4519,N_4520);
nand U4933 (N_4933,N_4731,N_4560);
nor U4934 (N_4934,N_4550,N_4646);
and U4935 (N_4935,N_4558,N_4624);
nor U4936 (N_4936,N_4597,N_4685);
and U4937 (N_4937,N_4720,N_4634);
nand U4938 (N_4938,N_4695,N_4533);
xnor U4939 (N_4939,N_4564,N_4701);
or U4940 (N_4940,N_4582,N_4523);
or U4941 (N_4941,N_4502,N_4618);
and U4942 (N_4942,N_4602,N_4736);
and U4943 (N_4943,N_4641,N_4732);
nand U4944 (N_4944,N_4559,N_4646);
nand U4945 (N_4945,N_4682,N_4743);
or U4946 (N_4946,N_4732,N_4702);
xnor U4947 (N_4947,N_4744,N_4722);
nor U4948 (N_4948,N_4709,N_4502);
nand U4949 (N_4949,N_4663,N_4582);
and U4950 (N_4950,N_4529,N_4622);
nor U4951 (N_4951,N_4709,N_4607);
and U4952 (N_4952,N_4544,N_4688);
or U4953 (N_4953,N_4646,N_4539);
and U4954 (N_4954,N_4578,N_4501);
nor U4955 (N_4955,N_4657,N_4697);
and U4956 (N_4956,N_4534,N_4744);
nor U4957 (N_4957,N_4735,N_4608);
or U4958 (N_4958,N_4562,N_4546);
xnor U4959 (N_4959,N_4732,N_4677);
or U4960 (N_4960,N_4555,N_4545);
and U4961 (N_4961,N_4721,N_4502);
nor U4962 (N_4962,N_4584,N_4593);
nor U4963 (N_4963,N_4645,N_4630);
or U4964 (N_4964,N_4659,N_4693);
and U4965 (N_4965,N_4664,N_4585);
nor U4966 (N_4966,N_4517,N_4716);
nor U4967 (N_4967,N_4594,N_4573);
nand U4968 (N_4968,N_4593,N_4706);
nor U4969 (N_4969,N_4561,N_4508);
nor U4970 (N_4970,N_4733,N_4549);
or U4971 (N_4971,N_4727,N_4539);
and U4972 (N_4972,N_4747,N_4568);
nand U4973 (N_4973,N_4665,N_4703);
or U4974 (N_4974,N_4510,N_4637);
xnor U4975 (N_4975,N_4543,N_4700);
nand U4976 (N_4976,N_4608,N_4592);
nor U4977 (N_4977,N_4506,N_4607);
nor U4978 (N_4978,N_4629,N_4565);
nor U4979 (N_4979,N_4710,N_4584);
and U4980 (N_4980,N_4566,N_4742);
xnor U4981 (N_4981,N_4587,N_4667);
and U4982 (N_4982,N_4601,N_4658);
and U4983 (N_4983,N_4664,N_4666);
nor U4984 (N_4984,N_4631,N_4614);
nor U4985 (N_4985,N_4524,N_4536);
nor U4986 (N_4986,N_4504,N_4618);
or U4987 (N_4987,N_4715,N_4729);
xnor U4988 (N_4988,N_4506,N_4603);
nand U4989 (N_4989,N_4510,N_4588);
nor U4990 (N_4990,N_4567,N_4585);
or U4991 (N_4991,N_4525,N_4555);
nand U4992 (N_4992,N_4694,N_4623);
nand U4993 (N_4993,N_4700,N_4609);
xor U4994 (N_4994,N_4716,N_4739);
nor U4995 (N_4995,N_4632,N_4561);
nand U4996 (N_4996,N_4734,N_4673);
nor U4997 (N_4997,N_4690,N_4522);
nand U4998 (N_4998,N_4703,N_4642);
or U4999 (N_4999,N_4556,N_4675);
or U5000 (N_5000,N_4775,N_4803);
or U5001 (N_5001,N_4819,N_4813);
or U5002 (N_5002,N_4917,N_4780);
nor U5003 (N_5003,N_4792,N_4930);
and U5004 (N_5004,N_4798,N_4883);
nor U5005 (N_5005,N_4990,N_4956);
nor U5006 (N_5006,N_4997,N_4827);
xnor U5007 (N_5007,N_4874,N_4943);
nand U5008 (N_5008,N_4824,N_4757);
nand U5009 (N_5009,N_4880,N_4876);
xor U5010 (N_5010,N_4981,N_4987);
nor U5011 (N_5011,N_4751,N_4994);
and U5012 (N_5012,N_4832,N_4758);
nand U5013 (N_5013,N_4753,N_4933);
and U5014 (N_5014,N_4769,N_4999);
nand U5015 (N_5015,N_4946,N_4841);
nor U5016 (N_5016,N_4783,N_4910);
or U5017 (N_5017,N_4977,N_4960);
nor U5018 (N_5018,N_4888,N_4844);
nand U5019 (N_5019,N_4834,N_4790);
and U5020 (N_5020,N_4872,N_4816);
nor U5021 (N_5021,N_4772,N_4965);
nand U5022 (N_5022,N_4750,N_4756);
or U5023 (N_5023,N_4825,N_4829);
nor U5024 (N_5024,N_4897,N_4856);
or U5025 (N_5025,N_4887,N_4864);
nor U5026 (N_5026,N_4967,N_4919);
or U5027 (N_5027,N_4858,N_4988);
nand U5028 (N_5028,N_4791,N_4935);
nor U5029 (N_5029,N_4848,N_4926);
or U5030 (N_5030,N_4823,N_4921);
xnor U5031 (N_5031,N_4770,N_4922);
or U5032 (N_5032,N_4854,N_4940);
xnor U5033 (N_5033,N_4972,N_4774);
and U5034 (N_5034,N_4773,N_4826);
nand U5035 (N_5035,N_4925,N_4948);
xor U5036 (N_5036,N_4971,N_4879);
xnor U5037 (N_5037,N_4916,N_4853);
or U5038 (N_5038,N_4920,N_4797);
nand U5039 (N_5039,N_4809,N_4914);
nor U5040 (N_5040,N_4942,N_4964);
nor U5041 (N_5041,N_4934,N_4955);
or U5042 (N_5042,N_4953,N_4855);
nor U5043 (N_5043,N_4982,N_4763);
nor U5044 (N_5044,N_4878,N_4839);
nand U5045 (N_5045,N_4966,N_4939);
nand U5046 (N_5046,N_4808,N_4898);
or U5047 (N_5047,N_4833,N_4998);
or U5048 (N_5048,N_4850,N_4995);
nor U5049 (N_5049,N_4800,N_4785);
or U5050 (N_5050,N_4868,N_4909);
xor U5051 (N_5051,N_4821,N_4820);
and U5052 (N_5052,N_4817,N_4822);
and U5053 (N_5053,N_4993,N_4895);
and U5054 (N_5054,N_4885,N_4985);
xnor U5055 (N_5055,N_4996,N_4802);
nor U5056 (N_5056,N_4899,N_4959);
or U5057 (N_5057,N_4900,N_4976);
and U5058 (N_5058,N_4860,N_4886);
and U5059 (N_5059,N_4947,N_4804);
and U5060 (N_5060,N_4840,N_4782);
xnor U5061 (N_5061,N_4866,N_4957);
nor U5062 (N_5062,N_4924,N_4784);
and U5063 (N_5063,N_4807,N_4811);
or U5064 (N_5064,N_4873,N_4755);
nor U5065 (N_5065,N_4903,N_4881);
nand U5066 (N_5066,N_4905,N_4944);
nor U5067 (N_5067,N_4845,N_4799);
or U5068 (N_5068,N_4892,N_4830);
or U5069 (N_5069,N_4768,N_4975);
nor U5070 (N_5070,N_4787,N_4893);
nand U5071 (N_5071,N_4989,N_4952);
or U5072 (N_5072,N_4950,N_4867);
or U5073 (N_5073,N_4901,N_4896);
xnor U5074 (N_5074,N_4894,N_4906);
or U5075 (N_5075,N_4777,N_4847);
nor U5076 (N_5076,N_4761,N_4870);
nor U5077 (N_5077,N_4961,N_4986);
nor U5078 (N_5078,N_4875,N_4983);
xor U5079 (N_5079,N_4907,N_4781);
nand U5080 (N_5080,N_4945,N_4932);
nor U5081 (N_5081,N_4857,N_4902);
and U5082 (N_5082,N_4871,N_4980);
or U5083 (N_5083,N_4764,N_4759);
or U5084 (N_5084,N_4915,N_4806);
or U5085 (N_5085,N_4937,N_4836);
xor U5086 (N_5086,N_4795,N_4978);
xor U5087 (N_5087,N_4936,N_4815);
nor U5088 (N_5088,N_4814,N_4812);
and U5089 (N_5089,N_4851,N_4890);
xnor U5090 (N_5090,N_4911,N_4818);
and U5091 (N_5091,N_4969,N_4954);
nand U5092 (N_5092,N_4970,N_4865);
and U5093 (N_5093,N_4929,N_4789);
nor U5094 (N_5094,N_4891,N_4863);
xor U5095 (N_5095,N_4928,N_4776);
nand U5096 (N_5096,N_4913,N_4831);
xnor U5097 (N_5097,N_4838,N_4778);
and U5098 (N_5098,N_4835,N_4918);
or U5099 (N_5099,N_4912,N_4752);
or U5100 (N_5100,N_4766,N_4882);
and U5101 (N_5101,N_4992,N_4767);
and U5102 (N_5102,N_4877,N_4762);
nor U5103 (N_5103,N_4810,N_4842);
xnor U5104 (N_5104,N_4968,N_4837);
nand U5105 (N_5105,N_4904,N_4771);
xor U5106 (N_5106,N_4931,N_4859);
xnor U5107 (N_5107,N_4793,N_4884);
nand U5108 (N_5108,N_4941,N_4786);
or U5109 (N_5109,N_4979,N_4796);
xnor U5110 (N_5110,N_4927,N_4849);
nand U5111 (N_5111,N_4794,N_4962);
xnor U5112 (N_5112,N_4938,N_4923);
nand U5113 (N_5113,N_4805,N_4779);
nor U5114 (N_5114,N_4908,N_4852);
or U5115 (N_5115,N_4974,N_4754);
or U5116 (N_5116,N_4958,N_4843);
and U5117 (N_5117,N_4963,N_4869);
xor U5118 (N_5118,N_4760,N_4801);
nor U5119 (N_5119,N_4861,N_4889);
xor U5120 (N_5120,N_4984,N_4973);
nor U5121 (N_5121,N_4765,N_4949);
nor U5122 (N_5122,N_4846,N_4991);
nor U5123 (N_5123,N_4828,N_4951);
nor U5124 (N_5124,N_4862,N_4788);
nand U5125 (N_5125,N_4830,N_4914);
xnor U5126 (N_5126,N_4815,N_4979);
and U5127 (N_5127,N_4805,N_4982);
nand U5128 (N_5128,N_4941,N_4784);
xnor U5129 (N_5129,N_4807,N_4953);
and U5130 (N_5130,N_4810,N_4915);
nand U5131 (N_5131,N_4823,N_4856);
xor U5132 (N_5132,N_4756,N_4781);
and U5133 (N_5133,N_4941,N_4902);
nor U5134 (N_5134,N_4750,N_4852);
and U5135 (N_5135,N_4976,N_4915);
and U5136 (N_5136,N_4876,N_4836);
and U5137 (N_5137,N_4856,N_4936);
nor U5138 (N_5138,N_4804,N_4993);
and U5139 (N_5139,N_4757,N_4844);
or U5140 (N_5140,N_4987,N_4866);
nor U5141 (N_5141,N_4821,N_4787);
xor U5142 (N_5142,N_4804,N_4906);
and U5143 (N_5143,N_4889,N_4801);
and U5144 (N_5144,N_4952,N_4808);
nor U5145 (N_5145,N_4951,N_4935);
xnor U5146 (N_5146,N_4917,N_4905);
or U5147 (N_5147,N_4816,N_4809);
xor U5148 (N_5148,N_4996,N_4927);
nor U5149 (N_5149,N_4861,N_4913);
nor U5150 (N_5150,N_4936,N_4930);
or U5151 (N_5151,N_4777,N_4759);
or U5152 (N_5152,N_4837,N_4977);
nor U5153 (N_5153,N_4967,N_4781);
and U5154 (N_5154,N_4913,N_4794);
nand U5155 (N_5155,N_4846,N_4915);
and U5156 (N_5156,N_4846,N_4894);
xor U5157 (N_5157,N_4846,N_4824);
nand U5158 (N_5158,N_4810,N_4968);
or U5159 (N_5159,N_4828,N_4986);
xor U5160 (N_5160,N_4804,N_4772);
and U5161 (N_5161,N_4954,N_4951);
or U5162 (N_5162,N_4793,N_4796);
nand U5163 (N_5163,N_4759,N_4904);
or U5164 (N_5164,N_4769,N_4922);
and U5165 (N_5165,N_4877,N_4823);
or U5166 (N_5166,N_4857,N_4812);
nor U5167 (N_5167,N_4932,N_4931);
nand U5168 (N_5168,N_4903,N_4914);
nor U5169 (N_5169,N_4850,N_4849);
nand U5170 (N_5170,N_4975,N_4961);
and U5171 (N_5171,N_4998,N_4805);
nand U5172 (N_5172,N_4991,N_4892);
xnor U5173 (N_5173,N_4755,N_4968);
or U5174 (N_5174,N_4796,N_4976);
nand U5175 (N_5175,N_4871,N_4894);
and U5176 (N_5176,N_4906,N_4910);
nand U5177 (N_5177,N_4776,N_4767);
and U5178 (N_5178,N_4956,N_4959);
nor U5179 (N_5179,N_4750,N_4783);
or U5180 (N_5180,N_4802,N_4988);
nor U5181 (N_5181,N_4852,N_4935);
and U5182 (N_5182,N_4816,N_4778);
or U5183 (N_5183,N_4882,N_4961);
or U5184 (N_5184,N_4766,N_4935);
and U5185 (N_5185,N_4970,N_4869);
nand U5186 (N_5186,N_4818,N_4762);
xor U5187 (N_5187,N_4795,N_4838);
nand U5188 (N_5188,N_4893,N_4808);
or U5189 (N_5189,N_4958,N_4985);
and U5190 (N_5190,N_4856,N_4923);
and U5191 (N_5191,N_4867,N_4777);
xor U5192 (N_5192,N_4938,N_4859);
xnor U5193 (N_5193,N_4900,N_4894);
and U5194 (N_5194,N_4899,N_4982);
nand U5195 (N_5195,N_4888,N_4801);
and U5196 (N_5196,N_4853,N_4851);
xor U5197 (N_5197,N_4934,N_4963);
nand U5198 (N_5198,N_4958,N_4780);
and U5199 (N_5199,N_4922,N_4930);
xor U5200 (N_5200,N_4809,N_4912);
nand U5201 (N_5201,N_4915,N_4939);
xor U5202 (N_5202,N_4802,N_4790);
or U5203 (N_5203,N_4802,N_4754);
and U5204 (N_5204,N_4969,N_4773);
or U5205 (N_5205,N_4815,N_4950);
nor U5206 (N_5206,N_4990,N_4866);
nand U5207 (N_5207,N_4920,N_4823);
nor U5208 (N_5208,N_4834,N_4974);
nor U5209 (N_5209,N_4847,N_4972);
or U5210 (N_5210,N_4770,N_4995);
xor U5211 (N_5211,N_4829,N_4792);
nand U5212 (N_5212,N_4811,N_4949);
nor U5213 (N_5213,N_4920,N_4980);
nand U5214 (N_5214,N_4825,N_4925);
and U5215 (N_5215,N_4963,N_4992);
xnor U5216 (N_5216,N_4950,N_4807);
nand U5217 (N_5217,N_4972,N_4818);
or U5218 (N_5218,N_4968,N_4893);
xnor U5219 (N_5219,N_4959,N_4753);
nand U5220 (N_5220,N_4978,N_4961);
and U5221 (N_5221,N_4992,N_4881);
xor U5222 (N_5222,N_4977,N_4886);
and U5223 (N_5223,N_4825,N_4919);
and U5224 (N_5224,N_4897,N_4807);
and U5225 (N_5225,N_4946,N_4778);
xnor U5226 (N_5226,N_4991,N_4997);
and U5227 (N_5227,N_4971,N_4803);
or U5228 (N_5228,N_4901,N_4965);
nand U5229 (N_5229,N_4813,N_4834);
xnor U5230 (N_5230,N_4882,N_4950);
or U5231 (N_5231,N_4993,N_4920);
nor U5232 (N_5232,N_4948,N_4995);
nor U5233 (N_5233,N_4932,N_4933);
or U5234 (N_5234,N_4951,N_4800);
and U5235 (N_5235,N_4753,N_4837);
nor U5236 (N_5236,N_4888,N_4815);
and U5237 (N_5237,N_4771,N_4892);
and U5238 (N_5238,N_4952,N_4940);
xor U5239 (N_5239,N_4919,N_4984);
nand U5240 (N_5240,N_4841,N_4911);
nor U5241 (N_5241,N_4932,N_4966);
nor U5242 (N_5242,N_4962,N_4933);
and U5243 (N_5243,N_4908,N_4981);
and U5244 (N_5244,N_4838,N_4915);
and U5245 (N_5245,N_4993,N_4915);
or U5246 (N_5246,N_4822,N_4851);
nor U5247 (N_5247,N_4839,N_4939);
and U5248 (N_5248,N_4881,N_4978);
nor U5249 (N_5249,N_4836,N_4933);
xor U5250 (N_5250,N_5208,N_5196);
and U5251 (N_5251,N_5005,N_5008);
xor U5252 (N_5252,N_5009,N_5175);
xnor U5253 (N_5253,N_5240,N_5126);
nand U5254 (N_5254,N_5099,N_5104);
nand U5255 (N_5255,N_5153,N_5167);
nor U5256 (N_5256,N_5101,N_5039);
xor U5257 (N_5257,N_5030,N_5195);
nand U5258 (N_5258,N_5166,N_5025);
xnor U5259 (N_5259,N_5011,N_5088);
and U5260 (N_5260,N_5220,N_5109);
and U5261 (N_5261,N_5181,N_5085);
xor U5262 (N_5262,N_5211,N_5115);
or U5263 (N_5263,N_5031,N_5243);
nor U5264 (N_5264,N_5040,N_5178);
or U5265 (N_5265,N_5065,N_5245);
or U5266 (N_5266,N_5189,N_5142);
and U5267 (N_5267,N_5094,N_5136);
nor U5268 (N_5268,N_5092,N_5097);
or U5269 (N_5269,N_5033,N_5093);
and U5270 (N_5270,N_5074,N_5044);
xnor U5271 (N_5271,N_5242,N_5236);
nand U5272 (N_5272,N_5235,N_5015);
and U5273 (N_5273,N_5123,N_5096);
nor U5274 (N_5274,N_5146,N_5132);
nand U5275 (N_5275,N_5177,N_5206);
xnor U5276 (N_5276,N_5125,N_5241);
nor U5277 (N_5277,N_5119,N_5098);
or U5278 (N_5278,N_5192,N_5003);
nor U5279 (N_5279,N_5113,N_5026);
nand U5280 (N_5280,N_5227,N_5029);
and U5281 (N_5281,N_5209,N_5165);
xor U5282 (N_5282,N_5226,N_5060);
xnor U5283 (N_5283,N_5051,N_5089);
or U5284 (N_5284,N_5246,N_5191);
nand U5285 (N_5285,N_5012,N_5197);
nor U5286 (N_5286,N_5018,N_5084);
nor U5287 (N_5287,N_5087,N_5002);
xnor U5288 (N_5288,N_5168,N_5214);
nand U5289 (N_5289,N_5000,N_5190);
nand U5290 (N_5290,N_5128,N_5054);
xor U5291 (N_5291,N_5057,N_5179);
nand U5292 (N_5292,N_5010,N_5038);
nor U5293 (N_5293,N_5134,N_5114);
xor U5294 (N_5294,N_5173,N_5032);
nand U5295 (N_5295,N_5120,N_5187);
and U5296 (N_5296,N_5022,N_5046);
nand U5297 (N_5297,N_5172,N_5052);
nor U5298 (N_5298,N_5130,N_5140);
nand U5299 (N_5299,N_5182,N_5107);
nand U5300 (N_5300,N_5091,N_5081);
xnor U5301 (N_5301,N_5204,N_5078);
nor U5302 (N_5302,N_5216,N_5004);
and U5303 (N_5303,N_5058,N_5176);
nand U5304 (N_5304,N_5161,N_5080);
xor U5305 (N_5305,N_5230,N_5072);
and U5306 (N_5306,N_5215,N_5174);
nand U5307 (N_5307,N_5169,N_5064);
and U5308 (N_5308,N_5152,N_5184);
xor U5309 (N_5309,N_5131,N_5076);
xnor U5310 (N_5310,N_5239,N_5063);
and U5311 (N_5311,N_5100,N_5129);
nor U5312 (N_5312,N_5116,N_5070);
or U5313 (N_5313,N_5073,N_5150);
nor U5314 (N_5314,N_5090,N_5223);
xnor U5315 (N_5315,N_5041,N_5056);
or U5316 (N_5316,N_5147,N_5210);
and U5317 (N_5317,N_5071,N_5069);
and U5318 (N_5318,N_5103,N_5198);
xor U5319 (N_5319,N_5151,N_5105);
nor U5320 (N_5320,N_5224,N_5013);
nor U5321 (N_5321,N_5157,N_5021);
and U5322 (N_5322,N_5218,N_5171);
nand U5323 (N_5323,N_5050,N_5001);
or U5324 (N_5324,N_5111,N_5049);
and U5325 (N_5325,N_5014,N_5156);
and U5326 (N_5326,N_5108,N_5117);
nor U5327 (N_5327,N_5007,N_5248);
nor U5328 (N_5328,N_5042,N_5149);
nor U5329 (N_5329,N_5238,N_5212);
and U5330 (N_5330,N_5028,N_5203);
or U5331 (N_5331,N_5023,N_5036);
nand U5332 (N_5332,N_5155,N_5035);
xnor U5333 (N_5333,N_5083,N_5201);
nand U5334 (N_5334,N_5062,N_5016);
xnor U5335 (N_5335,N_5194,N_5232);
and U5336 (N_5336,N_5186,N_5148);
nand U5337 (N_5337,N_5075,N_5024);
xor U5338 (N_5338,N_5106,N_5027);
nand U5339 (N_5339,N_5217,N_5020);
and U5340 (N_5340,N_5086,N_5247);
or U5341 (N_5341,N_5077,N_5154);
nand U5342 (N_5342,N_5199,N_5202);
nor U5343 (N_5343,N_5164,N_5162);
or U5344 (N_5344,N_5183,N_5234);
nand U5345 (N_5345,N_5059,N_5017);
xor U5346 (N_5346,N_5110,N_5158);
and U5347 (N_5347,N_5139,N_5228);
xnor U5348 (N_5348,N_5160,N_5244);
and U5349 (N_5349,N_5221,N_5019);
xor U5350 (N_5350,N_5055,N_5067);
nand U5351 (N_5351,N_5122,N_5037);
nor U5352 (N_5352,N_5225,N_5200);
nor U5353 (N_5353,N_5233,N_5207);
xnor U5354 (N_5354,N_5043,N_5141);
nand U5355 (N_5355,N_5127,N_5045);
xor U5356 (N_5356,N_5188,N_5061);
or U5357 (N_5357,N_5249,N_5193);
nor U5358 (N_5358,N_5229,N_5237);
nor U5359 (N_5359,N_5163,N_5068);
nor U5360 (N_5360,N_5102,N_5133);
and U5361 (N_5361,N_5231,N_5118);
or U5362 (N_5362,N_5213,N_5222);
and U5363 (N_5363,N_5219,N_5159);
and U5364 (N_5364,N_5180,N_5138);
xor U5365 (N_5365,N_5124,N_5143);
and U5366 (N_5366,N_5034,N_5082);
nand U5367 (N_5367,N_5095,N_5135);
and U5368 (N_5368,N_5137,N_5112);
or U5369 (N_5369,N_5053,N_5066);
or U5370 (N_5370,N_5121,N_5079);
or U5371 (N_5371,N_5185,N_5048);
or U5372 (N_5372,N_5145,N_5205);
nor U5373 (N_5373,N_5047,N_5144);
or U5374 (N_5374,N_5006,N_5170);
nand U5375 (N_5375,N_5035,N_5158);
nand U5376 (N_5376,N_5164,N_5104);
nor U5377 (N_5377,N_5000,N_5186);
xor U5378 (N_5378,N_5091,N_5193);
nor U5379 (N_5379,N_5042,N_5082);
and U5380 (N_5380,N_5198,N_5174);
xnor U5381 (N_5381,N_5184,N_5070);
or U5382 (N_5382,N_5068,N_5148);
xnor U5383 (N_5383,N_5149,N_5188);
xnor U5384 (N_5384,N_5184,N_5202);
nor U5385 (N_5385,N_5195,N_5172);
nor U5386 (N_5386,N_5092,N_5039);
nand U5387 (N_5387,N_5199,N_5136);
and U5388 (N_5388,N_5004,N_5214);
nor U5389 (N_5389,N_5209,N_5189);
and U5390 (N_5390,N_5125,N_5212);
nor U5391 (N_5391,N_5009,N_5086);
nor U5392 (N_5392,N_5126,N_5097);
or U5393 (N_5393,N_5175,N_5133);
nor U5394 (N_5394,N_5134,N_5096);
and U5395 (N_5395,N_5017,N_5220);
nand U5396 (N_5396,N_5137,N_5237);
nand U5397 (N_5397,N_5161,N_5249);
nor U5398 (N_5398,N_5154,N_5196);
or U5399 (N_5399,N_5100,N_5052);
xnor U5400 (N_5400,N_5063,N_5032);
or U5401 (N_5401,N_5202,N_5221);
or U5402 (N_5402,N_5234,N_5088);
nand U5403 (N_5403,N_5024,N_5130);
nand U5404 (N_5404,N_5093,N_5062);
or U5405 (N_5405,N_5106,N_5001);
or U5406 (N_5406,N_5047,N_5068);
xnor U5407 (N_5407,N_5006,N_5051);
nand U5408 (N_5408,N_5077,N_5025);
xnor U5409 (N_5409,N_5248,N_5008);
xor U5410 (N_5410,N_5133,N_5024);
and U5411 (N_5411,N_5076,N_5214);
nor U5412 (N_5412,N_5033,N_5135);
nor U5413 (N_5413,N_5060,N_5014);
and U5414 (N_5414,N_5093,N_5139);
xnor U5415 (N_5415,N_5089,N_5224);
and U5416 (N_5416,N_5003,N_5218);
and U5417 (N_5417,N_5226,N_5231);
and U5418 (N_5418,N_5128,N_5151);
xnor U5419 (N_5419,N_5005,N_5055);
and U5420 (N_5420,N_5121,N_5205);
nor U5421 (N_5421,N_5106,N_5098);
nand U5422 (N_5422,N_5139,N_5229);
nand U5423 (N_5423,N_5211,N_5202);
and U5424 (N_5424,N_5019,N_5177);
nor U5425 (N_5425,N_5164,N_5180);
xor U5426 (N_5426,N_5065,N_5100);
and U5427 (N_5427,N_5184,N_5164);
nand U5428 (N_5428,N_5033,N_5036);
and U5429 (N_5429,N_5184,N_5046);
or U5430 (N_5430,N_5112,N_5114);
nand U5431 (N_5431,N_5127,N_5041);
xor U5432 (N_5432,N_5096,N_5219);
nor U5433 (N_5433,N_5197,N_5089);
xnor U5434 (N_5434,N_5203,N_5148);
xor U5435 (N_5435,N_5188,N_5090);
nand U5436 (N_5436,N_5189,N_5000);
xor U5437 (N_5437,N_5188,N_5233);
nor U5438 (N_5438,N_5145,N_5040);
or U5439 (N_5439,N_5244,N_5023);
nand U5440 (N_5440,N_5101,N_5022);
and U5441 (N_5441,N_5204,N_5146);
and U5442 (N_5442,N_5082,N_5166);
nor U5443 (N_5443,N_5068,N_5004);
or U5444 (N_5444,N_5142,N_5093);
and U5445 (N_5445,N_5201,N_5049);
xnor U5446 (N_5446,N_5177,N_5090);
xor U5447 (N_5447,N_5183,N_5076);
and U5448 (N_5448,N_5236,N_5029);
nor U5449 (N_5449,N_5028,N_5004);
nor U5450 (N_5450,N_5095,N_5147);
xor U5451 (N_5451,N_5049,N_5230);
or U5452 (N_5452,N_5135,N_5030);
nand U5453 (N_5453,N_5033,N_5004);
and U5454 (N_5454,N_5177,N_5009);
nand U5455 (N_5455,N_5050,N_5104);
xnor U5456 (N_5456,N_5223,N_5120);
nor U5457 (N_5457,N_5205,N_5029);
xnor U5458 (N_5458,N_5064,N_5029);
nor U5459 (N_5459,N_5118,N_5142);
nor U5460 (N_5460,N_5153,N_5206);
or U5461 (N_5461,N_5179,N_5215);
xor U5462 (N_5462,N_5089,N_5081);
nand U5463 (N_5463,N_5246,N_5192);
or U5464 (N_5464,N_5193,N_5200);
or U5465 (N_5465,N_5065,N_5021);
and U5466 (N_5466,N_5169,N_5241);
and U5467 (N_5467,N_5168,N_5050);
nand U5468 (N_5468,N_5100,N_5089);
nor U5469 (N_5469,N_5147,N_5186);
nor U5470 (N_5470,N_5159,N_5025);
or U5471 (N_5471,N_5092,N_5178);
nor U5472 (N_5472,N_5181,N_5159);
nand U5473 (N_5473,N_5178,N_5198);
or U5474 (N_5474,N_5221,N_5119);
nor U5475 (N_5475,N_5207,N_5069);
nand U5476 (N_5476,N_5155,N_5047);
or U5477 (N_5477,N_5009,N_5021);
xnor U5478 (N_5478,N_5229,N_5233);
xnor U5479 (N_5479,N_5157,N_5068);
nand U5480 (N_5480,N_5093,N_5048);
xnor U5481 (N_5481,N_5230,N_5008);
nor U5482 (N_5482,N_5053,N_5123);
nand U5483 (N_5483,N_5211,N_5061);
xnor U5484 (N_5484,N_5245,N_5087);
xnor U5485 (N_5485,N_5221,N_5215);
nor U5486 (N_5486,N_5108,N_5148);
xor U5487 (N_5487,N_5182,N_5230);
nor U5488 (N_5488,N_5024,N_5041);
xor U5489 (N_5489,N_5149,N_5228);
xor U5490 (N_5490,N_5249,N_5182);
or U5491 (N_5491,N_5084,N_5111);
nor U5492 (N_5492,N_5162,N_5097);
or U5493 (N_5493,N_5007,N_5104);
and U5494 (N_5494,N_5224,N_5216);
xnor U5495 (N_5495,N_5209,N_5013);
nand U5496 (N_5496,N_5026,N_5141);
nor U5497 (N_5497,N_5197,N_5061);
nor U5498 (N_5498,N_5246,N_5239);
and U5499 (N_5499,N_5098,N_5138);
nand U5500 (N_5500,N_5257,N_5372);
and U5501 (N_5501,N_5346,N_5355);
xor U5502 (N_5502,N_5480,N_5336);
nand U5503 (N_5503,N_5305,N_5411);
or U5504 (N_5504,N_5350,N_5253);
and U5505 (N_5505,N_5339,N_5412);
or U5506 (N_5506,N_5453,N_5394);
xor U5507 (N_5507,N_5369,N_5345);
and U5508 (N_5508,N_5448,N_5340);
and U5509 (N_5509,N_5373,N_5400);
nand U5510 (N_5510,N_5290,N_5364);
nand U5511 (N_5511,N_5441,N_5337);
or U5512 (N_5512,N_5396,N_5371);
or U5513 (N_5513,N_5408,N_5335);
and U5514 (N_5514,N_5344,N_5283);
or U5515 (N_5515,N_5387,N_5489);
nor U5516 (N_5516,N_5289,N_5367);
nor U5517 (N_5517,N_5347,N_5494);
nand U5518 (N_5518,N_5426,N_5269);
xnor U5519 (N_5519,N_5381,N_5483);
nand U5520 (N_5520,N_5296,N_5284);
nand U5521 (N_5521,N_5285,N_5474);
xnor U5522 (N_5522,N_5302,N_5498);
xnor U5523 (N_5523,N_5431,N_5481);
nand U5524 (N_5524,N_5273,N_5445);
and U5525 (N_5525,N_5332,N_5386);
nand U5526 (N_5526,N_5295,N_5321);
nand U5527 (N_5527,N_5465,N_5376);
nand U5528 (N_5528,N_5306,N_5260);
or U5529 (N_5529,N_5360,N_5298);
nor U5530 (N_5530,N_5262,N_5402);
and U5531 (N_5531,N_5365,N_5294);
or U5532 (N_5532,N_5276,N_5352);
xnor U5533 (N_5533,N_5375,N_5363);
and U5534 (N_5534,N_5384,N_5310);
and U5535 (N_5535,N_5354,N_5460);
or U5536 (N_5536,N_5251,N_5325);
or U5537 (N_5537,N_5459,N_5383);
nor U5538 (N_5538,N_5432,N_5359);
nor U5539 (N_5539,N_5319,N_5293);
xnor U5540 (N_5540,N_5472,N_5404);
nor U5541 (N_5541,N_5437,N_5439);
or U5542 (N_5542,N_5392,N_5438);
xnor U5543 (N_5543,N_5309,N_5315);
nor U5544 (N_5544,N_5461,N_5322);
xor U5545 (N_5545,N_5265,N_5254);
and U5546 (N_5546,N_5434,N_5385);
nor U5547 (N_5547,N_5452,N_5368);
or U5548 (N_5548,N_5499,N_5420);
and U5549 (N_5549,N_5343,N_5318);
nor U5550 (N_5550,N_5324,N_5418);
xor U5551 (N_5551,N_5333,N_5388);
or U5552 (N_5552,N_5399,N_5421);
nor U5553 (N_5553,N_5451,N_5429);
or U5554 (N_5554,N_5397,N_5446);
and U5555 (N_5555,N_5312,N_5485);
nand U5556 (N_5556,N_5304,N_5362);
and U5557 (N_5557,N_5424,N_5490);
and U5558 (N_5558,N_5301,N_5270);
and U5559 (N_5559,N_5281,N_5264);
nand U5560 (N_5560,N_5491,N_5455);
and U5561 (N_5561,N_5390,N_5405);
and U5562 (N_5562,N_5415,N_5370);
and U5563 (N_5563,N_5331,N_5486);
xnor U5564 (N_5564,N_5379,N_5443);
nor U5565 (N_5565,N_5280,N_5377);
nand U5566 (N_5566,N_5287,N_5450);
or U5567 (N_5567,N_5275,N_5313);
nor U5568 (N_5568,N_5442,N_5341);
nand U5569 (N_5569,N_5497,N_5391);
and U5570 (N_5570,N_5409,N_5378);
nand U5571 (N_5571,N_5393,N_5488);
xor U5572 (N_5572,N_5259,N_5338);
nand U5573 (N_5573,N_5475,N_5271);
nor U5574 (N_5574,N_5348,N_5410);
and U5575 (N_5575,N_5433,N_5492);
or U5576 (N_5576,N_5416,N_5493);
and U5577 (N_5577,N_5414,N_5496);
xor U5578 (N_5578,N_5417,N_5456);
and U5579 (N_5579,N_5374,N_5477);
and U5580 (N_5580,N_5467,N_5326);
or U5581 (N_5581,N_5428,N_5462);
and U5582 (N_5582,N_5278,N_5449);
or U5583 (N_5583,N_5267,N_5479);
and U5584 (N_5584,N_5252,N_5423);
or U5585 (N_5585,N_5291,N_5484);
nor U5586 (N_5586,N_5323,N_5464);
or U5587 (N_5587,N_5401,N_5470);
nand U5588 (N_5588,N_5473,N_5292);
nor U5589 (N_5589,N_5250,N_5430);
and U5590 (N_5590,N_5329,N_5299);
and U5591 (N_5591,N_5279,N_5261);
and U5592 (N_5592,N_5366,N_5288);
and U5593 (N_5593,N_5314,N_5334);
nor U5594 (N_5594,N_5286,N_5406);
nand U5595 (N_5595,N_5468,N_5300);
xnor U5596 (N_5596,N_5478,N_5357);
or U5597 (N_5597,N_5358,N_5349);
xnor U5598 (N_5598,N_5255,N_5495);
or U5599 (N_5599,N_5317,N_5297);
nand U5600 (N_5600,N_5311,N_5425);
or U5601 (N_5601,N_5458,N_5487);
nor U5602 (N_5602,N_5457,N_5389);
and U5603 (N_5603,N_5440,N_5469);
and U5604 (N_5604,N_5303,N_5454);
and U5605 (N_5605,N_5447,N_5422);
and U5606 (N_5606,N_5272,N_5380);
nor U5607 (N_5607,N_5256,N_5444);
nor U5608 (N_5608,N_5316,N_5463);
and U5609 (N_5609,N_5398,N_5328);
or U5610 (N_5610,N_5308,N_5436);
nand U5611 (N_5611,N_5351,N_5419);
and U5612 (N_5612,N_5353,N_5435);
nor U5613 (N_5613,N_5471,N_5356);
nand U5614 (N_5614,N_5413,N_5268);
nand U5615 (N_5615,N_5327,N_5427);
nand U5616 (N_5616,N_5307,N_5330);
nor U5617 (N_5617,N_5263,N_5342);
or U5618 (N_5618,N_5395,N_5361);
xor U5619 (N_5619,N_5403,N_5274);
nand U5620 (N_5620,N_5382,N_5320);
or U5621 (N_5621,N_5476,N_5282);
and U5622 (N_5622,N_5277,N_5266);
nor U5623 (N_5623,N_5466,N_5482);
and U5624 (N_5624,N_5258,N_5407);
nor U5625 (N_5625,N_5331,N_5284);
xnor U5626 (N_5626,N_5343,N_5424);
xnor U5627 (N_5627,N_5403,N_5284);
and U5628 (N_5628,N_5269,N_5335);
and U5629 (N_5629,N_5352,N_5444);
nand U5630 (N_5630,N_5334,N_5270);
and U5631 (N_5631,N_5278,N_5430);
nand U5632 (N_5632,N_5257,N_5428);
nand U5633 (N_5633,N_5427,N_5413);
xnor U5634 (N_5634,N_5439,N_5407);
or U5635 (N_5635,N_5280,N_5449);
nand U5636 (N_5636,N_5386,N_5366);
or U5637 (N_5637,N_5463,N_5396);
nand U5638 (N_5638,N_5358,N_5430);
or U5639 (N_5639,N_5446,N_5300);
and U5640 (N_5640,N_5336,N_5403);
nand U5641 (N_5641,N_5439,N_5280);
nor U5642 (N_5642,N_5377,N_5379);
nor U5643 (N_5643,N_5481,N_5470);
or U5644 (N_5644,N_5293,N_5380);
nand U5645 (N_5645,N_5481,N_5456);
nand U5646 (N_5646,N_5395,N_5370);
xnor U5647 (N_5647,N_5491,N_5475);
xor U5648 (N_5648,N_5494,N_5423);
and U5649 (N_5649,N_5348,N_5391);
or U5650 (N_5650,N_5473,N_5400);
nor U5651 (N_5651,N_5377,N_5370);
xnor U5652 (N_5652,N_5432,N_5413);
nor U5653 (N_5653,N_5280,N_5457);
nand U5654 (N_5654,N_5369,N_5486);
or U5655 (N_5655,N_5443,N_5415);
or U5656 (N_5656,N_5285,N_5497);
xor U5657 (N_5657,N_5464,N_5385);
nor U5658 (N_5658,N_5344,N_5377);
nor U5659 (N_5659,N_5343,N_5460);
and U5660 (N_5660,N_5398,N_5490);
and U5661 (N_5661,N_5358,N_5436);
xor U5662 (N_5662,N_5300,N_5334);
xor U5663 (N_5663,N_5313,N_5409);
nor U5664 (N_5664,N_5438,N_5303);
and U5665 (N_5665,N_5435,N_5316);
nor U5666 (N_5666,N_5290,N_5292);
nor U5667 (N_5667,N_5476,N_5386);
nor U5668 (N_5668,N_5282,N_5465);
xor U5669 (N_5669,N_5437,N_5314);
nor U5670 (N_5670,N_5270,N_5386);
nand U5671 (N_5671,N_5292,N_5443);
nor U5672 (N_5672,N_5269,N_5406);
nand U5673 (N_5673,N_5410,N_5321);
nor U5674 (N_5674,N_5451,N_5321);
nand U5675 (N_5675,N_5360,N_5449);
and U5676 (N_5676,N_5304,N_5403);
xor U5677 (N_5677,N_5319,N_5469);
or U5678 (N_5678,N_5454,N_5397);
or U5679 (N_5679,N_5475,N_5428);
and U5680 (N_5680,N_5341,N_5396);
and U5681 (N_5681,N_5414,N_5470);
and U5682 (N_5682,N_5495,N_5466);
nor U5683 (N_5683,N_5386,N_5321);
or U5684 (N_5684,N_5291,N_5415);
and U5685 (N_5685,N_5369,N_5336);
nor U5686 (N_5686,N_5293,N_5496);
and U5687 (N_5687,N_5486,N_5279);
or U5688 (N_5688,N_5309,N_5339);
or U5689 (N_5689,N_5457,N_5361);
xor U5690 (N_5690,N_5286,N_5301);
nor U5691 (N_5691,N_5302,N_5422);
and U5692 (N_5692,N_5383,N_5256);
and U5693 (N_5693,N_5377,N_5383);
nor U5694 (N_5694,N_5301,N_5448);
or U5695 (N_5695,N_5432,N_5456);
or U5696 (N_5696,N_5398,N_5367);
and U5697 (N_5697,N_5492,N_5363);
nor U5698 (N_5698,N_5466,N_5373);
nor U5699 (N_5699,N_5376,N_5272);
nor U5700 (N_5700,N_5477,N_5268);
nand U5701 (N_5701,N_5270,N_5426);
xor U5702 (N_5702,N_5469,N_5354);
and U5703 (N_5703,N_5336,N_5262);
and U5704 (N_5704,N_5463,N_5373);
nor U5705 (N_5705,N_5417,N_5473);
nor U5706 (N_5706,N_5455,N_5392);
nor U5707 (N_5707,N_5297,N_5379);
xnor U5708 (N_5708,N_5465,N_5299);
and U5709 (N_5709,N_5296,N_5466);
or U5710 (N_5710,N_5340,N_5311);
xor U5711 (N_5711,N_5481,N_5451);
or U5712 (N_5712,N_5459,N_5398);
nand U5713 (N_5713,N_5295,N_5438);
nor U5714 (N_5714,N_5416,N_5319);
or U5715 (N_5715,N_5404,N_5322);
and U5716 (N_5716,N_5313,N_5393);
nor U5717 (N_5717,N_5408,N_5281);
nor U5718 (N_5718,N_5462,N_5256);
xnor U5719 (N_5719,N_5438,N_5470);
and U5720 (N_5720,N_5410,N_5378);
and U5721 (N_5721,N_5438,N_5268);
nor U5722 (N_5722,N_5462,N_5339);
nor U5723 (N_5723,N_5446,N_5302);
and U5724 (N_5724,N_5280,N_5403);
and U5725 (N_5725,N_5320,N_5461);
nand U5726 (N_5726,N_5421,N_5337);
and U5727 (N_5727,N_5476,N_5277);
or U5728 (N_5728,N_5445,N_5305);
or U5729 (N_5729,N_5403,N_5424);
nor U5730 (N_5730,N_5387,N_5281);
nand U5731 (N_5731,N_5325,N_5416);
nand U5732 (N_5732,N_5388,N_5461);
nor U5733 (N_5733,N_5484,N_5296);
nand U5734 (N_5734,N_5371,N_5329);
or U5735 (N_5735,N_5324,N_5342);
nand U5736 (N_5736,N_5277,N_5479);
nor U5737 (N_5737,N_5360,N_5289);
nor U5738 (N_5738,N_5461,N_5352);
xor U5739 (N_5739,N_5440,N_5308);
xnor U5740 (N_5740,N_5350,N_5357);
nor U5741 (N_5741,N_5281,N_5391);
nand U5742 (N_5742,N_5476,N_5486);
and U5743 (N_5743,N_5429,N_5313);
xnor U5744 (N_5744,N_5324,N_5334);
and U5745 (N_5745,N_5419,N_5462);
xnor U5746 (N_5746,N_5293,N_5469);
nand U5747 (N_5747,N_5256,N_5461);
xnor U5748 (N_5748,N_5336,N_5283);
or U5749 (N_5749,N_5344,N_5276);
xor U5750 (N_5750,N_5553,N_5654);
and U5751 (N_5751,N_5714,N_5584);
nor U5752 (N_5752,N_5636,N_5623);
nor U5753 (N_5753,N_5561,N_5609);
nor U5754 (N_5754,N_5722,N_5541);
and U5755 (N_5755,N_5583,N_5677);
and U5756 (N_5756,N_5612,N_5659);
nand U5757 (N_5757,N_5709,N_5526);
xor U5758 (N_5758,N_5557,N_5720);
or U5759 (N_5759,N_5540,N_5738);
xnor U5760 (N_5760,N_5749,N_5593);
and U5761 (N_5761,N_5743,N_5529);
nor U5762 (N_5762,N_5608,N_5517);
nand U5763 (N_5763,N_5666,N_5597);
or U5764 (N_5764,N_5549,N_5668);
or U5765 (N_5765,N_5680,N_5711);
or U5766 (N_5766,N_5552,N_5548);
nand U5767 (N_5767,N_5658,N_5707);
xnor U5768 (N_5768,N_5520,N_5513);
nand U5769 (N_5769,N_5535,N_5632);
xor U5770 (N_5770,N_5664,N_5576);
xnor U5771 (N_5771,N_5509,N_5566);
or U5772 (N_5772,N_5531,N_5629);
nand U5773 (N_5773,N_5705,N_5578);
nand U5774 (N_5774,N_5621,N_5594);
nor U5775 (N_5775,N_5596,N_5639);
xor U5776 (N_5776,N_5657,N_5665);
and U5777 (N_5777,N_5739,N_5554);
or U5778 (N_5778,N_5510,N_5701);
nor U5779 (N_5779,N_5533,N_5546);
nor U5780 (N_5780,N_5717,N_5511);
xnor U5781 (N_5781,N_5706,N_5688);
nand U5782 (N_5782,N_5579,N_5573);
nand U5783 (N_5783,N_5687,N_5699);
or U5784 (N_5784,N_5678,N_5581);
nor U5785 (N_5785,N_5641,N_5515);
or U5786 (N_5786,N_5560,N_5598);
nand U5787 (N_5787,N_5732,N_5518);
or U5788 (N_5788,N_5704,N_5726);
xor U5789 (N_5789,N_5656,N_5590);
nand U5790 (N_5790,N_5735,N_5730);
nor U5791 (N_5791,N_5672,N_5556);
nor U5792 (N_5792,N_5624,N_5626);
xor U5793 (N_5793,N_5559,N_5525);
xnor U5794 (N_5794,N_5622,N_5569);
nor U5795 (N_5795,N_5547,N_5615);
nor U5796 (N_5796,N_5521,N_5502);
or U5797 (N_5797,N_5697,N_5507);
xor U5798 (N_5798,N_5602,N_5628);
xor U5799 (N_5799,N_5631,N_5729);
and U5800 (N_5800,N_5550,N_5564);
nor U5801 (N_5801,N_5512,N_5610);
nand U5802 (N_5802,N_5508,N_5582);
nor U5803 (N_5803,N_5585,N_5587);
nand U5804 (N_5804,N_5731,N_5601);
and U5805 (N_5805,N_5663,N_5644);
and U5806 (N_5806,N_5645,N_5696);
and U5807 (N_5807,N_5646,N_5683);
and U5808 (N_5808,N_5613,N_5647);
or U5809 (N_5809,N_5700,N_5712);
nand U5810 (N_5810,N_5660,N_5643);
nor U5811 (N_5811,N_5505,N_5567);
and U5812 (N_5812,N_5742,N_5538);
nor U5813 (N_5813,N_5504,N_5648);
nand U5814 (N_5814,N_5682,N_5542);
xnor U5815 (N_5815,N_5721,N_5630);
nand U5816 (N_5816,N_5516,N_5501);
nor U5817 (N_5817,N_5570,N_5661);
and U5818 (N_5818,N_5519,N_5650);
xnor U5819 (N_5819,N_5703,N_5649);
nor U5820 (N_5820,N_5702,N_5617);
xnor U5821 (N_5821,N_5745,N_5637);
or U5822 (N_5822,N_5670,N_5572);
and U5823 (N_5823,N_5611,N_5551);
or U5824 (N_5824,N_5577,N_5747);
or U5825 (N_5825,N_5689,N_5595);
nand U5826 (N_5826,N_5600,N_5651);
nor U5827 (N_5827,N_5693,N_5638);
and U5828 (N_5828,N_5692,N_5627);
xnor U5829 (N_5829,N_5633,N_5724);
and U5830 (N_5830,N_5662,N_5652);
and U5831 (N_5831,N_5674,N_5728);
and U5832 (N_5832,N_5591,N_5718);
xnor U5833 (N_5833,N_5695,N_5606);
xnor U5834 (N_5834,N_5691,N_5574);
or U5835 (N_5835,N_5723,N_5620);
xor U5836 (N_5836,N_5737,N_5716);
or U5837 (N_5837,N_5733,N_5690);
and U5838 (N_5838,N_5736,N_5686);
and U5839 (N_5839,N_5575,N_5530);
or U5840 (N_5840,N_5684,N_5618);
xor U5841 (N_5841,N_5603,N_5614);
nand U5842 (N_5842,N_5588,N_5543);
xnor U5843 (N_5843,N_5744,N_5673);
and U5844 (N_5844,N_5698,N_5642);
and U5845 (N_5845,N_5746,N_5679);
or U5846 (N_5846,N_5605,N_5741);
or U5847 (N_5847,N_5580,N_5734);
nand U5848 (N_5848,N_5681,N_5685);
xor U5849 (N_5849,N_5635,N_5710);
nand U5850 (N_5850,N_5563,N_5545);
and U5851 (N_5851,N_5671,N_5655);
or U5852 (N_5852,N_5669,N_5586);
or U5853 (N_5853,N_5562,N_5740);
or U5854 (N_5854,N_5544,N_5719);
nor U5855 (N_5855,N_5667,N_5558);
nand U5856 (N_5856,N_5571,N_5537);
and U5857 (N_5857,N_5607,N_5708);
nand U5858 (N_5858,N_5713,N_5675);
nand U5859 (N_5859,N_5527,N_5536);
and U5860 (N_5860,N_5555,N_5532);
nand U5861 (N_5861,N_5725,N_5539);
nor U5862 (N_5862,N_5653,N_5534);
and U5863 (N_5863,N_5589,N_5528);
nand U5864 (N_5864,N_5599,N_5676);
and U5865 (N_5865,N_5715,N_5503);
nand U5866 (N_5866,N_5506,N_5568);
xor U5867 (N_5867,N_5524,N_5616);
nor U5868 (N_5868,N_5592,N_5619);
xnor U5869 (N_5869,N_5514,N_5748);
or U5870 (N_5870,N_5640,N_5694);
or U5871 (N_5871,N_5604,N_5634);
and U5872 (N_5872,N_5625,N_5522);
xnor U5873 (N_5873,N_5727,N_5523);
or U5874 (N_5874,N_5500,N_5565);
or U5875 (N_5875,N_5500,N_5562);
or U5876 (N_5876,N_5699,N_5735);
and U5877 (N_5877,N_5659,N_5624);
nand U5878 (N_5878,N_5611,N_5664);
nand U5879 (N_5879,N_5653,N_5624);
and U5880 (N_5880,N_5562,N_5648);
xnor U5881 (N_5881,N_5641,N_5533);
nor U5882 (N_5882,N_5549,N_5675);
nor U5883 (N_5883,N_5545,N_5530);
xnor U5884 (N_5884,N_5586,N_5747);
xor U5885 (N_5885,N_5683,N_5735);
xor U5886 (N_5886,N_5707,N_5657);
or U5887 (N_5887,N_5741,N_5583);
nand U5888 (N_5888,N_5611,N_5577);
and U5889 (N_5889,N_5504,N_5600);
nand U5890 (N_5890,N_5717,N_5586);
nand U5891 (N_5891,N_5630,N_5704);
nor U5892 (N_5892,N_5551,N_5712);
nor U5893 (N_5893,N_5532,N_5592);
nand U5894 (N_5894,N_5666,N_5547);
or U5895 (N_5895,N_5566,N_5651);
nor U5896 (N_5896,N_5583,N_5693);
nand U5897 (N_5897,N_5654,N_5608);
nor U5898 (N_5898,N_5506,N_5528);
nand U5899 (N_5899,N_5683,N_5502);
xnor U5900 (N_5900,N_5528,N_5693);
nand U5901 (N_5901,N_5714,N_5620);
nor U5902 (N_5902,N_5613,N_5678);
nor U5903 (N_5903,N_5570,N_5516);
nor U5904 (N_5904,N_5741,N_5658);
or U5905 (N_5905,N_5679,N_5537);
nand U5906 (N_5906,N_5662,N_5663);
or U5907 (N_5907,N_5515,N_5520);
and U5908 (N_5908,N_5547,N_5706);
xnor U5909 (N_5909,N_5738,N_5702);
or U5910 (N_5910,N_5655,N_5516);
or U5911 (N_5911,N_5693,N_5644);
xnor U5912 (N_5912,N_5673,N_5507);
nand U5913 (N_5913,N_5701,N_5598);
or U5914 (N_5914,N_5583,N_5680);
nand U5915 (N_5915,N_5703,N_5736);
xor U5916 (N_5916,N_5526,N_5698);
nand U5917 (N_5917,N_5514,N_5668);
and U5918 (N_5918,N_5718,N_5581);
or U5919 (N_5919,N_5718,N_5730);
nand U5920 (N_5920,N_5681,N_5748);
or U5921 (N_5921,N_5608,N_5748);
xor U5922 (N_5922,N_5748,N_5560);
xor U5923 (N_5923,N_5509,N_5713);
nor U5924 (N_5924,N_5541,N_5555);
or U5925 (N_5925,N_5554,N_5508);
nand U5926 (N_5926,N_5681,N_5552);
nand U5927 (N_5927,N_5505,N_5570);
and U5928 (N_5928,N_5723,N_5644);
xor U5929 (N_5929,N_5697,N_5529);
and U5930 (N_5930,N_5672,N_5514);
nand U5931 (N_5931,N_5548,N_5722);
xnor U5932 (N_5932,N_5644,N_5555);
nor U5933 (N_5933,N_5532,N_5627);
xor U5934 (N_5934,N_5526,N_5667);
nor U5935 (N_5935,N_5549,N_5671);
xnor U5936 (N_5936,N_5658,N_5576);
or U5937 (N_5937,N_5739,N_5571);
nor U5938 (N_5938,N_5545,N_5696);
or U5939 (N_5939,N_5666,N_5653);
and U5940 (N_5940,N_5593,N_5581);
or U5941 (N_5941,N_5660,N_5672);
or U5942 (N_5942,N_5656,N_5531);
nand U5943 (N_5943,N_5587,N_5609);
or U5944 (N_5944,N_5702,N_5696);
nand U5945 (N_5945,N_5612,N_5609);
nor U5946 (N_5946,N_5652,N_5539);
xnor U5947 (N_5947,N_5520,N_5569);
nand U5948 (N_5948,N_5721,N_5644);
nor U5949 (N_5949,N_5737,N_5508);
or U5950 (N_5950,N_5685,N_5643);
nor U5951 (N_5951,N_5576,N_5604);
or U5952 (N_5952,N_5740,N_5726);
nor U5953 (N_5953,N_5555,N_5698);
nor U5954 (N_5954,N_5671,N_5566);
nand U5955 (N_5955,N_5624,N_5727);
or U5956 (N_5956,N_5743,N_5694);
xor U5957 (N_5957,N_5744,N_5708);
nand U5958 (N_5958,N_5504,N_5739);
nand U5959 (N_5959,N_5635,N_5724);
nand U5960 (N_5960,N_5733,N_5593);
and U5961 (N_5961,N_5595,N_5591);
nand U5962 (N_5962,N_5653,N_5734);
nor U5963 (N_5963,N_5619,N_5578);
or U5964 (N_5964,N_5606,N_5566);
nor U5965 (N_5965,N_5543,N_5642);
nand U5966 (N_5966,N_5679,N_5698);
nor U5967 (N_5967,N_5684,N_5569);
nand U5968 (N_5968,N_5725,N_5714);
nor U5969 (N_5969,N_5636,N_5573);
nand U5970 (N_5970,N_5560,N_5719);
and U5971 (N_5971,N_5502,N_5542);
and U5972 (N_5972,N_5623,N_5614);
nand U5973 (N_5973,N_5506,N_5727);
and U5974 (N_5974,N_5640,N_5638);
nand U5975 (N_5975,N_5578,N_5618);
nor U5976 (N_5976,N_5565,N_5724);
and U5977 (N_5977,N_5744,N_5514);
nand U5978 (N_5978,N_5582,N_5513);
nand U5979 (N_5979,N_5563,N_5655);
or U5980 (N_5980,N_5652,N_5607);
or U5981 (N_5981,N_5503,N_5720);
or U5982 (N_5982,N_5583,N_5625);
nand U5983 (N_5983,N_5726,N_5552);
nand U5984 (N_5984,N_5698,N_5747);
or U5985 (N_5985,N_5666,N_5556);
xor U5986 (N_5986,N_5587,N_5693);
or U5987 (N_5987,N_5674,N_5725);
nor U5988 (N_5988,N_5719,N_5606);
or U5989 (N_5989,N_5660,N_5697);
nand U5990 (N_5990,N_5510,N_5636);
or U5991 (N_5991,N_5546,N_5742);
or U5992 (N_5992,N_5566,N_5543);
nor U5993 (N_5993,N_5707,N_5701);
xnor U5994 (N_5994,N_5729,N_5597);
and U5995 (N_5995,N_5646,N_5520);
nand U5996 (N_5996,N_5511,N_5652);
nand U5997 (N_5997,N_5577,N_5567);
or U5998 (N_5998,N_5528,N_5557);
or U5999 (N_5999,N_5553,N_5610);
or U6000 (N_6000,N_5944,N_5814);
xnor U6001 (N_6001,N_5996,N_5908);
nand U6002 (N_6002,N_5955,N_5932);
and U6003 (N_6003,N_5892,N_5920);
and U6004 (N_6004,N_5906,N_5937);
xnor U6005 (N_6005,N_5898,N_5921);
and U6006 (N_6006,N_5785,N_5816);
and U6007 (N_6007,N_5951,N_5979);
or U6008 (N_6008,N_5813,N_5991);
xnor U6009 (N_6009,N_5970,N_5826);
xnor U6010 (N_6010,N_5965,N_5988);
or U6011 (N_6011,N_5787,N_5771);
nand U6012 (N_6012,N_5842,N_5790);
or U6013 (N_6013,N_5775,N_5989);
or U6014 (N_6014,N_5935,N_5960);
or U6015 (N_6015,N_5945,N_5860);
xnor U6016 (N_6016,N_5885,N_5774);
xor U6017 (N_6017,N_5818,N_5819);
nor U6018 (N_6018,N_5983,N_5871);
nand U6019 (N_6019,N_5994,N_5980);
and U6020 (N_6020,N_5773,N_5999);
nand U6021 (N_6021,N_5878,N_5838);
nor U6022 (N_6022,N_5803,N_5897);
or U6023 (N_6023,N_5886,N_5879);
or U6024 (N_6024,N_5820,N_5966);
xnor U6025 (N_6025,N_5788,N_5830);
nor U6026 (N_6026,N_5863,N_5836);
or U6027 (N_6027,N_5903,N_5754);
nor U6028 (N_6028,N_5811,N_5828);
xor U6029 (N_6029,N_5783,N_5896);
or U6030 (N_6030,N_5971,N_5781);
and U6031 (N_6031,N_5969,N_5794);
nor U6032 (N_6032,N_5807,N_5913);
nor U6033 (N_6033,N_5793,N_5823);
or U6034 (N_6034,N_5856,N_5796);
and U6035 (N_6035,N_5938,N_5802);
or U6036 (N_6036,N_5873,N_5780);
nor U6037 (N_6037,N_5880,N_5952);
or U6038 (N_6038,N_5976,N_5911);
or U6039 (N_6039,N_5868,N_5872);
nor U6040 (N_6040,N_5844,N_5766);
and U6041 (N_6041,N_5964,N_5767);
nand U6042 (N_6042,N_5930,N_5992);
xnor U6043 (N_6043,N_5909,N_5875);
or U6044 (N_6044,N_5910,N_5997);
and U6045 (N_6045,N_5890,N_5751);
xor U6046 (N_6046,N_5756,N_5870);
and U6047 (N_6047,N_5953,N_5975);
xor U6048 (N_6048,N_5853,N_5889);
or U6049 (N_6049,N_5993,N_5835);
and U6050 (N_6050,N_5825,N_5987);
or U6051 (N_6051,N_5949,N_5998);
nand U6052 (N_6052,N_5939,N_5928);
nor U6053 (N_6053,N_5797,N_5974);
xnor U6054 (N_6054,N_5934,N_5902);
nand U6055 (N_6055,N_5808,N_5851);
nand U6056 (N_6056,N_5795,N_5900);
xnor U6057 (N_6057,N_5809,N_5887);
and U6058 (N_6058,N_5805,N_5968);
xor U6059 (N_6059,N_5986,N_5990);
and U6060 (N_6060,N_5926,N_5824);
xor U6061 (N_6061,N_5789,N_5772);
nand U6062 (N_6062,N_5854,N_5958);
and U6063 (N_6063,N_5876,N_5954);
xor U6064 (N_6064,N_5855,N_5973);
nand U6065 (N_6065,N_5786,N_5753);
nor U6066 (N_6066,N_5962,N_5961);
nor U6067 (N_6067,N_5815,N_5822);
xnor U6068 (N_6068,N_5915,N_5927);
and U6069 (N_6069,N_5812,N_5864);
nand U6070 (N_6070,N_5821,N_5959);
xnor U6071 (N_6071,N_5929,N_5752);
or U6072 (N_6072,N_5925,N_5760);
nor U6073 (N_6073,N_5852,N_5877);
nor U6074 (N_6074,N_5833,N_5948);
or U6075 (N_6075,N_5750,N_5799);
xor U6076 (N_6076,N_5763,N_5779);
nand U6077 (N_6077,N_5778,N_5762);
nand U6078 (N_6078,N_5755,N_5904);
or U6079 (N_6079,N_5784,N_5943);
nor U6080 (N_6080,N_5978,N_5977);
and U6081 (N_6081,N_5941,N_5905);
nor U6082 (N_6082,N_5982,N_5770);
or U6083 (N_6083,N_5942,N_5845);
nand U6084 (N_6084,N_5883,N_5895);
xnor U6085 (N_6085,N_5946,N_5882);
xnor U6086 (N_6086,N_5804,N_5867);
and U6087 (N_6087,N_5924,N_5843);
or U6088 (N_6088,N_5884,N_5901);
xor U6089 (N_6089,N_5765,N_5893);
nand U6090 (N_6090,N_5931,N_5847);
xnor U6091 (N_6091,N_5891,N_5899);
xor U6092 (N_6092,N_5792,N_5933);
xnor U6093 (N_6093,N_5874,N_5858);
nor U6094 (N_6094,N_5840,N_5777);
xor U6095 (N_6095,N_5850,N_5846);
or U6096 (N_6096,N_5985,N_5940);
xor U6097 (N_6097,N_5914,N_5848);
xnor U6098 (N_6098,N_5957,N_5866);
and U6099 (N_6099,N_5817,N_5806);
and U6100 (N_6100,N_5984,N_5841);
xnor U6101 (N_6101,N_5801,N_5936);
and U6102 (N_6102,N_5919,N_5758);
or U6103 (N_6103,N_5759,N_5950);
xnor U6104 (N_6104,N_5837,N_5917);
nor U6105 (N_6105,N_5869,N_5947);
nand U6106 (N_6106,N_5861,N_5888);
xnor U6107 (N_6107,N_5862,N_5981);
and U6108 (N_6108,N_5839,N_5881);
nand U6109 (N_6109,N_5972,N_5857);
xnor U6110 (N_6110,N_5956,N_5834);
and U6111 (N_6111,N_5918,N_5916);
and U6112 (N_6112,N_5963,N_5912);
or U6113 (N_6113,N_5782,N_5810);
and U6114 (N_6114,N_5894,N_5967);
xor U6115 (N_6115,N_5769,N_5791);
or U6116 (N_6116,N_5798,N_5829);
xnor U6117 (N_6117,N_5800,N_5923);
nand U6118 (N_6118,N_5832,N_5827);
or U6119 (N_6119,N_5764,N_5859);
or U6120 (N_6120,N_5907,N_5849);
nand U6121 (N_6121,N_5776,N_5768);
xnor U6122 (N_6122,N_5761,N_5922);
xnor U6123 (N_6123,N_5831,N_5865);
or U6124 (N_6124,N_5995,N_5757);
nand U6125 (N_6125,N_5787,N_5968);
nor U6126 (N_6126,N_5893,N_5777);
xor U6127 (N_6127,N_5826,N_5803);
and U6128 (N_6128,N_5757,N_5941);
nor U6129 (N_6129,N_5861,N_5941);
xnor U6130 (N_6130,N_5805,N_5770);
and U6131 (N_6131,N_5750,N_5930);
xnor U6132 (N_6132,N_5805,N_5902);
or U6133 (N_6133,N_5905,N_5879);
nor U6134 (N_6134,N_5837,N_5865);
nor U6135 (N_6135,N_5764,N_5865);
and U6136 (N_6136,N_5953,N_5750);
xor U6137 (N_6137,N_5811,N_5847);
xnor U6138 (N_6138,N_5805,N_5795);
nand U6139 (N_6139,N_5829,N_5993);
and U6140 (N_6140,N_5759,N_5991);
xnor U6141 (N_6141,N_5852,N_5805);
and U6142 (N_6142,N_5910,N_5818);
or U6143 (N_6143,N_5977,N_5765);
nand U6144 (N_6144,N_5797,N_5817);
xnor U6145 (N_6145,N_5874,N_5844);
and U6146 (N_6146,N_5786,N_5779);
xnor U6147 (N_6147,N_5998,N_5866);
xor U6148 (N_6148,N_5887,N_5814);
or U6149 (N_6149,N_5986,N_5970);
or U6150 (N_6150,N_5775,N_5988);
and U6151 (N_6151,N_5817,N_5825);
nor U6152 (N_6152,N_5953,N_5881);
xor U6153 (N_6153,N_5779,N_5953);
nor U6154 (N_6154,N_5757,N_5902);
and U6155 (N_6155,N_5766,N_5930);
nor U6156 (N_6156,N_5993,N_5798);
or U6157 (N_6157,N_5968,N_5800);
nand U6158 (N_6158,N_5757,N_5983);
nand U6159 (N_6159,N_5949,N_5807);
nor U6160 (N_6160,N_5915,N_5758);
nor U6161 (N_6161,N_5998,N_5971);
and U6162 (N_6162,N_5976,N_5868);
nor U6163 (N_6163,N_5997,N_5832);
xor U6164 (N_6164,N_5905,N_5792);
and U6165 (N_6165,N_5946,N_5957);
or U6166 (N_6166,N_5761,N_5814);
and U6167 (N_6167,N_5871,N_5773);
and U6168 (N_6168,N_5787,N_5961);
nand U6169 (N_6169,N_5788,N_5751);
nor U6170 (N_6170,N_5955,N_5891);
or U6171 (N_6171,N_5995,N_5842);
nand U6172 (N_6172,N_5948,N_5853);
nor U6173 (N_6173,N_5976,N_5964);
and U6174 (N_6174,N_5869,N_5770);
and U6175 (N_6175,N_5966,N_5789);
xor U6176 (N_6176,N_5957,N_5883);
nand U6177 (N_6177,N_5838,N_5961);
or U6178 (N_6178,N_5889,N_5787);
and U6179 (N_6179,N_5884,N_5978);
or U6180 (N_6180,N_5943,N_5979);
nand U6181 (N_6181,N_5973,N_5968);
xnor U6182 (N_6182,N_5761,N_5965);
xnor U6183 (N_6183,N_5861,N_5979);
nor U6184 (N_6184,N_5858,N_5928);
nor U6185 (N_6185,N_5815,N_5769);
xnor U6186 (N_6186,N_5917,N_5785);
nand U6187 (N_6187,N_5924,N_5910);
xor U6188 (N_6188,N_5913,N_5763);
nor U6189 (N_6189,N_5833,N_5932);
nor U6190 (N_6190,N_5914,N_5826);
nor U6191 (N_6191,N_5758,N_5844);
nor U6192 (N_6192,N_5993,N_5815);
nand U6193 (N_6193,N_5980,N_5836);
or U6194 (N_6194,N_5991,N_5878);
xnor U6195 (N_6195,N_5803,N_5900);
xor U6196 (N_6196,N_5943,N_5905);
xnor U6197 (N_6197,N_5908,N_5823);
nor U6198 (N_6198,N_5975,N_5905);
xnor U6199 (N_6199,N_5895,N_5885);
and U6200 (N_6200,N_5969,N_5964);
nor U6201 (N_6201,N_5758,N_5864);
xnor U6202 (N_6202,N_5990,N_5936);
and U6203 (N_6203,N_5881,N_5906);
xnor U6204 (N_6204,N_5869,N_5750);
and U6205 (N_6205,N_5974,N_5871);
and U6206 (N_6206,N_5764,N_5958);
nor U6207 (N_6207,N_5782,N_5944);
and U6208 (N_6208,N_5892,N_5882);
and U6209 (N_6209,N_5898,N_5900);
xor U6210 (N_6210,N_5780,N_5920);
nor U6211 (N_6211,N_5855,N_5840);
nand U6212 (N_6212,N_5857,N_5902);
or U6213 (N_6213,N_5964,N_5912);
nor U6214 (N_6214,N_5899,N_5855);
nor U6215 (N_6215,N_5881,N_5860);
and U6216 (N_6216,N_5939,N_5894);
xnor U6217 (N_6217,N_5935,N_5848);
or U6218 (N_6218,N_5817,N_5804);
nand U6219 (N_6219,N_5946,N_5779);
nor U6220 (N_6220,N_5844,N_5985);
nor U6221 (N_6221,N_5798,N_5902);
and U6222 (N_6222,N_5924,N_5802);
or U6223 (N_6223,N_5820,N_5867);
nor U6224 (N_6224,N_5877,N_5779);
nor U6225 (N_6225,N_5804,N_5989);
nand U6226 (N_6226,N_5963,N_5871);
nand U6227 (N_6227,N_5835,N_5760);
or U6228 (N_6228,N_5761,N_5986);
and U6229 (N_6229,N_5867,N_5959);
and U6230 (N_6230,N_5957,N_5848);
or U6231 (N_6231,N_5761,N_5797);
or U6232 (N_6232,N_5963,N_5820);
xor U6233 (N_6233,N_5783,N_5963);
nor U6234 (N_6234,N_5806,N_5801);
nand U6235 (N_6235,N_5809,N_5802);
xnor U6236 (N_6236,N_5914,N_5915);
xor U6237 (N_6237,N_5931,N_5937);
nand U6238 (N_6238,N_5872,N_5936);
and U6239 (N_6239,N_5843,N_5921);
nor U6240 (N_6240,N_5754,N_5927);
xor U6241 (N_6241,N_5845,N_5844);
and U6242 (N_6242,N_5782,N_5989);
or U6243 (N_6243,N_5849,N_5908);
nand U6244 (N_6244,N_5974,N_5875);
and U6245 (N_6245,N_5927,N_5987);
nand U6246 (N_6246,N_5900,N_5973);
xnor U6247 (N_6247,N_5905,N_5771);
and U6248 (N_6248,N_5832,N_5812);
and U6249 (N_6249,N_5915,N_5770);
nor U6250 (N_6250,N_6013,N_6163);
and U6251 (N_6251,N_6158,N_6128);
and U6252 (N_6252,N_6023,N_6177);
nand U6253 (N_6253,N_6109,N_6115);
xnor U6254 (N_6254,N_6239,N_6077);
nand U6255 (N_6255,N_6041,N_6153);
nand U6256 (N_6256,N_6096,N_6181);
and U6257 (N_6257,N_6069,N_6139);
or U6258 (N_6258,N_6084,N_6032);
or U6259 (N_6259,N_6097,N_6076);
and U6260 (N_6260,N_6233,N_6024);
and U6261 (N_6261,N_6112,N_6147);
nand U6262 (N_6262,N_6218,N_6092);
xnor U6263 (N_6263,N_6230,N_6043);
and U6264 (N_6264,N_6053,N_6197);
nand U6265 (N_6265,N_6065,N_6160);
xor U6266 (N_6266,N_6019,N_6120);
nor U6267 (N_6267,N_6007,N_6143);
xnor U6268 (N_6268,N_6093,N_6075);
xnor U6269 (N_6269,N_6101,N_6078);
and U6270 (N_6270,N_6190,N_6243);
and U6271 (N_6271,N_6142,N_6150);
xor U6272 (N_6272,N_6200,N_6237);
xor U6273 (N_6273,N_6136,N_6049);
nor U6274 (N_6274,N_6231,N_6079);
nand U6275 (N_6275,N_6073,N_6240);
xor U6276 (N_6276,N_6246,N_6220);
or U6277 (N_6277,N_6195,N_6014);
xor U6278 (N_6278,N_6038,N_6131);
nand U6279 (N_6279,N_6011,N_6026);
and U6280 (N_6280,N_6009,N_6247);
nor U6281 (N_6281,N_6234,N_6207);
nor U6282 (N_6282,N_6060,N_6185);
or U6283 (N_6283,N_6006,N_6151);
nand U6284 (N_6284,N_6114,N_6189);
nand U6285 (N_6285,N_6104,N_6054);
nor U6286 (N_6286,N_6125,N_6161);
nand U6287 (N_6287,N_6057,N_6241);
or U6288 (N_6288,N_6022,N_6118);
nand U6289 (N_6289,N_6148,N_6003);
nor U6290 (N_6290,N_6004,N_6074);
nor U6291 (N_6291,N_6132,N_6196);
nand U6292 (N_6292,N_6040,N_6106);
xor U6293 (N_6293,N_6113,N_6156);
or U6294 (N_6294,N_6063,N_6146);
nand U6295 (N_6295,N_6215,N_6082);
nor U6296 (N_6296,N_6030,N_6085);
nor U6297 (N_6297,N_6179,N_6225);
and U6298 (N_6298,N_6155,N_6058);
and U6299 (N_6299,N_6107,N_6224);
or U6300 (N_6300,N_6238,N_6042);
nor U6301 (N_6301,N_6081,N_6140);
xor U6302 (N_6302,N_6211,N_6090);
or U6303 (N_6303,N_6050,N_6087);
nand U6304 (N_6304,N_6100,N_6175);
nand U6305 (N_6305,N_6046,N_6229);
nor U6306 (N_6306,N_6135,N_6212);
nand U6307 (N_6307,N_6020,N_6236);
nor U6308 (N_6308,N_6203,N_6213);
xor U6309 (N_6309,N_6137,N_6249);
nor U6310 (N_6310,N_6176,N_6064);
nor U6311 (N_6311,N_6138,N_6037);
or U6312 (N_6312,N_6016,N_6015);
nand U6313 (N_6313,N_6048,N_6021);
and U6314 (N_6314,N_6012,N_6192);
nor U6315 (N_6315,N_6094,N_6091);
or U6316 (N_6316,N_6103,N_6198);
nor U6317 (N_6317,N_6129,N_6070);
and U6318 (N_6318,N_6056,N_6206);
nand U6319 (N_6319,N_6072,N_6000);
xor U6320 (N_6320,N_6183,N_6108);
nor U6321 (N_6321,N_6242,N_6086);
nor U6322 (N_6322,N_6111,N_6174);
xnor U6323 (N_6323,N_6002,N_6025);
or U6324 (N_6324,N_6235,N_6204);
xnor U6325 (N_6325,N_6039,N_6133);
nand U6326 (N_6326,N_6221,N_6099);
xnor U6327 (N_6327,N_6008,N_6062);
nor U6328 (N_6328,N_6191,N_6232);
nand U6329 (N_6329,N_6029,N_6066);
nand U6330 (N_6330,N_6244,N_6164);
nor U6331 (N_6331,N_6214,N_6216);
or U6332 (N_6332,N_6187,N_6144);
or U6333 (N_6333,N_6119,N_6031);
nor U6334 (N_6334,N_6035,N_6171);
nand U6335 (N_6335,N_6223,N_6027);
nor U6336 (N_6336,N_6051,N_6167);
xnor U6337 (N_6337,N_6245,N_6061);
nand U6338 (N_6338,N_6149,N_6033);
or U6339 (N_6339,N_6170,N_6123);
and U6340 (N_6340,N_6172,N_6166);
nor U6341 (N_6341,N_6184,N_6157);
nand U6342 (N_6342,N_6124,N_6210);
xnor U6343 (N_6343,N_6067,N_6152);
nand U6344 (N_6344,N_6001,N_6199);
xnor U6345 (N_6345,N_6162,N_6052);
and U6346 (N_6346,N_6127,N_6018);
xor U6347 (N_6347,N_6068,N_6194);
nand U6348 (N_6348,N_6209,N_6028);
xor U6349 (N_6349,N_6182,N_6010);
and U6350 (N_6350,N_6005,N_6110);
and U6351 (N_6351,N_6227,N_6219);
nand U6352 (N_6352,N_6188,N_6248);
nand U6353 (N_6353,N_6202,N_6205);
or U6354 (N_6354,N_6071,N_6034);
nor U6355 (N_6355,N_6165,N_6095);
or U6356 (N_6356,N_6217,N_6180);
xor U6357 (N_6357,N_6193,N_6226);
nor U6358 (N_6358,N_6141,N_6105);
nor U6359 (N_6359,N_6168,N_6045);
and U6360 (N_6360,N_6098,N_6059);
nor U6361 (N_6361,N_6121,N_6186);
and U6362 (N_6362,N_6017,N_6173);
nor U6363 (N_6363,N_6154,N_6044);
nand U6364 (N_6364,N_6080,N_6134);
nor U6365 (N_6365,N_6089,N_6178);
and U6366 (N_6366,N_6088,N_6036);
and U6367 (N_6367,N_6117,N_6208);
nand U6368 (N_6368,N_6145,N_6126);
and U6369 (N_6369,N_6130,N_6083);
nand U6370 (N_6370,N_6102,N_6201);
nand U6371 (N_6371,N_6228,N_6159);
xor U6372 (N_6372,N_6055,N_6047);
nor U6373 (N_6373,N_6122,N_6222);
or U6374 (N_6374,N_6169,N_6116);
and U6375 (N_6375,N_6061,N_6235);
nor U6376 (N_6376,N_6160,N_6067);
or U6377 (N_6377,N_6152,N_6105);
nand U6378 (N_6378,N_6096,N_6237);
nor U6379 (N_6379,N_6009,N_6002);
nand U6380 (N_6380,N_6218,N_6168);
and U6381 (N_6381,N_6239,N_6049);
nand U6382 (N_6382,N_6148,N_6157);
nand U6383 (N_6383,N_6224,N_6011);
or U6384 (N_6384,N_6095,N_6010);
or U6385 (N_6385,N_6211,N_6170);
xor U6386 (N_6386,N_6149,N_6168);
and U6387 (N_6387,N_6143,N_6220);
or U6388 (N_6388,N_6077,N_6017);
or U6389 (N_6389,N_6203,N_6241);
nand U6390 (N_6390,N_6190,N_6022);
nor U6391 (N_6391,N_6202,N_6148);
nor U6392 (N_6392,N_6066,N_6095);
or U6393 (N_6393,N_6102,N_6108);
and U6394 (N_6394,N_6241,N_6095);
and U6395 (N_6395,N_6031,N_6104);
xor U6396 (N_6396,N_6129,N_6063);
xnor U6397 (N_6397,N_6057,N_6132);
nor U6398 (N_6398,N_6176,N_6021);
and U6399 (N_6399,N_6064,N_6013);
or U6400 (N_6400,N_6117,N_6015);
or U6401 (N_6401,N_6060,N_6043);
or U6402 (N_6402,N_6017,N_6242);
and U6403 (N_6403,N_6150,N_6122);
nand U6404 (N_6404,N_6012,N_6169);
or U6405 (N_6405,N_6098,N_6128);
nor U6406 (N_6406,N_6052,N_6093);
and U6407 (N_6407,N_6115,N_6026);
or U6408 (N_6408,N_6074,N_6093);
xnor U6409 (N_6409,N_6109,N_6223);
nand U6410 (N_6410,N_6161,N_6244);
xnor U6411 (N_6411,N_6009,N_6096);
and U6412 (N_6412,N_6034,N_6104);
nand U6413 (N_6413,N_6089,N_6008);
nor U6414 (N_6414,N_6220,N_6108);
xor U6415 (N_6415,N_6003,N_6145);
nand U6416 (N_6416,N_6232,N_6159);
xor U6417 (N_6417,N_6244,N_6115);
xor U6418 (N_6418,N_6136,N_6206);
nand U6419 (N_6419,N_6100,N_6154);
nand U6420 (N_6420,N_6166,N_6185);
or U6421 (N_6421,N_6187,N_6199);
xnor U6422 (N_6422,N_6118,N_6219);
or U6423 (N_6423,N_6177,N_6025);
nor U6424 (N_6424,N_6164,N_6114);
xor U6425 (N_6425,N_6207,N_6106);
nor U6426 (N_6426,N_6070,N_6205);
nor U6427 (N_6427,N_6119,N_6203);
xor U6428 (N_6428,N_6223,N_6116);
nor U6429 (N_6429,N_6187,N_6120);
or U6430 (N_6430,N_6175,N_6220);
and U6431 (N_6431,N_6248,N_6241);
and U6432 (N_6432,N_6018,N_6168);
or U6433 (N_6433,N_6007,N_6055);
or U6434 (N_6434,N_6184,N_6111);
or U6435 (N_6435,N_6141,N_6242);
xor U6436 (N_6436,N_6134,N_6083);
nor U6437 (N_6437,N_6044,N_6226);
and U6438 (N_6438,N_6093,N_6149);
or U6439 (N_6439,N_6209,N_6111);
nand U6440 (N_6440,N_6152,N_6004);
nand U6441 (N_6441,N_6118,N_6187);
and U6442 (N_6442,N_6194,N_6071);
nand U6443 (N_6443,N_6025,N_6009);
and U6444 (N_6444,N_6007,N_6136);
nand U6445 (N_6445,N_6225,N_6208);
and U6446 (N_6446,N_6087,N_6248);
and U6447 (N_6447,N_6046,N_6083);
nand U6448 (N_6448,N_6144,N_6076);
or U6449 (N_6449,N_6163,N_6071);
nor U6450 (N_6450,N_6177,N_6238);
and U6451 (N_6451,N_6085,N_6084);
xor U6452 (N_6452,N_6164,N_6070);
nor U6453 (N_6453,N_6105,N_6186);
nor U6454 (N_6454,N_6186,N_6114);
xnor U6455 (N_6455,N_6180,N_6160);
xor U6456 (N_6456,N_6050,N_6184);
or U6457 (N_6457,N_6206,N_6238);
and U6458 (N_6458,N_6165,N_6189);
and U6459 (N_6459,N_6058,N_6032);
or U6460 (N_6460,N_6167,N_6073);
and U6461 (N_6461,N_6129,N_6208);
or U6462 (N_6462,N_6191,N_6023);
nand U6463 (N_6463,N_6240,N_6134);
xor U6464 (N_6464,N_6206,N_6102);
or U6465 (N_6465,N_6100,N_6006);
nand U6466 (N_6466,N_6047,N_6102);
nand U6467 (N_6467,N_6086,N_6247);
nand U6468 (N_6468,N_6061,N_6128);
nand U6469 (N_6469,N_6169,N_6074);
and U6470 (N_6470,N_6141,N_6122);
nor U6471 (N_6471,N_6165,N_6072);
or U6472 (N_6472,N_6159,N_6235);
and U6473 (N_6473,N_6167,N_6089);
or U6474 (N_6474,N_6171,N_6193);
nand U6475 (N_6475,N_6077,N_6111);
nand U6476 (N_6476,N_6060,N_6113);
xor U6477 (N_6477,N_6237,N_6228);
nor U6478 (N_6478,N_6038,N_6012);
or U6479 (N_6479,N_6248,N_6226);
nand U6480 (N_6480,N_6067,N_6214);
nand U6481 (N_6481,N_6208,N_6005);
nor U6482 (N_6482,N_6039,N_6212);
xor U6483 (N_6483,N_6243,N_6170);
and U6484 (N_6484,N_6066,N_6047);
and U6485 (N_6485,N_6111,N_6052);
and U6486 (N_6486,N_6128,N_6084);
nor U6487 (N_6487,N_6004,N_6219);
or U6488 (N_6488,N_6239,N_6041);
nor U6489 (N_6489,N_6043,N_6157);
or U6490 (N_6490,N_6121,N_6024);
or U6491 (N_6491,N_6181,N_6026);
nand U6492 (N_6492,N_6058,N_6125);
and U6493 (N_6493,N_6106,N_6005);
or U6494 (N_6494,N_6003,N_6241);
xor U6495 (N_6495,N_6141,N_6077);
and U6496 (N_6496,N_6107,N_6095);
nor U6497 (N_6497,N_6016,N_6185);
xnor U6498 (N_6498,N_6208,N_6122);
nor U6499 (N_6499,N_6109,N_6007);
or U6500 (N_6500,N_6365,N_6409);
nand U6501 (N_6501,N_6271,N_6332);
nand U6502 (N_6502,N_6465,N_6281);
nand U6503 (N_6503,N_6319,N_6385);
nor U6504 (N_6504,N_6287,N_6478);
nor U6505 (N_6505,N_6337,N_6393);
xnor U6506 (N_6506,N_6481,N_6480);
xor U6507 (N_6507,N_6426,N_6302);
xnor U6508 (N_6508,N_6402,N_6423);
and U6509 (N_6509,N_6380,N_6288);
xor U6510 (N_6510,N_6397,N_6286);
nand U6511 (N_6511,N_6311,N_6276);
nand U6512 (N_6512,N_6359,N_6340);
and U6513 (N_6513,N_6326,N_6432);
xnor U6514 (N_6514,N_6289,N_6491);
nor U6515 (N_6515,N_6394,N_6318);
xor U6516 (N_6516,N_6355,N_6327);
and U6517 (N_6517,N_6403,N_6382);
nand U6518 (N_6518,N_6298,N_6371);
and U6519 (N_6519,N_6396,N_6294);
xor U6520 (N_6520,N_6454,N_6277);
xor U6521 (N_6521,N_6368,N_6308);
nand U6522 (N_6522,N_6344,N_6448);
nand U6523 (N_6523,N_6364,N_6429);
xnor U6524 (N_6524,N_6456,N_6415);
and U6525 (N_6525,N_6291,N_6490);
nand U6526 (N_6526,N_6439,N_6485);
and U6527 (N_6527,N_6328,N_6341);
and U6528 (N_6528,N_6280,N_6436);
or U6529 (N_6529,N_6475,N_6353);
or U6530 (N_6530,N_6292,N_6401);
nand U6531 (N_6531,N_6453,N_6314);
and U6532 (N_6532,N_6321,N_6306);
and U6533 (N_6533,N_6483,N_6356);
xnor U6534 (N_6534,N_6305,N_6282);
xor U6535 (N_6535,N_6357,N_6455);
xnor U6536 (N_6536,N_6495,N_6474);
or U6537 (N_6537,N_6346,N_6461);
xor U6538 (N_6538,N_6378,N_6450);
nor U6539 (N_6539,N_6303,N_6384);
nand U6540 (N_6540,N_6431,N_6472);
xnor U6541 (N_6541,N_6320,N_6441);
xor U6542 (N_6542,N_6445,N_6343);
and U6543 (N_6543,N_6451,N_6304);
nand U6544 (N_6544,N_6492,N_6351);
nand U6545 (N_6545,N_6466,N_6388);
nand U6546 (N_6546,N_6416,N_6295);
nand U6547 (N_6547,N_6489,N_6443);
nor U6548 (N_6548,N_6331,N_6458);
nor U6549 (N_6549,N_6473,N_6285);
nor U6550 (N_6550,N_6470,N_6412);
nand U6551 (N_6551,N_6310,N_6421);
or U6552 (N_6552,N_6299,N_6354);
xnor U6553 (N_6553,N_6442,N_6376);
and U6554 (N_6554,N_6391,N_6379);
nand U6555 (N_6555,N_6381,N_6390);
xnor U6556 (N_6556,N_6283,N_6336);
nand U6557 (N_6557,N_6392,N_6476);
and U6558 (N_6558,N_6313,N_6496);
or U6559 (N_6559,N_6348,N_6422);
xnor U6560 (N_6560,N_6417,N_6437);
and U6561 (N_6561,N_6463,N_6316);
nand U6562 (N_6562,N_6352,N_6400);
nand U6563 (N_6563,N_6263,N_6279);
xor U6564 (N_6564,N_6251,N_6389);
xnor U6565 (N_6565,N_6301,N_6430);
xor U6566 (N_6566,N_6250,N_6494);
nand U6567 (N_6567,N_6372,N_6407);
xor U6568 (N_6568,N_6383,N_6497);
nor U6569 (N_6569,N_6484,N_6449);
xor U6570 (N_6570,N_6322,N_6387);
nand U6571 (N_6571,N_6469,N_6405);
nor U6572 (N_6572,N_6488,N_6427);
nand U6573 (N_6573,N_6452,N_6374);
xor U6574 (N_6574,N_6444,N_6375);
nor U6575 (N_6575,N_6425,N_6369);
xnor U6576 (N_6576,N_6404,N_6419);
nand U6577 (N_6577,N_6261,N_6339);
nand U6578 (N_6578,N_6307,N_6459);
and U6579 (N_6579,N_6269,N_6267);
xnor U6580 (N_6580,N_6462,N_6347);
xor U6581 (N_6581,N_6499,N_6350);
or U6582 (N_6582,N_6498,N_6256);
nor U6583 (N_6583,N_6254,N_6482);
nor U6584 (N_6584,N_6414,N_6424);
or U6585 (N_6585,N_6323,N_6366);
or U6586 (N_6586,N_6329,N_6438);
nand U6587 (N_6587,N_6428,N_6487);
or U6588 (N_6588,N_6486,N_6370);
xor U6589 (N_6589,N_6335,N_6258);
nor U6590 (N_6590,N_6260,N_6367);
xnor U6591 (N_6591,N_6358,N_6433);
nand U6592 (N_6592,N_6262,N_6408);
nand U6593 (N_6593,N_6398,N_6274);
and U6594 (N_6594,N_6278,N_6467);
or U6595 (N_6595,N_6296,N_6464);
nand U6596 (N_6596,N_6471,N_6373);
nand U6597 (N_6597,N_6457,N_6312);
and U6598 (N_6598,N_6293,N_6460);
or U6599 (N_6599,N_6255,N_6440);
or U6600 (N_6600,N_6363,N_6411);
or U6601 (N_6601,N_6317,N_6420);
nand U6602 (N_6602,N_6360,N_6290);
or U6603 (N_6603,N_6268,N_6309);
nor U6604 (N_6604,N_6333,N_6479);
xor U6605 (N_6605,N_6435,N_6253);
and U6606 (N_6606,N_6395,N_6434);
nor U6607 (N_6607,N_6264,N_6345);
and U6608 (N_6608,N_6266,N_6477);
nand U6609 (N_6609,N_6297,N_6273);
xor U6610 (N_6610,N_6493,N_6446);
nor U6611 (N_6611,N_6418,N_6300);
nand U6612 (N_6612,N_6406,N_6315);
xor U6613 (N_6613,N_6330,N_6265);
xnor U6614 (N_6614,N_6399,N_6447);
or U6615 (N_6615,N_6272,N_6342);
nand U6616 (N_6616,N_6362,N_6252);
and U6617 (N_6617,N_6386,N_6410);
nor U6618 (N_6618,N_6284,N_6324);
and U6619 (N_6619,N_6377,N_6270);
or U6620 (N_6620,N_6349,N_6325);
nor U6621 (N_6621,N_6259,N_6257);
xnor U6622 (N_6622,N_6275,N_6361);
and U6623 (N_6623,N_6413,N_6338);
or U6624 (N_6624,N_6468,N_6334);
xnor U6625 (N_6625,N_6268,N_6405);
xor U6626 (N_6626,N_6292,N_6344);
and U6627 (N_6627,N_6496,N_6363);
nor U6628 (N_6628,N_6285,N_6361);
nor U6629 (N_6629,N_6457,N_6305);
or U6630 (N_6630,N_6366,N_6469);
xor U6631 (N_6631,N_6263,N_6447);
nor U6632 (N_6632,N_6464,N_6437);
nor U6633 (N_6633,N_6332,N_6334);
nor U6634 (N_6634,N_6453,N_6312);
nand U6635 (N_6635,N_6336,N_6461);
nor U6636 (N_6636,N_6437,N_6300);
and U6637 (N_6637,N_6498,N_6364);
xnor U6638 (N_6638,N_6436,N_6474);
and U6639 (N_6639,N_6259,N_6311);
xor U6640 (N_6640,N_6454,N_6437);
xnor U6641 (N_6641,N_6301,N_6330);
or U6642 (N_6642,N_6389,N_6337);
and U6643 (N_6643,N_6304,N_6299);
nand U6644 (N_6644,N_6373,N_6353);
nand U6645 (N_6645,N_6268,N_6266);
xnor U6646 (N_6646,N_6271,N_6433);
nor U6647 (N_6647,N_6367,N_6275);
nor U6648 (N_6648,N_6369,N_6384);
and U6649 (N_6649,N_6291,N_6495);
or U6650 (N_6650,N_6302,N_6278);
xnor U6651 (N_6651,N_6253,N_6421);
nand U6652 (N_6652,N_6270,N_6299);
and U6653 (N_6653,N_6407,N_6402);
and U6654 (N_6654,N_6451,N_6417);
and U6655 (N_6655,N_6324,N_6398);
or U6656 (N_6656,N_6343,N_6357);
or U6657 (N_6657,N_6293,N_6378);
nor U6658 (N_6658,N_6441,N_6313);
nand U6659 (N_6659,N_6273,N_6415);
xnor U6660 (N_6660,N_6450,N_6411);
nor U6661 (N_6661,N_6458,N_6304);
nor U6662 (N_6662,N_6492,N_6368);
or U6663 (N_6663,N_6334,N_6457);
or U6664 (N_6664,N_6274,N_6381);
and U6665 (N_6665,N_6261,N_6432);
or U6666 (N_6666,N_6434,N_6333);
xnor U6667 (N_6667,N_6301,N_6356);
and U6668 (N_6668,N_6309,N_6399);
and U6669 (N_6669,N_6276,N_6301);
xor U6670 (N_6670,N_6350,N_6361);
nor U6671 (N_6671,N_6359,N_6264);
nand U6672 (N_6672,N_6491,N_6336);
nor U6673 (N_6673,N_6285,N_6483);
xor U6674 (N_6674,N_6446,N_6393);
and U6675 (N_6675,N_6257,N_6303);
and U6676 (N_6676,N_6471,N_6433);
xnor U6677 (N_6677,N_6457,N_6452);
nand U6678 (N_6678,N_6354,N_6486);
or U6679 (N_6679,N_6489,N_6307);
xnor U6680 (N_6680,N_6380,N_6445);
or U6681 (N_6681,N_6493,N_6320);
or U6682 (N_6682,N_6340,N_6401);
or U6683 (N_6683,N_6420,N_6405);
nor U6684 (N_6684,N_6471,N_6388);
xnor U6685 (N_6685,N_6290,N_6485);
xor U6686 (N_6686,N_6400,N_6309);
nand U6687 (N_6687,N_6251,N_6489);
nand U6688 (N_6688,N_6376,N_6315);
or U6689 (N_6689,N_6393,N_6290);
nor U6690 (N_6690,N_6434,N_6422);
nand U6691 (N_6691,N_6351,N_6346);
nor U6692 (N_6692,N_6493,N_6262);
xor U6693 (N_6693,N_6324,N_6353);
or U6694 (N_6694,N_6479,N_6388);
and U6695 (N_6695,N_6327,N_6254);
nor U6696 (N_6696,N_6413,N_6482);
nor U6697 (N_6697,N_6271,N_6297);
or U6698 (N_6698,N_6427,N_6313);
and U6699 (N_6699,N_6356,N_6320);
nand U6700 (N_6700,N_6398,N_6468);
xnor U6701 (N_6701,N_6476,N_6344);
nor U6702 (N_6702,N_6339,N_6251);
or U6703 (N_6703,N_6452,N_6497);
or U6704 (N_6704,N_6382,N_6308);
and U6705 (N_6705,N_6461,N_6260);
or U6706 (N_6706,N_6465,N_6376);
nand U6707 (N_6707,N_6413,N_6390);
or U6708 (N_6708,N_6317,N_6353);
and U6709 (N_6709,N_6422,N_6289);
nand U6710 (N_6710,N_6325,N_6251);
nand U6711 (N_6711,N_6286,N_6455);
nor U6712 (N_6712,N_6309,N_6421);
and U6713 (N_6713,N_6487,N_6381);
nor U6714 (N_6714,N_6487,N_6482);
and U6715 (N_6715,N_6320,N_6275);
nand U6716 (N_6716,N_6271,N_6256);
nor U6717 (N_6717,N_6392,N_6397);
and U6718 (N_6718,N_6378,N_6373);
xnor U6719 (N_6719,N_6357,N_6344);
and U6720 (N_6720,N_6429,N_6381);
xor U6721 (N_6721,N_6316,N_6416);
nor U6722 (N_6722,N_6399,N_6332);
xnor U6723 (N_6723,N_6375,N_6446);
xor U6724 (N_6724,N_6343,N_6423);
and U6725 (N_6725,N_6427,N_6446);
nand U6726 (N_6726,N_6307,N_6310);
and U6727 (N_6727,N_6450,N_6442);
nand U6728 (N_6728,N_6336,N_6449);
or U6729 (N_6729,N_6308,N_6267);
xnor U6730 (N_6730,N_6359,N_6327);
or U6731 (N_6731,N_6372,N_6441);
nand U6732 (N_6732,N_6495,N_6294);
xnor U6733 (N_6733,N_6362,N_6402);
nor U6734 (N_6734,N_6488,N_6315);
nand U6735 (N_6735,N_6407,N_6350);
or U6736 (N_6736,N_6304,N_6278);
xor U6737 (N_6737,N_6411,N_6264);
or U6738 (N_6738,N_6324,N_6419);
or U6739 (N_6739,N_6353,N_6282);
and U6740 (N_6740,N_6397,N_6367);
nor U6741 (N_6741,N_6481,N_6408);
nor U6742 (N_6742,N_6292,N_6479);
and U6743 (N_6743,N_6463,N_6266);
and U6744 (N_6744,N_6250,N_6324);
and U6745 (N_6745,N_6277,N_6368);
or U6746 (N_6746,N_6350,N_6420);
nand U6747 (N_6747,N_6342,N_6469);
or U6748 (N_6748,N_6325,N_6410);
and U6749 (N_6749,N_6250,N_6428);
nor U6750 (N_6750,N_6503,N_6646);
xnor U6751 (N_6751,N_6742,N_6687);
nor U6752 (N_6752,N_6634,N_6669);
and U6753 (N_6753,N_6746,N_6557);
nor U6754 (N_6754,N_6511,N_6610);
xnor U6755 (N_6755,N_6627,N_6533);
nand U6756 (N_6756,N_6692,N_6624);
xor U6757 (N_6757,N_6621,N_6611);
xor U6758 (N_6758,N_6714,N_6662);
or U6759 (N_6759,N_6561,N_6694);
or U6760 (N_6760,N_6528,N_6679);
xor U6761 (N_6761,N_6659,N_6600);
or U6762 (N_6762,N_6513,N_6631);
nand U6763 (N_6763,N_6520,N_6607);
nor U6764 (N_6764,N_6652,N_6717);
or U6765 (N_6765,N_6507,N_6743);
nor U6766 (N_6766,N_6550,N_6586);
and U6767 (N_6767,N_6749,N_6535);
or U6768 (N_6768,N_6551,N_6504);
or U6769 (N_6769,N_6565,N_6614);
nor U6770 (N_6770,N_6518,N_6726);
and U6771 (N_6771,N_6566,N_6649);
xnor U6772 (N_6772,N_6625,N_6602);
nand U6773 (N_6773,N_6695,N_6672);
or U6774 (N_6774,N_6530,N_6578);
or U6775 (N_6775,N_6623,N_6709);
or U6776 (N_6776,N_6597,N_6556);
or U6777 (N_6777,N_6689,N_6510);
nor U6778 (N_6778,N_6591,N_6590);
xnor U6779 (N_6779,N_6706,N_6571);
nor U6780 (N_6780,N_6554,N_6637);
and U6781 (N_6781,N_6502,N_6515);
xnor U6782 (N_6782,N_6526,N_6645);
and U6783 (N_6783,N_6710,N_6541);
xnor U6784 (N_6784,N_6639,N_6540);
nor U6785 (N_6785,N_6579,N_6673);
xor U6786 (N_6786,N_6643,N_6740);
and U6787 (N_6787,N_6638,N_6564);
xnor U6788 (N_6788,N_6674,N_6592);
nand U6789 (N_6789,N_6555,N_6720);
and U6790 (N_6790,N_6716,N_6676);
nand U6791 (N_6791,N_6626,N_6722);
or U6792 (N_6792,N_6707,N_6664);
nor U6793 (N_6793,N_6558,N_6713);
or U6794 (N_6794,N_6699,N_6567);
nor U6795 (N_6795,N_6516,N_6616);
nor U6796 (N_6796,N_6500,N_6609);
or U6797 (N_6797,N_6545,N_6577);
nand U6798 (N_6798,N_6527,N_6598);
xnor U6799 (N_6799,N_6543,N_6663);
nand U6800 (N_6800,N_6708,N_6678);
nor U6801 (N_6801,N_6568,N_6636);
nand U6802 (N_6802,N_6681,N_6622);
nand U6803 (N_6803,N_6601,N_6506);
and U6804 (N_6804,N_6712,N_6547);
nand U6805 (N_6805,N_6711,N_6501);
or U6806 (N_6806,N_6613,N_6514);
nand U6807 (N_6807,N_6732,N_6584);
xor U6808 (N_6808,N_6575,N_6635);
nor U6809 (N_6809,N_6683,N_6559);
and U6810 (N_6810,N_6741,N_6728);
or U6811 (N_6811,N_6606,N_6671);
and U6812 (N_6812,N_6724,N_6680);
and U6813 (N_6813,N_6594,N_6619);
xnor U6814 (N_6814,N_6542,N_6744);
and U6815 (N_6815,N_6719,N_6748);
xnor U6816 (N_6816,N_6560,N_6739);
xor U6817 (N_6817,N_6629,N_6675);
nor U6818 (N_6818,N_6529,N_6587);
xnor U6819 (N_6819,N_6546,N_6654);
nor U6820 (N_6820,N_6698,N_6553);
and U6821 (N_6821,N_6688,N_6736);
and U6822 (N_6822,N_6677,N_6697);
or U6823 (N_6823,N_6737,N_6653);
or U6824 (N_6824,N_6620,N_6604);
xnor U6825 (N_6825,N_6572,N_6523);
xor U6826 (N_6826,N_6632,N_6738);
xor U6827 (N_6827,N_6747,N_6524);
and U6828 (N_6828,N_6727,N_6605);
nand U6829 (N_6829,N_6603,N_6508);
nor U6830 (N_6830,N_6595,N_6721);
xnor U6831 (N_6831,N_6563,N_6648);
xor U6832 (N_6832,N_6618,N_6705);
xnor U6833 (N_6833,N_6667,N_6733);
nor U6834 (N_6834,N_6644,N_6641);
and U6835 (N_6835,N_6593,N_6682);
xnor U6836 (N_6836,N_6581,N_6745);
nand U6837 (N_6837,N_6525,N_6690);
and U6838 (N_6838,N_6723,N_6725);
nand U6839 (N_6839,N_6534,N_6655);
and U6840 (N_6840,N_6693,N_6651);
xnor U6841 (N_6841,N_6589,N_6574);
and U6842 (N_6842,N_6537,N_6701);
and U6843 (N_6843,N_6532,N_6617);
or U6844 (N_6844,N_6730,N_6596);
nand U6845 (N_6845,N_6647,N_6612);
xnor U6846 (N_6846,N_6583,N_6562);
or U6847 (N_6847,N_6715,N_6729);
or U6848 (N_6848,N_6585,N_6718);
xor U6849 (N_6849,N_6538,N_6657);
nor U6850 (N_6850,N_6633,N_6696);
or U6851 (N_6851,N_6734,N_6685);
nor U6852 (N_6852,N_6630,N_6656);
xnor U6853 (N_6853,N_6552,N_6544);
xnor U6854 (N_6854,N_6684,N_6608);
nor U6855 (N_6855,N_6569,N_6731);
nand U6856 (N_6856,N_6536,N_6522);
nand U6857 (N_6857,N_6512,N_6570);
xor U6858 (N_6858,N_6691,N_6599);
and U6859 (N_6859,N_6580,N_6573);
nand U6860 (N_6860,N_6700,N_6661);
nand U6861 (N_6861,N_6582,N_6642);
and U6862 (N_6862,N_6640,N_6549);
xnor U6863 (N_6863,N_6686,N_6668);
and U6864 (N_6864,N_6509,N_6666);
and U6865 (N_6865,N_6517,N_6539);
or U6866 (N_6866,N_6519,N_6704);
xnor U6867 (N_6867,N_6702,N_6521);
and U6868 (N_6868,N_6660,N_6588);
nor U6869 (N_6869,N_6665,N_6735);
or U6870 (N_6870,N_6628,N_6615);
nor U6871 (N_6871,N_6658,N_6703);
and U6872 (N_6872,N_6576,N_6531);
xnor U6873 (N_6873,N_6548,N_6505);
nand U6874 (N_6874,N_6650,N_6670);
xnor U6875 (N_6875,N_6579,N_6604);
nor U6876 (N_6876,N_6655,N_6707);
or U6877 (N_6877,N_6658,N_6526);
and U6878 (N_6878,N_6733,N_6701);
nand U6879 (N_6879,N_6685,N_6744);
and U6880 (N_6880,N_6566,N_6620);
or U6881 (N_6881,N_6680,N_6601);
or U6882 (N_6882,N_6516,N_6506);
or U6883 (N_6883,N_6579,N_6615);
nor U6884 (N_6884,N_6562,N_6673);
xor U6885 (N_6885,N_6565,N_6525);
or U6886 (N_6886,N_6572,N_6540);
nor U6887 (N_6887,N_6555,N_6525);
nand U6888 (N_6888,N_6546,N_6513);
and U6889 (N_6889,N_6566,N_6671);
and U6890 (N_6890,N_6594,N_6535);
or U6891 (N_6891,N_6647,N_6645);
nand U6892 (N_6892,N_6675,N_6661);
or U6893 (N_6893,N_6604,N_6501);
and U6894 (N_6894,N_6617,N_6542);
nand U6895 (N_6895,N_6635,N_6539);
nor U6896 (N_6896,N_6625,N_6731);
or U6897 (N_6897,N_6686,N_6683);
or U6898 (N_6898,N_6532,N_6530);
or U6899 (N_6899,N_6576,N_6720);
nand U6900 (N_6900,N_6512,N_6536);
or U6901 (N_6901,N_6585,N_6639);
nand U6902 (N_6902,N_6688,N_6714);
and U6903 (N_6903,N_6500,N_6550);
xnor U6904 (N_6904,N_6528,N_6653);
and U6905 (N_6905,N_6548,N_6534);
xnor U6906 (N_6906,N_6505,N_6740);
and U6907 (N_6907,N_6562,N_6684);
nand U6908 (N_6908,N_6676,N_6637);
or U6909 (N_6909,N_6685,N_6688);
and U6910 (N_6910,N_6601,N_6562);
nor U6911 (N_6911,N_6706,N_6608);
or U6912 (N_6912,N_6615,N_6675);
nor U6913 (N_6913,N_6693,N_6691);
and U6914 (N_6914,N_6651,N_6501);
nand U6915 (N_6915,N_6618,N_6743);
or U6916 (N_6916,N_6523,N_6727);
and U6917 (N_6917,N_6550,N_6668);
and U6918 (N_6918,N_6526,N_6628);
or U6919 (N_6919,N_6588,N_6734);
nand U6920 (N_6920,N_6748,N_6634);
or U6921 (N_6921,N_6694,N_6514);
nand U6922 (N_6922,N_6674,N_6571);
nand U6923 (N_6923,N_6589,N_6604);
and U6924 (N_6924,N_6608,N_6509);
or U6925 (N_6925,N_6617,N_6656);
nor U6926 (N_6926,N_6609,N_6729);
xnor U6927 (N_6927,N_6556,N_6551);
nand U6928 (N_6928,N_6686,N_6653);
or U6929 (N_6929,N_6656,N_6607);
or U6930 (N_6930,N_6730,N_6710);
xnor U6931 (N_6931,N_6557,N_6514);
xnor U6932 (N_6932,N_6516,N_6685);
nand U6933 (N_6933,N_6571,N_6605);
nor U6934 (N_6934,N_6648,N_6635);
nand U6935 (N_6935,N_6698,N_6726);
xor U6936 (N_6936,N_6725,N_6733);
and U6937 (N_6937,N_6748,N_6609);
nor U6938 (N_6938,N_6668,N_6746);
nor U6939 (N_6939,N_6594,N_6740);
nand U6940 (N_6940,N_6743,N_6690);
and U6941 (N_6941,N_6684,N_6631);
xnor U6942 (N_6942,N_6513,N_6609);
nor U6943 (N_6943,N_6706,N_6715);
and U6944 (N_6944,N_6583,N_6561);
nor U6945 (N_6945,N_6578,N_6700);
nand U6946 (N_6946,N_6584,N_6695);
or U6947 (N_6947,N_6569,N_6661);
nand U6948 (N_6948,N_6581,N_6504);
or U6949 (N_6949,N_6566,N_6504);
and U6950 (N_6950,N_6583,N_6683);
nand U6951 (N_6951,N_6543,N_6647);
nand U6952 (N_6952,N_6651,N_6638);
nand U6953 (N_6953,N_6744,N_6627);
nor U6954 (N_6954,N_6748,N_6547);
nand U6955 (N_6955,N_6580,N_6594);
xnor U6956 (N_6956,N_6674,N_6650);
or U6957 (N_6957,N_6561,N_6743);
nor U6958 (N_6958,N_6529,N_6579);
nor U6959 (N_6959,N_6608,N_6568);
nor U6960 (N_6960,N_6736,N_6505);
nand U6961 (N_6961,N_6677,N_6644);
or U6962 (N_6962,N_6661,N_6720);
or U6963 (N_6963,N_6628,N_6631);
and U6964 (N_6964,N_6656,N_6639);
or U6965 (N_6965,N_6518,N_6695);
or U6966 (N_6966,N_6532,N_6745);
and U6967 (N_6967,N_6720,N_6558);
or U6968 (N_6968,N_6513,N_6690);
xnor U6969 (N_6969,N_6502,N_6691);
or U6970 (N_6970,N_6520,N_6585);
xnor U6971 (N_6971,N_6616,N_6729);
xor U6972 (N_6972,N_6524,N_6655);
xnor U6973 (N_6973,N_6677,N_6682);
nor U6974 (N_6974,N_6596,N_6722);
or U6975 (N_6975,N_6620,N_6682);
xnor U6976 (N_6976,N_6712,N_6657);
nor U6977 (N_6977,N_6570,N_6649);
nand U6978 (N_6978,N_6700,N_6599);
and U6979 (N_6979,N_6679,N_6672);
xnor U6980 (N_6980,N_6515,N_6648);
nand U6981 (N_6981,N_6701,N_6650);
and U6982 (N_6982,N_6745,N_6537);
and U6983 (N_6983,N_6678,N_6703);
xnor U6984 (N_6984,N_6675,N_6501);
or U6985 (N_6985,N_6679,N_6564);
or U6986 (N_6986,N_6603,N_6621);
nor U6987 (N_6987,N_6642,N_6737);
xnor U6988 (N_6988,N_6555,N_6594);
xor U6989 (N_6989,N_6693,N_6631);
nand U6990 (N_6990,N_6670,N_6607);
and U6991 (N_6991,N_6723,N_6644);
nor U6992 (N_6992,N_6643,N_6739);
and U6993 (N_6993,N_6632,N_6586);
nand U6994 (N_6994,N_6603,N_6667);
or U6995 (N_6995,N_6642,N_6734);
nor U6996 (N_6996,N_6597,N_6532);
nor U6997 (N_6997,N_6519,N_6657);
xnor U6998 (N_6998,N_6634,N_6567);
nor U6999 (N_6999,N_6634,N_6514);
and U7000 (N_7000,N_6875,N_6958);
and U7001 (N_7001,N_6935,N_6985);
nand U7002 (N_7002,N_6786,N_6976);
nand U7003 (N_7003,N_6889,N_6913);
nand U7004 (N_7004,N_6772,N_6984);
nand U7005 (N_7005,N_6845,N_6816);
nor U7006 (N_7006,N_6957,N_6789);
or U7007 (N_7007,N_6812,N_6930);
nand U7008 (N_7008,N_6826,N_6847);
nand U7009 (N_7009,N_6782,N_6751);
and U7010 (N_7010,N_6840,N_6953);
nand U7011 (N_7011,N_6762,N_6983);
or U7012 (N_7012,N_6954,N_6823);
and U7013 (N_7013,N_6862,N_6902);
xnor U7014 (N_7014,N_6970,N_6821);
nor U7015 (N_7015,N_6947,N_6837);
nor U7016 (N_7016,N_6835,N_6820);
or U7017 (N_7017,N_6892,N_6886);
or U7018 (N_7018,N_6778,N_6885);
nor U7019 (N_7019,N_6859,N_6978);
nand U7020 (N_7020,N_6924,N_6829);
nor U7021 (N_7021,N_6941,N_6940);
or U7022 (N_7022,N_6931,N_6894);
nand U7023 (N_7023,N_6761,N_6766);
nand U7024 (N_7024,N_6819,N_6945);
and U7025 (N_7025,N_6896,N_6763);
nand U7026 (N_7026,N_6906,N_6877);
nor U7027 (N_7027,N_6998,N_6863);
nand U7028 (N_7028,N_6769,N_6815);
or U7029 (N_7029,N_6884,N_6839);
nand U7030 (N_7030,N_6943,N_6944);
or U7031 (N_7031,N_6880,N_6950);
nor U7032 (N_7032,N_6755,N_6759);
or U7033 (N_7033,N_6974,N_6929);
or U7034 (N_7034,N_6868,N_6911);
and U7035 (N_7035,N_6897,N_6919);
or U7036 (N_7036,N_6858,N_6901);
nand U7037 (N_7037,N_6948,N_6787);
nand U7038 (N_7038,N_6851,N_6914);
or U7039 (N_7039,N_6758,N_6836);
or U7040 (N_7040,N_6986,N_6883);
nor U7041 (N_7041,N_6770,N_6799);
or U7042 (N_7042,N_6952,N_6916);
or U7043 (N_7043,N_6971,N_6874);
or U7044 (N_7044,N_6951,N_6963);
or U7045 (N_7045,N_6895,N_6955);
nand U7046 (N_7046,N_6798,N_6779);
or U7047 (N_7047,N_6962,N_6818);
or U7048 (N_7048,N_6805,N_6804);
and U7049 (N_7049,N_6822,N_6824);
xor U7050 (N_7050,N_6866,N_6871);
nor U7051 (N_7051,N_6795,N_6961);
and U7052 (N_7052,N_6898,N_6933);
nand U7053 (N_7053,N_6873,N_6993);
or U7054 (N_7054,N_6942,N_6852);
nand U7055 (N_7055,N_6785,N_6838);
or U7056 (N_7056,N_6774,N_6999);
and U7057 (N_7057,N_6792,N_6988);
xnor U7058 (N_7058,N_6893,N_6876);
and U7059 (N_7059,N_6922,N_6910);
or U7060 (N_7060,N_6887,N_6832);
and U7061 (N_7061,N_6844,N_6938);
nor U7062 (N_7062,N_6752,N_6932);
xnor U7063 (N_7063,N_6807,N_6793);
or U7064 (N_7064,N_6834,N_6857);
and U7065 (N_7065,N_6926,N_6814);
nor U7066 (N_7066,N_6972,N_6989);
xnor U7067 (N_7067,N_6960,N_6881);
xnor U7068 (N_7068,N_6765,N_6977);
nand U7069 (N_7069,N_6760,N_6937);
or U7070 (N_7070,N_6810,N_6850);
nor U7071 (N_7071,N_6797,N_6927);
or U7072 (N_7072,N_6904,N_6968);
xor U7073 (N_7073,N_6949,N_6980);
nand U7074 (N_7074,N_6921,N_6920);
nor U7075 (N_7075,N_6788,N_6907);
nand U7076 (N_7076,N_6775,N_6771);
or U7077 (N_7077,N_6939,N_6806);
nor U7078 (N_7078,N_6833,N_6796);
or U7079 (N_7079,N_6861,N_6811);
or U7080 (N_7080,N_6917,N_6783);
xor U7081 (N_7081,N_6813,N_6888);
or U7082 (N_7082,N_6990,N_6825);
or U7083 (N_7083,N_6856,N_6860);
and U7084 (N_7084,N_6973,N_6891);
xnor U7085 (N_7085,N_6843,N_6870);
or U7086 (N_7086,N_6979,N_6905);
nor U7087 (N_7087,N_6967,N_6790);
nand U7088 (N_7088,N_6848,N_6841);
nor U7089 (N_7089,N_6773,N_6754);
nor U7090 (N_7090,N_6981,N_6764);
and U7091 (N_7091,N_6809,N_6784);
nand U7092 (N_7092,N_6801,N_6828);
and U7093 (N_7093,N_6777,N_6994);
nand U7094 (N_7094,N_6975,N_6956);
nor U7095 (N_7095,N_6915,N_6872);
nor U7096 (N_7096,N_6959,N_6890);
nor U7097 (N_7097,N_6800,N_6879);
or U7098 (N_7098,N_6853,N_6918);
nand U7099 (N_7099,N_6928,N_6756);
or U7100 (N_7100,N_6842,N_6849);
nor U7101 (N_7101,N_6831,N_6864);
and U7102 (N_7102,N_6912,N_6846);
xor U7103 (N_7103,N_6794,N_6923);
nor U7104 (N_7104,N_6909,N_6903);
or U7105 (N_7105,N_6934,N_6803);
nor U7106 (N_7106,N_6925,N_6855);
nor U7107 (N_7107,N_6987,N_6817);
or U7108 (N_7108,N_6964,N_6882);
and U7109 (N_7109,N_6780,N_6776);
xor U7110 (N_7110,N_6992,N_6865);
or U7111 (N_7111,N_6830,N_6753);
and U7112 (N_7112,N_6969,N_6991);
nand U7113 (N_7113,N_6767,N_6791);
or U7114 (N_7114,N_6867,N_6995);
and U7115 (N_7115,N_6900,N_6965);
and U7116 (N_7116,N_6908,N_6869);
xnor U7117 (N_7117,N_6878,N_6996);
xor U7118 (N_7118,N_6827,N_6997);
and U7119 (N_7119,N_6966,N_6750);
nor U7120 (N_7120,N_6946,N_6854);
and U7121 (N_7121,N_6936,N_6982);
or U7122 (N_7122,N_6781,N_6808);
nor U7123 (N_7123,N_6768,N_6757);
nand U7124 (N_7124,N_6899,N_6802);
or U7125 (N_7125,N_6894,N_6881);
xnor U7126 (N_7126,N_6822,N_6875);
nand U7127 (N_7127,N_6933,N_6801);
nand U7128 (N_7128,N_6882,N_6932);
and U7129 (N_7129,N_6973,N_6909);
nor U7130 (N_7130,N_6907,N_6778);
nand U7131 (N_7131,N_6977,N_6988);
nor U7132 (N_7132,N_6811,N_6803);
xor U7133 (N_7133,N_6863,N_6890);
nor U7134 (N_7134,N_6858,N_6756);
nor U7135 (N_7135,N_6934,N_6935);
or U7136 (N_7136,N_6913,N_6774);
or U7137 (N_7137,N_6886,N_6896);
and U7138 (N_7138,N_6842,N_6920);
and U7139 (N_7139,N_6811,N_6985);
xnor U7140 (N_7140,N_6869,N_6848);
nand U7141 (N_7141,N_6902,N_6964);
xor U7142 (N_7142,N_6752,N_6977);
nor U7143 (N_7143,N_6960,N_6860);
or U7144 (N_7144,N_6917,N_6969);
nand U7145 (N_7145,N_6771,N_6829);
or U7146 (N_7146,N_6809,N_6944);
xnor U7147 (N_7147,N_6907,N_6949);
nand U7148 (N_7148,N_6768,N_6976);
xor U7149 (N_7149,N_6909,N_6875);
nor U7150 (N_7150,N_6762,N_6836);
nand U7151 (N_7151,N_6857,N_6835);
xor U7152 (N_7152,N_6927,N_6830);
and U7153 (N_7153,N_6774,N_6956);
xnor U7154 (N_7154,N_6961,N_6823);
or U7155 (N_7155,N_6992,N_6881);
or U7156 (N_7156,N_6951,N_6984);
or U7157 (N_7157,N_6766,N_6859);
nand U7158 (N_7158,N_6934,N_6783);
nor U7159 (N_7159,N_6756,N_6856);
or U7160 (N_7160,N_6921,N_6775);
nor U7161 (N_7161,N_6819,N_6846);
nand U7162 (N_7162,N_6961,N_6793);
nor U7163 (N_7163,N_6890,N_6948);
and U7164 (N_7164,N_6789,N_6775);
nand U7165 (N_7165,N_6997,N_6986);
and U7166 (N_7166,N_6844,N_6872);
or U7167 (N_7167,N_6961,N_6902);
xnor U7168 (N_7168,N_6922,N_6832);
xor U7169 (N_7169,N_6812,N_6887);
xor U7170 (N_7170,N_6935,N_6829);
and U7171 (N_7171,N_6822,N_6955);
xnor U7172 (N_7172,N_6907,N_6934);
xnor U7173 (N_7173,N_6884,N_6833);
or U7174 (N_7174,N_6996,N_6824);
and U7175 (N_7175,N_6850,N_6875);
and U7176 (N_7176,N_6847,N_6884);
or U7177 (N_7177,N_6951,N_6755);
and U7178 (N_7178,N_6913,N_6786);
and U7179 (N_7179,N_6798,N_6841);
nand U7180 (N_7180,N_6976,N_6764);
xor U7181 (N_7181,N_6984,N_6839);
nand U7182 (N_7182,N_6847,N_6900);
nand U7183 (N_7183,N_6884,N_6987);
nand U7184 (N_7184,N_6837,N_6930);
and U7185 (N_7185,N_6838,N_6935);
xor U7186 (N_7186,N_6854,N_6993);
nand U7187 (N_7187,N_6895,N_6909);
xor U7188 (N_7188,N_6895,N_6863);
and U7189 (N_7189,N_6938,N_6902);
nor U7190 (N_7190,N_6828,N_6798);
nand U7191 (N_7191,N_6760,N_6999);
nor U7192 (N_7192,N_6812,N_6863);
nor U7193 (N_7193,N_6995,N_6918);
nand U7194 (N_7194,N_6998,N_6773);
nor U7195 (N_7195,N_6992,N_6835);
and U7196 (N_7196,N_6934,N_6878);
or U7197 (N_7197,N_6956,N_6808);
and U7198 (N_7198,N_6918,N_6930);
nand U7199 (N_7199,N_6917,N_6806);
nor U7200 (N_7200,N_6777,N_6965);
nand U7201 (N_7201,N_6772,N_6751);
nor U7202 (N_7202,N_6762,N_6890);
or U7203 (N_7203,N_6894,N_6887);
or U7204 (N_7204,N_6900,N_6996);
nor U7205 (N_7205,N_6964,N_6796);
and U7206 (N_7206,N_6835,N_6917);
nor U7207 (N_7207,N_6937,N_6866);
xnor U7208 (N_7208,N_6927,N_6837);
and U7209 (N_7209,N_6755,N_6859);
and U7210 (N_7210,N_6773,N_6988);
nor U7211 (N_7211,N_6902,N_6995);
or U7212 (N_7212,N_6906,N_6836);
or U7213 (N_7213,N_6813,N_6964);
nand U7214 (N_7214,N_6854,N_6870);
and U7215 (N_7215,N_6796,N_6994);
or U7216 (N_7216,N_6863,N_6839);
nor U7217 (N_7217,N_6958,N_6850);
nor U7218 (N_7218,N_6863,N_6754);
nor U7219 (N_7219,N_6864,N_6980);
nand U7220 (N_7220,N_6751,N_6983);
or U7221 (N_7221,N_6879,N_6788);
xnor U7222 (N_7222,N_6927,N_6770);
nand U7223 (N_7223,N_6756,N_6832);
nand U7224 (N_7224,N_6873,N_6957);
xnor U7225 (N_7225,N_6840,N_6896);
nand U7226 (N_7226,N_6945,N_6915);
or U7227 (N_7227,N_6889,N_6795);
nand U7228 (N_7228,N_6929,N_6920);
or U7229 (N_7229,N_6925,N_6848);
xor U7230 (N_7230,N_6838,N_6861);
xor U7231 (N_7231,N_6799,N_6889);
nand U7232 (N_7232,N_6864,N_6852);
xor U7233 (N_7233,N_6851,N_6827);
xnor U7234 (N_7234,N_6757,N_6776);
or U7235 (N_7235,N_6934,N_6813);
and U7236 (N_7236,N_6996,N_6953);
or U7237 (N_7237,N_6752,N_6785);
nor U7238 (N_7238,N_6814,N_6795);
nor U7239 (N_7239,N_6910,N_6752);
xnor U7240 (N_7240,N_6845,N_6846);
nand U7241 (N_7241,N_6764,N_6921);
nor U7242 (N_7242,N_6827,N_6751);
nor U7243 (N_7243,N_6809,N_6810);
or U7244 (N_7244,N_6977,N_6865);
nand U7245 (N_7245,N_6840,N_6886);
xor U7246 (N_7246,N_6895,N_6974);
or U7247 (N_7247,N_6764,N_6807);
xnor U7248 (N_7248,N_6893,N_6884);
nor U7249 (N_7249,N_6953,N_6961);
nand U7250 (N_7250,N_7194,N_7109);
xnor U7251 (N_7251,N_7073,N_7243);
nand U7252 (N_7252,N_7150,N_7038);
nand U7253 (N_7253,N_7024,N_7209);
or U7254 (N_7254,N_7146,N_7219);
nor U7255 (N_7255,N_7202,N_7106);
xnor U7256 (N_7256,N_7078,N_7061);
nor U7257 (N_7257,N_7077,N_7035);
and U7258 (N_7258,N_7220,N_7081);
nand U7259 (N_7259,N_7021,N_7165);
xnor U7260 (N_7260,N_7010,N_7217);
nand U7261 (N_7261,N_7245,N_7222);
xor U7262 (N_7262,N_7167,N_7029);
xor U7263 (N_7263,N_7231,N_7174);
xnor U7264 (N_7264,N_7225,N_7086);
xor U7265 (N_7265,N_7242,N_7173);
xnor U7266 (N_7266,N_7182,N_7006);
or U7267 (N_7267,N_7208,N_7183);
and U7268 (N_7268,N_7179,N_7026);
nor U7269 (N_7269,N_7060,N_7017);
nand U7270 (N_7270,N_7034,N_7135);
and U7271 (N_7271,N_7158,N_7016);
nor U7272 (N_7272,N_7198,N_7136);
nor U7273 (N_7273,N_7248,N_7049);
xor U7274 (N_7274,N_7129,N_7143);
xor U7275 (N_7275,N_7228,N_7224);
nand U7276 (N_7276,N_7004,N_7237);
and U7277 (N_7277,N_7175,N_7156);
nand U7278 (N_7278,N_7094,N_7070);
nand U7279 (N_7279,N_7047,N_7083);
xor U7280 (N_7280,N_7042,N_7119);
xnor U7281 (N_7281,N_7115,N_7062);
and U7282 (N_7282,N_7051,N_7023);
or U7283 (N_7283,N_7122,N_7171);
or U7284 (N_7284,N_7140,N_7155);
xor U7285 (N_7285,N_7043,N_7090);
and U7286 (N_7286,N_7247,N_7137);
xnor U7287 (N_7287,N_7113,N_7059);
xnor U7288 (N_7288,N_7238,N_7169);
and U7289 (N_7289,N_7056,N_7102);
and U7290 (N_7290,N_7246,N_7069);
or U7291 (N_7291,N_7065,N_7148);
nor U7292 (N_7292,N_7009,N_7221);
and U7293 (N_7293,N_7184,N_7002);
and U7294 (N_7294,N_7000,N_7084);
or U7295 (N_7295,N_7111,N_7011);
xnor U7296 (N_7296,N_7116,N_7160);
or U7297 (N_7297,N_7036,N_7048);
nor U7298 (N_7298,N_7147,N_7040);
and U7299 (N_7299,N_7014,N_7132);
nor U7300 (N_7300,N_7164,N_7152);
and U7301 (N_7301,N_7087,N_7207);
nand U7302 (N_7302,N_7071,N_7190);
nor U7303 (N_7303,N_7188,N_7210);
and U7304 (N_7304,N_7120,N_7142);
xnor U7305 (N_7305,N_7114,N_7153);
or U7306 (N_7306,N_7020,N_7180);
xnor U7307 (N_7307,N_7189,N_7012);
nand U7308 (N_7308,N_7064,N_7118);
nand U7309 (N_7309,N_7052,N_7110);
and U7310 (N_7310,N_7015,N_7008);
nand U7311 (N_7311,N_7177,N_7131);
xor U7312 (N_7312,N_7099,N_7058);
xnor U7313 (N_7313,N_7074,N_7240);
or U7314 (N_7314,N_7244,N_7151);
nand U7315 (N_7315,N_7172,N_7154);
or U7316 (N_7316,N_7204,N_7162);
nor U7317 (N_7317,N_7108,N_7191);
xnor U7318 (N_7318,N_7195,N_7033);
or U7319 (N_7319,N_7125,N_7145);
xnor U7320 (N_7320,N_7057,N_7127);
xnor U7321 (N_7321,N_7100,N_7236);
nand U7322 (N_7322,N_7032,N_7161);
or U7323 (N_7323,N_7185,N_7241);
xor U7324 (N_7324,N_7091,N_7193);
nor U7325 (N_7325,N_7031,N_7067);
or U7326 (N_7326,N_7226,N_7249);
and U7327 (N_7327,N_7170,N_7163);
nor U7328 (N_7328,N_7213,N_7103);
nor U7329 (N_7329,N_7068,N_7149);
nor U7330 (N_7330,N_7117,N_7139);
and U7331 (N_7331,N_7123,N_7128);
and U7332 (N_7332,N_7223,N_7001);
nor U7333 (N_7333,N_7168,N_7230);
xnor U7334 (N_7334,N_7215,N_7214);
xnor U7335 (N_7335,N_7200,N_7133);
nor U7336 (N_7336,N_7075,N_7199);
nand U7337 (N_7337,N_7098,N_7166);
and U7338 (N_7338,N_7003,N_7076);
nor U7339 (N_7339,N_7046,N_7055);
and U7340 (N_7340,N_7196,N_7211);
nor U7341 (N_7341,N_7178,N_7121);
nor U7342 (N_7342,N_7054,N_7203);
and U7343 (N_7343,N_7097,N_7104);
xor U7344 (N_7344,N_7141,N_7050);
or U7345 (N_7345,N_7124,N_7022);
or U7346 (N_7346,N_7159,N_7186);
or U7347 (N_7347,N_7206,N_7039);
nor U7348 (N_7348,N_7095,N_7030);
xnor U7349 (N_7349,N_7085,N_7101);
nor U7350 (N_7350,N_7134,N_7187);
and U7351 (N_7351,N_7176,N_7079);
xor U7352 (N_7352,N_7088,N_7205);
xnor U7353 (N_7353,N_7025,N_7007);
or U7354 (N_7354,N_7092,N_7027);
nand U7355 (N_7355,N_7028,N_7045);
and U7356 (N_7356,N_7044,N_7197);
or U7357 (N_7357,N_7096,N_7234);
nor U7358 (N_7358,N_7089,N_7229);
and U7359 (N_7359,N_7157,N_7235);
nor U7360 (N_7360,N_7105,N_7181);
nand U7361 (N_7361,N_7218,N_7066);
nor U7362 (N_7362,N_7233,N_7232);
and U7363 (N_7363,N_7126,N_7018);
nand U7364 (N_7364,N_7041,N_7192);
or U7365 (N_7365,N_7072,N_7107);
nand U7366 (N_7366,N_7144,N_7005);
and U7367 (N_7367,N_7053,N_7080);
or U7368 (N_7368,N_7201,N_7013);
nor U7369 (N_7369,N_7216,N_7063);
or U7370 (N_7370,N_7037,N_7239);
nor U7371 (N_7371,N_7082,N_7138);
or U7372 (N_7372,N_7112,N_7130);
and U7373 (N_7373,N_7212,N_7227);
and U7374 (N_7374,N_7093,N_7019);
and U7375 (N_7375,N_7165,N_7110);
and U7376 (N_7376,N_7119,N_7050);
nand U7377 (N_7377,N_7069,N_7192);
nor U7378 (N_7378,N_7059,N_7147);
or U7379 (N_7379,N_7020,N_7153);
or U7380 (N_7380,N_7085,N_7033);
and U7381 (N_7381,N_7175,N_7158);
or U7382 (N_7382,N_7108,N_7000);
and U7383 (N_7383,N_7065,N_7127);
xor U7384 (N_7384,N_7034,N_7056);
xor U7385 (N_7385,N_7045,N_7231);
nor U7386 (N_7386,N_7200,N_7217);
and U7387 (N_7387,N_7027,N_7084);
xor U7388 (N_7388,N_7032,N_7003);
or U7389 (N_7389,N_7221,N_7050);
and U7390 (N_7390,N_7224,N_7157);
xnor U7391 (N_7391,N_7174,N_7016);
xnor U7392 (N_7392,N_7030,N_7070);
or U7393 (N_7393,N_7040,N_7004);
nand U7394 (N_7394,N_7152,N_7175);
xor U7395 (N_7395,N_7142,N_7021);
nand U7396 (N_7396,N_7024,N_7121);
xnor U7397 (N_7397,N_7138,N_7108);
nand U7398 (N_7398,N_7083,N_7182);
and U7399 (N_7399,N_7089,N_7151);
nor U7400 (N_7400,N_7028,N_7103);
nor U7401 (N_7401,N_7199,N_7014);
nor U7402 (N_7402,N_7114,N_7071);
and U7403 (N_7403,N_7232,N_7009);
and U7404 (N_7404,N_7196,N_7153);
nand U7405 (N_7405,N_7008,N_7245);
and U7406 (N_7406,N_7010,N_7109);
and U7407 (N_7407,N_7050,N_7067);
xor U7408 (N_7408,N_7192,N_7073);
xnor U7409 (N_7409,N_7139,N_7005);
nand U7410 (N_7410,N_7002,N_7230);
or U7411 (N_7411,N_7085,N_7128);
xnor U7412 (N_7412,N_7172,N_7054);
xnor U7413 (N_7413,N_7242,N_7019);
nor U7414 (N_7414,N_7206,N_7009);
or U7415 (N_7415,N_7044,N_7165);
nand U7416 (N_7416,N_7136,N_7027);
and U7417 (N_7417,N_7080,N_7234);
nand U7418 (N_7418,N_7026,N_7204);
nor U7419 (N_7419,N_7010,N_7175);
and U7420 (N_7420,N_7201,N_7227);
nand U7421 (N_7421,N_7213,N_7117);
xnor U7422 (N_7422,N_7170,N_7082);
nor U7423 (N_7423,N_7181,N_7034);
or U7424 (N_7424,N_7246,N_7081);
xnor U7425 (N_7425,N_7137,N_7147);
and U7426 (N_7426,N_7210,N_7227);
nand U7427 (N_7427,N_7209,N_7139);
nor U7428 (N_7428,N_7151,N_7094);
xor U7429 (N_7429,N_7152,N_7008);
xor U7430 (N_7430,N_7238,N_7154);
nor U7431 (N_7431,N_7126,N_7121);
xnor U7432 (N_7432,N_7217,N_7004);
or U7433 (N_7433,N_7028,N_7095);
nor U7434 (N_7434,N_7093,N_7087);
nand U7435 (N_7435,N_7219,N_7242);
or U7436 (N_7436,N_7089,N_7238);
xor U7437 (N_7437,N_7040,N_7200);
nor U7438 (N_7438,N_7075,N_7036);
nor U7439 (N_7439,N_7077,N_7162);
nand U7440 (N_7440,N_7167,N_7219);
nand U7441 (N_7441,N_7008,N_7237);
xnor U7442 (N_7442,N_7072,N_7133);
and U7443 (N_7443,N_7021,N_7036);
or U7444 (N_7444,N_7134,N_7059);
or U7445 (N_7445,N_7185,N_7097);
and U7446 (N_7446,N_7098,N_7159);
xnor U7447 (N_7447,N_7238,N_7048);
xnor U7448 (N_7448,N_7001,N_7198);
or U7449 (N_7449,N_7205,N_7228);
or U7450 (N_7450,N_7141,N_7075);
or U7451 (N_7451,N_7043,N_7047);
or U7452 (N_7452,N_7152,N_7061);
nand U7453 (N_7453,N_7137,N_7046);
nor U7454 (N_7454,N_7129,N_7239);
or U7455 (N_7455,N_7131,N_7217);
nor U7456 (N_7456,N_7009,N_7241);
or U7457 (N_7457,N_7145,N_7048);
nor U7458 (N_7458,N_7066,N_7247);
nor U7459 (N_7459,N_7204,N_7038);
xor U7460 (N_7460,N_7180,N_7156);
or U7461 (N_7461,N_7172,N_7158);
nor U7462 (N_7462,N_7023,N_7219);
or U7463 (N_7463,N_7113,N_7148);
nor U7464 (N_7464,N_7013,N_7029);
nor U7465 (N_7465,N_7235,N_7125);
or U7466 (N_7466,N_7055,N_7032);
nor U7467 (N_7467,N_7005,N_7199);
and U7468 (N_7468,N_7075,N_7191);
nand U7469 (N_7469,N_7074,N_7225);
nor U7470 (N_7470,N_7102,N_7243);
or U7471 (N_7471,N_7149,N_7159);
nand U7472 (N_7472,N_7223,N_7129);
xnor U7473 (N_7473,N_7236,N_7164);
xnor U7474 (N_7474,N_7118,N_7244);
or U7475 (N_7475,N_7064,N_7031);
nor U7476 (N_7476,N_7067,N_7123);
or U7477 (N_7477,N_7094,N_7012);
nor U7478 (N_7478,N_7218,N_7006);
and U7479 (N_7479,N_7103,N_7186);
nor U7480 (N_7480,N_7021,N_7248);
or U7481 (N_7481,N_7009,N_7104);
xnor U7482 (N_7482,N_7090,N_7246);
xor U7483 (N_7483,N_7183,N_7018);
xnor U7484 (N_7484,N_7057,N_7038);
or U7485 (N_7485,N_7107,N_7043);
or U7486 (N_7486,N_7133,N_7225);
and U7487 (N_7487,N_7230,N_7162);
xnor U7488 (N_7488,N_7104,N_7059);
and U7489 (N_7489,N_7066,N_7025);
or U7490 (N_7490,N_7060,N_7124);
and U7491 (N_7491,N_7048,N_7130);
and U7492 (N_7492,N_7086,N_7194);
and U7493 (N_7493,N_7159,N_7168);
nand U7494 (N_7494,N_7052,N_7122);
and U7495 (N_7495,N_7166,N_7197);
nor U7496 (N_7496,N_7175,N_7177);
and U7497 (N_7497,N_7094,N_7205);
xnor U7498 (N_7498,N_7088,N_7113);
nand U7499 (N_7499,N_7174,N_7104);
or U7500 (N_7500,N_7351,N_7304);
xnor U7501 (N_7501,N_7449,N_7267);
nor U7502 (N_7502,N_7281,N_7260);
nand U7503 (N_7503,N_7377,N_7400);
or U7504 (N_7504,N_7468,N_7479);
xnor U7505 (N_7505,N_7321,N_7290);
nor U7506 (N_7506,N_7424,N_7346);
or U7507 (N_7507,N_7431,N_7356);
xnor U7508 (N_7508,N_7336,N_7358);
xnor U7509 (N_7509,N_7385,N_7367);
nand U7510 (N_7510,N_7444,N_7443);
or U7511 (N_7511,N_7323,N_7275);
nand U7512 (N_7512,N_7492,N_7446);
and U7513 (N_7513,N_7481,N_7314);
or U7514 (N_7514,N_7438,N_7398);
xor U7515 (N_7515,N_7308,N_7452);
nor U7516 (N_7516,N_7470,N_7369);
nor U7517 (N_7517,N_7456,N_7319);
nand U7518 (N_7518,N_7399,N_7343);
and U7519 (N_7519,N_7416,N_7422);
and U7520 (N_7520,N_7317,N_7407);
and U7521 (N_7521,N_7439,N_7373);
nand U7522 (N_7522,N_7276,N_7262);
and U7523 (N_7523,N_7279,N_7383);
or U7524 (N_7524,N_7345,N_7331);
nor U7525 (N_7525,N_7355,N_7394);
xnor U7526 (N_7526,N_7261,N_7310);
and U7527 (N_7527,N_7389,N_7427);
nand U7528 (N_7528,N_7469,N_7381);
nand U7529 (N_7529,N_7418,N_7288);
nor U7530 (N_7530,N_7357,N_7359);
xor U7531 (N_7531,N_7423,N_7312);
nor U7532 (N_7532,N_7485,N_7437);
or U7533 (N_7533,N_7445,N_7412);
nor U7534 (N_7534,N_7284,N_7337);
nand U7535 (N_7535,N_7305,N_7382);
xnor U7536 (N_7536,N_7297,N_7387);
nand U7537 (N_7537,N_7482,N_7498);
and U7538 (N_7538,N_7453,N_7316);
nand U7539 (N_7539,N_7436,N_7303);
or U7540 (N_7540,N_7366,N_7473);
or U7541 (N_7541,N_7402,N_7397);
nor U7542 (N_7542,N_7268,N_7360);
or U7543 (N_7543,N_7464,N_7457);
nor U7544 (N_7544,N_7461,N_7497);
and U7545 (N_7545,N_7392,N_7333);
xor U7546 (N_7546,N_7306,N_7440);
nor U7547 (N_7547,N_7368,N_7463);
or U7548 (N_7548,N_7415,N_7301);
xnor U7549 (N_7549,N_7414,N_7480);
and U7550 (N_7550,N_7488,N_7264);
or U7551 (N_7551,N_7477,N_7256);
nor U7552 (N_7552,N_7471,N_7362);
or U7553 (N_7553,N_7250,N_7393);
and U7554 (N_7554,N_7404,N_7315);
and U7555 (N_7555,N_7434,N_7348);
xor U7556 (N_7556,N_7287,N_7350);
nand U7557 (N_7557,N_7325,N_7465);
nand U7558 (N_7558,N_7409,N_7390);
nor U7559 (N_7559,N_7257,N_7340);
xnor U7560 (N_7560,N_7411,N_7293);
xnor U7561 (N_7561,N_7354,N_7442);
nand U7562 (N_7562,N_7255,N_7253);
and U7563 (N_7563,N_7380,N_7349);
nor U7564 (N_7564,N_7493,N_7455);
xnor U7565 (N_7565,N_7483,N_7417);
xnor U7566 (N_7566,N_7426,N_7298);
xor U7567 (N_7567,N_7272,N_7296);
nor U7568 (N_7568,N_7344,N_7467);
and U7569 (N_7569,N_7313,N_7274);
nor U7570 (N_7570,N_7347,N_7252);
xor U7571 (N_7571,N_7406,N_7302);
nand U7572 (N_7572,N_7273,N_7484);
and U7573 (N_7573,N_7489,N_7283);
xnor U7574 (N_7574,N_7289,N_7263);
nor U7575 (N_7575,N_7459,N_7277);
and U7576 (N_7576,N_7490,N_7478);
or U7577 (N_7577,N_7282,N_7254);
and U7578 (N_7578,N_7462,N_7420);
or U7579 (N_7579,N_7408,N_7458);
xor U7580 (N_7580,N_7460,N_7454);
nor U7581 (N_7581,N_7396,N_7428);
or U7582 (N_7582,N_7403,N_7370);
and U7583 (N_7583,N_7496,N_7330);
or U7584 (N_7584,N_7342,N_7421);
xor U7585 (N_7585,N_7259,N_7425);
and U7586 (N_7586,N_7395,N_7410);
nand U7587 (N_7587,N_7378,N_7365);
nand U7588 (N_7588,N_7413,N_7332);
or U7589 (N_7589,N_7363,N_7472);
xnor U7590 (N_7590,N_7375,N_7430);
nand U7591 (N_7591,N_7324,N_7328);
nand U7592 (N_7592,N_7476,N_7309);
xor U7593 (N_7593,N_7429,N_7352);
and U7594 (N_7594,N_7361,N_7487);
nand U7595 (N_7595,N_7335,N_7278);
or U7596 (N_7596,N_7300,N_7294);
xor U7597 (N_7597,N_7339,N_7447);
and U7598 (N_7598,N_7286,N_7491);
nor U7599 (N_7599,N_7499,N_7269);
nand U7600 (N_7600,N_7405,N_7384);
xnor U7601 (N_7601,N_7388,N_7280);
xnor U7602 (N_7602,N_7320,N_7386);
and U7603 (N_7603,N_7353,N_7475);
nor U7604 (N_7604,N_7329,N_7435);
xor U7605 (N_7605,N_7372,N_7401);
or U7606 (N_7606,N_7326,N_7334);
and U7607 (N_7607,N_7295,N_7251);
nor U7608 (N_7608,N_7450,N_7338);
xnor U7609 (N_7609,N_7311,N_7270);
or U7610 (N_7610,N_7292,N_7374);
and U7611 (N_7611,N_7474,N_7391);
and U7612 (N_7612,N_7495,N_7307);
xor U7613 (N_7613,N_7466,N_7486);
or U7614 (N_7614,N_7364,N_7258);
xor U7615 (N_7615,N_7271,N_7285);
nor U7616 (N_7616,N_7432,N_7419);
nor U7617 (N_7617,N_7448,N_7371);
nor U7618 (N_7618,N_7441,N_7451);
and U7619 (N_7619,N_7494,N_7322);
and U7620 (N_7620,N_7291,N_7266);
nor U7621 (N_7621,N_7379,N_7341);
nand U7622 (N_7622,N_7327,N_7376);
and U7623 (N_7623,N_7265,N_7318);
nand U7624 (N_7624,N_7299,N_7433);
and U7625 (N_7625,N_7360,N_7342);
or U7626 (N_7626,N_7488,N_7292);
and U7627 (N_7627,N_7289,N_7285);
and U7628 (N_7628,N_7430,N_7428);
xor U7629 (N_7629,N_7330,N_7395);
nand U7630 (N_7630,N_7499,N_7458);
or U7631 (N_7631,N_7257,N_7480);
or U7632 (N_7632,N_7386,N_7406);
and U7633 (N_7633,N_7375,N_7318);
nor U7634 (N_7634,N_7449,N_7361);
nand U7635 (N_7635,N_7271,N_7378);
nor U7636 (N_7636,N_7487,N_7390);
and U7637 (N_7637,N_7459,N_7334);
nor U7638 (N_7638,N_7357,N_7321);
nand U7639 (N_7639,N_7284,N_7467);
or U7640 (N_7640,N_7284,N_7323);
nand U7641 (N_7641,N_7310,N_7313);
nand U7642 (N_7642,N_7399,N_7337);
and U7643 (N_7643,N_7484,N_7491);
nand U7644 (N_7644,N_7367,N_7337);
nor U7645 (N_7645,N_7322,N_7254);
xor U7646 (N_7646,N_7294,N_7250);
nand U7647 (N_7647,N_7433,N_7422);
and U7648 (N_7648,N_7365,N_7474);
or U7649 (N_7649,N_7421,N_7388);
and U7650 (N_7650,N_7272,N_7367);
nand U7651 (N_7651,N_7491,N_7328);
and U7652 (N_7652,N_7409,N_7417);
or U7653 (N_7653,N_7471,N_7405);
and U7654 (N_7654,N_7409,N_7275);
xnor U7655 (N_7655,N_7279,N_7328);
xor U7656 (N_7656,N_7354,N_7341);
nand U7657 (N_7657,N_7470,N_7253);
xnor U7658 (N_7658,N_7320,N_7441);
nor U7659 (N_7659,N_7494,N_7457);
nand U7660 (N_7660,N_7436,N_7484);
or U7661 (N_7661,N_7490,N_7443);
nor U7662 (N_7662,N_7283,N_7435);
or U7663 (N_7663,N_7415,N_7382);
nand U7664 (N_7664,N_7346,N_7437);
or U7665 (N_7665,N_7357,N_7469);
nand U7666 (N_7666,N_7487,N_7333);
xnor U7667 (N_7667,N_7314,N_7427);
or U7668 (N_7668,N_7435,N_7431);
xnor U7669 (N_7669,N_7359,N_7326);
xnor U7670 (N_7670,N_7402,N_7480);
and U7671 (N_7671,N_7328,N_7291);
nand U7672 (N_7672,N_7295,N_7305);
and U7673 (N_7673,N_7376,N_7364);
or U7674 (N_7674,N_7389,N_7378);
xor U7675 (N_7675,N_7397,N_7319);
xor U7676 (N_7676,N_7429,N_7268);
or U7677 (N_7677,N_7362,N_7292);
or U7678 (N_7678,N_7341,N_7287);
nor U7679 (N_7679,N_7338,N_7314);
nor U7680 (N_7680,N_7459,N_7473);
nor U7681 (N_7681,N_7250,N_7470);
xor U7682 (N_7682,N_7474,N_7347);
nor U7683 (N_7683,N_7450,N_7332);
nor U7684 (N_7684,N_7380,N_7264);
and U7685 (N_7685,N_7484,N_7489);
or U7686 (N_7686,N_7395,N_7348);
xnor U7687 (N_7687,N_7271,N_7375);
nor U7688 (N_7688,N_7349,N_7396);
nor U7689 (N_7689,N_7353,N_7267);
xor U7690 (N_7690,N_7458,N_7288);
nand U7691 (N_7691,N_7276,N_7365);
or U7692 (N_7692,N_7387,N_7459);
xnor U7693 (N_7693,N_7317,N_7318);
nor U7694 (N_7694,N_7400,N_7390);
or U7695 (N_7695,N_7277,N_7260);
nor U7696 (N_7696,N_7404,N_7485);
and U7697 (N_7697,N_7353,N_7459);
nor U7698 (N_7698,N_7385,N_7481);
nand U7699 (N_7699,N_7283,N_7436);
nor U7700 (N_7700,N_7467,N_7482);
and U7701 (N_7701,N_7360,N_7408);
nor U7702 (N_7702,N_7448,N_7336);
xor U7703 (N_7703,N_7403,N_7445);
nand U7704 (N_7704,N_7413,N_7292);
or U7705 (N_7705,N_7384,N_7458);
and U7706 (N_7706,N_7461,N_7474);
nor U7707 (N_7707,N_7250,N_7391);
nand U7708 (N_7708,N_7340,N_7319);
nand U7709 (N_7709,N_7302,N_7305);
and U7710 (N_7710,N_7362,N_7364);
nand U7711 (N_7711,N_7474,N_7422);
or U7712 (N_7712,N_7356,N_7324);
or U7713 (N_7713,N_7374,N_7376);
nor U7714 (N_7714,N_7392,N_7336);
and U7715 (N_7715,N_7332,N_7256);
nor U7716 (N_7716,N_7475,N_7357);
or U7717 (N_7717,N_7420,N_7413);
xnor U7718 (N_7718,N_7326,N_7494);
or U7719 (N_7719,N_7329,N_7358);
nand U7720 (N_7720,N_7349,N_7405);
nand U7721 (N_7721,N_7253,N_7481);
or U7722 (N_7722,N_7352,N_7293);
nand U7723 (N_7723,N_7418,N_7410);
xnor U7724 (N_7724,N_7479,N_7365);
and U7725 (N_7725,N_7463,N_7320);
or U7726 (N_7726,N_7336,N_7489);
xor U7727 (N_7727,N_7494,N_7458);
nor U7728 (N_7728,N_7301,N_7353);
and U7729 (N_7729,N_7252,N_7306);
nand U7730 (N_7730,N_7257,N_7315);
nor U7731 (N_7731,N_7286,N_7415);
nand U7732 (N_7732,N_7433,N_7285);
and U7733 (N_7733,N_7496,N_7449);
nor U7734 (N_7734,N_7414,N_7306);
nor U7735 (N_7735,N_7381,N_7402);
or U7736 (N_7736,N_7386,N_7352);
nand U7737 (N_7737,N_7320,N_7269);
and U7738 (N_7738,N_7386,N_7361);
xnor U7739 (N_7739,N_7285,N_7345);
nor U7740 (N_7740,N_7377,N_7451);
xor U7741 (N_7741,N_7493,N_7288);
and U7742 (N_7742,N_7372,N_7289);
nand U7743 (N_7743,N_7362,N_7355);
nand U7744 (N_7744,N_7301,N_7444);
nand U7745 (N_7745,N_7259,N_7403);
xor U7746 (N_7746,N_7281,N_7348);
and U7747 (N_7747,N_7366,N_7418);
and U7748 (N_7748,N_7454,N_7393);
nor U7749 (N_7749,N_7402,N_7466);
or U7750 (N_7750,N_7543,N_7554);
xor U7751 (N_7751,N_7591,N_7620);
and U7752 (N_7752,N_7691,N_7606);
or U7753 (N_7753,N_7626,N_7612);
nor U7754 (N_7754,N_7646,N_7516);
or U7755 (N_7755,N_7537,N_7529);
nor U7756 (N_7756,N_7611,N_7693);
and U7757 (N_7757,N_7631,N_7512);
nor U7758 (N_7758,N_7643,N_7619);
nor U7759 (N_7759,N_7561,N_7695);
and U7760 (N_7760,N_7617,N_7656);
xor U7761 (N_7761,N_7724,N_7578);
nor U7762 (N_7762,N_7501,N_7649);
nor U7763 (N_7763,N_7660,N_7652);
xnor U7764 (N_7764,N_7655,N_7719);
nand U7765 (N_7765,N_7678,N_7671);
nand U7766 (N_7766,N_7599,N_7514);
or U7767 (N_7767,N_7734,N_7544);
or U7768 (N_7768,N_7579,N_7566);
or U7769 (N_7769,N_7613,N_7745);
and U7770 (N_7770,N_7594,N_7665);
xnor U7771 (N_7771,N_7739,N_7556);
xor U7772 (N_7772,N_7707,N_7712);
xnor U7773 (N_7773,N_7698,N_7571);
xnor U7774 (N_7774,N_7681,N_7670);
xor U7775 (N_7775,N_7720,N_7662);
or U7776 (N_7776,N_7568,N_7511);
nor U7777 (N_7777,N_7634,N_7639);
nor U7778 (N_7778,N_7565,N_7697);
xnor U7779 (N_7779,N_7675,N_7551);
and U7780 (N_7780,N_7597,N_7685);
nor U7781 (N_7781,N_7540,N_7558);
nand U7782 (N_7782,N_7648,N_7641);
xor U7783 (N_7783,N_7608,N_7650);
nor U7784 (N_7784,N_7531,N_7555);
or U7785 (N_7785,N_7673,N_7583);
xnor U7786 (N_7786,N_7593,N_7500);
and U7787 (N_7787,N_7716,N_7689);
and U7788 (N_7788,N_7528,N_7694);
nand U7789 (N_7789,N_7687,N_7533);
and U7790 (N_7790,N_7517,N_7709);
nand U7791 (N_7791,N_7515,N_7507);
nand U7792 (N_7792,N_7723,N_7651);
and U7793 (N_7793,N_7610,N_7557);
nor U7794 (N_7794,N_7627,N_7600);
nor U7795 (N_7795,N_7504,N_7667);
nand U7796 (N_7796,N_7732,N_7576);
or U7797 (N_7797,N_7588,N_7744);
nand U7798 (N_7798,N_7527,N_7736);
nand U7799 (N_7799,N_7553,N_7690);
nand U7800 (N_7800,N_7748,N_7635);
nor U7801 (N_7801,N_7521,N_7563);
and U7802 (N_7802,N_7539,N_7609);
or U7803 (N_7803,N_7513,N_7622);
and U7804 (N_7804,N_7721,N_7562);
nor U7805 (N_7805,N_7630,N_7711);
or U7806 (N_7806,N_7573,N_7523);
xor U7807 (N_7807,N_7705,N_7672);
nor U7808 (N_7808,N_7522,N_7542);
and U7809 (N_7809,N_7726,N_7710);
xor U7810 (N_7810,N_7519,N_7725);
nor U7811 (N_7811,N_7584,N_7598);
nor U7812 (N_7812,N_7666,N_7676);
xnor U7813 (N_7813,N_7536,N_7728);
and U7814 (N_7814,N_7580,N_7601);
nand U7815 (N_7815,N_7526,N_7592);
or U7816 (N_7816,N_7505,N_7577);
xor U7817 (N_7817,N_7605,N_7743);
nor U7818 (N_7818,N_7625,N_7741);
xnor U7819 (N_7819,N_7653,N_7548);
nor U7820 (N_7820,N_7703,N_7682);
and U7821 (N_7821,N_7549,N_7683);
nand U7822 (N_7822,N_7589,N_7629);
nand U7823 (N_7823,N_7602,N_7623);
or U7824 (N_7824,N_7607,N_7510);
nand U7825 (N_7825,N_7679,N_7704);
nand U7826 (N_7826,N_7596,N_7647);
xor U7827 (N_7827,N_7664,N_7508);
xor U7828 (N_7828,N_7506,N_7686);
and U7829 (N_7829,N_7737,N_7644);
and U7830 (N_7830,N_7636,N_7530);
or U7831 (N_7831,N_7525,N_7552);
nand U7832 (N_7832,N_7654,N_7722);
and U7833 (N_7833,N_7518,N_7642);
nor U7834 (N_7834,N_7603,N_7714);
nor U7835 (N_7835,N_7702,N_7633);
nor U7836 (N_7836,N_7560,N_7718);
nor U7837 (N_7837,N_7546,N_7582);
xnor U7838 (N_7838,N_7632,N_7669);
nor U7839 (N_7839,N_7564,N_7740);
xor U7840 (N_7840,N_7715,N_7535);
xor U7841 (N_7841,N_7735,N_7708);
nor U7842 (N_7842,N_7746,N_7574);
and U7843 (N_7843,N_7731,N_7729);
or U7844 (N_7844,N_7659,N_7706);
or U7845 (N_7845,N_7677,N_7700);
and U7846 (N_7846,N_7645,N_7585);
nand U7847 (N_7847,N_7587,N_7658);
nor U7848 (N_7848,N_7680,N_7575);
or U7849 (N_7849,N_7604,N_7668);
and U7850 (N_7850,N_7713,N_7699);
nor U7851 (N_7851,N_7738,N_7595);
or U7852 (N_7852,N_7688,N_7616);
or U7853 (N_7853,N_7503,N_7663);
xnor U7854 (N_7854,N_7717,N_7640);
xnor U7855 (N_7855,N_7572,N_7545);
nand U7856 (N_7856,N_7524,N_7661);
nor U7857 (N_7857,N_7590,N_7569);
and U7858 (N_7858,N_7509,N_7701);
and U7859 (N_7859,N_7538,N_7674);
xor U7860 (N_7860,N_7520,N_7727);
xor U7861 (N_7861,N_7749,N_7638);
nand U7862 (N_7862,N_7696,N_7618);
nor U7863 (N_7863,N_7624,N_7747);
nor U7864 (N_7864,N_7733,N_7657);
xnor U7865 (N_7865,N_7570,N_7550);
or U7866 (N_7866,N_7541,N_7614);
and U7867 (N_7867,N_7730,N_7684);
and U7868 (N_7868,N_7502,N_7547);
or U7869 (N_7869,N_7637,N_7586);
xnor U7870 (N_7870,N_7692,N_7532);
and U7871 (N_7871,N_7534,N_7567);
and U7872 (N_7872,N_7621,N_7742);
nor U7873 (N_7873,N_7559,N_7581);
or U7874 (N_7874,N_7615,N_7628);
or U7875 (N_7875,N_7627,N_7740);
nor U7876 (N_7876,N_7721,N_7651);
and U7877 (N_7877,N_7692,N_7659);
nand U7878 (N_7878,N_7666,N_7609);
nor U7879 (N_7879,N_7726,N_7622);
or U7880 (N_7880,N_7644,N_7594);
nand U7881 (N_7881,N_7537,N_7633);
and U7882 (N_7882,N_7617,N_7503);
nor U7883 (N_7883,N_7706,N_7515);
nor U7884 (N_7884,N_7702,N_7634);
xor U7885 (N_7885,N_7630,N_7683);
or U7886 (N_7886,N_7650,N_7665);
or U7887 (N_7887,N_7722,N_7625);
nand U7888 (N_7888,N_7745,N_7562);
or U7889 (N_7889,N_7559,N_7685);
or U7890 (N_7890,N_7503,N_7724);
nand U7891 (N_7891,N_7747,N_7701);
xnor U7892 (N_7892,N_7693,N_7591);
or U7893 (N_7893,N_7701,N_7630);
nand U7894 (N_7894,N_7573,N_7684);
or U7895 (N_7895,N_7644,N_7525);
nor U7896 (N_7896,N_7620,N_7677);
nand U7897 (N_7897,N_7686,N_7626);
and U7898 (N_7898,N_7585,N_7702);
or U7899 (N_7899,N_7644,N_7562);
nor U7900 (N_7900,N_7520,N_7730);
nand U7901 (N_7901,N_7710,N_7528);
nor U7902 (N_7902,N_7684,N_7571);
nand U7903 (N_7903,N_7604,N_7659);
or U7904 (N_7904,N_7629,N_7728);
nor U7905 (N_7905,N_7705,N_7719);
nor U7906 (N_7906,N_7597,N_7580);
nor U7907 (N_7907,N_7522,N_7666);
xnor U7908 (N_7908,N_7504,N_7627);
and U7909 (N_7909,N_7612,N_7641);
nor U7910 (N_7910,N_7676,N_7716);
nand U7911 (N_7911,N_7549,N_7547);
xnor U7912 (N_7912,N_7641,N_7568);
xor U7913 (N_7913,N_7571,N_7664);
nor U7914 (N_7914,N_7537,N_7712);
nand U7915 (N_7915,N_7529,N_7601);
xor U7916 (N_7916,N_7745,N_7634);
or U7917 (N_7917,N_7702,N_7531);
or U7918 (N_7918,N_7555,N_7678);
or U7919 (N_7919,N_7575,N_7559);
xor U7920 (N_7920,N_7639,N_7509);
and U7921 (N_7921,N_7601,N_7700);
nand U7922 (N_7922,N_7676,N_7719);
or U7923 (N_7923,N_7621,N_7610);
or U7924 (N_7924,N_7627,N_7649);
nor U7925 (N_7925,N_7610,N_7640);
or U7926 (N_7926,N_7719,N_7570);
nand U7927 (N_7927,N_7615,N_7712);
and U7928 (N_7928,N_7720,N_7633);
and U7929 (N_7929,N_7678,N_7562);
or U7930 (N_7930,N_7636,N_7614);
or U7931 (N_7931,N_7687,N_7685);
nor U7932 (N_7932,N_7733,N_7559);
or U7933 (N_7933,N_7508,N_7691);
xnor U7934 (N_7934,N_7619,N_7573);
and U7935 (N_7935,N_7646,N_7628);
xnor U7936 (N_7936,N_7695,N_7686);
xnor U7937 (N_7937,N_7617,N_7584);
nand U7938 (N_7938,N_7733,N_7615);
nor U7939 (N_7939,N_7564,N_7586);
nand U7940 (N_7940,N_7578,N_7587);
and U7941 (N_7941,N_7648,N_7620);
nor U7942 (N_7942,N_7619,N_7508);
or U7943 (N_7943,N_7553,N_7566);
nand U7944 (N_7944,N_7524,N_7526);
or U7945 (N_7945,N_7665,N_7680);
xnor U7946 (N_7946,N_7692,N_7620);
nor U7947 (N_7947,N_7562,N_7583);
xor U7948 (N_7948,N_7543,N_7510);
nor U7949 (N_7949,N_7566,N_7625);
nand U7950 (N_7950,N_7511,N_7746);
xnor U7951 (N_7951,N_7688,N_7721);
nor U7952 (N_7952,N_7520,N_7504);
nand U7953 (N_7953,N_7749,N_7651);
nor U7954 (N_7954,N_7637,N_7669);
or U7955 (N_7955,N_7639,N_7541);
xnor U7956 (N_7956,N_7632,N_7746);
and U7957 (N_7957,N_7685,N_7623);
xor U7958 (N_7958,N_7547,N_7703);
and U7959 (N_7959,N_7746,N_7559);
xnor U7960 (N_7960,N_7733,N_7661);
nor U7961 (N_7961,N_7663,N_7657);
and U7962 (N_7962,N_7652,N_7662);
or U7963 (N_7963,N_7712,N_7658);
nand U7964 (N_7964,N_7681,N_7620);
or U7965 (N_7965,N_7502,N_7696);
or U7966 (N_7966,N_7609,N_7743);
or U7967 (N_7967,N_7685,N_7689);
and U7968 (N_7968,N_7558,N_7604);
nand U7969 (N_7969,N_7515,N_7558);
nor U7970 (N_7970,N_7512,N_7567);
and U7971 (N_7971,N_7735,N_7690);
nor U7972 (N_7972,N_7520,N_7585);
nand U7973 (N_7973,N_7504,N_7546);
and U7974 (N_7974,N_7655,N_7511);
xor U7975 (N_7975,N_7577,N_7631);
and U7976 (N_7976,N_7515,N_7701);
nand U7977 (N_7977,N_7739,N_7679);
or U7978 (N_7978,N_7546,N_7609);
nor U7979 (N_7979,N_7632,N_7630);
xnor U7980 (N_7980,N_7638,N_7720);
nand U7981 (N_7981,N_7651,N_7617);
or U7982 (N_7982,N_7589,N_7538);
nand U7983 (N_7983,N_7565,N_7616);
or U7984 (N_7984,N_7637,N_7660);
xor U7985 (N_7985,N_7652,N_7618);
or U7986 (N_7986,N_7593,N_7586);
and U7987 (N_7987,N_7687,N_7503);
nor U7988 (N_7988,N_7699,N_7663);
and U7989 (N_7989,N_7653,N_7606);
xor U7990 (N_7990,N_7690,N_7585);
and U7991 (N_7991,N_7597,N_7541);
or U7992 (N_7992,N_7565,N_7507);
nor U7993 (N_7993,N_7630,N_7731);
nor U7994 (N_7994,N_7580,N_7723);
nor U7995 (N_7995,N_7584,N_7532);
nor U7996 (N_7996,N_7720,N_7714);
and U7997 (N_7997,N_7657,N_7647);
nand U7998 (N_7998,N_7742,N_7603);
nor U7999 (N_7999,N_7670,N_7525);
or U8000 (N_8000,N_7975,N_7883);
nand U8001 (N_8001,N_7982,N_7934);
xor U8002 (N_8002,N_7859,N_7953);
nor U8003 (N_8003,N_7796,N_7889);
nor U8004 (N_8004,N_7983,N_7904);
nand U8005 (N_8005,N_7961,N_7948);
xor U8006 (N_8006,N_7924,N_7808);
xnor U8007 (N_8007,N_7930,N_7978);
or U8008 (N_8008,N_7853,N_7907);
nor U8009 (N_8009,N_7903,N_7751);
nand U8010 (N_8010,N_7995,N_7988);
and U8011 (N_8011,N_7922,N_7756);
nor U8012 (N_8012,N_7985,N_7831);
and U8013 (N_8013,N_7974,N_7803);
and U8014 (N_8014,N_7750,N_7816);
and U8015 (N_8015,N_7917,N_7856);
nor U8016 (N_8016,N_7954,N_7980);
and U8017 (N_8017,N_7900,N_7827);
nand U8018 (N_8018,N_7817,N_7840);
or U8019 (N_8019,N_7802,N_7825);
nor U8020 (N_8020,N_7806,N_7902);
and U8021 (N_8021,N_7931,N_7855);
nor U8022 (N_8022,N_7848,N_7767);
nor U8023 (N_8023,N_7863,N_7788);
and U8024 (N_8024,N_7836,N_7925);
nor U8025 (N_8025,N_7832,N_7870);
nor U8026 (N_8026,N_7947,N_7968);
or U8027 (N_8027,N_7764,N_7799);
nand U8028 (N_8028,N_7795,N_7896);
nor U8029 (N_8029,N_7850,N_7981);
nand U8030 (N_8030,N_7857,N_7775);
and U8031 (N_8031,N_7997,N_7837);
nand U8032 (N_8032,N_7769,N_7885);
or U8033 (N_8033,N_7994,N_7842);
and U8034 (N_8034,N_7854,N_7860);
nand U8035 (N_8035,N_7835,N_7793);
nand U8036 (N_8036,N_7819,N_7834);
nand U8037 (N_8037,N_7916,N_7770);
nor U8038 (N_8038,N_7960,N_7880);
nand U8039 (N_8039,N_7933,N_7919);
nor U8040 (N_8040,N_7888,N_7754);
or U8041 (N_8041,N_7768,N_7787);
or U8042 (N_8042,N_7959,N_7777);
nand U8043 (N_8043,N_7923,N_7914);
nand U8044 (N_8044,N_7879,N_7890);
and U8045 (N_8045,N_7846,N_7894);
and U8046 (N_8046,N_7755,N_7752);
or U8047 (N_8047,N_7887,N_7818);
nand U8048 (N_8048,N_7895,N_7958);
and U8049 (N_8049,N_7881,N_7811);
and U8050 (N_8050,N_7866,N_7809);
nand U8051 (N_8051,N_7784,N_7949);
nor U8052 (N_8052,N_7946,N_7969);
or U8053 (N_8053,N_7973,N_7876);
xnor U8054 (N_8054,N_7971,N_7812);
nor U8055 (N_8055,N_7794,N_7776);
xor U8056 (N_8056,N_7822,N_7805);
xor U8057 (N_8057,N_7841,N_7972);
nand U8058 (N_8058,N_7852,N_7929);
and U8059 (N_8059,N_7928,N_7965);
nor U8060 (N_8060,N_7875,N_7936);
nand U8061 (N_8061,N_7804,N_7989);
xor U8062 (N_8062,N_7810,N_7792);
and U8063 (N_8063,N_7814,N_7830);
or U8064 (N_8064,N_7785,N_7932);
nor U8065 (N_8065,N_7865,N_7938);
xnor U8066 (N_8066,N_7905,N_7992);
and U8067 (N_8067,N_7868,N_7780);
and U8068 (N_8068,N_7843,N_7911);
nand U8069 (N_8069,N_7807,N_7999);
nand U8070 (N_8070,N_7912,N_7847);
or U8071 (N_8071,N_7952,N_7998);
nor U8072 (N_8072,N_7829,N_7790);
and U8073 (N_8073,N_7991,N_7763);
and U8074 (N_8074,N_7765,N_7979);
nor U8075 (N_8075,N_7976,N_7970);
nor U8076 (N_8076,N_7845,N_7906);
nor U8077 (N_8077,N_7977,N_7753);
and U8078 (N_8078,N_7964,N_7800);
nand U8079 (N_8079,N_7984,N_7955);
nand U8080 (N_8080,N_7833,N_7872);
nand U8081 (N_8081,N_7851,N_7801);
and U8082 (N_8082,N_7838,N_7918);
or U8083 (N_8083,N_7908,N_7878);
xor U8084 (N_8084,N_7937,N_7781);
xnor U8085 (N_8085,N_7966,N_7824);
or U8086 (N_8086,N_7874,N_7759);
and U8087 (N_8087,N_7957,N_7791);
xnor U8088 (N_8088,N_7993,N_7987);
xnor U8089 (N_8089,N_7913,N_7901);
xor U8090 (N_8090,N_7951,N_7963);
nor U8091 (N_8091,N_7921,N_7813);
nor U8092 (N_8092,N_7864,N_7886);
and U8093 (N_8093,N_7909,N_7990);
and U8094 (N_8094,N_7892,N_7897);
or U8095 (N_8095,N_7943,N_7967);
nor U8096 (N_8096,N_7826,N_7772);
or U8097 (N_8097,N_7761,N_7915);
or U8098 (N_8098,N_7873,N_7821);
or U8099 (N_8099,N_7839,N_7944);
or U8100 (N_8100,N_7789,N_7758);
xor U8101 (N_8101,N_7844,N_7786);
or U8102 (N_8102,N_7757,N_7815);
or U8103 (N_8103,N_7871,N_7762);
and U8104 (N_8104,N_7773,N_7950);
nand U8105 (N_8105,N_7771,N_7783);
xor U8106 (N_8106,N_7861,N_7862);
and U8107 (N_8107,N_7935,N_7899);
or U8108 (N_8108,N_7941,N_7766);
nor U8109 (N_8109,N_7774,N_7823);
nand U8110 (N_8110,N_7849,N_7858);
xor U8111 (N_8111,N_7778,N_7986);
and U8112 (N_8112,N_7882,N_7869);
xnor U8113 (N_8113,N_7867,N_7779);
and U8114 (N_8114,N_7891,N_7942);
or U8115 (N_8115,N_7760,N_7782);
xnor U8116 (N_8116,N_7797,N_7884);
and U8117 (N_8117,N_7939,N_7910);
or U8118 (N_8118,N_7945,N_7927);
nor U8119 (N_8119,N_7828,N_7920);
or U8120 (N_8120,N_7956,N_7877);
nor U8121 (N_8121,N_7940,N_7820);
xnor U8122 (N_8122,N_7893,N_7996);
or U8123 (N_8123,N_7898,N_7962);
and U8124 (N_8124,N_7926,N_7798);
xor U8125 (N_8125,N_7910,N_7800);
xor U8126 (N_8126,N_7915,N_7754);
xnor U8127 (N_8127,N_7874,N_7903);
xnor U8128 (N_8128,N_7872,N_7984);
nand U8129 (N_8129,N_7862,N_7856);
xor U8130 (N_8130,N_7826,N_7900);
nor U8131 (N_8131,N_7992,N_7803);
nor U8132 (N_8132,N_7767,N_7863);
nand U8133 (N_8133,N_7992,N_7993);
or U8134 (N_8134,N_7913,N_7868);
and U8135 (N_8135,N_7908,N_7885);
nand U8136 (N_8136,N_7812,N_7798);
and U8137 (N_8137,N_7932,N_7778);
xor U8138 (N_8138,N_7923,N_7789);
nor U8139 (N_8139,N_7829,N_7774);
or U8140 (N_8140,N_7904,N_7885);
xor U8141 (N_8141,N_7801,N_7934);
and U8142 (N_8142,N_7942,N_7790);
nor U8143 (N_8143,N_7911,N_7930);
xor U8144 (N_8144,N_7916,N_7812);
nand U8145 (N_8145,N_7924,N_7912);
xor U8146 (N_8146,N_7991,N_7861);
xnor U8147 (N_8147,N_7781,N_7839);
xor U8148 (N_8148,N_7870,N_7820);
and U8149 (N_8149,N_7806,N_7861);
or U8150 (N_8150,N_7863,N_7881);
nor U8151 (N_8151,N_7967,N_7817);
nor U8152 (N_8152,N_7806,N_7766);
xnor U8153 (N_8153,N_7966,N_7944);
and U8154 (N_8154,N_7941,N_7839);
or U8155 (N_8155,N_7900,N_7772);
or U8156 (N_8156,N_7820,N_7793);
and U8157 (N_8157,N_7981,N_7886);
and U8158 (N_8158,N_7841,N_7760);
xnor U8159 (N_8159,N_7968,N_7774);
and U8160 (N_8160,N_7979,N_7849);
or U8161 (N_8161,N_7968,N_7984);
and U8162 (N_8162,N_7826,N_7762);
nand U8163 (N_8163,N_7888,N_7853);
nor U8164 (N_8164,N_7980,N_7882);
xor U8165 (N_8165,N_7793,N_7869);
nand U8166 (N_8166,N_7857,N_7791);
or U8167 (N_8167,N_7997,N_7868);
nand U8168 (N_8168,N_7760,N_7946);
nand U8169 (N_8169,N_7892,N_7775);
or U8170 (N_8170,N_7793,N_7890);
nand U8171 (N_8171,N_7937,N_7938);
or U8172 (N_8172,N_7880,N_7779);
nand U8173 (N_8173,N_7890,N_7763);
nand U8174 (N_8174,N_7938,N_7836);
nor U8175 (N_8175,N_7893,N_7812);
nor U8176 (N_8176,N_7818,N_7871);
nand U8177 (N_8177,N_7890,N_7991);
or U8178 (N_8178,N_7980,N_7952);
nand U8179 (N_8179,N_7769,N_7826);
or U8180 (N_8180,N_7762,N_7933);
or U8181 (N_8181,N_7831,N_7780);
xnor U8182 (N_8182,N_7867,N_7822);
nor U8183 (N_8183,N_7920,N_7995);
nor U8184 (N_8184,N_7778,N_7923);
and U8185 (N_8185,N_7883,N_7908);
nand U8186 (N_8186,N_7878,N_7994);
and U8187 (N_8187,N_7842,N_7878);
and U8188 (N_8188,N_7923,N_7961);
or U8189 (N_8189,N_7818,N_7767);
nand U8190 (N_8190,N_7939,N_7925);
xor U8191 (N_8191,N_7823,N_7794);
nand U8192 (N_8192,N_7838,N_7793);
and U8193 (N_8193,N_7845,N_7955);
nor U8194 (N_8194,N_7860,N_7878);
or U8195 (N_8195,N_7896,N_7858);
xor U8196 (N_8196,N_7780,N_7922);
nor U8197 (N_8197,N_7819,N_7970);
or U8198 (N_8198,N_7771,N_7791);
xnor U8199 (N_8199,N_7872,N_7795);
or U8200 (N_8200,N_7778,N_7922);
xnor U8201 (N_8201,N_7853,N_7979);
nor U8202 (N_8202,N_7890,N_7765);
and U8203 (N_8203,N_7935,N_7922);
nor U8204 (N_8204,N_7768,N_7750);
and U8205 (N_8205,N_7984,N_7924);
nor U8206 (N_8206,N_7841,N_7856);
nand U8207 (N_8207,N_7987,N_7967);
nand U8208 (N_8208,N_7781,N_7962);
nor U8209 (N_8209,N_7993,N_7864);
nor U8210 (N_8210,N_7750,N_7838);
and U8211 (N_8211,N_7772,N_7882);
nor U8212 (N_8212,N_7854,N_7961);
or U8213 (N_8213,N_7965,N_7832);
nand U8214 (N_8214,N_7979,N_7781);
xnor U8215 (N_8215,N_7750,N_7803);
and U8216 (N_8216,N_7756,N_7971);
nand U8217 (N_8217,N_7979,N_7942);
xor U8218 (N_8218,N_7756,N_7996);
nand U8219 (N_8219,N_7803,N_7885);
nand U8220 (N_8220,N_7781,N_7759);
xor U8221 (N_8221,N_7857,N_7774);
and U8222 (N_8222,N_7997,N_7933);
or U8223 (N_8223,N_7764,N_7785);
xor U8224 (N_8224,N_7966,N_7876);
and U8225 (N_8225,N_7809,N_7900);
nand U8226 (N_8226,N_7929,N_7916);
and U8227 (N_8227,N_7773,N_7822);
and U8228 (N_8228,N_7951,N_7884);
and U8229 (N_8229,N_7778,N_7935);
or U8230 (N_8230,N_7787,N_7851);
nor U8231 (N_8231,N_7802,N_7960);
or U8232 (N_8232,N_7823,N_7868);
or U8233 (N_8233,N_7960,N_7817);
or U8234 (N_8234,N_7852,N_7811);
and U8235 (N_8235,N_7977,N_7787);
or U8236 (N_8236,N_7966,N_7960);
and U8237 (N_8237,N_7908,N_7750);
or U8238 (N_8238,N_7781,N_7919);
nand U8239 (N_8239,N_7961,N_7797);
or U8240 (N_8240,N_7754,N_7974);
nand U8241 (N_8241,N_7928,N_7937);
nand U8242 (N_8242,N_7767,N_7823);
nand U8243 (N_8243,N_7922,N_7959);
nor U8244 (N_8244,N_7931,N_7939);
and U8245 (N_8245,N_7832,N_7758);
nor U8246 (N_8246,N_7901,N_7805);
and U8247 (N_8247,N_7958,N_7961);
nand U8248 (N_8248,N_7833,N_7923);
nand U8249 (N_8249,N_7972,N_7893);
or U8250 (N_8250,N_8068,N_8205);
xor U8251 (N_8251,N_8038,N_8184);
or U8252 (N_8252,N_8082,N_8008);
nand U8253 (N_8253,N_8227,N_8210);
xnor U8254 (N_8254,N_8037,N_8125);
nand U8255 (N_8255,N_8151,N_8059);
nand U8256 (N_8256,N_8232,N_8192);
xor U8257 (N_8257,N_8017,N_8236);
xnor U8258 (N_8258,N_8161,N_8188);
and U8259 (N_8259,N_8035,N_8076);
nand U8260 (N_8260,N_8063,N_8244);
xor U8261 (N_8261,N_8090,N_8182);
nand U8262 (N_8262,N_8052,N_8087);
or U8263 (N_8263,N_8123,N_8055);
nand U8264 (N_8264,N_8166,N_8116);
nor U8265 (N_8265,N_8200,N_8249);
nand U8266 (N_8266,N_8095,N_8217);
and U8267 (N_8267,N_8067,N_8136);
nor U8268 (N_8268,N_8191,N_8100);
or U8269 (N_8269,N_8211,N_8153);
nor U8270 (N_8270,N_8208,N_8004);
nand U8271 (N_8271,N_8084,N_8110);
xnor U8272 (N_8272,N_8083,N_8107);
xor U8273 (N_8273,N_8178,N_8108);
nor U8274 (N_8274,N_8189,N_8117);
or U8275 (N_8275,N_8235,N_8047);
xor U8276 (N_8276,N_8088,N_8114);
xor U8277 (N_8277,N_8193,N_8034);
or U8278 (N_8278,N_8143,N_8072);
nand U8279 (N_8279,N_8077,N_8203);
nor U8280 (N_8280,N_8027,N_8020);
nor U8281 (N_8281,N_8156,N_8011);
nor U8282 (N_8282,N_8199,N_8176);
xnor U8283 (N_8283,N_8025,N_8238);
nor U8284 (N_8284,N_8006,N_8229);
and U8285 (N_8285,N_8042,N_8183);
or U8286 (N_8286,N_8225,N_8054);
xor U8287 (N_8287,N_8111,N_8045);
nor U8288 (N_8288,N_8102,N_8165);
or U8289 (N_8289,N_8133,N_8194);
nor U8290 (N_8290,N_8022,N_8150);
and U8291 (N_8291,N_8096,N_8186);
and U8292 (N_8292,N_8215,N_8226);
and U8293 (N_8293,N_8170,N_8075);
nand U8294 (N_8294,N_8169,N_8009);
xor U8295 (N_8295,N_8132,N_8240);
or U8296 (N_8296,N_8162,N_8173);
or U8297 (N_8297,N_8030,N_8222);
and U8298 (N_8298,N_8098,N_8018);
or U8299 (N_8299,N_8003,N_8180);
xor U8300 (N_8300,N_8148,N_8119);
xor U8301 (N_8301,N_8080,N_8130);
xor U8302 (N_8302,N_8032,N_8239);
xnor U8303 (N_8303,N_8033,N_8139);
nand U8304 (N_8304,N_8050,N_8079);
xnor U8305 (N_8305,N_8056,N_8127);
nand U8306 (N_8306,N_8094,N_8066);
xnor U8307 (N_8307,N_8069,N_8041);
nand U8308 (N_8308,N_8154,N_8099);
and U8309 (N_8309,N_8010,N_8073);
xor U8310 (N_8310,N_8112,N_8046);
or U8311 (N_8311,N_8219,N_8204);
nand U8312 (N_8312,N_8048,N_8036);
nor U8313 (N_8313,N_8230,N_8168);
nand U8314 (N_8314,N_8146,N_8134);
nor U8315 (N_8315,N_8214,N_8051);
nor U8316 (N_8316,N_8163,N_8092);
or U8317 (N_8317,N_8206,N_8109);
nor U8318 (N_8318,N_8044,N_8086);
and U8319 (N_8319,N_8040,N_8081);
or U8320 (N_8320,N_8216,N_8196);
nand U8321 (N_8321,N_8197,N_8005);
xor U8322 (N_8322,N_8031,N_8089);
and U8323 (N_8323,N_8071,N_8091);
and U8324 (N_8324,N_8135,N_8223);
xnor U8325 (N_8325,N_8187,N_8124);
nor U8326 (N_8326,N_8190,N_8157);
and U8327 (N_8327,N_8179,N_8198);
xnor U8328 (N_8328,N_8118,N_8172);
xor U8329 (N_8329,N_8175,N_8002);
and U8330 (N_8330,N_8158,N_8149);
xor U8331 (N_8331,N_8233,N_8057);
xor U8332 (N_8332,N_8106,N_8012);
or U8333 (N_8333,N_8185,N_8144);
nor U8334 (N_8334,N_8015,N_8128);
xnor U8335 (N_8335,N_8028,N_8171);
and U8336 (N_8336,N_8122,N_8085);
or U8337 (N_8337,N_8142,N_8220);
nor U8338 (N_8338,N_8065,N_8248);
and U8339 (N_8339,N_8016,N_8007);
and U8340 (N_8340,N_8078,N_8234);
xor U8341 (N_8341,N_8202,N_8247);
and U8342 (N_8342,N_8039,N_8074);
or U8343 (N_8343,N_8213,N_8137);
nor U8344 (N_8344,N_8145,N_8029);
xor U8345 (N_8345,N_8201,N_8121);
xor U8346 (N_8346,N_8101,N_8043);
and U8347 (N_8347,N_8070,N_8242);
nand U8348 (N_8348,N_8026,N_8152);
or U8349 (N_8349,N_8228,N_8062);
and U8350 (N_8350,N_8231,N_8140);
or U8351 (N_8351,N_8113,N_8115);
nand U8352 (N_8352,N_8049,N_8221);
nor U8353 (N_8353,N_8060,N_8064);
and U8354 (N_8354,N_8021,N_8129);
nand U8355 (N_8355,N_8131,N_8181);
xor U8356 (N_8356,N_8105,N_8023);
nand U8357 (N_8357,N_8155,N_8243);
nor U8358 (N_8358,N_8174,N_8218);
nand U8359 (N_8359,N_8159,N_8103);
xor U8360 (N_8360,N_8000,N_8120);
nand U8361 (N_8361,N_8093,N_8212);
and U8362 (N_8362,N_8246,N_8177);
nor U8363 (N_8363,N_8224,N_8058);
and U8364 (N_8364,N_8126,N_8104);
nor U8365 (N_8365,N_8160,N_8207);
or U8366 (N_8366,N_8014,N_8237);
nand U8367 (N_8367,N_8001,N_8061);
nor U8368 (N_8368,N_8141,N_8245);
or U8369 (N_8369,N_8241,N_8019);
xor U8370 (N_8370,N_8147,N_8013);
and U8371 (N_8371,N_8209,N_8097);
and U8372 (N_8372,N_8167,N_8164);
and U8373 (N_8373,N_8024,N_8053);
nor U8374 (N_8374,N_8138,N_8195);
or U8375 (N_8375,N_8052,N_8249);
or U8376 (N_8376,N_8040,N_8146);
nor U8377 (N_8377,N_8004,N_8046);
xor U8378 (N_8378,N_8002,N_8016);
nor U8379 (N_8379,N_8044,N_8021);
nand U8380 (N_8380,N_8048,N_8081);
or U8381 (N_8381,N_8180,N_8210);
xor U8382 (N_8382,N_8001,N_8164);
nor U8383 (N_8383,N_8054,N_8223);
and U8384 (N_8384,N_8201,N_8143);
xor U8385 (N_8385,N_8215,N_8125);
xnor U8386 (N_8386,N_8101,N_8049);
or U8387 (N_8387,N_8057,N_8066);
and U8388 (N_8388,N_8148,N_8206);
and U8389 (N_8389,N_8011,N_8049);
or U8390 (N_8390,N_8063,N_8131);
xor U8391 (N_8391,N_8047,N_8223);
and U8392 (N_8392,N_8132,N_8004);
nand U8393 (N_8393,N_8091,N_8026);
nand U8394 (N_8394,N_8172,N_8230);
nand U8395 (N_8395,N_8012,N_8218);
xnor U8396 (N_8396,N_8144,N_8181);
and U8397 (N_8397,N_8156,N_8176);
nor U8398 (N_8398,N_8235,N_8046);
xor U8399 (N_8399,N_8113,N_8178);
and U8400 (N_8400,N_8013,N_8200);
and U8401 (N_8401,N_8006,N_8067);
nand U8402 (N_8402,N_8173,N_8159);
or U8403 (N_8403,N_8093,N_8086);
nand U8404 (N_8404,N_8130,N_8068);
or U8405 (N_8405,N_8070,N_8041);
nor U8406 (N_8406,N_8101,N_8058);
or U8407 (N_8407,N_8221,N_8096);
or U8408 (N_8408,N_8094,N_8038);
or U8409 (N_8409,N_8167,N_8045);
nor U8410 (N_8410,N_8182,N_8154);
nand U8411 (N_8411,N_8219,N_8009);
nor U8412 (N_8412,N_8098,N_8218);
and U8413 (N_8413,N_8169,N_8039);
nand U8414 (N_8414,N_8217,N_8192);
or U8415 (N_8415,N_8049,N_8139);
and U8416 (N_8416,N_8113,N_8021);
nor U8417 (N_8417,N_8096,N_8138);
or U8418 (N_8418,N_8025,N_8071);
nor U8419 (N_8419,N_8203,N_8107);
nand U8420 (N_8420,N_8140,N_8115);
nand U8421 (N_8421,N_8015,N_8126);
nand U8422 (N_8422,N_8162,N_8050);
xnor U8423 (N_8423,N_8130,N_8196);
nand U8424 (N_8424,N_8118,N_8094);
nand U8425 (N_8425,N_8188,N_8210);
and U8426 (N_8426,N_8087,N_8088);
and U8427 (N_8427,N_8240,N_8114);
and U8428 (N_8428,N_8044,N_8005);
or U8429 (N_8429,N_8245,N_8160);
or U8430 (N_8430,N_8200,N_8230);
nand U8431 (N_8431,N_8058,N_8223);
nand U8432 (N_8432,N_8077,N_8048);
and U8433 (N_8433,N_8124,N_8099);
nand U8434 (N_8434,N_8151,N_8243);
nor U8435 (N_8435,N_8120,N_8110);
and U8436 (N_8436,N_8047,N_8129);
nand U8437 (N_8437,N_8079,N_8247);
xnor U8438 (N_8438,N_8119,N_8153);
and U8439 (N_8439,N_8037,N_8063);
nand U8440 (N_8440,N_8135,N_8226);
nor U8441 (N_8441,N_8010,N_8031);
or U8442 (N_8442,N_8080,N_8234);
nor U8443 (N_8443,N_8095,N_8045);
xnor U8444 (N_8444,N_8183,N_8049);
or U8445 (N_8445,N_8028,N_8085);
xnor U8446 (N_8446,N_8014,N_8063);
and U8447 (N_8447,N_8063,N_8111);
xnor U8448 (N_8448,N_8059,N_8208);
nand U8449 (N_8449,N_8169,N_8182);
nand U8450 (N_8450,N_8003,N_8002);
nand U8451 (N_8451,N_8113,N_8041);
nand U8452 (N_8452,N_8106,N_8168);
nand U8453 (N_8453,N_8047,N_8177);
nor U8454 (N_8454,N_8160,N_8120);
xnor U8455 (N_8455,N_8133,N_8075);
nand U8456 (N_8456,N_8102,N_8039);
nand U8457 (N_8457,N_8035,N_8140);
xnor U8458 (N_8458,N_8076,N_8071);
nor U8459 (N_8459,N_8062,N_8095);
xor U8460 (N_8460,N_8204,N_8147);
and U8461 (N_8461,N_8179,N_8108);
xnor U8462 (N_8462,N_8211,N_8049);
and U8463 (N_8463,N_8125,N_8123);
or U8464 (N_8464,N_8176,N_8027);
and U8465 (N_8465,N_8138,N_8199);
and U8466 (N_8466,N_8005,N_8056);
or U8467 (N_8467,N_8246,N_8197);
and U8468 (N_8468,N_8191,N_8110);
xor U8469 (N_8469,N_8191,N_8016);
and U8470 (N_8470,N_8228,N_8065);
and U8471 (N_8471,N_8232,N_8055);
nor U8472 (N_8472,N_8092,N_8054);
nor U8473 (N_8473,N_8097,N_8045);
nand U8474 (N_8474,N_8101,N_8105);
nand U8475 (N_8475,N_8218,N_8066);
and U8476 (N_8476,N_8089,N_8173);
or U8477 (N_8477,N_8155,N_8131);
xor U8478 (N_8478,N_8206,N_8158);
xnor U8479 (N_8479,N_8133,N_8174);
and U8480 (N_8480,N_8159,N_8248);
xnor U8481 (N_8481,N_8101,N_8002);
or U8482 (N_8482,N_8076,N_8110);
or U8483 (N_8483,N_8209,N_8085);
nor U8484 (N_8484,N_8005,N_8181);
nand U8485 (N_8485,N_8015,N_8145);
and U8486 (N_8486,N_8063,N_8059);
nor U8487 (N_8487,N_8053,N_8184);
and U8488 (N_8488,N_8117,N_8181);
and U8489 (N_8489,N_8120,N_8118);
xor U8490 (N_8490,N_8095,N_8100);
xnor U8491 (N_8491,N_8078,N_8210);
and U8492 (N_8492,N_8237,N_8077);
nand U8493 (N_8493,N_8143,N_8150);
or U8494 (N_8494,N_8121,N_8025);
or U8495 (N_8495,N_8058,N_8019);
nand U8496 (N_8496,N_8003,N_8207);
and U8497 (N_8497,N_8157,N_8208);
and U8498 (N_8498,N_8168,N_8191);
and U8499 (N_8499,N_8122,N_8191);
or U8500 (N_8500,N_8311,N_8472);
nand U8501 (N_8501,N_8361,N_8368);
or U8502 (N_8502,N_8348,N_8497);
nor U8503 (N_8503,N_8438,N_8336);
and U8504 (N_8504,N_8355,N_8376);
or U8505 (N_8505,N_8261,N_8269);
xnor U8506 (N_8506,N_8495,N_8468);
xnor U8507 (N_8507,N_8260,N_8447);
xnor U8508 (N_8508,N_8475,N_8334);
and U8509 (N_8509,N_8403,N_8317);
nor U8510 (N_8510,N_8288,N_8357);
and U8511 (N_8511,N_8346,N_8349);
or U8512 (N_8512,N_8370,N_8411);
nor U8513 (N_8513,N_8335,N_8390);
nand U8514 (N_8514,N_8496,N_8362);
and U8515 (N_8515,N_8427,N_8476);
nor U8516 (N_8516,N_8479,N_8493);
nand U8517 (N_8517,N_8270,N_8391);
nor U8518 (N_8518,N_8379,N_8259);
nand U8519 (N_8519,N_8393,N_8275);
xor U8520 (N_8520,N_8340,N_8462);
and U8521 (N_8521,N_8324,N_8265);
or U8522 (N_8522,N_8449,N_8486);
nand U8523 (N_8523,N_8441,N_8463);
or U8524 (N_8524,N_8351,N_8416);
nor U8525 (N_8525,N_8281,N_8380);
and U8526 (N_8526,N_8284,N_8296);
xor U8527 (N_8527,N_8470,N_8482);
nor U8528 (N_8528,N_8375,N_8268);
and U8529 (N_8529,N_8429,N_8484);
xnor U8530 (N_8530,N_8322,N_8446);
xor U8531 (N_8531,N_8253,N_8258);
and U8532 (N_8532,N_8491,N_8251);
xnor U8533 (N_8533,N_8323,N_8325);
nor U8534 (N_8534,N_8352,N_8499);
xor U8535 (N_8535,N_8272,N_8452);
xor U8536 (N_8536,N_8444,N_8287);
and U8537 (N_8537,N_8386,N_8487);
or U8538 (N_8538,N_8293,N_8459);
or U8539 (N_8539,N_8423,N_8289);
and U8540 (N_8540,N_8435,N_8458);
nor U8541 (N_8541,N_8399,N_8400);
nor U8542 (N_8542,N_8409,N_8356);
nand U8543 (N_8543,N_8398,N_8347);
nand U8544 (N_8544,N_8433,N_8498);
xnor U8545 (N_8545,N_8342,N_8267);
or U8546 (N_8546,N_8273,N_8254);
or U8547 (N_8547,N_8358,N_8445);
xnor U8548 (N_8548,N_8305,N_8374);
xnor U8549 (N_8549,N_8408,N_8350);
xnor U8550 (N_8550,N_8461,N_8315);
nor U8551 (N_8551,N_8250,N_8426);
or U8552 (N_8552,N_8405,N_8274);
nand U8553 (N_8553,N_8453,N_8443);
and U8554 (N_8554,N_8363,N_8313);
and U8555 (N_8555,N_8366,N_8279);
nand U8556 (N_8556,N_8280,N_8304);
nand U8557 (N_8557,N_8301,N_8292);
nor U8558 (N_8558,N_8488,N_8377);
nor U8559 (N_8559,N_8300,N_8432);
nand U8560 (N_8560,N_8417,N_8478);
xnor U8561 (N_8561,N_8307,N_8381);
or U8562 (N_8562,N_8407,N_8339);
nand U8563 (N_8563,N_8252,N_8312);
nor U8564 (N_8564,N_8450,N_8460);
nor U8565 (N_8565,N_8457,N_8278);
nand U8566 (N_8566,N_8303,N_8483);
xor U8567 (N_8567,N_8285,N_8420);
nor U8568 (N_8568,N_8337,N_8473);
nand U8569 (N_8569,N_8302,N_8321);
nand U8570 (N_8570,N_8290,N_8294);
xnor U8571 (N_8571,N_8434,N_8286);
nand U8572 (N_8572,N_8451,N_8365);
nand U8573 (N_8573,N_8424,N_8343);
and U8574 (N_8574,N_8422,N_8419);
and U8575 (N_8575,N_8466,N_8320);
and U8576 (N_8576,N_8364,N_8277);
nor U8577 (N_8577,N_8298,N_8257);
xnor U8578 (N_8578,N_8421,N_8314);
nor U8579 (N_8579,N_8338,N_8359);
nand U8580 (N_8580,N_8430,N_8297);
nor U8581 (N_8581,N_8266,N_8382);
nand U8582 (N_8582,N_8369,N_8282);
nor U8583 (N_8583,N_8326,N_8480);
or U8584 (N_8584,N_8471,N_8437);
or U8585 (N_8585,N_8360,N_8394);
or U8586 (N_8586,N_8436,N_8474);
or U8587 (N_8587,N_8308,N_8481);
or U8588 (N_8588,N_8378,N_8395);
nor U8589 (N_8589,N_8413,N_8271);
nor U8590 (N_8590,N_8319,N_8384);
xnor U8591 (N_8591,N_8344,N_8494);
nand U8592 (N_8592,N_8329,N_8341);
nor U8593 (N_8593,N_8389,N_8306);
and U8594 (N_8594,N_8283,N_8397);
nor U8595 (N_8595,N_8410,N_8402);
nor U8596 (N_8596,N_8477,N_8372);
and U8597 (N_8597,N_8418,N_8454);
xor U8598 (N_8598,N_8412,N_8440);
and U8599 (N_8599,N_8464,N_8295);
nor U8600 (N_8600,N_8256,N_8490);
and U8601 (N_8601,N_8262,N_8327);
nor U8602 (N_8602,N_8425,N_8263);
xor U8603 (N_8603,N_8309,N_8333);
or U8604 (N_8604,N_8439,N_8310);
nor U8605 (N_8605,N_8367,N_8388);
xnor U8606 (N_8606,N_8392,N_8492);
or U8607 (N_8607,N_8489,N_8371);
nand U8608 (N_8608,N_8414,N_8401);
or U8609 (N_8609,N_8387,N_8331);
nand U8610 (N_8610,N_8316,N_8291);
nand U8611 (N_8611,N_8442,N_8406);
nand U8612 (N_8612,N_8448,N_8345);
xnor U8613 (N_8613,N_8255,N_8385);
nor U8614 (N_8614,N_8383,N_8332);
nor U8615 (N_8615,N_8276,N_8465);
nor U8616 (N_8616,N_8318,N_8455);
and U8617 (N_8617,N_8396,N_8428);
nand U8618 (N_8618,N_8469,N_8456);
and U8619 (N_8619,N_8485,N_8353);
and U8620 (N_8620,N_8431,N_8415);
xnor U8621 (N_8621,N_8404,N_8330);
nand U8622 (N_8622,N_8264,N_8328);
xnor U8623 (N_8623,N_8467,N_8373);
or U8624 (N_8624,N_8354,N_8299);
nand U8625 (N_8625,N_8250,N_8414);
or U8626 (N_8626,N_8260,N_8485);
xnor U8627 (N_8627,N_8369,N_8332);
nor U8628 (N_8628,N_8491,N_8492);
or U8629 (N_8629,N_8356,N_8463);
nor U8630 (N_8630,N_8273,N_8297);
nor U8631 (N_8631,N_8275,N_8382);
nand U8632 (N_8632,N_8455,N_8399);
and U8633 (N_8633,N_8449,N_8393);
xnor U8634 (N_8634,N_8492,N_8302);
or U8635 (N_8635,N_8344,N_8464);
nand U8636 (N_8636,N_8356,N_8419);
and U8637 (N_8637,N_8335,N_8407);
xnor U8638 (N_8638,N_8434,N_8432);
nand U8639 (N_8639,N_8395,N_8480);
nand U8640 (N_8640,N_8478,N_8269);
xor U8641 (N_8641,N_8451,N_8469);
or U8642 (N_8642,N_8292,N_8321);
nor U8643 (N_8643,N_8490,N_8290);
xor U8644 (N_8644,N_8373,N_8256);
nand U8645 (N_8645,N_8288,N_8287);
or U8646 (N_8646,N_8383,N_8308);
nor U8647 (N_8647,N_8356,N_8289);
nand U8648 (N_8648,N_8356,N_8426);
and U8649 (N_8649,N_8323,N_8488);
nand U8650 (N_8650,N_8295,N_8268);
nand U8651 (N_8651,N_8441,N_8383);
and U8652 (N_8652,N_8354,N_8423);
xnor U8653 (N_8653,N_8306,N_8291);
nor U8654 (N_8654,N_8486,N_8331);
xnor U8655 (N_8655,N_8377,N_8342);
nor U8656 (N_8656,N_8427,N_8370);
nand U8657 (N_8657,N_8413,N_8289);
and U8658 (N_8658,N_8354,N_8335);
nand U8659 (N_8659,N_8480,N_8458);
and U8660 (N_8660,N_8451,N_8395);
and U8661 (N_8661,N_8265,N_8253);
nor U8662 (N_8662,N_8312,N_8338);
nor U8663 (N_8663,N_8353,N_8339);
or U8664 (N_8664,N_8442,N_8483);
nand U8665 (N_8665,N_8359,N_8345);
and U8666 (N_8666,N_8310,N_8411);
nand U8667 (N_8667,N_8487,N_8362);
nand U8668 (N_8668,N_8426,N_8447);
nand U8669 (N_8669,N_8257,N_8310);
xnor U8670 (N_8670,N_8464,N_8477);
nand U8671 (N_8671,N_8416,N_8426);
and U8672 (N_8672,N_8474,N_8255);
and U8673 (N_8673,N_8486,N_8419);
nand U8674 (N_8674,N_8301,N_8272);
or U8675 (N_8675,N_8304,N_8449);
nor U8676 (N_8676,N_8292,N_8257);
nand U8677 (N_8677,N_8443,N_8416);
and U8678 (N_8678,N_8433,N_8336);
xnor U8679 (N_8679,N_8371,N_8488);
and U8680 (N_8680,N_8267,N_8335);
nand U8681 (N_8681,N_8367,N_8349);
or U8682 (N_8682,N_8457,N_8413);
or U8683 (N_8683,N_8317,N_8481);
or U8684 (N_8684,N_8469,N_8382);
and U8685 (N_8685,N_8290,N_8406);
or U8686 (N_8686,N_8445,N_8304);
and U8687 (N_8687,N_8487,N_8393);
nor U8688 (N_8688,N_8299,N_8305);
nor U8689 (N_8689,N_8360,N_8480);
and U8690 (N_8690,N_8386,N_8353);
nor U8691 (N_8691,N_8464,N_8490);
xnor U8692 (N_8692,N_8280,N_8467);
nand U8693 (N_8693,N_8464,N_8461);
nor U8694 (N_8694,N_8413,N_8459);
nor U8695 (N_8695,N_8319,N_8387);
xor U8696 (N_8696,N_8269,N_8329);
nor U8697 (N_8697,N_8342,N_8432);
or U8698 (N_8698,N_8285,N_8313);
nor U8699 (N_8699,N_8255,N_8426);
and U8700 (N_8700,N_8437,N_8411);
or U8701 (N_8701,N_8427,N_8369);
nor U8702 (N_8702,N_8450,N_8262);
or U8703 (N_8703,N_8250,N_8422);
xnor U8704 (N_8704,N_8449,N_8342);
nor U8705 (N_8705,N_8278,N_8318);
xor U8706 (N_8706,N_8344,N_8396);
and U8707 (N_8707,N_8336,N_8424);
nand U8708 (N_8708,N_8321,N_8384);
nor U8709 (N_8709,N_8275,N_8469);
xnor U8710 (N_8710,N_8388,N_8324);
xor U8711 (N_8711,N_8265,N_8282);
xnor U8712 (N_8712,N_8404,N_8250);
nor U8713 (N_8713,N_8344,N_8381);
or U8714 (N_8714,N_8475,N_8482);
nor U8715 (N_8715,N_8283,N_8435);
nor U8716 (N_8716,N_8390,N_8487);
xnor U8717 (N_8717,N_8261,N_8256);
xor U8718 (N_8718,N_8344,N_8293);
nor U8719 (N_8719,N_8339,N_8341);
xnor U8720 (N_8720,N_8359,N_8326);
or U8721 (N_8721,N_8260,N_8444);
xor U8722 (N_8722,N_8317,N_8459);
and U8723 (N_8723,N_8387,N_8346);
nor U8724 (N_8724,N_8448,N_8467);
xnor U8725 (N_8725,N_8349,N_8347);
nor U8726 (N_8726,N_8432,N_8303);
and U8727 (N_8727,N_8423,N_8401);
or U8728 (N_8728,N_8337,N_8270);
xor U8729 (N_8729,N_8286,N_8469);
nor U8730 (N_8730,N_8403,N_8416);
nand U8731 (N_8731,N_8305,N_8458);
nor U8732 (N_8732,N_8497,N_8464);
or U8733 (N_8733,N_8435,N_8300);
xor U8734 (N_8734,N_8476,N_8455);
nor U8735 (N_8735,N_8450,N_8285);
and U8736 (N_8736,N_8318,N_8325);
or U8737 (N_8737,N_8375,N_8434);
or U8738 (N_8738,N_8342,N_8410);
xor U8739 (N_8739,N_8267,N_8303);
xor U8740 (N_8740,N_8441,N_8302);
and U8741 (N_8741,N_8294,N_8471);
and U8742 (N_8742,N_8353,N_8298);
xnor U8743 (N_8743,N_8425,N_8255);
and U8744 (N_8744,N_8348,N_8266);
and U8745 (N_8745,N_8489,N_8289);
and U8746 (N_8746,N_8443,N_8434);
nand U8747 (N_8747,N_8381,N_8406);
nand U8748 (N_8748,N_8437,N_8455);
and U8749 (N_8749,N_8420,N_8357);
nand U8750 (N_8750,N_8618,N_8683);
xnor U8751 (N_8751,N_8603,N_8673);
nor U8752 (N_8752,N_8616,N_8652);
or U8753 (N_8753,N_8634,N_8645);
or U8754 (N_8754,N_8522,N_8680);
and U8755 (N_8755,N_8587,N_8504);
nand U8756 (N_8756,N_8614,N_8611);
nor U8757 (N_8757,N_8586,N_8651);
nor U8758 (N_8758,N_8664,N_8696);
xnor U8759 (N_8759,N_8501,N_8737);
and U8760 (N_8760,N_8707,N_8677);
and U8761 (N_8761,N_8745,N_8602);
and U8762 (N_8762,N_8719,N_8689);
or U8763 (N_8763,N_8594,N_8559);
or U8764 (N_8764,N_8716,N_8609);
nand U8765 (N_8765,N_8549,N_8531);
nor U8766 (N_8766,N_8655,N_8599);
xnor U8767 (N_8767,N_8600,N_8523);
nor U8768 (N_8768,N_8511,N_8682);
and U8769 (N_8769,N_8540,N_8686);
and U8770 (N_8770,N_8519,N_8663);
nand U8771 (N_8771,N_8667,N_8713);
and U8772 (N_8772,N_8721,N_8518);
or U8773 (N_8773,N_8733,N_8581);
or U8774 (N_8774,N_8562,N_8650);
nor U8775 (N_8775,N_8711,N_8544);
or U8776 (N_8776,N_8654,N_8592);
xor U8777 (N_8777,N_8644,N_8700);
nand U8778 (N_8778,N_8672,N_8658);
nand U8779 (N_8779,N_8708,N_8515);
and U8780 (N_8780,N_8695,N_8573);
and U8781 (N_8781,N_8625,N_8726);
xnor U8782 (N_8782,N_8640,N_8722);
or U8783 (N_8783,N_8607,N_8589);
and U8784 (N_8784,N_8500,N_8653);
nand U8785 (N_8785,N_8521,N_8546);
xnor U8786 (N_8786,N_8665,N_8636);
xnor U8787 (N_8787,N_8561,N_8570);
xor U8788 (N_8788,N_8508,N_8572);
and U8789 (N_8789,N_8661,N_8660);
nor U8790 (N_8790,N_8533,N_8510);
nor U8791 (N_8791,N_8670,N_8738);
nor U8792 (N_8792,N_8718,N_8622);
nand U8793 (N_8793,N_8662,N_8605);
xor U8794 (N_8794,N_8554,N_8729);
or U8795 (N_8795,N_8727,N_8701);
xnor U8796 (N_8796,N_8598,N_8527);
nand U8797 (N_8797,N_8740,N_8582);
xor U8798 (N_8798,N_8747,N_8637);
xor U8799 (N_8799,N_8687,N_8635);
nor U8800 (N_8800,N_8743,N_8617);
and U8801 (N_8801,N_8615,N_8731);
or U8802 (N_8802,N_8741,N_8671);
nand U8803 (N_8803,N_8608,N_8541);
nand U8804 (N_8804,N_8529,N_8704);
or U8805 (N_8805,N_8593,N_8612);
nand U8806 (N_8806,N_8633,N_8623);
nand U8807 (N_8807,N_8698,N_8706);
and U8808 (N_8808,N_8628,N_8624);
and U8809 (N_8809,N_8532,N_8565);
or U8810 (N_8810,N_8555,N_8517);
or U8811 (N_8811,N_8638,N_8703);
xnor U8812 (N_8812,N_8601,N_8712);
and U8813 (N_8813,N_8674,N_8639);
and U8814 (N_8814,N_8621,N_8569);
nor U8815 (N_8815,N_8563,N_8659);
and U8816 (N_8816,N_8685,N_8530);
and U8817 (N_8817,N_8606,N_8724);
or U8818 (N_8818,N_8643,N_8545);
xor U8819 (N_8819,N_8619,N_8723);
nand U8820 (N_8820,N_8583,N_8710);
or U8821 (N_8821,N_8749,N_8604);
and U8822 (N_8822,N_8736,N_8692);
nor U8823 (N_8823,N_8613,N_8668);
and U8824 (N_8824,N_8728,N_8746);
nand U8825 (N_8825,N_8505,N_8675);
and U8826 (N_8826,N_8502,N_8538);
and U8827 (N_8827,N_8526,N_8597);
nand U8828 (N_8828,N_8647,N_8678);
or U8829 (N_8829,N_8566,N_8735);
nand U8830 (N_8830,N_8536,N_8543);
xor U8831 (N_8831,N_8577,N_8720);
and U8832 (N_8832,N_8620,N_8676);
nor U8833 (N_8833,N_8730,N_8535);
nand U8834 (N_8834,N_8688,N_8699);
and U8835 (N_8835,N_8509,N_8595);
nand U8836 (N_8836,N_8702,N_8550);
nor U8837 (N_8837,N_8556,N_8553);
or U8838 (N_8838,N_8537,N_8630);
or U8839 (N_8839,N_8524,N_8631);
or U8840 (N_8840,N_8714,N_8507);
or U8841 (N_8841,N_8564,N_8560);
xnor U8842 (N_8842,N_8520,N_8528);
nor U8843 (N_8843,N_8610,N_8516);
or U8844 (N_8844,N_8629,N_8715);
and U8845 (N_8845,N_8568,N_8669);
nand U8846 (N_8846,N_8547,N_8646);
nand U8847 (N_8847,N_8690,N_8575);
or U8848 (N_8848,N_8557,N_8739);
or U8849 (N_8849,N_8681,N_8506);
or U8850 (N_8850,N_8697,N_8748);
nor U8851 (N_8851,N_8590,N_8691);
and U8852 (N_8852,N_8684,N_8642);
nand U8853 (N_8853,N_8596,N_8694);
nor U8854 (N_8854,N_8539,N_8534);
xor U8855 (N_8855,N_8576,N_8744);
nand U8856 (N_8856,N_8588,N_8514);
nor U8857 (N_8857,N_8734,N_8585);
or U8858 (N_8858,N_8548,N_8632);
nand U8859 (N_8859,N_8503,N_8558);
nand U8860 (N_8860,N_8732,N_8578);
xnor U8861 (N_8861,N_8567,N_8580);
nor U8862 (N_8862,N_8693,N_8649);
and U8863 (N_8863,N_8709,N_8626);
or U8864 (N_8864,N_8552,N_8574);
or U8865 (N_8865,N_8679,N_8551);
nand U8866 (N_8866,N_8725,N_8513);
xnor U8867 (N_8867,N_8666,N_8656);
nor U8868 (N_8868,N_8525,N_8512);
nor U8869 (N_8869,N_8591,N_8742);
xnor U8870 (N_8870,N_8705,N_8641);
and U8871 (N_8871,N_8627,N_8579);
nand U8872 (N_8872,N_8571,N_8542);
and U8873 (N_8873,N_8657,N_8584);
nor U8874 (N_8874,N_8648,N_8717);
or U8875 (N_8875,N_8697,N_8732);
nand U8876 (N_8876,N_8532,N_8707);
or U8877 (N_8877,N_8662,N_8736);
nor U8878 (N_8878,N_8594,N_8519);
and U8879 (N_8879,N_8513,N_8685);
nor U8880 (N_8880,N_8690,N_8612);
and U8881 (N_8881,N_8502,N_8563);
nor U8882 (N_8882,N_8526,N_8535);
or U8883 (N_8883,N_8663,N_8556);
xnor U8884 (N_8884,N_8545,N_8576);
and U8885 (N_8885,N_8687,N_8743);
xor U8886 (N_8886,N_8636,N_8679);
nor U8887 (N_8887,N_8728,N_8691);
xor U8888 (N_8888,N_8716,N_8720);
nor U8889 (N_8889,N_8506,N_8581);
xnor U8890 (N_8890,N_8522,N_8648);
nor U8891 (N_8891,N_8641,N_8653);
xor U8892 (N_8892,N_8570,N_8632);
xnor U8893 (N_8893,N_8501,N_8586);
xnor U8894 (N_8894,N_8535,N_8729);
nand U8895 (N_8895,N_8601,N_8667);
or U8896 (N_8896,N_8642,N_8668);
nor U8897 (N_8897,N_8679,N_8614);
nor U8898 (N_8898,N_8676,N_8674);
xnor U8899 (N_8899,N_8588,N_8724);
xnor U8900 (N_8900,N_8743,N_8711);
xor U8901 (N_8901,N_8656,N_8695);
xor U8902 (N_8902,N_8582,N_8513);
nor U8903 (N_8903,N_8546,N_8681);
nand U8904 (N_8904,N_8610,N_8687);
or U8905 (N_8905,N_8636,N_8545);
and U8906 (N_8906,N_8629,N_8534);
and U8907 (N_8907,N_8570,N_8587);
xor U8908 (N_8908,N_8721,N_8559);
nor U8909 (N_8909,N_8548,N_8599);
or U8910 (N_8910,N_8516,N_8674);
nand U8911 (N_8911,N_8582,N_8707);
nor U8912 (N_8912,N_8536,N_8504);
xnor U8913 (N_8913,N_8667,N_8655);
or U8914 (N_8914,N_8688,N_8661);
and U8915 (N_8915,N_8601,N_8733);
xor U8916 (N_8916,N_8637,N_8679);
or U8917 (N_8917,N_8511,N_8573);
nor U8918 (N_8918,N_8744,N_8613);
nor U8919 (N_8919,N_8526,N_8557);
and U8920 (N_8920,N_8622,N_8562);
nor U8921 (N_8921,N_8561,N_8550);
nand U8922 (N_8922,N_8621,N_8681);
or U8923 (N_8923,N_8687,N_8706);
xor U8924 (N_8924,N_8642,N_8648);
nand U8925 (N_8925,N_8541,N_8661);
nand U8926 (N_8926,N_8660,N_8745);
nor U8927 (N_8927,N_8629,N_8524);
nor U8928 (N_8928,N_8632,N_8525);
xor U8929 (N_8929,N_8669,N_8567);
nand U8930 (N_8930,N_8684,N_8731);
or U8931 (N_8931,N_8549,N_8684);
and U8932 (N_8932,N_8614,N_8610);
nor U8933 (N_8933,N_8530,N_8711);
xor U8934 (N_8934,N_8612,N_8700);
nand U8935 (N_8935,N_8533,N_8742);
nor U8936 (N_8936,N_8636,N_8701);
xnor U8937 (N_8937,N_8644,N_8715);
xnor U8938 (N_8938,N_8642,N_8562);
and U8939 (N_8939,N_8589,N_8536);
or U8940 (N_8940,N_8701,N_8742);
and U8941 (N_8941,N_8644,N_8671);
nor U8942 (N_8942,N_8623,N_8679);
nand U8943 (N_8943,N_8707,N_8503);
xor U8944 (N_8944,N_8715,N_8516);
nor U8945 (N_8945,N_8655,N_8731);
nor U8946 (N_8946,N_8724,N_8602);
and U8947 (N_8947,N_8572,N_8578);
nor U8948 (N_8948,N_8561,N_8596);
nand U8949 (N_8949,N_8612,N_8696);
and U8950 (N_8950,N_8618,N_8622);
and U8951 (N_8951,N_8545,N_8583);
xnor U8952 (N_8952,N_8509,N_8646);
or U8953 (N_8953,N_8625,N_8695);
and U8954 (N_8954,N_8501,N_8554);
xor U8955 (N_8955,N_8685,N_8741);
nor U8956 (N_8956,N_8657,N_8607);
and U8957 (N_8957,N_8585,N_8727);
nor U8958 (N_8958,N_8664,N_8683);
and U8959 (N_8959,N_8590,N_8686);
xnor U8960 (N_8960,N_8719,N_8558);
nand U8961 (N_8961,N_8534,N_8660);
xnor U8962 (N_8962,N_8647,N_8527);
nor U8963 (N_8963,N_8727,N_8729);
nor U8964 (N_8964,N_8529,N_8649);
nand U8965 (N_8965,N_8505,N_8552);
nor U8966 (N_8966,N_8561,N_8724);
nand U8967 (N_8967,N_8511,N_8743);
nand U8968 (N_8968,N_8611,N_8515);
nand U8969 (N_8969,N_8566,N_8588);
nor U8970 (N_8970,N_8712,N_8529);
nor U8971 (N_8971,N_8596,N_8728);
nor U8972 (N_8972,N_8566,N_8641);
xor U8973 (N_8973,N_8714,N_8555);
or U8974 (N_8974,N_8515,N_8508);
and U8975 (N_8975,N_8624,N_8686);
nand U8976 (N_8976,N_8647,N_8661);
or U8977 (N_8977,N_8653,N_8729);
or U8978 (N_8978,N_8727,N_8645);
nand U8979 (N_8979,N_8565,N_8527);
nor U8980 (N_8980,N_8614,N_8553);
and U8981 (N_8981,N_8722,N_8638);
xor U8982 (N_8982,N_8598,N_8734);
and U8983 (N_8983,N_8506,N_8645);
or U8984 (N_8984,N_8723,N_8605);
xnor U8985 (N_8985,N_8732,N_8572);
or U8986 (N_8986,N_8557,N_8724);
or U8987 (N_8987,N_8554,N_8591);
nor U8988 (N_8988,N_8515,N_8724);
or U8989 (N_8989,N_8742,N_8578);
or U8990 (N_8990,N_8502,N_8550);
xnor U8991 (N_8991,N_8558,N_8538);
nor U8992 (N_8992,N_8554,N_8654);
nor U8993 (N_8993,N_8748,N_8732);
or U8994 (N_8994,N_8741,N_8689);
xor U8995 (N_8995,N_8742,N_8566);
xor U8996 (N_8996,N_8553,N_8583);
or U8997 (N_8997,N_8529,N_8599);
nor U8998 (N_8998,N_8737,N_8728);
or U8999 (N_8999,N_8696,N_8646);
and U9000 (N_9000,N_8819,N_8903);
xor U9001 (N_9001,N_8944,N_8970);
nand U9002 (N_9002,N_8849,N_8932);
nand U9003 (N_9003,N_8972,N_8825);
or U9004 (N_9004,N_8826,N_8981);
and U9005 (N_9005,N_8843,N_8909);
xnor U9006 (N_9006,N_8796,N_8942);
xnor U9007 (N_9007,N_8894,N_8862);
or U9008 (N_9008,N_8965,N_8791);
nand U9009 (N_9009,N_8812,N_8829);
xor U9010 (N_9010,N_8982,N_8848);
nand U9011 (N_9011,N_8879,N_8954);
nor U9012 (N_9012,N_8898,N_8931);
or U9013 (N_9013,N_8810,N_8856);
nor U9014 (N_9014,N_8824,N_8799);
nor U9015 (N_9015,N_8753,N_8927);
nor U9016 (N_9016,N_8989,N_8947);
nor U9017 (N_9017,N_8966,N_8871);
nand U9018 (N_9018,N_8919,N_8766);
and U9019 (N_9019,N_8850,N_8969);
xnor U9020 (N_9020,N_8764,N_8951);
or U9021 (N_9021,N_8789,N_8962);
and U9022 (N_9022,N_8797,N_8758);
nor U9023 (N_9023,N_8784,N_8937);
xor U9024 (N_9024,N_8977,N_8952);
nand U9025 (N_9025,N_8751,N_8876);
nand U9026 (N_9026,N_8974,N_8887);
xor U9027 (N_9027,N_8816,N_8908);
and U9028 (N_9028,N_8960,N_8756);
and U9029 (N_9029,N_8923,N_8990);
and U9030 (N_9030,N_8901,N_8983);
xor U9031 (N_9031,N_8866,N_8867);
and U9032 (N_9032,N_8897,N_8820);
and U9033 (N_9033,N_8997,N_8788);
nand U9034 (N_9034,N_8759,N_8993);
and U9035 (N_9035,N_8823,N_8750);
nor U9036 (N_9036,N_8940,N_8979);
or U9037 (N_9037,N_8853,N_8861);
or U9038 (N_9038,N_8805,N_8803);
xnor U9039 (N_9039,N_8831,N_8991);
xnor U9040 (N_9040,N_8775,N_8793);
nor U9041 (N_9041,N_8754,N_8815);
nand U9042 (N_9042,N_8811,N_8770);
xor U9043 (N_9043,N_8855,N_8837);
nor U9044 (N_9044,N_8808,N_8883);
and U9045 (N_9045,N_8978,N_8984);
xor U9046 (N_9046,N_8884,N_8762);
and U9047 (N_9047,N_8961,N_8941);
nor U9048 (N_9048,N_8905,N_8798);
nand U9049 (N_9049,N_8839,N_8918);
nand U9050 (N_9050,N_8920,N_8779);
nand U9051 (N_9051,N_8891,N_8928);
or U9052 (N_9052,N_8847,N_8773);
nand U9053 (N_9053,N_8841,N_8907);
nand U9054 (N_9054,N_8953,N_8889);
or U9055 (N_9055,N_8765,N_8801);
nor U9056 (N_9056,N_8921,N_8986);
nor U9057 (N_9057,N_8878,N_8963);
and U9058 (N_9058,N_8822,N_8769);
nand U9059 (N_9059,N_8911,N_8774);
nand U9060 (N_9060,N_8776,N_8895);
nor U9061 (N_9061,N_8948,N_8790);
nor U9062 (N_9062,N_8760,N_8994);
nor U9063 (N_9063,N_8992,N_8830);
nor U9064 (N_9064,N_8922,N_8783);
nor U9065 (N_9065,N_8834,N_8886);
nand U9066 (N_9066,N_8926,N_8869);
and U9067 (N_9067,N_8821,N_8802);
and U9068 (N_9068,N_8827,N_8781);
nor U9069 (N_9069,N_8755,N_8800);
and U9070 (N_9070,N_8971,N_8945);
and U9071 (N_9071,N_8868,N_8957);
xor U9072 (N_9072,N_8875,N_8881);
nor U9073 (N_9073,N_8842,N_8964);
and U9074 (N_9074,N_8845,N_8934);
or U9075 (N_9075,N_8930,N_8806);
nor U9076 (N_9076,N_8852,N_8864);
and U9077 (N_9077,N_8836,N_8767);
nand U9078 (N_9078,N_8778,N_8949);
nand U9079 (N_9079,N_8817,N_8840);
nor U9080 (N_9080,N_8795,N_8858);
nor U9081 (N_9081,N_8780,N_8863);
nor U9082 (N_9082,N_8777,N_8950);
and U9083 (N_9083,N_8936,N_8873);
nor U9084 (N_9084,N_8914,N_8757);
nand U9085 (N_9085,N_8851,N_8888);
nor U9086 (N_9086,N_8956,N_8935);
and U9087 (N_9087,N_8752,N_8859);
and U9088 (N_9088,N_8885,N_8860);
xnor U9089 (N_9089,N_8900,N_8917);
nor U9090 (N_9090,N_8814,N_8828);
xor U9091 (N_9091,N_8998,N_8771);
nand U9092 (N_9092,N_8786,N_8976);
nor U9093 (N_9093,N_8838,N_8761);
nor U9094 (N_9094,N_8782,N_8904);
and U9095 (N_9095,N_8890,N_8959);
nand U9096 (N_9096,N_8785,N_8955);
nand U9097 (N_9097,N_8763,N_8938);
nand U9098 (N_9098,N_8877,N_8995);
xnor U9099 (N_9099,N_8946,N_8833);
xor U9100 (N_9100,N_8893,N_8792);
nor U9101 (N_9101,N_8865,N_8844);
xnor U9102 (N_9102,N_8912,N_8999);
or U9103 (N_9103,N_8874,N_8902);
or U9104 (N_9104,N_8975,N_8925);
nor U9105 (N_9105,N_8880,N_8967);
and U9106 (N_9106,N_8813,N_8768);
and U9107 (N_9107,N_8933,N_8807);
or U9108 (N_9108,N_8943,N_8857);
nand U9109 (N_9109,N_8929,N_8916);
xor U9110 (N_9110,N_8915,N_8939);
nand U9111 (N_9111,N_8772,N_8804);
nand U9112 (N_9112,N_8968,N_8973);
or U9113 (N_9113,N_8899,N_8906);
or U9114 (N_9114,N_8958,N_8882);
nand U9115 (N_9115,N_8996,N_8913);
xnor U9116 (N_9116,N_8809,N_8985);
or U9117 (N_9117,N_8794,N_8988);
or U9118 (N_9118,N_8818,N_8835);
xor U9119 (N_9119,N_8892,N_8854);
nor U9120 (N_9120,N_8910,N_8832);
or U9121 (N_9121,N_8787,N_8846);
xnor U9122 (N_9122,N_8896,N_8987);
and U9123 (N_9123,N_8980,N_8870);
nor U9124 (N_9124,N_8872,N_8924);
nand U9125 (N_9125,N_8755,N_8956);
xor U9126 (N_9126,N_8817,N_8994);
nand U9127 (N_9127,N_8983,N_8948);
nor U9128 (N_9128,N_8773,N_8961);
nand U9129 (N_9129,N_8904,N_8913);
and U9130 (N_9130,N_8895,N_8844);
nand U9131 (N_9131,N_8842,N_8823);
nor U9132 (N_9132,N_8853,N_8827);
nor U9133 (N_9133,N_8951,N_8883);
nand U9134 (N_9134,N_8878,N_8962);
xnor U9135 (N_9135,N_8772,N_8791);
and U9136 (N_9136,N_8814,N_8858);
nor U9137 (N_9137,N_8809,N_8951);
and U9138 (N_9138,N_8808,N_8873);
nand U9139 (N_9139,N_8932,N_8756);
xnor U9140 (N_9140,N_8849,N_8845);
and U9141 (N_9141,N_8999,N_8831);
nor U9142 (N_9142,N_8806,N_8866);
or U9143 (N_9143,N_8845,N_8989);
nand U9144 (N_9144,N_8750,N_8769);
and U9145 (N_9145,N_8868,N_8967);
xnor U9146 (N_9146,N_8891,N_8837);
nand U9147 (N_9147,N_8996,N_8817);
and U9148 (N_9148,N_8776,N_8833);
and U9149 (N_9149,N_8845,N_8836);
or U9150 (N_9150,N_8982,N_8897);
xnor U9151 (N_9151,N_8982,N_8983);
or U9152 (N_9152,N_8963,N_8850);
and U9153 (N_9153,N_8795,N_8846);
nand U9154 (N_9154,N_8873,N_8844);
nor U9155 (N_9155,N_8810,N_8904);
nand U9156 (N_9156,N_8963,N_8811);
xnor U9157 (N_9157,N_8801,N_8920);
or U9158 (N_9158,N_8959,N_8942);
nor U9159 (N_9159,N_8768,N_8898);
or U9160 (N_9160,N_8809,N_8795);
nor U9161 (N_9161,N_8909,N_8778);
nand U9162 (N_9162,N_8802,N_8910);
and U9163 (N_9163,N_8978,N_8933);
nand U9164 (N_9164,N_8924,N_8766);
xor U9165 (N_9165,N_8799,N_8963);
xnor U9166 (N_9166,N_8936,N_8911);
and U9167 (N_9167,N_8839,N_8854);
and U9168 (N_9168,N_8882,N_8963);
xor U9169 (N_9169,N_8972,N_8926);
and U9170 (N_9170,N_8972,N_8787);
and U9171 (N_9171,N_8941,N_8857);
and U9172 (N_9172,N_8757,N_8945);
and U9173 (N_9173,N_8874,N_8944);
nand U9174 (N_9174,N_8866,N_8805);
or U9175 (N_9175,N_8929,N_8910);
and U9176 (N_9176,N_8826,N_8835);
or U9177 (N_9177,N_8884,N_8866);
nor U9178 (N_9178,N_8996,N_8867);
nor U9179 (N_9179,N_8904,N_8865);
and U9180 (N_9180,N_8877,N_8865);
xnor U9181 (N_9181,N_8873,N_8910);
nand U9182 (N_9182,N_8848,N_8935);
nor U9183 (N_9183,N_8786,N_8991);
nor U9184 (N_9184,N_8852,N_8842);
nand U9185 (N_9185,N_8781,N_8888);
xnor U9186 (N_9186,N_8778,N_8793);
xor U9187 (N_9187,N_8921,N_8886);
and U9188 (N_9188,N_8979,N_8810);
nand U9189 (N_9189,N_8794,N_8880);
or U9190 (N_9190,N_8965,N_8797);
xnor U9191 (N_9191,N_8786,N_8775);
nand U9192 (N_9192,N_8877,N_8948);
and U9193 (N_9193,N_8999,N_8923);
and U9194 (N_9194,N_8810,N_8854);
or U9195 (N_9195,N_8875,N_8952);
nand U9196 (N_9196,N_8781,N_8761);
xnor U9197 (N_9197,N_8753,N_8953);
nor U9198 (N_9198,N_8756,N_8901);
nor U9199 (N_9199,N_8915,N_8870);
xnor U9200 (N_9200,N_8783,N_8948);
nor U9201 (N_9201,N_8940,N_8779);
nand U9202 (N_9202,N_8919,N_8783);
and U9203 (N_9203,N_8856,N_8915);
or U9204 (N_9204,N_8821,N_8789);
nor U9205 (N_9205,N_8811,N_8841);
nand U9206 (N_9206,N_8947,N_8976);
and U9207 (N_9207,N_8869,N_8995);
nor U9208 (N_9208,N_8816,N_8754);
xor U9209 (N_9209,N_8941,N_8814);
nor U9210 (N_9210,N_8910,N_8999);
nand U9211 (N_9211,N_8996,N_8837);
nor U9212 (N_9212,N_8882,N_8877);
and U9213 (N_9213,N_8960,N_8980);
nand U9214 (N_9214,N_8960,N_8795);
xor U9215 (N_9215,N_8893,N_8891);
nor U9216 (N_9216,N_8965,N_8933);
or U9217 (N_9217,N_8965,N_8942);
nand U9218 (N_9218,N_8999,N_8927);
and U9219 (N_9219,N_8868,N_8896);
xnor U9220 (N_9220,N_8885,N_8872);
xor U9221 (N_9221,N_8759,N_8802);
and U9222 (N_9222,N_8755,N_8908);
nand U9223 (N_9223,N_8998,N_8853);
nand U9224 (N_9224,N_8852,N_8754);
and U9225 (N_9225,N_8815,N_8912);
xor U9226 (N_9226,N_8859,N_8852);
nand U9227 (N_9227,N_8966,N_8978);
or U9228 (N_9228,N_8948,N_8946);
or U9229 (N_9229,N_8939,N_8975);
and U9230 (N_9230,N_8894,N_8816);
nor U9231 (N_9231,N_8830,N_8997);
xnor U9232 (N_9232,N_8909,N_8827);
nor U9233 (N_9233,N_8826,N_8882);
nand U9234 (N_9234,N_8847,N_8933);
nand U9235 (N_9235,N_8853,N_8953);
nor U9236 (N_9236,N_8861,N_8863);
nand U9237 (N_9237,N_8771,N_8986);
or U9238 (N_9238,N_8930,N_8909);
xor U9239 (N_9239,N_8932,N_8838);
xor U9240 (N_9240,N_8947,N_8824);
xnor U9241 (N_9241,N_8965,N_8916);
nand U9242 (N_9242,N_8993,N_8979);
nand U9243 (N_9243,N_8862,N_8939);
and U9244 (N_9244,N_8930,N_8984);
and U9245 (N_9245,N_8921,N_8806);
nor U9246 (N_9246,N_8939,N_8964);
xnor U9247 (N_9247,N_8905,N_8925);
xnor U9248 (N_9248,N_8951,N_8802);
or U9249 (N_9249,N_8960,N_8946);
xnor U9250 (N_9250,N_9138,N_9139);
xnor U9251 (N_9251,N_9163,N_9122);
xor U9252 (N_9252,N_9158,N_9026);
nor U9253 (N_9253,N_9023,N_9191);
or U9254 (N_9254,N_9233,N_9142);
nand U9255 (N_9255,N_9228,N_9125);
xor U9256 (N_9256,N_9113,N_9220);
xnor U9257 (N_9257,N_9237,N_9080);
nand U9258 (N_9258,N_9189,N_9100);
xnor U9259 (N_9259,N_9239,N_9147);
xor U9260 (N_9260,N_9002,N_9104);
nor U9261 (N_9261,N_9036,N_9018);
xnor U9262 (N_9262,N_9157,N_9194);
and U9263 (N_9263,N_9004,N_9044);
nor U9264 (N_9264,N_9222,N_9094);
and U9265 (N_9265,N_9077,N_9082);
nor U9266 (N_9266,N_9008,N_9236);
and U9267 (N_9267,N_9196,N_9073);
or U9268 (N_9268,N_9148,N_9238);
and U9269 (N_9269,N_9035,N_9091);
nand U9270 (N_9270,N_9063,N_9133);
and U9271 (N_9271,N_9182,N_9150);
or U9272 (N_9272,N_9076,N_9223);
and U9273 (N_9273,N_9045,N_9198);
nand U9274 (N_9274,N_9211,N_9181);
xor U9275 (N_9275,N_9209,N_9168);
nand U9276 (N_9276,N_9090,N_9136);
nor U9277 (N_9277,N_9069,N_9056);
xnor U9278 (N_9278,N_9131,N_9192);
and U9279 (N_9279,N_9099,N_9112);
or U9280 (N_9280,N_9053,N_9123);
nor U9281 (N_9281,N_9021,N_9171);
and U9282 (N_9282,N_9014,N_9064);
xor U9283 (N_9283,N_9019,N_9137);
xor U9284 (N_9284,N_9241,N_9052);
and U9285 (N_9285,N_9143,N_9068);
nand U9286 (N_9286,N_9041,N_9006);
xnor U9287 (N_9287,N_9234,N_9025);
nor U9288 (N_9288,N_9200,N_9101);
xor U9289 (N_9289,N_9098,N_9127);
nand U9290 (N_9290,N_9121,N_9201);
and U9291 (N_9291,N_9226,N_9165);
or U9292 (N_9292,N_9183,N_9060);
nor U9293 (N_9293,N_9058,N_9034);
and U9294 (N_9294,N_9102,N_9174);
and U9295 (N_9295,N_9206,N_9040);
nor U9296 (N_9296,N_9205,N_9203);
or U9297 (N_9297,N_9166,N_9154);
nor U9298 (N_9298,N_9176,N_9245);
and U9299 (N_9299,N_9079,N_9027);
nor U9300 (N_9300,N_9081,N_9005);
xnor U9301 (N_9301,N_9075,N_9129);
or U9302 (N_9302,N_9193,N_9055);
nand U9303 (N_9303,N_9199,N_9010);
nand U9304 (N_9304,N_9061,N_9007);
or U9305 (N_9305,N_9132,N_9022);
xnor U9306 (N_9306,N_9086,N_9096);
xor U9307 (N_9307,N_9215,N_9126);
xor U9308 (N_9308,N_9095,N_9107);
nand U9309 (N_9309,N_9225,N_9180);
and U9310 (N_9310,N_9246,N_9167);
nand U9311 (N_9311,N_9031,N_9000);
nand U9312 (N_9312,N_9177,N_9070);
nor U9313 (N_9313,N_9207,N_9197);
nor U9314 (N_9314,N_9011,N_9156);
or U9315 (N_9315,N_9067,N_9092);
or U9316 (N_9316,N_9248,N_9243);
xnor U9317 (N_9317,N_9208,N_9161);
and U9318 (N_9318,N_9155,N_9146);
and U9319 (N_9319,N_9219,N_9172);
nor U9320 (N_9320,N_9048,N_9029);
nand U9321 (N_9321,N_9134,N_9124);
or U9322 (N_9322,N_9145,N_9232);
nand U9323 (N_9323,N_9003,N_9187);
xor U9324 (N_9324,N_9083,N_9151);
nor U9325 (N_9325,N_9097,N_9103);
or U9326 (N_9326,N_9235,N_9013);
nor U9327 (N_9327,N_9050,N_9184);
xnor U9328 (N_9328,N_9179,N_9074);
xnor U9329 (N_9329,N_9062,N_9242);
nand U9330 (N_9330,N_9159,N_9046);
and U9331 (N_9331,N_9160,N_9188);
and U9332 (N_9332,N_9175,N_9153);
or U9333 (N_9333,N_9020,N_9118);
xor U9334 (N_9334,N_9128,N_9185);
nor U9335 (N_9335,N_9015,N_9152);
nor U9336 (N_9336,N_9204,N_9162);
and U9337 (N_9337,N_9141,N_9231);
xor U9338 (N_9338,N_9247,N_9110);
and U9339 (N_9339,N_9178,N_9059);
and U9340 (N_9340,N_9216,N_9049);
xor U9341 (N_9341,N_9093,N_9089);
or U9342 (N_9342,N_9030,N_9221);
or U9343 (N_9343,N_9084,N_9140);
and U9344 (N_9344,N_9149,N_9195);
or U9345 (N_9345,N_9071,N_9227);
nand U9346 (N_9346,N_9117,N_9173);
and U9347 (N_9347,N_9057,N_9212);
and U9348 (N_9348,N_9037,N_9009);
nand U9349 (N_9349,N_9120,N_9087);
nor U9350 (N_9350,N_9190,N_9066);
and U9351 (N_9351,N_9054,N_9028);
or U9352 (N_9352,N_9024,N_9017);
or U9353 (N_9353,N_9164,N_9016);
or U9354 (N_9354,N_9144,N_9115);
nor U9355 (N_9355,N_9038,N_9065);
nand U9356 (N_9356,N_9230,N_9111);
xnor U9357 (N_9357,N_9108,N_9244);
xor U9358 (N_9358,N_9051,N_9130);
nor U9359 (N_9359,N_9033,N_9217);
xor U9360 (N_9360,N_9214,N_9202);
nand U9361 (N_9361,N_9249,N_9072);
nor U9362 (N_9362,N_9169,N_9039);
and U9363 (N_9363,N_9240,N_9043);
and U9364 (N_9364,N_9105,N_9213);
nor U9365 (N_9365,N_9218,N_9186);
and U9366 (N_9366,N_9114,N_9106);
nor U9367 (N_9367,N_9119,N_9229);
nand U9368 (N_9368,N_9170,N_9078);
xnor U9369 (N_9369,N_9224,N_9047);
xnor U9370 (N_9370,N_9116,N_9088);
nand U9371 (N_9371,N_9210,N_9109);
nand U9372 (N_9372,N_9012,N_9085);
and U9373 (N_9373,N_9135,N_9032);
xor U9374 (N_9374,N_9001,N_9042);
or U9375 (N_9375,N_9122,N_9031);
or U9376 (N_9376,N_9038,N_9099);
xnor U9377 (N_9377,N_9203,N_9215);
xnor U9378 (N_9378,N_9154,N_9056);
nor U9379 (N_9379,N_9116,N_9038);
and U9380 (N_9380,N_9239,N_9014);
or U9381 (N_9381,N_9193,N_9189);
and U9382 (N_9382,N_9075,N_9079);
xnor U9383 (N_9383,N_9080,N_9203);
nand U9384 (N_9384,N_9242,N_9081);
xnor U9385 (N_9385,N_9244,N_9007);
or U9386 (N_9386,N_9063,N_9097);
or U9387 (N_9387,N_9166,N_9230);
nor U9388 (N_9388,N_9107,N_9182);
or U9389 (N_9389,N_9208,N_9177);
nor U9390 (N_9390,N_9061,N_9058);
or U9391 (N_9391,N_9235,N_9139);
nor U9392 (N_9392,N_9070,N_9141);
and U9393 (N_9393,N_9191,N_9038);
or U9394 (N_9394,N_9144,N_9227);
nand U9395 (N_9395,N_9115,N_9050);
xor U9396 (N_9396,N_9216,N_9234);
nor U9397 (N_9397,N_9246,N_9213);
and U9398 (N_9398,N_9024,N_9243);
and U9399 (N_9399,N_9203,N_9154);
nor U9400 (N_9400,N_9074,N_9007);
nor U9401 (N_9401,N_9031,N_9005);
nand U9402 (N_9402,N_9011,N_9157);
and U9403 (N_9403,N_9164,N_9056);
and U9404 (N_9404,N_9201,N_9127);
nor U9405 (N_9405,N_9173,N_9193);
nand U9406 (N_9406,N_9179,N_9091);
nand U9407 (N_9407,N_9204,N_9145);
xor U9408 (N_9408,N_9184,N_9092);
xnor U9409 (N_9409,N_9206,N_9205);
nor U9410 (N_9410,N_9090,N_9080);
nand U9411 (N_9411,N_9069,N_9226);
or U9412 (N_9412,N_9146,N_9085);
nor U9413 (N_9413,N_9054,N_9074);
or U9414 (N_9414,N_9100,N_9215);
or U9415 (N_9415,N_9066,N_9233);
nand U9416 (N_9416,N_9101,N_9240);
and U9417 (N_9417,N_9180,N_9137);
nand U9418 (N_9418,N_9203,N_9115);
nor U9419 (N_9419,N_9232,N_9041);
or U9420 (N_9420,N_9070,N_9012);
or U9421 (N_9421,N_9054,N_9194);
xnor U9422 (N_9422,N_9149,N_9122);
xor U9423 (N_9423,N_9208,N_9077);
nand U9424 (N_9424,N_9206,N_9041);
and U9425 (N_9425,N_9246,N_9067);
or U9426 (N_9426,N_9238,N_9165);
nor U9427 (N_9427,N_9060,N_9123);
xnor U9428 (N_9428,N_9106,N_9177);
and U9429 (N_9429,N_9045,N_9248);
or U9430 (N_9430,N_9010,N_9234);
or U9431 (N_9431,N_9077,N_9055);
nor U9432 (N_9432,N_9177,N_9037);
and U9433 (N_9433,N_9034,N_9182);
or U9434 (N_9434,N_9067,N_9055);
xnor U9435 (N_9435,N_9035,N_9139);
or U9436 (N_9436,N_9156,N_9113);
or U9437 (N_9437,N_9120,N_9222);
and U9438 (N_9438,N_9151,N_9209);
nand U9439 (N_9439,N_9064,N_9167);
and U9440 (N_9440,N_9041,N_9096);
nor U9441 (N_9441,N_9146,N_9047);
xor U9442 (N_9442,N_9144,N_9176);
nand U9443 (N_9443,N_9060,N_9188);
or U9444 (N_9444,N_9199,N_9180);
nand U9445 (N_9445,N_9124,N_9126);
nand U9446 (N_9446,N_9099,N_9001);
xor U9447 (N_9447,N_9035,N_9095);
and U9448 (N_9448,N_9176,N_9147);
nand U9449 (N_9449,N_9193,N_9034);
xnor U9450 (N_9450,N_9060,N_9156);
nand U9451 (N_9451,N_9171,N_9081);
xnor U9452 (N_9452,N_9099,N_9030);
nand U9453 (N_9453,N_9186,N_9067);
or U9454 (N_9454,N_9076,N_9075);
nand U9455 (N_9455,N_9154,N_9233);
nand U9456 (N_9456,N_9023,N_9070);
nand U9457 (N_9457,N_9016,N_9234);
nand U9458 (N_9458,N_9196,N_9189);
and U9459 (N_9459,N_9181,N_9078);
nand U9460 (N_9460,N_9018,N_9043);
or U9461 (N_9461,N_9009,N_9136);
and U9462 (N_9462,N_9147,N_9152);
xnor U9463 (N_9463,N_9034,N_9232);
and U9464 (N_9464,N_9229,N_9064);
nand U9465 (N_9465,N_9113,N_9057);
nor U9466 (N_9466,N_9180,N_9006);
nor U9467 (N_9467,N_9180,N_9018);
or U9468 (N_9468,N_9085,N_9095);
nand U9469 (N_9469,N_9065,N_9196);
or U9470 (N_9470,N_9187,N_9135);
and U9471 (N_9471,N_9051,N_9097);
xnor U9472 (N_9472,N_9171,N_9227);
or U9473 (N_9473,N_9151,N_9060);
or U9474 (N_9474,N_9082,N_9015);
nand U9475 (N_9475,N_9172,N_9134);
and U9476 (N_9476,N_9244,N_9128);
and U9477 (N_9477,N_9207,N_9061);
or U9478 (N_9478,N_9161,N_9095);
nor U9479 (N_9479,N_9103,N_9003);
or U9480 (N_9480,N_9132,N_9182);
nor U9481 (N_9481,N_9032,N_9164);
xnor U9482 (N_9482,N_9029,N_9009);
xnor U9483 (N_9483,N_9221,N_9186);
nor U9484 (N_9484,N_9162,N_9244);
and U9485 (N_9485,N_9228,N_9108);
nand U9486 (N_9486,N_9125,N_9019);
and U9487 (N_9487,N_9049,N_9179);
nand U9488 (N_9488,N_9126,N_9220);
and U9489 (N_9489,N_9212,N_9176);
nand U9490 (N_9490,N_9181,N_9136);
xor U9491 (N_9491,N_9225,N_9170);
nor U9492 (N_9492,N_9025,N_9167);
nand U9493 (N_9493,N_9242,N_9122);
xnor U9494 (N_9494,N_9001,N_9061);
and U9495 (N_9495,N_9190,N_9237);
and U9496 (N_9496,N_9139,N_9085);
xor U9497 (N_9497,N_9170,N_9088);
nor U9498 (N_9498,N_9128,N_9148);
xor U9499 (N_9499,N_9239,N_9116);
nand U9500 (N_9500,N_9334,N_9279);
and U9501 (N_9501,N_9430,N_9385);
and U9502 (N_9502,N_9256,N_9319);
or U9503 (N_9503,N_9281,N_9446);
or U9504 (N_9504,N_9408,N_9358);
nand U9505 (N_9505,N_9255,N_9481);
or U9506 (N_9506,N_9463,N_9396);
nand U9507 (N_9507,N_9389,N_9304);
nand U9508 (N_9508,N_9283,N_9269);
xnor U9509 (N_9509,N_9404,N_9315);
nand U9510 (N_9510,N_9441,N_9376);
and U9511 (N_9511,N_9331,N_9388);
xnor U9512 (N_9512,N_9424,N_9291);
xor U9513 (N_9513,N_9412,N_9299);
xor U9514 (N_9514,N_9253,N_9305);
or U9515 (N_9515,N_9405,N_9455);
nand U9516 (N_9516,N_9250,N_9436);
nand U9517 (N_9517,N_9363,N_9369);
nor U9518 (N_9518,N_9414,N_9286);
xnor U9519 (N_9519,N_9333,N_9348);
nor U9520 (N_9520,N_9309,N_9438);
nand U9521 (N_9521,N_9415,N_9377);
xor U9522 (N_9522,N_9382,N_9409);
and U9523 (N_9523,N_9322,N_9459);
and U9524 (N_9524,N_9351,N_9393);
xnor U9525 (N_9525,N_9442,N_9311);
nand U9526 (N_9526,N_9476,N_9471);
xnor U9527 (N_9527,N_9372,N_9468);
nand U9528 (N_9528,N_9359,N_9312);
or U9529 (N_9529,N_9493,N_9294);
and U9530 (N_9530,N_9267,N_9298);
or U9531 (N_9531,N_9394,N_9306);
nand U9532 (N_9532,N_9303,N_9474);
nand U9533 (N_9533,N_9482,N_9375);
and U9534 (N_9534,N_9284,N_9433);
and U9535 (N_9535,N_9277,N_9371);
or U9536 (N_9536,N_9439,N_9460);
nand U9537 (N_9537,N_9308,N_9456);
nand U9538 (N_9538,N_9466,N_9307);
xnor U9539 (N_9539,N_9349,N_9383);
nand U9540 (N_9540,N_9258,N_9379);
and U9541 (N_9541,N_9448,N_9457);
or U9542 (N_9542,N_9338,N_9367);
nor U9543 (N_9543,N_9357,N_9260);
nand U9544 (N_9544,N_9346,N_9440);
xnor U9545 (N_9545,N_9452,N_9266);
and U9546 (N_9546,N_9332,N_9499);
and U9547 (N_9547,N_9340,N_9380);
xnor U9548 (N_9548,N_9453,N_9418);
and U9549 (N_9549,N_9313,N_9347);
xnor U9550 (N_9550,N_9352,N_9435);
or U9551 (N_9551,N_9330,N_9450);
or U9552 (N_9552,N_9310,N_9289);
and U9553 (N_9553,N_9287,N_9300);
nand U9554 (N_9554,N_9302,N_9496);
xor U9555 (N_9555,N_9278,N_9336);
and U9556 (N_9556,N_9406,N_9434);
and U9557 (N_9557,N_9323,N_9354);
xor U9558 (N_9558,N_9417,N_9282);
nand U9559 (N_9559,N_9373,N_9398);
and U9560 (N_9560,N_9270,N_9437);
or U9561 (N_9561,N_9397,N_9480);
and U9562 (N_9562,N_9462,N_9413);
nand U9563 (N_9563,N_9478,N_9273);
and U9564 (N_9564,N_9314,N_9264);
or U9565 (N_9565,N_9467,N_9420);
and U9566 (N_9566,N_9360,N_9350);
or U9567 (N_9567,N_9275,N_9479);
nor U9568 (N_9568,N_9262,N_9387);
or U9569 (N_9569,N_9419,N_9321);
and U9570 (N_9570,N_9489,N_9342);
or U9571 (N_9571,N_9491,N_9423);
nor U9572 (N_9572,N_9458,N_9259);
xor U9573 (N_9573,N_9401,N_9411);
nor U9574 (N_9574,N_9329,N_9384);
nand U9575 (N_9575,N_9390,N_9431);
nand U9576 (N_9576,N_9297,N_9252);
nand U9577 (N_9577,N_9427,N_9475);
nor U9578 (N_9578,N_9318,N_9301);
nand U9579 (N_9579,N_9407,N_9445);
xor U9580 (N_9580,N_9274,N_9386);
and U9581 (N_9581,N_9341,N_9449);
nor U9582 (N_9582,N_9251,N_9464);
nand U9583 (N_9583,N_9374,N_9402);
xnor U9584 (N_9584,N_9444,N_9381);
xor U9585 (N_9585,N_9324,N_9366);
or U9586 (N_9586,N_9343,N_9432);
or U9587 (N_9587,N_9485,N_9316);
xnor U9588 (N_9588,N_9272,N_9320);
nor U9589 (N_9589,N_9362,N_9477);
or U9590 (N_9590,N_9365,N_9425);
or U9591 (N_9591,N_9364,N_9483);
and U9592 (N_9592,N_9355,N_9490);
nand U9593 (N_9593,N_9265,N_9370);
and U9594 (N_9594,N_9400,N_9498);
and U9595 (N_9595,N_9378,N_9470);
nor U9596 (N_9596,N_9497,N_9392);
and U9597 (N_9597,N_9328,N_9454);
or U9598 (N_9598,N_9484,N_9361);
and U9599 (N_9599,N_9395,N_9326);
and U9600 (N_9600,N_9426,N_9288);
xnor U9601 (N_9601,N_9292,N_9403);
or U9602 (N_9602,N_9327,N_9261);
nand U9603 (N_9603,N_9317,N_9416);
xnor U9604 (N_9604,N_9353,N_9494);
xor U9605 (N_9605,N_9296,N_9472);
xor U9606 (N_9606,N_9421,N_9268);
or U9607 (N_9607,N_9280,N_9486);
nand U9608 (N_9608,N_9492,N_9368);
and U9609 (N_9609,N_9488,N_9356);
and U9610 (N_9610,N_9487,N_9447);
nand U9611 (N_9611,N_9290,N_9451);
nand U9612 (N_9612,N_9335,N_9276);
or U9613 (N_9613,N_9257,N_9461);
xnor U9614 (N_9614,N_9399,N_9345);
and U9615 (N_9615,N_9339,N_9428);
and U9616 (N_9616,N_9422,N_9410);
xor U9617 (N_9617,N_9271,N_9473);
xnor U9618 (N_9618,N_9285,N_9495);
nor U9619 (N_9619,N_9391,N_9263);
nand U9620 (N_9620,N_9469,N_9295);
or U9621 (N_9621,N_9293,N_9429);
xor U9622 (N_9622,N_9325,N_9443);
or U9623 (N_9623,N_9254,N_9465);
xnor U9624 (N_9624,N_9344,N_9337);
or U9625 (N_9625,N_9429,N_9497);
nand U9626 (N_9626,N_9492,N_9311);
nand U9627 (N_9627,N_9455,N_9295);
nor U9628 (N_9628,N_9367,N_9274);
or U9629 (N_9629,N_9446,N_9381);
nor U9630 (N_9630,N_9345,N_9453);
or U9631 (N_9631,N_9262,N_9395);
and U9632 (N_9632,N_9316,N_9312);
nor U9633 (N_9633,N_9452,N_9279);
xnor U9634 (N_9634,N_9256,N_9340);
or U9635 (N_9635,N_9308,N_9294);
nor U9636 (N_9636,N_9429,N_9399);
and U9637 (N_9637,N_9258,N_9318);
xor U9638 (N_9638,N_9439,N_9446);
xnor U9639 (N_9639,N_9322,N_9289);
or U9640 (N_9640,N_9370,N_9328);
nor U9641 (N_9641,N_9475,N_9368);
nand U9642 (N_9642,N_9262,N_9358);
or U9643 (N_9643,N_9405,N_9475);
xnor U9644 (N_9644,N_9489,N_9436);
nand U9645 (N_9645,N_9377,N_9459);
xnor U9646 (N_9646,N_9339,N_9422);
nand U9647 (N_9647,N_9426,N_9267);
or U9648 (N_9648,N_9252,N_9412);
nand U9649 (N_9649,N_9444,N_9311);
xor U9650 (N_9650,N_9457,N_9266);
or U9651 (N_9651,N_9395,N_9416);
nand U9652 (N_9652,N_9320,N_9296);
or U9653 (N_9653,N_9360,N_9315);
nor U9654 (N_9654,N_9357,N_9466);
or U9655 (N_9655,N_9482,N_9361);
and U9656 (N_9656,N_9450,N_9498);
or U9657 (N_9657,N_9340,N_9282);
and U9658 (N_9658,N_9373,N_9358);
nand U9659 (N_9659,N_9444,N_9408);
nand U9660 (N_9660,N_9445,N_9393);
and U9661 (N_9661,N_9491,N_9470);
nand U9662 (N_9662,N_9414,N_9445);
nor U9663 (N_9663,N_9255,N_9397);
and U9664 (N_9664,N_9358,N_9336);
nor U9665 (N_9665,N_9348,N_9438);
nand U9666 (N_9666,N_9302,N_9408);
nand U9667 (N_9667,N_9396,N_9253);
or U9668 (N_9668,N_9329,N_9379);
nand U9669 (N_9669,N_9435,N_9473);
or U9670 (N_9670,N_9303,N_9319);
nor U9671 (N_9671,N_9426,N_9316);
or U9672 (N_9672,N_9471,N_9289);
xor U9673 (N_9673,N_9310,N_9446);
and U9674 (N_9674,N_9345,N_9277);
nand U9675 (N_9675,N_9464,N_9271);
nand U9676 (N_9676,N_9263,N_9379);
and U9677 (N_9677,N_9430,N_9474);
and U9678 (N_9678,N_9358,N_9470);
and U9679 (N_9679,N_9297,N_9370);
and U9680 (N_9680,N_9474,N_9263);
or U9681 (N_9681,N_9420,N_9442);
nor U9682 (N_9682,N_9468,N_9414);
or U9683 (N_9683,N_9424,N_9462);
and U9684 (N_9684,N_9400,N_9462);
xnor U9685 (N_9685,N_9437,N_9337);
nor U9686 (N_9686,N_9271,N_9454);
xor U9687 (N_9687,N_9429,N_9423);
xor U9688 (N_9688,N_9383,N_9394);
nor U9689 (N_9689,N_9361,N_9304);
nor U9690 (N_9690,N_9400,N_9479);
nand U9691 (N_9691,N_9419,N_9390);
and U9692 (N_9692,N_9360,N_9314);
xnor U9693 (N_9693,N_9395,N_9350);
or U9694 (N_9694,N_9352,N_9317);
or U9695 (N_9695,N_9465,N_9270);
nand U9696 (N_9696,N_9391,N_9428);
and U9697 (N_9697,N_9497,N_9457);
nand U9698 (N_9698,N_9282,N_9392);
xnor U9699 (N_9699,N_9291,N_9471);
xnor U9700 (N_9700,N_9405,N_9472);
nand U9701 (N_9701,N_9343,N_9355);
nand U9702 (N_9702,N_9373,N_9314);
xnor U9703 (N_9703,N_9297,N_9488);
nor U9704 (N_9704,N_9330,N_9347);
nand U9705 (N_9705,N_9403,N_9457);
or U9706 (N_9706,N_9398,N_9275);
and U9707 (N_9707,N_9264,N_9306);
or U9708 (N_9708,N_9457,N_9380);
nor U9709 (N_9709,N_9259,N_9366);
and U9710 (N_9710,N_9452,N_9293);
and U9711 (N_9711,N_9270,N_9434);
nand U9712 (N_9712,N_9416,N_9441);
or U9713 (N_9713,N_9413,N_9494);
nor U9714 (N_9714,N_9489,N_9322);
nor U9715 (N_9715,N_9355,N_9474);
or U9716 (N_9716,N_9462,N_9272);
and U9717 (N_9717,N_9433,N_9324);
and U9718 (N_9718,N_9430,N_9370);
and U9719 (N_9719,N_9482,N_9485);
xnor U9720 (N_9720,N_9251,N_9284);
and U9721 (N_9721,N_9265,N_9432);
nor U9722 (N_9722,N_9397,N_9265);
or U9723 (N_9723,N_9453,N_9262);
and U9724 (N_9724,N_9385,N_9424);
or U9725 (N_9725,N_9402,N_9325);
and U9726 (N_9726,N_9338,N_9419);
nor U9727 (N_9727,N_9353,N_9303);
and U9728 (N_9728,N_9448,N_9324);
nor U9729 (N_9729,N_9289,N_9279);
xor U9730 (N_9730,N_9492,N_9283);
nand U9731 (N_9731,N_9486,N_9433);
and U9732 (N_9732,N_9316,N_9368);
and U9733 (N_9733,N_9351,N_9446);
and U9734 (N_9734,N_9427,N_9443);
xnor U9735 (N_9735,N_9376,N_9466);
or U9736 (N_9736,N_9289,N_9396);
nand U9737 (N_9737,N_9411,N_9368);
nor U9738 (N_9738,N_9468,N_9324);
nor U9739 (N_9739,N_9403,N_9269);
nor U9740 (N_9740,N_9258,N_9321);
or U9741 (N_9741,N_9398,N_9421);
or U9742 (N_9742,N_9252,N_9410);
and U9743 (N_9743,N_9347,N_9337);
nor U9744 (N_9744,N_9426,N_9467);
or U9745 (N_9745,N_9372,N_9386);
nand U9746 (N_9746,N_9377,N_9401);
and U9747 (N_9747,N_9307,N_9495);
nor U9748 (N_9748,N_9390,N_9492);
nor U9749 (N_9749,N_9479,N_9274);
or U9750 (N_9750,N_9517,N_9663);
or U9751 (N_9751,N_9646,N_9658);
nor U9752 (N_9752,N_9672,N_9509);
nand U9753 (N_9753,N_9541,N_9733);
nor U9754 (N_9754,N_9745,N_9701);
xnor U9755 (N_9755,N_9749,N_9522);
xnor U9756 (N_9756,N_9603,N_9530);
xnor U9757 (N_9757,N_9724,N_9671);
and U9758 (N_9758,N_9702,N_9503);
and U9759 (N_9759,N_9566,N_9626);
xnor U9760 (N_9760,N_9620,N_9562);
and U9761 (N_9761,N_9698,N_9655);
and U9762 (N_9762,N_9568,N_9644);
nor U9763 (N_9763,N_9681,N_9582);
xor U9764 (N_9764,N_9673,N_9540);
nand U9765 (N_9765,N_9521,N_9678);
or U9766 (N_9766,N_9527,N_9700);
and U9767 (N_9767,N_9748,N_9533);
and U9768 (N_9768,N_9682,N_9504);
nand U9769 (N_9769,N_9537,N_9640);
xor U9770 (N_9770,N_9691,N_9597);
nor U9771 (N_9771,N_9532,N_9716);
and U9772 (N_9772,N_9624,N_9534);
xor U9773 (N_9773,N_9548,N_9727);
or U9774 (N_9774,N_9637,N_9580);
nor U9775 (N_9775,N_9747,N_9543);
or U9776 (N_9776,N_9561,N_9668);
nand U9777 (N_9777,N_9652,N_9667);
nor U9778 (N_9778,N_9669,N_9583);
xnor U9779 (N_9779,N_9546,N_9559);
or U9780 (N_9780,N_9606,N_9524);
nor U9781 (N_9781,N_9690,N_9730);
nand U9782 (N_9782,N_9677,N_9665);
or U9783 (N_9783,N_9571,N_9746);
xnor U9784 (N_9784,N_9557,N_9656);
nand U9785 (N_9785,N_9588,N_9511);
nor U9786 (N_9786,N_9704,N_9500);
and U9787 (N_9787,N_9577,N_9590);
xor U9788 (N_9788,N_9585,N_9601);
nand U9789 (N_9789,N_9515,N_9570);
and U9790 (N_9790,N_9505,N_9619);
nand U9791 (N_9791,N_9726,N_9565);
xnor U9792 (N_9792,N_9736,N_9607);
nand U9793 (N_9793,N_9661,N_9718);
and U9794 (N_9794,N_9573,N_9553);
xnor U9795 (N_9795,N_9508,N_9609);
nand U9796 (N_9796,N_9728,N_9636);
or U9797 (N_9797,N_9703,N_9654);
nand U9798 (N_9798,N_9621,N_9689);
nor U9799 (N_9799,N_9618,N_9518);
and U9800 (N_9800,N_9731,N_9735);
nor U9801 (N_9801,N_9639,N_9643);
xor U9802 (N_9802,N_9594,N_9596);
and U9803 (N_9803,N_9502,N_9611);
and U9804 (N_9804,N_9551,N_9513);
xor U9805 (N_9805,N_9717,N_9721);
or U9806 (N_9806,N_9734,N_9598);
nand U9807 (N_9807,N_9719,N_9653);
xnor U9808 (N_9808,N_9694,N_9666);
or U9809 (N_9809,N_9708,N_9629);
and U9810 (N_9810,N_9574,N_9520);
and U9811 (N_9811,N_9630,N_9514);
and U9812 (N_9812,N_9645,N_9507);
nor U9813 (N_9813,N_9531,N_9710);
or U9814 (N_9814,N_9638,N_9600);
xnor U9815 (N_9815,N_9528,N_9579);
and U9816 (N_9816,N_9506,N_9675);
and U9817 (N_9817,N_9576,N_9615);
or U9818 (N_9818,N_9737,N_9519);
nor U9819 (N_9819,N_9742,N_9592);
nor U9820 (N_9820,N_9558,N_9697);
nor U9821 (N_9821,N_9563,N_9720);
nand U9822 (N_9822,N_9623,N_9538);
nand U9823 (N_9823,N_9605,N_9512);
and U9824 (N_9824,N_9684,N_9581);
and U9825 (N_9825,N_9599,N_9612);
xnor U9826 (N_9826,N_9632,N_9591);
and U9827 (N_9827,N_9659,N_9587);
or U9828 (N_9828,N_9713,N_9622);
and U9829 (N_9829,N_9692,N_9712);
nand U9830 (N_9830,N_9569,N_9578);
nand U9831 (N_9831,N_9740,N_9683);
and U9832 (N_9832,N_9660,N_9529);
nand U9833 (N_9833,N_9613,N_9604);
or U9834 (N_9834,N_9523,N_9688);
xnor U9835 (N_9835,N_9705,N_9510);
xnor U9836 (N_9836,N_9739,N_9634);
or U9837 (N_9837,N_9550,N_9516);
xor U9838 (N_9838,N_9608,N_9633);
nand U9839 (N_9839,N_9709,N_9555);
or U9840 (N_9840,N_9547,N_9715);
xnor U9841 (N_9841,N_9575,N_9696);
nor U9842 (N_9842,N_9647,N_9536);
xnor U9843 (N_9843,N_9625,N_9586);
xnor U9844 (N_9844,N_9706,N_9679);
and U9845 (N_9845,N_9526,N_9725);
xor U9846 (N_9846,N_9544,N_9539);
or U9847 (N_9847,N_9693,N_9627);
nand U9848 (N_9848,N_9657,N_9602);
nand U9849 (N_9849,N_9649,N_9635);
xor U9850 (N_9850,N_9572,N_9593);
and U9851 (N_9851,N_9664,N_9545);
or U9852 (N_9852,N_9556,N_9628);
and U9853 (N_9853,N_9662,N_9589);
xnor U9854 (N_9854,N_9616,N_9617);
nor U9855 (N_9855,N_9567,N_9595);
or U9856 (N_9856,N_9642,N_9714);
and U9857 (N_9857,N_9584,N_9680);
xor U9858 (N_9858,N_9552,N_9542);
and U9859 (N_9859,N_9564,N_9722);
or U9860 (N_9860,N_9651,N_9707);
nand U9861 (N_9861,N_9650,N_9711);
and U9862 (N_9862,N_9695,N_9674);
nor U9863 (N_9863,N_9670,N_9648);
xnor U9864 (N_9864,N_9741,N_9729);
nor U9865 (N_9865,N_9676,N_9723);
xor U9866 (N_9866,N_9614,N_9686);
nor U9867 (N_9867,N_9641,N_9560);
nor U9868 (N_9868,N_9687,N_9501);
and U9869 (N_9869,N_9554,N_9610);
or U9870 (N_9870,N_9699,N_9732);
and U9871 (N_9871,N_9744,N_9685);
nor U9872 (N_9872,N_9738,N_9631);
and U9873 (N_9873,N_9743,N_9525);
xnor U9874 (N_9874,N_9535,N_9549);
and U9875 (N_9875,N_9706,N_9586);
nor U9876 (N_9876,N_9584,N_9636);
and U9877 (N_9877,N_9537,N_9677);
nand U9878 (N_9878,N_9672,N_9612);
or U9879 (N_9879,N_9591,N_9511);
nand U9880 (N_9880,N_9646,N_9733);
nand U9881 (N_9881,N_9681,N_9607);
nand U9882 (N_9882,N_9699,N_9564);
xnor U9883 (N_9883,N_9668,N_9587);
xor U9884 (N_9884,N_9560,N_9506);
nor U9885 (N_9885,N_9677,N_9560);
nand U9886 (N_9886,N_9685,N_9725);
xor U9887 (N_9887,N_9643,N_9681);
nand U9888 (N_9888,N_9705,N_9665);
and U9889 (N_9889,N_9544,N_9741);
or U9890 (N_9890,N_9560,N_9574);
nand U9891 (N_9891,N_9530,N_9565);
or U9892 (N_9892,N_9551,N_9573);
nor U9893 (N_9893,N_9684,N_9569);
nand U9894 (N_9894,N_9707,N_9741);
xor U9895 (N_9895,N_9664,N_9612);
and U9896 (N_9896,N_9582,N_9736);
nand U9897 (N_9897,N_9569,N_9738);
and U9898 (N_9898,N_9560,N_9686);
xor U9899 (N_9899,N_9731,N_9531);
and U9900 (N_9900,N_9575,N_9670);
and U9901 (N_9901,N_9585,N_9711);
nor U9902 (N_9902,N_9665,N_9528);
nand U9903 (N_9903,N_9707,N_9570);
xor U9904 (N_9904,N_9746,N_9702);
and U9905 (N_9905,N_9614,N_9598);
nand U9906 (N_9906,N_9566,N_9584);
nand U9907 (N_9907,N_9538,N_9574);
nor U9908 (N_9908,N_9703,N_9600);
and U9909 (N_9909,N_9728,N_9680);
nor U9910 (N_9910,N_9596,N_9718);
xor U9911 (N_9911,N_9696,N_9503);
nand U9912 (N_9912,N_9666,N_9647);
xor U9913 (N_9913,N_9686,N_9743);
xnor U9914 (N_9914,N_9699,N_9561);
or U9915 (N_9915,N_9733,N_9578);
nand U9916 (N_9916,N_9550,N_9623);
nor U9917 (N_9917,N_9616,N_9732);
and U9918 (N_9918,N_9705,N_9570);
nor U9919 (N_9919,N_9708,N_9616);
and U9920 (N_9920,N_9638,N_9681);
nor U9921 (N_9921,N_9681,N_9550);
nor U9922 (N_9922,N_9513,N_9606);
nor U9923 (N_9923,N_9717,N_9508);
and U9924 (N_9924,N_9686,N_9508);
xor U9925 (N_9925,N_9582,N_9629);
nand U9926 (N_9926,N_9546,N_9726);
or U9927 (N_9927,N_9644,N_9736);
nand U9928 (N_9928,N_9586,N_9698);
xor U9929 (N_9929,N_9510,N_9722);
or U9930 (N_9930,N_9622,N_9731);
xnor U9931 (N_9931,N_9648,N_9549);
or U9932 (N_9932,N_9628,N_9721);
and U9933 (N_9933,N_9718,N_9573);
nor U9934 (N_9934,N_9642,N_9683);
or U9935 (N_9935,N_9630,N_9719);
nand U9936 (N_9936,N_9706,N_9507);
or U9937 (N_9937,N_9674,N_9717);
or U9938 (N_9938,N_9688,N_9660);
xnor U9939 (N_9939,N_9614,N_9645);
nand U9940 (N_9940,N_9630,N_9747);
or U9941 (N_9941,N_9527,N_9563);
xnor U9942 (N_9942,N_9594,N_9665);
or U9943 (N_9943,N_9731,N_9638);
and U9944 (N_9944,N_9632,N_9596);
xnor U9945 (N_9945,N_9573,N_9622);
and U9946 (N_9946,N_9725,N_9744);
nor U9947 (N_9947,N_9531,N_9564);
and U9948 (N_9948,N_9657,N_9634);
xor U9949 (N_9949,N_9739,N_9675);
and U9950 (N_9950,N_9676,N_9514);
nand U9951 (N_9951,N_9639,N_9699);
or U9952 (N_9952,N_9706,N_9688);
xnor U9953 (N_9953,N_9677,N_9597);
or U9954 (N_9954,N_9728,N_9713);
or U9955 (N_9955,N_9729,N_9638);
xnor U9956 (N_9956,N_9651,N_9527);
nand U9957 (N_9957,N_9681,N_9738);
xnor U9958 (N_9958,N_9586,N_9576);
and U9959 (N_9959,N_9747,N_9661);
xnor U9960 (N_9960,N_9735,N_9549);
xor U9961 (N_9961,N_9562,N_9634);
nor U9962 (N_9962,N_9703,N_9719);
nor U9963 (N_9963,N_9673,N_9740);
nand U9964 (N_9964,N_9667,N_9587);
and U9965 (N_9965,N_9652,N_9747);
nor U9966 (N_9966,N_9741,N_9624);
or U9967 (N_9967,N_9674,N_9688);
nor U9968 (N_9968,N_9728,N_9500);
and U9969 (N_9969,N_9629,N_9602);
or U9970 (N_9970,N_9681,N_9570);
nand U9971 (N_9971,N_9699,N_9696);
and U9972 (N_9972,N_9589,N_9739);
nor U9973 (N_9973,N_9747,N_9507);
xor U9974 (N_9974,N_9590,N_9655);
and U9975 (N_9975,N_9553,N_9740);
nand U9976 (N_9976,N_9628,N_9713);
or U9977 (N_9977,N_9639,N_9558);
and U9978 (N_9978,N_9701,N_9525);
and U9979 (N_9979,N_9640,N_9649);
xnor U9980 (N_9980,N_9621,N_9732);
or U9981 (N_9981,N_9552,N_9561);
or U9982 (N_9982,N_9724,N_9571);
nand U9983 (N_9983,N_9634,N_9730);
xnor U9984 (N_9984,N_9637,N_9589);
xor U9985 (N_9985,N_9732,N_9531);
xnor U9986 (N_9986,N_9551,N_9733);
or U9987 (N_9987,N_9573,N_9586);
xnor U9988 (N_9988,N_9512,N_9684);
nor U9989 (N_9989,N_9546,N_9631);
xnor U9990 (N_9990,N_9717,N_9526);
xor U9991 (N_9991,N_9511,N_9565);
and U9992 (N_9992,N_9665,N_9507);
or U9993 (N_9993,N_9545,N_9623);
or U9994 (N_9994,N_9521,N_9577);
or U9995 (N_9995,N_9674,N_9731);
nand U9996 (N_9996,N_9538,N_9661);
nand U9997 (N_9997,N_9683,N_9731);
nand U9998 (N_9998,N_9675,N_9527);
and U9999 (N_9999,N_9593,N_9635);
or U10000 (N_10000,N_9854,N_9773);
or U10001 (N_10001,N_9870,N_9882);
or U10002 (N_10002,N_9762,N_9916);
nand U10003 (N_10003,N_9959,N_9878);
xor U10004 (N_10004,N_9956,N_9822);
xnor U10005 (N_10005,N_9847,N_9823);
and U10006 (N_10006,N_9883,N_9778);
and U10007 (N_10007,N_9753,N_9947);
nand U10008 (N_10008,N_9999,N_9902);
and U10009 (N_10009,N_9988,N_9989);
or U10010 (N_10010,N_9937,N_9760);
nor U10011 (N_10011,N_9794,N_9751);
nand U10012 (N_10012,N_9763,N_9871);
nand U10013 (N_10013,N_9820,N_9899);
and U10014 (N_10014,N_9780,N_9993);
nor U10015 (N_10015,N_9757,N_9833);
or U10016 (N_10016,N_9968,N_9926);
and U10017 (N_10017,N_9836,N_9818);
and U10018 (N_10018,N_9858,N_9786);
or U10019 (N_10019,N_9933,N_9979);
nand U10020 (N_10020,N_9888,N_9772);
nand U10021 (N_10021,N_9980,N_9853);
nand U10022 (N_10022,N_9891,N_9932);
or U10023 (N_10023,N_9811,N_9910);
xnor U10024 (N_10024,N_9759,N_9785);
nand U10025 (N_10025,N_9830,N_9941);
or U10026 (N_10026,N_9921,N_9974);
nand U10027 (N_10027,N_9943,N_9962);
and U10028 (N_10028,N_9879,N_9877);
or U10029 (N_10029,N_9815,N_9790);
or U10030 (N_10030,N_9797,N_9918);
and U10031 (N_10031,N_9783,N_9948);
xor U10032 (N_10032,N_9934,N_9881);
xor U10033 (N_10033,N_9982,N_9880);
nand U10034 (N_10034,N_9816,N_9840);
xnor U10035 (N_10035,N_9821,N_9834);
nor U10036 (N_10036,N_9890,N_9842);
nand U10037 (N_10037,N_9832,N_9867);
and U10038 (N_10038,N_9781,N_9915);
and U10039 (N_10039,N_9907,N_9776);
xnor U10040 (N_10040,N_9930,N_9784);
nand U10041 (N_10041,N_9896,N_9938);
nand U10042 (N_10042,N_9909,N_9805);
nor U10043 (N_10043,N_9807,N_9925);
or U10044 (N_10044,N_9875,N_9767);
nor U10045 (N_10045,N_9843,N_9813);
nand U10046 (N_10046,N_9755,N_9868);
or U10047 (N_10047,N_9895,N_9861);
nor U10048 (N_10048,N_9764,N_9801);
nand U10049 (N_10049,N_9750,N_9994);
and U10050 (N_10050,N_9928,N_9960);
nor U10051 (N_10051,N_9990,N_9985);
and U10052 (N_10052,N_9991,N_9965);
and U10053 (N_10053,N_9791,N_9768);
xnor U10054 (N_10054,N_9898,N_9946);
nor U10055 (N_10055,N_9793,N_9939);
nand U10056 (N_10056,N_9856,N_9919);
nor U10057 (N_10057,N_9942,N_9796);
or U10058 (N_10058,N_9957,N_9998);
nor U10059 (N_10059,N_9849,N_9864);
and U10060 (N_10060,N_9809,N_9971);
nand U10061 (N_10061,N_9771,N_9931);
and U10062 (N_10062,N_9903,N_9792);
and U10063 (N_10063,N_9802,N_9770);
xor U10064 (N_10064,N_9826,N_9752);
and U10065 (N_10065,N_9936,N_9819);
and U10066 (N_10066,N_9817,N_9954);
xor U10067 (N_10067,N_9827,N_9837);
xnor U10068 (N_10068,N_9812,N_9754);
nor U10069 (N_10069,N_9824,N_9997);
xor U10070 (N_10070,N_9913,N_9970);
nand U10071 (N_10071,N_9857,N_9917);
nand U10072 (N_10072,N_9782,N_9855);
nand U10073 (N_10073,N_9844,N_9944);
nand U10074 (N_10074,N_9775,N_9838);
xor U10075 (N_10075,N_9955,N_9886);
nand U10076 (N_10076,N_9872,N_9927);
nand U10077 (N_10077,N_9992,N_9798);
nand U10078 (N_10078,N_9981,N_9774);
xor U10079 (N_10079,N_9884,N_9978);
or U10080 (N_10080,N_9779,N_9995);
and U10081 (N_10081,N_9924,N_9841);
and U10082 (N_10082,N_9846,N_9977);
nand U10083 (N_10083,N_9758,N_9845);
nand U10084 (N_10084,N_9969,N_9923);
xor U10085 (N_10085,N_9967,N_9761);
nor U10086 (N_10086,N_9894,N_9869);
or U10087 (N_10087,N_9808,N_9987);
nor U10088 (N_10088,N_9859,N_9950);
nand U10089 (N_10089,N_9766,N_9922);
or U10090 (N_10090,N_9862,N_9892);
xor U10091 (N_10091,N_9803,N_9789);
or U10092 (N_10092,N_9804,N_9828);
and U10093 (N_10093,N_9951,N_9865);
nand U10094 (N_10094,N_9839,N_9874);
and U10095 (N_10095,N_9945,N_9848);
xor U10096 (N_10096,N_9952,N_9860);
and U10097 (N_10097,N_9873,N_9831);
xor U10098 (N_10098,N_9966,N_9975);
and U10099 (N_10099,N_9893,N_9887);
xnor U10100 (N_10100,N_9889,N_9863);
and U10101 (N_10101,N_9905,N_9799);
xor U10102 (N_10102,N_9973,N_9900);
or U10103 (N_10103,N_9829,N_9914);
nor U10104 (N_10104,N_9963,N_9906);
nor U10105 (N_10105,N_9935,N_9787);
or U10106 (N_10106,N_9949,N_9825);
and U10107 (N_10107,N_9912,N_9929);
nor U10108 (N_10108,N_9835,N_9814);
nand U10109 (N_10109,N_9800,N_9806);
or U10110 (N_10110,N_9852,N_9911);
or U10111 (N_10111,N_9940,N_9777);
and U10112 (N_10112,N_9953,N_9765);
and U10113 (N_10113,N_9972,N_9996);
or U10114 (N_10114,N_9769,N_9986);
xnor U10115 (N_10115,N_9795,N_9984);
and U10116 (N_10116,N_9851,N_9961);
nand U10117 (N_10117,N_9876,N_9908);
nor U10118 (N_10118,N_9756,N_9788);
nand U10119 (N_10119,N_9866,N_9904);
or U10120 (N_10120,N_9964,N_9810);
nand U10121 (N_10121,N_9850,N_9958);
and U10122 (N_10122,N_9983,N_9920);
and U10123 (N_10123,N_9976,N_9897);
or U10124 (N_10124,N_9901,N_9885);
or U10125 (N_10125,N_9891,N_9791);
xor U10126 (N_10126,N_9917,N_9840);
and U10127 (N_10127,N_9945,N_9908);
nor U10128 (N_10128,N_9808,N_9779);
and U10129 (N_10129,N_9899,N_9788);
xnor U10130 (N_10130,N_9856,N_9923);
nand U10131 (N_10131,N_9949,N_9968);
and U10132 (N_10132,N_9808,N_9958);
or U10133 (N_10133,N_9989,N_9985);
or U10134 (N_10134,N_9851,N_9960);
and U10135 (N_10135,N_9795,N_9983);
or U10136 (N_10136,N_9866,N_9775);
or U10137 (N_10137,N_9882,N_9911);
xnor U10138 (N_10138,N_9820,N_9910);
or U10139 (N_10139,N_9841,N_9773);
and U10140 (N_10140,N_9848,N_9920);
nor U10141 (N_10141,N_9793,N_9969);
or U10142 (N_10142,N_9864,N_9844);
or U10143 (N_10143,N_9871,N_9901);
nor U10144 (N_10144,N_9984,N_9841);
or U10145 (N_10145,N_9947,N_9930);
and U10146 (N_10146,N_9808,N_9863);
nor U10147 (N_10147,N_9881,N_9786);
nor U10148 (N_10148,N_9954,N_9808);
xor U10149 (N_10149,N_9890,N_9780);
nand U10150 (N_10150,N_9788,N_9762);
nand U10151 (N_10151,N_9790,N_9908);
nand U10152 (N_10152,N_9977,N_9947);
xor U10153 (N_10153,N_9915,N_9991);
xnor U10154 (N_10154,N_9810,N_9996);
and U10155 (N_10155,N_9796,N_9916);
nor U10156 (N_10156,N_9870,N_9791);
or U10157 (N_10157,N_9851,N_9874);
nor U10158 (N_10158,N_9839,N_9761);
nor U10159 (N_10159,N_9977,N_9959);
xor U10160 (N_10160,N_9867,N_9774);
and U10161 (N_10161,N_9856,N_9956);
or U10162 (N_10162,N_9929,N_9905);
nand U10163 (N_10163,N_9756,N_9891);
and U10164 (N_10164,N_9815,N_9769);
and U10165 (N_10165,N_9779,N_9752);
nor U10166 (N_10166,N_9833,N_9911);
or U10167 (N_10167,N_9861,N_9791);
and U10168 (N_10168,N_9953,N_9922);
and U10169 (N_10169,N_9946,N_9951);
nor U10170 (N_10170,N_9751,N_9906);
xor U10171 (N_10171,N_9968,N_9783);
xnor U10172 (N_10172,N_9761,N_9961);
nor U10173 (N_10173,N_9787,N_9989);
or U10174 (N_10174,N_9975,N_9897);
and U10175 (N_10175,N_9842,N_9949);
and U10176 (N_10176,N_9900,N_9916);
xnor U10177 (N_10177,N_9982,N_9779);
nand U10178 (N_10178,N_9753,N_9757);
nor U10179 (N_10179,N_9863,N_9829);
nand U10180 (N_10180,N_9848,N_9975);
and U10181 (N_10181,N_9971,N_9764);
or U10182 (N_10182,N_9948,N_9907);
nor U10183 (N_10183,N_9877,N_9757);
xor U10184 (N_10184,N_9777,N_9842);
or U10185 (N_10185,N_9969,N_9869);
xor U10186 (N_10186,N_9973,N_9905);
nand U10187 (N_10187,N_9894,N_9780);
xor U10188 (N_10188,N_9968,N_9833);
nand U10189 (N_10189,N_9885,N_9992);
xor U10190 (N_10190,N_9813,N_9788);
or U10191 (N_10191,N_9766,N_9971);
nand U10192 (N_10192,N_9846,N_9901);
nand U10193 (N_10193,N_9986,N_9890);
and U10194 (N_10194,N_9988,N_9805);
or U10195 (N_10195,N_9762,N_9946);
or U10196 (N_10196,N_9875,N_9855);
and U10197 (N_10197,N_9877,N_9804);
or U10198 (N_10198,N_9914,N_9841);
nand U10199 (N_10199,N_9922,N_9885);
nor U10200 (N_10200,N_9893,N_9957);
or U10201 (N_10201,N_9992,N_9838);
and U10202 (N_10202,N_9852,N_9896);
or U10203 (N_10203,N_9967,N_9877);
xnor U10204 (N_10204,N_9750,N_9893);
and U10205 (N_10205,N_9847,N_9828);
or U10206 (N_10206,N_9765,N_9783);
or U10207 (N_10207,N_9752,N_9965);
or U10208 (N_10208,N_9969,N_9802);
xor U10209 (N_10209,N_9823,N_9994);
nor U10210 (N_10210,N_9869,N_9847);
nor U10211 (N_10211,N_9914,N_9882);
nor U10212 (N_10212,N_9939,N_9841);
nor U10213 (N_10213,N_9913,N_9764);
xor U10214 (N_10214,N_9916,N_9961);
nor U10215 (N_10215,N_9970,N_9944);
or U10216 (N_10216,N_9761,N_9809);
and U10217 (N_10217,N_9760,N_9849);
nand U10218 (N_10218,N_9896,N_9768);
nor U10219 (N_10219,N_9945,N_9924);
xnor U10220 (N_10220,N_9803,N_9754);
nor U10221 (N_10221,N_9822,N_9996);
nand U10222 (N_10222,N_9885,N_9840);
xor U10223 (N_10223,N_9798,N_9967);
nor U10224 (N_10224,N_9898,N_9781);
nor U10225 (N_10225,N_9808,N_9786);
nand U10226 (N_10226,N_9944,N_9948);
xnor U10227 (N_10227,N_9909,N_9939);
xor U10228 (N_10228,N_9915,N_9914);
and U10229 (N_10229,N_9938,N_9840);
nand U10230 (N_10230,N_9970,N_9846);
nor U10231 (N_10231,N_9991,N_9879);
or U10232 (N_10232,N_9946,N_9776);
nor U10233 (N_10233,N_9855,N_9969);
nor U10234 (N_10234,N_9800,N_9989);
xor U10235 (N_10235,N_9847,N_9954);
nor U10236 (N_10236,N_9919,N_9830);
nand U10237 (N_10237,N_9959,N_9834);
nand U10238 (N_10238,N_9894,N_9820);
and U10239 (N_10239,N_9985,N_9861);
or U10240 (N_10240,N_9983,N_9934);
and U10241 (N_10241,N_9910,N_9880);
nor U10242 (N_10242,N_9885,N_9958);
and U10243 (N_10243,N_9831,N_9807);
xor U10244 (N_10244,N_9947,N_9982);
or U10245 (N_10245,N_9978,N_9791);
xnor U10246 (N_10246,N_9989,N_9885);
or U10247 (N_10247,N_9838,N_9999);
or U10248 (N_10248,N_9759,N_9960);
nand U10249 (N_10249,N_9771,N_9898);
and U10250 (N_10250,N_10075,N_10093);
nor U10251 (N_10251,N_10237,N_10087);
xnor U10252 (N_10252,N_10103,N_10069);
xnor U10253 (N_10253,N_10105,N_10243);
nor U10254 (N_10254,N_10097,N_10008);
and U10255 (N_10255,N_10231,N_10193);
xor U10256 (N_10256,N_10106,N_10113);
xnor U10257 (N_10257,N_10187,N_10016);
nor U10258 (N_10258,N_10023,N_10025);
xor U10259 (N_10259,N_10125,N_10140);
nand U10260 (N_10260,N_10027,N_10213);
or U10261 (N_10261,N_10041,N_10145);
xnor U10262 (N_10262,N_10038,N_10164);
or U10263 (N_10263,N_10067,N_10055);
nor U10264 (N_10264,N_10096,N_10206);
and U10265 (N_10265,N_10168,N_10084);
nor U10266 (N_10266,N_10163,N_10198);
nand U10267 (N_10267,N_10200,N_10066);
or U10268 (N_10268,N_10162,N_10175);
xnor U10269 (N_10269,N_10049,N_10021);
nor U10270 (N_10270,N_10158,N_10020);
or U10271 (N_10271,N_10030,N_10060);
xnor U10272 (N_10272,N_10121,N_10144);
or U10273 (N_10273,N_10141,N_10234);
and U10274 (N_10274,N_10160,N_10005);
nor U10275 (N_10275,N_10058,N_10159);
or U10276 (N_10276,N_10204,N_10090);
or U10277 (N_10277,N_10152,N_10189);
or U10278 (N_10278,N_10249,N_10068);
nor U10279 (N_10279,N_10195,N_10071);
and U10280 (N_10280,N_10239,N_10235);
xor U10281 (N_10281,N_10129,N_10135);
or U10282 (N_10282,N_10029,N_10228);
xor U10283 (N_10283,N_10173,N_10079);
xnor U10284 (N_10284,N_10050,N_10196);
or U10285 (N_10285,N_10024,N_10065);
or U10286 (N_10286,N_10039,N_10004);
nand U10287 (N_10287,N_10156,N_10186);
or U10288 (N_10288,N_10150,N_10057);
and U10289 (N_10289,N_10081,N_10224);
and U10290 (N_10290,N_10114,N_10092);
nand U10291 (N_10291,N_10136,N_10147);
nand U10292 (N_10292,N_10244,N_10146);
nand U10293 (N_10293,N_10083,N_10155);
or U10294 (N_10294,N_10107,N_10233);
or U10295 (N_10295,N_10210,N_10044);
or U10296 (N_10296,N_10077,N_10190);
nand U10297 (N_10297,N_10133,N_10192);
and U10298 (N_10298,N_10072,N_10010);
nand U10299 (N_10299,N_10054,N_10127);
xnor U10300 (N_10300,N_10174,N_10085);
or U10301 (N_10301,N_10101,N_10171);
nor U10302 (N_10302,N_10134,N_10240);
xor U10303 (N_10303,N_10139,N_10132);
nor U10304 (N_10304,N_10091,N_10003);
nor U10305 (N_10305,N_10178,N_10184);
or U10306 (N_10306,N_10241,N_10033);
and U10307 (N_10307,N_10169,N_10166);
nor U10308 (N_10308,N_10154,N_10080);
xnor U10309 (N_10309,N_10056,N_10007);
xnor U10310 (N_10310,N_10046,N_10130);
or U10311 (N_10311,N_10078,N_10167);
nand U10312 (N_10312,N_10109,N_10032);
xnor U10313 (N_10313,N_10245,N_10119);
or U10314 (N_10314,N_10104,N_10151);
xnor U10315 (N_10315,N_10036,N_10179);
nand U10316 (N_10316,N_10165,N_10073);
or U10317 (N_10317,N_10001,N_10061);
nand U10318 (N_10318,N_10170,N_10100);
and U10319 (N_10319,N_10099,N_10000);
nor U10320 (N_10320,N_10161,N_10042);
nor U10321 (N_10321,N_10223,N_10123);
and U10322 (N_10322,N_10076,N_10126);
nor U10323 (N_10323,N_10182,N_10110);
and U10324 (N_10324,N_10172,N_10018);
nor U10325 (N_10325,N_10181,N_10118);
and U10326 (N_10326,N_10070,N_10086);
nand U10327 (N_10327,N_10225,N_10214);
and U10328 (N_10328,N_10216,N_10082);
or U10329 (N_10329,N_10040,N_10219);
or U10330 (N_10330,N_10246,N_10131);
xnor U10331 (N_10331,N_10052,N_10211);
xnor U10332 (N_10332,N_10188,N_10115);
and U10333 (N_10333,N_10063,N_10236);
xnor U10334 (N_10334,N_10035,N_10051);
xor U10335 (N_10335,N_10197,N_10124);
nor U10336 (N_10336,N_10026,N_10138);
xor U10337 (N_10337,N_10203,N_10009);
or U10338 (N_10338,N_10202,N_10111);
or U10339 (N_10339,N_10013,N_10015);
nor U10340 (N_10340,N_10102,N_10122);
or U10341 (N_10341,N_10226,N_10117);
nor U10342 (N_10342,N_10053,N_10221);
nand U10343 (N_10343,N_10017,N_10014);
or U10344 (N_10344,N_10180,N_10095);
nand U10345 (N_10345,N_10227,N_10012);
nand U10346 (N_10346,N_10208,N_10209);
xor U10347 (N_10347,N_10048,N_10185);
or U10348 (N_10348,N_10232,N_10176);
or U10349 (N_10349,N_10220,N_10137);
and U10350 (N_10350,N_10059,N_10183);
xor U10351 (N_10351,N_10002,N_10212);
nand U10352 (N_10352,N_10037,N_10098);
and U10353 (N_10353,N_10205,N_10230);
and U10354 (N_10354,N_10148,N_10088);
and U10355 (N_10355,N_10128,N_10142);
xor U10356 (N_10356,N_10064,N_10112);
or U10357 (N_10357,N_10011,N_10022);
nand U10358 (N_10358,N_10215,N_10108);
nor U10359 (N_10359,N_10194,N_10043);
or U10360 (N_10360,N_10201,N_10222);
and U10361 (N_10361,N_10019,N_10149);
xor U10362 (N_10362,N_10062,N_10047);
xor U10363 (N_10363,N_10242,N_10045);
nand U10364 (N_10364,N_10177,N_10143);
nor U10365 (N_10365,N_10120,N_10074);
nand U10366 (N_10366,N_10031,N_10248);
nand U10367 (N_10367,N_10247,N_10191);
nand U10368 (N_10368,N_10028,N_10199);
or U10369 (N_10369,N_10094,N_10207);
nand U10370 (N_10370,N_10157,N_10153);
xnor U10371 (N_10371,N_10218,N_10116);
nand U10372 (N_10372,N_10229,N_10217);
nand U10373 (N_10373,N_10089,N_10034);
nor U10374 (N_10374,N_10006,N_10238);
or U10375 (N_10375,N_10058,N_10248);
or U10376 (N_10376,N_10169,N_10122);
xor U10377 (N_10377,N_10120,N_10085);
nand U10378 (N_10378,N_10112,N_10106);
nand U10379 (N_10379,N_10156,N_10008);
nor U10380 (N_10380,N_10018,N_10202);
and U10381 (N_10381,N_10103,N_10216);
xor U10382 (N_10382,N_10029,N_10171);
or U10383 (N_10383,N_10117,N_10044);
nor U10384 (N_10384,N_10127,N_10114);
xor U10385 (N_10385,N_10143,N_10169);
xor U10386 (N_10386,N_10138,N_10104);
nor U10387 (N_10387,N_10000,N_10188);
xor U10388 (N_10388,N_10048,N_10047);
or U10389 (N_10389,N_10021,N_10112);
nand U10390 (N_10390,N_10021,N_10134);
or U10391 (N_10391,N_10219,N_10130);
and U10392 (N_10392,N_10205,N_10079);
nor U10393 (N_10393,N_10036,N_10008);
nand U10394 (N_10394,N_10075,N_10076);
nor U10395 (N_10395,N_10228,N_10018);
and U10396 (N_10396,N_10227,N_10102);
xor U10397 (N_10397,N_10067,N_10241);
xor U10398 (N_10398,N_10192,N_10234);
and U10399 (N_10399,N_10201,N_10217);
nand U10400 (N_10400,N_10213,N_10204);
or U10401 (N_10401,N_10059,N_10225);
nor U10402 (N_10402,N_10206,N_10195);
or U10403 (N_10403,N_10198,N_10084);
nand U10404 (N_10404,N_10102,N_10056);
nor U10405 (N_10405,N_10074,N_10062);
or U10406 (N_10406,N_10103,N_10114);
and U10407 (N_10407,N_10033,N_10031);
or U10408 (N_10408,N_10241,N_10238);
or U10409 (N_10409,N_10172,N_10219);
nor U10410 (N_10410,N_10034,N_10102);
or U10411 (N_10411,N_10244,N_10147);
xnor U10412 (N_10412,N_10070,N_10089);
nor U10413 (N_10413,N_10232,N_10105);
xnor U10414 (N_10414,N_10047,N_10103);
or U10415 (N_10415,N_10106,N_10226);
nor U10416 (N_10416,N_10235,N_10047);
nand U10417 (N_10417,N_10131,N_10008);
xor U10418 (N_10418,N_10061,N_10236);
and U10419 (N_10419,N_10173,N_10156);
or U10420 (N_10420,N_10222,N_10033);
and U10421 (N_10421,N_10039,N_10082);
nand U10422 (N_10422,N_10005,N_10001);
nor U10423 (N_10423,N_10182,N_10027);
nor U10424 (N_10424,N_10032,N_10098);
nand U10425 (N_10425,N_10164,N_10147);
or U10426 (N_10426,N_10206,N_10036);
nor U10427 (N_10427,N_10043,N_10150);
and U10428 (N_10428,N_10112,N_10114);
xor U10429 (N_10429,N_10168,N_10054);
nor U10430 (N_10430,N_10138,N_10238);
nor U10431 (N_10431,N_10232,N_10200);
nand U10432 (N_10432,N_10084,N_10100);
or U10433 (N_10433,N_10149,N_10063);
nand U10434 (N_10434,N_10195,N_10089);
nor U10435 (N_10435,N_10200,N_10211);
and U10436 (N_10436,N_10148,N_10146);
nor U10437 (N_10437,N_10049,N_10169);
or U10438 (N_10438,N_10015,N_10078);
nand U10439 (N_10439,N_10212,N_10145);
or U10440 (N_10440,N_10203,N_10200);
and U10441 (N_10441,N_10125,N_10050);
and U10442 (N_10442,N_10184,N_10169);
and U10443 (N_10443,N_10022,N_10210);
and U10444 (N_10444,N_10207,N_10178);
xnor U10445 (N_10445,N_10206,N_10196);
or U10446 (N_10446,N_10158,N_10150);
nand U10447 (N_10447,N_10072,N_10040);
xor U10448 (N_10448,N_10049,N_10243);
and U10449 (N_10449,N_10129,N_10070);
xor U10450 (N_10450,N_10153,N_10038);
nor U10451 (N_10451,N_10142,N_10016);
and U10452 (N_10452,N_10187,N_10163);
and U10453 (N_10453,N_10110,N_10237);
xnor U10454 (N_10454,N_10169,N_10146);
and U10455 (N_10455,N_10244,N_10187);
nand U10456 (N_10456,N_10112,N_10169);
and U10457 (N_10457,N_10247,N_10089);
nor U10458 (N_10458,N_10163,N_10220);
nand U10459 (N_10459,N_10248,N_10216);
and U10460 (N_10460,N_10060,N_10194);
nand U10461 (N_10461,N_10073,N_10245);
and U10462 (N_10462,N_10018,N_10125);
and U10463 (N_10463,N_10178,N_10077);
or U10464 (N_10464,N_10007,N_10006);
or U10465 (N_10465,N_10074,N_10059);
and U10466 (N_10466,N_10224,N_10229);
xor U10467 (N_10467,N_10052,N_10070);
xor U10468 (N_10468,N_10153,N_10019);
nand U10469 (N_10469,N_10124,N_10021);
or U10470 (N_10470,N_10030,N_10049);
nor U10471 (N_10471,N_10228,N_10188);
xnor U10472 (N_10472,N_10027,N_10101);
or U10473 (N_10473,N_10079,N_10004);
or U10474 (N_10474,N_10211,N_10240);
or U10475 (N_10475,N_10232,N_10111);
xnor U10476 (N_10476,N_10007,N_10068);
or U10477 (N_10477,N_10198,N_10050);
nand U10478 (N_10478,N_10135,N_10222);
nand U10479 (N_10479,N_10235,N_10042);
nor U10480 (N_10480,N_10100,N_10104);
xor U10481 (N_10481,N_10024,N_10114);
nor U10482 (N_10482,N_10138,N_10012);
or U10483 (N_10483,N_10066,N_10044);
nor U10484 (N_10484,N_10131,N_10018);
nor U10485 (N_10485,N_10000,N_10194);
nor U10486 (N_10486,N_10155,N_10115);
nor U10487 (N_10487,N_10217,N_10181);
xor U10488 (N_10488,N_10235,N_10143);
xnor U10489 (N_10489,N_10179,N_10065);
xor U10490 (N_10490,N_10125,N_10130);
or U10491 (N_10491,N_10136,N_10146);
nor U10492 (N_10492,N_10165,N_10206);
and U10493 (N_10493,N_10045,N_10015);
nor U10494 (N_10494,N_10009,N_10045);
nor U10495 (N_10495,N_10240,N_10248);
nand U10496 (N_10496,N_10089,N_10147);
or U10497 (N_10497,N_10187,N_10237);
nor U10498 (N_10498,N_10206,N_10090);
nand U10499 (N_10499,N_10237,N_10019);
nand U10500 (N_10500,N_10489,N_10468);
xor U10501 (N_10501,N_10443,N_10483);
xor U10502 (N_10502,N_10314,N_10261);
nor U10503 (N_10503,N_10465,N_10356);
nand U10504 (N_10504,N_10300,N_10448);
or U10505 (N_10505,N_10394,N_10321);
nand U10506 (N_10506,N_10334,N_10382);
xor U10507 (N_10507,N_10464,N_10326);
xor U10508 (N_10508,N_10404,N_10350);
nand U10509 (N_10509,N_10390,N_10376);
and U10510 (N_10510,N_10458,N_10446);
nand U10511 (N_10511,N_10269,N_10330);
or U10512 (N_10512,N_10267,N_10408);
or U10513 (N_10513,N_10431,N_10413);
nor U10514 (N_10514,N_10459,N_10405);
and U10515 (N_10515,N_10371,N_10438);
nor U10516 (N_10516,N_10332,N_10393);
nor U10517 (N_10517,N_10399,N_10362);
or U10518 (N_10518,N_10481,N_10425);
nor U10519 (N_10519,N_10339,N_10329);
or U10520 (N_10520,N_10265,N_10336);
and U10521 (N_10521,N_10412,N_10328);
and U10522 (N_10522,N_10259,N_10319);
nand U10523 (N_10523,N_10427,N_10294);
nor U10524 (N_10524,N_10355,N_10273);
and U10525 (N_10525,N_10411,N_10450);
or U10526 (N_10526,N_10307,N_10485);
or U10527 (N_10527,N_10287,N_10442);
xnor U10528 (N_10528,N_10434,N_10260);
and U10529 (N_10529,N_10291,N_10370);
or U10530 (N_10530,N_10445,N_10272);
nand U10531 (N_10531,N_10423,N_10263);
or U10532 (N_10532,N_10324,N_10388);
xor U10533 (N_10533,N_10387,N_10478);
nor U10534 (N_10534,N_10360,N_10416);
nand U10535 (N_10535,N_10354,N_10415);
nand U10536 (N_10536,N_10286,N_10447);
nand U10537 (N_10537,N_10302,N_10398);
nand U10538 (N_10538,N_10374,N_10397);
and U10539 (N_10539,N_10357,N_10365);
or U10540 (N_10540,N_10496,N_10422);
or U10541 (N_10541,N_10395,N_10424);
xor U10542 (N_10542,N_10317,N_10497);
nor U10543 (N_10543,N_10476,N_10407);
nand U10544 (N_10544,N_10344,N_10296);
xor U10545 (N_10545,N_10322,N_10274);
xor U10546 (N_10546,N_10375,N_10310);
nand U10547 (N_10547,N_10392,N_10313);
nand U10548 (N_10548,N_10472,N_10482);
nand U10549 (N_10549,N_10460,N_10479);
xor U10550 (N_10550,N_10396,N_10435);
nand U10551 (N_10551,N_10299,N_10305);
nand U10552 (N_10552,N_10403,N_10283);
or U10553 (N_10553,N_10301,N_10323);
nand U10554 (N_10554,N_10421,N_10311);
nand U10555 (N_10555,N_10297,N_10280);
nand U10556 (N_10556,N_10469,N_10417);
nand U10557 (N_10557,N_10380,N_10312);
nor U10558 (N_10558,N_10252,N_10488);
nand U10559 (N_10559,N_10277,N_10409);
xor U10560 (N_10560,N_10281,N_10359);
nand U10561 (N_10561,N_10251,N_10491);
and U10562 (N_10562,N_10257,N_10318);
nor U10563 (N_10563,N_10303,N_10391);
nand U10564 (N_10564,N_10298,N_10254);
nor U10565 (N_10565,N_10270,N_10320);
xnor U10566 (N_10566,N_10414,N_10499);
or U10567 (N_10567,N_10293,N_10340);
nand U10568 (N_10568,N_10406,N_10255);
nand U10569 (N_10569,N_10428,N_10351);
nor U10570 (N_10570,N_10295,N_10377);
xor U10571 (N_10571,N_10282,N_10361);
or U10572 (N_10572,N_10401,N_10256);
nand U10573 (N_10573,N_10429,N_10418);
xnor U10574 (N_10574,N_10366,N_10315);
nand U10575 (N_10575,N_10343,N_10471);
nand U10576 (N_10576,N_10470,N_10495);
or U10577 (N_10577,N_10333,N_10342);
and U10578 (N_10578,N_10304,N_10266);
or U10579 (N_10579,N_10289,N_10346);
or U10580 (N_10580,N_10379,N_10466);
nand U10581 (N_10581,N_10341,N_10275);
and U10582 (N_10582,N_10383,N_10347);
or U10583 (N_10583,N_10327,N_10452);
nand U10584 (N_10584,N_10419,N_10473);
nand U10585 (N_10585,N_10349,N_10290);
xnor U10586 (N_10586,N_10439,N_10335);
or U10587 (N_10587,N_10258,N_10386);
or U10588 (N_10588,N_10353,N_10306);
xnor U10589 (N_10589,N_10250,N_10480);
and U10590 (N_10590,N_10378,N_10331);
xor U10591 (N_10591,N_10288,N_10278);
nand U10592 (N_10592,N_10348,N_10264);
nor U10593 (N_10593,N_10437,N_10451);
nor U10594 (N_10594,N_10279,N_10487);
and U10595 (N_10595,N_10454,N_10308);
nor U10596 (N_10596,N_10440,N_10292);
or U10597 (N_10597,N_10433,N_10345);
nand U10598 (N_10598,N_10352,N_10337);
nor U10599 (N_10599,N_10364,N_10463);
nand U10600 (N_10600,N_10436,N_10363);
or U10601 (N_10601,N_10367,N_10325);
nand U10602 (N_10602,N_10309,N_10284);
nor U10603 (N_10603,N_10372,N_10493);
nand U10604 (N_10604,N_10368,N_10316);
and U10605 (N_10605,N_10444,N_10456);
nand U10606 (N_10606,N_10271,N_10369);
nor U10607 (N_10607,N_10490,N_10381);
and U10608 (N_10608,N_10338,N_10426);
or U10609 (N_10609,N_10432,N_10268);
xnor U10610 (N_10610,N_10384,N_10498);
nand U10611 (N_10611,N_10477,N_10253);
xnor U10612 (N_10612,N_10475,N_10373);
and U10613 (N_10613,N_10285,N_10461);
xor U10614 (N_10614,N_10358,N_10467);
nand U10615 (N_10615,N_10457,N_10453);
nand U10616 (N_10616,N_10276,N_10494);
and U10617 (N_10617,N_10262,N_10385);
xnor U10618 (N_10618,N_10462,N_10402);
nand U10619 (N_10619,N_10486,N_10492);
or U10620 (N_10620,N_10474,N_10441);
xor U10621 (N_10621,N_10400,N_10455);
and U10622 (N_10622,N_10430,N_10420);
and U10623 (N_10623,N_10449,N_10389);
and U10624 (N_10624,N_10484,N_10410);
and U10625 (N_10625,N_10485,N_10315);
xnor U10626 (N_10626,N_10466,N_10432);
xor U10627 (N_10627,N_10292,N_10448);
xnor U10628 (N_10628,N_10440,N_10359);
nand U10629 (N_10629,N_10292,N_10427);
nor U10630 (N_10630,N_10270,N_10328);
and U10631 (N_10631,N_10313,N_10370);
nor U10632 (N_10632,N_10329,N_10286);
nor U10633 (N_10633,N_10425,N_10361);
and U10634 (N_10634,N_10415,N_10343);
or U10635 (N_10635,N_10387,N_10452);
nor U10636 (N_10636,N_10325,N_10292);
xor U10637 (N_10637,N_10346,N_10394);
xor U10638 (N_10638,N_10394,N_10400);
xor U10639 (N_10639,N_10307,N_10384);
or U10640 (N_10640,N_10427,N_10385);
or U10641 (N_10641,N_10285,N_10431);
nor U10642 (N_10642,N_10466,N_10386);
nand U10643 (N_10643,N_10282,N_10310);
xnor U10644 (N_10644,N_10478,N_10359);
and U10645 (N_10645,N_10261,N_10410);
or U10646 (N_10646,N_10377,N_10404);
xor U10647 (N_10647,N_10316,N_10330);
nand U10648 (N_10648,N_10408,N_10288);
and U10649 (N_10649,N_10466,N_10408);
or U10650 (N_10650,N_10299,N_10416);
nand U10651 (N_10651,N_10293,N_10294);
xnor U10652 (N_10652,N_10468,N_10450);
nor U10653 (N_10653,N_10435,N_10366);
and U10654 (N_10654,N_10389,N_10400);
nor U10655 (N_10655,N_10386,N_10401);
xor U10656 (N_10656,N_10352,N_10475);
nor U10657 (N_10657,N_10326,N_10395);
xor U10658 (N_10658,N_10470,N_10440);
xnor U10659 (N_10659,N_10309,N_10459);
xnor U10660 (N_10660,N_10258,N_10277);
or U10661 (N_10661,N_10489,N_10288);
nor U10662 (N_10662,N_10262,N_10481);
xor U10663 (N_10663,N_10433,N_10370);
or U10664 (N_10664,N_10413,N_10331);
and U10665 (N_10665,N_10344,N_10479);
nor U10666 (N_10666,N_10435,N_10383);
and U10667 (N_10667,N_10463,N_10388);
nor U10668 (N_10668,N_10455,N_10404);
and U10669 (N_10669,N_10317,N_10492);
nor U10670 (N_10670,N_10422,N_10327);
or U10671 (N_10671,N_10492,N_10371);
xor U10672 (N_10672,N_10342,N_10360);
nor U10673 (N_10673,N_10497,N_10478);
and U10674 (N_10674,N_10395,N_10338);
nand U10675 (N_10675,N_10458,N_10433);
nand U10676 (N_10676,N_10330,N_10459);
and U10677 (N_10677,N_10338,N_10258);
or U10678 (N_10678,N_10321,N_10485);
xnor U10679 (N_10679,N_10316,N_10289);
nand U10680 (N_10680,N_10257,N_10389);
xor U10681 (N_10681,N_10467,N_10426);
xor U10682 (N_10682,N_10412,N_10435);
xnor U10683 (N_10683,N_10391,N_10345);
nand U10684 (N_10684,N_10439,N_10316);
and U10685 (N_10685,N_10256,N_10422);
nand U10686 (N_10686,N_10269,N_10310);
xor U10687 (N_10687,N_10339,N_10394);
and U10688 (N_10688,N_10348,N_10472);
nor U10689 (N_10689,N_10302,N_10425);
nand U10690 (N_10690,N_10395,N_10361);
or U10691 (N_10691,N_10316,N_10284);
and U10692 (N_10692,N_10288,N_10400);
nor U10693 (N_10693,N_10262,N_10498);
xor U10694 (N_10694,N_10351,N_10462);
and U10695 (N_10695,N_10256,N_10376);
nor U10696 (N_10696,N_10378,N_10315);
nor U10697 (N_10697,N_10299,N_10444);
or U10698 (N_10698,N_10377,N_10291);
and U10699 (N_10699,N_10397,N_10414);
xor U10700 (N_10700,N_10412,N_10294);
xor U10701 (N_10701,N_10459,N_10386);
and U10702 (N_10702,N_10431,N_10450);
nand U10703 (N_10703,N_10281,N_10370);
or U10704 (N_10704,N_10394,N_10312);
and U10705 (N_10705,N_10265,N_10308);
nand U10706 (N_10706,N_10351,N_10493);
nand U10707 (N_10707,N_10398,N_10493);
xnor U10708 (N_10708,N_10270,N_10485);
or U10709 (N_10709,N_10299,N_10373);
or U10710 (N_10710,N_10305,N_10359);
nor U10711 (N_10711,N_10311,N_10407);
nor U10712 (N_10712,N_10269,N_10343);
nand U10713 (N_10713,N_10415,N_10435);
xnor U10714 (N_10714,N_10426,N_10303);
nand U10715 (N_10715,N_10353,N_10450);
or U10716 (N_10716,N_10312,N_10418);
or U10717 (N_10717,N_10438,N_10301);
xnor U10718 (N_10718,N_10275,N_10423);
or U10719 (N_10719,N_10433,N_10304);
or U10720 (N_10720,N_10498,N_10308);
and U10721 (N_10721,N_10345,N_10339);
xnor U10722 (N_10722,N_10340,N_10349);
nand U10723 (N_10723,N_10459,N_10454);
or U10724 (N_10724,N_10263,N_10489);
nor U10725 (N_10725,N_10428,N_10483);
nor U10726 (N_10726,N_10474,N_10252);
nor U10727 (N_10727,N_10379,N_10368);
or U10728 (N_10728,N_10443,N_10357);
nand U10729 (N_10729,N_10252,N_10293);
nor U10730 (N_10730,N_10296,N_10460);
or U10731 (N_10731,N_10354,N_10292);
or U10732 (N_10732,N_10301,N_10480);
and U10733 (N_10733,N_10457,N_10252);
and U10734 (N_10734,N_10363,N_10410);
nor U10735 (N_10735,N_10469,N_10489);
nand U10736 (N_10736,N_10400,N_10252);
nor U10737 (N_10737,N_10330,N_10291);
nand U10738 (N_10738,N_10383,N_10299);
xnor U10739 (N_10739,N_10367,N_10488);
nor U10740 (N_10740,N_10257,N_10499);
and U10741 (N_10741,N_10457,N_10381);
nor U10742 (N_10742,N_10329,N_10335);
or U10743 (N_10743,N_10429,N_10408);
or U10744 (N_10744,N_10280,N_10477);
nand U10745 (N_10745,N_10482,N_10447);
or U10746 (N_10746,N_10274,N_10388);
and U10747 (N_10747,N_10440,N_10490);
xnor U10748 (N_10748,N_10370,N_10426);
or U10749 (N_10749,N_10351,N_10429);
and U10750 (N_10750,N_10520,N_10740);
or U10751 (N_10751,N_10694,N_10624);
nand U10752 (N_10752,N_10524,N_10707);
xnor U10753 (N_10753,N_10655,N_10528);
xor U10754 (N_10754,N_10680,N_10716);
and U10755 (N_10755,N_10526,N_10614);
nand U10756 (N_10756,N_10661,N_10568);
and U10757 (N_10757,N_10611,N_10737);
nor U10758 (N_10758,N_10579,N_10552);
xnor U10759 (N_10759,N_10563,N_10710);
or U10760 (N_10760,N_10717,N_10708);
or U10761 (N_10761,N_10660,N_10733);
xor U10762 (N_10762,N_10695,N_10630);
xor U10763 (N_10763,N_10683,N_10651);
nor U10764 (N_10764,N_10731,N_10502);
and U10765 (N_10765,N_10510,N_10506);
nand U10766 (N_10766,N_10743,N_10561);
or U10767 (N_10767,N_10514,N_10523);
nor U10768 (N_10768,N_10719,N_10530);
nor U10769 (N_10769,N_10650,N_10726);
xor U10770 (N_10770,N_10503,N_10622);
nand U10771 (N_10771,N_10612,N_10557);
nor U10772 (N_10772,N_10629,N_10747);
nand U10773 (N_10773,N_10544,N_10541);
or U10774 (N_10774,N_10543,N_10516);
and U10775 (N_10775,N_10635,N_10511);
and U10776 (N_10776,N_10537,N_10572);
nor U10777 (N_10777,N_10625,N_10539);
xor U10778 (N_10778,N_10678,N_10674);
or U10779 (N_10779,N_10592,N_10636);
xor U10780 (N_10780,N_10648,N_10598);
and U10781 (N_10781,N_10555,N_10679);
nor U10782 (N_10782,N_10685,N_10748);
and U10783 (N_10783,N_10613,N_10741);
xor U10784 (N_10784,N_10595,N_10704);
and U10785 (N_10785,N_10601,N_10712);
or U10786 (N_10786,N_10631,N_10736);
and U10787 (N_10787,N_10522,N_10730);
nand U10788 (N_10788,N_10647,N_10692);
xor U10789 (N_10789,N_10597,N_10633);
nand U10790 (N_10790,N_10681,N_10585);
and U10791 (N_10791,N_10735,N_10628);
xnor U10792 (N_10792,N_10582,N_10697);
nand U10793 (N_10793,N_10723,N_10593);
and U10794 (N_10794,N_10594,N_10641);
nor U10795 (N_10795,N_10643,N_10721);
xor U10796 (N_10796,N_10682,N_10724);
nor U10797 (N_10797,N_10659,N_10556);
and U10798 (N_10798,N_10727,N_10702);
nor U10799 (N_10799,N_10604,N_10550);
and U10800 (N_10800,N_10696,N_10646);
xnor U10801 (N_10801,N_10621,N_10618);
nor U10802 (N_10802,N_10616,N_10548);
nor U10803 (N_10803,N_10599,N_10684);
nand U10804 (N_10804,N_10742,N_10638);
or U10805 (N_10805,N_10690,N_10688);
or U10806 (N_10806,N_10518,N_10645);
xnor U10807 (N_10807,N_10590,N_10700);
xnor U10808 (N_10808,N_10619,N_10567);
nor U10809 (N_10809,N_10517,N_10734);
nand U10810 (N_10810,N_10637,N_10553);
xor U10811 (N_10811,N_10578,N_10686);
xnor U10812 (N_10812,N_10536,N_10535);
and U10813 (N_10813,N_10709,N_10657);
and U10814 (N_10814,N_10559,N_10698);
xor U10815 (N_10815,N_10505,N_10722);
xnor U10816 (N_10816,N_10632,N_10658);
nand U10817 (N_10817,N_10689,N_10519);
or U10818 (N_10818,N_10521,N_10603);
nor U10819 (N_10819,N_10589,N_10554);
xor U10820 (N_10820,N_10720,N_10665);
and U10821 (N_10821,N_10738,N_10558);
nand U10822 (N_10822,N_10501,N_10718);
or U10823 (N_10823,N_10666,N_10623);
or U10824 (N_10824,N_10706,N_10607);
xor U10825 (N_10825,N_10513,N_10639);
and U10826 (N_10826,N_10673,N_10570);
nor U10827 (N_10827,N_10566,N_10652);
nand U10828 (N_10828,N_10617,N_10500);
xor U10829 (N_10829,N_10671,N_10642);
or U10830 (N_10830,N_10507,N_10549);
nor U10831 (N_10831,N_10703,N_10732);
nand U10832 (N_10832,N_10531,N_10654);
xnor U10833 (N_10833,N_10699,N_10746);
xor U10834 (N_10834,N_10596,N_10605);
nand U10835 (N_10835,N_10653,N_10586);
nor U10836 (N_10836,N_10615,N_10569);
nor U10837 (N_10837,N_10608,N_10609);
or U10838 (N_10838,N_10532,N_10551);
and U10839 (N_10839,N_10739,N_10508);
and U10840 (N_10840,N_10668,N_10580);
and U10841 (N_10841,N_10527,N_10729);
or U10842 (N_10842,N_10687,N_10573);
nand U10843 (N_10843,N_10542,N_10562);
or U10844 (N_10844,N_10564,N_10565);
and U10845 (N_10845,N_10525,N_10588);
and U10846 (N_10846,N_10644,N_10606);
and U10847 (N_10847,N_10538,N_10509);
or U10848 (N_10848,N_10675,N_10693);
and U10849 (N_10849,N_10571,N_10534);
and U10850 (N_10850,N_10705,N_10728);
and U10851 (N_10851,N_10670,N_10667);
xnor U10852 (N_10852,N_10512,N_10676);
nor U10853 (N_10853,N_10749,N_10574);
xor U10854 (N_10854,N_10610,N_10591);
and U10855 (N_10855,N_10662,N_10745);
nand U10856 (N_10856,N_10634,N_10713);
nand U10857 (N_10857,N_10672,N_10533);
xnor U10858 (N_10858,N_10529,N_10649);
and U10859 (N_10859,N_10560,N_10701);
and U10860 (N_10860,N_10584,N_10602);
nand U10861 (N_10861,N_10600,N_10620);
and U10862 (N_10862,N_10515,N_10626);
or U10863 (N_10863,N_10546,N_10587);
nor U10864 (N_10864,N_10627,N_10504);
and U10865 (N_10865,N_10744,N_10669);
and U10866 (N_10866,N_10715,N_10677);
xnor U10867 (N_10867,N_10583,N_10575);
and U10868 (N_10868,N_10725,N_10711);
nand U10869 (N_10869,N_10545,N_10581);
or U10870 (N_10870,N_10691,N_10547);
and U10871 (N_10871,N_10540,N_10577);
or U10872 (N_10872,N_10656,N_10640);
nand U10873 (N_10873,N_10576,N_10663);
or U10874 (N_10874,N_10664,N_10714);
or U10875 (N_10875,N_10531,N_10541);
or U10876 (N_10876,N_10657,N_10603);
nand U10877 (N_10877,N_10519,N_10627);
nand U10878 (N_10878,N_10551,N_10627);
and U10879 (N_10879,N_10598,N_10571);
nor U10880 (N_10880,N_10515,N_10595);
xor U10881 (N_10881,N_10564,N_10529);
and U10882 (N_10882,N_10542,N_10531);
and U10883 (N_10883,N_10664,N_10512);
xor U10884 (N_10884,N_10578,N_10747);
nor U10885 (N_10885,N_10690,N_10563);
nand U10886 (N_10886,N_10626,N_10611);
nand U10887 (N_10887,N_10593,N_10625);
nor U10888 (N_10888,N_10586,N_10665);
or U10889 (N_10889,N_10622,N_10612);
xor U10890 (N_10890,N_10615,N_10598);
or U10891 (N_10891,N_10612,N_10593);
nor U10892 (N_10892,N_10515,N_10638);
xor U10893 (N_10893,N_10729,N_10569);
or U10894 (N_10894,N_10503,N_10689);
xor U10895 (N_10895,N_10730,N_10617);
xor U10896 (N_10896,N_10516,N_10528);
nor U10897 (N_10897,N_10665,N_10694);
xor U10898 (N_10898,N_10596,N_10675);
nand U10899 (N_10899,N_10595,N_10565);
xnor U10900 (N_10900,N_10717,N_10526);
or U10901 (N_10901,N_10712,N_10637);
or U10902 (N_10902,N_10513,N_10665);
xor U10903 (N_10903,N_10570,N_10525);
nor U10904 (N_10904,N_10584,N_10585);
and U10905 (N_10905,N_10617,N_10534);
or U10906 (N_10906,N_10625,N_10740);
nand U10907 (N_10907,N_10605,N_10575);
xnor U10908 (N_10908,N_10741,N_10692);
or U10909 (N_10909,N_10586,N_10559);
nand U10910 (N_10910,N_10667,N_10629);
nand U10911 (N_10911,N_10593,N_10547);
nand U10912 (N_10912,N_10603,N_10676);
nand U10913 (N_10913,N_10642,N_10550);
or U10914 (N_10914,N_10693,N_10570);
xnor U10915 (N_10915,N_10651,N_10521);
nor U10916 (N_10916,N_10715,N_10739);
nand U10917 (N_10917,N_10675,N_10647);
nand U10918 (N_10918,N_10633,N_10506);
nand U10919 (N_10919,N_10524,N_10737);
nor U10920 (N_10920,N_10641,N_10667);
xnor U10921 (N_10921,N_10747,N_10726);
nand U10922 (N_10922,N_10642,N_10708);
xnor U10923 (N_10923,N_10536,N_10531);
nand U10924 (N_10924,N_10716,N_10500);
and U10925 (N_10925,N_10504,N_10636);
nor U10926 (N_10926,N_10599,N_10593);
or U10927 (N_10927,N_10514,N_10683);
or U10928 (N_10928,N_10691,N_10717);
nand U10929 (N_10929,N_10536,N_10538);
and U10930 (N_10930,N_10712,N_10642);
or U10931 (N_10931,N_10574,N_10721);
or U10932 (N_10932,N_10702,N_10726);
nand U10933 (N_10933,N_10538,N_10504);
nor U10934 (N_10934,N_10703,N_10549);
xor U10935 (N_10935,N_10699,N_10518);
nand U10936 (N_10936,N_10678,N_10664);
nand U10937 (N_10937,N_10674,N_10569);
nand U10938 (N_10938,N_10741,N_10556);
xor U10939 (N_10939,N_10646,N_10707);
and U10940 (N_10940,N_10601,N_10568);
xnor U10941 (N_10941,N_10566,N_10605);
xnor U10942 (N_10942,N_10673,N_10705);
and U10943 (N_10943,N_10720,N_10712);
nor U10944 (N_10944,N_10748,N_10744);
nor U10945 (N_10945,N_10532,N_10545);
nand U10946 (N_10946,N_10673,N_10541);
and U10947 (N_10947,N_10642,N_10503);
xor U10948 (N_10948,N_10688,N_10657);
nor U10949 (N_10949,N_10539,N_10657);
xnor U10950 (N_10950,N_10613,N_10683);
nand U10951 (N_10951,N_10723,N_10686);
nor U10952 (N_10952,N_10599,N_10627);
xnor U10953 (N_10953,N_10746,N_10721);
nor U10954 (N_10954,N_10516,N_10557);
xor U10955 (N_10955,N_10695,N_10613);
nor U10956 (N_10956,N_10707,N_10553);
xnor U10957 (N_10957,N_10696,N_10714);
xnor U10958 (N_10958,N_10716,N_10732);
xor U10959 (N_10959,N_10713,N_10512);
nand U10960 (N_10960,N_10710,N_10628);
and U10961 (N_10961,N_10517,N_10609);
or U10962 (N_10962,N_10653,N_10623);
nor U10963 (N_10963,N_10619,N_10535);
and U10964 (N_10964,N_10565,N_10502);
nor U10965 (N_10965,N_10661,N_10588);
nand U10966 (N_10966,N_10685,N_10609);
nand U10967 (N_10967,N_10726,N_10562);
and U10968 (N_10968,N_10577,N_10680);
nand U10969 (N_10969,N_10679,N_10591);
xnor U10970 (N_10970,N_10682,N_10669);
xor U10971 (N_10971,N_10630,N_10742);
xnor U10972 (N_10972,N_10581,N_10625);
or U10973 (N_10973,N_10640,N_10542);
and U10974 (N_10974,N_10527,N_10568);
nor U10975 (N_10975,N_10727,N_10708);
or U10976 (N_10976,N_10646,N_10596);
nor U10977 (N_10977,N_10654,N_10676);
or U10978 (N_10978,N_10619,N_10546);
xnor U10979 (N_10979,N_10644,N_10593);
and U10980 (N_10980,N_10572,N_10640);
and U10981 (N_10981,N_10673,N_10664);
xor U10982 (N_10982,N_10529,N_10584);
nand U10983 (N_10983,N_10708,N_10605);
nand U10984 (N_10984,N_10539,N_10563);
and U10985 (N_10985,N_10694,N_10560);
nor U10986 (N_10986,N_10719,N_10727);
or U10987 (N_10987,N_10734,N_10696);
or U10988 (N_10988,N_10540,N_10738);
and U10989 (N_10989,N_10690,N_10582);
xnor U10990 (N_10990,N_10507,N_10503);
nor U10991 (N_10991,N_10567,N_10741);
and U10992 (N_10992,N_10578,N_10617);
and U10993 (N_10993,N_10538,N_10527);
or U10994 (N_10994,N_10733,N_10551);
nor U10995 (N_10995,N_10530,N_10624);
or U10996 (N_10996,N_10574,N_10511);
xor U10997 (N_10997,N_10521,N_10711);
xor U10998 (N_10998,N_10624,N_10742);
and U10999 (N_10999,N_10579,N_10728);
nand U11000 (N_11000,N_10784,N_10963);
nand U11001 (N_11001,N_10959,N_10929);
xor U11002 (N_11002,N_10758,N_10868);
xnor U11003 (N_11003,N_10806,N_10791);
nor U11004 (N_11004,N_10986,N_10948);
nor U11005 (N_11005,N_10964,N_10955);
nor U11006 (N_11006,N_10821,N_10858);
or U11007 (N_11007,N_10870,N_10914);
nor U11008 (N_11008,N_10942,N_10980);
or U11009 (N_11009,N_10864,N_10916);
xor U11010 (N_11010,N_10968,N_10876);
nor U11011 (N_11011,N_10899,N_10969);
xnor U11012 (N_11012,N_10975,N_10895);
and U11013 (N_11013,N_10953,N_10800);
and U11014 (N_11014,N_10880,N_10844);
and U11015 (N_11015,N_10897,N_10911);
nand U11016 (N_11016,N_10863,N_10952);
nand U11017 (N_11017,N_10935,N_10773);
or U11018 (N_11018,N_10967,N_10869);
nor U11019 (N_11019,N_10789,N_10988);
xnor U11020 (N_11020,N_10941,N_10946);
xor U11021 (N_11021,N_10756,N_10814);
and U11022 (N_11022,N_10878,N_10875);
or U11023 (N_11023,N_10796,N_10910);
nand U11024 (N_11024,N_10932,N_10904);
and U11025 (N_11025,N_10859,N_10985);
and U11026 (N_11026,N_10830,N_10798);
xnor U11027 (N_11027,N_10768,N_10882);
nand U11028 (N_11028,N_10804,N_10797);
xnor U11029 (N_11029,N_10930,N_10908);
or U11030 (N_11030,N_10794,N_10823);
or U11031 (N_11031,N_10865,N_10767);
nor U11032 (N_11032,N_10822,N_10936);
xnor U11033 (N_11033,N_10818,N_10927);
and U11034 (N_11034,N_10838,N_10802);
and U11035 (N_11035,N_10901,N_10807);
nor U11036 (N_11036,N_10944,N_10873);
nor U11037 (N_11037,N_10752,N_10771);
xor U11038 (N_11038,N_10765,N_10801);
nor U11039 (N_11039,N_10779,N_10851);
nor U11040 (N_11040,N_10984,N_10759);
and U11041 (N_11041,N_10907,N_10898);
and U11042 (N_11042,N_10762,N_10855);
xor U11043 (N_11043,N_10778,N_10799);
and U11044 (N_11044,N_10939,N_10937);
and U11045 (N_11045,N_10862,N_10894);
nand U11046 (N_11046,N_10788,N_10774);
nand U11047 (N_11047,N_10833,N_10871);
nand U11048 (N_11048,N_10813,N_10976);
nor U11049 (N_11049,N_10999,N_10850);
xnor U11050 (N_11050,N_10861,N_10888);
and U11051 (N_11051,N_10820,N_10884);
and U11052 (N_11052,N_10761,N_10921);
or U11053 (N_11053,N_10962,N_10912);
or U11054 (N_11054,N_10934,N_10816);
xor U11055 (N_11055,N_10812,N_10866);
nor U11056 (N_11056,N_10931,N_10811);
nand U11057 (N_11057,N_10991,N_10775);
xnor U11058 (N_11058,N_10994,N_10996);
and U11059 (N_11059,N_10849,N_10772);
and U11060 (N_11060,N_10841,N_10848);
and U11061 (N_11061,N_10776,N_10909);
nand U11062 (N_11062,N_10970,N_10764);
or U11063 (N_11063,N_10961,N_10890);
xor U11064 (N_11064,N_10893,N_10956);
and U11065 (N_11065,N_10872,N_10896);
nand U11066 (N_11066,N_10874,N_10808);
xnor U11067 (N_11067,N_10965,N_10781);
or U11068 (N_11068,N_10995,N_10840);
and U11069 (N_11069,N_10795,N_10977);
nand U11070 (N_11070,N_10786,N_10825);
xnor U11071 (N_11071,N_10792,N_10993);
xnor U11072 (N_11072,N_10782,N_10867);
or U11073 (N_11073,N_10928,N_10925);
nand U11074 (N_11074,N_10889,N_10815);
and U11075 (N_11075,N_10966,N_10973);
nor U11076 (N_11076,N_10983,N_10857);
and U11077 (N_11077,N_10949,N_10951);
nor U11078 (N_11078,N_10892,N_10785);
nor U11079 (N_11079,N_10954,N_10923);
and U11080 (N_11080,N_10913,N_10978);
nand U11081 (N_11081,N_10979,N_10924);
nand U11082 (N_11082,N_10829,N_10905);
nor U11083 (N_11083,N_10918,N_10831);
nor U11084 (N_11084,N_10860,N_10835);
or U11085 (N_11085,N_10981,N_10922);
nand U11086 (N_11086,N_10834,N_10920);
and U11087 (N_11087,N_10883,N_10847);
nand U11088 (N_11088,N_10902,N_10832);
xor U11089 (N_11089,N_10777,N_10943);
and U11090 (N_11090,N_10803,N_10886);
nor U11091 (N_11091,N_10839,N_10900);
nand U11092 (N_11092,N_10760,N_10992);
nand U11093 (N_11093,N_10787,N_10828);
nor U11094 (N_11094,N_10987,N_10809);
and U11095 (N_11095,N_10766,N_10906);
nor U11096 (N_11096,N_10877,N_10837);
nor U11097 (N_11097,N_10885,N_10971);
and U11098 (N_11098,N_10853,N_10826);
nand U11099 (N_11099,N_10770,N_10945);
xor U11100 (N_11100,N_10933,N_10843);
or U11101 (N_11101,N_10887,N_10754);
or U11102 (N_11102,N_10856,N_10917);
xor U11103 (N_11103,N_10810,N_10836);
xnor U11104 (N_11104,N_10972,N_10974);
nand U11105 (N_11105,N_10819,N_10926);
or U11106 (N_11106,N_10769,N_10919);
nand U11107 (N_11107,N_10750,N_10757);
xor U11108 (N_11108,N_10982,N_10881);
xnor U11109 (N_11109,N_10783,N_10824);
nand U11110 (N_11110,N_10938,N_10846);
nor U11111 (N_11111,N_10958,N_10805);
xor U11112 (N_11112,N_10879,N_10960);
xnor U11113 (N_11113,N_10827,N_10950);
nand U11114 (N_11114,N_10854,N_10842);
xor U11115 (N_11115,N_10780,N_10790);
or U11116 (N_11116,N_10989,N_10845);
or U11117 (N_11117,N_10940,N_10990);
nor U11118 (N_11118,N_10891,N_10817);
nand U11119 (N_11119,N_10763,N_10793);
or U11120 (N_11120,N_10998,N_10957);
and U11121 (N_11121,N_10903,N_10751);
and U11122 (N_11122,N_10753,N_10852);
nand U11123 (N_11123,N_10755,N_10997);
or U11124 (N_11124,N_10947,N_10915);
and U11125 (N_11125,N_10936,N_10816);
nand U11126 (N_11126,N_10877,N_10854);
xnor U11127 (N_11127,N_10925,N_10890);
nand U11128 (N_11128,N_10937,N_10995);
nand U11129 (N_11129,N_10895,N_10989);
nand U11130 (N_11130,N_10956,N_10759);
nand U11131 (N_11131,N_10849,N_10933);
nand U11132 (N_11132,N_10991,N_10874);
nand U11133 (N_11133,N_10811,N_10754);
xor U11134 (N_11134,N_10989,N_10953);
or U11135 (N_11135,N_10779,N_10775);
nand U11136 (N_11136,N_10879,N_10968);
nand U11137 (N_11137,N_10907,N_10877);
xnor U11138 (N_11138,N_10992,N_10856);
and U11139 (N_11139,N_10861,N_10968);
or U11140 (N_11140,N_10798,N_10755);
xor U11141 (N_11141,N_10832,N_10796);
nand U11142 (N_11142,N_10937,N_10836);
nand U11143 (N_11143,N_10989,N_10784);
xor U11144 (N_11144,N_10910,N_10751);
nand U11145 (N_11145,N_10965,N_10923);
nor U11146 (N_11146,N_10909,N_10862);
and U11147 (N_11147,N_10895,N_10875);
xor U11148 (N_11148,N_10766,N_10803);
or U11149 (N_11149,N_10846,N_10958);
and U11150 (N_11150,N_10856,N_10807);
nand U11151 (N_11151,N_10926,N_10980);
nor U11152 (N_11152,N_10890,N_10980);
nand U11153 (N_11153,N_10970,N_10990);
or U11154 (N_11154,N_10843,N_10937);
xor U11155 (N_11155,N_10858,N_10755);
and U11156 (N_11156,N_10887,N_10991);
nor U11157 (N_11157,N_10968,N_10858);
and U11158 (N_11158,N_10981,N_10923);
or U11159 (N_11159,N_10933,N_10970);
and U11160 (N_11160,N_10807,N_10934);
nor U11161 (N_11161,N_10824,N_10993);
xnor U11162 (N_11162,N_10886,N_10974);
nor U11163 (N_11163,N_10803,N_10869);
xor U11164 (N_11164,N_10966,N_10810);
or U11165 (N_11165,N_10942,N_10848);
nor U11166 (N_11166,N_10974,N_10828);
and U11167 (N_11167,N_10825,N_10788);
nand U11168 (N_11168,N_10835,N_10873);
xor U11169 (N_11169,N_10995,N_10956);
or U11170 (N_11170,N_10939,N_10751);
nand U11171 (N_11171,N_10998,N_10790);
nand U11172 (N_11172,N_10977,N_10967);
nor U11173 (N_11173,N_10952,N_10872);
nand U11174 (N_11174,N_10980,N_10832);
and U11175 (N_11175,N_10989,N_10930);
nor U11176 (N_11176,N_10811,N_10962);
nand U11177 (N_11177,N_10932,N_10868);
and U11178 (N_11178,N_10939,N_10759);
or U11179 (N_11179,N_10986,N_10958);
and U11180 (N_11180,N_10887,N_10968);
and U11181 (N_11181,N_10909,N_10895);
nand U11182 (N_11182,N_10960,N_10868);
nand U11183 (N_11183,N_10968,N_10755);
nor U11184 (N_11184,N_10882,N_10857);
and U11185 (N_11185,N_10794,N_10948);
xor U11186 (N_11186,N_10993,N_10851);
or U11187 (N_11187,N_10916,N_10800);
or U11188 (N_11188,N_10815,N_10901);
and U11189 (N_11189,N_10891,N_10951);
or U11190 (N_11190,N_10952,N_10849);
or U11191 (N_11191,N_10799,N_10817);
nand U11192 (N_11192,N_10862,N_10979);
nor U11193 (N_11193,N_10980,N_10872);
and U11194 (N_11194,N_10990,N_10890);
nand U11195 (N_11195,N_10800,N_10889);
xor U11196 (N_11196,N_10971,N_10770);
or U11197 (N_11197,N_10922,N_10802);
and U11198 (N_11198,N_10786,N_10919);
and U11199 (N_11199,N_10923,N_10840);
and U11200 (N_11200,N_10787,N_10814);
or U11201 (N_11201,N_10992,N_10776);
nand U11202 (N_11202,N_10852,N_10772);
nor U11203 (N_11203,N_10879,N_10832);
nor U11204 (N_11204,N_10966,N_10867);
nand U11205 (N_11205,N_10803,N_10980);
or U11206 (N_11206,N_10884,N_10910);
xor U11207 (N_11207,N_10789,N_10786);
or U11208 (N_11208,N_10937,N_10954);
nor U11209 (N_11209,N_10943,N_10958);
nand U11210 (N_11210,N_10839,N_10792);
nand U11211 (N_11211,N_10753,N_10964);
nand U11212 (N_11212,N_10887,N_10766);
xor U11213 (N_11213,N_10841,N_10786);
or U11214 (N_11214,N_10918,N_10974);
nand U11215 (N_11215,N_10830,N_10813);
nand U11216 (N_11216,N_10844,N_10811);
nand U11217 (N_11217,N_10750,N_10852);
nand U11218 (N_11218,N_10925,N_10895);
xor U11219 (N_11219,N_10948,N_10884);
nor U11220 (N_11220,N_10981,N_10869);
nand U11221 (N_11221,N_10763,N_10970);
or U11222 (N_11222,N_10977,N_10861);
nand U11223 (N_11223,N_10948,N_10957);
nand U11224 (N_11224,N_10976,N_10908);
nor U11225 (N_11225,N_10907,N_10841);
nor U11226 (N_11226,N_10996,N_10897);
nor U11227 (N_11227,N_10792,N_10936);
xor U11228 (N_11228,N_10800,N_10942);
nor U11229 (N_11229,N_10786,N_10899);
or U11230 (N_11230,N_10958,N_10984);
xor U11231 (N_11231,N_10877,N_10957);
nand U11232 (N_11232,N_10813,N_10836);
and U11233 (N_11233,N_10866,N_10827);
and U11234 (N_11234,N_10928,N_10951);
and U11235 (N_11235,N_10819,N_10938);
nand U11236 (N_11236,N_10840,N_10788);
nor U11237 (N_11237,N_10965,N_10907);
nand U11238 (N_11238,N_10928,N_10849);
nor U11239 (N_11239,N_10820,N_10813);
xor U11240 (N_11240,N_10794,N_10937);
and U11241 (N_11241,N_10932,N_10801);
and U11242 (N_11242,N_10834,N_10916);
or U11243 (N_11243,N_10955,N_10786);
or U11244 (N_11244,N_10794,N_10936);
or U11245 (N_11245,N_10913,N_10875);
nor U11246 (N_11246,N_10917,N_10835);
nand U11247 (N_11247,N_10846,N_10753);
nor U11248 (N_11248,N_10914,N_10937);
xor U11249 (N_11249,N_10940,N_10936);
nor U11250 (N_11250,N_11041,N_11138);
xor U11251 (N_11251,N_11120,N_11222);
nand U11252 (N_11252,N_11227,N_11155);
nor U11253 (N_11253,N_11075,N_11144);
nand U11254 (N_11254,N_11081,N_11195);
or U11255 (N_11255,N_11171,N_11172);
nand U11256 (N_11256,N_11135,N_11108);
nand U11257 (N_11257,N_11057,N_11249);
xor U11258 (N_11258,N_11140,N_11116);
nor U11259 (N_11259,N_11213,N_11058);
xor U11260 (N_11260,N_11221,N_11111);
and U11261 (N_11261,N_11173,N_11022);
or U11262 (N_11262,N_11244,N_11190);
or U11263 (N_11263,N_11113,N_11093);
or U11264 (N_11264,N_11228,N_11127);
nor U11265 (N_11265,N_11198,N_11086);
or U11266 (N_11266,N_11042,N_11072);
xor U11267 (N_11267,N_11009,N_11176);
xnor U11268 (N_11268,N_11174,N_11117);
nor U11269 (N_11269,N_11211,N_11010);
nor U11270 (N_11270,N_11078,N_11157);
nand U11271 (N_11271,N_11018,N_11153);
nor U11272 (N_11272,N_11148,N_11114);
nand U11273 (N_11273,N_11030,N_11133);
nand U11274 (N_11274,N_11092,N_11008);
and U11275 (N_11275,N_11131,N_11082);
and U11276 (N_11276,N_11197,N_11205);
xnor U11277 (N_11277,N_11019,N_11181);
or U11278 (N_11278,N_11007,N_11214);
nor U11279 (N_11279,N_11103,N_11161);
or U11280 (N_11280,N_11217,N_11015);
or U11281 (N_11281,N_11162,N_11179);
and U11282 (N_11282,N_11106,N_11166);
nor U11283 (N_11283,N_11132,N_11164);
or U11284 (N_11284,N_11090,N_11187);
or U11285 (N_11285,N_11071,N_11234);
nand U11286 (N_11286,N_11165,N_11121);
nor U11287 (N_11287,N_11033,N_11077);
xnor U11288 (N_11288,N_11073,N_11087);
or U11289 (N_11289,N_11137,N_11115);
or U11290 (N_11290,N_11185,N_11056);
nor U11291 (N_11291,N_11067,N_11031);
and U11292 (N_11292,N_11223,N_11066);
xnor U11293 (N_11293,N_11200,N_11230);
xor U11294 (N_11294,N_11012,N_11158);
nand U11295 (N_11295,N_11156,N_11054);
or U11296 (N_11296,N_11143,N_11177);
or U11297 (N_11297,N_11063,N_11020);
xnor U11298 (N_11298,N_11122,N_11237);
and U11299 (N_11299,N_11003,N_11220);
nand U11300 (N_11300,N_11112,N_11246);
xor U11301 (N_11301,N_11076,N_11101);
nand U11302 (N_11302,N_11088,N_11040);
and U11303 (N_11303,N_11189,N_11100);
xor U11304 (N_11304,N_11248,N_11027);
and U11305 (N_11305,N_11050,N_11049);
xnor U11306 (N_11306,N_11184,N_11046);
or U11307 (N_11307,N_11139,N_11145);
nand U11308 (N_11308,N_11229,N_11091);
nor U11309 (N_11309,N_11017,N_11005);
or U11310 (N_11310,N_11104,N_11002);
nor U11311 (N_11311,N_11098,N_11242);
nand U11312 (N_11312,N_11136,N_11001);
nor U11313 (N_11313,N_11247,N_11240);
nand U11314 (N_11314,N_11194,N_11011);
nor U11315 (N_11315,N_11102,N_11210);
nand U11316 (N_11316,N_11159,N_11235);
xnor U11317 (N_11317,N_11188,N_11224);
nand U11318 (N_11318,N_11149,N_11037);
nand U11319 (N_11319,N_11062,N_11048);
xnor U11320 (N_11320,N_11036,N_11209);
nand U11321 (N_11321,N_11192,N_11207);
and U11322 (N_11322,N_11055,N_11029);
or U11323 (N_11323,N_11238,N_11163);
and U11324 (N_11324,N_11044,N_11226);
or U11325 (N_11325,N_11241,N_11169);
xnor U11326 (N_11326,N_11193,N_11096);
or U11327 (N_11327,N_11013,N_11070);
and U11328 (N_11328,N_11119,N_11107);
nand U11329 (N_11329,N_11069,N_11160);
nor U11330 (N_11330,N_11225,N_11128);
nor U11331 (N_11331,N_11097,N_11061);
nor U11332 (N_11332,N_11168,N_11196);
nand U11333 (N_11333,N_11038,N_11124);
or U11334 (N_11334,N_11231,N_11126);
nand U11335 (N_11335,N_11035,N_11216);
or U11336 (N_11336,N_11167,N_11178);
nand U11337 (N_11337,N_11130,N_11129);
nor U11338 (N_11338,N_11052,N_11023);
nor U11339 (N_11339,N_11191,N_11045);
and U11340 (N_11340,N_11233,N_11186);
nand U11341 (N_11341,N_11059,N_11006);
xnor U11342 (N_11342,N_11134,N_11079);
nor U11343 (N_11343,N_11021,N_11146);
xnor U11344 (N_11344,N_11043,N_11094);
nor U11345 (N_11345,N_11147,N_11109);
nand U11346 (N_11346,N_11074,N_11034);
nor U11347 (N_11347,N_11219,N_11016);
xor U11348 (N_11348,N_11239,N_11204);
nand U11349 (N_11349,N_11060,N_11110);
nor U11350 (N_11350,N_11141,N_11175);
xnor U11351 (N_11351,N_11080,N_11218);
or U11352 (N_11352,N_11202,N_11084);
or U11353 (N_11353,N_11182,N_11039);
nand U11354 (N_11354,N_11064,N_11051);
and U11355 (N_11355,N_11065,N_11206);
or U11356 (N_11356,N_11026,N_11024);
nand U11357 (N_11357,N_11245,N_11099);
nor U11358 (N_11358,N_11232,N_11243);
or U11359 (N_11359,N_11025,N_11170);
and U11360 (N_11360,N_11047,N_11151);
and U11361 (N_11361,N_11199,N_11203);
xor U11362 (N_11362,N_11004,N_11142);
nand U11363 (N_11363,N_11095,N_11236);
and U11364 (N_11364,N_11180,N_11083);
xor U11365 (N_11365,N_11068,N_11000);
or U11366 (N_11366,N_11123,N_11125);
nor U11367 (N_11367,N_11085,N_11201);
nor U11368 (N_11368,N_11089,N_11212);
xor U11369 (N_11369,N_11150,N_11152);
or U11370 (N_11370,N_11053,N_11215);
and U11371 (N_11371,N_11183,N_11028);
or U11372 (N_11372,N_11118,N_11208);
nor U11373 (N_11373,N_11154,N_11032);
nor U11374 (N_11374,N_11014,N_11105);
nand U11375 (N_11375,N_11182,N_11242);
or U11376 (N_11376,N_11074,N_11168);
nand U11377 (N_11377,N_11147,N_11077);
nor U11378 (N_11378,N_11135,N_11087);
and U11379 (N_11379,N_11139,N_11163);
or U11380 (N_11380,N_11069,N_11232);
and U11381 (N_11381,N_11040,N_11089);
xor U11382 (N_11382,N_11245,N_11108);
and U11383 (N_11383,N_11054,N_11212);
or U11384 (N_11384,N_11055,N_11022);
xor U11385 (N_11385,N_11028,N_11074);
nand U11386 (N_11386,N_11074,N_11199);
and U11387 (N_11387,N_11110,N_11102);
nor U11388 (N_11388,N_11097,N_11159);
nor U11389 (N_11389,N_11242,N_11165);
nand U11390 (N_11390,N_11013,N_11050);
nand U11391 (N_11391,N_11102,N_11030);
nand U11392 (N_11392,N_11128,N_11144);
xnor U11393 (N_11393,N_11175,N_11103);
nand U11394 (N_11394,N_11203,N_11084);
and U11395 (N_11395,N_11246,N_11115);
and U11396 (N_11396,N_11218,N_11224);
nor U11397 (N_11397,N_11190,N_11083);
xnor U11398 (N_11398,N_11214,N_11203);
or U11399 (N_11399,N_11030,N_11013);
and U11400 (N_11400,N_11019,N_11060);
and U11401 (N_11401,N_11109,N_11209);
xnor U11402 (N_11402,N_11077,N_11080);
xnor U11403 (N_11403,N_11174,N_11043);
nand U11404 (N_11404,N_11112,N_11205);
or U11405 (N_11405,N_11235,N_11183);
and U11406 (N_11406,N_11062,N_11068);
xnor U11407 (N_11407,N_11106,N_11048);
xor U11408 (N_11408,N_11146,N_11016);
and U11409 (N_11409,N_11127,N_11043);
nand U11410 (N_11410,N_11029,N_11139);
xnor U11411 (N_11411,N_11152,N_11177);
or U11412 (N_11412,N_11224,N_11052);
xnor U11413 (N_11413,N_11177,N_11122);
or U11414 (N_11414,N_11098,N_11189);
or U11415 (N_11415,N_11130,N_11016);
xnor U11416 (N_11416,N_11118,N_11216);
and U11417 (N_11417,N_11006,N_11132);
and U11418 (N_11418,N_11204,N_11144);
xor U11419 (N_11419,N_11017,N_11004);
nand U11420 (N_11420,N_11145,N_11235);
or U11421 (N_11421,N_11051,N_11033);
nor U11422 (N_11422,N_11209,N_11011);
nand U11423 (N_11423,N_11235,N_11166);
nand U11424 (N_11424,N_11061,N_11009);
nor U11425 (N_11425,N_11008,N_11169);
or U11426 (N_11426,N_11215,N_11236);
and U11427 (N_11427,N_11186,N_11038);
xor U11428 (N_11428,N_11211,N_11220);
nor U11429 (N_11429,N_11000,N_11025);
nand U11430 (N_11430,N_11018,N_11080);
xor U11431 (N_11431,N_11097,N_11199);
nand U11432 (N_11432,N_11120,N_11034);
xor U11433 (N_11433,N_11159,N_11183);
and U11434 (N_11434,N_11214,N_11074);
and U11435 (N_11435,N_11067,N_11232);
xnor U11436 (N_11436,N_11216,N_11026);
and U11437 (N_11437,N_11099,N_11218);
nand U11438 (N_11438,N_11240,N_11030);
or U11439 (N_11439,N_11055,N_11046);
xnor U11440 (N_11440,N_11025,N_11248);
nor U11441 (N_11441,N_11142,N_11023);
xor U11442 (N_11442,N_11070,N_11081);
or U11443 (N_11443,N_11189,N_11017);
and U11444 (N_11444,N_11242,N_11066);
and U11445 (N_11445,N_11001,N_11000);
xnor U11446 (N_11446,N_11098,N_11013);
or U11447 (N_11447,N_11083,N_11025);
nor U11448 (N_11448,N_11206,N_11079);
nand U11449 (N_11449,N_11106,N_11039);
xnor U11450 (N_11450,N_11183,N_11177);
and U11451 (N_11451,N_11176,N_11118);
nor U11452 (N_11452,N_11030,N_11243);
xor U11453 (N_11453,N_11190,N_11192);
and U11454 (N_11454,N_11201,N_11142);
and U11455 (N_11455,N_11058,N_11184);
xnor U11456 (N_11456,N_11179,N_11127);
or U11457 (N_11457,N_11094,N_11121);
and U11458 (N_11458,N_11224,N_11102);
nand U11459 (N_11459,N_11001,N_11042);
nand U11460 (N_11460,N_11014,N_11182);
xor U11461 (N_11461,N_11057,N_11095);
or U11462 (N_11462,N_11183,N_11097);
nand U11463 (N_11463,N_11090,N_11081);
and U11464 (N_11464,N_11182,N_11224);
or U11465 (N_11465,N_11241,N_11084);
and U11466 (N_11466,N_11084,N_11159);
xnor U11467 (N_11467,N_11079,N_11221);
nand U11468 (N_11468,N_11072,N_11001);
or U11469 (N_11469,N_11058,N_11114);
nor U11470 (N_11470,N_11247,N_11191);
nand U11471 (N_11471,N_11150,N_11186);
and U11472 (N_11472,N_11239,N_11082);
xor U11473 (N_11473,N_11229,N_11163);
nand U11474 (N_11474,N_11005,N_11034);
or U11475 (N_11475,N_11088,N_11198);
and U11476 (N_11476,N_11145,N_11056);
xnor U11477 (N_11477,N_11248,N_11165);
nor U11478 (N_11478,N_11108,N_11045);
nor U11479 (N_11479,N_11072,N_11153);
nand U11480 (N_11480,N_11092,N_11011);
nor U11481 (N_11481,N_11045,N_11168);
or U11482 (N_11482,N_11177,N_11157);
or U11483 (N_11483,N_11162,N_11158);
xnor U11484 (N_11484,N_11048,N_11123);
nand U11485 (N_11485,N_11185,N_11220);
nand U11486 (N_11486,N_11173,N_11120);
nand U11487 (N_11487,N_11063,N_11073);
nand U11488 (N_11488,N_11183,N_11196);
xor U11489 (N_11489,N_11214,N_11112);
nand U11490 (N_11490,N_11127,N_11042);
xnor U11491 (N_11491,N_11027,N_11082);
or U11492 (N_11492,N_11103,N_11112);
nor U11493 (N_11493,N_11128,N_11209);
nand U11494 (N_11494,N_11094,N_11211);
or U11495 (N_11495,N_11203,N_11024);
xnor U11496 (N_11496,N_11151,N_11230);
nand U11497 (N_11497,N_11057,N_11122);
xnor U11498 (N_11498,N_11249,N_11019);
or U11499 (N_11499,N_11051,N_11235);
xor U11500 (N_11500,N_11324,N_11296);
nor U11501 (N_11501,N_11299,N_11266);
xor U11502 (N_11502,N_11430,N_11273);
xnor U11503 (N_11503,N_11347,N_11252);
and U11504 (N_11504,N_11307,N_11354);
nor U11505 (N_11505,N_11353,N_11436);
or U11506 (N_11506,N_11297,N_11407);
or U11507 (N_11507,N_11253,N_11272);
xnor U11508 (N_11508,N_11348,N_11270);
or U11509 (N_11509,N_11326,N_11455);
xnor U11510 (N_11510,N_11300,N_11284);
and U11511 (N_11511,N_11325,N_11370);
xor U11512 (N_11512,N_11308,N_11342);
xnor U11513 (N_11513,N_11495,N_11489);
and U11514 (N_11514,N_11352,N_11408);
nand U11515 (N_11515,N_11496,N_11264);
nor U11516 (N_11516,N_11334,N_11360);
nor U11517 (N_11517,N_11323,N_11446);
and U11518 (N_11518,N_11403,N_11485);
nand U11519 (N_11519,N_11406,N_11368);
xor U11520 (N_11520,N_11410,N_11311);
xnor U11521 (N_11521,N_11423,N_11336);
or U11522 (N_11522,N_11305,N_11490);
nor U11523 (N_11523,N_11271,N_11429);
and U11524 (N_11524,N_11498,N_11391);
nor U11525 (N_11525,N_11465,N_11486);
and U11526 (N_11526,N_11442,N_11255);
and U11527 (N_11527,N_11349,N_11285);
or U11528 (N_11528,N_11369,N_11474);
xor U11529 (N_11529,N_11457,N_11383);
xnor U11530 (N_11530,N_11394,N_11427);
and U11531 (N_11531,N_11425,N_11293);
or U11532 (N_11532,N_11361,N_11301);
nand U11533 (N_11533,N_11364,N_11363);
nor U11534 (N_11534,N_11335,N_11276);
xnor U11535 (N_11535,N_11473,N_11309);
and U11536 (N_11536,N_11450,N_11268);
xor U11537 (N_11537,N_11393,N_11290);
nor U11538 (N_11538,N_11413,N_11351);
nand U11539 (N_11539,N_11447,N_11438);
xor U11540 (N_11540,N_11404,N_11289);
nor U11541 (N_11541,N_11357,N_11390);
and U11542 (N_11542,N_11459,N_11461);
and U11543 (N_11543,N_11462,N_11437);
and U11544 (N_11544,N_11366,N_11345);
nor U11545 (N_11545,N_11322,N_11350);
and U11546 (N_11546,N_11303,N_11478);
xnor U11547 (N_11547,N_11471,N_11267);
xor U11548 (N_11548,N_11260,N_11392);
nor U11549 (N_11549,N_11286,N_11330);
xor U11550 (N_11550,N_11332,N_11338);
or U11551 (N_11551,N_11416,N_11304);
and U11552 (N_11552,N_11463,N_11343);
xnor U11553 (N_11553,N_11374,N_11379);
nand U11554 (N_11554,N_11265,N_11414);
nor U11555 (N_11555,N_11439,N_11456);
or U11556 (N_11556,N_11470,N_11451);
or U11557 (N_11557,N_11420,N_11306);
nand U11558 (N_11558,N_11344,N_11275);
and U11559 (N_11559,N_11281,N_11481);
nand U11560 (N_11560,N_11313,N_11399);
nand U11561 (N_11561,N_11431,N_11328);
nor U11562 (N_11562,N_11458,N_11402);
or U11563 (N_11563,N_11319,N_11434);
or U11564 (N_11564,N_11411,N_11251);
nor U11565 (N_11565,N_11445,N_11375);
xnor U11566 (N_11566,N_11405,N_11460);
nand U11567 (N_11567,N_11254,N_11329);
and U11568 (N_11568,N_11466,N_11278);
nand U11569 (N_11569,N_11424,N_11356);
or U11570 (N_11570,N_11483,N_11387);
nor U11571 (N_11571,N_11441,N_11401);
or U11572 (N_11572,N_11341,N_11422);
or U11573 (N_11573,N_11380,N_11453);
or U11574 (N_11574,N_11487,N_11385);
nand U11575 (N_11575,N_11476,N_11475);
nor U11576 (N_11576,N_11372,N_11454);
nand U11577 (N_11577,N_11378,N_11467);
or U11578 (N_11578,N_11321,N_11362);
and U11579 (N_11579,N_11376,N_11283);
or U11580 (N_11580,N_11365,N_11440);
xor U11581 (N_11581,N_11274,N_11320);
nand U11582 (N_11582,N_11432,N_11256);
and U11583 (N_11583,N_11409,N_11398);
nor U11584 (N_11584,N_11250,N_11288);
and U11585 (N_11585,N_11400,N_11417);
nor U11586 (N_11586,N_11371,N_11415);
and U11587 (N_11587,N_11295,N_11488);
and U11588 (N_11588,N_11479,N_11384);
nor U11589 (N_11589,N_11314,N_11279);
or U11590 (N_11590,N_11449,N_11492);
xor U11591 (N_11591,N_11317,N_11382);
or U11592 (N_11592,N_11358,N_11497);
or U11593 (N_11593,N_11426,N_11386);
xor U11594 (N_11594,N_11355,N_11421);
and U11595 (N_11595,N_11294,N_11482);
or U11596 (N_11596,N_11395,N_11277);
nand U11597 (N_11597,N_11477,N_11396);
nand U11598 (N_11598,N_11418,N_11412);
xor U11599 (N_11599,N_11339,N_11315);
nand U11600 (N_11600,N_11428,N_11263);
nand U11601 (N_11601,N_11359,N_11435);
xnor U11602 (N_11602,N_11494,N_11291);
and U11603 (N_11603,N_11302,N_11484);
and U11604 (N_11604,N_11397,N_11389);
and U11605 (N_11605,N_11333,N_11377);
and U11606 (N_11606,N_11327,N_11282);
xor U11607 (N_11607,N_11257,N_11337);
nand U11608 (N_11608,N_11310,N_11318);
nand U11609 (N_11609,N_11381,N_11443);
nand U11610 (N_11610,N_11452,N_11448);
and U11611 (N_11611,N_11388,N_11499);
and U11612 (N_11612,N_11493,N_11261);
and U11613 (N_11613,N_11491,N_11269);
and U11614 (N_11614,N_11258,N_11469);
or U11615 (N_11615,N_11346,N_11340);
and U11616 (N_11616,N_11367,N_11262);
and U11617 (N_11617,N_11312,N_11464);
nor U11618 (N_11618,N_11287,N_11433);
and U11619 (N_11619,N_11292,N_11419);
or U11620 (N_11620,N_11373,N_11444);
xor U11621 (N_11621,N_11316,N_11331);
nand U11622 (N_11622,N_11480,N_11472);
or U11623 (N_11623,N_11280,N_11259);
or U11624 (N_11624,N_11468,N_11298);
nand U11625 (N_11625,N_11423,N_11434);
or U11626 (N_11626,N_11291,N_11387);
and U11627 (N_11627,N_11348,N_11315);
nand U11628 (N_11628,N_11438,N_11381);
and U11629 (N_11629,N_11358,N_11303);
nor U11630 (N_11630,N_11386,N_11350);
nor U11631 (N_11631,N_11288,N_11419);
nand U11632 (N_11632,N_11436,N_11449);
or U11633 (N_11633,N_11264,N_11469);
nor U11634 (N_11634,N_11498,N_11463);
nand U11635 (N_11635,N_11381,N_11399);
and U11636 (N_11636,N_11312,N_11320);
or U11637 (N_11637,N_11275,N_11456);
nor U11638 (N_11638,N_11343,N_11250);
nand U11639 (N_11639,N_11266,N_11398);
nor U11640 (N_11640,N_11293,N_11421);
and U11641 (N_11641,N_11349,N_11389);
nand U11642 (N_11642,N_11411,N_11252);
and U11643 (N_11643,N_11464,N_11403);
nand U11644 (N_11644,N_11447,N_11321);
nor U11645 (N_11645,N_11445,N_11385);
or U11646 (N_11646,N_11430,N_11256);
and U11647 (N_11647,N_11259,N_11482);
nor U11648 (N_11648,N_11266,N_11344);
nand U11649 (N_11649,N_11337,N_11497);
nor U11650 (N_11650,N_11266,N_11491);
nand U11651 (N_11651,N_11414,N_11267);
nor U11652 (N_11652,N_11418,N_11272);
nor U11653 (N_11653,N_11450,N_11498);
nand U11654 (N_11654,N_11463,N_11435);
nand U11655 (N_11655,N_11380,N_11335);
and U11656 (N_11656,N_11475,N_11281);
nor U11657 (N_11657,N_11341,N_11340);
nor U11658 (N_11658,N_11467,N_11344);
and U11659 (N_11659,N_11459,N_11302);
nand U11660 (N_11660,N_11351,N_11268);
nor U11661 (N_11661,N_11398,N_11450);
or U11662 (N_11662,N_11468,N_11417);
and U11663 (N_11663,N_11395,N_11334);
xor U11664 (N_11664,N_11460,N_11293);
nand U11665 (N_11665,N_11391,N_11269);
xor U11666 (N_11666,N_11311,N_11381);
or U11667 (N_11667,N_11321,N_11275);
and U11668 (N_11668,N_11396,N_11258);
nor U11669 (N_11669,N_11443,N_11402);
nand U11670 (N_11670,N_11490,N_11373);
xor U11671 (N_11671,N_11336,N_11486);
or U11672 (N_11672,N_11403,N_11380);
or U11673 (N_11673,N_11449,N_11441);
nand U11674 (N_11674,N_11288,N_11357);
xor U11675 (N_11675,N_11430,N_11373);
nor U11676 (N_11676,N_11369,N_11456);
and U11677 (N_11677,N_11467,N_11357);
nor U11678 (N_11678,N_11386,N_11377);
or U11679 (N_11679,N_11257,N_11327);
xnor U11680 (N_11680,N_11331,N_11262);
or U11681 (N_11681,N_11288,N_11428);
and U11682 (N_11682,N_11418,N_11316);
nand U11683 (N_11683,N_11364,N_11486);
nor U11684 (N_11684,N_11441,N_11313);
nand U11685 (N_11685,N_11290,N_11427);
nand U11686 (N_11686,N_11267,N_11346);
and U11687 (N_11687,N_11313,N_11469);
xor U11688 (N_11688,N_11419,N_11450);
nor U11689 (N_11689,N_11459,N_11254);
and U11690 (N_11690,N_11471,N_11343);
or U11691 (N_11691,N_11416,N_11462);
and U11692 (N_11692,N_11431,N_11446);
nor U11693 (N_11693,N_11367,N_11321);
or U11694 (N_11694,N_11383,N_11277);
or U11695 (N_11695,N_11275,N_11411);
nand U11696 (N_11696,N_11328,N_11286);
nor U11697 (N_11697,N_11325,N_11279);
nor U11698 (N_11698,N_11410,N_11388);
xnor U11699 (N_11699,N_11472,N_11481);
xnor U11700 (N_11700,N_11401,N_11402);
nand U11701 (N_11701,N_11251,N_11300);
nor U11702 (N_11702,N_11443,N_11280);
nor U11703 (N_11703,N_11384,N_11408);
or U11704 (N_11704,N_11488,N_11414);
or U11705 (N_11705,N_11445,N_11443);
xnor U11706 (N_11706,N_11421,N_11335);
xnor U11707 (N_11707,N_11330,N_11407);
and U11708 (N_11708,N_11257,N_11306);
nor U11709 (N_11709,N_11404,N_11297);
nor U11710 (N_11710,N_11308,N_11323);
and U11711 (N_11711,N_11372,N_11387);
nor U11712 (N_11712,N_11411,N_11304);
and U11713 (N_11713,N_11277,N_11263);
xnor U11714 (N_11714,N_11421,N_11369);
nor U11715 (N_11715,N_11322,N_11374);
or U11716 (N_11716,N_11354,N_11315);
xnor U11717 (N_11717,N_11364,N_11465);
nor U11718 (N_11718,N_11269,N_11380);
or U11719 (N_11719,N_11450,N_11438);
or U11720 (N_11720,N_11365,N_11470);
and U11721 (N_11721,N_11448,N_11360);
nor U11722 (N_11722,N_11367,N_11383);
nand U11723 (N_11723,N_11366,N_11464);
xor U11724 (N_11724,N_11490,N_11277);
and U11725 (N_11725,N_11275,N_11493);
nand U11726 (N_11726,N_11423,N_11256);
nand U11727 (N_11727,N_11350,N_11440);
or U11728 (N_11728,N_11417,N_11367);
or U11729 (N_11729,N_11480,N_11415);
and U11730 (N_11730,N_11463,N_11399);
or U11731 (N_11731,N_11393,N_11442);
and U11732 (N_11732,N_11388,N_11441);
nor U11733 (N_11733,N_11431,N_11450);
xnor U11734 (N_11734,N_11464,N_11381);
xnor U11735 (N_11735,N_11284,N_11430);
or U11736 (N_11736,N_11451,N_11458);
and U11737 (N_11737,N_11344,N_11428);
and U11738 (N_11738,N_11257,N_11253);
nor U11739 (N_11739,N_11408,N_11292);
nor U11740 (N_11740,N_11332,N_11303);
nor U11741 (N_11741,N_11397,N_11441);
nor U11742 (N_11742,N_11398,N_11376);
or U11743 (N_11743,N_11316,N_11401);
nand U11744 (N_11744,N_11260,N_11383);
and U11745 (N_11745,N_11371,N_11388);
nor U11746 (N_11746,N_11310,N_11400);
or U11747 (N_11747,N_11331,N_11416);
nor U11748 (N_11748,N_11405,N_11468);
and U11749 (N_11749,N_11447,N_11414);
nor U11750 (N_11750,N_11550,N_11706);
or U11751 (N_11751,N_11566,N_11675);
nand U11752 (N_11752,N_11739,N_11563);
xnor U11753 (N_11753,N_11527,N_11578);
or U11754 (N_11754,N_11510,N_11542);
or U11755 (N_11755,N_11579,N_11624);
nor U11756 (N_11756,N_11569,N_11680);
nand U11757 (N_11757,N_11657,N_11714);
nand U11758 (N_11758,N_11523,N_11532);
nor U11759 (N_11759,N_11695,N_11726);
nor U11760 (N_11760,N_11520,N_11728);
or U11761 (N_11761,N_11685,N_11522);
and U11762 (N_11762,N_11646,N_11678);
nand U11763 (N_11763,N_11628,N_11727);
and U11764 (N_11764,N_11537,N_11749);
nand U11765 (N_11765,N_11744,N_11748);
nor U11766 (N_11766,N_11591,N_11610);
nor U11767 (N_11767,N_11570,N_11576);
and U11768 (N_11768,N_11588,N_11710);
nor U11769 (N_11769,N_11590,N_11604);
and U11770 (N_11770,N_11630,N_11546);
and U11771 (N_11771,N_11572,N_11717);
nor U11772 (N_11772,N_11612,N_11666);
xnor U11773 (N_11773,N_11650,N_11512);
or U11774 (N_11774,N_11691,N_11644);
or U11775 (N_11775,N_11557,N_11683);
or U11776 (N_11776,N_11515,N_11559);
or U11777 (N_11777,N_11554,N_11609);
xor U11778 (N_11778,N_11519,N_11545);
nand U11779 (N_11779,N_11541,N_11525);
nand U11780 (N_11780,N_11614,N_11524);
nor U11781 (N_11781,N_11551,N_11712);
or U11782 (N_11782,N_11533,N_11705);
or U11783 (N_11783,N_11632,N_11703);
or U11784 (N_11784,N_11702,N_11692);
xnor U11785 (N_11785,N_11682,N_11643);
nand U11786 (N_11786,N_11668,N_11608);
nand U11787 (N_11787,N_11679,N_11531);
xor U11788 (N_11788,N_11638,N_11677);
or U11789 (N_11789,N_11742,N_11645);
nor U11790 (N_11790,N_11556,N_11656);
or U11791 (N_11791,N_11725,N_11652);
nand U11792 (N_11792,N_11582,N_11599);
nor U11793 (N_11793,N_11504,N_11711);
or U11794 (N_11794,N_11697,N_11625);
nand U11795 (N_11795,N_11740,N_11509);
xnor U11796 (N_11796,N_11659,N_11704);
and U11797 (N_11797,N_11672,N_11639);
or U11798 (N_11798,N_11693,N_11687);
or U11799 (N_11799,N_11664,N_11626);
nand U11800 (N_11800,N_11513,N_11539);
nor U11801 (N_11801,N_11648,N_11611);
or U11802 (N_11802,N_11634,N_11535);
nor U11803 (N_11803,N_11631,N_11745);
nand U11804 (N_11804,N_11660,N_11642);
and U11805 (N_11805,N_11686,N_11589);
and U11806 (N_11806,N_11577,N_11701);
xor U11807 (N_11807,N_11681,N_11688);
nor U11808 (N_11808,N_11731,N_11581);
nand U11809 (N_11809,N_11637,N_11501);
or U11810 (N_11810,N_11586,N_11720);
or U11811 (N_11811,N_11561,N_11508);
nand U11812 (N_11812,N_11615,N_11698);
xor U11813 (N_11813,N_11558,N_11635);
or U11814 (N_11814,N_11506,N_11584);
or U11815 (N_11815,N_11516,N_11735);
or U11816 (N_11816,N_11700,N_11517);
nand U11817 (N_11817,N_11560,N_11732);
xnor U11818 (N_11818,N_11548,N_11596);
nand U11819 (N_11819,N_11715,N_11647);
xnor U11820 (N_11820,N_11721,N_11511);
or U11821 (N_11821,N_11674,N_11734);
and U11822 (N_11822,N_11503,N_11518);
and U11823 (N_11823,N_11594,N_11676);
nand U11824 (N_11824,N_11738,N_11724);
and U11825 (N_11825,N_11514,N_11536);
or U11826 (N_11826,N_11661,N_11730);
or U11827 (N_11827,N_11694,N_11530);
xor U11828 (N_11828,N_11529,N_11593);
xnor U11829 (N_11829,N_11587,N_11565);
nor U11830 (N_11830,N_11592,N_11607);
nand U11831 (N_11831,N_11708,N_11633);
and U11832 (N_11832,N_11696,N_11667);
nand U11833 (N_11833,N_11616,N_11665);
and U11834 (N_11834,N_11621,N_11567);
xnor U11835 (N_11835,N_11534,N_11719);
and U11836 (N_11836,N_11640,N_11574);
nor U11837 (N_11837,N_11620,N_11543);
nand U11838 (N_11838,N_11601,N_11619);
and U11839 (N_11839,N_11564,N_11746);
nor U11840 (N_11840,N_11636,N_11658);
or U11841 (N_11841,N_11617,N_11598);
or U11842 (N_11842,N_11709,N_11741);
xnor U11843 (N_11843,N_11583,N_11654);
nor U11844 (N_11844,N_11690,N_11733);
nand U11845 (N_11845,N_11549,N_11526);
and U11846 (N_11846,N_11653,N_11505);
nand U11847 (N_11847,N_11575,N_11580);
or U11848 (N_11848,N_11718,N_11544);
xor U11849 (N_11849,N_11613,N_11605);
and U11850 (N_11850,N_11600,N_11538);
nor U11851 (N_11851,N_11670,N_11671);
and U11852 (N_11852,N_11540,N_11716);
or U11853 (N_11853,N_11618,N_11562);
xnor U11854 (N_11854,N_11622,N_11585);
xnor U11855 (N_11855,N_11673,N_11736);
xor U11856 (N_11856,N_11651,N_11713);
nand U11857 (N_11857,N_11722,N_11729);
nand U11858 (N_11858,N_11603,N_11553);
xnor U11859 (N_11859,N_11547,N_11552);
or U11860 (N_11860,N_11571,N_11663);
nor U11861 (N_11861,N_11723,N_11502);
xor U11862 (N_11862,N_11606,N_11595);
xor U11863 (N_11863,N_11655,N_11555);
nor U11864 (N_11864,N_11641,N_11623);
or U11865 (N_11865,N_11662,N_11507);
nand U11866 (N_11866,N_11684,N_11707);
and U11867 (N_11867,N_11528,N_11568);
nor U11868 (N_11868,N_11573,N_11627);
and U11869 (N_11869,N_11737,N_11689);
nand U11870 (N_11870,N_11747,N_11699);
and U11871 (N_11871,N_11743,N_11649);
or U11872 (N_11872,N_11629,N_11597);
xor U11873 (N_11873,N_11521,N_11602);
xnor U11874 (N_11874,N_11500,N_11669);
xor U11875 (N_11875,N_11510,N_11601);
xor U11876 (N_11876,N_11730,N_11728);
and U11877 (N_11877,N_11601,N_11706);
xor U11878 (N_11878,N_11616,N_11551);
nor U11879 (N_11879,N_11662,N_11603);
and U11880 (N_11880,N_11736,N_11524);
nor U11881 (N_11881,N_11706,N_11500);
nand U11882 (N_11882,N_11544,N_11652);
nand U11883 (N_11883,N_11741,N_11730);
or U11884 (N_11884,N_11533,N_11728);
xnor U11885 (N_11885,N_11729,N_11584);
nor U11886 (N_11886,N_11550,N_11530);
or U11887 (N_11887,N_11616,N_11684);
nand U11888 (N_11888,N_11573,N_11602);
and U11889 (N_11889,N_11535,N_11567);
and U11890 (N_11890,N_11541,N_11659);
and U11891 (N_11891,N_11706,N_11684);
and U11892 (N_11892,N_11665,N_11745);
nor U11893 (N_11893,N_11632,N_11598);
nor U11894 (N_11894,N_11560,N_11702);
or U11895 (N_11895,N_11538,N_11618);
nand U11896 (N_11896,N_11702,N_11589);
or U11897 (N_11897,N_11534,N_11559);
or U11898 (N_11898,N_11679,N_11621);
nor U11899 (N_11899,N_11630,N_11713);
xnor U11900 (N_11900,N_11575,N_11739);
or U11901 (N_11901,N_11746,N_11653);
and U11902 (N_11902,N_11613,N_11688);
nand U11903 (N_11903,N_11546,N_11731);
and U11904 (N_11904,N_11504,N_11598);
or U11905 (N_11905,N_11582,N_11547);
xnor U11906 (N_11906,N_11525,N_11679);
xnor U11907 (N_11907,N_11695,N_11574);
xnor U11908 (N_11908,N_11557,N_11591);
nand U11909 (N_11909,N_11606,N_11655);
nand U11910 (N_11910,N_11670,N_11548);
xor U11911 (N_11911,N_11654,N_11670);
nor U11912 (N_11912,N_11508,N_11644);
or U11913 (N_11913,N_11527,N_11519);
or U11914 (N_11914,N_11634,N_11637);
xnor U11915 (N_11915,N_11705,N_11608);
nor U11916 (N_11916,N_11559,N_11563);
and U11917 (N_11917,N_11539,N_11527);
or U11918 (N_11918,N_11717,N_11748);
or U11919 (N_11919,N_11587,N_11518);
or U11920 (N_11920,N_11566,N_11734);
xor U11921 (N_11921,N_11643,N_11679);
xor U11922 (N_11922,N_11523,N_11698);
and U11923 (N_11923,N_11524,N_11521);
and U11924 (N_11924,N_11632,N_11669);
nor U11925 (N_11925,N_11563,N_11687);
or U11926 (N_11926,N_11694,N_11586);
xor U11927 (N_11927,N_11630,N_11553);
and U11928 (N_11928,N_11639,N_11589);
and U11929 (N_11929,N_11521,N_11713);
nor U11930 (N_11930,N_11647,N_11623);
nor U11931 (N_11931,N_11711,N_11609);
or U11932 (N_11932,N_11593,N_11626);
and U11933 (N_11933,N_11634,N_11742);
xnor U11934 (N_11934,N_11694,N_11650);
or U11935 (N_11935,N_11593,N_11670);
nor U11936 (N_11936,N_11740,N_11624);
nor U11937 (N_11937,N_11596,N_11727);
or U11938 (N_11938,N_11739,N_11617);
or U11939 (N_11939,N_11621,N_11534);
xor U11940 (N_11940,N_11725,N_11551);
xnor U11941 (N_11941,N_11700,N_11643);
and U11942 (N_11942,N_11729,N_11554);
xor U11943 (N_11943,N_11574,N_11680);
xor U11944 (N_11944,N_11686,N_11515);
xor U11945 (N_11945,N_11673,N_11611);
or U11946 (N_11946,N_11559,N_11651);
xor U11947 (N_11947,N_11732,N_11601);
nand U11948 (N_11948,N_11583,N_11744);
xnor U11949 (N_11949,N_11602,N_11628);
xnor U11950 (N_11950,N_11581,N_11500);
xor U11951 (N_11951,N_11555,N_11554);
or U11952 (N_11952,N_11738,N_11607);
xor U11953 (N_11953,N_11531,N_11600);
or U11954 (N_11954,N_11595,N_11738);
nand U11955 (N_11955,N_11525,N_11565);
xor U11956 (N_11956,N_11606,N_11604);
and U11957 (N_11957,N_11617,N_11628);
xnor U11958 (N_11958,N_11721,N_11677);
or U11959 (N_11959,N_11692,N_11555);
and U11960 (N_11960,N_11706,N_11638);
nand U11961 (N_11961,N_11595,N_11727);
xnor U11962 (N_11962,N_11616,N_11618);
xor U11963 (N_11963,N_11589,N_11713);
and U11964 (N_11964,N_11688,N_11521);
xnor U11965 (N_11965,N_11564,N_11683);
or U11966 (N_11966,N_11704,N_11747);
nand U11967 (N_11967,N_11631,N_11652);
nor U11968 (N_11968,N_11511,N_11610);
nor U11969 (N_11969,N_11647,N_11620);
or U11970 (N_11970,N_11569,N_11662);
or U11971 (N_11971,N_11612,N_11594);
or U11972 (N_11972,N_11696,N_11636);
or U11973 (N_11973,N_11584,N_11720);
nand U11974 (N_11974,N_11536,N_11589);
or U11975 (N_11975,N_11659,N_11557);
xnor U11976 (N_11976,N_11708,N_11677);
nor U11977 (N_11977,N_11621,N_11525);
nor U11978 (N_11978,N_11506,N_11740);
and U11979 (N_11979,N_11539,N_11664);
and U11980 (N_11980,N_11683,N_11735);
nor U11981 (N_11981,N_11643,N_11740);
or U11982 (N_11982,N_11699,N_11671);
xnor U11983 (N_11983,N_11724,N_11630);
xnor U11984 (N_11984,N_11574,N_11525);
xor U11985 (N_11985,N_11535,N_11655);
nor U11986 (N_11986,N_11544,N_11517);
nand U11987 (N_11987,N_11605,N_11739);
nand U11988 (N_11988,N_11559,N_11655);
nor U11989 (N_11989,N_11652,N_11684);
or U11990 (N_11990,N_11576,N_11716);
and U11991 (N_11991,N_11636,N_11703);
or U11992 (N_11992,N_11729,N_11626);
or U11993 (N_11993,N_11742,N_11726);
xnor U11994 (N_11994,N_11637,N_11554);
and U11995 (N_11995,N_11623,N_11595);
or U11996 (N_11996,N_11672,N_11533);
xor U11997 (N_11997,N_11560,N_11656);
nand U11998 (N_11998,N_11578,N_11628);
or U11999 (N_11999,N_11667,N_11510);
nor U12000 (N_12000,N_11880,N_11973);
or U12001 (N_12001,N_11947,N_11783);
nand U12002 (N_12002,N_11954,N_11891);
or U12003 (N_12003,N_11917,N_11799);
nand U12004 (N_12004,N_11923,N_11805);
and U12005 (N_12005,N_11931,N_11804);
nor U12006 (N_12006,N_11769,N_11786);
nor U12007 (N_12007,N_11965,N_11844);
xnor U12008 (N_12008,N_11985,N_11918);
and U12009 (N_12009,N_11991,N_11776);
nor U12010 (N_12010,N_11790,N_11757);
and U12011 (N_12011,N_11955,N_11910);
nand U12012 (N_12012,N_11766,N_11849);
nand U12013 (N_12013,N_11946,N_11868);
nand U12014 (N_12014,N_11759,N_11814);
or U12015 (N_12015,N_11861,N_11831);
nand U12016 (N_12016,N_11961,N_11881);
or U12017 (N_12017,N_11984,N_11960);
nor U12018 (N_12018,N_11934,N_11884);
nor U12019 (N_12019,N_11981,N_11808);
nor U12020 (N_12020,N_11887,N_11930);
nor U12021 (N_12021,N_11760,N_11850);
or U12022 (N_12022,N_11939,N_11969);
xor U12023 (N_12023,N_11926,N_11924);
nor U12024 (N_12024,N_11854,N_11911);
or U12025 (N_12025,N_11784,N_11837);
nor U12026 (N_12026,N_11750,N_11990);
nor U12027 (N_12027,N_11879,N_11885);
xnor U12028 (N_12028,N_11865,N_11864);
nand U12029 (N_12029,N_11975,N_11795);
nand U12030 (N_12030,N_11839,N_11970);
nand U12031 (N_12031,N_11972,N_11945);
xnor U12032 (N_12032,N_11978,N_11919);
nand U12033 (N_12033,N_11904,N_11830);
or U12034 (N_12034,N_11895,N_11983);
xnor U12035 (N_12035,N_11761,N_11798);
or U12036 (N_12036,N_11986,N_11922);
or U12037 (N_12037,N_11883,N_11770);
nor U12038 (N_12038,N_11936,N_11998);
nor U12039 (N_12039,N_11807,N_11822);
nor U12040 (N_12040,N_11820,N_11901);
or U12041 (N_12041,N_11905,N_11863);
nor U12042 (N_12042,N_11828,N_11894);
nand U12043 (N_12043,N_11855,N_11823);
or U12044 (N_12044,N_11779,N_11796);
or U12045 (N_12045,N_11780,N_11900);
xor U12046 (N_12046,N_11815,N_11942);
and U12047 (N_12047,N_11778,N_11755);
nor U12048 (N_12048,N_11812,N_11834);
and U12049 (N_12049,N_11892,N_11829);
or U12050 (N_12050,N_11912,N_11940);
nor U12051 (N_12051,N_11857,N_11789);
nand U12052 (N_12052,N_11771,N_11943);
nand U12053 (N_12053,N_11791,N_11897);
or U12054 (N_12054,N_11803,N_11772);
or U12055 (N_12055,N_11836,N_11764);
nand U12056 (N_12056,N_11751,N_11874);
nor U12057 (N_12057,N_11898,N_11792);
nor U12058 (N_12058,N_11956,N_11997);
and U12059 (N_12059,N_11852,N_11754);
nor U12060 (N_12060,N_11915,N_11878);
nor U12061 (N_12061,N_11862,N_11979);
nand U12062 (N_12062,N_11909,N_11976);
and U12063 (N_12063,N_11818,N_11843);
and U12064 (N_12064,N_11993,N_11819);
nor U12065 (N_12065,N_11873,N_11841);
xor U12066 (N_12066,N_11999,N_11925);
or U12067 (N_12067,N_11952,N_11893);
and U12068 (N_12068,N_11914,N_11968);
nor U12069 (N_12069,N_11860,N_11949);
and U12070 (N_12070,N_11788,N_11962);
xnor U12071 (N_12071,N_11906,N_11963);
or U12072 (N_12072,N_11869,N_11756);
xor U12073 (N_12073,N_11765,N_11775);
nor U12074 (N_12074,N_11762,N_11948);
xnor U12075 (N_12075,N_11838,N_11957);
and U12076 (N_12076,N_11824,N_11802);
nor U12077 (N_12077,N_11980,N_11890);
nand U12078 (N_12078,N_11982,N_11781);
and U12079 (N_12079,N_11950,N_11817);
and U12080 (N_12080,N_11937,N_11842);
and U12081 (N_12081,N_11899,N_11995);
and U12082 (N_12082,N_11951,N_11964);
or U12083 (N_12083,N_11959,N_11845);
or U12084 (N_12084,N_11941,N_11929);
or U12085 (N_12085,N_11816,N_11763);
nor U12086 (N_12086,N_11938,N_11928);
xor U12087 (N_12087,N_11867,N_11787);
xnor U12088 (N_12088,N_11859,N_11967);
xnor U12089 (N_12089,N_11752,N_11886);
xnor U12090 (N_12090,N_11870,N_11992);
nand U12091 (N_12091,N_11858,N_11987);
and U12092 (N_12092,N_11913,N_11903);
nor U12093 (N_12093,N_11908,N_11801);
and U12094 (N_12094,N_11809,N_11825);
nor U12095 (N_12095,N_11793,N_11971);
or U12096 (N_12096,N_11996,N_11932);
and U12097 (N_12097,N_11933,N_11773);
and U12098 (N_12098,N_11944,N_11927);
or U12099 (N_12099,N_11835,N_11768);
nor U12100 (N_12100,N_11810,N_11827);
nor U12101 (N_12101,N_11866,N_11774);
and U12102 (N_12102,N_11935,N_11920);
xor U12103 (N_12103,N_11907,N_11851);
nor U12104 (N_12104,N_11758,N_11856);
or U12105 (N_12105,N_11902,N_11953);
nor U12106 (N_12106,N_11958,N_11888);
nor U12107 (N_12107,N_11800,N_11875);
nor U12108 (N_12108,N_11811,N_11797);
and U12109 (N_12109,N_11785,N_11876);
nor U12110 (N_12110,N_11753,N_11989);
and U12111 (N_12111,N_11848,N_11782);
xor U12112 (N_12112,N_11872,N_11794);
and U12113 (N_12113,N_11833,N_11832);
nor U12114 (N_12114,N_11977,N_11840);
or U12115 (N_12115,N_11882,N_11826);
and U12116 (N_12116,N_11853,N_11813);
xor U12117 (N_12117,N_11777,N_11974);
or U12118 (N_12118,N_11988,N_11896);
nand U12119 (N_12119,N_11966,N_11846);
nor U12120 (N_12120,N_11889,N_11994);
nand U12121 (N_12121,N_11847,N_11916);
or U12122 (N_12122,N_11871,N_11921);
or U12123 (N_12123,N_11821,N_11877);
xnor U12124 (N_12124,N_11767,N_11806);
nand U12125 (N_12125,N_11811,N_11862);
xnor U12126 (N_12126,N_11761,N_11961);
and U12127 (N_12127,N_11993,N_11833);
xor U12128 (N_12128,N_11793,N_11963);
nand U12129 (N_12129,N_11971,N_11800);
nand U12130 (N_12130,N_11765,N_11887);
or U12131 (N_12131,N_11829,N_11998);
nor U12132 (N_12132,N_11768,N_11827);
xor U12133 (N_12133,N_11832,N_11766);
nand U12134 (N_12134,N_11872,N_11790);
nor U12135 (N_12135,N_11832,N_11856);
and U12136 (N_12136,N_11944,N_11970);
and U12137 (N_12137,N_11963,N_11842);
xor U12138 (N_12138,N_11896,N_11908);
nor U12139 (N_12139,N_11991,N_11999);
xnor U12140 (N_12140,N_11950,N_11908);
nor U12141 (N_12141,N_11768,N_11956);
nand U12142 (N_12142,N_11847,N_11943);
nand U12143 (N_12143,N_11802,N_11775);
and U12144 (N_12144,N_11945,N_11904);
and U12145 (N_12145,N_11765,N_11795);
and U12146 (N_12146,N_11788,N_11775);
xor U12147 (N_12147,N_11883,N_11938);
or U12148 (N_12148,N_11788,N_11955);
nor U12149 (N_12149,N_11829,N_11910);
or U12150 (N_12150,N_11810,N_11954);
nor U12151 (N_12151,N_11775,N_11764);
nor U12152 (N_12152,N_11999,N_11928);
xor U12153 (N_12153,N_11863,N_11950);
nor U12154 (N_12154,N_11968,N_11886);
nor U12155 (N_12155,N_11974,N_11760);
and U12156 (N_12156,N_11874,N_11817);
and U12157 (N_12157,N_11811,N_11950);
nor U12158 (N_12158,N_11773,N_11830);
xnor U12159 (N_12159,N_11957,N_11882);
xnor U12160 (N_12160,N_11934,N_11946);
nand U12161 (N_12161,N_11871,N_11982);
xnor U12162 (N_12162,N_11770,N_11845);
nor U12163 (N_12163,N_11786,N_11946);
and U12164 (N_12164,N_11877,N_11838);
xor U12165 (N_12165,N_11957,N_11825);
or U12166 (N_12166,N_11957,N_11778);
nand U12167 (N_12167,N_11760,N_11781);
nand U12168 (N_12168,N_11937,N_11979);
and U12169 (N_12169,N_11990,N_11758);
or U12170 (N_12170,N_11790,N_11902);
and U12171 (N_12171,N_11874,N_11832);
nand U12172 (N_12172,N_11842,N_11942);
and U12173 (N_12173,N_11888,N_11910);
and U12174 (N_12174,N_11897,N_11844);
nand U12175 (N_12175,N_11953,N_11954);
and U12176 (N_12176,N_11999,N_11982);
and U12177 (N_12177,N_11977,N_11918);
and U12178 (N_12178,N_11956,N_11763);
nor U12179 (N_12179,N_11872,N_11768);
xnor U12180 (N_12180,N_11914,N_11769);
and U12181 (N_12181,N_11894,N_11792);
xnor U12182 (N_12182,N_11887,N_11828);
xor U12183 (N_12183,N_11962,N_11927);
nand U12184 (N_12184,N_11882,N_11906);
nand U12185 (N_12185,N_11936,N_11860);
xor U12186 (N_12186,N_11867,N_11854);
nand U12187 (N_12187,N_11753,N_11978);
nand U12188 (N_12188,N_11954,N_11977);
nor U12189 (N_12189,N_11763,N_11992);
xor U12190 (N_12190,N_11929,N_11763);
nor U12191 (N_12191,N_11857,N_11866);
nor U12192 (N_12192,N_11797,N_11972);
or U12193 (N_12193,N_11793,N_11878);
or U12194 (N_12194,N_11910,N_11892);
nand U12195 (N_12195,N_11789,N_11876);
or U12196 (N_12196,N_11910,N_11846);
nand U12197 (N_12197,N_11946,N_11864);
or U12198 (N_12198,N_11919,N_11871);
and U12199 (N_12199,N_11818,N_11883);
and U12200 (N_12200,N_11928,N_11873);
and U12201 (N_12201,N_11866,N_11785);
or U12202 (N_12202,N_11818,N_11890);
and U12203 (N_12203,N_11889,N_11778);
nand U12204 (N_12204,N_11915,N_11764);
xnor U12205 (N_12205,N_11985,N_11947);
nor U12206 (N_12206,N_11861,N_11845);
nor U12207 (N_12207,N_11831,N_11844);
xnor U12208 (N_12208,N_11855,N_11903);
nand U12209 (N_12209,N_11872,N_11754);
xnor U12210 (N_12210,N_11934,N_11963);
and U12211 (N_12211,N_11796,N_11753);
xor U12212 (N_12212,N_11875,N_11804);
and U12213 (N_12213,N_11869,N_11914);
xor U12214 (N_12214,N_11764,N_11807);
or U12215 (N_12215,N_11816,N_11850);
nor U12216 (N_12216,N_11936,N_11907);
or U12217 (N_12217,N_11849,N_11884);
and U12218 (N_12218,N_11762,N_11972);
nand U12219 (N_12219,N_11929,N_11858);
or U12220 (N_12220,N_11965,N_11979);
nand U12221 (N_12221,N_11966,N_11773);
nand U12222 (N_12222,N_11803,N_11755);
nor U12223 (N_12223,N_11868,N_11998);
nor U12224 (N_12224,N_11790,N_11888);
xor U12225 (N_12225,N_11882,N_11935);
xor U12226 (N_12226,N_11883,N_11988);
nand U12227 (N_12227,N_11836,N_11935);
nand U12228 (N_12228,N_11969,N_11914);
xnor U12229 (N_12229,N_11948,N_11766);
or U12230 (N_12230,N_11905,N_11802);
or U12231 (N_12231,N_11865,N_11896);
nor U12232 (N_12232,N_11825,N_11981);
nor U12233 (N_12233,N_11887,N_11848);
xnor U12234 (N_12234,N_11909,N_11777);
or U12235 (N_12235,N_11802,N_11887);
nor U12236 (N_12236,N_11931,N_11837);
or U12237 (N_12237,N_11908,N_11930);
or U12238 (N_12238,N_11958,N_11752);
or U12239 (N_12239,N_11943,N_11938);
nand U12240 (N_12240,N_11819,N_11955);
nand U12241 (N_12241,N_11799,N_11866);
xnor U12242 (N_12242,N_11850,N_11970);
nor U12243 (N_12243,N_11931,N_11752);
nor U12244 (N_12244,N_11843,N_11939);
and U12245 (N_12245,N_11816,N_11827);
nor U12246 (N_12246,N_11756,N_11805);
nand U12247 (N_12247,N_11932,N_11788);
and U12248 (N_12248,N_11916,N_11942);
or U12249 (N_12249,N_11937,N_11787);
and U12250 (N_12250,N_12041,N_12110);
and U12251 (N_12251,N_12117,N_12078);
xnor U12252 (N_12252,N_12176,N_12099);
nand U12253 (N_12253,N_12192,N_12040);
or U12254 (N_12254,N_12243,N_12164);
or U12255 (N_12255,N_12057,N_12096);
or U12256 (N_12256,N_12198,N_12014);
nand U12257 (N_12257,N_12240,N_12068);
or U12258 (N_12258,N_12087,N_12021);
xor U12259 (N_12259,N_12215,N_12002);
or U12260 (N_12260,N_12009,N_12107);
xnor U12261 (N_12261,N_12030,N_12058);
nand U12262 (N_12262,N_12154,N_12184);
and U12263 (N_12263,N_12049,N_12221);
nor U12264 (N_12264,N_12042,N_12100);
xnor U12265 (N_12265,N_12060,N_12241);
nor U12266 (N_12266,N_12234,N_12134);
and U12267 (N_12267,N_12151,N_12238);
and U12268 (N_12268,N_12064,N_12138);
or U12269 (N_12269,N_12102,N_12061);
nand U12270 (N_12270,N_12195,N_12210);
nand U12271 (N_12271,N_12051,N_12201);
or U12272 (N_12272,N_12166,N_12065);
or U12273 (N_12273,N_12032,N_12018);
nand U12274 (N_12274,N_12031,N_12092);
nand U12275 (N_12275,N_12098,N_12045);
nor U12276 (N_12276,N_12153,N_12122);
and U12277 (N_12277,N_12205,N_12054);
or U12278 (N_12278,N_12070,N_12039);
and U12279 (N_12279,N_12088,N_12161);
and U12280 (N_12280,N_12026,N_12189);
nand U12281 (N_12281,N_12128,N_12175);
and U12282 (N_12282,N_12015,N_12233);
xor U12283 (N_12283,N_12181,N_12135);
xor U12284 (N_12284,N_12144,N_12199);
xor U12285 (N_12285,N_12187,N_12237);
or U12286 (N_12286,N_12126,N_12007);
xnor U12287 (N_12287,N_12033,N_12095);
nand U12288 (N_12288,N_12114,N_12245);
nor U12289 (N_12289,N_12156,N_12246);
nand U12290 (N_12290,N_12093,N_12071);
nand U12291 (N_12291,N_12214,N_12044);
and U12292 (N_12292,N_12178,N_12216);
and U12293 (N_12293,N_12050,N_12244);
nand U12294 (N_12294,N_12226,N_12196);
xnor U12295 (N_12295,N_12141,N_12121);
or U12296 (N_12296,N_12228,N_12197);
xor U12297 (N_12297,N_12118,N_12011);
or U12298 (N_12298,N_12115,N_12248);
or U12299 (N_12299,N_12174,N_12235);
or U12300 (N_12300,N_12016,N_12206);
xnor U12301 (N_12301,N_12207,N_12162);
and U12302 (N_12302,N_12150,N_12202);
xor U12303 (N_12303,N_12089,N_12209);
nor U12304 (N_12304,N_12193,N_12046);
xnor U12305 (N_12305,N_12085,N_12143);
and U12306 (N_12306,N_12017,N_12230);
and U12307 (N_12307,N_12133,N_12082);
or U12308 (N_12308,N_12113,N_12147);
xor U12309 (N_12309,N_12167,N_12059);
and U12310 (N_12310,N_12169,N_12097);
or U12311 (N_12311,N_12188,N_12010);
xnor U12312 (N_12312,N_12218,N_12006);
xnor U12313 (N_12313,N_12101,N_12180);
xor U12314 (N_12314,N_12223,N_12236);
or U12315 (N_12315,N_12140,N_12247);
xnor U12316 (N_12316,N_12106,N_12047);
nor U12317 (N_12317,N_12112,N_12146);
nand U12318 (N_12318,N_12225,N_12168);
or U12319 (N_12319,N_12079,N_12003);
xor U12320 (N_12320,N_12103,N_12119);
nand U12321 (N_12321,N_12086,N_12022);
xor U12322 (N_12322,N_12067,N_12171);
nand U12323 (N_12323,N_12053,N_12142);
nor U12324 (N_12324,N_12165,N_12173);
nand U12325 (N_12325,N_12159,N_12094);
nand U12326 (N_12326,N_12072,N_12019);
nor U12327 (N_12327,N_12183,N_12105);
or U12328 (N_12328,N_12194,N_12208);
nor U12329 (N_12329,N_12029,N_12091);
nor U12330 (N_12330,N_12231,N_12163);
nor U12331 (N_12331,N_12052,N_12123);
nand U12332 (N_12332,N_12077,N_12001);
or U12333 (N_12333,N_12063,N_12027);
or U12334 (N_12334,N_12043,N_12108);
xnor U12335 (N_12335,N_12037,N_12170);
nand U12336 (N_12336,N_12212,N_12035);
xnor U12337 (N_12337,N_12155,N_12177);
or U12338 (N_12338,N_12149,N_12129);
nand U12339 (N_12339,N_12190,N_12012);
xnor U12340 (N_12340,N_12127,N_12139);
nor U12341 (N_12341,N_12073,N_12081);
nand U12342 (N_12342,N_12203,N_12211);
xor U12343 (N_12343,N_12200,N_12109);
or U12344 (N_12344,N_12083,N_12084);
nand U12345 (N_12345,N_12239,N_12069);
nor U12346 (N_12346,N_12023,N_12186);
or U12347 (N_12347,N_12229,N_12179);
nand U12348 (N_12348,N_12232,N_12048);
nand U12349 (N_12349,N_12242,N_12075);
nor U12350 (N_12350,N_12004,N_12204);
nor U12351 (N_12351,N_12055,N_12132);
nor U12352 (N_12352,N_12008,N_12182);
nand U12353 (N_12353,N_12104,N_12024);
nand U12354 (N_12354,N_12137,N_12130);
or U12355 (N_12355,N_12158,N_12172);
or U12356 (N_12356,N_12120,N_12066);
or U12357 (N_12357,N_12148,N_12136);
and U12358 (N_12358,N_12224,N_12111);
or U12359 (N_12359,N_12056,N_12124);
and U12360 (N_12360,N_12217,N_12145);
or U12361 (N_12361,N_12157,N_12220);
or U12362 (N_12362,N_12125,N_12160);
nor U12363 (N_12363,N_12025,N_12116);
xnor U12364 (N_12364,N_12131,N_12028);
nor U12365 (N_12365,N_12034,N_12074);
xor U12366 (N_12366,N_12062,N_12249);
or U12367 (N_12367,N_12005,N_12090);
nor U12368 (N_12368,N_12219,N_12020);
and U12369 (N_12369,N_12080,N_12213);
and U12370 (N_12370,N_12227,N_12036);
xnor U12371 (N_12371,N_12222,N_12000);
nand U12372 (N_12372,N_12185,N_12076);
and U12373 (N_12373,N_12152,N_12038);
nand U12374 (N_12374,N_12191,N_12013);
nand U12375 (N_12375,N_12036,N_12136);
nand U12376 (N_12376,N_12052,N_12143);
nor U12377 (N_12377,N_12032,N_12219);
or U12378 (N_12378,N_12106,N_12175);
nand U12379 (N_12379,N_12183,N_12238);
xor U12380 (N_12380,N_12071,N_12008);
and U12381 (N_12381,N_12082,N_12191);
and U12382 (N_12382,N_12128,N_12026);
xnor U12383 (N_12383,N_12022,N_12188);
nand U12384 (N_12384,N_12242,N_12099);
xnor U12385 (N_12385,N_12025,N_12141);
and U12386 (N_12386,N_12046,N_12008);
nand U12387 (N_12387,N_12245,N_12248);
xnor U12388 (N_12388,N_12006,N_12109);
and U12389 (N_12389,N_12029,N_12024);
or U12390 (N_12390,N_12025,N_12208);
xnor U12391 (N_12391,N_12052,N_12189);
nor U12392 (N_12392,N_12203,N_12028);
nand U12393 (N_12393,N_12054,N_12168);
xnor U12394 (N_12394,N_12243,N_12215);
nand U12395 (N_12395,N_12209,N_12005);
and U12396 (N_12396,N_12200,N_12130);
xnor U12397 (N_12397,N_12169,N_12073);
or U12398 (N_12398,N_12110,N_12130);
nand U12399 (N_12399,N_12009,N_12219);
nand U12400 (N_12400,N_12037,N_12163);
and U12401 (N_12401,N_12194,N_12214);
nor U12402 (N_12402,N_12093,N_12064);
nor U12403 (N_12403,N_12244,N_12018);
nand U12404 (N_12404,N_12044,N_12000);
xnor U12405 (N_12405,N_12115,N_12087);
nor U12406 (N_12406,N_12189,N_12077);
nor U12407 (N_12407,N_12149,N_12181);
nor U12408 (N_12408,N_12039,N_12095);
xor U12409 (N_12409,N_12132,N_12020);
nand U12410 (N_12410,N_12188,N_12178);
nor U12411 (N_12411,N_12112,N_12228);
or U12412 (N_12412,N_12152,N_12068);
nor U12413 (N_12413,N_12121,N_12110);
nand U12414 (N_12414,N_12132,N_12054);
nand U12415 (N_12415,N_12248,N_12045);
xor U12416 (N_12416,N_12147,N_12027);
or U12417 (N_12417,N_12131,N_12161);
or U12418 (N_12418,N_12247,N_12028);
and U12419 (N_12419,N_12108,N_12140);
and U12420 (N_12420,N_12203,N_12163);
nor U12421 (N_12421,N_12216,N_12191);
nor U12422 (N_12422,N_12101,N_12185);
and U12423 (N_12423,N_12171,N_12227);
or U12424 (N_12424,N_12110,N_12098);
nor U12425 (N_12425,N_12137,N_12139);
nand U12426 (N_12426,N_12249,N_12212);
and U12427 (N_12427,N_12214,N_12112);
and U12428 (N_12428,N_12039,N_12117);
nor U12429 (N_12429,N_12126,N_12066);
and U12430 (N_12430,N_12079,N_12075);
xnor U12431 (N_12431,N_12161,N_12035);
nor U12432 (N_12432,N_12119,N_12074);
xnor U12433 (N_12433,N_12104,N_12218);
nand U12434 (N_12434,N_12071,N_12042);
xor U12435 (N_12435,N_12245,N_12156);
nor U12436 (N_12436,N_12033,N_12214);
and U12437 (N_12437,N_12210,N_12235);
or U12438 (N_12438,N_12109,N_12185);
or U12439 (N_12439,N_12155,N_12026);
and U12440 (N_12440,N_12178,N_12161);
xor U12441 (N_12441,N_12216,N_12134);
nor U12442 (N_12442,N_12022,N_12068);
xor U12443 (N_12443,N_12096,N_12243);
nand U12444 (N_12444,N_12059,N_12229);
and U12445 (N_12445,N_12037,N_12116);
or U12446 (N_12446,N_12210,N_12181);
and U12447 (N_12447,N_12189,N_12106);
xnor U12448 (N_12448,N_12073,N_12083);
nand U12449 (N_12449,N_12080,N_12041);
nor U12450 (N_12450,N_12146,N_12030);
xor U12451 (N_12451,N_12070,N_12177);
nand U12452 (N_12452,N_12082,N_12021);
or U12453 (N_12453,N_12008,N_12204);
xor U12454 (N_12454,N_12122,N_12214);
or U12455 (N_12455,N_12217,N_12223);
xor U12456 (N_12456,N_12019,N_12115);
xnor U12457 (N_12457,N_12033,N_12002);
xor U12458 (N_12458,N_12149,N_12134);
or U12459 (N_12459,N_12105,N_12209);
nor U12460 (N_12460,N_12192,N_12033);
nor U12461 (N_12461,N_12190,N_12209);
xor U12462 (N_12462,N_12003,N_12223);
xor U12463 (N_12463,N_12003,N_12095);
xor U12464 (N_12464,N_12087,N_12192);
nand U12465 (N_12465,N_12089,N_12124);
or U12466 (N_12466,N_12017,N_12114);
or U12467 (N_12467,N_12188,N_12198);
and U12468 (N_12468,N_12018,N_12126);
nand U12469 (N_12469,N_12243,N_12174);
nand U12470 (N_12470,N_12037,N_12245);
xor U12471 (N_12471,N_12129,N_12231);
or U12472 (N_12472,N_12016,N_12112);
nor U12473 (N_12473,N_12148,N_12135);
or U12474 (N_12474,N_12014,N_12062);
or U12475 (N_12475,N_12229,N_12086);
or U12476 (N_12476,N_12230,N_12198);
or U12477 (N_12477,N_12223,N_12180);
nand U12478 (N_12478,N_12099,N_12037);
and U12479 (N_12479,N_12057,N_12218);
nor U12480 (N_12480,N_12189,N_12065);
or U12481 (N_12481,N_12143,N_12077);
and U12482 (N_12482,N_12128,N_12140);
and U12483 (N_12483,N_12104,N_12229);
xor U12484 (N_12484,N_12158,N_12242);
or U12485 (N_12485,N_12188,N_12129);
and U12486 (N_12486,N_12172,N_12054);
xnor U12487 (N_12487,N_12152,N_12027);
nand U12488 (N_12488,N_12031,N_12239);
nor U12489 (N_12489,N_12235,N_12012);
xnor U12490 (N_12490,N_12075,N_12161);
xnor U12491 (N_12491,N_12160,N_12059);
nor U12492 (N_12492,N_12199,N_12128);
or U12493 (N_12493,N_12039,N_12238);
nand U12494 (N_12494,N_12037,N_12024);
nand U12495 (N_12495,N_12138,N_12168);
and U12496 (N_12496,N_12141,N_12066);
and U12497 (N_12497,N_12029,N_12230);
nor U12498 (N_12498,N_12003,N_12115);
nand U12499 (N_12499,N_12111,N_12098);
nor U12500 (N_12500,N_12298,N_12338);
or U12501 (N_12501,N_12314,N_12378);
or U12502 (N_12502,N_12252,N_12320);
and U12503 (N_12503,N_12441,N_12339);
xor U12504 (N_12504,N_12418,N_12353);
nor U12505 (N_12505,N_12313,N_12377);
nand U12506 (N_12506,N_12358,N_12348);
or U12507 (N_12507,N_12375,N_12489);
xnor U12508 (N_12508,N_12469,N_12437);
nand U12509 (N_12509,N_12372,N_12488);
and U12510 (N_12510,N_12302,N_12495);
or U12511 (N_12511,N_12317,N_12286);
xnor U12512 (N_12512,N_12267,N_12264);
nor U12513 (N_12513,N_12420,N_12394);
and U12514 (N_12514,N_12265,N_12496);
xor U12515 (N_12515,N_12455,N_12304);
and U12516 (N_12516,N_12402,N_12474);
nor U12517 (N_12517,N_12368,N_12274);
and U12518 (N_12518,N_12276,N_12475);
nor U12519 (N_12519,N_12443,N_12250);
or U12520 (N_12520,N_12391,N_12432);
or U12521 (N_12521,N_12433,N_12306);
and U12522 (N_12522,N_12283,N_12260);
and U12523 (N_12523,N_12261,N_12430);
or U12524 (N_12524,N_12476,N_12340);
xnor U12525 (N_12525,N_12292,N_12397);
and U12526 (N_12526,N_12266,N_12341);
xor U12527 (N_12527,N_12407,N_12381);
nor U12528 (N_12528,N_12279,N_12386);
and U12529 (N_12529,N_12392,N_12434);
nor U12530 (N_12530,N_12413,N_12263);
xor U12531 (N_12531,N_12308,N_12492);
xor U12532 (N_12532,N_12349,N_12466);
xor U12533 (N_12533,N_12429,N_12427);
xor U12534 (N_12534,N_12484,N_12417);
xnor U12535 (N_12535,N_12270,N_12440);
xor U12536 (N_12536,N_12327,N_12334);
or U12537 (N_12537,N_12384,N_12342);
nand U12538 (N_12538,N_12347,N_12382);
nand U12539 (N_12539,N_12410,N_12345);
nand U12540 (N_12540,N_12256,N_12460);
and U12541 (N_12541,N_12419,N_12486);
nor U12542 (N_12542,N_12373,N_12477);
xor U12543 (N_12543,N_12388,N_12409);
nor U12544 (N_12544,N_12360,N_12387);
nor U12545 (N_12545,N_12284,N_12403);
or U12546 (N_12546,N_12465,N_12493);
xor U12547 (N_12547,N_12452,N_12406);
xor U12548 (N_12548,N_12271,N_12350);
nand U12549 (N_12549,N_12344,N_12312);
nand U12550 (N_12550,N_12472,N_12445);
xnor U12551 (N_12551,N_12294,N_12385);
and U12552 (N_12552,N_12396,N_12404);
and U12553 (N_12553,N_12325,N_12468);
nor U12554 (N_12554,N_12322,N_12405);
xnor U12555 (N_12555,N_12389,N_12285);
nand U12556 (N_12556,N_12311,N_12422);
and U12557 (N_12557,N_12331,N_12473);
and U12558 (N_12558,N_12303,N_12498);
or U12559 (N_12559,N_12451,N_12467);
nor U12560 (N_12560,N_12416,N_12426);
nand U12561 (N_12561,N_12436,N_12251);
xnor U12562 (N_12562,N_12280,N_12254);
nor U12563 (N_12563,N_12258,N_12272);
nor U12564 (N_12564,N_12369,N_12257);
nor U12565 (N_12565,N_12371,N_12295);
nor U12566 (N_12566,N_12262,N_12357);
or U12567 (N_12567,N_12332,N_12379);
and U12568 (N_12568,N_12435,N_12365);
nand U12569 (N_12569,N_12310,N_12329);
and U12570 (N_12570,N_12290,N_12447);
nor U12571 (N_12571,N_12352,N_12330);
nor U12572 (N_12572,N_12362,N_12268);
or U12573 (N_12573,N_12335,N_12363);
nand U12574 (N_12574,N_12454,N_12305);
and U12575 (N_12575,N_12390,N_12269);
xor U12576 (N_12576,N_12494,N_12464);
and U12577 (N_12577,N_12478,N_12483);
and U12578 (N_12578,N_12355,N_12364);
xnor U12579 (N_12579,N_12398,N_12356);
xnor U12580 (N_12580,N_12450,N_12366);
xor U12581 (N_12581,N_12444,N_12343);
nor U12582 (N_12582,N_12380,N_12289);
or U12583 (N_12583,N_12453,N_12287);
xor U12584 (N_12584,N_12456,N_12288);
xor U12585 (N_12585,N_12299,N_12490);
xnor U12586 (N_12586,N_12480,N_12315);
xor U12587 (N_12587,N_12414,N_12463);
and U12588 (N_12588,N_12497,N_12401);
xor U12589 (N_12589,N_12282,N_12400);
xnor U12590 (N_12590,N_12481,N_12333);
nand U12591 (N_12591,N_12411,N_12318);
and U12592 (N_12592,N_12415,N_12412);
xor U12593 (N_12593,N_12301,N_12383);
and U12594 (N_12594,N_12424,N_12278);
nor U12595 (N_12595,N_12438,N_12462);
or U12596 (N_12596,N_12485,N_12277);
nand U12597 (N_12597,N_12336,N_12324);
xnor U12598 (N_12598,N_12367,N_12421);
or U12599 (N_12599,N_12351,N_12309);
xor U12600 (N_12600,N_12255,N_12448);
nor U12601 (N_12601,N_12359,N_12296);
xor U12602 (N_12602,N_12374,N_12487);
nand U12603 (N_12603,N_12376,N_12273);
nand U12604 (N_12604,N_12459,N_12281);
nand U12605 (N_12605,N_12337,N_12439);
and U12606 (N_12606,N_12479,N_12297);
xnor U12607 (N_12607,N_12471,N_12354);
xor U12608 (N_12608,N_12321,N_12482);
nand U12609 (N_12609,N_12361,N_12291);
nor U12610 (N_12610,N_12449,N_12461);
nor U12611 (N_12611,N_12499,N_12457);
or U12612 (N_12612,N_12326,N_12319);
nor U12613 (N_12613,N_12370,N_12408);
nand U12614 (N_12614,N_12346,N_12253);
or U12615 (N_12615,N_12399,N_12470);
and U12616 (N_12616,N_12428,N_12458);
nor U12617 (N_12617,N_12446,N_12431);
xnor U12618 (N_12618,N_12393,N_12423);
nand U12619 (N_12619,N_12275,N_12316);
and U12620 (N_12620,N_12300,N_12425);
or U12621 (N_12621,N_12307,N_12328);
nand U12622 (N_12622,N_12395,N_12491);
nor U12623 (N_12623,N_12442,N_12259);
or U12624 (N_12624,N_12293,N_12323);
nor U12625 (N_12625,N_12356,N_12387);
and U12626 (N_12626,N_12353,N_12409);
xnor U12627 (N_12627,N_12426,N_12258);
and U12628 (N_12628,N_12456,N_12330);
and U12629 (N_12629,N_12399,N_12395);
nor U12630 (N_12630,N_12390,N_12253);
xor U12631 (N_12631,N_12265,N_12405);
xnor U12632 (N_12632,N_12315,N_12489);
and U12633 (N_12633,N_12264,N_12497);
nand U12634 (N_12634,N_12297,N_12456);
xnor U12635 (N_12635,N_12254,N_12346);
and U12636 (N_12636,N_12335,N_12384);
nor U12637 (N_12637,N_12373,N_12427);
nor U12638 (N_12638,N_12294,N_12252);
or U12639 (N_12639,N_12329,N_12313);
nor U12640 (N_12640,N_12268,N_12337);
and U12641 (N_12641,N_12261,N_12398);
nand U12642 (N_12642,N_12436,N_12268);
or U12643 (N_12643,N_12431,N_12327);
xor U12644 (N_12644,N_12470,N_12306);
and U12645 (N_12645,N_12340,N_12322);
or U12646 (N_12646,N_12381,N_12460);
and U12647 (N_12647,N_12453,N_12302);
or U12648 (N_12648,N_12498,N_12398);
xor U12649 (N_12649,N_12436,N_12468);
or U12650 (N_12650,N_12358,N_12355);
and U12651 (N_12651,N_12288,N_12338);
and U12652 (N_12652,N_12404,N_12325);
and U12653 (N_12653,N_12303,N_12412);
nor U12654 (N_12654,N_12388,N_12372);
nor U12655 (N_12655,N_12261,N_12388);
nand U12656 (N_12656,N_12370,N_12263);
and U12657 (N_12657,N_12446,N_12365);
nor U12658 (N_12658,N_12326,N_12359);
and U12659 (N_12659,N_12383,N_12325);
nand U12660 (N_12660,N_12492,N_12345);
xnor U12661 (N_12661,N_12282,N_12364);
or U12662 (N_12662,N_12481,N_12254);
nor U12663 (N_12663,N_12333,N_12297);
xor U12664 (N_12664,N_12395,N_12446);
and U12665 (N_12665,N_12255,N_12440);
or U12666 (N_12666,N_12289,N_12406);
xnor U12667 (N_12667,N_12324,N_12385);
nand U12668 (N_12668,N_12463,N_12449);
nor U12669 (N_12669,N_12259,N_12293);
and U12670 (N_12670,N_12328,N_12463);
or U12671 (N_12671,N_12441,N_12451);
nor U12672 (N_12672,N_12311,N_12464);
nor U12673 (N_12673,N_12287,N_12493);
or U12674 (N_12674,N_12480,N_12347);
xor U12675 (N_12675,N_12385,N_12361);
xnor U12676 (N_12676,N_12265,N_12447);
and U12677 (N_12677,N_12372,N_12251);
or U12678 (N_12678,N_12279,N_12295);
and U12679 (N_12679,N_12465,N_12384);
or U12680 (N_12680,N_12443,N_12436);
xnor U12681 (N_12681,N_12285,N_12310);
or U12682 (N_12682,N_12386,N_12410);
nor U12683 (N_12683,N_12472,N_12385);
or U12684 (N_12684,N_12390,N_12403);
or U12685 (N_12685,N_12251,N_12407);
nand U12686 (N_12686,N_12432,N_12264);
xnor U12687 (N_12687,N_12426,N_12298);
and U12688 (N_12688,N_12342,N_12433);
nand U12689 (N_12689,N_12298,N_12439);
or U12690 (N_12690,N_12429,N_12323);
nand U12691 (N_12691,N_12390,N_12497);
xnor U12692 (N_12692,N_12252,N_12434);
and U12693 (N_12693,N_12253,N_12321);
or U12694 (N_12694,N_12487,N_12492);
nand U12695 (N_12695,N_12261,N_12312);
nand U12696 (N_12696,N_12381,N_12399);
or U12697 (N_12697,N_12325,N_12375);
and U12698 (N_12698,N_12449,N_12345);
or U12699 (N_12699,N_12404,N_12312);
nand U12700 (N_12700,N_12287,N_12411);
nand U12701 (N_12701,N_12271,N_12365);
or U12702 (N_12702,N_12499,N_12343);
and U12703 (N_12703,N_12283,N_12411);
nand U12704 (N_12704,N_12304,N_12383);
or U12705 (N_12705,N_12452,N_12320);
nand U12706 (N_12706,N_12337,N_12444);
nor U12707 (N_12707,N_12371,N_12367);
xnor U12708 (N_12708,N_12304,N_12473);
xnor U12709 (N_12709,N_12349,N_12455);
nand U12710 (N_12710,N_12375,N_12320);
or U12711 (N_12711,N_12401,N_12289);
xor U12712 (N_12712,N_12419,N_12494);
nand U12713 (N_12713,N_12305,N_12269);
xor U12714 (N_12714,N_12329,N_12486);
and U12715 (N_12715,N_12307,N_12256);
and U12716 (N_12716,N_12274,N_12340);
nand U12717 (N_12717,N_12485,N_12315);
nor U12718 (N_12718,N_12340,N_12310);
nand U12719 (N_12719,N_12252,N_12412);
nand U12720 (N_12720,N_12447,N_12435);
xnor U12721 (N_12721,N_12276,N_12459);
or U12722 (N_12722,N_12484,N_12286);
nand U12723 (N_12723,N_12251,N_12275);
xor U12724 (N_12724,N_12456,N_12347);
and U12725 (N_12725,N_12309,N_12392);
or U12726 (N_12726,N_12388,N_12481);
nand U12727 (N_12727,N_12290,N_12273);
xnor U12728 (N_12728,N_12348,N_12408);
or U12729 (N_12729,N_12317,N_12436);
xnor U12730 (N_12730,N_12287,N_12459);
xor U12731 (N_12731,N_12404,N_12280);
xor U12732 (N_12732,N_12474,N_12442);
xor U12733 (N_12733,N_12283,N_12439);
or U12734 (N_12734,N_12432,N_12464);
and U12735 (N_12735,N_12427,N_12355);
or U12736 (N_12736,N_12431,N_12426);
xnor U12737 (N_12737,N_12442,N_12306);
and U12738 (N_12738,N_12389,N_12371);
nor U12739 (N_12739,N_12342,N_12318);
and U12740 (N_12740,N_12407,N_12258);
or U12741 (N_12741,N_12301,N_12429);
or U12742 (N_12742,N_12257,N_12407);
and U12743 (N_12743,N_12470,N_12308);
nand U12744 (N_12744,N_12299,N_12418);
and U12745 (N_12745,N_12441,N_12299);
or U12746 (N_12746,N_12388,N_12440);
nor U12747 (N_12747,N_12268,N_12423);
nand U12748 (N_12748,N_12340,N_12430);
xor U12749 (N_12749,N_12396,N_12478);
or U12750 (N_12750,N_12655,N_12662);
or U12751 (N_12751,N_12510,N_12543);
xor U12752 (N_12752,N_12702,N_12545);
nor U12753 (N_12753,N_12676,N_12649);
nand U12754 (N_12754,N_12696,N_12719);
nor U12755 (N_12755,N_12692,N_12657);
and U12756 (N_12756,N_12598,N_12516);
xor U12757 (N_12757,N_12555,N_12581);
or U12758 (N_12758,N_12551,N_12612);
nor U12759 (N_12759,N_12747,N_12671);
or U12760 (N_12760,N_12541,N_12678);
or U12761 (N_12761,N_12506,N_12568);
nor U12762 (N_12762,N_12668,N_12695);
and U12763 (N_12763,N_12567,N_12505);
or U12764 (N_12764,N_12539,N_12528);
nand U12765 (N_12765,N_12698,N_12615);
nand U12766 (N_12766,N_12582,N_12617);
nor U12767 (N_12767,N_12621,N_12652);
or U12768 (N_12768,N_12590,N_12643);
nor U12769 (N_12769,N_12500,N_12630);
or U12770 (N_12770,N_12550,N_12704);
or U12771 (N_12771,N_12736,N_12563);
nor U12772 (N_12772,N_12647,N_12554);
or U12773 (N_12773,N_12586,N_12663);
xnor U12774 (N_12774,N_12527,N_12712);
nor U12775 (N_12775,N_12574,N_12690);
or U12776 (N_12776,N_12691,N_12659);
xor U12777 (N_12777,N_12656,N_12660);
xor U12778 (N_12778,N_12522,N_12687);
nand U12779 (N_12779,N_12749,N_12608);
nand U12780 (N_12780,N_12675,N_12537);
xor U12781 (N_12781,N_12644,N_12531);
xor U12782 (N_12782,N_12714,N_12625);
or U12783 (N_12783,N_12746,N_12706);
xnor U12784 (N_12784,N_12629,N_12593);
and U12785 (N_12785,N_12523,N_12705);
or U12786 (N_12786,N_12648,N_12573);
and U12787 (N_12787,N_12616,N_12507);
nor U12788 (N_12788,N_12564,N_12583);
xnor U12789 (N_12789,N_12632,N_12618);
nand U12790 (N_12790,N_12666,N_12673);
or U12791 (N_12791,N_12589,N_12658);
nor U12792 (N_12792,N_12599,N_12699);
and U12793 (N_12793,N_12602,N_12742);
nor U12794 (N_12794,N_12743,N_12511);
and U12795 (N_12795,N_12639,N_12501);
or U12796 (N_12796,N_12641,N_12595);
and U12797 (N_12797,N_12606,N_12619);
nand U12798 (N_12798,N_12703,N_12721);
and U12799 (N_12799,N_12620,N_12680);
nand U12800 (N_12800,N_12728,N_12627);
xor U12801 (N_12801,N_12709,N_12536);
or U12802 (N_12802,N_12524,N_12674);
nor U12803 (N_12803,N_12587,N_12701);
or U12804 (N_12804,N_12634,N_12513);
and U12805 (N_12805,N_12733,N_12650);
and U12806 (N_12806,N_12519,N_12729);
nor U12807 (N_12807,N_12614,N_12596);
and U12808 (N_12808,N_12628,N_12626);
and U12809 (N_12809,N_12745,N_12578);
or U12810 (N_12810,N_12585,N_12645);
nor U12811 (N_12811,N_12600,N_12518);
nor U12812 (N_12812,N_12651,N_12509);
xor U12813 (N_12813,N_12653,N_12694);
and U12814 (N_12814,N_12569,N_12515);
xor U12815 (N_12815,N_12514,N_12670);
and U12816 (N_12816,N_12664,N_12560);
nand U12817 (N_12817,N_12533,N_12716);
nor U12818 (N_12818,N_12558,N_12732);
and U12819 (N_12819,N_12594,N_12734);
nand U12820 (N_12820,N_12685,N_12744);
nand U12821 (N_12821,N_12526,N_12566);
or U12822 (N_12822,N_12542,N_12723);
nand U12823 (N_12823,N_12635,N_12597);
or U12824 (N_12824,N_12683,N_12686);
nor U12825 (N_12825,N_12584,N_12570);
or U12826 (N_12826,N_12559,N_12603);
and U12827 (N_12827,N_12684,N_12613);
nor U12828 (N_12828,N_12740,N_12609);
nor U12829 (N_12829,N_12741,N_12640);
or U12830 (N_12830,N_12737,N_12708);
nor U12831 (N_12831,N_12535,N_12504);
nand U12832 (N_12832,N_12715,N_12730);
nor U12833 (N_12833,N_12718,N_12553);
or U12834 (N_12834,N_12646,N_12622);
nor U12835 (N_12835,N_12738,N_12546);
and U12836 (N_12836,N_12688,N_12682);
or U12837 (N_12837,N_12624,N_12735);
nor U12838 (N_12838,N_12611,N_12576);
or U12839 (N_12839,N_12552,N_12547);
and U12840 (N_12840,N_12538,N_12530);
or U12841 (N_12841,N_12579,N_12575);
nand U12842 (N_12842,N_12739,N_12572);
or U12843 (N_12843,N_12588,N_12642);
or U12844 (N_12844,N_12548,N_12711);
xnor U12845 (N_12845,N_12577,N_12592);
and U12846 (N_12846,N_12610,N_12679);
nor U12847 (N_12847,N_12565,N_12726);
nand U12848 (N_12848,N_12534,N_12669);
nand U12849 (N_12849,N_12713,N_12748);
or U12850 (N_12850,N_12532,N_12604);
nor U12851 (N_12851,N_12722,N_12521);
nor U12852 (N_12852,N_12707,N_12724);
xnor U12853 (N_12853,N_12529,N_12623);
xnor U12854 (N_12854,N_12720,N_12731);
or U12855 (N_12855,N_12561,N_12502);
and U12856 (N_12856,N_12693,N_12672);
nor U12857 (N_12857,N_12727,N_12689);
nand U12858 (N_12858,N_12636,N_12525);
and U12859 (N_12859,N_12633,N_12665);
or U12860 (N_12860,N_12571,N_12717);
or U12861 (N_12861,N_12677,N_12503);
or U12862 (N_12862,N_12631,N_12605);
xnor U12863 (N_12863,N_12607,N_12540);
and U12864 (N_12864,N_12697,N_12508);
or U12865 (N_12865,N_12700,N_12638);
and U12866 (N_12866,N_12556,N_12512);
xnor U12867 (N_12867,N_12520,N_12557);
and U12868 (N_12868,N_12591,N_12549);
xor U12869 (N_12869,N_12580,N_12637);
xor U12870 (N_12870,N_12654,N_12517);
nand U12871 (N_12871,N_12544,N_12601);
nor U12872 (N_12872,N_12681,N_12725);
xnor U12873 (N_12873,N_12661,N_12562);
or U12874 (N_12874,N_12710,N_12667);
or U12875 (N_12875,N_12595,N_12645);
nand U12876 (N_12876,N_12747,N_12706);
and U12877 (N_12877,N_12624,N_12666);
xor U12878 (N_12878,N_12639,N_12633);
xor U12879 (N_12879,N_12533,N_12539);
nor U12880 (N_12880,N_12704,N_12685);
nand U12881 (N_12881,N_12711,N_12648);
and U12882 (N_12882,N_12579,N_12631);
or U12883 (N_12883,N_12541,N_12521);
or U12884 (N_12884,N_12748,N_12508);
xnor U12885 (N_12885,N_12720,N_12506);
nor U12886 (N_12886,N_12560,N_12638);
or U12887 (N_12887,N_12581,N_12515);
nand U12888 (N_12888,N_12733,N_12511);
or U12889 (N_12889,N_12504,N_12648);
and U12890 (N_12890,N_12502,N_12544);
xnor U12891 (N_12891,N_12656,N_12695);
nor U12892 (N_12892,N_12600,N_12554);
nor U12893 (N_12893,N_12684,N_12735);
or U12894 (N_12894,N_12637,N_12620);
or U12895 (N_12895,N_12658,N_12601);
nand U12896 (N_12896,N_12653,N_12608);
xnor U12897 (N_12897,N_12721,N_12687);
nor U12898 (N_12898,N_12644,N_12706);
or U12899 (N_12899,N_12719,N_12677);
or U12900 (N_12900,N_12643,N_12545);
and U12901 (N_12901,N_12621,N_12679);
nand U12902 (N_12902,N_12666,N_12519);
xnor U12903 (N_12903,N_12735,N_12714);
or U12904 (N_12904,N_12560,N_12556);
nor U12905 (N_12905,N_12674,N_12621);
nor U12906 (N_12906,N_12541,N_12745);
nand U12907 (N_12907,N_12682,N_12518);
or U12908 (N_12908,N_12531,N_12715);
xnor U12909 (N_12909,N_12705,N_12550);
nor U12910 (N_12910,N_12584,N_12691);
and U12911 (N_12911,N_12656,N_12591);
nor U12912 (N_12912,N_12682,N_12577);
or U12913 (N_12913,N_12741,N_12519);
nand U12914 (N_12914,N_12550,N_12715);
and U12915 (N_12915,N_12504,N_12594);
nand U12916 (N_12916,N_12736,N_12671);
and U12917 (N_12917,N_12700,N_12530);
and U12918 (N_12918,N_12701,N_12577);
or U12919 (N_12919,N_12694,N_12605);
or U12920 (N_12920,N_12599,N_12514);
nor U12921 (N_12921,N_12568,N_12521);
or U12922 (N_12922,N_12592,N_12693);
xor U12923 (N_12923,N_12699,N_12595);
and U12924 (N_12924,N_12529,N_12713);
or U12925 (N_12925,N_12747,N_12627);
nand U12926 (N_12926,N_12533,N_12634);
nor U12927 (N_12927,N_12593,N_12650);
nor U12928 (N_12928,N_12520,N_12570);
nand U12929 (N_12929,N_12639,N_12590);
or U12930 (N_12930,N_12701,N_12676);
and U12931 (N_12931,N_12631,N_12730);
xor U12932 (N_12932,N_12657,N_12554);
xor U12933 (N_12933,N_12669,N_12686);
nor U12934 (N_12934,N_12577,N_12618);
or U12935 (N_12935,N_12626,N_12545);
and U12936 (N_12936,N_12517,N_12532);
nor U12937 (N_12937,N_12625,N_12705);
nand U12938 (N_12938,N_12540,N_12531);
and U12939 (N_12939,N_12540,N_12720);
nand U12940 (N_12940,N_12549,N_12536);
and U12941 (N_12941,N_12540,N_12624);
or U12942 (N_12942,N_12691,N_12605);
xnor U12943 (N_12943,N_12730,N_12533);
or U12944 (N_12944,N_12710,N_12614);
xnor U12945 (N_12945,N_12681,N_12519);
or U12946 (N_12946,N_12729,N_12675);
or U12947 (N_12947,N_12691,N_12744);
xnor U12948 (N_12948,N_12696,N_12525);
and U12949 (N_12949,N_12603,N_12513);
or U12950 (N_12950,N_12670,N_12572);
nor U12951 (N_12951,N_12578,N_12658);
xnor U12952 (N_12952,N_12565,N_12611);
nand U12953 (N_12953,N_12585,N_12682);
nor U12954 (N_12954,N_12501,N_12565);
nor U12955 (N_12955,N_12673,N_12582);
nand U12956 (N_12956,N_12646,N_12679);
xor U12957 (N_12957,N_12639,N_12661);
nor U12958 (N_12958,N_12618,N_12731);
nand U12959 (N_12959,N_12590,N_12522);
nand U12960 (N_12960,N_12578,N_12500);
or U12961 (N_12961,N_12584,N_12695);
nor U12962 (N_12962,N_12509,N_12547);
and U12963 (N_12963,N_12500,N_12656);
xor U12964 (N_12964,N_12747,N_12594);
nand U12965 (N_12965,N_12578,N_12743);
nand U12966 (N_12966,N_12506,N_12576);
nand U12967 (N_12967,N_12716,N_12745);
and U12968 (N_12968,N_12587,N_12670);
and U12969 (N_12969,N_12507,N_12543);
nor U12970 (N_12970,N_12538,N_12591);
and U12971 (N_12971,N_12564,N_12545);
and U12972 (N_12972,N_12520,N_12738);
and U12973 (N_12973,N_12504,N_12627);
nand U12974 (N_12974,N_12556,N_12565);
or U12975 (N_12975,N_12652,N_12678);
nand U12976 (N_12976,N_12603,N_12608);
and U12977 (N_12977,N_12637,N_12578);
xor U12978 (N_12978,N_12676,N_12516);
and U12979 (N_12979,N_12683,N_12541);
or U12980 (N_12980,N_12617,N_12741);
and U12981 (N_12981,N_12652,N_12646);
nand U12982 (N_12982,N_12567,N_12690);
nand U12983 (N_12983,N_12692,N_12738);
xor U12984 (N_12984,N_12738,N_12515);
nand U12985 (N_12985,N_12578,N_12687);
nor U12986 (N_12986,N_12591,N_12673);
xor U12987 (N_12987,N_12665,N_12613);
or U12988 (N_12988,N_12585,N_12699);
xor U12989 (N_12989,N_12730,N_12651);
nand U12990 (N_12990,N_12542,N_12652);
nor U12991 (N_12991,N_12551,N_12650);
xor U12992 (N_12992,N_12580,N_12743);
nand U12993 (N_12993,N_12571,N_12558);
nand U12994 (N_12994,N_12637,N_12563);
xor U12995 (N_12995,N_12512,N_12693);
and U12996 (N_12996,N_12613,N_12601);
and U12997 (N_12997,N_12558,N_12722);
xor U12998 (N_12998,N_12542,N_12709);
and U12999 (N_12999,N_12520,N_12536);
and U13000 (N_13000,N_12958,N_12951);
and U13001 (N_13001,N_12850,N_12766);
nor U13002 (N_13002,N_12874,N_12841);
nand U13003 (N_13003,N_12948,N_12889);
xnor U13004 (N_13004,N_12903,N_12811);
xor U13005 (N_13005,N_12756,N_12885);
nor U13006 (N_13006,N_12990,N_12788);
nor U13007 (N_13007,N_12828,N_12761);
nand U13008 (N_13008,N_12805,N_12823);
nor U13009 (N_13009,N_12926,N_12853);
or U13010 (N_13010,N_12978,N_12825);
and U13011 (N_13011,N_12770,N_12804);
or U13012 (N_13012,N_12963,N_12773);
and U13013 (N_13013,N_12778,N_12839);
nor U13014 (N_13014,N_12918,N_12912);
nand U13015 (N_13015,N_12763,N_12999);
nor U13016 (N_13016,N_12939,N_12813);
or U13017 (N_13017,N_12835,N_12758);
nand U13018 (N_13018,N_12959,N_12900);
nor U13019 (N_13019,N_12847,N_12754);
nor U13020 (N_13020,N_12865,N_12934);
and U13021 (N_13021,N_12777,N_12976);
xor U13022 (N_13022,N_12946,N_12924);
and U13023 (N_13023,N_12809,N_12907);
xor U13024 (N_13024,N_12843,N_12919);
nor U13025 (N_13025,N_12960,N_12981);
nand U13026 (N_13026,N_12833,N_12972);
xor U13027 (N_13027,N_12859,N_12973);
or U13028 (N_13028,N_12937,N_12969);
or U13029 (N_13029,N_12769,N_12970);
nand U13030 (N_13030,N_12916,N_12817);
nor U13031 (N_13031,N_12944,N_12938);
xnor U13032 (N_13032,N_12895,N_12849);
or U13033 (N_13033,N_12751,N_12979);
nand U13034 (N_13034,N_12952,N_12868);
and U13035 (N_13035,N_12857,N_12755);
xor U13036 (N_13036,N_12925,N_12995);
nor U13037 (N_13037,N_12820,N_12826);
and U13038 (N_13038,N_12871,N_12984);
and U13039 (N_13039,N_12795,N_12863);
xnor U13040 (N_13040,N_12797,N_12877);
xor U13041 (N_13041,N_12838,N_12818);
nor U13042 (N_13042,N_12909,N_12914);
and U13043 (N_13043,N_12760,N_12893);
nand U13044 (N_13044,N_12856,N_12852);
nor U13045 (N_13045,N_12832,N_12915);
and U13046 (N_13046,N_12931,N_12971);
nor U13047 (N_13047,N_12815,N_12928);
nand U13048 (N_13048,N_12792,N_12870);
nand U13049 (N_13049,N_12997,N_12869);
nor U13050 (N_13050,N_12993,N_12779);
xor U13051 (N_13051,N_12930,N_12822);
xnor U13052 (N_13052,N_12898,N_12796);
xnor U13053 (N_13053,N_12789,N_12932);
nand U13054 (N_13054,N_12955,N_12967);
and U13055 (N_13055,N_12784,N_12782);
and U13056 (N_13056,N_12872,N_12992);
xor U13057 (N_13057,N_12883,N_12791);
and U13058 (N_13058,N_12980,N_12917);
or U13059 (N_13059,N_12882,N_12757);
nor U13060 (N_13060,N_12837,N_12892);
xnor U13061 (N_13061,N_12807,N_12989);
nand U13062 (N_13062,N_12798,N_12765);
nand U13063 (N_13063,N_12860,N_12904);
or U13064 (N_13064,N_12962,N_12940);
and U13065 (N_13065,N_12975,N_12986);
or U13066 (N_13066,N_12793,N_12861);
nor U13067 (N_13067,N_12768,N_12921);
nand U13068 (N_13068,N_12836,N_12824);
nand U13069 (N_13069,N_12816,N_12879);
nor U13070 (N_13070,N_12949,N_12886);
and U13071 (N_13071,N_12941,N_12950);
xnor U13072 (N_13072,N_12845,N_12913);
and U13073 (N_13073,N_12964,N_12956);
nor U13074 (N_13074,N_12772,N_12876);
nand U13075 (N_13075,N_12831,N_12827);
nor U13076 (N_13076,N_12810,N_12750);
or U13077 (N_13077,N_12819,N_12942);
nor U13078 (N_13078,N_12787,N_12968);
or U13079 (N_13079,N_12808,N_12897);
nor U13080 (N_13080,N_12806,N_12759);
xnor U13081 (N_13081,N_12906,N_12775);
xnor U13082 (N_13082,N_12801,N_12994);
nand U13083 (N_13083,N_12890,N_12764);
nor U13084 (N_13084,N_12776,N_12901);
xor U13085 (N_13085,N_12899,N_12966);
nand U13086 (N_13086,N_12753,N_12974);
or U13087 (N_13087,N_12996,N_12927);
and U13088 (N_13088,N_12774,N_12982);
or U13089 (N_13089,N_12799,N_12781);
and U13090 (N_13090,N_12991,N_12884);
xnor U13091 (N_13091,N_12923,N_12985);
nor U13092 (N_13092,N_12834,N_12780);
xor U13093 (N_13093,N_12953,N_12790);
and U13094 (N_13094,N_12922,N_12908);
or U13095 (N_13095,N_12965,N_12910);
and U13096 (N_13096,N_12851,N_12848);
or U13097 (N_13097,N_12830,N_12911);
nand U13098 (N_13098,N_12802,N_12875);
and U13099 (N_13099,N_12794,N_12786);
and U13100 (N_13100,N_12998,N_12881);
xor U13101 (N_13101,N_12896,N_12803);
xor U13102 (N_13102,N_12945,N_12864);
xnor U13103 (N_13103,N_12935,N_12862);
or U13104 (N_13104,N_12977,N_12812);
or U13105 (N_13105,N_12854,N_12767);
or U13106 (N_13106,N_12800,N_12752);
nand U13107 (N_13107,N_12762,N_12888);
nand U13108 (N_13108,N_12947,N_12821);
and U13109 (N_13109,N_12936,N_12842);
and U13110 (N_13110,N_12866,N_12983);
and U13111 (N_13111,N_12846,N_12905);
and U13112 (N_13112,N_12840,N_12858);
nand U13113 (N_13113,N_12880,N_12987);
xnor U13114 (N_13114,N_12814,N_12988);
or U13115 (N_13115,N_12873,N_12961);
or U13116 (N_13116,N_12867,N_12957);
xnor U13117 (N_13117,N_12783,N_12771);
nand U13118 (N_13118,N_12829,N_12920);
nand U13119 (N_13119,N_12894,N_12855);
nor U13120 (N_13120,N_12902,N_12954);
nand U13121 (N_13121,N_12891,N_12929);
xnor U13122 (N_13122,N_12878,N_12785);
xor U13123 (N_13123,N_12844,N_12887);
xor U13124 (N_13124,N_12933,N_12943);
xor U13125 (N_13125,N_12795,N_12948);
nand U13126 (N_13126,N_12904,N_12990);
and U13127 (N_13127,N_12939,N_12876);
nand U13128 (N_13128,N_12885,N_12882);
xnor U13129 (N_13129,N_12827,N_12838);
and U13130 (N_13130,N_12824,N_12785);
or U13131 (N_13131,N_12794,N_12972);
xnor U13132 (N_13132,N_12991,N_12815);
and U13133 (N_13133,N_12935,N_12791);
or U13134 (N_13134,N_12795,N_12786);
and U13135 (N_13135,N_12843,N_12887);
nand U13136 (N_13136,N_12858,N_12836);
nor U13137 (N_13137,N_12933,N_12889);
or U13138 (N_13138,N_12979,N_12886);
nand U13139 (N_13139,N_12764,N_12935);
or U13140 (N_13140,N_12847,N_12750);
nand U13141 (N_13141,N_12810,N_12968);
xor U13142 (N_13142,N_12985,N_12995);
or U13143 (N_13143,N_12909,N_12821);
nand U13144 (N_13144,N_12992,N_12842);
or U13145 (N_13145,N_12996,N_12798);
nor U13146 (N_13146,N_12846,N_12763);
and U13147 (N_13147,N_12849,N_12949);
nor U13148 (N_13148,N_12779,N_12891);
or U13149 (N_13149,N_12780,N_12837);
xor U13150 (N_13150,N_12820,N_12750);
or U13151 (N_13151,N_12795,N_12865);
and U13152 (N_13152,N_12775,N_12984);
nor U13153 (N_13153,N_12962,N_12751);
nand U13154 (N_13154,N_12885,N_12896);
xnor U13155 (N_13155,N_12929,N_12775);
xnor U13156 (N_13156,N_12986,N_12951);
and U13157 (N_13157,N_12966,N_12874);
nor U13158 (N_13158,N_12876,N_12964);
or U13159 (N_13159,N_12813,N_12830);
nand U13160 (N_13160,N_12787,N_12946);
nand U13161 (N_13161,N_12976,N_12963);
nor U13162 (N_13162,N_12874,N_12855);
or U13163 (N_13163,N_12956,N_12843);
or U13164 (N_13164,N_12913,N_12802);
xor U13165 (N_13165,N_12940,N_12775);
and U13166 (N_13166,N_12767,N_12915);
xor U13167 (N_13167,N_12792,N_12875);
nand U13168 (N_13168,N_12929,N_12909);
xnor U13169 (N_13169,N_12840,N_12913);
nand U13170 (N_13170,N_12929,N_12941);
nand U13171 (N_13171,N_12814,N_12826);
or U13172 (N_13172,N_12777,N_12832);
nor U13173 (N_13173,N_12766,N_12784);
xnor U13174 (N_13174,N_12771,N_12939);
and U13175 (N_13175,N_12837,N_12973);
and U13176 (N_13176,N_12945,N_12752);
or U13177 (N_13177,N_12881,N_12878);
and U13178 (N_13178,N_12865,N_12764);
or U13179 (N_13179,N_12820,N_12901);
nand U13180 (N_13180,N_12859,N_12857);
nand U13181 (N_13181,N_12895,N_12792);
xnor U13182 (N_13182,N_12903,N_12978);
or U13183 (N_13183,N_12792,N_12979);
nand U13184 (N_13184,N_12865,N_12778);
and U13185 (N_13185,N_12917,N_12911);
nor U13186 (N_13186,N_12750,N_12770);
xnor U13187 (N_13187,N_12902,N_12765);
or U13188 (N_13188,N_12822,N_12893);
and U13189 (N_13189,N_12778,N_12883);
or U13190 (N_13190,N_12750,N_12756);
nor U13191 (N_13191,N_12904,N_12972);
or U13192 (N_13192,N_12902,N_12933);
xor U13193 (N_13193,N_12786,N_12972);
nor U13194 (N_13194,N_12942,N_12846);
nand U13195 (N_13195,N_12752,N_12868);
xnor U13196 (N_13196,N_12888,N_12785);
nor U13197 (N_13197,N_12918,N_12791);
or U13198 (N_13198,N_12879,N_12990);
and U13199 (N_13199,N_12835,N_12999);
nand U13200 (N_13200,N_12826,N_12825);
xnor U13201 (N_13201,N_12767,N_12940);
nand U13202 (N_13202,N_12782,N_12839);
or U13203 (N_13203,N_12884,N_12867);
nand U13204 (N_13204,N_12802,N_12845);
xor U13205 (N_13205,N_12937,N_12896);
and U13206 (N_13206,N_12783,N_12917);
and U13207 (N_13207,N_12826,N_12902);
or U13208 (N_13208,N_12863,N_12837);
nor U13209 (N_13209,N_12914,N_12846);
and U13210 (N_13210,N_12982,N_12936);
or U13211 (N_13211,N_12925,N_12977);
nor U13212 (N_13212,N_12752,N_12782);
or U13213 (N_13213,N_12878,N_12972);
and U13214 (N_13214,N_12824,N_12956);
and U13215 (N_13215,N_12920,N_12957);
or U13216 (N_13216,N_12819,N_12833);
nand U13217 (N_13217,N_12985,N_12851);
xnor U13218 (N_13218,N_12983,N_12949);
nand U13219 (N_13219,N_12762,N_12825);
nor U13220 (N_13220,N_12816,N_12954);
nor U13221 (N_13221,N_12886,N_12802);
nand U13222 (N_13222,N_12871,N_12824);
and U13223 (N_13223,N_12806,N_12927);
nor U13224 (N_13224,N_12954,N_12989);
nor U13225 (N_13225,N_12944,N_12962);
or U13226 (N_13226,N_12891,N_12790);
or U13227 (N_13227,N_12966,N_12766);
or U13228 (N_13228,N_12788,N_12881);
or U13229 (N_13229,N_12857,N_12985);
xor U13230 (N_13230,N_12842,N_12986);
nand U13231 (N_13231,N_12750,N_12859);
or U13232 (N_13232,N_12934,N_12977);
xor U13233 (N_13233,N_12881,N_12860);
nor U13234 (N_13234,N_12953,N_12777);
nor U13235 (N_13235,N_12845,N_12947);
or U13236 (N_13236,N_12988,N_12943);
or U13237 (N_13237,N_12917,N_12772);
nor U13238 (N_13238,N_12853,N_12959);
nor U13239 (N_13239,N_12938,N_12943);
nand U13240 (N_13240,N_12860,N_12882);
and U13241 (N_13241,N_12881,N_12774);
nor U13242 (N_13242,N_12828,N_12865);
nor U13243 (N_13243,N_12880,N_12918);
xor U13244 (N_13244,N_12931,N_12932);
nor U13245 (N_13245,N_12802,N_12883);
or U13246 (N_13246,N_12804,N_12964);
xor U13247 (N_13247,N_12960,N_12854);
nand U13248 (N_13248,N_12968,N_12818);
and U13249 (N_13249,N_12784,N_12881);
or U13250 (N_13250,N_13008,N_13017);
and U13251 (N_13251,N_13188,N_13165);
xnor U13252 (N_13252,N_13013,N_13241);
nand U13253 (N_13253,N_13187,N_13189);
xor U13254 (N_13254,N_13006,N_13193);
nand U13255 (N_13255,N_13054,N_13098);
and U13256 (N_13256,N_13103,N_13076);
nand U13257 (N_13257,N_13102,N_13005);
xnor U13258 (N_13258,N_13124,N_13221);
and U13259 (N_13259,N_13222,N_13195);
or U13260 (N_13260,N_13121,N_13063);
nor U13261 (N_13261,N_13247,N_13055);
nand U13262 (N_13262,N_13060,N_13171);
or U13263 (N_13263,N_13248,N_13153);
nor U13264 (N_13264,N_13068,N_13020);
or U13265 (N_13265,N_13021,N_13071);
or U13266 (N_13266,N_13002,N_13082);
nor U13267 (N_13267,N_13242,N_13035);
xnor U13268 (N_13268,N_13166,N_13186);
and U13269 (N_13269,N_13125,N_13133);
nor U13270 (N_13270,N_13000,N_13105);
nor U13271 (N_13271,N_13224,N_13137);
nand U13272 (N_13272,N_13096,N_13225);
nor U13273 (N_13273,N_13040,N_13173);
and U13274 (N_13274,N_13205,N_13119);
nor U13275 (N_13275,N_13232,N_13025);
nand U13276 (N_13276,N_13135,N_13163);
nor U13277 (N_13277,N_13145,N_13080);
or U13278 (N_13278,N_13052,N_13238);
xor U13279 (N_13279,N_13095,N_13059);
xor U13280 (N_13280,N_13118,N_13162);
or U13281 (N_13281,N_13149,N_13034);
xnor U13282 (N_13282,N_13010,N_13159);
nand U13283 (N_13283,N_13164,N_13061);
nand U13284 (N_13284,N_13139,N_13074);
nor U13285 (N_13285,N_13069,N_13246);
or U13286 (N_13286,N_13231,N_13038);
nand U13287 (N_13287,N_13219,N_13203);
xnor U13288 (N_13288,N_13182,N_13104);
xor U13289 (N_13289,N_13051,N_13218);
xor U13290 (N_13290,N_13049,N_13113);
and U13291 (N_13291,N_13023,N_13101);
nor U13292 (N_13292,N_13147,N_13243);
xor U13293 (N_13293,N_13152,N_13122);
nor U13294 (N_13294,N_13200,N_13184);
nand U13295 (N_13295,N_13183,N_13198);
or U13296 (N_13296,N_13202,N_13086);
xnor U13297 (N_13297,N_13097,N_13141);
and U13298 (N_13298,N_13046,N_13026);
nand U13299 (N_13299,N_13134,N_13047);
nor U13300 (N_13300,N_13204,N_13024);
xor U13301 (N_13301,N_13110,N_13078);
or U13302 (N_13302,N_13111,N_13011);
xor U13303 (N_13303,N_13131,N_13199);
and U13304 (N_13304,N_13083,N_13037);
and U13305 (N_13305,N_13053,N_13123);
and U13306 (N_13306,N_13003,N_13245);
nor U13307 (N_13307,N_13239,N_13197);
and U13308 (N_13308,N_13213,N_13072);
nor U13309 (N_13309,N_13108,N_13227);
xnor U13310 (N_13310,N_13033,N_13235);
xor U13311 (N_13311,N_13176,N_13027);
xnor U13312 (N_13312,N_13009,N_13174);
nor U13313 (N_13313,N_13081,N_13158);
xor U13314 (N_13314,N_13144,N_13223);
xnor U13315 (N_13315,N_13194,N_13154);
nand U13316 (N_13316,N_13178,N_13177);
nand U13317 (N_13317,N_13093,N_13240);
xor U13318 (N_13318,N_13128,N_13062);
nand U13319 (N_13319,N_13042,N_13018);
xnor U13320 (N_13320,N_13136,N_13206);
and U13321 (N_13321,N_13112,N_13032);
nand U13322 (N_13322,N_13016,N_13126);
nand U13323 (N_13323,N_13129,N_13015);
xnor U13324 (N_13324,N_13155,N_13211);
and U13325 (N_13325,N_13022,N_13120);
and U13326 (N_13326,N_13036,N_13099);
or U13327 (N_13327,N_13043,N_13161);
xor U13328 (N_13328,N_13192,N_13181);
nand U13329 (N_13329,N_13116,N_13220);
or U13330 (N_13330,N_13100,N_13210);
and U13331 (N_13331,N_13212,N_13207);
xor U13332 (N_13332,N_13065,N_13115);
nor U13333 (N_13333,N_13057,N_13226);
and U13334 (N_13334,N_13169,N_13019);
nand U13335 (N_13335,N_13185,N_13058);
and U13336 (N_13336,N_13170,N_13090);
and U13337 (N_13337,N_13091,N_13175);
nor U13338 (N_13338,N_13044,N_13109);
nor U13339 (N_13339,N_13031,N_13039);
nor U13340 (N_13340,N_13014,N_13216);
nor U13341 (N_13341,N_13012,N_13067);
xnor U13342 (N_13342,N_13208,N_13114);
or U13343 (N_13343,N_13070,N_13087);
xor U13344 (N_13344,N_13196,N_13088);
xor U13345 (N_13345,N_13004,N_13030);
xnor U13346 (N_13346,N_13138,N_13092);
and U13347 (N_13347,N_13094,N_13230);
and U13348 (N_13348,N_13064,N_13146);
or U13349 (N_13349,N_13191,N_13179);
xnor U13350 (N_13350,N_13156,N_13107);
or U13351 (N_13351,N_13130,N_13127);
nor U13352 (N_13352,N_13150,N_13249);
and U13353 (N_13353,N_13229,N_13048);
and U13354 (N_13354,N_13079,N_13140);
nand U13355 (N_13355,N_13132,N_13106);
nor U13356 (N_13356,N_13157,N_13045);
nor U13357 (N_13357,N_13172,N_13180);
or U13358 (N_13358,N_13244,N_13234);
nand U13359 (N_13359,N_13084,N_13041);
or U13360 (N_13360,N_13056,N_13236);
xnor U13361 (N_13361,N_13075,N_13117);
and U13362 (N_13362,N_13201,N_13228);
nand U13363 (N_13363,N_13001,N_13151);
or U13364 (N_13364,N_13077,N_13143);
or U13365 (N_13365,N_13028,N_13237);
xor U13366 (N_13366,N_13066,N_13217);
or U13367 (N_13367,N_13050,N_13215);
or U13368 (N_13368,N_13007,N_13085);
nor U13369 (N_13369,N_13148,N_13233);
xor U13370 (N_13370,N_13214,N_13089);
and U13371 (N_13371,N_13168,N_13167);
nand U13372 (N_13372,N_13160,N_13142);
nor U13373 (N_13373,N_13029,N_13073);
or U13374 (N_13374,N_13190,N_13209);
and U13375 (N_13375,N_13057,N_13078);
xnor U13376 (N_13376,N_13241,N_13074);
or U13377 (N_13377,N_13233,N_13094);
nand U13378 (N_13378,N_13063,N_13190);
or U13379 (N_13379,N_13061,N_13092);
and U13380 (N_13380,N_13196,N_13106);
or U13381 (N_13381,N_13075,N_13085);
or U13382 (N_13382,N_13092,N_13188);
and U13383 (N_13383,N_13091,N_13181);
nand U13384 (N_13384,N_13016,N_13249);
xor U13385 (N_13385,N_13013,N_13025);
or U13386 (N_13386,N_13195,N_13187);
and U13387 (N_13387,N_13104,N_13247);
nand U13388 (N_13388,N_13111,N_13093);
xnor U13389 (N_13389,N_13010,N_13084);
and U13390 (N_13390,N_13013,N_13102);
xnor U13391 (N_13391,N_13098,N_13103);
nor U13392 (N_13392,N_13066,N_13182);
or U13393 (N_13393,N_13227,N_13127);
or U13394 (N_13394,N_13058,N_13234);
xnor U13395 (N_13395,N_13055,N_13161);
xnor U13396 (N_13396,N_13018,N_13121);
nor U13397 (N_13397,N_13144,N_13012);
nand U13398 (N_13398,N_13017,N_13182);
nand U13399 (N_13399,N_13187,N_13063);
xnor U13400 (N_13400,N_13096,N_13033);
or U13401 (N_13401,N_13045,N_13195);
and U13402 (N_13402,N_13151,N_13057);
or U13403 (N_13403,N_13005,N_13176);
xor U13404 (N_13404,N_13036,N_13101);
xor U13405 (N_13405,N_13011,N_13212);
nor U13406 (N_13406,N_13113,N_13191);
or U13407 (N_13407,N_13044,N_13024);
xor U13408 (N_13408,N_13088,N_13092);
and U13409 (N_13409,N_13162,N_13205);
and U13410 (N_13410,N_13006,N_13135);
or U13411 (N_13411,N_13182,N_13162);
and U13412 (N_13412,N_13226,N_13149);
and U13413 (N_13413,N_13247,N_13110);
nand U13414 (N_13414,N_13152,N_13017);
nor U13415 (N_13415,N_13008,N_13144);
or U13416 (N_13416,N_13220,N_13074);
xnor U13417 (N_13417,N_13093,N_13177);
xnor U13418 (N_13418,N_13068,N_13218);
nand U13419 (N_13419,N_13178,N_13223);
xnor U13420 (N_13420,N_13005,N_13014);
or U13421 (N_13421,N_13110,N_13217);
xor U13422 (N_13422,N_13203,N_13025);
xnor U13423 (N_13423,N_13168,N_13130);
and U13424 (N_13424,N_13130,N_13154);
or U13425 (N_13425,N_13013,N_13038);
or U13426 (N_13426,N_13066,N_13104);
or U13427 (N_13427,N_13046,N_13168);
nand U13428 (N_13428,N_13109,N_13178);
nand U13429 (N_13429,N_13225,N_13077);
xor U13430 (N_13430,N_13191,N_13164);
xnor U13431 (N_13431,N_13063,N_13248);
xnor U13432 (N_13432,N_13186,N_13146);
xor U13433 (N_13433,N_13188,N_13213);
and U13434 (N_13434,N_13087,N_13175);
nand U13435 (N_13435,N_13220,N_13005);
or U13436 (N_13436,N_13208,N_13055);
and U13437 (N_13437,N_13153,N_13182);
xnor U13438 (N_13438,N_13048,N_13215);
or U13439 (N_13439,N_13129,N_13237);
or U13440 (N_13440,N_13075,N_13011);
nor U13441 (N_13441,N_13108,N_13125);
xnor U13442 (N_13442,N_13135,N_13122);
nor U13443 (N_13443,N_13231,N_13113);
or U13444 (N_13444,N_13136,N_13127);
nor U13445 (N_13445,N_13202,N_13227);
or U13446 (N_13446,N_13120,N_13110);
and U13447 (N_13447,N_13018,N_13192);
nand U13448 (N_13448,N_13086,N_13058);
and U13449 (N_13449,N_13167,N_13134);
and U13450 (N_13450,N_13103,N_13190);
nand U13451 (N_13451,N_13102,N_13077);
and U13452 (N_13452,N_13047,N_13125);
and U13453 (N_13453,N_13182,N_13222);
or U13454 (N_13454,N_13205,N_13123);
nand U13455 (N_13455,N_13187,N_13209);
nand U13456 (N_13456,N_13214,N_13038);
nor U13457 (N_13457,N_13186,N_13128);
nor U13458 (N_13458,N_13058,N_13233);
nand U13459 (N_13459,N_13005,N_13101);
or U13460 (N_13460,N_13249,N_13226);
nor U13461 (N_13461,N_13186,N_13249);
and U13462 (N_13462,N_13137,N_13027);
or U13463 (N_13463,N_13017,N_13200);
and U13464 (N_13464,N_13096,N_13183);
xor U13465 (N_13465,N_13186,N_13169);
or U13466 (N_13466,N_13179,N_13174);
nor U13467 (N_13467,N_13054,N_13141);
and U13468 (N_13468,N_13069,N_13012);
and U13469 (N_13469,N_13006,N_13166);
xnor U13470 (N_13470,N_13025,N_13207);
or U13471 (N_13471,N_13184,N_13031);
and U13472 (N_13472,N_13187,N_13046);
and U13473 (N_13473,N_13051,N_13054);
or U13474 (N_13474,N_13131,N_13130);
xor U13475 (N_13475,N_13238,N_13128);
and U13476 (N_13476,N_13153,N_13208);
nand U13477 (N_13477,N_13035,N_13115);
nor U13478 (N_13478,N_13093,N_13054);
and U13479 (N_13479,N_13095,N_13201);
nor U13480 (N_13480,N_13179,N_13202);
or U13481 (N_13481,N_13019,N_13125);
or U13482 (N_13482,N_13050,N_13074);
nor U13483 (N_13483,N_13238,N_13184);
nor U13484 (N_13484,N_13193,N_13232);
or U13485 (N_13485,N_13078,N_13241);
or U13486 (N_13486,N_13208,N_13210);
and U13487 (N_13487,N_13040,N_13138);
or U13488 (N_13488,N_13213,N_13073);
nor U13489 (N_13489,N_13196,N_13082);
and U13490 (N_13490,N_13018,N_13112);
nor U13491 (N_13491,N_13146,N_13172);
nand U13492 (N_13492,N_13249,N_13171);
or U13493 (N_13493,N_13023,N_13235);
or U13494 (N_13494,N_13190,N_13232);
and U13495 (N_13495,N_13187,N_13049);
xor U13496 (N_13496,N_13214,N_13180);
nand U13497 (N_13497,N_13029,N_13008);
nor U13498 (N_13498,N_13108,N_13174);
or U13499 (N_13499,N_13065,N_13210);
xor U13500 (N_13500,N_13392,N_13447);
nand U13501 (N_13501,N_13271,N_13301);
xnor U13502 (N_13502,N_13329,N_13395);
or U13503 (N_13503,N_13302,N_13410);
or U13504 (N_13504,N_13379,N_13378);
or U13505 (N_13505,N_13261,N_13473);
xor U13506 (N_13506,N_13364,N_13334);
or U13507 (N_13507,N_13460,N_13403);
or U13508 (N_13508,N_13297,N_13282);
xor U13509 (N_13509,N_13421,N_13402);
or U13510 (N_13510,N_13435,N_13423);
nor U13511 (N_13511,N_13414,N_13448);
or U13512 (N_13512,N_13331,N_13474);
nand U13513 (N_13513,N_13366,N_13468);
nand U13514 (N_13514,N_13283,N_13461);
xor U13515 (N_13515,N_13493,N_13259);
or U13516 (N_13516,N_13312,N_13342);
xnor U13517 (N_13517,N_13360,N_13376);
or U13518 (N_13518,N_13340,N_13477);
and U13519 (N_13519,N_13464,N_13452);
and U13520 (N_13520,N_13308,N_13499);
nor U13521 (N_13521,N_13272,N_13491);
or U13522 (N_13522,N_13482,N_13253);
xnor U13523 (N_13523,N_13412,N_13257);
and U13524 (N_13524,N_13390,N_13486);
xnor U13525 (N_13525,N_13305,N_13455);
or U13526 (N_13526,N_13432,N_13325);
or U13527 (N_13527,N_13362,N_13319);
xor U13528 (N_13528,N_13451,N_13462);
or U13529 (N_13529,N_13408,N_13430);
nand U13530 (N_13530,N_13459,N_13489);
nand U13531 (N_13531,N_13300,N_13442);
xor U13532 (N_13532,N_13295,N_13434);
nor U13533 (N_13533,N_13490,N_13268);
nor U13534 (N_13534,N_13481,N_13384);
nor U13535 (N_13535,N_13438,N_13327);
nand U13536 (N_13536,N_13391,N_13393);
nand U13537 (N_13537,N_13396,N_13496);
nor U13538 (N_13538,N_13322,N_13356);
or U13539 (N_13539,N_13266,N_13250);
or U13540 (N_13540,N_13280,N_13483);
xor U13541 (N_13541,N_13457,N_13404);
nand U13542 (N_13542,N_13344,N_13478);
nand U13543 (N_13543,N_13353,N_13374);
xor U13544 (N_13544,N_13277,N_13424);
or U13545 (N_13545,N_13357,N_13270);
xor U13546 (N_13546,N_13429,N_13497);
xnor U13547 (N_13547,N_13258,N_13389);
nand U13548 (N_13548,N_13400,N_13467);
and U13549 (N_13549,N_13426,N_13458);
nor U13550 (N_13550,N_13273,N_13354);
nor U13551 (N_13551,N_13341,N_13407);
and U13552 (N_13552,N_13278,N_13363);
nand U13553 (N_13553,N_13454,N_13425);
nand U13554 (N_13554,N_13355,N_13323);
or U13555 (N_13555,N_13262,N_13388);
and U13556 (N_13556,N_13446,N_13326);
or U13557 (N_13557,N_13351,N_13383);
nor U13558 (N_13558,N_13399,N_13381);
nor U13559 (N_13559,N_13313,N_13370);
nand U13560 (N_13560,N_13321,N_13416);
or U13561 (N_13561,N_13494,N_13449);
xor U13562 (N_13562,N_13328,N_13309);
and U13563 (N_13563,N_13263,N_13445);
and U13564 (N_13564,N_13398,N_13317);
and U13565 (N_13565,N_13385,N_13456);
and U13566 (N_13566,N_13469,N_13346);
nand U13567 (N_13567,N_13413,N_13476);
or U13568 (N_13568,N_13251,N_13420);
nor U13569 (N_13569,N_13475,N_13394);
nor U13570 (N_13570,N_13397,N_13372);
or U13571 (N_13571,N_13289,N_13359);
or U13572 (N_13572,N_13304,N_13316);
or U13573 (N_13573,N_13286,N_13350);
nand U13574 (N_13574,N_13288,N_13495);
nand U13575 (N_13575,N_13433,N_13307);
nor U13576 (N_13576,N_13336,N_13401);
and U13577 (N_13577,N_13439,N_13252);
or U13578 (N_13578,N_13338,N_13419);
nand U13579 (N_13579,N_13443,N_13298);
or U13580 (N_13580,N_13260,N_13367);
and U13581 (N_13581,N_13275,N_13311);
or U13582 (N_13582,N_13352,N_13256);
nor U13583 (N_13583,N_13290,N_13373);
nand U13584 (N_13584,N_13267,N_13371);
xor U13585 (N_13585,N_13382,N_13294);
nor U13586 (N_13586,N_13436,N_13492);
nor U13587 (N_13587,N_13296,N_13337);
nand U13588 (N_13588,N_13314,N_13406);
nand U13589 (N_13589,N_13409,N_13318);
and U13590 (N_13590,N_13377,N_13293);
and U13591 (N_13591,N_13343,N_13437);
or U13592 (N_13592,N_13466,N_13292);
nor U13593 (N_13593,N_13361,N_13265);
and U13594 (N_13594,N_13375,N_13345);
nand U13595 (N_13595,N_13417,N_13450);
nor U13596 (N_13596,N_13369,N_13387);
or U13597 (N_13597,N_13485,N_13349);
nand U13598 (N_13598,N_13330,N_13324);
or U13599 (N_13599,N_13358,N_13471);
nand U13600 (N_13600,N_13276,N_13418);
nor U13601 (N_13601,N_13310,N_13422);
or U13602 (N_13602,N_13333,N_13415);
nand U13603 (N_13603,N_13405,N_13264);
nor U13604 (N_13604,N_13303,N_13484);
nand U13605 (N_13605,N_13480,N_13441);
xor U13606 (N_13606,N_13281,N_13299);
nand U13607 (N_13607,N_13320,N_13453);
or U13608 (N_13608,N_13488,N_13440);
nor U13609 (N_13609,N_13315,N_13335);
xnor U13610 (N_13610,N_13487,N_13285);
nor U13611 (N_13611,N_13306,N_13470);
and U13612 (N_13612,N_13368,N_13255);
nor U13613 (N_13613,N_13284,N_13347);
xnor U13614 (N_13614,N_13348,N_13428);
nand U13615 (N_13615,N_13287,N_13365);
nor U13616 (N_13616,N_13386,N_13444);
nand U13617 (N_13617,N_13279,N_13411);
nor U13618 (N_13618,N_13463,N_13269);
nand U13619 (N_13619,N_13274,N_13380);
nor U13620 (N_13620,N_13291,N_13498);
nor U13621 (N_13621,N_13431,N_13427);
nand U13622 (N_13622,N_13472,N_13254);
nand U13623 (N_13623,N_13332,N_13339);
and U13624 (N_13624,N_13465,N_13479);
and U13625 (N_13625,N_13474,N_13295);
nand U13626 (N_13626,N_13365,N_13451);
xnor U13627 (N_13627,N_13269,N_13481);
nor U13628 (N_13628,N_13434,N_13369);
nor U13629 (N_13629,N_13285,N_13469);
or U13630 (N_13630,N_13398,N_13492);
and U13631 (N_13631,N_13487,N_13350);
and U13632 (N_13632,N_13379,N_13479);
nand U13633 (N_13633,N_13325,N_13482);
and U13634 (N_13634,N_13423,N_13495);
and U13635 (N_13635,N_13353,N_13313);
or U13636 (N_13636,N_13413,N_13389);
and U13637 (N_13637,N_13262,N_13323);
xnor U13638 (N_13638,N_13409,N_13283);
nand U13639 (N_13639,N_13462,N_13311);
nand U13640 (N_13640,N_13344,N_13445);
nor U13641 (N_13641,N_13377,N_13308);
and U13642 (N_13642,N_13323,N_13472);
or U13643 (N_13643,N_13253,N_13430);
and U13644 (N_13644,N_13386,N_13394);
and U13645 (N_13645,N_13258,N_13252);
nand U13646 (N_13646,N_13331,N_13276);
nand U13647 (N_13647,N_13410,N_13424);
and U13648 (N_13648,N_13329,N_13298);
and U13649 (N_13649,N_13492,N_13469);
nor U13650 (N_13650,N_13339,N_13491);
xnor U13651 (N_13651,N_13412,N_13483);
xnor U13652 (N_13652,N_13484,N_13300);
nand U13653 (N_13653,N_13336,N_13304);
nand U13654 (N_13654,N_13489,N_13365);
nand U13655 (N_13655,N_13328,N_13266);
and U13656 (N_13656,N_13297,N_13261);
xnor U13657 (N_13657,N_13288,N_13472);
nor U13658 (N_13658,N_13380,N_13429);
and U13659 (N_13659,N_13275,N_13397);
or U13660 (N_13660,N_13499,N_13411);
xnor U13661 (N_13661,N_13457,N_13263);
or U13662 (N_13662,N_13445,N_13498);
and U13663 (N_13663,N_13444,N_13301);
xor U13664 (N_13664,N_13481,N_13372);
xor U13665 (N_13665,N_13313,N_13392);
and U13666 (N_13666,N_13424,N_13284);
nor U13667 (N_13667,N_13332,N_13405);
or U13668 (N_13668,N_13330,N_13476);
and U13669 (N_13669,N_13437,N_13253);
or U13670 (N_13670,N_13446,N_13490);
and U13671 (N_13671,N_13275,N_13369);
xnor U13672 (N_13672,N_13411,N_13399);
and U13673 (N_13673,N_13297,N_13456);
nand U13674 (N_13674,N_13265,N_13435);
nand U13675 (N_13675,N_13373,N_13487);
nor U13676 (N_13676,N_13294,N_13407);
nor U13677 (N_13677,N_13335,N_13393);
xnor U13678 (N_13678,N_13408,N_13328);
xnor U13679 (N_13679,N_13404,N_13492);
nand U13680 (N_13680,N_13416,N_13423);
nand U13681 (N_13681,N_13467,N_13435);
xnor U13682 (N_13682,N_13447,N_13475);
or U13683 (N_13683,N_13478,N_13408);
nor U13684 (N_13684,N_13340,N_13492);
and U13685 (N_13685,N_13330,N_13272);
and U13686 (N_13686,N_13328,N_13322);
nor U13687 (N_13687,N_13301,N_13427);
xnor U13688 (N_13688,N_13408,N_13275);
nor U13689 (N_13689,N_13320,N_13251);
or U13690 (N_13690,N_13266,N_13332);
and U13691 (N_13691,N_13322,N_13436);
nor U13692 (N_13692,N_13337,N_13458);
or U13693 (N_13693,N_13268,N_13453);
nand U13694 (N_13694,N_13463,N_13419);
nand U13695 (N_13695,N_13442,N_13294);
xnor U13696 (N_13696,N_13381,N_13426);
or U13697 (N_13697,N_13481,N_13415);
xor U13698 (N_13698,N_13256,N_13252);
nand U13699 (N_13699,N_13451,N_13397);
nor U13700 (N_13700,N_13463,N_13444);
or U13701 (N_13701,N_13306,N_13316);
or U13702 (N_13702,N_13402,N_13418);
and U13703 (N_13703,N_13277,N_13324);
and U13704 (N_13704,N_13425,N_13464);
and U13705 (N_13705,N_13302,N_13365);
nor U13706 (N_13706,N_13276,N_13488);
nand U13707 (N_13707,N_13362,N_13468);
and U13708 (N_13708,N_13342,N_13268);
or U13709 (N_13709,N_13279,N_13294);
nand U13710 (N_13710,N_13452,N_13294);
nand U13711 (N_13711,N_13286,N_13378);
or U13712 (N_13712,N_13323,N_13361);
nand U13713 (N_13713,N_13389,N_13453);
nand U13714 (N_13714,N_13343,N_13430);
and U13715 (N_13715,N_13343,N_13449);
nand U13716 (N_13716,N_13365,N_13370);
or U13717 (N_13717,N_13440,N_13317);
nand U13718 (N_13718,N_13271,N_13279);
nor U13719 (N_13719,N_13314,N_13298);
and U13720 (N_13720,N_13305,N_13395);
nand U13721 (N_13721,N_13254,N_13497);
and U13722 (N_13722,N_13315,N_13366);
and U13723 (N_13723,N_13448,N_13472);
nor U13724 (N_13724,N_13393,N_13445);
nor U13725 (N_13725,N_13476,N_13376);
nand U13726 (N_13726,N_13469,N_13289);
nor U13727 (N_13727,N_13315,N_13392);
and U13728 (N_13728,N_13384,N_13456);
xor U13729 (N_13729,N_13477,N_13303);
nor U13730 (N_13730,N_13268,N_13324);
nor U13731 (N_13731,N_13367,N_13294);
nand U13732 (N_13732,N_13490,N_13468);
nand U13733 (N_13733,N_13451,N_13327);
or U13734 (N_13734,N_13268,N_13445);
nor U13735 (N_13735,N_13287,N_13254);
and U13736 (N_13736,N_13437,N_13387);
xor U13737 (N_13737,N_13319,N_13415);
and U13738 (N_13738,N_13412,N_13473);
nor U13739 (N_13739,N_13348,N_13297);
or U13740 (N_13740,N_13273,N_13264);
xnor U13741 (N_13741,N_13261,N_13332);
and U13742 (N_13742,N_13416,N_13364);
or U13743 (N_13743,N_13458,N_13285);
xnor U13744 (N_13744,N_13447,N_13335);
nand U13745 (N_13745,N_13291,N_13423);
xor U13746 (N_13746,N_13290,N_13292);
or U13747 (N_13747,N_13381,N_13457);
xor U13748 (N_13748,N_13373,N_13330);
or U13749 (N_13749,N_13349,N_13297);
nand U13750 (N_13750,N_13607,N_13576);
and U13751 (N_13751,N_13728,N_13634);
xnor U13752 (N_13752,N_13549,N_13726);
nand U13753 (N_13753,N_13725,N_13727);
and U13754 (N_13754,N_13526,N_13633);
and U13755 (N_13755,N_13595,N_13560);
nand U13756 (N_13756,N_13567,N_13628);
and U13757 (N_13757,N_13653,N_13661);
nand U13758 (N_13758,N_13647,N_13699);
nand U13759 (N_13759,N_13606,N_13627);
and U13760 (N_13760,N_13702,N_13742);
xor U13761 (N_13761,N_13687,N_13671);
nand U13762 (N_13762,N_13617,N_13692);
xnor U13763 (N_13763,N_13676,N_13685);
xnor U13764 (N_13764,N_13715,N_13650);
and U13765 (N_13765,N_13580,N_13528);
or U13766 (N_13766,N_13645,N_13609);
and U13767 (N_13767,N_13613,N_13679);
nand U13768 (N_13768,N_13590,N_13736);
nor U13769 (N_13769,N_13608,N_13629);
nand U13770 (N_13770,N_13536,N_13593);
xnor U13771 (N_13771,N_13743,N_13641);
or U13772 (N_13772,N_13698,N_13573);
xor U13773 (N_13773,N_13550,N_13731);
nand U13774 (N_13774,N_13594,N_13582);
and U13775 (N_13775,N_13733,N_13616);
xnor U13776 (N_13776,N_13561,N_13714);
and U13777 (N_13777,N_13600,N_13720);
nand U13778 (N_13778,N_13730,N_13552);
and U13779 (N_13779,N_13626,N_13522);
or U13780 (N_13780,N_13555,N_13525);
nand U13781 (N_13781,N_13716,N_13683);
nand U13782 (N_13782,N_13507,N_13677);
nor U13783 (N_13783,N_13592,N_13689);
xor U13784 (N_13784,N_13533,N_13579);
nand U13785 (N_13785,N_13691,N_13568);
and U13786 (N_13786,N_13631,N_13669);
and U13787 (N_13787,N_13710,N_13625);
or U13788 (N_13788,N_13635,N_13638);
or U13789 (N_13789,N_13734,N_13547);
or U13790 (N_13790,N_13610,N_13519);
xnor U13791 (N_13791,N_13705,N_13503);
nor U13792 (N_13792,N_13707,N_13701);
and U13793 (N_13793,N_13672,N_13680);
nand U13794 (N_13794,N_13735,N_13575);
nand U13795 (N_13795,N_13603,N_13581);
nand U13796 (N_13796,N_13623,N_13660);
xor U13797 (N_13797,N_13697,N_13696);
or U13798 (N_13798,N_13515,N_13674);
nand U13799 (N_13799,N_13518,N_13663);
nand U13800 (N_13800,N_13665,N_13597);
nor U13801 (N_13801,N_13570,N_13658);
or U13802 (N_13802,N_13695,N_13614);
and U13803 (N_13803,N_13723,N_13513);
nor U13804 (N_13804,N_13618,N_13559);
xor U13805 (N_13805,N_13521,N_13530);
nand U13806 (N_13806,N_13646,N_13502);
and U13807 (N_13807,N_13557,N_13583);
xnor U13808 (N_13808,N_13682,N_13666);
xor U13809 (N_13809,N_13588,N_13585);
or U13810 (N_13810,N_13640,N_13556);
or U13811 (N_13811,N_13621,N_13572);
nand U13812 (N_13812,N_13668,N_13688);
xor U13813 (N_13813,N_13748,N_13694);
nand U13814 (N_13814,N_13745,N_13541);
nand U13815 (N_13815,N_13520,N_13622);
nand U13816 (N_13816,N_13577,N_13620);
and U13817 (N_13817,N_13574,N_13708);
nor U13818 (N_13818,N_13670,N_13554);
nand U13819 (N_13819,N_13558,N_13690);
xor U13820 (N_13820,N_13605,N_13721);
nand U13821 (N_13821,N_13540,N_13667);
xor U13822 (N_13822,N_13543,N_13589);
or U13823 (N_13823,N_13739,N_13706);
xor U13824 (N_13824,N_13601,N_13532);
nor U13825 (N_13825,N_13531,N_13704);
nor U13826 (N_13826,N_13678,N_13504);
nor U13827 (N_13827,N_13612,N_13713);
nor U13828 (N_13828,N_13615,N_13534);
nor U13829 (N_13829,N_13586,N_13546);
and U13830 (N_13830,N_13569,N_13539);
xnor U13831 (N_13831,N_13587,N_13566);
nor U13832 (N_13832,N_13722,N_13740);
and U13833 (N_13833,N_13508,N_13738);
nand U13834 (N_13834,N_13724,N_13524);
xor U13835 (N_13835,N_13505,N_13654);
or U13836 (N_13836,N_13675,N_13510);
nand U13837 (N_13837,N_13729,N_13564);
nor U13838 (N_13838,N_13516,N_13604);
and U13839 (N_13839,N_13718,N_13624);
nor U13840 (N_13840,N_13664,N_13709);
or U13841 (N_13841,N_13749,N_13644);
nor U13842 (N_13842,N_13686,N_13542);
and U13843 (N_13843,N_13662,N_13717);
and U13844 (N_13844,N_13512,N_13591);
and U13845 (N_13845,N_13642,N_13548);
nor U13846 (N_13846,N_13719,N_13632);
nor U13847 (N_13847,N_13712,N_13596);
and U13848 (N_13848,N_13732,N_13700);
and U13849 (N_13849,N_13500,N_13703);
xnor U13850 (N_13850,N_13655,N_13538);
and U13851 (N_13851,N_13648,N_13649);
or U13852 (N_13852,N_13673,N_13527);
nor U13853 (N_13853,N_13684,N_13602);
and U13854 (N_13854,N_13501,N_13611);
nor U13855 (N_13855,N_13565,N_13529);
nand U13856 (N_13856,N_13514,N_13659);
nand U13857 (N_13857,N_13657,N_13509);
xnor U13858 (N_13858,N_13523,N_13746);
and U13859 (N_13859,N_13741,N_13711);
nor U13860 (N_13860,N_13630,N_13639);
or U13861 (N_13861,N_13744,N_13643);
nand U13862 (N_13862,N_13652,N_13544);
nor U13863 (N_13863,N_13506,N_13656);
xnor U13864 (N_13864,N_13551,N_13598);
and U13865 (N_13865,N_13599,N_13517);
nand U13866 (N_13866,N_13636,N_13537);
nand U13867 (N_13867,N_13562,N_13747);
or U13868 (N_13868,N_13651,N_13619);
or U13869 (N_13869,N_13637,N_13578);
and U13870 (N_13870,N_13681,N_13693);
or U13871 (N_13871,N_13545,N_13584);
and U13872 (N_13872,N_13553,N_13563);
nor U13873 (N_13873,N_13511,N_13571);
and U13874 (N_13874,N_13737,N_13535);
nor U13875 (N_13875,N_13520,N_13748);
and U13876 (N_13876,N_13692,N_13570);
nor U13877 (N_13877,N_13608,N_13645);
nor U13878 (N_13878,N_13701,N_13548);
nor U13879 (N_13879,N_13538,N_13598);
nand U13880 (N_13880,N_13546,N_13697);
nor U13881 (N_13881,N_13689,N_13602);
or U13882 (N_13882,N_13633,N_13583);
or U13883 (N_13883,N_13545,N_13578);
and U13884 (N_13884,N_13549,N_13530);
or U13885 (N_13885,N_13714,N_13590);
xnor U13886 (N_13886,N_13601,N_13594);
nand U13887 (N_13887,N_13556,N_13539);
xor U13888 (N_13888,N_13600,N_13724);
and U13889 (N_13889,N_13732,N_13513);
and U13890 (N_13890,N_13531,N_13502);
nand U13891 (N_13891,N_13599,N_13641);
xor U13892 (N_13892,N_13683,N_13619);
nand U13893 (N_13893,N_13701,N_13666);
nor U13894 (N_13894,N_13514,N_13687);
and U13895 (N_13895,N_13687,N_13559);
and U13896 (N_13896,N_13619,N_13544);
or U13897 (N_13897,N_13656,N_13563);
and U13898 (N_13898,N_13695,N_13570);
xnor U13899 (N_13899,N_13549,N_13746);
nor U13900 (N_13900,N_13714,N_13693);
nor U13901 (N_13901,N_13534,N_13504);
and U13902 (N_13902,N_13596,N_13577);
nand U13903 (N_13903,N_13554,N_13651);
xnor U13904 (N_13904,N_13548,N_13569);
xor U13905 (N_13905,N_13672,N_13684);
nor U13906 (N_13906,N_13673,N_13688);
or U13907 (N_13907,N_13728,N_13595);
xor U13908 (N_13908,N_13704,N_13728);
nor U13909 (N_13909,N_13557,N_13737);
or U13910 (N_13910,N_13719,N_13537);
and U13911 (N_13911,N_13700,N_13661);
nor U13912 (N_13912,N_13542,N_13575);
and U13913 (N_13913,N_13556,N_13537);
or U13914 (N_13914,N_13708,N_13597);
nand U13915 (N_13915,N_13741,N_13594);
nor U13916 (N_13916,N_13610,N_13591);
nand U13917 (N_13917,N_13598,N_13507);
and U13918 (N_13918,N_13606,N_13667);
and U13919 (N_13919,N_13500,N_13631);
and U13920 (N_13920,N_13674,N_13671);
nor U13921 (N_13921,N_13604,N_13724);
or U13922 (N_13922,N_13719,N_13593);
and U13923 (N_13923,N_13698,N_13520);
and U13924 (N_13924,N_13725,N_13666);
xnor U13925 (N_13925,N_13709,N_13567);
nand U13926 (N_13926,N_13571,N_13537);
and U13927 (N_13927,N_13536,N_13609);
nand U13928 (N_13928,N_13544,N_13519);
and U13929 (N_13929,N_13539,N_13689);
nor U13930 (N_13930,N_13558,N_13580);
nand U13931 (N_13931,N_13675,N_13516);
or U13932 (N_13932,N_13661,N_13684);
and U13933 (N_13933,N_13514,N_13640);
nand U13934 (N_13934,N_13579,N_13604);
or U13935 (N_13935,N_13531,N_13629);
xnor U13936 (N_13936,N_13674,N_13737);
xnor U13937 (N_13937,N_13707,N_13733);
nand U13938 (N_13938,N_13736,N_13653);
nor U13939 (N_13939,N_13647,N_13548);
or U13940 (N_13940,N_13620,N_13730);
or U13941 (N_13941,N_13606,N_13713);
xnor U13942 (N_13942,N_13628,N_13739);
or U13943 (N_13943,N_13701,N_13748);
or U13944 (N_13944,N_13665,N_13602);
nand U13945 (N_13945,N_13651,N_13578);
or U13946 (N_13946,N_13683,N_13519);
xor U13947 (N_13947,N_13604,N_13670);
or U13948 (N_13948,N_13573,N_13740);
nor U13949 (N_13949,N_13616,N_13748);
nor U13950 (N_13950,N_13695,N_13653);
nand U13951 (N_13951,N_13631,N_13651);
nand U13952 (N_13952,N_13592,N_13627);
nand U13953 (N_13953,N_13691,N_13538);
and U13954 (N_13954,N_13539,N_13645);
xor U13955 (N_13955,N_13701,N_13519);
or U13956 (N_13956,N_13692,N_13658);
and U13957 (N_13957,N_13516,N_13520);
nor U13958 (N_13958,N_13546,N_13667);
or U13959 (N_13959,N_13559,N_13518);
nor U13960 (N_13960,N_13663,N_13509);
nand U13961 (N_13961,N_13536,N_13565);
xor U13962 (N_13962,N_13686,N_13628);
xor U13963 (N_13963,N_13625,N_13571);
or U13964 (N_13964,N_13731,N_13748);
and U13965 (N_13965,N_13637,N_13728);
xnor U13966 (N_13966,N_13649,N_13542);
nor U13967 (N_13967,N_13746,N_13660);
nand U13968 (N_13968,N_13667,N_13701);
nand U13969 (N_13969,N_13505,N_13713);
xnor U13970 (N_13970,N_13704,N_13559);
and U13971 (N_13971,N_13549,N_13616);
xnor U13972 (N_13972,N_13502,N_13696);
nand U13973 (N_13973,N_13505,N_13649);
nand U13974 (N_13974,N_13541,N_13519);
or U13975 (N_13975,N_13642,N_13736);
nor U13976 (N_13976,N_13502,N_13718);
or U13977 (N_13977,N_13681,N_13591);
nor U13978 (N_13978,N_13746,N_13628);
or U13979 (N_13979,N_13508,N_13743);
nand U13980 (N_13980,N_13626,N_13656);
nor U13981 (N_13981,N_13555,N_13690);
or U13982 (N_13982,N_13500,N_13501);
xnor U13983 (N_13983,N_13733,N_13734);
and U13984 (N_13984,N_13531,N_13551);
nand U13985 (N_13985,N_13693,N_13640);
xor U13986 (N_13986,N_13513,N_13696);
or U13987 (N_13987,N_13595,N_13655);
and U13988 (N_13988,N_13676,N_13575);
or U13989 (N_13989,N_13521,N_13606);
nor U13990 (N_13990,N_13740,N_13741);
nand U13991 (N_13991,N_13568,N_13668);
nand U13992 (N_13992,N_13517,N_13620);
or U13993 (N_13993,N_13669,N_13533);
nor U13994 (N_13994,N_13554,N_13690);
or U13995 (N_13995,N_13536,N_13733);
or U13996 (N_13996,N_13677,N_13573);
nand U13997 (N_13997,N_13661,N_13697);
nand U13998 (N_13998,N_13552,N_13546);
or U13999 (N_13999,N_13746,N_13722);
and U14000 (N_14000,N_13908,N_13922);
nor U14001 (N_14001,N_13881,N_13931);
nand U14002 (N_14002,N_13975,N_13890);
or U14003 (N_14003,N_13869,N_13898);
xnor U14004 (N_14004,N_13929,N_13937);
nor U14005 (N_14005,N_13820,N_13767);
nand U14006 (N_14006,N_13834,N_13813);
nand U14007 (N_14007,N_13943,N_13879);
nor U14008 (N_14008,N_13936,N_13807);
nand U14009 (N_14009,N_13829,N_13946);
and U14010 (N_14010,N_13885,N_13839);
or U14011 (N_14011,N_13751,N_13785);
and U14012 (N_14012,N_13873,N_13967);
and U14013 (N_14013,N_13808,N_13769);
xnor U14014 (N_14014,N_13985,N_13948);
and U14015 (N_14015,N_13994,N_13880);
nand U14016 (N_14016,N_13914,N_13989);
and U14017 (N_14017,N_13801,N_13832);
nor U14018 (N_14018,N_13805,N_13852);
nand U14019 (N_14019,N_13945,N_13845);
or U14020 (N_14020,N_13979,N_13770);
and U14021 (N_14021,N_13900,N_13958);
nand U14022 (N_14022,N_13878,N_13983);
or U14023 (N_14023,N_13786,N_13778);
nand U14024 (N_14024,N_13783,N_13949);
nand U14025 (N_14025,N_13806,N_13874);
or U14026 (N_14026,N_13951,N_13865);
xnor U14027 (N_14027,N_13823,N_13753);
xnor U14028 (N_14028,N_13906,N_13836);
or U14029 (N_14029,N_13954,N_13850);
xor U14030 (N_14030,N_13831,N_13991);
or U14031 (N_14031,N_13952,N_13755);
xor U14032 (N_14032,N_13856,N_13893);
and U14033 (N_14033,N_13780,N_13844);
and U14034 (N_14034,N_13827,N_13837);
or U14035 (N_14035,N_13897,N_13795);
nor U14036 (N_14036,N_13848,N_13966);
and U14037 (N_14037,N_13911,N_13761);
nand U14038 (N_14038,N_13798,N_13833);
xnor U14039 (N_14039,N_13970,N_13814);
xor U14040 (N_14040,N_13884,N_13886);
nor U14041 (N_14041,N_13877,N_13972);
nor U14042 (N_14042,N_13899,N_13875);
or U14043 (N_14043,N_13861,N_13842);
nor U14044 (N_14044,N_13920,N_13982);
nand U14045 (N_14045,N_13782,N_13830);
or U14046 (N_14046,N_13773,N_13800);
xor U14047 (N_14047,N_13959,N_13819);
nor U14048 (N_14048,N_13796,N_13903);
or U14049 (N_14049,N_13888,N_13926);
nand U14050 (N_14050,N_13964,N_13940);
or U14051 (N_14051,N_13758,N_13938);
and U14052 (N_14052,N_13928,N_13997);
nor U14053 (N_14053,N_13930,N_13826);
nor U14054 (N_14054,N_13953,N_13913);
xor U14055 (N_14055,N_13788,N_13968);
or U14056 (N_14056,N_13777,N_13846);
or U14057 (N_14057,N_13891,N_13978);
or U14058 (N_14058,N_13784,N_13990);
or U14059 (N_14059,N_13939,N_13812);
nand U14060 (N_14060,N_13871,N_13981);
nand U14061 (N_14061,N_13776,N_13762);
xnor U14062 (N_14062,N_13955,N_13824);
nand U14063 (N_14063,N_13901,N_13759);
nand U14064 (N_14064,N_13774,N_13915);
xnor U14065 (N_14065,N_13904,N_13754);
or U14066 (N_14066,N_13793,N_13750);
nand U14067 (N_14067,N_13858,N_13804);
xor U14068 (N_14068,N_13916,N_13987);
nand U14069 (N_14069,N_13789,N_13912);
nand U14070 (N_14070,N_13960,N_13924);
nor U14071 (N_14071,N_13870,N_13811);
and U14072 (N_14072,N_13976,N_13772);
and U14073 (N_14073,N_13941,N_13797);
xnor U14074 (N_14074,N_13999,N_13752);
or U14075 (N_14075,N_13794,N_13971);
and U14076 (N_14076,N_13992,N_13935);
xnor U14077 (N_14077,N_13894,N_13969);
nor U14078 (N_14078,N_13757,N_13822);
nor U14079 (N_14079,N_13816,N_13917);
nand U14080 (N_14080,N_13872,N_13840);
or U14081 (N_14081,N_13925,N_13995);
nor U14082 (N_14082,N_13843,N_13957);
xnor U14083 (N_14083,N_13876,N_13760);
nand U14084 (N_14084,N_13864,N_13933);
nor U14085 (N_14085,N_13756,N_13895);
xor U14086 (N_14086,N_13923,N_13835);
xor U14087 (N_14087,N_13947,N_13919);
xnor U14088 (N_14088,N_13866,N_13818);
xnor U14089 (N_14089,N_13825,N_13809);
xnor U14090 (N_14090,N_13984,N_13921);
or U14091 (N_14091,N_13907,N_13766);
or U14092 (N_14092,N_13765,N_13855);
nor U14093 (N_14093,N_13902,N_13918);
nand U14094 (N_14094,N_13892,N_13942);
or U14095 (N_14095,N_13905,N_13847);
nor U14096 (N_14096,N_13781,N_13956);
xnor U14097 (N_14097,N_13973,N_13998);
nand U14098 (N_14098,N_13787,N_13962);
or U14099 (N_14099,N_13934,N_13857);
xor U14100 (N_14100,N_13867,N_13779);
or U14101 (N_14101,N_13932,N_13851);
nand U14102 (N_14102,N_13790,N_13927);
and U14103 (N_14103,N_13996,N_13909);
xnor U14104 (N_14104,N_13803,N_13849);
nor U14105 (N_14105,N_13817,N_13988);
xor U14106 (N_14106,N_13792,N_13815);
xnor U14107 (N_14107,N_13859,N_13802);
nor U14108 (N_14108,N_13883,N_13896);
and U14109 (N_14109,N_13810,N_13974);
xnor U14110 (N_14110,N_13841,N_13882);
xor U14111 (N_14111,N_13853,N_13910);
nand U14112 (N_14112,N_13961,N_13977);
xor U14113 (N_14113,N_13821,N_13854);
and U14114 (N_14114,N_13887,N_13799);
or U14115 (N_14115,N_13791,N_13889);
xnor U14116 (N_14116,N_13993,N_13838);
xor U14117 (N_14117,N_13862,N_13764);
xnor U14118 (N_14118,N_13860,N_13828);
and U14119 (N_14119,N_13965,N_13771);
and U14120 (N_14120,N_13963,N_13863);
and U14121 (N_14121,N_13868,N_13950);
or U14122 (N_14122,N_13775,N_13768);
nand U14123 (N_14123,N_13986,N_13944);
nor U14124 (N_14124,N_13980,N_13763);
xor U14125 (N_14125,N_13897,N_13907);
xor U14126 (N_14126,N_13780,N_13896);
nand U14127 (N_14127,N_13847,N_13806);
or U14128 (N_14128,N_13954,N_13894);
or U14129 (N_14129,N_13759,N_13842);
or U14130 (N_14130,N_13862,N_13813);
nor U14131 (N_14131,N_13962,N_13833);
nand U14132 (N_14132,N_13867,N_13876);
nand U14133 (N_14133,N_13809,N_13900);
nor U14134 (N_14134,N_13873,N_13775);
and U14135 (N_14135,N_13838,N_13758);
or U14136 (N_14136,N_13872,N_13878);
xor U14137 (N_14137,N_13805,N_13813);
and U14138 (N_14138,N_13991,N_13964);
nor U14139 (N_14139,N_13803,N_13862);
and U14140 (N_14140,N_13793,N_13897);
nand U14141 (N_14141,N_13946,N_13922);
or U14142 (N_14142,N_13942,N_13846);
nand U14143 (N_14143,N_13852,N_13991);
xnor U14144 (N_14144,N_13916,N_13798);
or U14145 (N_14145,N_13897,N_13997);
and U14146 (N_14146,N_13789,N_13959);
nand U14147 (N_14147,N_13956,N_13780);
or U14148 (N_14148,N_13878,N_13978);
xnor U14149 (N_14149,N_13962,N_13859);
nor U14150 (N_14150,N_13775,N_13798);
xor U14151 (N_14151,N_13903,N_13939);
xor U14152 (N_14152,N_13800,N_13867);
xor U14153 (N_14153,N_13846,N_13758);
nor U14154 (N_14154,N_13908,N_13791);
and U14155 (N_14155,N_13898,N_13877);
or U14156 (N_14156,N_13775,N_13913);
or U14157 (N_14157,N_13895,N_13854);
nor U14158 (N_14158,N_13796,N_13941);
nor U14159 (N_14159,N_13928,N_13898);
nor U14160 (N_14160,N_13873,N_13914);
and U14161 (N_14161,N_13780,N_13807);
xnor U14162 (N_14162,N_13764,N_13754);
nor U14163 (N_14163,N_13915,N_13842);
xor U14164 (N_14164,N_13840,N_13764);
nor U14165 (N_14165,N_13987,N_13800);
nor U14166 (N_14166,N_13802,N_13969);
nand U14167 (N_14167,N_13839,N_13783);
xnor U14168 (N_14168,N_13894,N_13807);
xnor U14169 (N_14169,N_13950,N_13813);
nand U14170 (N_14170,N_13799,N_13983);
nor U14171 (N_14171,N_13963,N_13846);
nand U14172 (N_14172,N_13929,N_13998);
and U14173 (N_14173,N_13941,N_13863);
or U14174 (N_14174,N_13869,N_13965);
xnor U14175 (N_14175,N_13812,N_13799);
xnor U14176 (N_14176,N_13865,N_13919);
or U14177 (N_14177,N_13775,N_13751);
or U14178 (N_14178,N_13860,N_13919);
nand U14179 (N_14179,N_13830,N_13971);
or U14180 (N_14180,N_13809,N_13818);
or U14181 (N_14181,N_13806,N_13989);
or U14182 (N_14182,N_13926,N_13840);
xnor U14183 (N_14183,N_13979,N_13938);
nor U14184 (N_14184,N_13942,N_13920);
and U14185 (N_14185,N_13862,N_13913);
and U14186 (N_14186,N_13775,N_13792);
or U14187 (N_14187,N_13845,N_13819);
or U14188 (N_14188,N_13906,N_13947);
xor U14189 (N_14189,N_13933,N_13940);
xnor U14190 (N_14190,N_13857,N_13919);
nor U14191 (N_14191,N_13883,N_13964);
nor U14192 (N_14192,N_13964,N_13989);
xor U14193 (N_14193,N_13826,N_13822);
xor U14194 (N_14194,N_13813,N_13767);
or U14195 (N_14195,N_13995,N_13808);
nand U14196 (N_14196,N_13941,N_13756);
nand U14197 (N_14197,N_13869,N_13803);
nor U14198 (N_14198,N_13933,N_13822);
nor U14199 (N_14199,N_13769,N_13939);
and U14200 (N_14200,N_13778,N_13884);
nor U14201 (N_14201,N_13827,N_13852);
nor U14202 (N_14202,N_13757,N_13884);
or U14203 (N_14203,N_13876,N_13892);
and U14204 (N_14204,N_13799,N_13809);
nand U14205 (N_14205,N_13831,N_13880);
nand U14206 (N_14206,N_13760,N_13958);
and U14207 (N_14207,N_13771,N_13984);
nor U14208 (N_14208,N_13988,N_13888);
xor U14209 (N_14209,N_13839,N_13832);
xor U14210 (N_14210,N_13913,N_13848);
and U14211 (N_14211,N_13989,N_13917);
or U14212 (N_14212,N_13930,N_13993);
nand U14213 (N_14213,N_13758,N_13890);
xnor U14214 (N_14214,N_13853,N_13866);
nor U14215 (N_14215,N_13788,N_13825);
nand U14216 (N_14216,N_13761,N_13997);
xnor U14217 (N_14217,N_13820,N_13907);
or U14218 (N_14218,N_13817,N_13931);
or U14219 (N_14219,N_13843,N_13962);
nor U14220 (N_14220,N_13813,N_13777);
xnor U14221 (N_14221,N_13830,N_13882);
xnor U14222 (N_14222,N_13868,N_13807);
nand U14223 (N_14223,N_13792,N_13993);
nand U14224 (N_14224,N_13919,N_13872);
nor U14225 (N_14225,N_13945,N_13879);
and U14226 (N_14226,N_13947,N_13918);
and U14227 (N_14227,N_13863,N_13968);
xor U14228 (N_14228,N_13816,N_13878);
and U14229 (N_14229,N_13752,N_13806);
xor U14230 (N_14230,N_13982,N_13790);
or U14231 (N_14231,N_13784,N_13903);
nand U14232 (N_14232,N_13999,N_13802);
nor U14233 (N_14233,N_13995,N_13755);
nor U14234 (N_14234,N_13853,N_13861);
and U14235 (N_14235,N_13946,N_13927);
nor U14236 (N_14236,N_13945,N_13870);
or U14237 (N_14237,N_13883,N_13933);
nor U14238 (N_14238,N_13934,N_13996);
and U14239 (N_14239,N_13785,N_13951);
xnor U14240 (N_14240,N_13967,N_13780);
or U14241 (N_14241,N_13874,N_13921);
xor U14242 (N_14242,N_13963,N_13898);
or U14243 (N_14243,N_13836,N_13919);
nor U14244 (N_14244,N_13994,N_13764);
nor U14245 (N_14245,N_13988,N_13800);
xnor U14246 (N_14246,N_13909,N_13751);
nor U14247 (N_14247,N_13830,N_13844);
and U14248 (N_14248,N_13874,N_13988);
xor U14249 (N_14249,N_13879,N_13794);
nand U14250 (N_14250,N_14188,N_14026);
or U14251 (N_14251,N_14016,N_14249);
and U14252 (N_14252,N_14152,N_14178);
or U14253 (N_14253,N_14171,N_14110);
nand U14254 (N_14254,N_14069,N_14047);
nor U14255 (N_14255,N_14079,N_14133);
and U14256 (N_14256,N_14019,N_14107);
nand U14257 (N_14257,N_14063,N_14183);
and U14258 (N_14258,N_14229,N_14052);
nor U14259 (N_14259,N_14168,N_14078);
xnor U14260 (N_14260,N_14066,N_14111);
nor U14261 (N_14261,N_14137,N_14029);
nor U14262 (N_14262,N_14220,N_14008);
xor U14263 (N_14263,N_14000,N_14185);
nor U14264 (N_14264,N_14020,N_14238);
and U14265 (N_14265,N_14085,N_14009);
nor U14266 (N_14266,N_14046,N_14245);
nor U14267 (N_14267,N_14094,N_14037);
nor U14268 (N_14268,N_14098,N_14215);
xnor U14269 (N_14269,N_14032,N_14126);
nor U14270 (N_14270,N_14140,N_14148);
and U14271 (N_14271,N_14053,N_14170);
xnor U14272 (N_14272,N_14217,N_14210);
nand U14273 (N_14273,N_14073,N_14011);
or U14274 (N_14274,N_14236,N_14247);
and U14275 (N_14275,N_14030,N_14181);
and U14276 (N_14276,N_14114,N_14156);
and U14277 (N_14277,N_14169,N_14061);
or U14278 (N_14278,N_14102,N_14106);
or U14279 (N_14279,N_14092,N_14246);
nand U14280 (N_14280,N_14097,N_14088);
nand U14281 (N_14281,N_14205,N_14175);
xor U14282 (N_14282,N_14162,N_14112);
nand U14283 (N_14283,N_14243,N_14043);
nand U14284 (N_14284,N_14232,N_14196);
or U14285 (N_14285,N_14151,N_14059);
or U14286 (N_14286,N_14143,N_14223);
or U14287 (N_14287,N_14074,N_14248);
nand U14288 (N_14288,N_14024,N_14237);
or U14289 (N_14289,N_14153,N_14145);
or U14290 (N_14290,N_14113,N_14040);
nor U14291 (N_14291,N_14087,N_14072);
xnor U14292 (N_14292,N_14154,N_14028);
nor U14293 (N_14293,N_14214,N_14197);
nor U14294 (N_14294,N_14051,N_14136);
and U14295 (N_14295,N_14182,N_14184);
nor U14296 (N_14296,N_14057,N_14002);
nand U14297 (N_14297,N_14076,N_14075);
and U14298 (N_14298,N_14099,N_14095);
nor U14299 (N_14299,N_14129,N_14005);
or U14300 (N_14300,N_14058,N_14209);
nand U14301 (N_14301,N_14022,N_14155);
nor U14302 (N_14302,N_14045,N_14070);
nor U14303 (N_14303,N_14015,N_14064);
and U14304 (N_14304,N_14100,N_14163);
or U14305 (N_14305,N_14165,N_14118);
xor U14306 (N_14306,N_14242,N_14234);
nor U14307 (N_14307,N_14125,N_14180);
nand U14308 (N_14308,N_14139,N_14123);
nor U14309 (N_14309,N_14160,N_14159);
xnor U14310 (N_14310,N_14093,N_14115);
and U14311 (N_14311,N_14201,N_14212);
and U14312 (N_14312,N_14012,N_14167);
and U14313 (N_14313,N_14189,N_14124);
nor U14314 (N_14314,N_14239,N_14080);
nand U14315 (N_14315,N_14056,N_14240);
xnor U14316 (N_14316,N_14142,N_14204);
and U14317 (N_14317,N_14135,N_14222);
and U14318 (N_14318,N_14207,N_14067);
nor U14319 (N_14319,N_14001,N_14233);
nor U14320 (N_14320,N_14035,N_14027);
nand U14321 (N_14321,N_14105,N_14108);
xnor U14322 (N_14322,N_14157,N_14041);
xor U14323 (N_14323,N_14213,N_14049);
nor U14324 (N_14324,N_14089,N_14174);
or U14325 (N_14325,N_14219,N_14090);
and U14326 (N_14326,N_14241,N_14187);
nand U14327 (N_14327,N_14050,N_14228);
xnor U14328 (N_14328,N_14193,N_14176);
xnor U14329 (N_14329,N_14144,N_14039);
nor U14330 (N_14330,N_14007,N_14065);
and U14331 (N_14331,N_14173,N_14186);
nor U14332 (N_14332,N_14091,N_14060);
nor U14333 (N_14333,N_14226,N_14131);
nor U14334 (N_14334,N_14084,N_14013);
and U14335 (N_14335,N_14224,N_14235);
xnor U14336 (N_14336,N_14161,N_14218);
xnor U14337 (N_14337,N_14231,N_14014);
and U14338 (N_14338,N_14048,N_14116);
nand U14339 (N_14339,N_14190,N_14192);
xnor U14340 (N_14340,N_14221,N_14179);
and U14341 (N_14341,N_14244,N_14120);
nand U14342 (N_14342,N_14134,N_14195);
nor U14343 (N_14343,N_14062,N_14119);
and U14344 (N_14344,N_14054,N_14147);
and U14345 (N_14345,N_14031,N_14006);
nand U14346 (N_14346,N_14004,N_14225);
xnor U14347 (N_14347,N_14191,N_14121);
or U14348 (N_14348,N_14141,N_14122);
or U14349 (N_14349,N_14227,N_14103);
nand U14350 (N_14350,N_14166,N_14202);
nand U14351 (N_14351,N_14082,N_14172);
nor U14352 (N_14352,N_14018,N_14164);
or U14353 (N_14353,N_14200,N_14194);
and U14354 (N_14354,N_14206,N_14127);
nand U14355 (N_14355,N_14128,N_14077);
nor U14356 (N_14356,N_14042,N_14044);
nand U14357 (N_14357,N_14150,N_14081);
nand U14358 (N_14358,N_14034,N_14211);
xor U14359 (N_14359,N_14132,N_14096);
xor U14360 (N_14360,N_14104,N_14208);
nor U14361 (N_14361,N_14068,N_14216);
nor U14362 (N_14362,N_14117,N_14033);
xnor U14363 (N_14363,N_14177,N_14017);
and U14364 (N_14364,N_14158,N_14138);
nor U14365 (N_14365,N_14038,N_14199);
nor U14366 (N_14366,N_14198,N_14149);
nand U14367 (N_14367,N_14010,N_14083);
and U14368 (N_14368,N_14101,N_14025);
nand U14369 (N_14369,N_14036,N_14230);
and U14370 (N_14370,N_14055,N_14003);
and U14371 (N_14371,N_14021,N_14146);
xnor U14372 (N_14372,N_14071,N_14086);
and U14373 (N_14373,N_14023,N_14203);
and U14374 (N_14374,N_14130,N_14109);
or U14375 (N_14375,N_14151,N_14164);
nor U14376 (N_14376,N_14198,N_14231);
nor U14377 (N_14377,N_14021,N_14076);
nor U14378 (N_14378,N_14243,N_14132);
and U14379 (N_14379,N_14129,N_14041);
nand U14380 (N_14380,N_14152,N_14213);
or U14381 (N_14381,N_14026,N_14162);
and U14382 (N_14382,N_14001,N_14148);
nand U14383 (N_14383,N_14197,N_14137);
nor U14384 (N_14384,N_14002,N_14200);
nor U14385 (N_14385,N_14007,N_14203);
and U14386 (N_14386,N_14054,N_14083);
nand U14387 (N_14387,N_14027,N_14179);
nand U14388 (N_14388,N_14243,N_14048);
xnor U14389 (N_14389,N_14045,N_14148);
nand U14390 (N_14390,N_14002,N_14146);
xor U14391 (N_14391,N_14030,N_14056);
and U14392 (N_14392,N_14108,N_14063);
or U14393 (N_14393,N_14019,N_14176);
xnor U14394 (N_14394,N_14055,N_14168);
nand U14395 (N_14395,N_14248,N_14055);
nand U14396 (N_14396,N_14122,N_14161);
xnor U14397 (N_14397,N_14222,N_14009);
and U14398 (N_14398,N_14170,N_14095);
or U14399 (N_14399,N_14150,N_14063);
and U14400 (N_14400,N_14015,N_14103);
and U14401 (N_14401,N_14149,N_14185);
and U14402 (N_14402,N_14068,N_14171);
and U14403 (N_14403,N_14135,N_14133);
nor U14404 (N_14404,N_14151,N_14008);
xnor U14405 (N_14405,N_14210,N_14085);
nand U14406 (N_14406,N_14109,N_14131);
or U14407 (N_14407,N_14209,N_14000);
and U14408 (N_14408,N_14091,N_14195);
or U14409 (N_14409,N_14030,N_14157);
or U14410 (N_14410,N_14038,N_14212);
nand U14411 (N_14411,N_14002,N_14053);
nor U14412 (N_14412,N_14003,N_14222);
nor U14413 (N_14413,N_14110,N_14243);
nor U14414 (N_14414,N_14220,N_14230);
nand U14415 (N_14415,N_14113,N_14056);
or U14416 (N_14416,N_14010,N_14098);
or U14417 (N_14417,N_14094,N_14160);
nor U14418 (N_14418,N_14041,N_14245);
nand U14419 (N_14419,N_14133,N_14234);
xnor U14420 (N_14420,N_14012,N_14149);
or U14421 (N_14421,N_14102,N_14146);
and U14422 (N_14422,N_14247,N_14107);
and U14423 (N_14423,N_14212,N_14156);
nand U14424 (N_14424,N_14172,N_14094);
nor U14425 (N_14425,N_14175,N_14077);
xnor U14426 (N_14426,N_14088,N_14144);
and U14427 (N_14427,N_14171,N_14148);
nand U14428 (N_14428,N_14226,N_14056);
nor U14429 (N_14429,N_14200,N_14126);
nand U14430 (N_14430,N_14247,N_14132);
nand U14431 (N_14431,N_14077,N_14232);
xnor U14432 (N_14432,N_14133,N_14030);
and U14433 (N_14433,N_14038,N_14125);
nor U14434 (N_14434,N_14227,N_14135);
and U14435 (N_14435,N_14210,N_14019);
nand U14436 (N_14436,N_14093,N_14100);
or U14437 (N_14437,N_14240,N_14047);
nand U14438 (N_14438,N_14044,N_14015);
nand U14439 (N_14439,N_14237,N_14159);
or U14440 (N_14440,N_14215,N_14042);
or U14441 (N_14441,N_14063,N_14092);
and U14442 (N_14442,N_14037,N_14188);
nor U14443 (N_14443,N_14241,N_14054);
or U14444 (N_14444,N_14047,N_14230);
or U14445 (N_14445,N_14206,N_14094);
nor U14446 (N_14446,N_14074,N_14048);
or U14447 (N_14447,N_14044,N_14032);
nand U14448 (N_14448,N_14242,N_14001);
or U14449 (N_14449,N_14225,N_14150);
or U14450 (N_14450,N_14244,N_14027);
nor U14451 (N_14451,N_14135,N_14024);
or U14452 (N_14452,N_14211,N_14100);
xnor U14453 (N_14453,N_14021,N_14150);
or U14454 (N_14454,N_14205,N_14090);
nand U14455 (N_14455,N_14219,N_14151);
or U14456 (N_14456,N_14196,N_14040);
xnor U14457 (N_14457,N_14195,N_14114);
xnor U14458 (N_14458,N_14147,N_14117);
nand U14459 (N_14459,N_14237,N_14037);
nor U14460 (N_14460,N_14090,N_14228);
or U14461 (N_14461,N_14154,N_14214);
nand U14462 (N_14462,N_14053,N_14142);
xor U14463 (N_14463,N_14180,N_14153);
nand U14464 (N_14464,N_14061,N_14000);
and U14465 (N_14465,N_14118,N_14014);
and U14466 (N_14466,N_14174,N_14211);
xor U14467 (N_14467,N_14045,N_14223);
nor U14468 (N_14468,N_14030,N_14110);
xor U14469 (N_14469,N_14036,N_14076);
nand U14470 (N_14470,N_14091,N_14037);
or U14471 (N_14471,N_14103,N_14235);
xor U14472 (N_14472,N_14175,N_14009);
nor U14473 (N_14473,N_14241,N_14068);
nand U14474 (N_14474,N_14154,N_14113);
and U14475 (N_14475,N_14049,N_14011);
and U14476 (N_14476,N_14194,N_14000);
and U14477 (N_14477,N_14147,N_14030);
and U14478 (N_14478,N_14009,N_14131);
xor U14479 (N_14479,N_14047,N_14049);
nand U14480 (N_14480,N_14066,N_14009);
and U14481 (N_14481,N_14244,N_14159);
nor U14482 (N_14482,N_14103,N_14091);
or U14483 (N_14483,N_14213,N_14052);
nand U14484 (N_14484,N_14173,N_14063);
xnor U14485 (N_14485,N_14235,N_14069);
and U14486 (N_14486,N_14202,N_14122);
or U14487 (N_14487,N_14197,N_14210);
and U14488 (N_14488,N_14059,N_14026);
nand U14489 (N_14489,N_14165,N_14120);
nand U14490 (N_14490,N_14093,N_14057);
and U14491 (N_14491,N_14046,N_14052);
nor U14492 (N_14492,N_14081,N_14169);
nand U14493 (N_14493,N_14244,N_14102);
and U14494 (N_14494,N_14096,N_14027);
nand U14495 (N_14495,N_14126,N_14013);
or U14496 (N_14496,N_14132,N_14218);
nand U14497 (N_14497,N_14130,N_14148);
nand U14498 (N_14498,N_14074,N_14159);
and U14499 (N_14499,N_14000,N_14227);
and U14500 (N_14500,N_14441,N_14263);
or U14501 (N_14501,N_14336,N_14477);
nand U14502 (N_14502,N_14476,N_14385);
or U14503 (N_14503,N_14322,N_14352);
or U14504 (N_14504,N_14338,N_14365);
xnor U14505 (N_14505,N_14303,N_14301);
nor U14506 (N_14506,N_14399,N_14341);
nor U14507 (N_14507,N_14425,N_14382);
or U14508 (N_14508,N_14280,N_14410);
or U14509 (N_14509,N_14393,N_14475);
or U14510 (N_14510,N_14487,N_14418);
xnor U14511 (N_14511,N_14268,N_14276);
nand U14512 (N_14512,N_14455,N_14428);
xor U14513 (N_14513,N_14386,N_14287);
nor U14514 (N_14514,N_14277,N_14423);
xnor U14515 (N_14515,N_14494,N_14383);
nor U14516 (N_14516,N_14306,N_14465);
nand U14517 (N_14517,N_14327,N_14286);
nand U14518 (N_14518,N_14316,N_14409);
nand U14519 (N_14519,N_14359,N_14252);
and U14520 (N_14520,N_14310,N_14373);
nor U14521 (N_14521,N_14363,N_14495);
or U14522 (N_14522,N_14312,N_14361);
or U14523 (N_14523,N_14463,N_14388);
xor U14524 (N_14524,N_14490,N_14362);
xnor U14525 (N_14525,N_14379,N_14292);
nor U14526 (N_14526,N_14479,N_14358);
and U14527 (N_14527,N_14319,N_14456);
nand U14528 (N_14528,N_14294,N_14346);
or U14529 (N_14529,N_14339,N_14491);
xnor U14530 (N_14530,N_14360,N_14289);
and U14531 (N_14531,N_14275,N_14253);
nand U14532 (N_14532,N_14272,N_14305);
xnor U14533 (N_14533,N_14329,N_14406);
nand U14534 (N_14534,N_14401,N_14480);
nor U14535 (N_14535,N_14485,N_14427);
nand U14536 (N_14536,N_14351,N_14282);
and U14537 (N_14537,N_14438,N_14394);
nor U14538 (N_14538,N_14278,N_14343);
or U14539 (N_14539,N_14326,N_14446);
xor U14540 (N_14540,N_14376,N_14364);
and U14541 (N_14541,N_14396,N_14387);
or U14542 (N_14542,N_14370,N_14309);
nor U14543 (N_14543,N_14481,N_14260);
and U14544 (N_14544,N_14274,N_14342);
or U14545 (N_14545,N_14350,N_14473);
xnor U14546 (N_14546,N_14251,N_14458);
and U14547 (N_14547,N_14355,N_14429);
or U14548 (N_14548,N_14417,N_14345);
nand U14549 (N_14549,N_14408,N_14405);
nor U14550 (N_14550,N_14390,N_14493);
and U14551 (N_14551,N_14496,N_14380);
nand U14552 (N_14552,N_14354,N_14432);
and U14553 (N_14553,N_14255,N_14332);
xnor U14554 (N_14554,N_14257,N_14313);
nand U14555 (N_14555,N_14483,N_14435);
or U14556 (N_14556,N_14412,N_14497);
or U14557 (N_14557,N_14330,N_14334);
nand U14558 (N_14558,N_14457,N_14357);
nor U14559 (N_14559,N_14482,N_14397);
nand U14560 (N_14560,N_14295,N_14353);
xor U14561 (N_14561,N_14281,N_14430);
xnor U14562 (N_14562,N_14299,N_14344);
nor U14563 (N_14563,N_14377,N_14348);
xor U14564 (N_14564,N_14470,N_14250);
nand U14565 (N_14565,N_14411,N_14265);
nor U14566 (N_14566,N_14356,N_14266);
nor U14567 (N_14567,N_14462,N_14381);
nor U14568 (N_14568,N_14279,N_14384);
and U14569 (N_14569,N_14499,N_14311);
xor U14570 (N_14570,N_14447,N_14413);
or U14571 (N_14571,N_14421,N_14283);
xnor U14572 (N_14572,N_14367,N_14261);
or U14573 (N_14573,N_14267,N_14460);
or U14574 (N_14574,N_14271,N_14290);
nor U14575 (N_14575,N_14403,N_14372);
nor U14576 (N_14576,N_14454,N_14471);
nor U14577 (N_14577,N_14461,N_14415);
nor U14578 (N_14578,N_14439,N_14371);
xnor U14579 (N_14579,N_14437,N_14416);
and U14580 (N_14580,N_14469,N_14426);
xnor U14581 (N_14581,N_14366,N_14315);
nor U14582 (N_14582,N_14442,N_14314);
xor U14583 (N_14583,N_14450,N_14395);
xnor U14584 (N_14584,N_14424,N_14374);
nand U14585 (N_14585,N_14273,N_14431);
nand U14586 (N_14586,N_14349,N_14307);
and U14587 (N_14587,N_14404,N_14414);
nor U14588 (N_14588,N_14308,N_14324);
and U14589 (N_14589,N_14402,N_14448);
or U14590 (N_14590,N_14256,N_14440);
and U14591 (N_14591,N_14284,N_14340);
or U14592 (N_14592,N_14443,N_14368);
xnor U14593 (N_14593,N_14269,N_14453);
nor U14594 (N_14594,N_14258,N_14391);
and U14595 (N_14595,N_14347,N_14297);
or U14596 (N_14596,N_14304,N_14419);
nor U14597 (N_14597,N_14398,N_14320);
xnor U14598 (N_14598,N_14466,N_14262);
xnor U14599 (N_14599,N_14293,N_14492);
xnor U14600 (N_14600,N_14392,N_14331);
nor U14601 (N_14601,N_14467,N_14288);
nand U14602 (N_14602,N_14434,N_14254);
nand U14603 (N_14603,N_14296,N_14468);
nor U14604 (N_14604,N_14337,N_14464);
nor U14605 (N_14605,N_14422,N_14451);
nand U14606 (N_14606,N_14478,N_14335);
or U14607 (N_14607,N_14389,N_14472);
and U14608 (N_14608,N_14333,N_14484);
nand U14609 (N_14609,N_14318,N_14400);
nand U14610 (N_14610,N_14270,N_14285);
or U14611 (N_14611,N_14328,N_14444);
nor U14612 (N_14612,N_14452,N_14300);
nor U14613 (N_14613,N_14321,N_14291);
nor U14614 (N_14614,N_14498,N_14459);
nand U14615 (N_14615,N_14407,N_14488);
nor U14616 (N_14616,N_14445,N_14436);
nor U14617 (N_14617,N_14317,N_14264);
nor U14618 (N_14618,N_14378,N_14259);
nor U14619 (N_14619,N_14302,N_14489);
and U14620 (N_14620,N_14486,N_14298);
and U14621 (N_14621,N_14420,N_14433);
and U14622 (N_14622,N_14449,N_14325);
or U14623 (N_14623,N_14323,N_14375);
nor U14624 (N_14624,N_14369,N_14474);
nand U14625 (N_14625,N_14476,N_14300);
and U14626 (N_14626,N_14300,N_14496);
xor U14627 (N_14627,N_14416,N_14411);
xor U14628 (N_14628,N_14427,N_14407);
nor U14629 (N_14629,N_14313,N_14435);
and U14630 (N_14630,N_14281,N_14270);
xor U14631 (N_14631,N_14473,N_14417);
nor U14632 (N_14632,N_14422,N_14440);
and U14633 (N_14633,N_14462,N_14423);
nor U14634 (N_14634,N_14487,N_14295);
nor U14635 (N_14635,N_14409,N_14264);
nor U14636 (N_14636,N_14342,N_14376);
xor U14637 (N_14637,N_14467,N_14304);
or U14638 (N_14638,N_14451,N_14337);
nor U14639 (N_14639,N_14370,N_14396);
nor U14640 (N_14640,N_14466,N_14250);
or U14641 (N_14641,N_14301,N_14313);
xnor U14642 (N_14642,N_14390,N_14344);
or U14643 (N_14643,N_14458,N_14274);
nand U14644 (N_14644,N_14429,N_14279);
or U14645 (N_14645,N_14497,N_14258);
xor U14646 (N_14646,N_14254,N_14306);
xor U14647 (N_14647,N_14256,N_14493);
and U14648 (N_14648,N_14268,N_14317);
and U14649 (N_14649,N_14399,N_14363);
xor U14650 (N_14650,N_14427,N_14436);
xor U14651 (N_14651,N_14444,N_14372);
and U14652 (N_14652,N_14412,N_14263);
nor U14653 (N_14653,N_14411,N_14264);
xnor U14654 (N_14654,N_14428,N_14351);
or U14655 (N_14655,N_14365,N_14297);
nor U14656 (N_14656,N_14295,N_14450);
nand U14657 (N_14657,N_14393,N_14367);
xnor U14658 (N_14658,N_14350,N_14421);
or U14659 (N_14659,N_14308,N_14441);
nand U14660 (N_14660,N_14299,N_14279);
and U14661 (N_14661,N_14496,N_14257);
and U14662 (N_14662,N_14490,N_14409);
nor U14663 (N_14663,N_14440,N_14483);
nor U14664 (N_14664,N_14489,N_14332);
nor U14665 (N_14665,N_14341,N_14378);
and U14666 (N_14666,N_14306,N_14480);
nor U14667 (N_14667,N_14313,N_14399);
xnor U14668 (N_14668,N_14337,N_14262);
xnor U14669 (N_14669,N_14342,N_14488);
xnor U14670 (N_14670,N_14379,N_14366);
and U14671 (N_14671,N_14473,N_14283);
or U14672 (N_14672,N_14481,N_14263);
and U14673 (N_14673,N_14441,N_14416);
nand U14674 (N_14674,N_14270,N_14278);
or U14675 (N_14675,N_14448,N_14451);
nand U14676 (N_14676,N_14499,N_14496);
xor U14677 (N_14677,N_14283,N_14324);
nor U14678 (N_14678,N_14483,N_14430);
or U14679 (N_14679,N_14394,N_14273);
xor U14680 (N_14680,N_14284,N_14468);
or U14681 (N_14681,N_14321,N_14351);
or U14682 (N_14682,N_14438,N_14449);
and U14683 (N_14683,N_14330,N_14341);
nand U14684 (N_14684,N_14476,N_14392);
xnor U14685 (N_14685,N_14295,N_14261);
and U14686 (N_14686,N_14338,N_14452);
nand U14687 (N_14687,N_14354,N_14302);
nor U14688 (N_14688,N_14495,N_14324);
nand U14689 (N_14689,N_14278,N_14263);
or U14690 (N_14690,N_14349,N_14449);
xor U14691 (N_14691,N_14438,N_14361);
xnor U14692 (N_14692,N_14312,N_14304);
nand U14693 (N_14693,N_14350,N_14462);
nand U14694 (N_14694,N_14280,N_14268);
nor U14695 (N_14695,N_14377,N_14381);
or U14696 (N_14696,N_14342,N_14418);
nand U14697 (N_14697,N_14442,N_14475);
and U14698 (N_14698,N_14491,N_14318);
or U14699 (N_14699,N_14312,N_14427);
or U14700 (N_14700,N_14412,N_14377);
xor U14701 (N_14701,N_14259,N_14303);
or U14702 (N_14702,N_14467,N_14404);
xnor U14703 (N_14703,N_14469,N_14390);
nor U14704 (N_14704,N_14254,N_14471);
nor U14705 (N_14705,N_14374,N_14259);
xor U14706 (N_14706,N_14378,N_14481);
nand U14707 (N_14707,N_14282,N_14388);
xnor U14708 (N_14708,N_14451,N_14497);
and U14709 (N_14709,N_14348,N_14349);
and U14710 (N_14710,N_14314,N_14255);
nor U14711 (N_14711,N_14302,N_14418);
xnor U14712 (N_14712,N_14302,N_14411);
or U14713 (N_14713,N_14281,N_14488);
nor U14714 (N_14714,N_14391,N_14296);
xnor U14715 (N_14715,N_14478,N_14290);
nor U14716 (N_14716,N_14449,N_14338);
nand U14717 (N_14717,N_14400,N_14448);
xor U14718 (N_14718,N_14466,N_14463);
xnor U14719 (N_14719,N_14417,N_14478);
xor U14720 (N_14720,N_14404,N_14465);
xor U14721 (N_14721,N_14437,N_14342);
nor U14722 (N_14722,N_14360,N_14288);
xor U14723 (N_14723,N_14374,N_14397);
and U14724 (N_14724,N_14294,N_14336);
nor U14725 (N_14725,N_14492,N_14413);
nand U14726 (N_14726,N_14419,N_14273);
xor U14727 (N_14727,N_14434,N_14361);
xnor U14728 (N_14728,N_14374,N_14490);
and U14729 (N_14729,N_14412,N_14447);
xnor U14730 (N_14730,N_14309,N_14349);
and U14731 (N_14731,N_14313,N_14462);
nand U14732 (N_14732,N_14411,N_14391);
or U14733 (N_14733,N_14406,N_14402);
and U14734 (N_14734,N_14491,N_14255);
xnor U14735 (N_14735,N_14416,N_14401);
nand U14736 (N_14736,N_14282,N_14366);
nor U14737 (N_14737,N_14414,N_14282);
and U14738 (N_14738,N_14259,N_14401);
and U14739 (N_14739,N_14263,N_14443);
or U14740 (N_14740,N_14263,N_14350);
nor U14741 (N_14741,N_14495,N_14450);
or U14742 (N_14742,N_14434,N_14380);
nand U14743 (N_14743,N_14332,N_14356);
nand U14744 (N_14744,N_14497,N_14460);
nand U14745 (N_14745,N_14387,N_14358);
nor U14746 (N_14746,N_14405,N_14295);
or U14747 (N_14747,N_14292,N_14353);
and U14748 (N_14748,N_14407,N_14372);
or U14749 (N_14749,N_14287,N_14328);
nand U14750 (N_14750,N_14692,N_14671);
xor U14751 (N_14751,N_14619,N_14522);
xnor U14752 (N_14752,N_14554,N_14676);
xor U14753 (N_14753,N_14540,N_14713);
xor U14754 (N_14754,N_14598,N_14673);
nand U14755 (N_14755,N_14720,N_14573);
or U14756 (N_14756,N_14582,N_14654);
or U14757 (N_14757,N_14506,N_14595);
nand U14758 (N_14758,N_14639,N_14531);
or U14759 (N_14759,N_14605,N_14659);
or U14760 (N_14760,N_14677,N_14613);
nor U14761 (N_14761,N_14636,N_14572);
nor U14762 (N_14762,N_14689,N_14525);
nand U14763 (N_14763,N_14682,N_14538);
and U14764 (N_14764,N_14717,N_14644);
or U14765 (N_14765,N_14704,N_14674);
nand U14766 (N_14766,N_14647,N_14643);
nor U14767 (N_14767,N_14546,N_14507);
nand U14768 (N_14768,N_14610,N_14615);
xor U14769 (N_14769,N_14627,N_14560);
nor U14770 (N_14770,N_14743,N_14588);
or U14771 (N_14771,N_14716,N_14660);
nand U14772 (N_14772,N_14731,N_14548);
nor U14773 (N_14773,N_14536,N_14509);
nor U14774 (N_14774,N_14718,N_14736);
or U14775 (N_14775,N_14719,N_14634);
or U14776 (N_14776,N_14519,N_14730);
nor U14777 (N_14777,N_14597,N_14699);
or U14778 (N_14778,N_14667,N_14528);
nand U14779 (N_14779,N_14524,N_14591);
nor U14780 (N_14780,N_14558,N_14656);
nand U14781 (N_14781,N_14621,N_14672);
xor U14782 (N_14782,N_14709,N_14612);
nand U14783 (N_14783,N_14665,N_14724);
and U14784 (N_14784,N_14521,N_14715);
xor U14785 (N_14785,N_14511,N_14629);
xnor U14786 (N_14786,N_14744,N_14729);
xor U14787 (N_14787,N_14520,N_14600);
and U14788 (N_14788,N_14734,N_14611);
nand U14789 (N_14789,N_14529,N_14574);
nand U14790 (N_14790,N_14628,N_14728);
and U14791 (N_14791,N_14543,N_14745);
xnor U14792 (N_14792,N_14534,N_14586);
nor U14793 (N_14793,N_14504,N_14658);
xor U14794 (N_14794,N_14514,N_14710);
and U14795 (N_14795,N_14642,N_14593);
nor U14796 (N_14796,N_14670,N_14669);
and U14797 (N_14797,N_14695,N_14622);
and U14798 (N_14798,N_14609,N_14510);
nand U14799 (N_14799,N_14696,N_14706);
nor U14800 (N_14800,N_14726,N_14500);
xor U14801 (N_14801,N_14575,N_14581);
nand U14802 (N_14802,N_14678,N_14614);
nand U14803 (N_14803,N_14617,N_14501);
xnor U14804 (N_14804,N_14623,N_14596);
or U14805 (N_14805,N_14723,N_14701);
and U14806 (N_14806,N_14566,N_14517);
and U14807 (N_14807,N_14637,N_14631);
and U14808 (N_14808,N_14583,N_14662);
nand U14809 (N_14809,N_14714,N_14516);
and U14810 (N_14810,N_14604,N_14578);
or U14811 (N_14811,N_14570,N_14607);
nor U14812 (N_14812,N_14652,N_14552);
nor U14813 (N_14813,N_14741,N_14576);
xnor U14814 (N_14814,N_14561,N_14685);
nand U14815 (N_14815,N_14742,N_14589);
nor U14816 (N_14816,N_14545,N_14648);
nand U14817 (N_14817,N_14563,N_14638);
xor U14818 (N_14818,N_14749,N_14721);
and U14819 (N_14819,N_14539,N_14577);
and U14820 (N_14820,N_14567,N_14722);
nor U14821 (N_14821,N_14544,N_14556);
nand U14822 (N_14822,N_14748,N_14502);
xnor U14823 (N_14823,N_14703,N_14657);
and U14824 (N_14824,N_14565,N_14740);
xor U14825 (N_14825,N_14735,N_14681);
xor U14826 (N_14826,N_14702,N_14738);
nor U14827 (N_14827,N_14518,N_14698);
xor U14828 (N_14828,N_14680,N_14679);
or U14829 (N_14829,N_14568,N_14630);
nor U14830 (N_14830,N_14587,N_14569);
xor U14831 (N_14831,N_14603,N_14503);
nor U14832 (N_14832,N_14562,N_14512);
nand U14833 (N_14833,N_14616,N_14505);
and U14834 (N_14834,N_14564,N_14585);
nor U14835 (N_14835,N_14661,N_14533);
nand U14836 (N_14836,N_14747,N_14690);
nand U14837 (N_14837,N_14697,N_14532);
or U14838 (N_14838,N_14555,N_14515);
nor U14839 (N_14839,N_14606,N_14513);
or U14840 (N_14840,N_14625,N_14693);
or U14841 (N_14841,N_14664,N_14620);
xnor U14842 (N_14842,N_14541,N_14653);
nand U14843 (N_14843,N_14590,N_14632);
and U14844 (N_14844,N_14550,N_14523);
or U14845 (N_14845,N_14599,N_14687);
xnor U14846 (N_14846,N_14739,N_14535);
nor U14847 (N_14847,N_14571,N_14691);
or U14848 (N_14848,N_14650,N_14640);
and U14849 (N_14849,N_14618,N_14727);
or U14850 (N_14850,N_14746,N_14707);
nor U14851 (N_14851,N_14666,N_14633);
nor U14852 (N_14852,N_14683,N_14655);
xnor U14853 (N_14853,N_14601,N_14712);
or U14854 (N_14854,N_14711,N_14530);
nand U14855 (N_14855,N_14635,N_14602);
nor U14856 (N_14856,N_14542,N_14732);
xor U14857 (N_14857,N_14705,N_14733);
xor U14858 (N_14858,N_14624,N_14508);
nand U14859 (N_14859,N_14547,N_14668);
nand U14860 (N_14860,N_14684,N_14549);
nand U14861 (N_14861,N_14526,N_14584);
or U14862 (N_14862,N_14580,N_14708);
nor U14863 (N_14863,N_14688,N_14649);
xnor U14864 (N_14864,N_14725,N_14579);
nand U14865 (N_14865,N_14645,N_14553);
and U14866 (N_14866,N_14592,N_14559);
or U14867 (N_14867,N_14694,N_14608);
or U14868 (N_14868,N_14626,N_14641);
or U14869 (N_14869,N_14651,N_14557);
nor U14870 (N_14870,N_14737,N_14646);
or U14871 (N_14871,N_14700,N_14551);
nand U14872 (N_14872,N_14594,N_14527);
and U14873 (N_14873,N_14663,N_14686);
nand U14874 (N_14874,N_14537,N_14675);
and U14875 (N_14875,N_14688,N_14505);
or U14876 (N_14876,N_14648,N_14655);
nor U14877 (N_14877,N_14701,N_14742);
nor U14878 (N_14878,N_14515,N_14672);
and U14879 (N_14879,N_14726,N_14527);
xor U14880 (N_14880,N_14654,N_14630);
or U14881 (N_14881,N_14588,N_14537);
and U14882 (N_14882,N_14540,N_14689);
nand U14883 (N_14883,N_14619,N_14661);
nand U14884 (N_14884,N_14588,N_14544);
or U14885 (N_14885,N_14619,N_14561);
nor U14886 (N_14886,N_14566,N_14652);
nor U14887 (N_14887,N_14744,N_14562);
and U14888 (N_14888,N_14647,N_14595);
nor U14889 (N_14889,N_14736,N_14692);
and U14890 (N_14890,N_14683,N_14598);
or U14891 (N_14891,N_14697,N_14648);
xor U14892 (N_14892,N_14630,N_14677);
nor U14893 (N_14893,N_14628,N_14664);
and U14894 (N_14894,N_14515,N_14656);
nand U14895 (N_14895,N_14607,N_14679);
nand U14896 (N_14896,N_14644,N_14556);
or U14897 (N_14897,N_14536,N_14531);
and U14898 (N_14898,N_14502,N_14594);
nor U14899 (N_14899,N_14535,N_14561);
or U14900 (N_14900,N_14635,N_14525);
xnor U14901 (N_14901,N_14705,N_14724);
xor U14902 (N_14902,N_14633,N_14649);
or U14903 (N_14903,N_14525,N_14663);
or U14904 (N_14904,N_14721,N_14665);
xor U14905 (N_14905,N_14710,N_14530);
or U14906 (N_14906,N_14668,N_14725);
nand U14907 (N_14907,N_14691,N_14687);
xnor U14908 (N_14908,N_14690,N_14645);
and U14909 (N_14909,N_14658,N_14693);
nor U14910 (N_14910,N_14532,N_14729);
xor U14911 (N_14911,N_14540,N_14661);
nand U14912 (N_14912,N_14606,N_14602);
and U14913 (N_14913,N_14625,N_14746);
and U14914 (N_14914,N_14621,N_14689);
or U14915 (N_14915,N_14538,N_14619);
nor U14916 (N_14916,N_14622,N_14652);
or U14917 (N_14917,N_14708,N_14511);
nor U14918 (N_14918,N_14623,N_14599);
nor U14919 (N_14919,N_14507,N_14650);
nor U14920 (N_14920,N_14733,N_14687);
or U14921 (N_14921,N_14613,N_14598);
nand U14922 (N_14922,N_14666,N_14611);
xnor U14923 (N_14923,N_14624,N_14604);
and U14924 (N_14924,N_14732,N_14644);
nand U14925 (N_14925,N_14545,N_14605);
or U14926 (N_14926,N_14510,N_14516);
xnor U14927 (N_14927,N_14667,N_14612);
or U14928 (N_14928,N_14652,N_14661);
nand U14929 (N_14929,N_14534,N_14720);
nor U14930 (N_14930,N_14557,N_14655);
nor U14931 (N_14931,N_14501,N_14708);
and U14932 (N_14932,N_14715,N_14672);
xnor U14933 (N_14933,N_14548,N_14738);
nand U14934 (N_14934,N_14543,N_14735);
or U14935 (N_14935,N_14708,N_14736);
xnor U14936 (N_14936,N_14734,N_14595);
nand U14937 (N_14937,N_14648,N_14667);
or U14938 (N_14938,N_14500,N_14634);
xnor U14939 (N_14939,N_14500,N_14589);
and U14940 (N_14940,N_14671,N_14606);
nor U14941 (N_14941,N_14700,N_14515);
and U14942 (N_14942,N_14740,N_14692);
nor U14943 (N_14943,N_14568,N_14540);
xor U14944 (N_14944,N_14570,N_14737);
nand U14945 (N_14945,N_14640,N_14696);
or U14946 (N_14946,N_14700,N_14502);
nand U14947 (N_14947,N_14520,N_14737);
or U14948 (N_14948,N_14693,N_14611);
xnor U14949 (N_14949,N_14710,N_14724);
nor U14950 (N_14950,N_14581,N_14608);
nand U14951 (N_14951,N_14567,N_14512);
and U14952 (N_14952,N_14552,N_14545);
nand U14953 (N_14953,N_14669,N_14716);
nor U14954 (N_14954,N_14688,N_14736);
xor U14955 (N_14955,N_14527,N_14623);
xor U14956 (N_14956,N_14724,N_14597);
xor U14957 (N_14957,N_14628,N_14599);
and U14958 (N_14958,N_14528,N_14605);
and U14959 (N_14959,N_14591,N_14581);
xnor U14960 (N_14960,N_14587,N_14724);
xnor U14961 (N_14961,N_14533,N_14745);
xor U14962 (N_14962,N_14572,N_14590);
nor U14963 (N_14963,N_14553,N_14699);
nor U14964 (N_14964,N_14735,N_14658);
nor U14965 (N_14965,N_14742,N_14514);
and U14966 (N_14966,N_14502,N_14580);
nor U14967 (N_14967,N_14720,N_14531);
nand U14968 (N_14968,N_14597,N_14558);
xor U14969 (N_14969,N_14539,N_14536);
nand U14970 (N_14970,N_14536,N_14571);
nor U14971 (N_14971,N_14706,N_14714);
and U14972 (N_14972,N_14522,N_14649);
and U14973 (N_14973,N_14599,N_14519);
nor U14974 (N_14974,N_14711,N_14510);
or U14975 (N_14975,N_14696,N_14648);
nand U14976 (N_14976,N_14692,N_14578);
nor U14977 (N_14977,N_14621,N_14735);
or U14978 (N_14978,N_14683,N_14692);
or U14979 (N_14979,N_14581,N_14611);
and U14980 (N_14980,N_14669,N_14613);
nand U14981 (N_14981,N_14707,N_14530);
nor U14982 (N_14982,N_14724,N_14685);
or U14983 (N_14983,N_14578,N_14523);
or U14984 (N_14984,N_14665,N_14595);
nand U14985 (N_14985,N_14652,N_14709);
and U14986 (N_14986,N_14692,N_14667);
and U14987 (N_14987,N_14536,N_14506);
and U14988 (N_14988,N_14527,N_14660);
and U14989 (N_14989,N_14660,N_14645);
nor U14990 (N_14990,N_14669,N_14569);
and U14991 (N_14991,N_14638,N_14516);
nor U14992 (N_14992,N_14508,N_14571);
nand U14993 (N_14993,N_14531,N_14731);
nor U14994 (N_14994,N_14508,N_14599);
nor U14995 (N_14995,N_14665,N_14563);
and U14996 (N_14996,N_14672,N_14530);
and U14997 (N_14997,N_14664,N_14624);
and U14998 (N_14998,N_14692,N_14727);
xor U14999 (N_14999,N_14680,N_14654);
and U15000 (N_15000,N_14858,N_14758);
and U15001 (N_15001,N_14864,N_14873);
or U15002 (N_15002,N_14831,N_14884);
xnor U15003 (N_15003,N_14988,N_14806);
xor U15004 (N_15004,N_14970,N_14991);
nor U15005 (N_15005,N_14801,N_14824);
and U15006 (N_15006,N_14766,N_14832);
and U15007 (N_15007,N_14881,N_14963);
nand U15008 (N_15008,N_14779,N_14962);
nor U15009 (N_15009,N_14827,N_14756);
nor U15010 (N_15010,N_14867,N_14793);
or U15011 (N_15011,N_14961,N_14948);
and U15012 (N_15012,N_14949,N_14938);
xor U15013 (N_15013,N_14753,N_14854);
or U15014 (N_15014,N_14840,N_14856);
nor U15015 (N_15015,N_14800,N_14876);
and U15016 (N_15016,N_14907,N_14956);
nor U15017 (N_15017,N_14828,N_14857);
and U15018 (N_15018,N_14814,N_14787);
nand U15019 (N_15019,N_14791,N_14983);
xor U15020 (N_15020,N_14768,N_14982);
xor U15021 (N_15021,N_14880,N_14958);
and U15022 (N_15022,N_14789,N_14941);
nor U15023 (N_15023,N_14936,N_14860);
nor U15024 (N_15024,N_14946,N_14959);
nor U15025 (N_15025,N_14843,N_14917);
nand U15026 (N_15026,N_14821,N_14759);
and U15027 (N_15027,N_14790,N_14967);
or U15028 (N_15028,N_14829,N_14803);
nand U15029 (N_15029,N_14998,N_14819);
xnor U15030 (N_15030,N_14862,N_14834);
nor U15031 (N_15031,N_14947,N_14833);
and U15032 (N_15032,N_14909,N_14934);
or U15033 (N_15033,N_14925,N_14937);
nor U15034 (N_15034,N_14751,N_14839);
and U15035 (N_15035,N_14808,N_14830);
nand U15036 (N_15036,N_14866,N_14969);
xnor U15037 (N_15037,N_14823,N_14841);
and U15038 (N_15038,N_14820,N_14945);
nor U15039 (N_15039,N_14942,N_14782);
and U15040 (N_15040,N_14986,N_14811);
or U15041 (N_15041,N_14897,N_14900);
nand U15042 (N_15042,N_14794,N_14853);
or U15043 (N_15043,N_14943,N_14906);
xor U15044 (N_15044,N_14773,N_14874);
or U15045 (N_15045,N_14926,N_14971);
nor U15046 (N_15046,N_14780,N_14930);
nor U15047 (N_15047,N_14771,N_14836);
or U15048 (N_15048,N_14763,N_14918);
nor U15049 (N_15049,N_14885,N_14972);
xor U15050 (N_15050,N_14888,N_14848);
nand U15051 (N_15051,N_14895,N_14877);
nand U15052 (N_15052,N_14929,N_14996);
or U15053 (N_15053,N_14919,N_14902);
nor U15054 (N_15054,N_14985,N_14898);
xnor U15055 (N_15055,N_14966,N_14924);
xor U15056 (N_15056,N_14990,N_14810);
and U15057 (N_15057,N_14783,N_14765);
xor U15058 (N_15058,N_14863,N_14932);
nand U15059 (N_15059,N_14792,N_14788);
or U15060 (N_15060,N_14802,N_14978);
or U15061 (N_15061,N_14825,N_14950);
nor U15062 (N_15062,N_14980,N_14994);
and U15063 (N_15063,N_14894,N_14842);
and U15064 (N_15064,N_14981,N_14807);
xnor U15065 (N_15065,N_14844,N_14754);
nand U15066 (N_15066,N_14775,N_14769);
nor U15067 (N_15067,N_14940,N_14855);
and U15068 (N_15068,N_14975,N_14851);
xnor U15069 (N_15069,N_14837,N_14822);
nor U15070 (N_15070,N_14955,N_14987);
nor U15071 (N_15071,N_14799,N_14984);
xnor U15072 (N_15072,N_14838,N_14939);
nand U15073 (N_15073,N_14952,N_14847);
xor U15074 (N_15074,N_14868,N_14915);
xor U15075 (N_15075,N_14770,N_14908);
or U15076 (N_15076,N_14933,N_14826);
xor U15077 (N_15077,N_14977,N_14797);
and U15078 (N_15078,N_14974,N_14859);
nor U15079 (N_15079,N_14910,N_14953);
or U15080 (N_15080,N_14992,N_14879);
or U15081 (N_15081,N_14812,N_14813);
and U15082 (N_15082,N_14935,N_14944);
or U15083 (N_15083,N_14761,N_14968);
nor U15084 (N_15084,N_14784,N_14786);
xor U15085 (N_15085,N_14989,N_14951);
or U15086 (N_15086,N_14889,N_14960);
nand U15087 (N_15087,N_14916,N_14928);
xnor U15088 (N_15088,N_14922,N_14817);
nor U15089 (N_15089,N_14999,N_14809);
nand U15090 (N_15090,N_14805,N_14890);
xor U15091 (N_15091,N_14954,N_14870);
nand U15092 (N_15092,N_14965,N_14816);
nand U15093 (N_15093,N_14912,N_14875);
or U15094 (N_15094,N_14893,N_14796);
or U15095 (N_15095,N_14976,N_14750);
nor U15096 (N_15096,N_14845,N_14869);
or U15097 (N_15097,N_14997,N_14767);
xor U15098 (N_15098,N_14896,N_14891);
or U15099 (N_15099,N_14887,N_14849);
nor U15100 (N_15100,N_14850,N_14852);
and U15101 (N_15101,N_14979,N_14911);
and U15102 (N_15102,N_14993,N_14927);
or U15103 (N_15103,N_14872,N_14755);
nand U15104 (N_15104,N_14904,N_14774);
nor U15105 (N_15105,N_14760,N_14964);
and U15106 (N_15106,N_14764,N_14776);
nand U15107 (N_15107,N_14995,N_14762);
nor U15108 (N_15108,N_14901,N_14804);
nor U15109 (N_15109,N_14921,N_14777);
xnor U15110 (N_15110,N_14957,N_14871);
nor U15111 (N_15111,N_14886,N_14899);
and U15112 (N_15112,N_14778,N_14883);
nor U15113 (N_15113,N_14757,N_14903);
nand U15114 (N_15114,N_14835,N_14846);
nor U15115 (N_15115,N_14892,N_14865);
xnor U15116 (N_15116,N_14905,N_14798);
and U15117 (N_15117,N_14785,N_14752);
or U15118 (N_15118,N_14920,N_14913);
or U15119 (N_15119,N_14973,N_14878);
nand U15120 (N_15120,N_14931,N_14795);
nor U15121 (N_15121,N_14923,N_14818);
or U15122 (N_15122,N_14914,N_14781);
xnor U15123 (N_15123,N_14772,N_14815);
nand U15124 (N_15124,N_14882,N_14861);
nor U15125 (N_15125,N_14997,N_14766);
nand U15126 (N_15126,N_14876,N_14813);
nor U15127 (N_15127,N_14869,N_14821);
xor U15128 (N_15128,N_14839,N_14907);
and U15129 (N_15129,N_14769,N_14844);
and U15130 (N_15130,N_14880,N_14932);
nand U15131 (N_15131,N_14783,N_14823);
nor U15132 (N_15132,N_14786,N_14948);
and U15133 (N_15133,N_14796,N_14858);
nand U15134 (N_15134,N_14803,N_14786);
and U15135 (N_15135,N_14755,N_14843);
xor U15136 (N_15136,N_14876,N_14952);
nor U15137 (N_15137,N_14919,N_14814);
or U15138 (N_15138,N_14786,N_14878);
nand U15139 (N_15139,N_14869,N_14814);
nor U15140 (N_15140,N_14764,N_14903);
and U15141 (N_15141,N_14967,N_14752);
nand U15142 (N_15142,N_14928,N_14955);
or U15143 (N_15143,N_14968,N_14922);
or U15144 (N_15144,N_14807,N_14792);
xnor U15145 (N_15145,N_14863,N_14781);
nor U15146 (N_15146,N_14893,N_14982);
and U15147 (N_15147,N_14877,N_14802);
xnor U15148 (N_15148,N_14954,N_14772);
xor U15149 (N_15149,N_14905,N_14814);
nor U15150 (N_15150,N_14917,N_14890);
nor U15151 (N_15151,N_14985,N_14991);
and U15152 (N_15152,N_14893,N_14788);
and U15153 (N_15153,N_14960,N_14979);
and U15154 (N_15154,N_14790,N_14787);
and U15155 (N_15155,N_14980,N_14945);
nor U15156 (N_15156,N_14854,N_14921);
xor U15157 (N_15157,N_14840,N_14946);
or U15158 (N_15158,N_14804,N_14911);
nor U15159 (N_15159,N_14861,N_14837);
and U15160 (N_15160,N_14826,N_14880);
nand U15161 (N_15161,N_14948,N_14886);
nor U15162 (N_15162,N_14871,N_14900);
and U15163 (N_15163,N_14929,N_14793);
nand U15164 (N_15164,N_14907,N_14826);
and U15165 (N_15165,N_14774,N_14967);
nor U15166 (N_15166,N_14763,N_14770);
or U15167 (N_15167,N_14985,N_14970);
nand U15168 (N_15168,N_14806,N_14952);
and U15169 (N_15169,N_14948,N_14814);
or U15170 (N_15170,N_14766,N_14806);
nor U15171 (N_15171,N_14949,N_14896);
and U15172 (N_15172,N_14755,N_14762);
nand U15173 (N_15173,N_14912,N_14878);
nor U15174 (N_15174,N_14848,N_14825);
and U15175 (N_15175,N_14992,N_14908);
nor U15176 (N_15176,N_14990,N_14757);
xnor U15177 (N_15177,N_14912,N_14871);
nor U15178 (N_15178,N_14831,N_14930);
nand U15179 (N_15179,N_14895,N_14848);
xnor U15180 (N_15180,N_14955,N_14822);
nor U15181 (N_15181,N_14863,N_14771);
nor U15182 (N_15182,N_14904,N_14764);
or U15183 (N_15183,N_14860,N_14944);
xor U15184 (N_15184,N_14962,N_14955);
xnor U15185 (N_15185,N_14849,N_14928);
nor U15186 (N_15186,N_14944,N_14814);
nand U15187 (N_15187,N_14924,N_14940);
xor U15188 (N_15188,N_14995,N_14776);
or U15189 (N_15189,N_14906,N_14771);
nor U15190 (N_15190,N_14957,N_14997);
nand U15191 (N_15191,N_14917,N_14784);
nor U15192 (N_15192,N_14900,N_14818);
nor U15193 (N_15193,N_14778,N_14900);
nand U15194 (N_15194,N_14757,N_14939);
nand U15195 (N_15195,N_14944,N_14807);
and U15196 (N_15196,N_14967,N_14876);
xor U15197 (N_15197,N_14828,N_14790);
and U15198 (N_15198,N_14846,N_14975);
and U15199 (N_15199,N_14771,N_14860);
nor U15200 (N_15200,N_14830,N_14978);
or U15201 (N_15201,N_14962,N_14973);
xor U15202 (N_15202,N_14979,N_14794);
and U15203 (N_15203,N_14927,N_14844);
nand U15204 (N_15204,N_14881,N_14937);
nor U15205 (N_15205,N_14799,N_14854);
and U15206 (N_15206,N_14817,N_14931);
xnor U15207 (N_15207,N_14787,N_14967);
and U15208 (N_15208,N_14874,N_14949);
xor U15209 (N_15209,N_14832,N_14972);
and U15210 (N_15210,N_14913,N_14888);
or U15211 (N_15211,N_14907,N_14775);
and U15212 (N_15212,N_14818,N_14984);
xnor U15213 (N_15213,N_14766,N_14972);
nor U15214 (N_15214,N_14873,N_14834);
nor U15215 (N_15215,N_14935,N_14919);
nand U15216 (N_15216,N_14857,N_14874);
xor U15217 (N_15217,N_14840,N_14933);
or U15218 (N_15218,N_14799,N_14866);
nor U15219 (N_15219,N_14786,N_14830);
nor U15220 (N_15220,N_14945,N_14908);
nor U15221 (N_15221,N_14808,N_14870);
and U15222 (N_15222,N_14890,N_14950);
and U15223 (N_15223,N_14789,N_14808);
nor U15224 (N_15224,N_14997,N_14949);
nor U15225 (N_15225,N_14841,N_14991);
nand U15226 (N_15226,N_14755,N_14833);
and U15227 (N_15227,N_14856,N_14819);
xnor U15228 (N_15228,N_14842,N_14812);
nand U15229 (N_15229,N_14947,N_14807);
and U15230 (N_15230,N_14848,N_14872);
nor U15231 (N_15231,N_14886,N_14924);
nor U15232 (N_15232,N_14825,N_14800);
nand U15233 (N_15233,N_14999,N_14864);
nand U15234 (N_15234,N_14948,N_14873);
and U15235 (N_15235,N_14976,N_14905);
nand U15236 (N_15236,N_14930,N_14844);
or U15237 (N_15237,N_14897,N_14803);
nand U15238 (N_15238,N_14832,N_14879);
xor U15239 (N_15239,N_14972,N_14760);
and U15240 (N_15240,N_14750,N_14771);
xnor U15241 (N_15241,N_14976,N_14892);
nor U15242 (N_15242,N_14987,N_14905);
and U15243 (N_15243,N_14998,N_14978);
and U15244 (N_15244,N_14904,N_14966);
xnor U15245 (N_15245,N_14939,N_14896);
or U15246 (N_15246,N_14945,N_14951);
or U15247 (N_15247,N_14853,N_14831);
nor U15248 (N_15248,N_14823,N_14835);
and U15249 (N_15249,N_14891,N_14820);
nand U15250 (N_15250,N_15160,N_15036);
or U15251 (N_15251,N_15122,N_15235);
nor U15252 (N_15252,N_15123,N_15118);
xor U15253 (N_15253,N_15127,N_15230);
nor U15254 (N_15254,N_15059,N_15001);
and U15255 (N_15255,N_15194,N_15078);
and U15256 (N_15256,N_15208,N_15172);
and U15257 (N_15257,N_15136,N_15093);
nand U15258 (N_15258,N_15096,N_15198);
or U15259 (N_15259,N_15181,N_15120);
and U15260 (N_15260,N_15183,N_15132);
nand U15261 (N_15261,N_15023,N_15197);
and U15262 (N_15262,N_15141,N_15081);
or U15263 (N_15263,N_15089,N_15018);
nor U15264 (N_15264,N_15114,N_15144);
nand U15265 (N_15265,N_15157,N_15206);
and U15266 (N_15266,N_15241,N_15137);
or U15267 (N_15267,N_15050,N_15091);
and U15268 (N_15268,N_15138,N_15038);
xnor U15269 (N_15269,N_15193,N_15066);
nor U15270 (N_15270,N_15151,N_15043);
nand U15271 (N_15271,N_15247,N_15051);
nand U15272 (N_15272,N_15164,N_15039);
nor U15273 (N_15273,N_15025,N_15006);
nor U15274 (N_15274,N_15130,N_15178);
and U15275 (N_15275,N_15228,N_15248);
nor U15276 (N_15276,N_15162,N_15209);
and U15277 (N_15277,N_15238,N_15147);
or U15278 (N_15278,N_15163,N_15010);
and U15279 (N_15279,N_15040,N_15180);
or U15280 (N_15280,N_15155,N_15104);
and U15281 (N_15281,N_15105,N_15071);
xor U15282 (N_15282,N_15037,N_15200);
and U15283 (N_15283,N_15218,N_15046);
and U15284 (N_15284,N_15220,N_15211);
or U15285 (N_15285,N_15229,N_15214);
nor U15286 (N_15286,N_15210,N_15012);
nand U15287 (N_15287,N_15140,N_15126);
nand U15288 (N_15288,N_15034,N_15222);
nor U15289 (N_15289,N_15226,N_15148);
nor U15290 (N_15290,N_15237,N_15005);
nand U15291 (N_15291,N_15027,N_15143);
xor U15292 (N_15292,N_15075,N_15170);
and U15293 (N_15293,N_15191,N_15113);
nand U15294 (N_15294,N_15103,N_15233);
xor U15295 (N_15295,N_15047,N_15174);
and U15296 (N_15296,N_15240,N_15003);
nor U15297 (N_15297,N_15195,N_15024);
and U15298 (N_15298,N_15074,N_15135);
nor U15299 (N_15299,N_15020,N_15227);
or U15300 (N_15300,N_15186,N_15219);
nand U15301 (N_15301,N_15205,N_15041);
and U15302 (N_15302,N_15000,N_15097);
nand U15303 (N_15303,N_15142,N_15095);
nor U15304 (N_15304,N_15225,N_15029);
nor U15305 (N_15305,N_15079,N_15058);
and U15306 (N_15306,N_15080,N_15030);
nand U15307 (N_15307,N_15112,N_15125);
or U15308 (N_15308,N_15249,N_15086);
nand U15309 (N_15309,N_15007,N_15028);
nor U15310 (N_15310,N_15049,N_15070);
and U15311 (N_15311,N_15201,N_15109);
nand U15312 (N_15312,N_15062,N_15239);
and U15313 (N_15313,N_15108,N_15173);
nor U15314 (N_15314,N_15221,N_15026);
and U15315 (N_15315,N_15053,N_15152);
xnor U15316 (N_15316,N_15016,N_15159);
nand U15317 (N_15317,N_15176,N_15084);
and U15318 (N_15318,N_15196,N_15192);
nand U15319 (N_15319,N_15085,N_15110);
xor U15320 (N_15320,N_15098,N_15061);
xnor U15321 (N_15321,N_15116,N_15242);
xnor U15322 (N_15322,N_15231,N_15213);
or U15323 (N_15323,N_15002,N_15131);
nand U15324 (N_15324,N_15014,N_15133);
xnor U15325 (N_15325,N_15063,N_15128);
or U15326 (N_15326,N_15184,N_15232);
nor U15327 (N_15327,N_15179,N_15045);
or U15328 (N_15328,N_15124,N_15011);
and U15329 (N_15329,N_15150,N_15008);
xor U15330 (N_15330,N_15044,N_15154);
xnor U15331 (N_15331,N_15129,N_15202);
and U15332 (N_15332,N_15244,N_15065);
nand U15333 (N_15333,N_15019,N_15056);
and U15334 (N_15334,N_15153,N_15013);
xnor U15335 (N_15335,N_15111,N_15171);
and U15336 (N_15336,N_15033,N_15067);
or U15337 (N_15337,N_15161,N_15100);
nand U15338 (N_15338,N_15055,N_15117);
xor U15339 (N_15339,N_15064,N_15057);
and U15340 (N_15340,N_15015,N_15060);
or U15341 (N_15341,N_15189,N_15145);
xnor U15342 (N_15342,N_15243,N_15004);
and U15343 (N_15343,N_15092,N_15169);
or U15344 (N_15344,N_15199,N_15156);
nand U15345 (N_15345,N_15077,N_15094);
nand U15346 (N_15346,N_15099,N_15035);
nand U15347 (N_15347,N_15009,N_15182);
and U15348 (N_15348,N_15236,N_15021);
and U15349 (N_15349,N_15102,N_15134);
xor U15350 (N_15350,N_15106,N_15223);
or U15351 (N_15351,N_15217,N_15207);
xor U15352 (N_15352,N_15088,N_15073);
xnor U15353 (N_15353,N_15168,N_15187);
or U15354 (N_15354,N_15017,N_15101);
xnor U15355 (N_15355,N_15224,N_15119);
nor U15356 (N_15356,N_15146,N_15177);
nor U15357 (N_15357,N_15022,N_15166);
nand U15358 (N_15358,N_15076,N_15139);
or U15359 (N_15359,N_15069,N_15032);
or U15360 (N_15360,N_15082,N_15054);
or U15361 (N_15361,N_15052,N_15175);
nand U15362 (N_15362,N_15216,N_15188);
or U15363 (N_15363,N_15190,N_15090);
or U15364 (N_15364,N_15031,N_15068);
xnor U15365 (N_15365,N_15107,N_15204);
xor U15366 (N_15366,N_15121,N_15215);
nand U15367 (N_15367,N_15234,N_15203);
xor U15368 (N_15368,N_15042,N_15048);
nand U15369 (N_15369,N_15246,N_15245);
nand U15370 (N_15370,N_15087,N_15165);
nand U15371 (N_15371,N_15072,N_15167);
nor U15372 (N_15372,N_15185,N_15149);
nor U15373 (N_15373,N_15212,N_15115);
and U15374 (N_15374,N_15083,N_15158);
nand U15375 (N_15375,N_15109,N_15053);
nand U15376 (N_15376,N_15198,N_15159);
and U15377 (N_15377,N_15086,N_15157);
and U15378 (N_15378,N_15156,N_15180);
or U15379 (N_15379,N_15076,N_15174);
nand U15380 (N_15380,N_15000,N_15195);
and U15381 (N_15381,N_15173,N_15164);
nand U15382 (N_15382,N_15020,N_15224);
xor U15383 (N_15383,N_15036,N_15208);
nand U15384 (N_15384,N_15237,N_15075);
xnor U15385 (N_15385,N_15105,N_15013);
xnor U15386 (N_15386,N_15077,N_15125);
and U15387 (N_15387,N_15018,N_15001);
xor U15388 (N_15388,N_15123,N_15115);
xor U15389 (N_15389,N_15136,N_15103);
and U15390 (N_15390,N_15211,N_15025);
and U15391 (N_15391,N_15172,N_15037);
nand U15392 (N_15392,N_15080,N_15110);
xnor U15393 (N_15393,N_15059,N_15063);
nor U15394 (N_15394,N_15112,N_15070);
or U15395 (N_15395,N_15248,N_15062);
nand U15396 (N_15396,N_15138,N_15192);
nor U15397 (N_15397,N_15194,N_15133);
xnor U15398 (N_15398,N_15170,N_15165);
and U15399 (N_15399,N_15220,N_15191);
nor U15400 (N_15400,N_15201,N_15179);
or U15401 (N_15401,N_15115,N_15160);
nor U15402 (N_15402,N_15202,N_15009);
xor U15403 (N_15403,N_15192,N_15181);
nand U15404 (N_15404,N_15064,N_15183);
nor U15405 (N_15405,N_15222,N_15082);
or U15406 (N_15406,N_15126,N_15179);
and U15407 (N_15407,N_15089,N_15122);
xnor U15408 (N_15408,N_15083,N_15220);
nand U15409 (N_15409,N_15179,N_15090);
nor U15410 (N_15410,N_15102,N_15021);
and U15411 (N_15411,N_15203,N_15236);
or U15412 (N_15412,N_15047,N_15245);
nand U15413 (N_15413,N_15174,N_15123);
nor U15414 (N_15414,N_15153,N_15016);
nand U15415 (N_15415,N_15141,N_15186);
xor U15416 (N_15416,N_15003,N_15008);
xnor U15417 (N_15417,N_15153,N_15231);
nand U15418 (N_15418,N_15141,N_15136);
nor U15419 (N_15419,N_15181,N_15210);
or U15420 (N_15420,N_15231,N_15114);
and U15421 (N_15421,N_15194,N_15105);
xnor U15422 (N_15422,N_15134,N_15116);
nor U15423 (N_15423,N_15128,N_15067);
nor U15424 (N_15424,N_15103,N_15246);
or U15425 (N_15425,N_15152,N_15157);
nor U15426 (N_15426,N_15100,N_15191);
or U15427 (N_15427,N_15178,N_15179);
and U15428 (N_15428,N_15003,N_15058);
xnor U15429 (N_15429,N_15142,N_15086);
or U15430 (N_15430,N_15111,N_15038);
nand U15431 (N_15431,N_15142,N_15222);
or U15432 (N_15432,N_15150,N_15067);
nor U15433 (N_15433,N_15164,N_15013);
nor U15434 (N_15434,N_15083,N_15096);
nor U15435 (N_15435,N_15023,N_15005);
xor U15436 (N_15436,N_15013,N_15233);
nand U15437 (N_15437,N_15039,N_15195);
xnor U15438 (N_15438,N_15169,N_15086);
nor U15439 (N_15439,N_15089,N_15054);
nand U15440 (N_15440,N_15176,N_15219);
nand U15441 (N_15441,N_15143,N_15035);
or U15442 (N_15442,N_15114,N_15093);
nand U15443 (N_15443,N_15000,N_15091);
and U15444 (N_15444,N_15124,N_15047);
and U15445 (N_15445,N_15024,N_15000);
xnor U15446 (N_15446,N_15184,N_15249);
nor U15447 (N_15447,N_15074,N_15188);
and U15448 (N_15448,N_15032,N_15132);
and U15449 (N_15449,N_15199,N_15115);
nand U15450 (N_15450,N_15048,N_15211);
nand U15451 (N_15451,N_15195,N_15111);
nand U15452 (N_15452,N_15198,N_15080);
xnor U15453 (N_15453,N_15221,N_15034);
and U15454 (N_15454,N_15176,N_15089);
nand U15455 (N_15455,N_15143,N_15039);
and U15456 (N_15456,N_15168,N_15034);
nand U15457 (N_15457,N_15049,N_15222);
and U15458 (N_15458,N_15206,N_15138);
nor U15459 (N_15459,N_15233,N_15036);
and U15460 (N_15460,N_15021,N_15206);
or U15461 (N_15461,N_15101,N_15224);
nand U15462 (N_15462,N_15108,N_15048);
and U15463 (N_15463,N_15091,N_15245);
or U15464 (N_15464,N_15054,N_15163);
xnor U15465 (N_15465,N_15056,N_15236);
and U15466 (N_15466,N_15158,N_15233);
and U15467 (N_15467,N_15128,N_15247);
xor U15468 (N_15468,N_15194,N_15192);
xor U15469 (N_15469,N_15191,N_15230);
or U15470 (N_15470,N_15016,N_15196);
nor U15471 (N_15471,N_15041,N_15031);
xnor U15472 (N_15472,N_15207,N_15040);
and U15473 (N_15473,N_15173,N_15174);
nor U15474 (N_15474,N_15062,N_15016);
or U15475 (N_15475,N_15227,N_15088);
or U15476 (N_15476,N_15078,N_15005);
and U15477 (N_15477,N_15191,N_15004);
and U15478 (N_15478,N_15120,N_15003);
and U15479 (N_15479,N_15165,N_15043);
or U15480 (N_15480,N_15225,N_15209);
or U15481 (N_15481,N_15139,N_15035);
nand U15482 (N_15482,N_15056,N_15079);
or U15483 (N_15483,N_15060,N_15037);
and U15484 (N_15484,N_15168,N_15083);
and U15485 (N_15485,N_15176,N_15137);
xnor U15486 (N_15486,N_15238,N_15190);
and U15487 (N_15487,N_15028,N_15094);
nand U15488 (N_15488,N_15192,N_15070);
or U15489 (N_15489,N_15026,N_15174);
xnor U15490 (N_15490,N_15240,N_15032);
xor U15491 (N_15491,N_15172,N_15141);
xor U15492 (N_15492,N_15043,N_15091);
nor U15493 (N_15493,N_15133,N_15185);
xnor U15494 (N_15494,N_15157,N_15149);
and U15495 (N_15495,N_15063,N_15090);
nand U15496 (N_15496,N_15063,N_15186);
nor U15497 (N_15497,N_15121,N_15035);
and U15498 (N_15498,N_15153,N_15041);
nand U15499 (N_15499,N_15087,N_15020);
nand U15500 (N_15500,N_15375,N_15273);
or U15501 (N_15501,N_15268,N_15308);
or U15502 (N_15502,N_15442,N_15413);
xor U15503 (N_15503,N_15400,N_15383);
nand U15504 (N_15504,N_15275,N_15347);
nor U15505 (N_15505,N_15491,N_15422);
xor U15506 (N_15506,N_15495,N_15387);
xor U15507 (N_15507,N_15298,N_15267);
or U15508 (N_15508,N_15465,N_15306);
and U15509 (N_15509,N_15489,N_15282);
and U15510 (N_15510,N_15264,N_15434);
xor U15511 (N_15511,N_15300,N_15263);
nor U15512 (N_15512,N_15470,N_15497);
and U15513 (N_15513,N_15295,N_15418);
xnor U15514 (N_15514,N_15441,N_15485);
nand U15515 (N_15515,N_15254,N_15419);
and U15516 (N_15516,N_15468,N_15457);
and U15517 (N_15517,N_15374,N_15394);
nor U15518 (N_15518,N_15493,N_15321);
nand U15519 (N_15519,N_15367,N_15487);
or U15520 (N_15520,N_15408,N_15381);
xnor U15521 (N_15521,N_15437,N_15463);
and U15522 (N_15522,N_15483,N_15490);
and U15523 (N_15523,N_15399,N_15471);
and U15524 (N_15524,N_15351,N_15378);
and U15525 (N_15525,N_15499,N_15426);
or U15526 (N_15526,N_15265,N_15309);
nand U15527 (N_15527,N_15409,N_15476);
nand U15528 (N_15528,N_15281,N_15481);
xnor U15529 (N_15529,N_15395,N_15352);
nor U15530 (N_15530,N_15360,N_15388);
nor U15531 (N_15531,N_15432,N_15416);
nand U15532 (N_15532,N_15301,N_15317);
or U15533 (N_15533,N_15252,N_15278);
xor U15534 (N_15534,N_15276,N_15405);
nor U15535 (N_15535,N_15285,N_15448);
and U15536 (N_15536,N_15447,N_15337);
or U15537 (N_15537,N_15255,N_15456);
or U15538 (N_15538,N_15289,N_15404);
xor U15539 (N_15539,N_15326,N_15461);
nand U15540 (N_15540,N_15488,N_15294);
or U15541 (N_15541,N_15435,N_15496);
xnor U15542 (N_15542,N_15407,N_15284);
and U15543 (N_15543,N_15296,N_15303);
xor U15544 (N_15544,N_15323,N_15458);
xor U15545 (N_15545,N_15477,N_15357);
and U15546 (N_15546,N_15396,N_15454);
and U15547 (N_15547,N_15322,N_15312);
and U15548 (N_15548,N_15258,N_15302);
nand U15549 (N_15549,N_15433,N_15266);
and U15550 (N_15550,N_15443,N_15260);
nand U15551 (N_15551,N_15256,N_15333);
nor U15552 (N_15552,N_15286,N_15444);
nand U15553 (N_15553,N_15462,N_15412);
nor U15554 (N_15554,N_15425,N_15349);
or U15555 (N_15555,N_15459,N_15280);
xnor U15556 (N_15556,N_15403,N_15320);
or U15557 (N_15557,N_15393,N_15368);
nand U15558 (N_15558,N_15385,N_15406);
nand U15559 (N_15559,N_15314,N_15401);
and U15560 (N_15560,N_15327,N_15449);
or U15561 (N_15561,N_15494,N_15377);
nand U15562 (N_15562,N_15464,N_15346);
and U15563 (N_15563,N_15420,N_15369);
nand U15564 (N_15564,N_15460,N_15427);
or U15565 (N_15565,N_15328,N_15279);
nor U15566 (N_15566,N_15479,N_15363);
xor U15567 (N_15567,N_15257,N_15430);
nand U15568 (N_15568,N_15411,N_15397);
xnor U15569 (N_15569,N_15474,N_15292);
xnor U15570 (N_15570,N_15451,N_15318);
and U15571 (N_15571,N_15384,N_15299);
nand U15572 (N_15572,N_15251,N_15277);
nand U15573 (N_15573,N_15339,N_15469);
nor U15574 (N_15574,N_15358,N_15431);
xor U15575 (N_15575,N_15475,N_15336);
or U15576 (N_15576,N_15472,N_15271);
nor U15577 (N_15577,N_15386,N_15445);
nand U15578 (N_15578,N_15353,N_15373);
and U15579 (N_15579,N_15417,N_15421);
or U15580 (N_15580,N_15283,N_15455);
nor U15581 (N_15581,N_15342,N_15261);
nand U15582 (N_15582,N_15316,N_15324);
nor U15583 (N_15583,N_15361,N_15453);
nor U15584 (N_15584,N_15272,N_15429);
nor U15585 (N_15585,N_15325,N_15259);
or U15586 (N_15586,N_15344,N_15398);
nand U15587 (N_15587,N_15440,N_15366);
nor U15588 (N_15588,N_15450,N_15372);
xnor U15589 (N_15589,N_15446,N_15355);
nand U15590 (N_15590,N_15428,N_15274);
or U15591 (N_15591,N_15253,N_15438);
nor U15592 (N_15592,N_15313,N_15370);
nand U15593 (N_15593,N_15498,N_15291);
and U15594 (N_15594,N_15382,N_15376);
or U15595 (N_15595,N_15362,N_15262);
nor U15596 (N_15596,N_15343,N_15293);
and U15597 (N_15597,N_15250,N_15338);
nor U15598 (N_15598,N_15329,N_15423);
or U15599 (N_15599,N_15332,N_15305);
nor U15600 (N_15600,N_15350,N_15482);
nor U15601 (N_15601,N_15341,N_15330);
nor U15602 (N_15602,N_15334,N_15389);
nand U15603 (N_15603,N_15484,N_15356);
or U15604 (N_15604,N_15424,N_15410);
nor U15605 (N_15605,N_15348,N_15473);
or U15606 (N_15606,N_15315,N_15390);
xor U15607 (N_15607,N_15478,N_15492);
nor U15608 (N_15608,N_15392,N_15379);
or U15609 (N_15609,N_15354,N_15486);
xor U15610 (N_15610,N_15466,N_15331);
xor U15611 (N_15611,N_15319,N_15340);
xnor U15612 (N_15612,N_15414,N_15290);
nand U15613 (N_15613,N_15359,N_15402);
nor U15614 (N_15614,N_15310,N_15269);
nor U15615 (N_15615,N_15380,N_15467);
and U15616 (N_15616,N_15288,N_15287);
or U15617 (N_15617,N_15304,N_15297);
and U15618 (N_15618,N_15415,N_15480);
and U15619 (N_15619,N_15436,N_15391);
nand U15620 (N_15620,N_15335,N_15311);
nor U15621 (N_15621,N_15270,N_15307);
nand U15622 (N_15622,N_15439,N_15364);
nand U15623 (N_15623,N_15371,N_15365);
and U15624 (N_15624,N_15345,N_15452);
xnor U15625 (N_15625,N_15291,N_15330);
and U15626 (N_15626,N_15321,N_15273);
nand U15627 (N_15627,N_15403,N_15462);
and U15628 (N_15628,N_15421,N_15483);
nor U15629 (N_15629,N_15425,N_15279);
and U15630 (N_15630,N_15367,N_15384);
or U15631 (N_15631,N_15308,N_15287);
or U15632 (N_15632,N_15381,N_15278);
xor U15633 (N_15633,N_15423,N_15364);
and U15634 (N_15634,N_15251,N_15473);
and U15635 (N_15635,N_15363,N_15288);
nor U15636 (N_15636,N_15418,N_15401);
nand U15637 (N_15637,N_15419,N_15317);
and U15638 (N_15638,N_15356,N_15438);
xor U15639 (N_15639,N_15451,N_15299);
and U15640 (N_15640,N_15423,N_15321);
xor U15641 (N_15641,N_15405,N_15474);
nand U15642 (N_15642,N_15453,N_15475);
nand U15643 (N_15643,N_15415,N_15391);
nor U15644 (N_15644,N_15380,N_15313);
and U15645 (N_15645,N_15455,N_15301);
xor U15646 (N_15646,N_15374,N_15378);
xnor U15647 (N_15647,N_15346,N_15474);
and U15648 (N_15648,N_15499,N_15456);
nand U15649 (N_15649,N_15376,N_15264);
or U15650 (N_15650,N_15426,N_15393);
xnor U15651 (N_15651,N_15310,N_15314);
or U15652 (N_15652,N_15482,N_15469);
xor U15653 (N_15653,N_15272,N_15288);
xnor U15654 (N_15654,N_15392,N_15345);
and U15655 (N_15655,N_15457,N_15455);
and U15656 (N_15656,N_15430,N_15301);
nor U15657 (N_15657,N_15267,N_15280);
xor U15658 (N_15658,N_15381,N_15496);
nand U15659 (N_15659,N_15281,N_15458);
xor U15660 (N_15660,N_15401,N_15438);
nor U15661 (N_15661,N_15405,N_15305);
or U15662 (N_15662,N_15387,N_15281);
and U15663 (N_15663,N_15300,N_15479);
and U15664 (N_15664,N_15406,N_15428);
xnor U15665 (N_15665,N_15337,N_15308);
or U15666 (N_15666,N_15324,N_15291);
xnor U15667 (N_15667,N_15325,N_15294);
nor U15668 (N_15668,N_15420,N_15385);
nand U15669 (N_15669,N_15445,N_15291);
nand U15670 (N_15670,N_15264,N_15418);
nor U15671 (N_15671,N_15288,N_15368);
or U15672 (N_15672,N_15271,N_15426);
xnor U15673 (N_15673,N_15281,N_15452);
and U15674 (N_15674,N_15358,N_15424);
and U15675 (N_15675,N_15282,N_15294);
nand U15676 (N_15676,N_15276,N_15401);
nor U15677 (N_15677,N_15391,N_15331);
or U15678 (N_15678,N_15282,N_15412);
or U15679 (N_15679,N_15411,N_15492);
nand U15680 (N_15680,N_15270,N_15496);
nand U15681 (N_15681,N_15359,N_15343);
or U15682 (N_15682,N_15274,N_15486);
nor U15683 (N_15683,N_15440,N_15374);
nor U15684 (N_15684,N_15455,N_15492);
xnor U15685 (N_15685,N_15470,N_15495);
nor U15686 (N_15686,N_15275,N_15259);
nand U15687 (N_15687,N_15264,N_15379);
or U15688 (N_15688,N_15255,N_15328);
xnor U15689 (N_15689,N_15484,N_15488);
nor U15690 (N_15690,N_15458,N_15348);
or U15691 (N_15691,N_15369,N_15275);
or U15692 (N_15692,N_15359,N_15451);
xor U15693 (N_15693,N_15298,N_15329);
xnor U15694 (N_15694,N_15275,N_15341);
or U15695 (N_15695,N_15358,N_15252);
nand U15696 (N_15696,N_15339,N_15460);
nor U15697 (N_15697,N_15335,N_15366);
or U15698 (N_15698,N_15423,N_15485);
xor U15699 (N_15699,N_15449,N_15346);
xnor U15700 (N_15700,N_15265,N_15417);
nor U15701 (N_15701,N_15418,N_15466);
or U15702 (N_15702,N_15296,N_15446);
nor U15703 (N_15703,N_15456,N_15266);
or U15704 (N_15704,N_15466,N_15478);
and U15705 (N_15705,N_15255,N_15483);
nor U15706 (N_15706,N_15489,N_15283);
nand U15707 (N_15707,N_15362,N_15432);
or U15708 (N_15708,N_15386,N_15337);
nand U15709 (N_15709,N_15309,N_15307);
xnor U15710 (N_15710,N_15272,N_15352);
or U15711 (N_15711,N_15459,N_15294);
and U15712 (N_15712,N_15357,N_15482);
and U15713 (N_15713,N_15319,N_15430);
or U15714 (N_15714,N_15311,N_15347);
nor U15715 (N_15715,N_15269,N_15378);
or U15716 (N_15716,N_15374,N_15292);
nand U15717 (N_15717,N_15321,N_15454);
or U15718 (N_15718,N_15378,N_15300);
and U15719 (N_15719,N_15407,N_15442);
xor U15720 (N_15720,N_15346,N_15424);
and U15721 (N_15721,N_15453,N_15458);
or U15722 (N_15722,N_15315,N_15477);
or U15723 (N_15723,N_15355,N_15321);
nor U15724 (N_15724,N_15406,N_15278);
nor U15725 (N_15725,N_15372,N_15409);
or U15726 (N_15726,N_15406,N_15422);
nor U15727 (N_15727,N_15257,N_15292);
and U15728 (N_15728,N_15275,N_15299);
xnor U15729 (N_15729,N_15337,N_15460);
nor U15730 (N_15730,N_15376,N_15381);
or U15731 (N_15731,N_15272,N_15422);
nor U15732 (N_15732,N_15419,N_15435);
xnor U15733 (N_15733,N_15449,N_15337);
or U15734 (N_15734,N_15300,N_15310);
xor U15735 (N_15735,N_15436,N_15489);
nor U15736 (N_15736,N_15358,N_15286);
or U15737 (N_15737,N_15440,N_15491);
xor U15738 (N_15738,N_15446,N_15482);
xnor U15739 (N_15739,N_15420,N_15307);
or U15740 (N_15740,N_15282,N_15391);
xnor U15741 (N_15741,N_15375,N_15472);
or U15742 (N_15742,N_15420,N_15450);
nand U15743 (N_15743,N_15277,N_15381);
nor U15744 (N_15744,N_15312,N_15494);
xor U15745 (N_15745,N_15307,N_15423);
and U15746 (N_15746,N_15475,N_15356);
or U15747 (N_15747,N_15449,N_15279);
or U15748 (N_15748,N_15325,N_15293);
and U15749 (N_15749,N_15437,N_15280);
xor U15750 (N_15750,N_15606,N_15532);
nor U15751 (N_15751,N_15506,N_15738);
or U15752 (N_15752,N_15740,N_15674);
nor U15753 (N_15753,N_15624,N_15646);
nand U15754 (N_15754,N_15745,N_15502);
xnor U15755 (N_15755,N_15693,N_15523);
and U15756 (N_15756,N_15656,N_15650);
or U15757 (N_15757,N_15635,N_15616);
xor U15758 (N_15758,N_15726,N_15552);
xnor U15759 (N_15759,N_15717,N_15588);
and U15760 (N_15760,N_15632,N_15556);
xor U15761 (N_15761,N_15739,N_15682);
nand U15762 (N_15762,N_15633,N_15603);
or U15763 (N_15763,N_15659,N_15602);
or U15764 (N_15764,N_15510,N_15694);
nand U15765 (N_15765,N_15539,N_15604);
or U15766 (N_15766,N_15504,N_15714);
and U15767 (N_15767,N_15695,N_15660);
and U15768 (N_15768,N_15541,N_15508);
nor U15769 (N_15769,N_15654,N_15550);
xor U15770 (N_15770,N_15645,N_15651);
or U15771 (N_15771,N_15628,N_15696);
xor U15772 (N_15772,N_15505,N_15689);
or U15773 (N_15773,N_15643,N_15546);
or U15774 (N_15774,N_15509,N_15743);
or U15775 (N_15775,N_15730,N_15615);
nand U15776 (N_15776,N_15573,N_15563);
and U15777 (N_15777,N_15585,N_15749);
nand U15778 (N_15778,N_15511,N_15564);
nand U15779 (N_15779,N_15710,N_15720);
nor U15780 (N_15780,N_15538,N_15529);
or U15781 (N_15781,N_15637,N_15562);
nor U15782 (N_15782,N_15512,N_15549);
xnor U15783 (N_15783,N_15702,N_15697);
nor U15784 (N_15784,N_15680,N_15729);
nand U15785 (N_15785,N_15568,N_15578);
xnor U15786 (N_15786,N_15727,N_15566);
nand U15787 (N_15787,N_15600,N_15630);
xor U15788 (N_15788,N_15589,N_15705);
nor U15789 (N_15789,N_15609,N_15707);
or U15790 (N_15790,N_15676,N_15690);
nand U15791 (N_15791,N_15531,N_15692);
nand U15792 (N_15792,N_15734,N_15728);
nand U15793 (N_15793,N_15594,N_15537);
xnor U15794 (N_15794,N_15618,N_15548);
or U15795 (N_15795,N_15547,N_15518);
and U15796 (N_15796,N_15642,N_15742);
nand U15797 (N_15797,N_15555,N_15699);
and U15798 (N_15798,N_15688,N_15669);
xor U15799 (N_15799,N_15744,N_15653);
nand U15800 (N_15800,N_15735,N_15583);
and U15801 (N_15801,N_15587,N_15601);
nor U15802 (N_15802,N_15647,N_15672);
and U15803 (N_15803,N_15535,N_15686);
and U15804 (N_15804,N_15684,N_15747);
nand U15805 (N_15805,N_15652,N_15617);
and U15806 (N_15806,N_15644,N_15698);
xnor U15807 (N_15807,N_15599,N_15677);
or U15808 (N_15808,N_15675,N_15554);
or U15809 (N_15809,N_15596,N_15703);
xnor U15810 (N_15810,N_15716,N_15526);
xnor U15811 (N_15811,N_15673,N_15608);
and U15812 (N_15812,N_15691,N_15700);
xor U15813 (N_15813,N_15513,N_15634);
nor U15814 (N_15814,N_15607,N_15665);
nor U15815 (N_15815,N_15721,N_15520);
or U15816 (N_15816,N_15528,N_15576);
or U15817 (N_15817,N_15595,N_15517);
nor U15818 (N_15818,N_15515,N_15641);
nor U15819 (N_15819,N_15663,N_15725);
or U15820 (N_15820,N_15557,N_15706);
or U15821 (N_15821,N_15649,N_15575);
and U15822 (N_15822,N_15558,N_15519);
nor U15823 (N_15823,N_15620,N_15522);
xnor U15824 (N_15824,N_15561,N_15621);
nor U15825 (N_15825,N_15670,N_15627);
nor U15826 (N_15826,N_15708,N_15683);
xor U15827 (N_15827,N_15590,N_15500);
xnor U15828 (N_15828,N_15521,N_15533);
or U15829 (N_15829,N_15638,N_15732);
nor U15830 (N_15830,N_15733,N_15605);
and U15831 (N_15831,N_15625,N_15619);
and U15832 (N_15832,N_15613,N_15636);
nand U15833 (N_15833,N_15543,N_15525);
and U15834 (N_15834,N_15681,N_15661);
nand U15835 (N_15835,N_15580,N_15724);
or U15836 (N_15836,N_15569,N_15584);
and U15837 (N_15837,N_15524,N_15722);
and U15838 (N_15838,N_15639,N_15551);
and U15839 (N_15839,N_15614,N_15597);
or U15840 (N_15840,N_15567,N_15553);
xor U15841 (N_15841,N_15540,N_15593);
and U15842 (N_15842,N_15516,N_15657);
nor U15843 (N_15843,N_15623,N_15741);
and U15844 (N_15844,N_15582,N_15542);
and U15845 (N_15845,N_15592,N_15711);
xnor U15846 (N_15846,N_15612,N_15704);
nand U15847 (N_15847,N_15679,N_15577);
or U15848 (N_15848,N_15640,N_15530);
xor U15849 (N_15849,N_15514,N_15737);
xor U15850 (N_15850,N_15668,N_15622);
nand U15851 (N_15851,N_15713,N_15545);
nand U15852 (N_15852,N_15671,N_15591);
or U15853 (N_15853,N_15678,N_15565);
nor U15854 (N_15854,N_15610,N_15662);
nand U15855 (N_15855,N_15559,N_15648);
nand U15856 (N_15856,N_15574,N_15746);
nor U15857 (N_15857,N_15701,N_15571);
nand U15858 (N_15858,N_15598,N_15685);
and U15859 (N_15859,N_15507,N_15736);
nor U15860 (N_15860,N_15723,N_15631);
xnor U15861 (N_15861,N_15712,N_15658);
nor U15862 (N_15862,N_15687,N_15664);
and U15863 (N_15863,N_15536,N_15748);
xnor U15864 (N_15864,N_15544,N_15560);
xor U15865 (N_15865,N_15503,N_15579);
and U15866 (N_15866,N_15666,N_15667);
or U15867 (N_15867,N_15534,N_15626);
or U15868 (N_15868,N_15572,N_15719);
or U15869 (N_15869,N_15718,N_15586);
or U15870 (N_15870,N_15581,N_15527);
and U15871 (N_15871,N_15655,N_15715);
and U15872 (N_15872,N_15501,N_15570);
nor U15873 (N_15873,N_15709,N_15611);
nor U15874 (N_15874,N_15731,N_15629);
nand U15875 (N_15875,N_15660,N_15724);
and U15876 (N_15876,N_15549,N_15574);
nor U15877 (N_15877,N_15605,N_15639);
nor U15878 (N_15878,N_15692,N_15712);
nor U15879 (N_15879,N_15678,N_15579);
nor U15880 (N_15880,N_15598,N_15642);
nor U15881 (N_15881,N_15665,N_15508);
nor U15882 (N_15882,N_15660,N_15708);
xnor U15883 (N_15883,N_15579,N_15727);
xnor U15884 (N_15884,N_15713,N_15544);
and U15885 (N_15885,N_15537,N_15547);
or U15886 (N_15886,N_15681,N_15570);
and U15887 (N_15887,N_15578,N_15686);
or U15888 (N_15888,N_15693,N_15640);
or U15889 (N_15889,N_15578,N_15605);
nand U15890 (N_15890,N_15555,N_15549);
and U15891 (N_15891,N_15560,N_15605);
and U15892 (N_15892,N_15681,N_15554);
and U15893 (N_15893,N_15734,N_15737);
or U15894 (N_15894,N_15668,N_15539);
nand U15895 (N_15895,N_15643,N_15594);
or U15896 (N_15896,N_15510,N_15530);
and U15897 (N_15897,N_15684,N_15659);
xor U15898 (N_15898,N_15572,N_15594);
nor U15899 (N_15899,N_15637,N_15740);
and U15900 (N_15900,N_15519,N_15556);
and U15901 (N_15901,N_15637,N_15615);
nor U15902 (N_15902,N_15614,N_15579);
nor U15903 (N_15903,N_15633,N_15597);
nor U15904 (N_15904,N_15734,N_15678);
and U15905 (N_15905,N_15659,N_15726);
or U15906 (N_15906,N_15683,N_15723);
nor U15907 (N_15907,N_15608,N_15658);
xnor U15908 (N_15908,N_15586,N_15623);
or U15909 (N_15909,N_15595,N_15596);
nor U15910 (N_15910,N_15704,N_15638);
nor U15911 (N_15911,N_15700,N_15555);
xnor U15912 (N_15912,N_15678,N_15716);
and U15913 (N_15913,N_15640,N_15573);
and U15914 (N_15914,N_15642,N_15575);
or U15915 (N_15915,N_15530,N_15735);
nand U15916 (N_15916,N_15587,N_15654);
nor U15917 (N_15917,N_15624,N_15603);
or U15918 (N_15918,N_15510,N_15534);
nand U15919 (N_15919,N_15597,N_15552);
and U15920 (N_15920,N_15740,N_15634);
and U15921 (N_15921,N_15556,N_15660);
nor U15922 (N_15922,N_15566,N_15615);
or U15923 (N_15923,N_15579,N_15572);
and U15924 (N_15924,N_15658,N_15538);
and U15925 (N_15925,N_15666,N_15583);
xor U15926 (N_15926,N_15639,N_15618);
and U15927 (N_15927,N_15541,N_15722);
and U15928 (N_15928,N_15735,N_15548);
or U15929 (N_15929,N_15523,N_15740);
nand U15930 (N_15930,N_15516,N_15602);
and U15931 (N_15931,N_15500,N_15688);
nor U15932 (N_15932,N_15737,N_15741);
nor U15933 (N_15933,N_15652,N_15546);
nor U15934 (N_15934,N_15551,N_15620);
and U15935 (N_15935,N_15730,N_15560);
nor U15936 (N_15936,N_15664,N_15676);
xnor U15937 (N_15937,N_15573,N_15557);
nor U15938 (N_15938,N_15583,N_15545);
nand U15939 (N_15939,N_15656,N_15581);
nand U15940 (N_15940,N_15722,N_15728);
nor U15941 (N_15941,N_15572,N_15544);
nand U15942 (N_15942,N_15554,N_15672);
nand U15943 (N_15943,N_15691,N_15749);
and U15944 (N_15944,N_15515,N_15518);
nand U15945 (N_15945,N_15663,N_15735);
nand U15946 (N_15946,N_15742,N_15588);
nor U15947 (N_15947,N_15624,N_15735);
xnor U15948 (N_15948,N_15725,N_15651);
or U15949 (N_15949,N_15575,N_15590);
or U15950 (N_15950,N_15741,N_15722);
and U15951 (N_15951,N_15658,N_15522);
and U15952 (N_15952,N_15618,N_15704);
and U15953 (N_15953,N_15636,N_15573);
or U15954 (N_15954,N_15735,N_15635);
nand U15955 (N_15955,N_15749,N_15566);
nand U15956 (N_15956,N_15748,N_15631);
and U15957 (N_15957,N_15605,N_15745);
nor U15958 (N_15958,N_15697,N_15741);
nand U15959 (N_15959,N_15694,N_15708);
xnor U15960 (N_15960,N_15610,N_15749);
or U15961 (N_15961,N_15727,N_15648);
nand U15962 (N_15962,N_15543,N_15694);
nand U15963 (N_15963,N_15575,N_15604);
nand U15964 (N_15964,N_15531,N_15743);
nand U15965 (N_15965,N_15646,N_15737);
nor U15966 (N_15966,N_15567,N_15609);
xnor U15967 (N_15967,N_15591,N_15727);
xor U15968 (N_15968,N_15532,N_15665);
nor U15969 (N_15969,N_15683,N_15641);
xor U15970 (N_15970,N_15677,N_15610);
and U15971 (N_15971,N_15637,N_15628);
nor U15972 (N_15972,N_15570,N_15592);
or U15973 (N_15973,N_15686,N_15659);
or U15974 (N_15974,N_15541,N_15637);
nor U15975 (N_15975,N_15737,N_15569);
and U15976 (N_15976,N_15681,N_15510);
nor U15977 (N_15977,N_15535,N_15646);
and U15978 (N_15978,N_15592,N_15633);
or U15979 (N_15979,N_15515,N_15748);
xor U15980 (N_15980,N_15700,N_15719);
nor U15981 (N_15981,N_15569,N_15554);
and U15982 (N_15982,N_15648,N_15529);
or U15983 (N_15983,N_15699,N_15505);
nor U15984 (N_15984,N_15642,N_15701);
nand U15985 (N_15985,N_15658,N_15505);
and U15986 (N_15986,N_15537,N_15688);
xnor U15987 (N_15987,N_15564,N_15720);
nand U15988 (N_15988,N_15564,N_15684);
or U15989 (N_15989,N_15559,N_15639);
xnor U15990 (N_15990,N_15567,N_15508);
and U15991 (N_15991,N_15519,N_15719);
and U15992 (N_15992,N_15715,N_15677);
or U15993 (N_15993,N_15533,N_15537);
or U15994 (N_15994,N_15662,N_15571);
or U15995 (N_15995,N_15503,N_15673);
nand U15996 (N_15996,N_15540,N_15569);
nor U15997 (N_15997,N_15593,N_15628);
xor U15998 (N_15998,N_15519,N_15557);
nor U15999 (N_15999,N_15556,N_15524);
nand U16000 (N_16000,N_15926,N_15750);
xnor U16001 (N_16001,N_15843,N_15848);
nand U16002 (N_16002,N_15970,N_15900);
or U16003 (N_16003,N_15946,N_15813);
and U16004 (N_16004,N_15937,N_15863);
xnor U16005 (N_16005,N_15763,N_15780);
xnor U16006 (N_16006,N_15940,N_15807);
nand U16007 (N_16007,N_15927,N_15952);
and U16008 (N_16008,N_15822,N_15767);
or U16009 (N_16009,N_15985,N_15845);
nor U16010 (N_16010,N_15886,N_15999);
and U16011 (N_16011,N_15989,N_15849);
nand U16012 (N_16012,N_15768,N_15980);
or U16013 (N_16013,N_15800,N_15953);
xor U16014 (N_16014,N_15933,N_15788);
xnor U16015 (N_16015,N_15932,N_15955);
xnor U16016 (N_16016,N_15973,N_15760);
or U16017 (N_16017,N_15784,N_15819);
nand U16018 (N_16018,N_15797,N_15809);
nand U16019 (N_16019,N_15770,N_15778);
xnor U16020 (N_16020,N_15939,N_15846);
or U16021 (N_16021,N_15979,N_15816);
xor U16022 (N_16022,N_15850,N_15918);
nand U16023 (N_16023,N_15908,N_15917);
xor U16024 (N_16024,N_15976,N_15892);
and U16025 (N_16025,N_15839,N_15798);
and U16026 (N_16026,N_15995,N_15988);
nand U16027 (N_16027,N_15752,N_15837);
nor U16028 (N_16028,N_15875,N_15975);
xor U16029 (N_16029,N_15823,N_15847);
or U16030 (N_16030,N_15872,N_15907);
xnor U16031 (N_16031,N_15965,N_15925);
xnor U16032 (N_16032,N_15966,N_15934);
and U16033 (N_16033,N_15873,N_15827);
nand U16034 (N_16034,N_15777,N_15916);
or U16035 (N_16035,N_15758,N_15877);
or U16036 (N_16036,N_15783,N_15832);
nor U16037 (N_16037,N_15992,N_15874);
xnor U16038 (N_16038,N_15781,N_15885);
xnor U16039 (N_16039,N_15864,N_15901);
and U16040 (N_16040,N_15785,N_15817);
xnor U16041 (N_16041,N_15844,N_15757);
nand U16042 (N_16042,N_15812,N_15782);
nand U16043 (N_16043,N_15871,N_15861);
or U16044 (N_16044,N_15990,N_15876);
nor U16045 (N_16045,N_15870,N_15968);
and U16046 (N_16046,N_15942,N_15754);
and U16047 (N_16047,N_15772,N_15801);
and U16048 (N_16048,N_15759,N_15997);
nor U16049 (N_16049,N_15944,N_15841);
xnor U16050 (N_16050,N_15821,N_15833);
xor U16051 (N_16051,N_15826,N_15924);
nand U16052 (N_16052,N_15906,N_15789);
and U16053 (N_16053,N_15806,N_15804);
nand U16054 (N_16054,N_15824,N_15792);
and U16055 (N_16055,N_15972,N_15795);
and U16056 (N_16056,N_15862,N_15967);
nand U16057 (N_16057,N_15909,N_15775);
xnor U16058 (N_16058,N_15854,N_15828);
or U16059 (N_16059,N_15962,N_15912);
nand U16060 (N_16060,N_15830,N_15765);
and U16061 (N_16061,N_15774,N_15884);
and U16062 (N_16062,N_15919,N_15954);
xor U16063 (N_16063,N_15762,N_15882);
nor U16064 (N_16064,N_15779,N_15755);
nor U16065 (N_16065,N_15829,N_15898);
or U16066 (N_16066,N_15996,N_15982);
and U16067 (N_16067,N_15974,N_15959);
nand U16068 (N_16068,N_15814,N_15984);
xor U16069 (N_16069,N_15950,N_15805);
nor U16070 (N_16070,N_15981,N_15834);
nand U16071 (N_16071,N_15978,N_15856);
nor U16072 (N_16072,N_15904,N_15914);
xnor U16073 (N_16073,N_15929,N_15969);
or U16074 (N_16074,N_15986,N_15935);
or U16075 (N_16075,N_15931,N_15991);
and U16076 (N_16076,N_15913,N_15949);
or U16077 (N_16077,N_15897,N_15887);
and U16078 (N_16078,N_15868,N_15756);
xor U16079 (N_16079,N_15960,N_15936);
or U16080 (N_16080,N_15853,N_15920);
nor U16081 (N_16081,N_15889,N_15851);
xor U16082 (N_16082,N_15771,N_15857);
xor U16083 (N_16083,N_15825,N_15852);
xor U16084 (N_16084,N_15793,N_15893);
nor U16085 (N_16085,N_15958,N_15859);
xor U16086 (N_16086,N_15855,N_15860);
nand U16087 (N_16087,N_15842,N_15983);
xnor U16088 (N_16088,N_15803,N_15956);
xor U16089 (N_16089,N_15815,N_15977);
xnor U16090 (N_16090,N_15891,N_15883);
or U16091 (N_16091,N_15987,N_15769);
xnor U16092 (N_16092,N_15796,N_15880);
xnor U16093 (N_16093,N_15776,N_15894);
and U16094 (N_16094,N_15888,N_15971);
nor U16095 (N_16095,N_15911,N_15895);
nand U16096 (N_16096,N_15964,N_15896);
xnor U16097 (N_16097,N_15902,N_15947);
nor U16098 (N_16098,N_15836,N_15790);
or U16099 (N_16099,N_15957,N_15951);
nor U16100 (N_16100,N_15766,N_15961);
and U16101 (N_16101,N_15903,N_15879);
nor U16102 (N_16102,N_15773,N_15963);
and U16103 (N_16103,N_15921,N_15865);
or U16104 (N_16104,N_15791,N_15802);
xnor U16105 (N_16105,N_15787,N_15835);
nor U16106 (N_16106,N_15878,N_15993);
xor U16107 (N_16107,N_15923,N_15881);
and U16108 (N_16108,N_15867,N_15808);
and U16109 (N_16109,N_15905,N_15998);
xor U16110 (N_16110,N_15810,N_15943);
and U16111 (N_16111,N_15840,N_15930);
nor U16112 (N_16112,N_15866,N_15751);
nor U16113 (N_16113,N_15794,N_15818);
nand U16114 (N_16114,N_15948,N_15820);
nor U16115 (N_16115,N_15811,N_15890);
nand U16116 (N_16116,N_15941,N_15753);
xor U16117 (N_16117,N_15831,N_15928);
and U16118 (N_16118,N_15922,N_15786);
xnor U16119 (N_16119,N_15910,N_15838);
xnor U16120 (N_16120,N_15869,N_15799);
and U16121 (N_16121,N_15764,N_15915);
xor U16122 (N_16122,N_15858,N_15761);
and U16123 (N_16123,N_15899,N_15938);
or U16124 (N_16124,N_15945,N_15994);
xor U16125 (N_16125,N_15752,N_15961);
nor U16126 (N_16126,N_15981,N_15816);
xor U16127 (N_16127,N_15777,N_15902);
nor U16128 (N_16128,N_15823,N_15879);
nor U16129 (N_16129,N_15946,N_15993);
nor U16130 (N_16130,N_15917,N_15963);
nor U16131 (N_16131,N_15909,N_15818);
nand U16132 (N_16132,N_15967,N_15988);
and U16133 (N_16133,N_15965,N_15904);
xnor U16134 (N_16134,N_15860,N_15937);
and U16135 (N_16135,N_15919,N_15917);
xnor U16136 (N_16136,N_15840,N_15897);
or U16137 (N_16137,N_15799,N_15809);
and U16138 (N_16138,N_15961,N_15783);
nand U16139 (N_16139,N_15826,N_15871);
or U16140 (N_16140,N_15852,N_15774);
or U16141 (N_16141,N_15765,N_15774);
nor U16142 (N_16142,N_15762,N_15920);
and U16143 (N_16143,N_15795,N_15942);
nand U16144 (N_16144,N_15768,N_15971);
nand U16145 (N_16145,N_15780,N_15860);
nand U16146 (N_16146,N_15832,N_15964);
xnor U16147 (N_16147,N_15995,N_15784);
nor U16148 (N_16148,N_15936,N_15996);
nand U16149 (N_16149,N_15925,N_15932);
and U16150 (N_16150,N_15878,N_15824);
nand U16151 (N_16151,N_15827,N_15912);
nor U16152 (N_16152,N_15762,N_15804);
nand U16153 (N_16153,N_15785,N_15821);
nand U16154 (N_16154,N_15752,N_15827);
or U16155 (N_16155,N_15949,N_15854);
or U16156 (N_16156,N_15907,N_15999);
or U16157 (N_16157,N_15832,N_15895);
and U16158 (N_16158,N_15851,N_15770);
nand U16159 (N_16159,N_15884,N_15805);
and U16160 (N_16160,N_15939,N_15873);
or U16161 (N_16161,N_15777,N_15899);
or U16162 (N_16162,N_15769,N_15953);
nor U16163 (N_16163,N_15982,N_15942);
xor U16164 (N_16164,N_15959,N_15874);
and U16165 (N_16165,N_15968,N_15920);
or U16166 (N_16166,N_15943,N_15946);
xor U16167 (N_16167,N_15797,N_15857);
nor U16168 (N_16168,N_15864,N_15777);
xnor U16169 (N_16169,N_15975,N_15913);
or U16170 (N_16170,N_15871,N_15929);
and U16171 (N_16171,N_15763,N_15839);
nand U16172 (N_16172,N_15959,N_15912);
xnor U16173 (N_16173,N_15873,N_15879);
nand U16174 (N_16174,N_15894,N_15809);
nor U16175 (N_16175,N_15888,N_15779);
or U16176 (N_16176,N_15924,N_15754);
xnor U16177 (N_16177,N_15979,N_15752);
or U16178 (N_16178,N_15830,N_15981);
xor U16179 (N_16179,N_15859,N_15973);
xnor U16180 (N_16180,N_15868,N_15998);
nor U16181 (N_16181,N_15949,N_15818);
nand U16182 (N_16182,N_15819,N_15837);
xor U16183 (N_16183,N_15859,N_15962);
and U16184 (N_16184,N_15963,N_15931);
nor U16185 (N_16185,N_15855,N_15937);
and U16186 (N_16186,N_15996,N_15931);
nor U16187 (N_16187,N_15881,N_15831);
nand U16188 (N_16188,N_15830,N_15935);
and U16189 (N_16189,N_15953,N_15992);
nor U16190 (N_16190,N_15939,N_15756);
and U16191 (N_16191,N_15846,N_15802);
nand U16192 (N_16192,N_15915,N_15992);
or U16193 (N_16193,N_15770,N_15875);
or U16194 (N_16194,N_15801,N_15754);
or U16195 (N_16195,N_15959,N_15804);
and U16196 (N_16196,N_15953,N_15811);
xnor U16197 (N_16197,N_15914,N_15779);
or U16198 (N_16198,N_15979,N_15955);
and U16199 (N_16199,N_15818,N_15903);
xnor U16200 (N_16200,N_15849,N_15951);
nand U16201 (N_16201,N_15841,N_15815);
xor U16202 (N_16202,N_15855,N_15783);
nand U16203 (N_16203,N_15849,N_15775);
or U16204 (N_16204,N_15899,N_15936);
xor U16205 (N_16205,N_15987,N_15855);
xnor U16206 (N_16206,N_15770,N_15880);
and U16207 (N_16207,N_15932,N_15959);
xor U16208 (N_16208,N_15949,N_15758);
or U16209 (N_16209,N_15926,N_15784);
nand U16210 (N_16210,N_15948,N_15797);
xor U16211 (N_16211,N_15997,N_15978);
nand U16212 (N_16212,N_15816,N_15788);
nor U16213 (N_16213,N_15946,N_15882);
and U16214 (N_16214,N_15961,N_15784);
nor U16215 (N_16215,N_15753,N_15907);
nor U16216 (N_16216,N_15790,N_15851);
or U16217 (N_16217,N_15846,N_15961);
nor U16218 (N_16218,N_15974,N_15821);
nor U16219 (N_16219,N_15931,N_15982);
or U16220 (N_16220,N_15750,N_15846);
xor U16221 (N_16221,N_15830,N_15797);
or U16222 (N_16222,N_15862,N_15899);
nor U16223 (N_16223,N_15972,N_15861);
nor U16224 (N_16224,N_15886,N_15807);
and U16225 (N_16225,N_15790,N_15974);
xnor U16226 (N_16226,N_15982,N_15950);
nor U16227 (N_16227,N_15989,N_15851);
and U16228 (N_16228,N_15865,N_15769);
nand U16229 (N_16229,N_15878,N_15882);
nand U16230 (N_16230,N_15807,N_15908);
xor U16231 (N_16231,N_15968,N_15837);
nor U16232 (N_16232,N_15919,N_15786);
nand U16233 (N_16233,N_15866,N_15993);
xor U16234 (N_16234,N_15884,N_15862);
and U16235 (N_16235,N_15900,N_15801);
and U16236 (N_16236,N_15955,N_15909);
nor U16237 (N_16237,N_15815,N_15931);
xnor U16238 (N_16238,N_15906,N_15818);
and U16239 (N_16239,N_15929,N_15752);
or U16240 (N_16240,N_15857,N_15861);
xor U16241 (N_16241,N_15798,N_15827);
nor U16242 (N_16242,N_15954,N_15985);
nand U16243 (N_16243,N_15797,N_15776);
xor U16244 (N_16244,N_15768,N_15841);
or U16245 (N_16245,N_15849,N_15860);
nand U16246 (N_16246,N_15761,N_15830);
or U16247 (N_16247,N_15968,N_15781);
xor U16248 (N_16248,N_15822,N_15979);
xor U16249 (N_16249,N_15898,N_15867);
nand U16250 (N_16250,N_16003,N_16165);
nor U16251 (N_16251,N_16072,N_16023);
and U16252 (N_16252,N_16224,N_16062);
or U16253 (N_16253,N_16210,N_16092);
or U16254 (N_16254,N_16087,N_16235);
or U16255 (N_16255,N_16083,N_16058);
nand U16256 (N_16256,N_16216,N_16007);
and U16257 (N_16257,N_16021,N_16155);
nand U16258 (N_16258,N_16115,N_16154);
nand U16259 (N_16259,N_16002,N_16212);
nand U16260 (N_16260,N_16242,N_16071);
nor U16261 (N_16261,N_16042,N_16167);
xnor U16262 (N_16262,N_16215,N_16075);
or U16263 (N_16263,N_16031,N_16022);
and U16264 (N_16264,N_16001,N_16059);
and U16265 (N_16265,N_16117,N_16178);
nor U16266 (N_16266,N_16009,N_16151);
xor U16267 (N_16267,N_16146,N_16027);
nor U16268 (N_16268,N_16140,N_16056);
nand U16269 (N_16269,N_16012,N_16202);
nor U16270 (N_16270,N_16116,N_16095);
nor U16271 (N_16271,N_16109,N_16104);
xnor U16272 (N_16272,N_16247,N_16111);
nand U16273 (N_16273,N_16190,N_16240);
nand U16274 (N_16274,N_16160,N_16137);
nor U16275 (N_16275,N_16051,N_16166);
or U16276 (N_16276,N_16054,N_16123);
nor U16277 (N_16277,N_16013,N_16236);
nor U16278 (N_16278,N_16246,N_16041);
or U16279 (N_16279,N_16050,N_16174);
nor U16280 (N_16280,N_16164,N_16203);
nand U16281 (N_16281,N_16209,N_16034);
and U16282 (N_16282,N_16204,N_16227);
nand U16283 (N_16283,N_16000,N_16110);
nand U16284 (N_16284,N_16035,N_16122);
or U16285 (N_16285,N_16015,N_16177);
or U16286 (N_16286,N_16020,N_16066);
xnor U16287 (N_16287,N_16089,N_16052);
nor U16288 (N_16288,N_16085,N_16149);
nand U16289 (N_16289,N_16182,N_16081);
nor U16290 (N_16290,N_16082,N_16096);
xnor U16291 (N_16291,N_16150,N_16249);
and U16292 (N_16292,N_16008,N_16016);
or U16293 (N_16293,N_16130,N_16171);
and U16294 (N_16294,N_16097,N_16172);
or U16295 (N_16295,N_16205,N_16094);
or U16296 (N_16296,N_16135,N_16077);
xnor U16297 (N_16297,N_16118,N_16219);
and U16298 (N_16298,N_16119,N_16107);
nand U16299 (N_16299,N_16191,N_16142);
or U16300 (N_16300,N_16187,N_16222);
nor U16301 (N_16301,N_16176,N_16014);
nor U16302 (N_16302,N_16076,N_16103);
xnor U16303 (N_16303,N_16189,N_16004);
and U16304 (N_16304,N_16011,N_16038);
xnor U16305 (N_16305,N_16173,N_16148);
or U16306 (N_16306,N_16170,N_16136);
xor U16307 (N_16307,N_16238,N_16217);
nand U16308 (N_16308,N_16046,N_16057);
xor U16309 (N_16309,N_16044,N_16192);
and U16310 (N_16310,N_16145,N_16070);
nor U16311 (N_16311,N_16153,N_16231);
or U16312 (N_16312,N_16045,N_16053);
xnor U16313 (N_16313,N_16237,N_16124);
xnor U16314 (N_16314,N_16152,N_16063);
xnor U16315 (N_16315,N_16181,N_16218);
xor U16316 (N_16316,N_16006,N_16055);
nand U16317 (N_16317,N_16228,N_16244);
nor U16318 (N_16318,N_16141,N_16157);
xnor U16319 (N_16319,N_16245,N_16033);
nand U16320 (N_16320,N_16126,N_16175);
and U16321 (N_16321,N_16026,N_16121);
xor U16322 (N_16322,N_16084,N_16114);
or U16323 (N_16323,N_16019,N_16214);
nand U16324 (N_16324,N_16248,N_16199);
or U16325 (N_16325,N_16120,N_16159);
and U16326 (N_16326,N_16230,N_16113);
nand U16327 (N_16327,N_16106,N_16101);
and U16328 (N_16328,N_16198,N_16005);
nor U16329 (N_16329,N_16188,N_16169);
nor U16330 (N_16330,N_16102,N_16079);
or U16331 (N_16331,N_16090,N_16229);
nand U16332 (N_16332,N_16105,N_16029);
or U16333 (N_16333,N_16074,N_16239);
nor U16334 (N_16334,N_16206,N_16028);
xnor U16335 (N_16335,N_16195,N_16200);
or U16336 (N_16336,N_16213,N_16049);
and U16337 (N_16337,N_16134,N_16223);
or U16338 (N_16338,N_16221,N_16067);
nor U16339 (N_16339,N_16147,N_16099);
or U16340 (N_16340,N_16010,N_16163);
or U16341 (N_16341,N_16080,N_16158);
and U16342 (N_16342,N_16132,N_16128);
and U16343 (N_16343,N_16201,N_16232);
xnor U16344 (N_16344,N_16144,N_16220);
nor U16345 (N_16345,N_16138,N_16156);
or U16346 (N_16346,N_16061,N_16168);
nor U16347 (N_16347,N_16093,N_16139);
nand U16348 (N_16348,N_16018,N_16241);
nor U16349 (N_16349,N_16043,N_16068);
xnor U16350 (N_16350,N_16047,N_16032);
or U16351 (N_16351,N_16048,N_16112);
nor U16352 (N_16352,N_16143,N_16179);
or U16353 (N_16353,N_16180,N_16193);
or U16354 (N_16354,N_16017,N_16091);
or U16355 (N_16355,N_16036,N_16183);
nor U16356 (N_16356,N_16133,N_16069);
xnor U16357 (N_16357,N_16185,N_16086);
nand U16358 (N_16358,N_16233,N_16088);
nor U16359 (N_16359,N_16030,N_16039);
and U16360 (N_16360,N_16131,N_16025);
and U16361 (N_16361,N_16225,N_16196);
or U16362 (N_16362,N_16226,N_16207);
and U16363 (N_16363,N_16078,N_16197);
nand U16364 (N_16364,N_16060,N_16040);
nand U16365 (N_16365,N_16098,N_16243);
and U16366 (N_16366,N_16161,N_16100);
and U16367 (N_16367,N_16184,N_16024);
xor U16368 (N_16368,N_16234,N_16037);
nand U16369 (N_16369,N_16129,N_16065);
nor U16370 (N_16370,N_16127,N_16125);
nand U16371 (N_16371,N_16108,N_16162);
or U16372 (N_16372,N_16073,N_16194);
and U16373 (N_16373,N_16186,N_16208);
and U16374 (N_16374,N_16064,N_16211);
xnor U16375 (N_16375,N_16070,N_16199);
nor U16376 (N_16376,N_16191,N_16230);
nand U16377 (N_16377,N_16091,N_16095);
xnor U16378 (N_16378,N_16143,N_16226);
nand U16379 (N_16379,N_16145,N_16095);
or U16380 (N_16380,N_16024,N_16125);
or U16381 (N_16381,N_16096,N_16221);
xnor U16382 (N_16382,N_16234,N_16131);
or U16383 (N_16383,N_16235,N_16148);
and U16384 (N_16384,N_16198,N_16203);
xnor U16385 (N_16385,N_16230,N_16244);
nor U16386 (N_16386,N_16177,N_16191);
nor U16387 (N_16387,N_16073,N_16197);
nand U16388 (N_16388,N_16165,N_16222);
nor U16389 (N_16389,N_16234,N_16132);
and U16390 (N_16390,N_16083,N_16203);
nand U16391 (N_16391,N_16092,N_16000);
nor U16392 (N_16392,N_16143,N_16025);
nor U16393 (N_16393,N_16138,N_16012);
or U16394 (N_16394,N_16095,N_16008);
xor U16395 (N_16395,N_16016,N_16108);
nor U16396 (N_16396,N_16140,N_16099);
or U16397 (N_16397,N_16140,N_16065);
and U16398 (N_16398,N_16112,N_16070);
or U16399 (N_16399,N_16094,N_16017);
nand U16400 (N_16400,N_16188,N_16161);
nand U16401 (N_16401,N_16121,N_16144);
or U16402 (N_16402,N_16218,N_16187);
and U16403 (N_16403,N_16163,N_16225);
xnor U16404 (N_16404,N_16054,N_16149);
and U16405 (N_16405,N_16179,N_16198);
xnor U16406 (N_16406,N_16021,N_16145);
or U16407 (N_16407,N_16019,N_16075);
nand U16408 (N_16408,N_16021,N_16103);
and U16409 (N_16409,N_16221,N_16227);
and U16410 (N_16410,N_16226,N_16022);
nand U16411 (N_16411,N_16249,N_16034);
nand U16412 (N_16412,N_16230,N_16160);
xnor U16413 (N_16413,N_16037,N_16137);
xnor U16414 (N_16414,N_16043,N_16021);
and U16415 (N_16415,N_16196,N_16168);
nor U16416 (N_16416,N_16082,N_16150);
nand U16417 (N_16417,N_16048,N_16087);
xnor U16418 (N_16418,N_16152,N_16084);
xnor U16419 (N_16419,N_16170,N_16162);
and U16420 (N_16420,N_16237,N_16013);
and U16421 (N_16421,N_16044,N_16240);
nand U16422 (N_16422,N_16030,N_16172);
xnor U16423 (N_16423,N_16009,N_16185);
or U16424 (N_16424,N_16192,N_16026);
nor U16425 (N_16425,N_16007,N_16101);
nor U16426 (N_16426,N_16102,N_16241);
xnor U16427 (N_16427,N_16164,N_16199);
xnor U16428 (N_16428,N_16111,N_16018);
nand U16429 (N_16429,N_16030,N_16233);
nor U16430 (N_16430,N_16248,N_16200);
nand U16431 (N_16431,N_16046,N_16191);
or U16432 (N_16432,N_16013,N_16038);
and U16433 (N_16433,N_16215,N_16228);
and U16434 (N_16434,N_16198,N_16130);
xnor U16435 (N_16435,N_16147,N_16233);
nor U16436 (N_16436,N_16057,N_16135);
nand U16437 (N_16437,N_16114,N_16197);
xnor U16438 (N_16438,N_16050,N_16097);
xor U16439 (N_16439,N_16063,N_16164);
or U16440 (N_16440,N_16150,N_16032);
or U16441 (N_16441,N_16027,N_16205);
and U16442 (N_16442,N_16056,N_16169);
xor U16443 (N_16443,N_16233,N_16226);
nor U16444 (N_16444,N_16071,N_16095);
xor U16445 (N_16445,N_16002,N_16167);
nor U16446 (N_16446,N_16244,N_16238);
nor U16447 (N_16447,N_16194,N_16084);
or U16448 (N_16448,N_16125,N_16050);
nand U16449 (N_16449,N_16061,N_16120);
nor U16450 (N_16450,N_16143,N_16063);
xnor U16451 (N_16451,N_16002,N_16034);
or U16452 (N_16452,N_16193,N_16134);
nor U16453 (N_16453,N_16145,N_16156);
and U16454 (N_16454,N_16064,N_16068);
nor U16455 (N_16455,N_16041,N_16214);
nor U16456 (N_16456,N_16028,N_16047);
nand U16457 (N_16457,N_16018,N_16010);
nand U16458 (N_16458,N_16086,N_16115);
and U16459 (N_16459,N_16166,N_16022);
xor U16460 (N_16460,N_16050,N_16173);
and U16461 (N_16461,N_16099,N_16044);
or U16462 (N_16462,N_16240,N_16070);
nor U16463 (N_16463,N_16224,N_16211);
or U16464 (N_16464,N_16146,N_16182);
xor U16465 (N_16465,N_16159,N_16091);
nor U16466 (N_16466,N_16170,N_16002);
and U16467 (N_16467,N_16198,N_16206);
xor U16468 (N_16468,N_16055,N_16059);
nand U16469 (N_16469,N_16128,N_16125);
and U16470 (N_16470,N_16203,N_16147);
or U16471 (N_16471,N_16066,N_16160);
and U16472 (N_16472,N_16056,N_16058);
and U16473 (N_16473,N_16063,N_16121);
and U16474 (N_16474,N_16199,N_16167);
nand U16475 (N_16475,N_16226,N_16042);
nor U16476 (N_16476,N_16042,N_16214);
nand U16477 (N_16477,N_16126,N_16118);
nor U16478 (N_16478,N_16147,N_16232);
nor U16479 (N_16479,N_16099,N_16148);
or U16480 (N_16480,N_16044,N_16003);
or U16481 (N_16481,N_16113,N_16158);
or U16482 (N_16482,N_16221,N_16010);
nand U16483 (N_16483,N_16196,N_16220);
or U16484 (N_16484,N_16207,N_16004);
nand U16485 (N_16485,N_16059,N_16218);
nand U16486 (N_16486,N_16230,N_16216);
or U16487 (N_16487,N_16112,N_16040);
nor U16488 (N_16488,N_16106,N_16123);
or U16489 (N_16489,N_16112,N_16161);
and U16490 (N_16490,N_16147,N_16074);
and U16491 (N_16491,N_16177,N_16172);
and U16492 (N_16492,N_16098,N_16081);
or U16493 (N_16493,N_16166,N_16239);
or U16494 (N_16494,N_16116,N_16224);
xnor U16495 (N_16495,N_16120,N_16057);
xor U16496 (N_16496,N_16152,N_16087);
or U16497 (N_16497,N_16200,N_16015);
or U16498 (N_16498,N_16123,N_16067);
nand U16499 (N_16499,N_16190,N_16046);
or U16500 (N_16500,N_16425,N_16429);
xnor U16501 (N_16501,N_16318,N_16304);
xnor U16502 (N_16502,N_16255,N_16407);
nand U16503 (N_16503,N_16430,N_16380);
xnor U16504 (N_16504,N_16283,N_16329);
nand U16505 (N_16505,N_16491,N_16275);
xor U16506 (N_16506,N_16433,N_16485);
xnor U16507 (N_16507,N_16482,N_16466);
nor U16508 (N_16508,N_16293,N_16458);
nand U16509 (N_16509,N_16375,N_16441);
nor U16510 (N_16510,N_16442,N_16373);
nor U16511 (N_16511,N_16324,N_16473);
nand U16512 (N_16512,N_16376,N_16401);
and U16513 (N_16513,N_16261,N_16477);
or U16514 (N_16514,N_16278,N_16451);
nand U16515 (N_16515,N_16302,N_16287);
or U16516 (N_16516,N_16438,N_16445);
nor U16517 (N_16517,N_16332,N_16274);
and U16518 (N_16518,N_16454,N_16481);
xnor U16519 (N_16519,N_16369,N_16259);
nand U16520 (N_16520,N_16457,N_16410);
nand U16521 (N_16521,N_16415,N_16434);
nand U16522 (N_16522,N_16272,N_16495);
xor U16523 (N_16523,N_16319,N_16371);
nor U16524 (N_16524,N_16340,N_16417);
or U16525 (N_16525,N_16475,N_16269);
nand U16526 (N_16526,N_16471,N_16294);
nand U16527 (N_16527,N_16467,N_16443);
nor U16528 (N_16528,N_16455,N_16322);
xnor U16529 (N_16529,N_16363,N_16388);
or U16530 (N_16530,N_16306,N_16398);
nand U16531 (N_16531,N_16422,N_16374);
nand U16532 (N_16532,N_16483,N_16356);
nand U16533 (N_16533,N_16300,N_16346);
xor U16534 (N_16534,N_16428,N_16291);
nor U16535 (N_16535,N_16309,N_16265);
nor U16536 (N_16536,N_16449,N_16290);
and U16537 (N_16537,N_16366,N_16311);
and U16538 (N_16538,N_16260,N_16253);
xnor U16539 (N_16539,N_16280,N_16459);
xor U16540 (N_16540,N_16431,N_16386);
and U16541 (N_16541,N_16297,N_16270);
nand U16542 (N_16542,N_16258,N_16406);
and U16543 (N_16543,N_16305,N_16333);
nand U16544 (N_16544,N_16416,N_16472);
and U16545 (N_16545,N_16492,N_16321);
and U16546 (N_16546,N_16404,N_16279);
nor U16547 (N_16547,N_16350,N_16489);
nor U16548 (N_16548,N_16385,N_16353);
nor U16549 (N_16549,N_16354,N_16381);
nor U16550 (N_16550,N_16468,N_16336);
and U16551 (N_16551,N_16408,N_16362);
or U16552 (N_16552,N_16469,N_16310);
nand U16553 (N_16553,N_16264,N_16383);
nand U16554 (N_16554,N_16476,N_16341);
nor U16555 (N_16555,N_16478,N_16316);
nand U16556 (N_16556,N_16320,N_16301);
nand U16557 (N_16557,N_16420,N_16326);
nor U16558 (N_16558,N_16395,N_16393);
or U16559 (N_16559,N_16414,N_16251);
nand U16560 (N_16560,N_16338,N_16282);
or U16561 (N_16561,N_16327,N_16440);
and U16562 (N_16562,N_16285,N_16387);
nand U16563 (N_16563,N_16389,N_16367);
xnor U16564 (N_16564,N_16368,N_16288);
or U16565 (N_16565,N_16384,N_16418);
nor U16566 (N_16566,N_16273,N_16358);
nand U16567 (N_16567,N_16360,N_16463);
or U16568 (N_16568,N_16343,N_16337);
and U16569 (N_16569,N_16487,N_16413);
nor U16570 (N_16570,N_16335,N_16446);
xnor U16571 (N_16571,N_16490,N_16361);
and U16572 (N_16572,N_16252,N_16392);
xor U16573 (N_16573,N_16464,N_16372);
nor U16574 (N_16574,N_16267,N_16352);
xor U16575 (N_16575,N_16325,N_16462);
xnor U16576 (N_16576,N_16289,N_16480);
or U16577 (N_16577,N_16379,N_16439);
and U16578 (N_16578,N_16357,N_16263);
or U16579 (N_16579,N_16403,N_16437);
nand U16580 (N_16580,N_16447,N_16461);
nand U16581 (N_16581,N_16390,N_16497);
or U16582 (N_16582,N_16470,N_16342);
nand U16583 (N_16583,N_16323,N_16498);
nor U16584 (N_16584,N_16378,N_16496);
and U16585 (N_16585,N_16339,N_16370);
nand U16586 (N_16586,N_16331,N_16421);
nor U16587 (N_16587,N_16411,N_16276);
nand U16588 (N_16588,N_16365,N_16493);
and U16589 (N_16589,N_16298,N_16399);
and U16590 (N_16590,N_16423,N_16412);
and U16591 (N_16591,N_16486,N_16292);
nand U16592 (N_16592,N_16499,N_16479);
or U16593 (N_16593,N_16400,N_16317);
nor U16594 (N_16594,N_16277,N_16452);
and U16595 (N_16595,N_16494,N_16303);
nand U16596 (N_16596,N_16344,N_16271);
nor U16597 (N_16597,N_16436,N_16250);
nor U16598 (N_16598,N_16453,N_16460);
xnor U16599 (N_16599,N_16296,N_16450);
nor U16600 (N_16600,N_16488,N_16426);
nand U16601 (N_16601,N_16262,N_16444);
nor U16602 (N_16602,N_16397,N_16474);
xnor U16603 (N_16603,N_16382,N_16284);
and U16604 (N_16604,N_16359,N_16465);
nor U16605 (N_16605,N_16394,N_16409);
nor U16606 (N_16606,N_16351,N_16377);
or U16607 (N_16607,N_16312,N_16402);
nand U16608 (N_16608,N_16345,N_16348);
nor U16609 (N_16609,N_16257,N_16405);
nand U16610 (N_16610,N_16435,N_16313);
xor U16611 (N_16611,N_16396,N_16484);
or U16612 (N_16612,N_16330,N_16281);
or U16613 (N_16613,N_16456,N_16334);
nand U16614 (N_16614,N_16448,N_16256);
and U16615 (N_16615,N_16391,N_16266);
nor U16616 (N_16616,N_16286,N_16349);
or U16617 (N_16617,N_16268,N_16424);
or U16618 (N_16618,N_16307,N_16328);
or U16619 (N_16619,N_16364,N_16315);
or U16620 (N_16620,N_16419,N_16427);
xnor U16621 (N_16621,N_16432,N_16254);
and U16622 (N_16622,N_16299,N_16314);
nor U16623 (N_16623,N_16347,N_16295);
xor U16624 (N_16624,N_16308,N_16355);
nor U16625 (N_16625,N_16338,N_16304);
xor U16626 (N_16626,N_16253,N_16306);
nor U16627 (N_16627,N_16255,N_16475);
nand U16628 (N_16628,N_16371,N_16309);
nand U16629 (N_16629,N_16488,N_16330);
or U16630 (N_16630,N_16271,N_16270);
or U16631 (N_16631,N_16406,N_16342);
or U16632 (N_16632,N_16366,N_16287);
and U16633 (N_16633,N_16444,N_16378);
nand U16634 (N_16634,N_16327,N_16346);
xnor U16635 (N_16635,N_16308,N_16432);
nand U16636 (N_16636,N_16291,N_16453);
xor U16637 (N_16637,N_16296,N_16302);
xnor U16638 (N_16638,N_16490,N_16335);
nor U16639 (N_16639,N_16340,N_16402);
xnor U16640 (N_16640,N_16320,N_16327);
nor U16641 (N_16641,N_16400,N_16498);
xnor U16642 (N_16642,N_16362,N_16448);
xor U16643 (N_16643,N_16456,N_16383);
nand U16644 (N_16644,N_16259,N_16363);
xnor U16645 (N_16645,N_16285,N_16362);
nor U16646 (N_16646,N_16317,N_16413);
nor U16647 (N_16647,N_16308,N_16371);
nor U16648 (N_16648,N_16375,N_16488);
and U16649 (N_16649,N_16490,N_16432);
and U16650 (N_16650,N_16495,N_16317);
or U16651 (N_16651,N_16359,N_16438);
or U16652 (N_16652,N_16405,N_16401);
xor U16653 (N_16653,N_16270,N_16455);
or U16654 (N_16654,N_16486,N_16443);
or U16655 (N_16655,N_16364,N_16283);
nor U16656 (N_16656,N_16270,N_16415);
nand U16657 (N_16657,N_16284,N_16376);
nor U16658 (N_16658,N_16278,N_16392);
nor U16659 (N_16659,N_16428,N_16295);
and U16660 (N_16660,N_16382,N_16292);
nand U16661 (N_16661,N_16340,N_16392);
xor U16662 (N_16662,N_16295,N_16294);
and U16663 (N_16663,N_16470,N_16354);
and U16664 (N_16664,N_16364,N_16488);
or U16665 (N_16665,N_16315,N_16374);
and U16666 (N_16666,N_16425,N_16370);
or U16667 (N_16667,N_16331,N_16250);
nor U16668 (N_16668,N_16269,N_16283);
or U16669 (N_16669,N_16422,N_16360);
or U16670 (N_16670,N_16374,N_16303);
nand U16671 (N_16671,N_16261,N_16468);
nand U16672 (N_16672,N_16484,N_16410);
or U16673 (N_16673,N_16345,N_16496);
nor U16674 (N_16674,N_16342,N_16438);
and U16675 (N_16675,N_16268,N_16350);
nor U16676 (N_16676,N_16351,N_16311);
and U16677 (N_16677,N_16465,N_16384);
or U16678 (N_16678,N_16489,N_16337);
or U16679 (N_16679,N_16416,N_16494);
nand U16680 (N_16680,N_16315,N_16253);
nand U16681 (N_16681,N_16303,N_16344);
or U16682 (N_16682,N_16399,N_16492);
xor U16683 (N_16683,N_16386,N_16383);
nor U16684 (N_16684,N_16411,N_16350);
or U16685 (N_16685,N_16298,N_16404);
and U16686 (N_16686,N_16444,N_16359);
and U16687 (N_16687,N_16404,N_16320);
and U16688 (N_16688,N_16387,N_16388);
nor U16689 (N_16689,N_16398,N_16402);
nor U16690 (N_16690,N_16260,N_16444);
xor U16691 (N_16691,N_16424,N_16325);
and U16692 (N_16692,N_16457,N_16346);
nand U16693 (N_16693,N_16446,N_16392);
nor U16694 (N_16694,N_16279,N_16259);
xor U16695 (N_16695,N_16455,N_16382);
or U16696 (N_16696,N_16370,N_16266);
and U16697 (N_16697,N_16267,N_16343);
nor U16698 (N_16698,N_16400,N_16289);
xnor U16699 (N_16699,N_16312,N_16356);
or U16700 (N_16700,N_16475,N_16471);
xnor U16701 (N_16701,N_16475,N_16478);
or U16702 (N_16702,N_16388,N_16277);
xor U16703 (N_16703,N_16438,N_16326);
xor U16704 (N_16704,N_16272,N_16423);
xnor U16705 (N_16705,N_16406,N_16418);
nor U16706 (N_16706,N_16476,N_16273);
and U16707 (N_16707,N_16467,N_16271);
xor U16708 (N_16708,N_16334,N_16476);
xnor U16709 (N_16709,N_16463,N_16398);
nand U16710 (N_16710,N_16464,N_16477);
and U16711 (N_16711,N_16437,N_16289);
or U16712 (N_16712,N_16314,N_16307);
nand U16713 (N_16713,N_16306,N_16495);
and U16714 (N_16714,N_16372,N_16478);
xor U16715 (N_16715,N_16395,N_16487);
and U16716 (N_16716,N_16318,N_16448);
xnor U16717 (N_16717,N_16429,N_16366);
or U16718 (N_16718,N_16472,N_16279);
nand U16719 (N_16719,N_16440,N_16410);
nand U16720 (N_16720,N_16382,N_16463);
or U16721 (N_16721,N_16419,N_16461);
nand U16722 (N_16722,N_16286,N_16301);
and U16723 (N_16723,N_16314,N_16442);
or U16724 (N_16724,N_16270,N_16333);
nor U16725 (N_16725,N_16498,N_16304);
nand U16726 (N_16726,N_16331,N_16314);
nor U16727 (N_16727,N_16323,N_16404);
and U16728 (N_16728,N_16300,N_16451);
or U16729 (N_16729,N_16259,N_16447);
nor U16730 (N_16730,N_16290,N_16482);
and U16731 (N_16731,N_16422,N_16341);
nor U16732 (N_16732,N_16366,N_16480);
nor U16733 (N_16733,N_16366,N_16493);
xnor U16734 (N_16734,N_16395,N_16403);
or U16735 (N_16735,N_16353,N_16403);
nor U16736 (N_16736,N_16279,N_16296);
or U16737 (N_16737,N_16342,N_16471);
nor U16738 (N_16738,N_16342,N_16417);
nand U16739 (N_16739,N_16426,N_16462);
nor U16740 (N_16740,N_16361,N_16416);
or U16741 (N_16741,N_16470,N_16461);
nand U16742 (N_16742,N_16405,N_16354);
nand U16743 (N_16743,N_16370,N_16352);
or U16744 (N_16744,N_16274,N_16489);
nor U16745 (N_16745,N_16377,N_16295);
or U16746 (N_16746,N_16321,N_16434);
and U16747 (N_16747,N_16408,N_16315);
xnor U16748 (N_16748,N_16412,N_16440);
nor U16749 (N_16749,N_16313,N_16410);
and U16750 (N_16750,N_16611,N_16501);
nand U16751 (N_16751,N_16609,N_16726);
and U16752 (N_16752,N_16602,N_16530);
or U16753 (N_16753,N_16705,N_16581);
nand U16754 (N_16754,N_16606,N_16585);
and U16755 (N_16755,N_16560,N_16500);
xnor U16756 (N_16756,N_16564,N_16590);
and U16757 (N_16757,N_16553,N_16698);
xor U16758 (N_16758,N_16637,N_16510);
nor U16759 (N_16759,N_16523,N_16638);
nand U16760 (N_16760,N_16742,N_16628);
nand U16761 (N_16761,N_16616,N_16556);
nor U16762 (N_16762,N_16506,N_16620);
nand U16763 (N_16763,N_16540,N_16548);
nor U16764 (N_16764,N_16708,N_16626);
nor U16765 (N_16765,N_16593,N_16549);
xnor U16766 (N_16766,N_16656,N_16588);
nand U16767 (N_16767,N_16517,N_16610);
nand U16768 (N_16768,N_16583,N_16561);
nand U16769 (N_16769,N_16614,N_16687);
xor U16770 (N_16770,N_16557,N_16694);
xor U16771 (N_16771,N_16675,N_16571);
nand U16772 (N_16772,N_16728,N_16711);
nor U16773 (N_16773,N_16743,N_16684);
or U16774 (N_16774,N_16587,N_16736);
or U16775 (N_16775,N_16550,N_16543);
nor U16776 (N_16776,N_16563,N_16525);
and U16777 (N_16777,N_16535,N_16701);
nor U16778 (N_16778,N_16720,N_16686);
nand U16779 (N_16779,N_16747,N_16661);
xnor U16780 (N_16780,N_16714,N_16624);
or U16781 (N_16781,N_16601,N_16539);
or U16782 (N_16782,N_16635,N_16679);
nand U16783 (N_16783,N_16666,N_16580);
nor U16784 (N_16784,N_16740,N_16589);
nor U16785 (N_16785,N_16645,N_16572);
nand U16786 (N_16786,N_16668,N_16534);
and U16787 (N_16787,N_16651,N_16691);
nand U16788 (N_16788,N_16622,N_16677);
or U16789 (N_16789,N_16575,N_16715);
and U16790 (N_16790,N_16554,N_16703);
nor U16791 (N_16791,N_16612,N_16591);
or U16792 (N_16792,N_16745,N_16707);
nor U16793 (N_16793,N_16737,N_16644);
nor U16794 (N_16794,N_16657,N_16710);
nor U16795 (N_16795,N_16502,N_16746);
nand U16796 (N_16796,N_16536,N_16749);
nand U16797 (N_16797,N_16521,N_16515);
or U16798 (N_16798,N_16735,N_16692);
xor U16799 (N_16799,N_16717,N_16505);
and U16800 (N_16800,N_16531,N_16649);
xor U16801 (N_16801,N_16532,N_16689);
xnor U16802 (N_16802,N_16570,N_16600);
and U16803 (N_16803,N_16704,N_16568);
nor U16804 (N_16804,N_16509,N_16518);
and U16805 (N_16805,N_16594,N_16648);
xnor U16806 (N_16806,N_16706,N_16725);
xnor U16807 (N_16807,N_16538,N_16596);
and U16808 (N_16808,N_16663,N_16507);
nor U16809 (N_16809,N_16730,N_16617);
nand U16810 (N_16810,N_16662,N_16603);
and U16811 (N_16811,N_16697,N_16630);
and U16812 (N_16812,N_16695,N_16627);
and U16813 (N_16813,N_16597,N_16709);
xnor U16814 (N_16814,N_16653,N_16723);
xor U16815 (N_16815,N_16607,N_16551);
xnor U16816 (N_16816,N_16744,N_16696);
nor U16817 (N_16817,N_16524,N_16579);
nand U16818 (N_16818,N_16618,N_16567);
xor U16819 (N_16819,N_16672,N_16647);
nor U16820 (N_16820,N_16546,N_16660);
nor U16821 (N_16821,N_16576,N_16727);
nand U16822 (N_16822,N_16503,N_16673);
xnor U16823 (N_16823,N_16682,N_16573);
or U16824 (N_16824,N_16513,N_16693);
nor U16825 (N_16825,N_16658,N_16674);
and U16826 (N_16826,N_16562,N_16639);
nand U16827 (N_16827,N_16729,N_16699);
nor U16828 (N_16828,N_16731,N_16512);
and U16829 (N_16829,N_16718,N_16641);
nor U16830 (N_16830,N_16566,N_16688);
nand U16831 (N_16831,N_16748,N_16592);
and U16832 (N_16832,N_16640,N_16632);
nand U16833 (N_16833,N_16719,N_16508);
nor U16834 (N_16834,N_16741,N_16529);
xor U16835 (N_16835,N_16613,N_16646);
nor U16836 (N_16836,N_16631,N_16516);
or U16837 (N_16837,N_16724,N_16669);
nand U16838 (N_16838,N_16514,N_16511);
and U16839 (N_16839,N_16685,N_16713);
and U16840 (N_16840,N_16528,N_16667);
nand U16841 (N_16841,N_16636,N_16683);
nor U16842 (N_16842,N_16526,N_16544);
xnor U16843 (N_16843,N_16598,N_16738);
or U16844 (N_16844,N_16665,N_16599);
xor U16845 (N_16845,N_16520,N_16605);
nand U16846 (N_16846,N_16615,N_16739);
nor U16847 (N_16847,N_16732,N_16574);
nand U16848 (N_16848,N_16504,N_16608);
xnor U16849 (N_16849,N_16569,N_16537);
xnor U16850 (N_16850,N_16712,N_16533);
or U16851 (N_16851,N_16678,N_16633);
or U16852 (N_16852,N_16643,N_16676);
and U16853 (N_16853,N_16582,N_16604);
nor U16854 (N_16854,N_16652,N_16664);
nand U16855 (N_16855,N_16733,N_16519);
or U16856 (N_16856,N_16595,N_16642);
xnor U16857 (N_16857,N_16629,N_16680);
nor U16858 (N_16858,N_16552,N_16654);
and U16859 (N_16859,N_16681,N_16545);
xnor U16860 (N_16860,N_16734,N_16650);
and U16861 (N_16861,N_16702,N_16659);
nand U16862 (N_16862,N_16578,N_16621);
xor U16863 (N_16863,N_16655,N_16690);
xor U16864 (N_16864,N_16559,N_16542);
or U16865 (N_16865,N_16558,N_16619);
and U16866 (N_16866,N_16722,N_16577);
xnor U16867 (N_16867,N_16623,N_16634);
nand U16868 (N_16868,N_16625,N_16671);
and U16869 (N_16869,N_16716,N_16527);
or U16870 (N_16870,N_16670,N_16547);
and U16871 (N_16871,N_16586,N_16522);
xor U16872 (N_16872,N_16700,N_16555);
xor U16873 (N_16873,N_16565,N_16721);
xor U16874 (N_16874,N_16584,N_16541);
xnor U16875 (N_16875,N_16602,N_16624);
nand U16876 (N_16876,N_16517,N_16638);
or U16877 (N_16877,N_16690,N_16534);
and U16878 (N_16878,N_16529,N_16574);
and U16879 (N_16879,N_16599,N_16598);
xor U16880 (N_16880,N_16688,N_16518);
nor U16881 (N_16881,N_16614,N_16685);
nor U16882 (N_16882,N_16576,N_16597);
or U16883 (N_16883,N_16749,N_16671);
or U16884 (N_16884,N_16614,N_16632);
and U16885 (N_16885,N_16634,N_16744);
nor U16886 (N_16886,N_16553,N_16747);
or U16887 (N_16887,N_16587,N_16679);
and U16888 (N_16888,N_16587,N_16543);
xor U16889 (N_16889,N_16632,N_16626);
xor U16890 (N_16890,N_16722,N_16639);
and U16891 (N_16891,N_16672,N_16634);
nor U16892 (N_16892,N_16516,N_16517);
or U16893 (N_16893,N_16695,N_16616);
nand U16894 (N_16894,N_16744,N_16610);
and U16895 (N_16895,N_16620,N_16543);
xnor U16896 (N_16896,N_16560,N_16521);
nor U16897 (N_16897,N_16518,N_16696);
or U16898 (N_16898,N_16502,N_16529);
xor U16899 (N_16899,N_16624,N_16645);
nand U16900 (N_16900,N_16607,N_16721);
nor U16901 (N_16901,N_16715,N_16735);
nand U16902 (N_16902,N_16507,N_16571);
nor U16903 (N_16903,N_16689,N_16692);
and U16904 (N_16904,N_16739,N_16643);
or U16905 (N_16905,N_16614,N_16651);
or U16906 (N_16906,N_16671,N_16663);
xor U16907 (N_16907,N_16737,N_16588);
xor U16908 (N_16908,N_16550,N_16625);
nor U16909 (N_16909,N_16633,N_16560);
and U16910 (N_16910,N_16739,N_16725);
xor U16911 (N_16911,N_16690,N_16537);
or U16912 (N_16912,N_16656,N_16506);
or U16913 (N_16913,N_16734,N_16690);
xor U16914 (N_16914,N_16594,N_16700);
nand U16915 (N_16915,N_16707,N_16599);
nand U16916 (N_16916,N_16557,N_16561);
or U16917 (N_16917,N_16647,N_16668);
or U16918 (N_16918,N_16511,N_16717);
or U16919 (N_16919,N_16607,N_16715);
xor U16920 (N_16920,N_16536,N_16504);
or U16921 (N_16921,N_16654,N_16663);
nor U16922 (N_16922,N_16694,N_16525);
and U16923 (N_16923,N_16579,N_16608);
and U16924 (N_16924,N_16507,N_16570);
or U16925 (N_16925,N_16552,N_16572);
xor U16926 (N_16926,N_16615,N_16566);
xor U16927 (N_16927,N_16640,N_16696);
nand U16928 (N_16928,N_16541,N_16743);
or U16929 (N_16929,N_16564,N_16650);
and U16930 (N_16930,N_16729,N_16710);
nand U16931 (N_16931,N_16528,N_16715);
and U16932 (N_16932,N_16611,N_16552);
nor U16933 (N_16933,N_16519,N_16535);
xnor U16934 (N_16934,N_16653,N_16691);
nor U16935 (N_16935,N_16584,N_16598);
nor U16936 (N_16936,N_16642,N_16599);
or U16937 (N_16937,N_16664,N_16639);
xor U16938 (N_16938,N_16554,N_16714);
or U16939 (N_16939,N_16505,N_16573);
or U16940 (N_16940,N_16509,N_16702);
nor U16941 (N_16941,N_16704,N_16712);
nand U16942 (N_16942,N_16582,N_16668);
or U16943 (N_16943,N_16608,N_16549);
nor U16944 (N_16944,N_16551,N_16710);
and U16945 (N_16945,N_16634,N_16559);
and U16946 (N_16946,N_16663,N_16574);
nand U16947 (N_16947,N_16674,N_16749);
and U16948 (N_16948,N_16627,N_16619);
nand U16949 (N_16949,N_16634,N_16628);
xor U16950 (N_16950,N_16672,N_16567);
nor U16951 (N_16951,N_16595,N_16589);
and U16952 (N_16952,N_16622,N_16684);
xnor U16953 (N_16953,N_16641,N_16663);
nand U16954 (N_16954,N_16625,N_16529);
nor U16955 (N_16955,N_16573,N_16531);
or U16956 (N_16956,N_16681,N_16649);
or U16957 (N_16957,N_16527,N_16627);
nor U16958 (N_16958,N_16721,N_16653);
nand U16959 (N_16959,N_16609,N_16548);
xor U16960 (N_16960,N_16673,N_16708);
nor U16961 (N_16961,N_16539,N_16500);
nor U16962 (N_16962,N_16695,N_16665);
or U16963 (N_16963,N_16584,N_16664);
xor U16964 (N_16964,N_16736,N_16703);
xor U16965 (N_16965,N_16749,N_16622);
and U16966 (N_16966,N_16521,N_16730);
and U16967 (N_16967,N_16610,N_16672);
nand U16968 (N_16968,N_16700,N_16622);
and U16969 (N_16969,N_16645,N_16573);
nor U16970 (N_16970,N_16627,N_16722);
and U16971 (N_16971,N_16628,N_16538);
and U16972 (N_16972,N_16748,N_16700);
xnor U16973 (N_16973,N_16665,N_16540);
xnor U16974 (N_16974,N_16643,N_16503);
nor U16975 (N_16975,N_16699,N_16530);
nor U16976 (N_16976,N_16708,N_16615);
and U16977 (N_16977,N_16606,N_16611);
or U16978 (N_16978,N_16622,N_16698);
xor U16979 (N_16979,N_16583,N_16552);
nand U16980 (N_16980,N_16544,N_16716);
nor U16981 (N_16981,N_16553,N_16543);
xnor U16982 (N_16982,N_16628,N_16696);
xor U16983 (N_16983,N_16624,N_16666);
xor U16984 (N_16984,N_16748,N_16686);
and U16985 (N_16985,N_16563,N_16724);
xnor U16986 (N_16986,N_16591,N_16627);
and U16987 (N_16987,N_16655,N_16596);
xor U16988 (N_16988,N_16594,N_16730);
xnor U16989 (N_16989,N_16690,N_16583);
nand U16990 (N_16990,N_16669,N_16665);
nand U16991 (N_16991,N_16707,N_16653);
or U16992 (N_16992,N_16710,N_16559);
or U16993 (N_16993,N_16705,N_16613);
and U16994 (N_16994,N_16626,N_16559);
and U16995 (N_16995,N_16705,N_16646);
or U16996 (N_16996,N_16574,N_16677);
xor U16997 (N_16997,N_16637,N_16590);
nor U16998 (N_16998,N_16544,N_16612);
nor U16999 (N_16999,N_16629,N_16613);
and U17000 (N_17000,N_16824,N_16972);
or U17001 (N_17001,N_16942,N_16919);
or U17002 (N_17002,N_16799,N_16950);
xnor U17003 (N_17003,N_16957,N_16829);
and U17004 (N_17004,N_16768,N_16977);
or U17005 (N_17005,N_16995,N_16764);
and U17006 (N_17006,N_16795,N_16853);
nor U17007 (N_17007,N_16828,N_16976);
xnor U17008 (N_17008,N_16939,N_16763);
nor U17009 (N_17009,N_16931,N_16888);
and U17010 (N_17010,N_16982,N_16994);
xnor U17011 (N_17011,N_16883,N_16997);
xor U17012 (N_17012,N_16865,N_16958);
xor U17013 (N_17013,N_16776,N_16999);
xnor U17014 (N_17014,N_16819,N_16875);
or U17015 (N_17015,N_16936,N_16849);
xor U17016 (N_17016,N_16884,N_16761);
xor U17017 (N_17017,N_16793,N_16953);
or U17018 (N_17018,N_16855,N_16991);
nor U17019 (N_17019,N_16765,N_16815);
or U17020 (N_17020,N_16965,N_16927);
or U17021 (N_17021,N_16978,N_16962);
xor U17022 (N_17022,N_16791,N_16868);
and U17023 (N_17023,N_16970,N_16785);
or U17024 (N_17024,N_16794,N_16760);
xor U17025 (N_17025,N_16968,N_16906);
xor U17026 (N_17026,N_16837,N_16803);
xor U17027 (N_17027,N_16992,N_16832);
or U17028 (N_17028,N_16983,N_16891);
or U17029 (N_17029,N_16933,N_16897);
nor U17030 (N_17030,N_16893,N_16870);
or U17031 (N_17031,N_16759,N_16781);
or U17032 (N_17032,N_16964,N_16812);
and U17033 (N_17033,N_16998,N_16881);
and U17034 (N_17034,N_16887,N_16873);
nor U17035 (N_17035,N_16802,N_16782);
nor U17036 (N_17036,N_16834,N_16894);
nor U17037 (N_17037,N_16949,N_16818);
or U17038 (N_17038,N_16825,N_16928);
and U17039 (N_17039,N_16833,N_16923);
xor U17040 (N_17040,N_16902,N_16912);
nand U17041 (N_17041,N_16984,N_16753);
and U17042 (N_17042,N_16806,N_16915);
nand U17043 (N_17043,N_16948,N_16770);
nand U17044 (N_17044,N_16911,N_16941);
nor U17045 (N_17045,N_16905,N_16916);
nand U17046 (N_17046,N_16775,N_16839);
nor U17047 (N_17047,N_16798,N_16898);
or U17048 (N_17048,N_16867,N_16751);
or U17049 (N_17049,N_16845,N_16773);
nor U17050 (N_17050,N_16967,N_16856);
and U17051 (N_17051,N_16988,N_16841);
or U17052 (N_17052,N_16935,N_16771);
and U17053 (N_17053,N_16981,N_16779);
or U17054 (N_17054,N_16811,N_16940);
nand U17055 (N_17055,N_16838,N_16857);
nor U17056 (N_17056,N_16872,N_16844);
or U17057 (N_17057,N_16947,N_16861);
or U17058 (N_17058,N_16980,N_16787);
and U17059 (N_17059,N_16914,N_16859);
or U17060 (N_17060,N_16769,N_16896);
nor U17061 (N_17061,N_16821,N_16890);
nor U17062 (N_17062,N_16974,N_16926);
xor U17063 (N_17063,N_16805,N_16880);
nand U17064 (N_17064,N_16847,N_16752);
and U17065 (N_17065,N_16943,N_16971);
nand U17066 (N_17066,N_16777,N_16944);
or U17067 (N_17067,N_16985,N_16850);
nor U17068 (N_17068,N_16796,N_16929);
nor U17069 (N_17069,N_16809,N_16904);
nand U17070 (N_17070,N_16879,N_16774);
nor U17071 (N_17071,N_16808,N_16804);
and U17072 (N_17072,N_16784,N_16973);
nor U17073 (N_17073,N_16755,N_16917);
nand U17074 (N_17074,N_16956,N_16959);
or U17075 (N_17075,N_16756,N_16786);
or U17076 (N_17076,N_16816,N_16899);
or U17077 (N_17077,N_16934,N_16930);
or U17078 (N_17078,N_16869,N_16862);
or U17079 (N_17079,N_16979,N_16963);
xnor U17080 (N_17080,N_16848,N_16827);
nor U17081 (N_17081,N_16987,N_16820);
nor U17082 (N_17082,N_16750,N_16840);
nor U17083 (N_17083,N_16907,N_16797);
or U17084 (N_17084,N_16858,N_16780);
nand U17085 (N_17085,N_16801,N_16903);
and U17086 (N_17086,N_16792,N_16854);
nand U17087 (N_17087,N_16975,N_16932);
xor U17088 (N_17088,N_16989,N_16789);
or U17089 (N_17089,N_16996,N_16910);
nand U17090 (N_17090,N_16826,N_16835);
nor U17091 (N_17091,N_16900,N_16871);
or U17092 (N_17092,N_16754,N_16758);
nor U17093 (N_17093,N_16955,N_16922);
nand U17094 (N_17094,N_16924,N_16966);
or U17095 (N_17095,N_16954,N_16843);
or U17096 (N_17096,N_16790,N_16895);
nand U17097 (N_17097,N_16757,N_16990);
or U17098 (N_17098,N_16772,N_16866);
xor U17099 (N_17099,N_16766,N_16778);
nand U17100 (N_17100,N_16961,N_16960);
or U17101 (N_17101,N_16908,N_16945);
xnor U17102 (N_17102,N_16851,N_16813);
and U17103 (N_17103,N_16882,N_16800);
and U17104 (N_17104,N_16864,N_16993);
xor U17105 (N_17105,N_16852,N_16886);
nand U17106 (N_17106,N_16822,N_16909);
nand U17107 (N_17107,N_16901,N_16952);
xor U17108 (N_17108,N_16986,N_16913);
and U17109 (N_17109,N_16885,N_16876);
or U17110 (N_17110,N_16937,N_16920);
xnor U17111 (N_17111,N_16877,N_16874);
or U17112 (N_17112,N_16938,N_16842);
or U17113 (N_17113,N_16892,N_16921);
nand U17114 (N_17114,N_16846,N_16863);
nor U17115 (N_17115,N_16946,N_16951);
nand U17116 (N_17116,N_16889,N_16830);
nor U17117 (N_17117,N_16807,N_16925);
nand U17118 (N_17118,N_16783,N_16831);
or U17119 (N_17119,N_16969,N_16788);
nor U17120 (N_17120,N_16814,N_16918);
nand U17121 (N_17121,N_16767,N_16817);
or U17122 (N_17122,N_16860,N_16836);
or U17123 (N_17123,N_16762,N_16810);
or U17124 (N_17124,N_16823,N_16878);
xor U17125 (N_17125,N_16825,N_16860);
and U17126 (N_17126,N_16892,N_16887);
or U17127 (N_17127,N_16937,N_16950);
and U17128 (N_17128,N_16831,N_16884);
xor U17129 (N_17129,N_16767,N_16953);
nor U17130 (N_17130,N_16959,N_16914);
nor U17131 (N_17131,N_16961,N_16803);
nand U17132 (N_17132,N_16891,N_16885);
or U17133 (N_17133,N_16846,N_16956);
nor U17134 (N_17134,N_16841,N_16766);
nand U17135 (N_17135,N_16839,N_16762);
nand U17136 (N_17136,N_16806,N_16896);
and U17137 (N_17137,N_16822,N_16923);
nor U17138 (N_17138,N_16952,N_16883);
xor U17139 (N_17139,N_16927,N_16941);
xor U17140 (N_17140,N_16971,N_16857);
nand U17141 (N_17141,N_16908,N_16833);
xnor U17142 (N_17142,N_16842,N_16862);
nor U17143 (N_17143,N_16781,N_16863);
nand U17144 (N_17144,N_16921,N_16880);
xnor U17145 (N_17145,N_16923,N_16924);
nand U17146 (N_17146,N_16775,N_16805);
xor U17147 (N_17147,N_16953,N_16969);
and U17148 (N_17148,N_16786,N_16750);
nor U17149 (N_17149,N_16807,N_16760);
nand U17150 (N_17150,N_16968,N_16987);
nand U17151 (N_17151,N_16892,N_16881);
or U17152 (N_17152,N_16996,N_16758);
xor U17153 (N_17153,N_16817,N_16963);
and U17154 (N_17154,N_16943,N_16999);
nor U17155 (N_17155,N_16785,N_16777);
nor U17156 (N_17156,N_16971,N_16768);
nand U17157 (N_17157,N_16815,N_16792);
nand U17158 (N_17158,N_16854,N_16911);
or U17159 (N_17159,N_16949,N_16973);
xnor U17160 (N_17160,N_16963,N_16961);
nand U17161 (N_17161,N_16959,N_16750);
or U17162 (N_17162,N_16837,N_16986);
xnor U17163 (N_17163,N_16959,N_16934);
and U17164 (N_17164,N_16957,N_16941);
nor U17165 (N_17165,N_16941,N_16960);
nand U17166 (N_17166,N_16826,N_16804);
or U17167 (N_17167,N_16886,N_16978);
xnor U17168 (N_17168,N_16784,N_16915);
and U17169 (N_17169,N_16933,N_16779);
nand U17170 (N_17170,N_16947,N_16996);
or U17171 (N_17171,N_16865,N_16918);
or U17172 (N_17172,N_16930,N_16771);
nor U17173 (N_17173,N_16889,N_16754);
nand U17174 (N_17174,N_16891,N_16862);
nor U17175 (N_17175,N_16981,N_16965);
nand U17176 (N_17176,N_16787,N_16972);
and U17177 (N_17177,N_16920,N_16951);
or U17178 (N_17178,N_16785,N_16854);
xor U17179 (N_17179,N_16912,N_16819);
nor U17180 (N_17180,N_16830,N_16751);
and U17181 (N_17181,N_16830,N_16809);
or U17182 (N_17182,N_16932,N_16757);
nand U17183 (N_17183,N_16933,N_16758);
nor U17184 (N_17184,N_16881,N_16852);
xnor U17185 (N_17185,N_16953,N_16802);
xnor U17186 (N_17186,N_16830,N_16769);
or U17187 (N_17187,N_16830,N_16789);
nor U17188 (N_17188,N_16866,N_16894);
nand U17189 (N_17189,N_16900,N_16947);
nor U17190 (N_17190,N_16985,N_16845);
or U17191 (N_17191,N_16848,N_16821);
nor U17192 (N_17192,N_16929,N_16987);
nand U17193 (N_17193,N_16990,N_16987);
xor U17194 (N_17194,N_16763,N_16928);
xnor U17195 (N_17195,N_16907,N_16871);
and U17196 (N_17196,N_16974,N_16903);
or U17197 (N_17197,N_16804,N_16905);
nand U17198 (N_17198,N_16781,N_16906);
nor U17199 (N_17199,N_16826,N_16807);
and U17200 (N_17200,N_16772,N_16923);
xor U17201 (N_17201,N_16824,N_16917);
and U17202 (N_17202,N_16848,N_16941);
nand U17203 (N_17203,N_16971,N_16750);
and U17204 (N_17204,N_16841,N_16969);
nor U17205 (N_17205,N_16831,N_16868);
xnor U17206 (N_17206,N_16769,N_16932);
nor U17207 (N_17207,N_16847,N_16882);
xor U17208 (N_17208,N_16822,N_16869);
xor U17209 (N_17209,N_16770,N_16877);
xnor U17210 (N_17210,N_16765,N_16965);
nand U17211 (N_17211,N_16905,N_16862);
xor U17212 (N_17212,N_16961,N_16932);
nand U17213 (N_17213,N_16839,N_16991);
or U17214 (N_17214,N_16813,N_16854);
nor U17215 (N_17215,N_16921,N_16750);
or U17216 (N_17216,N_16913,N_16892);
nor U17217 (N_17217,N_16811,N_16884);
nor U17218 (N_17218,N_16949,N_16828);
xnor U17219 (N_17219,N_16750,N_16999);
nand U17220 (N_17220,N_16844,N_16984);
xnor U17221 (N_17221,N_16969,N_16821);
xor U17222 (N_17222,N_16918,N_16990);
xnor U17223 (N_17223,N_16940,N_16770);
or U17224 (N_17224,N_16950,N_16862);
xnor U17225 (N_17225,N_16922,N_16941);
or U17226 (N_17226,N_16867,N_16876);
or U17227 (N_17227,N_16969,N_16760);
nand U17228 (N_17228,N_16933,N_16926);
nor U17229 (N_17229,N_16808,N_16849);
nor U17230 (N_17230,N_16788,N_16892);
or U17231 (N_17231,N_16878,N_16956);
and U17232 (N_17232,N_16827,N_16974);
nor U17233 (N_17233,N_16948,N_16797);
nor U17234 (N_17234,N_16816,N_16843);
nand U17235 (N_17235,N_16917,N_16998);
nor U17236 (N_17236,N_16974,N_16882);
xnor U17237 (N_17237,N_16987,N_16844);
and U17238 (N_17238,N_16903,N_16888);
nor U17239 (N_17239,N_16771,N_16869);
and U17240 (N_17240,N_16996,N_16984);
xor U17241 (N_17241,N_16772,N_16829);
xnor U17242 (N_17242,N_16946,N_16939);
nor U17243 (N_17243,N_16830,N_16804);
xnor U17244 (N_17244,N_16757,N_16969);
xor U17245 (N_17245,N_16773,N_16907);
nor U17246 (N_17246,N_16912,N_16934);
nand U17247 (N_17247,N_16929,N_16839);
or U17248 (N_17248,N_16847,N_16872);
and U17249 (N_17249,N_16801,N_16827);
nand U17250 (N_17250,N_17071,N_17028);
or U17251 (N_17251,N_17099,N_17031);
xor U17252 (N_17252,N_17013,N_17107);
and U17253 (N_17253,N_17244,N_17236);
nor U17254 (N_17254,N_17082,N_17232);
and U17255 (N_17255,N_17227,N_17179);
nand U17256 (N_17256,N_17027,N_17036);
nor U17257 (N_17257,N_17170,N_17194);
and U17258 (N_17258,N_17054,N_17133);
and U17259 (N_17259,N_17122,N_17080);
nor U17260 (N_17260,N_17212,N_17016);
or U17261 (N_17261,N_17172,N_17109);
xnor U17262 (N_17262,N_17238,N_17117);
or U17263 (N_17263,N_17022,N_17111);
nor U17264 (N_17264,N_17011,N_17216);
xnor U17265 (N_17265,N_17202,N_17229);
or U17266 (N_17266,N_17167,N_17168);
xor U17267 (N_17267,N_17088,N_17035);
nor U17268 (N_17268,N_17215,N_17019);
or U17269 (N_17269,N_17075,N_17199);
xor U17270 (N_17270,N_17131,N_17037);
nand U17271 (N_17271,N_17151,N_17164);
and U17272 (N_17272,N_17163,N_17145);
and U17273 (N_17273,N_17120,N_17073);
nand U17274 (N_17274,N_17051,N_17079);
nor U17275 (N_17275,N_17030,N_17014);
xor U17276 (N_17276,N_17039,N_17192);
nand U17277 (N_17277,N_17091,N_17137);
or U17278 (N_17278,N_17057,N_17032);
or U17279 (N_17279,N_17041,N_17144);
xnor U17280 (N_17280,N_17042,N_17113);
nor U17281 (N_17281,N_17095,N_17147);
or U17282 (N_17282,N_17115,N_17094);
nand U17283 (N_17283,N_17235,N_17093);
or U17284 (N_17284,N_17004,N_17006);
and U17285 (N_17285,N_17247,N_17204);
and U17286 (N_17286,N_17070,N_17024);
and U17287 (N_17287,N_17017,N_17210);
xor U17288 (N_17288,N_17203,N_17092);
nor U17289 (N_17289,N_17208,N_17052);
or U17290 (N_17290,N_17062,N_17007);
and U17291 (N_17291,N_17118,N_17184);
and U17292 (N_17292,N_17124,N_17034);
nor U17293 (N_17293,N_17008,N_17101);
xor U17294 (N_17294,N_17178,N_17197);
nor U17295 (N_17295,N_17181,N_17249);
xnor U17296 (N_17296,N_17000,N_17018);
nor U17297 (N_17297,N_17200,N_17185);
xor U17298 (N_17298,N_17020,N_17048);
xor U17299 (N_17299,N_17242,N_17023);
nor U17300 (N_17300,N_17043,N_17174);
nand U17301 (N_17301,N_17159,N_17241);
xor U17302 (N_17302,N_17246,N_17045);
and U17303 (N_17303,N_17096,N_17127);
and U17304 (N_17304,N_17029,N_17047);
nand U17305 (N_17305,N_17155,N_17191);
nand U17306 (N_17306,N_17050,N_17165);
nand U17307 (N_17307,N_17003,N_17220);
or U17308 (N_17308,N_17044,N_17106);
nor U17309 (N_17309,N_17234,N_17195);
nor U17310 (N_17310,N_17056,N_17245);
and U17311 (N_17311,N_17143,N_17160);
nor U17312 (N_17312,N_17128,N_17012);
nand U17313 (N_17313,N_17121,N_17136);
xnor U17314 (N_17314,N_17169,N_17105);
or U17315 (N_17315,N_17112,N_17066);
or U17316 (N_17316,N_17207,N_17058);
or U17317 (N_17317,N_17223,N_17065);
or U17318 (N_17318,N_17214,N_17140);
and U17319 (N_17319,N_17108,N_17193);
or U17320 (N_17320,N_17221,N_17243);
xor U17321 (N_17321,N_17248,N_17205);
nor U17322 (N_17322,N_17190,N_17084);
and U17323 (N_17323,N_17153,N_17150);
xor U17324 (N_17324,N_17177,N_17240);
and U17325 (N_17325,N_17069,N_17175);
xnor U17326 (N_17326,N_17089,N_17157);
and U17327 (N_17327,N_17219,N_17225);
and U17328 (N_17328,N_17224,N_17110);
nor U17329 (N_17329,N_17100,N_17010);
and U17330 (N_17330,N_17156,N_17116);
and U17331 (N_17331,N_17049,N_17123);
nor U17332 (N_17332,N_17217,N_17083);
nor U17333 (N_17333,N_17125,N_17187);
xnor U17334 (N_17334,N_17218,N_17040);
nand U17335 (N_17335,N_17138,N_17228);
nor U17336 (N_17336,N_17149,N_17186);
nand U17337 (N_17337,N_17076,N_17188);
and U17338 (N_17338,N_17237,N_17072);
nor U17339 (N_17339,N_17090,N_17103);
or U17340 (N_17340,N_17183,N_17213);
xnor U17341 (N_17341,N_17162,N_17114);
or U17342 (N_17342,N_17139,N_17129);
or U17343 (N_17343,N_17055,N_17158);
and U17344 (N_17344,N_17005,N_17209);
and U17345 (N_17345,N_17211,N_17196);
nand U17346 (N_17346,N_17231,N_17002);
and U17347 (N_17347,N_17053,N_17239);
and U17348 (N_17348,N_17189,N_17135);
xnor U17349 (N_17349,N_17074,N_17009);
xor U17350 (N_17350,N_17226,N_17148);
and U17351 (N_17351,N_17126,N_17015);
or U17352 (N_17352,N_17142,N_17038);
nand U17353 (N_17353,N_17180,N_17102);
xnor U17354 (N_17354,N_17198,N_17061);
nor U17355 (N_17355,N_17182,N_17046);
nor U17356 (N_17356,N_17104,N_17201);
and U17357 (N_17357,N_17230,N_17026);
or U17358 (N_17358,N_17068,N_17025);
xnor U17359 (N_17359,N_17087,N_17081);
and U17360 (N_17360,N_17021,N_17033);
xor U17361 (N_17361,N_17166,N_17060);
nor U17362 (N_17362,N_17097,N_17134);
xnor U17363 (N_17363,N_17233,N_17206);
and U17364 (N_17364,N_17001,N_17130);
xnor U17365 (N_17365,N_17141,N_17078);
and U17366 (N_17366,N_17086,N_17161);
and U17367 (N_17367,N_17132,N_17085);
nor U17368 (N_17368,N_17067,N_17063);
xor U17369 (N_17369,N_17146,N_17173);
nand U17370 (N_17370,N_17119,N_17171);
nand U17371 (N_17371,N_17152,N_17176);
nand U17372 (N_17372,N_17098,N_17059);
nand U17373 (N_17373,N_17064,N_17154);
or U17374 (N_17374,N_17077,N_17222);
or U17375 (N_17375,N_17220,N_17158);
nand U17376 (N_17376,N_17143,N_17078);
nor U17377 (N_17377,N_17211,N_17108);
nand U17378 (N_17378,N_17187,N_17178);
or U17379 (N_17379,N_17176,N_17066);
and U17380 (N_17380,N_17179,N_17125);
xnor U17381 (N_17381,N_17081,N_17002);
or U17382 (N_17382,N_17107,N_17081);
or U17383 (N_17383,N_17193,N_17180);
xnor U17384 (N_17384,N_17227,N_17231);
nor U17385 (N_17385,N_17044,N_17155);
xnor U17386 (N_17386,N_17009,N_17174);
xor U17387 (N_17387,N_17137,N_17085);
xor U17388 (N_17388,N_17234,N_17186);
xor U17389 (N_17389,N_17056,N_17036);
nand U17390 (N_17390,N_17238,N_17118);
and U17391 (N_17391,N_17174,N_17094);
and U17392 (N_17392,N_17124,N_17210);
xnor U17393 (N_17393,N_17240,N_17012);
xor U17394 (N_17394,N_17050,N_17065);
xor U17395 (N_17395,N_17163,N_17230);
and U17396 (N_17396,N_17075,N_17122);
and U17397 (N_17397,N_17049,N_17202);
nand U17398 (N_17398,N_17022,N_17206);
nor U17399 (N_17399,N_17100,N_17211);
and U17400 (N_17400,N_17179,N_17055);
xor U17401 (N_17401,N_17211,N_17053);
and U17402 (N_17402,N_17038,N_17116);
nand U17403 (N_17403,N_17209,N_17065);
and U17404 (N_17404,N_17028,N_17108);
or U17405 (N_17405,N_17135,N_17034);
and U17406 (N_17406,N_17194,N_17134);
xor U17407 (N_17407,N_17003,N_17158);
nand U17408 (N_17408,N_17000,N_17103);
nor U17409 (N_17409,N_17170,N_17164);
and U17410 (N_17410,N_17180,N_17050);
or U17411 (N_17411,N_17247,N_17124);
or U17412 (N_17412,N_17135,N_17071);
nand U17413 (N_17413,N_17191,N_17070);
or U17414 (N_17414,N_17199,N_17240);
nand U17415 (N_17415,N_17119,N_17107);
nor U17416 (N_17416,N_17233,N_17187);
xnor U17417 (N_17417,N_17062,N_17152);
xnor U17418 (N_17418,N_17026,N_17057);
and U17419 (N_17419,N_17135,N_17021);
xnor U17420 (N_17420,N_17188,N_17145);
and U17421 (N_17421,N_17227,N_17069);
xnor U17422 (N_17422,N_17136,N_17020);
or U17423 (N_17423,N_17033,N_17241);
and U17424 (N_17424,N_17005,N_17183);
nor U17425 (N_17425,N_17153,N_17039);
or U17426 (N_17426,N_17144,N_17225);
and U17427 (N_17427,N_17242,N_17064);
xor U17428 (N_17428,N_17127,N_17227);
nand U17429 (N_17429,N_17093,N_17233);
nand U17430 (N_17430,N_17136,N_17033);
or U17431 (N_17431,N_17008,N_17049);
or U17432 (N_17432,N_17062,N_17039);
nor U17433 (N_17433,N_17249,N_17246);
or U17434 (N_17434,N_17164,N_17195);
and U17435 (N_17435,N_17111,N_17160);
or U17436 (N_17436,N_17190,N_17141);
nor U17437 (N_17437,N_17205,N_17107);
nand U17438 (N_17438,N_17244,N_17189);
or U17439 (N_17439,N_17088,N_17192);
or U17440 (N_17440,N_17164,N_17059);
or U17441 (N_17441,N_17237,N_17114);
and U17442 (N_17442,N_17110,N_17019);
xnor U17443 (N_17443,N_17174,N_17018);
xnor U17444 (N_17444,N_17242,N_17142);
and U17445 (N_17445,N_17024,N_17120);
xnor U17446 (N_17446,N_17185,N_17077);
and U17447 (N_17447,N_17101,N_17052);
nor U17448 (N_17448,N_17060,N_17206);
nor U17449 (N_17449,N_17046,N_17168);
and U17450 (N_17450,N_17184,N_17080);
nand U17451 (N_17451,N_17124,N_17234);
and U17452 (N_17452,N_17013,N_17087);
nand U17453 (N_17453,N_17128,N_17187);
nor U17454 (N_17454,N_17188,N_17016);
or U17455 (N_17455,N_17207,N_17067);
or U17456 (N_17456,N_17204,N_17145);
xnor U17457 (N_17457,N_17236,N_17211);
nand U17458 (N_17458,N_17191,N_17036);
nor U17459 (N_17459,N_17009,N_17098);
xnor U17460 (N_17460,N_17195,N_17208);
xor U17461 (N_17461,N_17228,N_17166);
or U17462 (N_17462,N_17216,N_17208);
nand U17463 (N_17463,N_17178,N_17150);
xnor U17464 (N_17464,N_17192,N_17103);
nor U17465 (N_17465,N_17035,N_17207);
nor U17466 (N_17466,N_17086,N_17053);
nand U17467 (N_17467,N_17085,N_17187);
and U17468 (N_17468,N_17137,N_17126);
xor U17469 (N_17469,N_17058,N_17190);
nand U17470 (N_17470,N_17231,N_17149);
nor U17471 (N_17471,N_17227,N_17089);
and U17472 (N_17472,N_17145,N_17192);
xnor U17473 (N_17473,N_17018,N_17067);
or U17474 (N_17474,N_17235,N_17069);
and U17475 (N_17475,N_17193,N_17040);
or U17476 (N_17476,N_17091,N_17047);
or U17477 (N_17477,N_17071,N_17155);
nor U17478 (N_17478,N_17124,N_17037);
xnor U17479 (N_17479,N_17187,N_17077);
xnor U17480 (N_17480,N_17052,N_17029);
nand U17481 (N_17481,N_17121,N_17059);
nor U17482 (N_17482,N_17072,N_17084);
and U17483 (N_17483,N_17084,N_17024);
nand U17484 (N_17484,N_17185,N_17004);
xnor U17485 (N_17485,N_17048,N_17121);
nor U17486 (N_17486,N_17120,N_17092);
xnor U17487 (N_17487,N_17200,N_17075);
and U17488 (N_17488,N_17205,N_17112);
or U17489 (N_17489,N_17018,N_17119);
or U17490 (N_17490,N_17165,N_17116);
or U17491 (N_17491,N_17138,N_17061);
nand U17492 (N_17492,N_17006,N_17208);
nand U17493 (N_17493,N_17034,N_17088);
xor U17494 (N_17494,N_17151,N_17200);
and U17495 (N_17495,N_17031,N_17098);
xor U17496 (N_17496,N_17012,N_17033);
and U17497 (N_17497,N_17013,N_17010);
xnor U17498 (N_17498,N_17119,N_17082);
and U17499 (N_17499,N_17142,N_17163);
xor U17500 (N_17500,N_17457,N_17365);
nand U17501 (N_17501,N_17319,N_17477);
or U17502 (N_17502,N_17422,N_17333);
or U17503 (N_17503,N_17262,N_17356);
or U17504 (N_17504,N_17466,N_17468);
xnor U17505 (N_17505,N_17346,N_17398);
xor U17506 (N_17506,N_17251,N_17412);
or U17507 (N_17507,N_17417,N_17261);
xor U17508 (N_17508,N_17476,N_17275);
or U17509 (N_17509,N_17350,N_17304);
xnor U17510 (N_17510,N_17371,N_17306);
nor U17511 (N_17511,N_17458,N_17462);
xor U17512 (N_17512,N_17443,N_17393);
nor U17513 (N_17513,N_17380,N_17258);
nor U17514 (N_17514,N_17452,N_17354);
xor U17515 (N_17515,N_17449,N_17447);
or U17516 (N_17516,N_17439,N_17271);
and U17517 (N_17517,N_17483,N_17289);
nand U17518 (N_17518,N_17392,N_17499);
and U17519 (N_17519,N_17423,N_17397);
xor U17520 (N_17520,N_17484,N_17283);
nor U17521 (N_17521,N_17292,N_17385);
and U17522 (N_17522,N_17363,N_17268);
and U17523 (N_17523,N_17311,N_17294);
and U17524 (N_17524,N_17374,N_17366);
and U17525 (N_17525,N_17470,N_17254);
xnor U17526 (N_17526,N_17314,N_17345);
or U17527 (N_17527,N_17303,N_17302);
nand U17528 (N_17528,N_17485,N_17436);
nand U17529 (N_17529,N_17322,N_17373);
or U17530 (N_17530,N_17433,N_17370);
nand U17531 (N_17531,N_17325,N_17253);
nor U17532 (N_17532,N_17324,N_17432);
xnor U17533 (N_17533,N_17344,N_17478);
xor U17534 (N_17534,N_17358,N_17493);
and U17535 (N_17535,N_17390,N_17342);
xor U17536 (N_17536,N_17479,N_17286);
and U17537 (N_17537,N_17329,N_17274);
or U17538 (N_17538,N_17475,N_17353);
and U17539 (N_17539,N_17320,N_17280);
or U17540 (N_17540,N_17288,N_17343);
nor U17541 (N_17541,N_17307,N_17260);
and U17542 (N_17542,N_17265,N_17317);
nand U17543 (N_17543,N_17362,N_17386);
nor U17544 (N_17544,N_17308,N_17339);
and U17545 (N_17545,N_17338,N_17347);
nand U17546 (N_17546,N_17349,N_17318);
and U17547 (N_17547,N_17418,N_17402);
nor U17548 (N_17548,N_17357,N_17377);
xnor U17549 (N_17549,N_17263,N_17336);
nand U17550 (N_17550,N_17473,N_17420);
or U17551 (N_17551,N_17267,N_17332);
nor U17552 (N_17552,N_17472,N_17257);
or U17553 (N_17553,N_17327,N_17293);
and U17554 (N_17554,N_17299,N_17467);
and U17555 (N_17555,N_17295,N_17351);
nand U17556 (N_17556,N_17471,N_17376);
nor U17557 (N_17557,N_17388,N_17456);
nand U17558 (N_17558,N_17334,N_17360);
xnor U17559 (N_17559,N_17448,N_17284);
and U17560 (N_17560,N_17369,N_17413);
xor U17561 (N_17561,N_17340,N_17469);
nand U17562 (N_17562,N_17463,N_17312);
xor U17563 (N_17563,N_17434,N_17375);
or U17564 (N_17564,N_17273,N_17282);
or U17565 (N_17565,N_17330,N_17438);
or U17566 (N_17566,N_17498,N_17269);
nor U17567 (N_17567,N_17429,N_17446);
nand U17568 (N_17568,N_17291,N_17450);
and U17569 (N_17569,N_17337,N_17278);
nor U17570 (N_17570,N_17427,N_17321);
nor U17571 (N_17571,N_17415,N_17464);
and U17572 (N_17572,N_17444,N_17445);
xor U17573 (N_17573,N_17297,N_17272);
and U17574 (N_17574,N_17255,N_17394);
xor U17575 (N_17575,N_17480,N_17454);
nand U17576 (N_17576,N_17313,N_17474);
nand U17577 (N_17577,N_17451,N_17400);
nand U17578 (N_17578,N_17409,N_17379);
or U17579 (N_17579,N_17378,N_17287);
nor U17580 (N_17580,N_17431,N_17492);
and U17581 (N_17581,N_17410,N_17323);
nor U17582 (N_17582,N_17411,N_17406);
and U17583 (N_17583,N_17465,N_17355);
nor U17584 (N_17584,N_17316,N_17270);
nand U17585 (N_17585,N_17488,N_17487);
nand U17586 (N_17586,N_17437,N_17399);
and U17587 (N_17587,N_17486,N_17326);
or U17588 (N_17588,N_17368,N_17404);
nand U17589 (N_17589,N_17305,N_17279);
and U17590 (N_17590,N_17300,N_17309);
xor U17591 (N_17591,N_17348,N_17364);
xnor U17592 (N_17592,N_17416,N_17264);
or U17593 (N_17593,N_17494,N_17426);
xor U17594 (N_17594,N_17331,N_17252);
or U17595 (N_17595,N_17256,N_17442);
or U17596 (N_17596,N_17405,N_17381);
and U17597 (N_17597,N_17315,N_17341);
xnor U17598 (N_17598,N_17395,N_17335);
or U17599 (N_17599,N_17461,N_17396);
xnor U17600 (N_17600,N_17310,N_17391);
xor U17601 (N_17601,N_17407,N_17290);
nand U17602 (N_17602,N_17497,N_17481);
and U17603 (N_17603,N_17459,N_17361);
nand U17604 (N_17604,N_17440,N_17482);
xnor U17605 (N_17605,N_17352,N_17453);
xor U17606 (N_17606,N_17301,N_17383);
and U17607 (N_17607,N_17384,N_17489);
and U17608 (N_17608,N_17372,N_17428);
and U17609 (N_17609,N_17425,N_17328);
nor U17610 (N_17610,N_17285,N_17276);
or U17611 (N_17611,N_17259,N_17491);
nor U17612 (N_17612,N_17382,N_17298);
xnor U17613 (N_17613,N_17389,N_17460);
xor U17614 (N_17614,N_17266,N_17421);
nand U17615 (N_17615,N_17495,N_17430);
nand U17616 (N_17616,N_17496,N_17367);
nand U17617 (N_17617,N_17277,N_17296);
nand U17618 (N_17618,N_17490,N_17408);
or U17619 (N_17619,N_17403,N_17441);
and U17620 (N_17620,N_17250,N_17387);
xnor U17621 (N_17621,N_17424,N_17281);
or U17622 (N_17622,N_17414,N_17359);
nor U17623 (N_17623,N_17401,N_17419);
nand U17624 (N_17624,N_17435,N_17455);
and U17625 (N_17625,N_17281,N_17379);
and U17626 (N_17626,N_17481,N_17260);
and U17627 (N_17627,N_17285,N_17445);
nor U17628 (N_17628,N_17411,N_17306);
xnor U17629 (N_17629,N_17309,N_17419);
and U17630 (N_17630,N_17380,N_17261);
or U17631 (N_17631,N_17453,N_17413);
nor U17632 (N_17632,N_17391,N_17373);
nand U17633 (N_17633,N_17273,N_17383);
xnor U17634 (N_17634,N_17449,N_17299);
or U17635 (N_17635,N_17415,N_17301);
and U17636 (N_17636,N_17489,N_17368);
and U17637 (N_17637,N_17438,N_17251);
or U17638 (N_17638,N_17297,N_17465);
xor U17639 (N_17639,N_17480,N_17335);
nand U17640 (N_17640,N_17334,N_17292);
nor U17641 (N_17641,N_17291,N_17297);
or U17642 (N_17642,N_17474,N_17404);
or U17643 (N_17643,N_17375,N_17349);
nand U17644 (N_17644,N_17447,N_17278);
nand U17645 (N_17645,N_17253,N_17276);
xor U17646 (N_17646,N_17474,N_17303);
and U17647 (N_17647,N_17403,N_17494);
and U17648 (N_17648,N_17299,N_17428);
xnor U17649 (N_17649,N_17485,N_17263);
xor U17650 (N_17650,N_17479,N_17285);
xnor U17651 (N_17651,N_17274,N_17262);
and U17652 (N_17652,N_17371,N_17393);
and U17653 (N_17653,N_17422,N_17377);
xor U17654 (N_17654,N_17316,N_17419);
or U17655 (N_17655,N_17438,N_17252);
and U17656 (N_17656,N_17394,N_17496);
xnor U17657 (N_17657,N_17431,N_17438);
and U17658 (N_17658,N_17423,N_17470);
nor U17659 (N_17659,N_17363,N_17359);
nand U17660 (N_17660,N_17440,N_17285);
nor U17661 (N_17661,N_17351,N_17291);
and U17662 (N_17662,N_17315,N_17323);
or U17663 (N_17663,N_17292,N_17451);
or U17664 (N_17664,N_17261,N_17300);
xnor U17665 (N_17665,N_17494,N_17301);
nand U17666 (N_17666,N_17358,N_17478);
nand U17667 (N_17667,N_17458,N_17400);
xor U17668 (N_17668,N_17316,N_17394);
nor U17669 (N_17669,N_17335,N_17469);
nand U17670 (N_17670,N_17472,N_17485);
or U17671 (N_17671,N_17463,N_17409);
and U17672 (N_17672,N_17484,N_17486);
and U17673 (N_17673,N_17439,N_17438);
or U17674 (N_17674,N_17371,N_17399);
nor U17675 (N_17675,N_17453,N_17277);
nand U17676 (N_17676,N_17389,N_17417);
xnor U17677 (N_17677,N_17296,N_17493);
or U17678 (N_17678,N_17391,N_17351);
and U17679 (N_17679,N_17360,N_17354);
nand U17680 (N_17680,N_17290,N_17383);
nor U17681 (N_17681,N_17479,N_17432);
and U17682 (N_17682,N_17263,N_17400);
nand U17683 (N_17683,N_17396,N_17364);
and U17684 (N_17684,N_17386,N_17412);
and U17685 (N_17685,N_17290,N_17449);
or U17686 (N_17686,N_17468,N_17297);
nor U17687 (N_17687,N_17392,N_17361);
nor U17688 (N_17688,N_17283,N_17351);
xnor U17689 (N_17689,N_17289,N_17274);
nand U17690 (N_17690,N_17471,N_17469);
and U17691 (N_17691,N_17459,N_17299);
and U17692 (N_17692,N_17481,N_17376);
and U17693 (N_17693,N_17382,N_17277);
nor U17694 (N_17694,N_17256,N_17347);
and U17695 (N_17695,N_17430,N_17274);
nor U17696 (N_17696,N_17443,N_17286);
or U17697 (N_17697,N_17310,N_17485);
xor U17698 (N_17698,N_17437,N_17381);
or U17699 (N_17699,N_17497,N_17393);
or U17700 (N_17700,N_17269,N_17270);
nand U17701 (N_17701,N_17413,N_17405);
xor U17702 (N_17702,N_17411,N_17430);
or U17703 (N_17703,N_17370,N_17298);
xnor U17704 (N_17704,N_17416,N_17369);
or U17705 (N_17705,N_17366,N_17476);
nand U17706 (N_17706,N_17475,N_17309);
xor U17707 (N_17707,N_17252,N_17364);
nand U17708 (N_17708,N_17370,N_17400);
or U17709 (N_17709,N_17435,N_17353);
xnor U17710 (N_17710,N_17484,N_17258);
nor U17711 (N_17711,N_17496,N_17395);
and U17712 (N_17712,N_17394,N_17411);
xor U17713 (N_17713,N_17474,N_17266);
nor U17714 (N_17714,N_17416,N_17314);
and U17715 (N_17715,N_17327,N_17478);
nor U17716 (N_17716,N_17384,N_17347);
nand U17717 (N_17717,N_17412,N_17260);
or U17718 (N_17718,N_17445,N_17263);
nand U17719 (N_17719,N_17296,N_17372);
xor U17720 (N_17720,N_17469,N_17311);
xor U17721 (N_17721,N_17367,N_17308);
or U17722 (N_17722,N_17387,N_17480);
nand U17723 (N_17723,N_17350,N_17386);
nor U17724 (N_17724,N_17322,N_17428);
xnor U17725 (N_17725,N_17258,N_17476);
xor U17726 (N_17726,N_17278,N_17391);
xnor U17727 (N_17727,N_17486,N_17458);
or U17728 (N_17728,N_17407,N_17405);
and U17729 (N_17729,N_17348,N_17391);
nand U17730 (N_17730,N_17335,N_17315);
nand U17731 (N_17731,N_17350,N_17404);
nor U17732 (N_17732,N_17285,N_17346);
xor U17733 (N_17733,N_17302,N_17415);
xnor U17734 (N_17734,N_17294,N_17470);
and U17735 (N_17735,N_17293,N_17411);
nor U17736 (N_17736,N_17414,N_17347);
xor U17737 (N_17737,N_17400,N_17295);
xnor U17738 (N_17738,N_17390,N_17346);
xnor U17739 (N_17739,N_17450,N_17398);
or U17740 (N_17740,N_17378,N_17354);
nand U17741 (N_17741,N_17478,N_17413);
nor U17742 (N_17742,N_17322,N_17251);
nand U17743 (N_17743,N_17393,N_17394);
nor U17744 (N_17744,N_17293,N_17271);
nor U17745 (N_17745,N_17456,N_17264);
nor U17746 (N_17746,N_17337,N_17386);
or U17747 (N_17747,N_17428,N_17258);
and U17748 (N_17748,N_17316,N_17475);
nand U17749 (N_17749,N_17334,N_17463);
xnor U17750 (N_17750,N_17686,N_17745);
xnor U17751 (N_17751,N_17659,N_17657);
and U17752 (N_17752,N_17719,N_17520);
and U17753 (N_17753,N_17566,N_17557);
xnor U17754 (N_17754,N_17621,N_17727);
nand U17755 (N_17755,N_17718,N_17548);
nand U17756 (N_17756,N_17635,N_17724);
nor U17757 (N_17757,N_17558,N_17681);
xor U17758 (N_17758,N_17533,N_17600);
nand U17759 (N_17759,N_17511,N_17714);
or U17760 (N_17760,N_17679,N_17666);
and U17761 (N_17761,N_17656,N_17601);
and U17762 (N_17762,N_17532,N_17609);
or U17763 (N_17763,N_17623,N_17583);
nor U17764 (N_17764,N_17704,N_17651);
or U17765 (N_17765,N_17603,N_17574);
xor U17766 (N_17766,N_17720,N_17709);
and U17767 (N_17767,N_17508,N_17652);
nand U17768 (N_17768,N_17604,N_17747);
and U17769 (N_17769,N_17605,N_17692);
xnor U17770 (N_17770,N_17564,N_17700);
and U17771 (N_17771,N_17640,N_17741);
or U17772 (N_17772,N_17726,N_17694);
or U17773 (N_17773,N_17544,N_17626);
and U17774 (N_17774,N_17671,N_17575);
and U17775 (N_17775,N_17644,N_17586);
nor U17776 (N_17776,N_17736,N_17639);
xnor U17777 (N_17777,N_17592,N_17665);
nand U17778 (N_17778,N_17573,N_17742);
xnor U17779 (N_17779,N_17624,N_17530);
or U17780 (N_17780,N_17569,N_17571);
and U17781 (N_17781,N_17632,N_17510);
or U17782 (N_17782,N_17570,N_17509);
xnor U17783 (N_17783,N_17534,N_17588);
or U17784 (N_17784,N_17585,N_17687);
and U17785 (N_17785,N_17522,N_17634);
xnor U17786 (N_17786,N_17563,N_17645);
xnor U17787 (N_17787,N_17501,N_17646);
xor U17788 (N_17788,N_17521,N_17734);
or U17789 (N_17789,N_17662,N_17721);
and U17790 (N_17790,N_17708,N_17518);
xor U17791 (N_17791,N_17680,N_17608);
nor U17792 (N_17792,N_17673,N_17581);
or U17793 (N_17793,N_17744,N_17531);
nor U17794 (N_17794,N_17589,N_17560);
nor U17795 (N_17795,N_17732,N_17684);
or U17796 (N_17796,N_17553,N_17636);
or U17797 (N_17797,N_17660,N_17504);
nand U17798 (N_17798,N_17715,N_17688);
or U17799 (N_17799,N_17554,N_17703);
nand U17800 (N_17800,N_17716,N_17723);
or U17801 (N_17801,N_17528,N_17722);
nand U17802 (N_17802,N_17713,N_17625);
and U17803 (N_17803,N_17540,N_17587);
xnor U17804 (N_17804,N_17582,N_17593);
nand U17805 (N_17805,N_17706,N_17606);
or U17806 (N_17806,N_17539,N_17678);
and U17807 (N_17807,N_17629,N_17602);
nor U17808 (N_17808,N_17641,N_17670);
or U17809 (N_17809,N_17515,N_17561);
and U17810 (N_17810,N_17505,N_17572);
and U17811 (N_17811,N_17682,N_17523);
and U17812 (N_17812,N_17630,N_17565);
nor U17813 (N_17813,N_17730,N_17507);
or U17814 (N_17814,N_17697,N_17567);
nand U17815 (N_17815,N_17705,N_17696);
xnor U17816 (N_17816,N_17611,N_17546);
nand U17817 (N_17817,N_17578,N_17710);
or U17818 (N_17818,N_17607,N_17595);
nor U17819 (N_17819,N_17695,N_17535);
or U17820 (N_17820,N_17517,N_17690);
and U17821 (N_17821,N_17672,N_17576);
or U17822 (N_17822,N_17503,N_17537);
xor U17823 (N_17823,N_17525,N_17739);
nor U17824 (N_17824,N_17619,N_17725);
and U17825 (N_17825,N_17516,N_17663);
and U17826 (N_17826,N_17617,N_17677);
xor U17827 (N_17827,N_17568,N_17735);
nor U17828 (N_17828,N_17702,N_17647);
nand U17829 (N_17829,N_17613,N_17514);
and U17830 (N_17830,N_17654,N_17731);
nand U17831 (N_17831,N_17599,N_17549);
nor U17832 (N_17832,N_17538,N_17614);
nor U17833 (N_17833,N_17661,N_17627);
nor U17834 (N_17834,N_17633,N_17683);
xnor U17835 (N_17835,N_17693,N_17685);
nor U17836 (N_17836,N_17650,N_17555);
nor U17837 (N_17837,N_17711,N_17653);
nor U17838 (N_17838,N_17598,N_17590);
nand U17839 (N_17839,N_17707,N_17618);
xnor U17840 (N_17840,N_17597,N_17664);
and U17841 (N_17841,N_17580,N_17676);
xnor U17842 (N_17842,N_17500,N_17596);
and U17843 (N_17843,N_17529,N_17701);
and U17844 (N_17844,N_17612,N_17551);
or U17845 (N_17845,N_17638,N_17674);
or U17846 (N_17846,N_17506,N_17628);
nor U17847 (N_17847,N_17728,N_17740);
nor U17848 (N_17848,N_17737,N_17591);
and U17849 (N_17849,N_17556,N_17552);
nor U17850 (N_17850,N_17543,N_17643);
nor U17851 (N_17851,N_17616,N_17668);
nor U17852 (N_17852,N_17655,N_17577);
nor U17853 (N_17853,N_17733,N_17649);
nor U17854 (N_17854,N_17648,N_17748);
nor U17855 (N_17855,N_17712,N_17689);
and U17856 (N_17856,N_17594,N_17579);
nand U17857 (N_17857,N_17637,N_17631);
nand U17858 (N_17858,N_17717,N_17746);
nor U17859 (N_17859,N_17658,N_17729);
nand U17860 (N_17860,N_17519,N_17527);
nand U17861 (N_17861,N_17502,N_17541);
xor U17862 (N_17862,N_17642,N_17526);
and U17863 (N_17863,N_17542,N_17669);
nand U17864 (N_17864,N_17545,N_17620);
or U17865 (N_17865,N_17536,N_17699);
or U17866 (N_17866,N_17667,N_17610);
xnor U17867 (N_17867,N_17524,N_17743);
xor U17868 (N_17868,N_17691,N_17622);
or U17869 (N_17869,N_17562,N_17698);
nand U17870 (N_17870,N_17675,N_17547);
and U17871 (N_17871,N_17559,N_17749);
or U17872 (N_17872,N_17550,N_17513);
or U17873 (N_17873,N_17584,N_17615);
or U17874 (N_17874,N_17512,N_17738);
and U17875 (N_17875,N_17559,N_17536);
or U17876 (N_17876,N_17646,N_17595);
and U17877 (N_17877,N_17613,N_17585);
nor U17878 (N_17878,N_17715,N_17668);
and U17879 (N_17879,N_17531,N_17601);
and U17880 (N_17880,N_17657,N_17704);
nand U17881 (N_17881,N_17627,N_17741);
xor U17882 (N_17882,N_17569,N_17574);
xnor U17883 (N_17883,N_17658,N_17684);
nor U17884 (N_17884,N_17549,N_17546);
nand U17885 (N_17885,N_17578,N_17732);
nor U17886 (N_17886,N_17726,N_17744);
xnor U17887 (N_17887,N_17671,N_17643);
nand U17888 (N_17888,N_17611,N_17559);
nand U17889 (N_17889,N_17533,N_17712);
or U17890 (N_17890,N_17508,N_17640);
nand U17891 (N_17891,N_17618,N_17657);
xor U17892 (N_17892,N_17504,N_17742);
and U17893 (N_17893,N_17562,N_17617);
or U17894 (N_17894,N_17714,N_17544);
and U17895 (N_17895,N_17699,N_17681);
xnor U17896 (N_17896,N_17721,N_17675);
and U17897 (N_17897,N_17699,N_17690);
and U17898 (N_17898,N_17695,N_17638);
nand U17899 (N_17899,N_17717,N_17725);
and U17900 (N_17900,N_17574,N_17711);
nand U17901 (N_17901,N_17527,N_17686);
xnor U17902 (N_17902,N_17744,N_17653);
and U17903 (N_17903,N_17628,N_17678);
or U17904 (N_17904,N_17732,N_17521);
or U17905 (N_17905,N_17531,N_17501);
xor U17906 (N_17906,N_17706,N_17628);
and U17907 (N_17907,N_17517,N_17700);
nand U17908 (N_17908,N_17645,N_17694);
nand U17909 (N_17909,N_17647,N_17605);
and U17910 (N_17910,N_17740,N_17706);
nor U17911 (N_17911,N_17715,N_17563);
xnor U17912 (N_17912,N_17636,N_17550);
nand U17913 (N_17913,N_17562,N_17629);
and U17914 (N_17914,N_17593,N_17744);
nand U17915 (N_17915,N_17675,N_17629);
xnor U17916 (N_17916,N_17655,N_17530);
nand U17917 (N_17917,N_17556,N_17535);
nor U17918 (N_17918,N_17746,N_17567);
or U17919 (N_17919,N_17551,N_17575);
xor U17920 (N_17920,N_17546,N_17729);
nand U17921 (N_17921,N_17694,N_17534);
xnor U17922 (N_17922,N_17559,N_17610);
xor U17923 (N_17923,N_17723,N_17589);
nor U17924 (N_17924,N_17711,N_17629);
nor U17925 (N_17925,N_17510,N_17670);
nand U17926 (N_17926,N_17537,N_17670);
or U17927 (N_17927,N_17558,N_17664);
or U17928 (N_17928,N_17522,N_17720);
nand U17929 (N_17929,N_17677,N_17600);
and U17930 (N_17930,N_17676,N_17696);
nor U17931 (N_17931,N_17608,N_17573);
xor U17932 (N_17932,N_17712,N_17634);
xor U17933 (N_17933,N_17664,N_17680);
and U17934 (N_17934,N_17724,N_17677);
or U17935 (N_17935,N_17710,N_17509);
nor U17936 (N_17936,N_17696,N_17584);
nand U17937 (N_17937,N_17543,N_17730);
nor U17938 (N_17938,N_17641,N_17721);
and U17939 (N_17939,N_17554,N_17594);
nand U17940 (N_17940,N_17571,N_17643);
or U17941 (N_17941,N_17569,N_17724);
nor U17942 (N_17942,N_17504,N_17508);
nor U17943 (N_17943,N_17697,N_17562);
nor U17944 (N_17944,N_17671,N_17535);
or U17945 (N_17945,N_17732,N_17705);
and U17946 (N_17946,N_17569,N_17743);
or U17947 (N_17947,N_17644,N_17507);
xnor U17948 (N_17948,N_17687,N_17536);
or U17949 (N_17949,N_17551,N_17659);
or U17950 (N_17950,N_17712,N_17559);
or U17951 (N_17951,N_17528,N_17560);
nor U17952 (N_17952,N_17652,N_17718);
and U17953 (N_17953,N_17712,N_17635);
nand U17954 (N_17954,N_17626,N_17673);
nor U17955 (N_17955,N_17699,N_17666);
and U17956 (N_17956,N_17588,N_17523);
xnor U17957 (N_17957,N_17511,N_17670);
nor U17958 (N_17958,N_17624,N_17660);
and U17959 (N_17959,N_17514,N_17745);
or U17960 (N_17960,N_17657,N_17702);
and U17961 (N_17961,N_17735,N_17695);
xor U17962 (N_17962,N_17648,N_17555);
or U17963 (N_17963,N_17703,N_17698);
xor U17964 (N_17964,N_17566,N_17622);
nor U17965 (N_17965,N_17507,N_17548);
nand U17966 (N_17966,N_17562,N_17564);
nor U17967 (N_17967,N_17639,N_17602);
nand U17968 (N_17968,N_17522,N_17568);
nor U17969 (N_17969,N_17555,N_17748);
nand U17970 (N_17970,N_17608,N_17633);
and U17971 (N_17971,N_17504,N_17595);
nor U17972 (N_17972,N_17677,N_17599);
and U17973 (N_17973,N_17547,N_17510);
and U17974 (N_17974,N_17596,N_17539);
xnor U17975 (N_17975,N_17723,N_17708);
xor U17976 (N_17976,N_17587,N_17523);
nor U17977 (N_17977,N_17656,N_17557);
or U17978 (N_17978,N_17690,N_17591);
or U17979 (N_17979,N_17598,N_17664);
nor U17980 (N_17980,N_17621,N_17588);
xnor U17981 (N_17981,N_17572,N_17576);
nor U17982 (N_17982,N_17511,N_17602);
nor U17983 (N_17983,N_17515,N_17568);
xnor U17984 (N_17984,N_17589,N_17689);
nand U17985 (N_17985,N_17520,N_17590);
xor U17986 (N_17986,N_17658,N_17502);
xor U17987 (N_17987,N_17603,N_17676);
or U17988 (N_17988,N_17531,N_17547);
nand U17989 (N_17989,N_17735,N_17606);
nor U17990 (N_17990,N_17627,N_17578);
nand U17991 (N_17991,N_17548,N_17601);
or U17992 (N_17992,N_17740,N_17722);
nand U17993 (N_17993,N_17683,N_17616);
nand U17994 (N_17994,N_17537,N_17521);
xnor U17995 (N_17995,N_17731,N_17569);
or U17996 (N_17996,N_17518,N_17728);
nor U17997 (N_17997,N_17701,N_17592);
nor U17998 (N_17998,N_17526,N_17608);
or U17999 (N_17999,N_17638,N_17531);
and U18000 (N_18000,N_17996,N_17896);
nor U18001 (N_18001,N_17760,N_17956);
or U18002 (N_18002,N_17950,N_17938);
nor U18003 (N_18003,N_17812,N_17759);
xnor U18004 (N_18004,N_17894,N_17977);
xnor U18005 (N_18005,N_17828,N_17786);
and U18006 (N_18006,N_17825,N_17832);
or U18007 (N_18007,N_17911,N_17919);
and U18008 (N_18008,N_17949,N_17936);
nor U18009 (N_18009,N_17978,N_17829);
or U18010 (N_18010,N_17973,N_17943);
nor U18011 (N_18011,N_17774,N_17816);
nor U18012 (N_18012,N_17903,N_17827);
and U18013 (N_18013,N_17927,N_17989);
xor U18014 (N_18014,N_17820,N_17854);
xnor U18015 (N_18015,N_17848,N_17803);
nor U18016 (N_18016,N_17758,N_17857);
or U18017 (N_18017,N_17859,N_17830);
or U18018 (N_18018,N_17966,N_17761);
or U18019 (N_18019,N_17775,N_17969);
nor U18020 (N_18020,N_17754,N_17844);
nor U18021 (N_18021,N_17778,N_17984);
nand U18022 (N_18022,N_17959,N_17779);
and U18023 (N_18023,N_17924,N_17841);
nand U18024 (N_18024,N_17809,N_17899);
or U18025 (N_18025,N_17751,N_17845);
nand U18026 (N_18026,N_17752,N_17842);
xnor U18027 (N_18027,N_17824,N_17791);
nand U18028 (N_18028,N_17815,N_17994);
and U18029 (N_18029,N_17930,N_17790);
nand U18030 (N_18030,N_17870,N_17921);
nand U18031 (N_18031,N_17990,N_17908);
nand U18032 (N_18032,N_17788,N_17783);
or U18033 (N_18033,N_17798,N_17850);
xnor U18034 (N_18034,N_17905,N_17819);
and U18035 (N_18035,N_17968,N_17757);
and U18036 (N_18036,N_17768,N_17856);
or U18037 (N_18037,N_17946,N_17954);
nand U18038 (N_18038,N_17887,N_17773);
nor U18039 (N_18039,N_17792,N_17861);
or U18040 (N_18040,N_17868,N_17878);
nand U18041 (N_18041,N_17869,N_17986);
xor U18042 (N_18042,N_17948,N_17886);
nand U18043 (N_18043,N_17982,N_17912);
or U18044 (N_18044,N_17953,N_17769);
nor U18045 (N_18045,N_17882,N_17764);
and U18046 (N_18046,N_17814,N_17895);
and U18047 (N_18047,N_17874,N_17811);
and U18048 (N_18048,N_17972,N_17897);
nor U18049 (N_18049,N_17767,N_17756);
nand U18050 (N_18050,N_17926,N_17916);
and U18051 (N_18051,N_17920,N_17780);
nor U18052 (N_18052,N_17822,N_17843);
nor U18053 (N_18053,N_17838,N_17913);
nor U18054 (N_18054,N_17917,N_17763);
nand U18055 (N_18055,N_17889,N_17907);
and U18056 (N_18056,N_17784,N_17823);
or U18057 (N_18057,N_17813,N_17960);
or U18058 (N_18058,N_17879,N_17902);
xnor U18059 (N_18059,N_17770,N_17952);
or U18060 (N_18060,N_17796,N_17955);
xor U18061 (N_18061,N_17964,N_17765);
and U18062 (N_18062,N_17835,N_17833);
and U18063 (N_18063,N_17962,N_17781);
xnor U18064 (N_18064,N_17890,N_17772);
or U18065 (N_18065,N_17925,N_17951);
and U18066 (N_18066,N_17993,N_17851);
and U18067 (N_18067,N_17928,N_17883);
or U18068 (N_18068,N_17834,N_17991);
nand U18069 (N_18069,N_17802,N_17863);
or U18070 (N_18070,N_17970,N_17942);
or U18071 (N_18071,N_17901,N_17817);
or U18072 (N_18072,N_17975,N_17777);
or U18073 (N_18073,N_17888,N_17983);
xnor U18074 (N_18074,N_17821,N_17846);
nand U18075 (N_18075,N_17876,N_17979);
and U18076 (N_18076,N_17914,N_17900);
or U18077 (N_18077,N_17875,N_17963);
nor U18078 (N_18078,N_17789,N_17836);
and U18079 (N_18079,N_17853,N_17794);
xor U18080 (N_18080,N_17957,N_17753);
nand U18081 (N_18081,N_17918,N_17818);
xor U18082 (N_18082,N_17871,N_17880);
nand U18083 (N_18083,N_17797,N_17947);
xor U18084 (N_18084,N_17800,N_17934);
xnor U18085 (N_18085,N_17945,N_17937);
and U18086 (N_18086,N_17933,N_17799);
nand U18087 (N_18087,N_17807,N_17961);
and U18088 (N_18088,N_17971,N_17785);
nor U18089 (N_18089,N_17755,N_17801);
nand U18090 (N_18090,N_17931,N_17847);
or U18091 (N_18091,N_17997,N_17965);
or U18092 (N_18092,N_17941,N_17929);
or U18093 (N_18093,N_17750,N_17992);
nor U18094 (N_18094,N_17795,N_17766);
nor U18095 (N_18095,N_17985,N_17771);
nor U18096 (N_18096,N_17776,N_17855);
and U18097 (N_18097,N_17839,N_17915);
xnor U18098 (N_18098,N_17885,N_17909);
and U18099 (N_18099,N_17849,N_17987);
and U18100 (N_18100,N_17884,N_17995);
nand U18101 (N_18101,N_17976,N_17998);
xor U18102 (N_18102,N_17958,N_17860);
nor U18103 (N_18103,N_17873,N_17762);
xor U18104 (N_18104,N_17906,N_17867);
or U18105 (N_18105,N_17980,N_17988);
xor U18106 (N_18106,N_17805,N_17852);
or U18107 (N_18107,N_17837,N_17944);
nor U18108 (N_18108,N_17881,N_17872);
xnor U18109 (N_18109,N_17967,N_17831);
or U18110 (N_18110,N_17940,N_17840);
xor U18111 (N_18111,N_17804,N_17865);
or U18112 (N_18112,N_17932,N_17864);
and U18113 (N_18113,N_17826,N_17893);
or U18114 (N_18114,N_17910,N_17782);
xor U18115 (N_18115,N_17922,N_17981);
nor U18116 (N_18116,N_17866,N_17923);
and U18117 (N_18117,N_17892,N_17891);
nor U18118 (N_18118,N_17862,N_17808);
and U18119 (N_18119,N_17877,N_17793);
nand U18120 (N_18120,N_17935,N_17974);
xnor U18121 (N_18121,N_17810,N_17898);
and U18122 (N_18122,N_17939,N_17858);
nor U18123 (N_18123,N_17787,N_17806);
nor U18124 (N_18124,N_17904,N_17999);
nor U18125 (N_18125,N_17781,N_17927);
and U18126 (N_18126,N_17984,N_17786);
xor U18127 (N_18127,N_17992,N_17946);
and U18128 (N_18128,N_17771,N_17872);
or U18129 (N_18129,N_17932,N_17841);
and U18130 (N_18130,N_17806,N_17939);
xnor U18131 (N_18131,N_17768,N_17758);
or U18132 (N_18132,N_17899,N_17779);
nand U18133 (N_18133,N_17929,N_17832);
and U18134 (N_18134,N_17847,N_17920);
or U18135 (N_18135,N_17974,N_17957);
xor U18136 (N_18136,N_17875,N_17907);
nor U18137 (N_18137,N_17780,N_17753);
or U18138 (N_18138,N_17846,N_17855);
nor U18139 (N_18139,N_17810,N_17786);
nand U18140 (N_18140,N_17760,N_17894);
or U18141 (N_18141,N_17993,N_17870);
nor U18142 (N_18142,N_17864,N_17868);
and U18143 (N_18143,N_17840,N_17846);
or U18144 (N_18144,N_17937,N_17997);
or U18145 (N_18145,N_17961,N_17951);
and U18146 (N_18146,N_17895,N_17778);
xnor U18147 (N_18147,N_17822,N_17945);
nand U18148 (N_18148,N_17779,N_17994);
xnor U18149 (N_18149,N_17850,N_17900);
or U18150 (N_18150,N_17936,N_17836);
and U18151 (N_18151,N_17860,N_17961);
or U18152 (N_18152,N_17813,N_17971);
and U18153 (N_18153,N_17873,N_17939);
and U18154 (N_18154,N_17885,N_17768);
xor U18155 (N_18155,N_17972,N_17955);
or U18156 (N_18156,N_17840,N_17819);
xor U18157 (N_18157,N_17858,N_17875);
or U18158 (N_18158,N_17897,N_17869);
nor U18159 (N_18159,N_17972,N_17880);
xor U18160 (N_18160,N_17755,N_17944);
or U18161 (N_18161,N_17790,N_17818);
nor U18162 (N_18162,N_17783,N_17838);
xor U18163 (N_18163,N_17770,N_17970);
and U18164 (N_18164,N_17993,N_17949);
xnor U18165 (N_18165,N_17922,N_17883);
xor U18166 (N_18166,N_17856,N_17853);
and U18167 (N_18167,N_17974,N_17796);
or U18168 (N_18168,N_17925,N_17920);
xnor U18169 (N_18169,N_17921,N_17899);
nand U18170 (N_18170,N_17835,N_17841);
nand U18171 (N_18171,N_17794,N_17758);
nor U18172 (N_18172,N_17998,N_17918);
or U18173 (N_18173,N_17963,N_17775);
nor U18174 (N_18174,N_17812,N_17985);
nor U18175 (N_18175,N_17840,N_17778);
nand U18176 (N_18176,N_17885,N_17969);
xor U18177 (N_18177,N_17820,N_17879);
xor U18178 (N_18178,N_17812,N_17906);
xnor U18179 (N_18179,N_17856,N_17996);
and U18180 (N_18180,N_17996,N_17875);
nand U18181 (N_18181,N_17905,N_17868);
and U18182 (N_18182,N_17775,N_17833);
nand U18183 (N_18183,N_17824,N_17771);
nand U18184 (N_18184,N_17897,N_17992);
nand U18185 (N_18185,N_17898,N_17865);
nand U18186 (N_18186,N_17926,N_17774);
nor U18187 (N_18187,N_17933,N_17954);
xnor U18188 (N_18188,N_17770,N_17775);
and U18189 (N_18189,N_17913,N_17987);
or U18190 (N_18190,N_17903,N_17964);
or U18191 (N_18191,N_17832,N_17806);
xnor U18192 (N_18192,N_17837,N_17965);
nand U18193 (N_18193,N_17883,N_17930);
and U18194 (N_18194,N_17788,N_17881);
nand U18195 (N_18195,N_17895,N_17958);
and U18196 (N_18196,N_17797,N_17758);
and U18197 (N_18197,N_17820,N_17948);
nand U18198 (N_18198,N_17884,N_17873);
or U18199 (N_18199,N_17902,N_17810);
nor U18200 (N_18200,N_17767,N_17819);
nor U18201 (N_18201,N_17835,N_17935);
nand U18202 (N_18202,N_17816,N_17975);
nor U18203 (N_18203,N_17975,N_17909);
and U18204 (N_18204,N_17881,N_17843);
or U18205 (N_18205,N_17847,N_17907);
xor U18206 (N_18206,N_17898,N_17772);
or U18207 (N_18207,N_17842,N_17770);
and U18208 (N_18208,N_17876,N_17835);
nand U18209 (N_18209,N_17894,N_17954);
xnor U18210 (N_18210,N_17753,N_17891);
xnor U18211 (N_18211,N_17802,N_17895);
nor U18212 (N_18212,N_17812,N_17858);
nand U18213 (N_18213,N_17843,N_17819);
xor U18214 (N_18214,N_17789,N_17758);
nor U18215 (N_18215,N_17927,N_17965);
nor U18216 (N_18216,N_17774,N_17789);
nor U18217 (N_18217,N_17906,N_17887);
nor U18218 (N_18218,N_17996,N_17785);
and U18219 (N_18219,N_17911,N_17904);
nand U18220 (N_18220,N_17925,N_17851);
and U18221 (N_18221,N_17968,N_17838);
nor U18222 (N_18222,N_17914,N_17907);
nor U18223 (N_18223,N_17957,N_17956);
nor U18224 (N_18224,N_17821,N_17942);
or U18225 (N_18225,N_17865,N_17949);
nor U18226 (N_18226,N_17996,N_17889);
xnor U18227 (N_18227,N_17946,N_17877);
nor U18228 (N_18228,N_17977,N_17932);
or U18229 (N_18229,N_17821,N_17892);
and U18230 (N_18230,N_17791,N_17769);
nand U18231 (N_18231,N_17832,N_17861);
or U18232 (N_18232,N_17996,N_17965);
and U18233 (N_18233,N_17906,N_17798);
xor U18234 (N_18234,N_17977,N_17763);
nor U18235 (N_18235,N_17862,N_17944);
or U18236 (N_18236,N_17920,N_17818);
nand U18237 (N_18237,N_17832,N_17916);
and U18238 (N_18238,N_17862,N_17933);
xor U18239 (N_18239,N_17816,N_17986);
xor U18240 (N_18240,N_17993,N_17885);
or U18241 (N_18241,N_17757,N_17831);
nor U18242 (N_18242,N_17823,N_17912);
and U18243 (N_18243,N_17835,N_17923);
or U18244 (N_18244,N_17852,N_17803);
and U18245 (N_18245,N_17823,N_17774);
nand U18246 (N_18246,N_17990,N_17988);
or U18247 (N_18247,N_17779,N_17764);
nand U18248 (N_18248,N_17819,N_17751);
nand U18249 (N_18249,N_17779,N_17979);
nand U18250 (N_18250,N_18186,N_18107);
xnor U18251 (N_18251,N_18109,N_18231);
nor U18252 (N_18252,N_18175,N_18026);
and U18253 (N_18253,N_18010,N_18183);
xnor U18254 (N_18254,N_18153,N_18158);
or U18255 (N_18255,N_18156,N_18233);
nor U18256 (N_18256,N_18170,N_18194);
nand U18257 (N_18257,N_18027,N_18116);
xor U18258 (N_18258,N_18097,N_18179);
xnor U18259 (N_18259,N_18047,N_18172);
or U18260 (N_18260,N_18148,N_18035);
nor U18261 (N_18261,N_18131,N_18248);
or U18262 (N_18262,N_18200,N_18155);
nor U18263 (N_18263,N_18143,N_18145);
and U18264 (N_18264,N_18236,N_18157);
or U18265 (N_18265,N_18210,N_18081);
and U18266 (N_18266,N_18220,N_18247);
and U18267 (N_18267,N_18168,N_18087);
nand U18268 (N_18268,N_18188,N_18065);
xnor U18269 (N_18269,N_18096,N_18075);
and U18270 (N_18270,N_18139,N_18038);
or U18271 (N_18271,N_18106,N_18084);
xor U18272 (N_18272,N_18062,N_18103);
xnor U18273 (N_18273,N_18083,N_18135);
nand U18274 (N_18274,N_18147,N_18070);
xor U18275 (N_18275,N_18076,N_18063);
xnor U18276 (N_18276,N_18078,N_18119);
nand U18277 (N_18277,N_18021,N_18074);
nand U18278 (N_18278,N_18060,N_18234);
xor U18279 (N_18279,N_18245,N_18144);
or U18280 (N_18280,N_18112,N_18137);
nor U18281 (N_18281,N_18014,N_18031);
xnor U18282 (N_18282,N_18192,N_18048);
or U18283 (N_18283,N_18006,N_18237);
and U18284 (N_18284,N_18044,N_18114);
xnor U18285 (N_18285,N_18053,N_18129);
nand U18286 (N_18286,N_18046,N_18187);
or U18287 (N_18287,N_18197,N_18196);
nand U18288 (N_18288,N_18141,N_18176);
or U18289 (N_18289,N_18163,N_18056);
nor U18290 (N_18290,N_18110,N_18189);
nor U18291 (N_18291,N_18102,N_18128);
and U18292 (N_18292,N_18177,N_18217);
nand U18293 (N_18293,N_18151,N_18016);
xor U18294 (N_18294,N_18167,N_18066);
nor U18295 (N_18295,N_18086,N_18132);
or U18296 (N_18296,N_18182,N_18199);
xor U18297 (N_18297,N_18240,N_18039);
or U18298 (N_18298,N_18222,N_18165);
and U18299 (N_18299,N_18160,N_18124);
xor U18300 (N_18300,N_18079,N_18218);
nand U18301 (N_18301,N_18029,N_18040);
nand U18302 (N_18302,N_18017,N_18052);
xnor U18303 (N_18303,N_18152,N_18204);
nor U18304 (N_18304,N_18050,N_18214);
or U18305 (N_18305,N_18012,N_18091);
and U18306 (N_18306,N_18211,N_18054);
or U18307 (N_18307,N_18082,N_18073);
xor U18308 (N_18308,N_18013,N_18174);
nor U18309 (N_18309,N_18125,N_18127);
nor U18310 (N_18310,N_18008,N_18232);
nand U18311 (N_18311,N_18191,N_18111);
xor U18312 (N_18312,N_18100,N_18215);
nand U18313 (N_18313,N_18241,N_18042);
nand U18314 (N_18314,N_18059,N_18193);
nand U18315 (N_18315,N_18166,N_18045);
or U18316 (N_18316,N_18181,N_18004);
xor U18317 (N_18317,N_18018,N_18180);
nor U18318 (N_18318,N_18037,N_18227);
and U18319 (N_18319,N_18134,N_18088);
or U18320 (N_18320,N_18022,N_18120);
nand U18321 (N_18321,N_18001,N_18229);
xnor U18322 (N_18322,N_18239,N_18077);
nand U18323 (N_18323,N_18136,N_18028);
and U18324 (N_18324,N_18205,N_18089);
and U18325 (N_18325,N_18000,N_18146);
and U18326 (N_18326,N_18202,N_18169);
xor U18327 (N_18327,N_18093,N_18178);
nand U18328 (N_18328,N_18138,N_18159);
or U18329 (N_18329,N_18171,N_18243);
nand U18330 (N_18330,N_18019,N_18108);
and U18331 (N_18331,N_18064,N_18095);
or U18332 (N_18332,N_18104,N_18190);
xor U18333 (N_18333,N_18249,N_18161);
nor U18334 (N_18334,N_18235,N_18150);
and U18335 (N_18335,N_18023,N_18126);
and U18336 (N_18336,N_18185,N_18219);
and U18337 (N_18337,N_18090,N_18041);
nor U18338 (N_18338,N_18009,N_18113);
and U18339 (N_18339,N_18094,N_18003);
xor U18340 (N_18340,N_18154,N_18133);
nor U18341 (N_18341,N_18226,N_18020);
and U18342 (N_18342,N_18142,N_18242);
xnor U18343 (N_18343,N_18195,N_18030);
or U18344 (N_18344,N_18072,N_18115);
nand U18345 (N_18345,N_18061,N_18213);
or U18346 (N_18346,N_18043,N_18080);
xor U18347 (N_18347,N_18173,N_18033);
xor U18348 (N_18348,N_18206,N_18025);
and U18349 (N_18349,N_18149,N_18230);
nand U18350 (N_18350,N_18055,N_18221);
and U18351 (N_18351,N_18099,N_18238);
xnor U18352 (N_18352,N_18224,N_18092);
xor U18353 (N_18353,N_18216,N_18067);
xor U18354 (N_18354,N_18032,N_18198);
and U18355 (N_18355,N_18069,N_18058);
nor U18356 (N_18356,N_18140,N_18209);
xor U18357 (N_18357,N_18002,N_18117);
and U18358 (N_18358,N_18228,N_18011);
nand U18359 (N_18359,N_18162,N_18071);
or U18360 (N_18360,N_18121,N_18015);
nand U18361 (N_18361,N_18007,N_18212);
xnor U18362 (N_18362,N_18034,N_18098);
nor U18363 (N_18363,N_18123,N_18223);
or U18364 (N_18364,N_18118,N_18036);
nor U18365 (N_18365,N_18049,N_18184);
nor U18366 (N_18366,N_18207,N_18005);
nand U18367 (N_18367,N_18122,N_18024);
nor U18368 (N_18368,N_18203,N_18105);
nor U18369 (N_18369,N_18068,N_18051);
xor U18370 (N_18370,N_18201,N_18057);
nand U18371 (N_18371,N_18130,N_18244);
and U18372 (N_18372,N_18164,N_18085);
and U18373 (N_18373,N_18101,N_18225);
nor U18374 (N_18374,N_18208,N_18246);
or U18375 (N_18375,N_18220,N_18227);
nor U18376 (N_18376,N_18220,N_18143);
xor U18377 (N_18377,N_18035,N_18088);
and U18378 (N_18378,N_18148,N_18143);
or U18379 (N_18379,N_18180,N_18164);
nor U18380 (N_18380,N_18105,N_18102);
or U18381 (N_18381,N_18189,N_18180);
nor U18382 (N_18382,N_18167,N_18111);
nand U18383 (N_18383,N_18142,N_18126);
xnor U18384 (N_18384,N_18184,N_18004);
nand U18385 (N_18385,N_18140,N_18000);
or U18386 (N_18386,N_18126,N_18039);
or U18387 (N_18387,N_18000,N_18185);
xnor U18388 (N_18388,N_18143,N_18200);
and U18389 (N_18389,N_18127,N_18038);
nand U18390 (N_18390,N_18117,N_18162);
nand U18391 (N_18391,N_18166,N_18047);
or U18392 (N_18392,N_18023,N_18108);
nor U18393 (N_18393,N_18030,N_18024);
xnor U18394 (N_18394,N_18105,N_18154);
xnor U18395 (N_18395,N_18134,N_18209);
xor U18396 (N_18396,N_18166,N_18115);
or U18397 (N_18397,N_18127,N_18235);
nand U18398 (N_18398,N_18131,N_18194);
nand U18399 (N_18399,N_18214,N_18213);
nor U18400 (N_18400,N_18131,N_18146);
xnor U18401 (N_18401,N_18201,N_18000);
nor U18402 (N_18402,N_18172,N_18162);
nor U18403 (N_18403,N_18199,N_18101);
nor U18404 (N_18404,N_18246,N_18059);
xor U18405 (N_18405,N_18009,N_18102);
or U18406 (N_18406,N_18012,N_18174);
and U18407 (N_18407,N_18035,N_18078);
xor U18408 (N_18408,N_18086,N_18026);
nand U18409 (N_18409,N_18020,N_18239);
nor U18410 (N_18410,N_18089,N_18118);
xnor U18411 (N_18411,N_18174,N_18230);
and U18412 (N_18412,N_18077,N_18187);
nor U18413 (N_18413,N_18099,N_18246);
and U18414 (N_18414,N_18172,N_18035);
nand U18415 (N_18415,N_18027,N_18232);
and U18416 (N_18416,N_18158,N_18055);
xor U18417 (N_18417,N_18099,N_18104);
and U18418 (N_18418,N_18226,N_18095);
or U18419 (N_18419,N_18182,N_18083);
nand U18420 (N_18420,N_18172,N_18214);
xnor U18421 (N_18421,N_18187,N_18065);
or U18422 (N_18422,N_18020,N_18096);
and U18423 (N_18423,N_18129,N_18234);
xor U18424 (N_18424,N_18004,N_18081);
nor U18425 (N_18425,N_18020,N_18209);
nand U18426 (N_18426,N_18136,N_18245);
nor U18427 (N_18427,N_18149,N_18192);
xnor U18428 (N_18428,N_18153,N_18147);
xnor U18429 (N_18429,N_18046,N_18165);
xnor U18430 (N_18430,N_18177,N_18229);
nor U18431 (N_18431,N_18153,N_18063);
and U18432 (N_18432,N_18215,N_18213);
or U18433 (N_18433,N_18231,N_18199);
or U18434 (N_18434,N_18188,N_18224);
or U18435 (N_18435,N_18099,N_18229);
and U18436 (N_18436,N_18161,N_18019);
xnor U18437 (N_18437,N_18194,N_18173);
and U18438 (N_18438,N_18089,N_18160);
and U18439 (N_18439,N_18212,N_18202);
nand U18440 (N_18440,N_18012,N_18141);
or U18441 (N_18441,N_18139,N_18178);
nor U18442 (N_18442,N_18176,N_18001);
and U18443 (N_18443,N_18172,N_18245);
nand U18444 (N_18444,N_18243,N_18041);
nand U18445 (N_18445,N_18069,N_18087);
xor U18446 (N_18446,N_18109,N_18129);
xnor U18447 (N_18447,N_18006,N_18158);
and U18448 (N_18448,N_18180,N_18127);
or U18449 (N_18449,N_18231,N_18030);
or U18450 (N_18450,N_18054,N_18055);
nand U18451 (N_18451,N_18010,N_18240);
or U18452 (N_18452,N_18187,N_18058);
or U18453 (N_18453,N_18169,N_18035);
or U18454 (N_18454,N_18105,N_18075);
nand U18455 (N_18455,N_18202,N_18130);
or U18456 (N_18456,N_18214,N_18099);
xor U18457 (N_18457,N_18165,N_18209);
nand U18458 (N_18458,N_18123,N_18010);
nor U18459 (N_18459,N_18235,N_18218);
nor U18460 (N_18460,N_18045,N_18235);
and U18461 (N_18461,N_18066,N_18109);
or U18462 (N_18462,N_18167,N_18204);
and U18463 (N_18463,N_18175,N_18205);
and U18464 (N_18464,N_18150,N_18097);
and U18465 (N_18465,N_18233,N_18196);
nand U18466 (N_18466,N_18119,N_18083);
nand U18467 (N_18467,N_18232,N_18247);
nor U18468 (N_18468,N_18148,N_18185);
and U18469 (N_18469,N_18148,N_18081);
nand U18470 (N_18470,N_18107,N_18025);
or U18471 (N_18471,N_18000,N_18199);
xnor U18472 (N_18472,N_18080,N_18050);
nand U18473 (N_18473,N_18047,N_18220);
xor U18474 (N_18474,N_18104,N_18071);
and U18475 (N_18475,N_18208,N_18063);
nand U18476 (N_18476,N_18213,N_18100);
nor U18477 (N_18477,N_18242,N_18092);
nor U18478 (N_18478,N_18084,N_18026);
nor U18479 (N_18479,N_18172,N_18163);
nand U18480 (N_18480,N_18242,N_18012);
nand U18481 (N_18481,N_18216,N_18218);
nand U18482 (N_18482,N_18188,N_18070);
nand U18483 (N_18483,N_18199,N_18167);
nor U18484 (N_18484,N_18230,N_18165);
nand U18485 (N_18485,N_18229,N_18166);
or U18486 (N_18486,N_18180,N_18212);
or U18487 (N_18487,N_18145,N_18190);
xor U18488 (N_18488,N_18230,N_18012);
nor U18489 (N_18489,N_18165,N_18126);
nor U18490 (N_18490,N_18133,N_18236);
and U18491 (N_18491,N_18229,N_18184);
or U18492 (N_18492,N_18153,N_18117);
or U18493 (N_18493,N_18070,N_18031);
and U18494 (N_18494,N_18223,N_18015);
nand U18495 (N_18495,N_18077,N_18132);
xor U18496 (N_18496,N_18140,N_18203);
nand U18497 (N_18497,N_18011,N_18136);
xnor U18498 (N_18498,N_18032,N_18154);
and U18499 (N_18499,N_18090,N_18218);
or U18500 (N_18500,N_18437,N_18474);
and U18501 (N_18501,N_18341,N_18354);
or U18502 (N_18502,N_18498,N_18471);
nand U18503 (N_18503,N_18459,N_18297);
xnor U18504 (N_18504,N_18385,N_18335);
nor U18505 (N_18505,N_18321,N_18311);
xor U18506 (N_18506,N_18304,N_18334);
or U18507 (N_18507,N_18336,N_18340);
nand U18508 (N_18508,N_18472,N_18346);
or U18509 (N_18509,N_18475,N_18374);
or U18510 (N_18510,N_18382,N_18309);
nand U18511 (N_18511,N_18455,N_18273);
and U18512 (N_18512,N_18404,N_18255);
nand U18513 (N_18513,N_18417,N_18323);
nand U18514 (N_18514,N_18351,N_18337);
and U18515 (N_18515,N_18443,N_18305);
nor U18516 (N_18516,N_18313,N_18258);
nand U18517 (N_18517,N_18429,N_18369);
nand U18518 (N_18518,N_18262,N_18410);
nor U18519 (N_18519,N_18444,N_18407);
and U18520 (N_18520,N_18491,N_18328);
nor U18521 (N_18521,N_18329,N_18485);
nor U18522 (N_18522,N_18431,N_18421);
and U18523 (N_18523,N_18257,N_18386);
xnor U18524 (N_18524,N_18299,N_18473);
nor U18525 (N_18525,N_18468,N_18364);
nor U18526 (N_18526,N_18449,N_18342);
and U18527 (N_18527,N_18415,N_18390);
nor U18528 (N_18528,N_18486,N_18463);
nand U18529 (N_18529,N_18401,N_18447);
or U18530 (N_18530,N_18457,N_18344);
xor U18531 (N_18531,N_18379,N_18306);
nor U18532 (N_18532,N_18488,N_18363);
nor U18533 (N_18533,N_18484,N_18263);
xnor U18534 (N_18534,N_18458,N_18439);
xor U18535 (N_18535,N_18413,N_18419);
nand U18536 (N_18536,N_18256,N_18274);
nor U18537 (N_18537,N_18435,N_18389);
or U18538 (N_18538,N_18295,N_18312);
nor U18539 (N_18539,N_18322,N_18367);
nor U18540 (N_18540,N_18302,N_18405);
nor U18541 (N_18541,N_18264,N_18418);
xnor U18542 (N_18542,N_18261,N_18427);
and U18543 (N_18543,N_18403,N_18260);
and U18544 (N_18544,N_18284,N_18350);
or U18545 (N_18545,N_18453,N_18448);
or U18546 (N_18546,N_18310,N_18398);
nor U18547 (N_18547,N_18432,N_18366);
and U18548 (N_18548,N_18440,N_18275);
and U18549 (N_18549,N_18450,N_18276);
nand U18550 (N_18550,N_18481,N_18317);
nand U18551 (N_18551,N_18378,N_18361);
and U18552 (N_18552,N_18283,N_18412);
nor U18553 (N_18553,N_18308,N_18339);
or U18554 (N_18554,N_18254,N_18406);
and U18555 (N_18555,N_18315,N_18290);
nand U18556 (N_18556,N_18288,N_18372);
and U18557 (N_18557,N_18371,N_18461);
xor U18558 (N_18558,N_18436,N_18469);
and U18559 (N_18559,N_18253,N_18482);
nor U18560 (N_18560,N_18259,N_18286);
nand U18561 (N_18561,N_18345,N_18483);
or U18562 (N_18562,N_18392,N_18296);
nand U18563 (N_18563,N_18338,N_18320);
nand U18564 (N_18564,N_18269,N_18442);
nand U18565 (N_18565,N_18266,N_18285);
nor U18566 (N_18566,N_18353,N_18377);
and U18567 (N_18567,N_18362,N_18307);
xnor U18568 (N_18568,N_18327,N_18375);
nand U18569 (N_18569,N_18497,N_18496);
or U18570 (N_18570,N_18303,N_18325);
nand U18571 (N_18571,N_18278,N_18438);
nor U18572 (N_18572,N_18479,N_18318);
nor U18573 (N_18573,N_18426,N_18281);
and U18574 (N_18574,N_18470,N_18466);
xnor U18575 (N_18575,N_18424,N_18454);
nand U18576 (N_18576,N_18411,N_18282);
xor U18577 (N_18577,N_18316,N_18359);
xor U18578 (N_18578,N_18330,N_18465);
and U18579 (N_18579,N_18476,N_18358);
and U18580 (N_18580,N_18343,N_18477);
nor U18581 (N_18581,N_18271,N_18287);
nor U18582 (N_18582,N_18399,N_18393);
nand U18583 (N_18583,N_18445,N_18396);
nor U18584 (N_18584,N_18409,N_18387);
or U18585 (N_18585,N_18480,N_18467);
nor U18586 (N_18586,N_18397,N_18490);
and U18587 (N_18587,N_18289,N_18433);
nor U18588 (N_18588,N_18402,N_18324);
nor U18589 (N_18589,N_18265,N_18425);
or U18590 (N_18590,N_18270,N_18478);
xor U18591 (N_18591,N_18456,N_18331);
nand U18592 (N_18592,N_18384,N_18391);
and U18593 (N_18593,N_18422,N_18388);
nor U18594 (N_18594,N_18492,N_18298);
nor U18595 (N_18595,N_18356,N_18268);
nor U18596 (N_18596,N_18280,N_18464);
and U18597 (N_18597,N_18383,N_18332);
xor U18598 (N_18598,N_18370,N_18250);
nand U18599 (N_18599,N_18400,N_18499);
xor U18600 (N_18600,N_18416,N_18376);
and U18601 (N_18601,N_18368,N_18460);
and U18602 (N_18602,N_18349,N_18495);
and U18603 (N_18603,N_18446,N_18381);
xor U18604 (N_18604,N_18423,N_18326);
nor U18605 (N_18605,N_18394,N_18252);
nand U18606 (N_18606,N_18452,N_18493);
nor U18607 (N_18607,N_18360,N_18319);
nor U18608 (N_18608,N_18357,N_18434);
xor U18609 (N_18609,N_18277,N_18489);
nor U18610 (N_18610,N_18314,N_18279);
xnor U18611 (N_18611,N_18365,N_18352);
nor U18612 (N_18612,N_18428,N_18380);
or U18613 (N_18613,N_18301,N_18441);
or U18614 (N_18614,N_18251,N_18462);
and U18615 (N_18615,N_18294,N_18430);
and U18616 (N_18616,N_18272,N_18451);
nor U18617 (N_18617,N_18291,N_18420);
nand U18618 (N_18618,N_18348,N_18347);
nand U18619 (N_18619,N_18355,N_18373);
and U18620 (N_18620,N_18414,N_18333);
nand U18621 (N_18621,N_18487,N_18293);
nand U18622 (N_18622,N_18408,N_18292);
or U18623 (N_18623,N_18300,N_18395);
nand U18624 (N_18624,N_18267,N_18494);
or U18625 (N_18625,N_18392,N_18391);
nor U18626 (N_18626,N_18460,N_18292);
xnor U18627 (N_18627,N_18370,N_18412);
xnor U18628 (N_18628,N_18342,N_18287);
and U18629 (N_18629,N_18301,N_18470);
nor U18630 (N_18630,N_18484,N_18353);
xnor U18631 (N_18631,N_18401,N_18436);
or U18632 (N_18632,N_18250,N_18316);
and U18633 (N_18633,N_18372,N_18337);
nand U18634 (N_18634,N_18407,N_18283);
nand U18635 (N_18635,N_18344,N_18419);
or U18636 (N_18636,N_18471,N_18327);
and U18637 (N_18637,N_18281,N_18326);
or U18638 (N_18638,N_18289,N_18348);
and U18639 (N_18639,N_18259,N_18266);
nand U18640 (N_18640,N_18473,N_18324);
nand U18641 (N_18641,N_18421,N_18483);
and U18642 (N_18642,N_18369,N_18475);
nand U18643 (N_18643,N_18328,N_18254);
and U18644 (N_18644,N_18269,N_18490);
nand U18645 (N_18645,N_18345,N_18499);
and U18646 (N_18646,N_18427,N_18331);
nor U18647 (N_18647,N_18407,N_18412);
nand U18648 (N_18648,N_18444,N_18411);
nand U18649 (N_18649,N_18339,N_18492);
and U18650 (N_18650,N_18289,N_18397);
xor U18651 (N_18651,N_18257,N_18418);
and U18652 (N_18652,N_18332,N_18311);
or U18653 (N_18653,N_18295,N_18406);
nor U18654 (N_18654,N_18342,N_18469);
xor U18655 (N_18655,N_18369,N_18314);
or U18656 (N_18656,N_18363,N_18293);
nand U18657 (N_18657,N_18330,N_18440);
nand U18658 (N_18658,N_18320,N_18411);
nor U18659 (N_18659,N_18443,N_18273);
nand U18660 (N_18660,N_18260,N_18289);
or U18661 (N_18661,N_18493,N_18389);
xnor U18662 (N_18662,N_18495,N_18455);
nand U18663 (N_18663,N_18425,N_18356);
or U18664 (N_18664,N_18266,N_18292);
xnor U18665 (N_18665,N_18324,N_18416);
xnor U18666 (N_18666,N_18347,N_18442);
or U18667 (N_18667,N_18327,N_18281);
or U18668 (N_18668,N_18470,N_18345);
xor U18669 (N_18669,N_18364,N_18347);
nor U18670 (N_18670,N_18390,N_18342);
and U18671 (N_18671,N_18366,N_18456);
and U18672 (N_18672,N_18264,N_18376);
nor U18673 (N_18673,N_18351,N_18359);
and U18674 (N_18674,N_18368,N_18296);
nor U18675 (N_18675,N_18347,N_18252);
or U18676 (N_18676,N_18490,N_18454);
nor U18677 (N_18677,N_18416,N_18435);
nor U18678 (N_18678,N_18294,N_18267);
or U18679 (N_18679,N_18293,N_18421);
nand U18680 (N_18680,N_18329,N_18402);
xor U18681 (N_18681,N_18375,N_18381);
nand U18682 (N_18682,N_18474,N_18305);
nand U18683 (N_18683,N_18448,N_18334);
and U18684 (N_18684,N_18462,N_18299);
xor U18685 (N_18685,N_18322,N_18299);
or U18686 (N_18686,N_18398,N_18325);
and U18687 (N_18687,N_18276,N_18302);
nor U18688 (N_18688,N_18333,N_18270);
nor U18689 (N_18689,N_18498,N_18443);
and U18690 (N_18690,N_18458,N_18349);
and U18691 (N_18691,N_18472,N_18251);
and U18692 (N_18692,N_18260,N_18339);
nand U18693 (N_18693,N_18449,N_18396);
nand U18694 (N_18694,N_18324,N_18453);
and U18695 (N_18695,N_18466,N_18371);
xnor U18696 (N_18696,N_18447,N_18452);
nand U18697 (N_18697,N_18461,N_18266);
nor U18698 (N_18698,N_18291,N_18295);
nand U18699 (N_18699,N_18306,N_18375);
xor U18700 (N_18700,N_18273,N_18396);
and U18701 (N_18701,N_18493,N_18351);
nand U18702 (N_18702,N_18495,N_18385);
and U18703 (N_18703,N_18307,N_18463);
nor U18704 (N_18704,N_18467,N_18499);
nor U18705 (N_18705,N_18328,N_18375);
nand U18706 (N_18706,N_18289,N_18496);
nand U18707 (N_18707,N_18444,N_18418);
nand U18708 (N_18708,N_18343,N_18460);
nor U18709 (N_18709,N_18261,N_18437);
and U18710 (N_18710,N_18274,N_18357);
xnor U18711 (N_18711,N_18373,N_18311);
and U18712 (N_18712,N_18492,N_18290);
nor U18713 (N_18713,N_18267,N_18257);
xor U18714 (N_18714,N_18446,N_18343);
or U18715 (N_18715,N_18294,N_18397);
xor U18716 (N_18716,N_18411,N_18416);
nand U18717 (N_18717,N_18476,N_18351);
nor U18718 (N_18718,N_18309,N_18365);
or U18719 (N_18719,N_18485,N_18420);
nor U18720 (N_18720,N_18431,N_18354);
nor U18721 (N_18721,N_18348,N_18337);
nor U18722 (N_18722,N_18288,N_18370);
nor U18723 (N_18723,N_18314,N_18313);
xnor U18724 (N_18724,N_18387,N_18462);
and U18725 (N_18725,N_18462,N_18327);
or U18726 (N_18726,N_18313,N_18307);
xnor U18727 (N_18727,N_18491,N_18269);
and U18728 (N_18728,N_18279,N_18276);
and U18729 (N_18729,N_18411,N_18429);
nand U18730 (N_18730,N_18312,N_18336);
and U18731 (N_18731,N_18401,N_18365);
or U18732 (N_18732,N_18462,N_18293);
nor U18733 (N_18733,N_18304,N_18356);
nand U18734 (N_18734,N_18351,N_18392);
xnor U18735 (N_18735,N_18345,N_18422);
and U18736 (N_18736,N_18492,N_18320);
nand U18737 (N_18737,N_18278,N_18480);
or U18738 (N_18738,N_18348,N_18293);
nor U18739 (N_18739,N_18457,N_18453);
and U18740 (N_18740,N_18290,N_18408);
or U18741 (N_18741,N_18396,N_18417);
or U18742 (N_18742,N_18291,N_18303);
and U18743 (N_18743,N_18322,N_18467);
nor U18744 (N_18744,N_18261,N_18252);
nand U18745 (N_18745,N_18365,N_18287);
and U18746 (N_18746,N_18384,N_18443);
or U18747 (N_18747,N_18277,N_18333);
and U18748 (N_18748,N_18365,N_18423);
xnor U18749 (N_18749,N_18441,N_18287);
xnor U18750 (N_18750,N_18721,N_18525);
nand U18751 (N_18751,N_18738,N_18555);
and U18752 (N_18752,N_18746,N_18697);
nand U18753 (N_18753,N_18609,N_18704);
nor U18754 (N_18754,N_18570,N_18518);
xnor U18755 (N_18755,N_18584,N_18623);
or U18756 (N_18756,N_18695,N_18568);
xor U18757 (N_18757,N_18578,N_18514);
nor U18758 (N_18758,N_18612,N_18732);
nor U18759 (N_18759,N_18714,N_18660);
nor U18760 (N_18760,N_18506,N_18505);
nor U18761 (N_18761,N_18583,N_18647);
xnor U18762 (N_18762,N_18736,N_18724);
and U18763 (N_18763,N_18743,N_18662);
nand U18764 (N_18764,N_18577,N_18579);
and U18765 (N_18765,N_18571,N_18679);
xnor U18766 (N_18766,N_18676,N_18620);
nand U18767 (N_18767,N_18547,N_18566);
nor U18768 (N_18768,N_18698,N_18646);
or U18769 (N_18769,N_18531,N_18587);
or U18770 (N_18770,N_18546,N_18633);
nand U18771 (N_18771,N_18558,N_18628);
nor U18772 (N_18772,N_18708,N_18635);
xnor U18773 (N_18773,N_18630,N_18717);
nand U18774 (N_18774,N_18601,N_18634);
nand U18775 (N_18775,N_18520,N_18552);
xor U18776 (N_18776,N_18618,N_18632);
and U18777 (N_18777,N_18699,N_18530);
nand U18778 (N_18778,N_18709,N_18517);
nand U18779 (N_18779,N_18688,N_18681);
or U18780 (N_18780,N_18575,N_18561);
nor U18781 (N_18781,N_18533,N_18507);
nor U18782 (N_18782,N_18564,N_18509);
and U18783 (N_18783,N_18692,N_18508);
nand U18784 (N_18784,N_18621,N_18730);
nor U18785 (N_18785,N_18614,N_18742);
and U18786 (N_18786,N_18576,N_18607);
nor U18787 (N_18787,N_18745,N_18683);
xnor U18788 (N_18788,N_18636,N_18663);
xor U18789 (N_18789,N_18696,N_18669);
nor U18790 (N_18790,N_18710,N_18656);
or U18791 (N_18791,N_18522,N_18668);
and U18792 (N_18792,N_18666,N_18739);
and U18793 (N_18793,N_18649,N_18574);
and U18794 (N_18794,N_18526,N_18673);
and U18795 (N_18795,N_18733,N_18741);
nor U18796 (N_18796,N_18549,N_18554);
and U18797 (N_18797,N_18648,N_18731);
nor U18798 (N_18798,N_18585,N_18503);
nand U18799 (N_18799,N_18643,N_18582);
nand U18800 (N_18800,N_18586,N_18567);
and U18801 (N_18801,N_18653,N_18705);
xnor U18802 (N_18802,N_18548,N_18703);
nor U18803 (N_18803,N_18678,N_18545);
and U18804 (N_18804,N_18672,N_18674);
xor U18805 (N_18805,N_18563,N_18611);
nor U18806 (N_18806,N_18625,N_18686);
xnor U18807 (N_18807,N_18535,N_18543);
nand U18808 (N_18808,N_18675,N_18627);
nor U18809 (N_18809,N_18671,N_18670);
nor U18810 (N_18810,N_18734,N_18685);
or U18811 (N_18811,N_18718,N_18640);
nand U18812 (N_18812,N_18713,N_18622);
xor U18813 (N_18813,N_18581,N_18510);
and U18814 (N_18814,N_18631,N_18608);
or U18815 (N_18815,N_18598,N_18701);
xor U18816 (N_18816,N_18613,N_18599);
nand U18817 (N_18817,N_18544,N_18716);
nor U18818 (N_18818,N_18638,N_18610);
and U18819 (N_18819,N_18565,N_18593);
or U18820 (N_18820,N_18528,N_18682);
or U18821 (N_18821,N_18605,N_18641);
and U18822 (N_18822,N_18560,N_18600);
or U18823 (N_18823,N_18728,N_18619);
or U18824 (N_18824,N_18589,N_18502);
nor U18825 (N_18825,N_18711,N_18616);
nand U18826 (N_18826,N_18521,N_18665);
xor U18827 (N_18827,N_18513,N_18726);
nand U18828 (N_18828,N_18748,N_18542);
xnor U18829 (N_18829,N_18689,N_18624);
nor U18830 (N_18830,N_18725,N_18693);
and U18831 (N_18831,N_18715,N_18597);
or U18832 (N_18832,N_18596,N_18556);
nor U18833 (N_18833,N_18626,N_18747);
nor U18834 (N_18834,N_18532,N_18720);
nand U18835 (N_18835,N_18537,N_18500);
or U18836 (N_18836,N_18642,N_18690);
nand U18837 (N_18837,N_18562,N_18534);
or U18838 (N_18838,N_18588,N_18539);
and U18839 (N_18839,N_18538,N_18604);
or U18840 (N_18840,N_18603,N_18652);
nand U18841 (N_18841,N_18559,N_18645);
xnor U18842 (N_18842,N_18637,N_18557);
and U18843 (N_18843,N_18524,N_18606);
xor U18844 (N_18844,N_18515,N_18684);
nor U18845 (N_18845,N_18615,N_18523);
and U18846 (N_18846,N_18664,N_18536);
nand U18847 (N_18847,N_18654,N_18629);
or U18848 (N_18848,N_18694,N_18553);
nand U18849 (N_18849,N_18617,N_18591);
and U18850 (N_18850,N_18512,N_18529);
and U18851 (N_18851,N_18740,N_18650);
xnor U18852 (N_18852,N_18592,N_18651);
nand U18853 (N_18853,N_18655,N_18722);
nand U18854 (N_18854,N_18659,N_18661);
xor U18855 (N_18855,N_18712,N_18737);
and U18856 (N_18856,N_18519,N_18719);
or U18857 (N_18857,N_18550,N_18516);
and U18858 (N_18858,N_18573,N_18707);
or U18859 (N_18859,N_18658,N_18691);
or U18860 (N_18860,N_18723,N_18749);
nor U18861 (N_18861,N_18572,N_18677);
or U18862 (N_18862,N_18580,N_18501);
nor U18863 (N_18863,N_18729,N_18595);
and U18864 (N_18864,N_18702,N_18680);
or U18865 (N_18865,N_18569,N_18744);
nand U18866 (N_18866,N_18541,N_18639);
and U18867 (N_18867,N_18527,N_18727);
xor U18868 (N_18868,N_18735,N_18551);
nor U18869 (N_18869,N_18644,N_18590);
or U18870 (N_18870,N_18700,N_18594);
nand U18871 (N_18871,N_18667,N_18504);
nand U18872 (N_18872,N_18706,N_18657);
or U18873 (N_18873,N_18602,N_18687);
xnor U18874 (N_18874,N_18540,N_18511);
and U18875 (N_18875,N_18662,N_18727);
nand U18876 (N_18876,N_18723,N_18715);
nor U18877 (N_18877,N_18556,N_18680);
or U18878 (N_18878,N_18617,N_18732);
nand U18879 (N_18879,N_18614,N_18637);
or U18880 (N_18880,N_18645,N_18582);
nor U18881 (N_18881,N_18644,N_18616);
or U18882 (N_18882,N_18645,N_18718);
or U18883 (N_18883,N_18636,N_18640);
nand U18884 (N_18884,N_18730,N_18725);
or U18885 (N_18885,N_18502,N_18526);
nor U18886 (N_18886,N_18581,N_18508);
nand U18887 (N_18887,N_18564,N_18569);
and U18888 (N_18888,N_18725,N_18614);
nand U18889 (N_18889,N_18711,N_18523);
or U18890 (N_18890,N_18742,N_18564);
or U18891 (N_18891,N_18538,N_18725);
nand U18892 (N_18892,N_18578,N_18635);
and U18893 (N_18893,N_18734,N_18636);
nor U18894 (N_18894,N_18509,N_18726);
nor U18895 (N_18895,N_18587,N_18666);
or U18896 (N_18896,N_18688,N_18704);
nand U18897 (N_18897,N_18603,N_18646);
nor U18898 (N_18898,N_18637,N_18572);
or U18899 (N_18899,N_18545,N_18700);
nand U18900 (N_18900,N_18620,N_18617);
or U18901 (N_18901,N_18722,N_18557);
nor U18902 (N_18902,N_18705,N_18646);
nand U18903 (N_18903,N_18605,N_18705);
and U18904 (N_18904,N_18555,N_18649);
xor U18905 (N_18905,N_18595,N_18722);
and U18906 (N_18906,N_18621,N_18553);
or U18907 (N_18907,N_18528,N_18571);
or U18908 (N_18908,N_18622,N_18610);
xnor U18909 (N_18909,N_18675,N_18516);
or U18910 (N_18910,N_18679,N_18504);
and U18911 (N_18911,N_18630,N_18606);
xor U18912 (N_18912,N_18626,N_18508);
nand U18913 (N_18913,N_18520,N_18511);
xor U18914 (N_18914,N_18619,N_18722);
nor U18915 (N_18915,N_18581,N_18691);
nor U18916 (N_18916,N_18583,N_18602);
and U18917 (N_18917,N_18683,N_18638);
xnor U18918 (N_18918,N_18667,N_18658);
nand U18919 (N_18919,N_18617,N_18505);
nand U18920 (N_18920,N_18669,N_18603);
and U18921 (N_18921,N_18527,N_18575);
nor U18922 (N_18922,N_18579,N_18715);
nor U18923 (N_18923,N_18627,N_18600);
nand U18924 (N_18924,N_18683,N_18525);
nand U18925 (N_18925,N_18731,N_18612);
xor U18926 (N_18926,N_18516,N_18582);
nor U18927 (N_18927,N_18539,N_18582);
nand U18928 (N_18928,N_18587,N_18603);
xnor U18929 (N_18929,N_18618,N_18658);
nor U18930 (N_18930,N_18710,N_18719);
nand U18931 (N_18931,N_18568,N_18638);
or U18932 (N_18932,N_18709,N_18749);
nand U18933 (N_18933,N_18613,N_18528);
or U18934 (N_18934,N_18677,N_18500);
nand U18935 (N_18935,N_18551,N_18710);
nor U18936 (N_18936,N_18542,N_18576);
nand U18937 (N_18937,N_18692,N_18730);
nor U18938 (N_18938,N_18633,N_18558);
nand U18939 (N_18939,N_18544,N_18541);
nor U18940 (N_18940,N_18542,N_18591);
or U18941 (N_18941,N_18574,N_18664);
or U18942 (N_18942,N_18728,N_18679);
nand U18943 (N_18943,N_18628,N_18645);
and U18944 (N_18944,N_18548,N_18735);
nand U18945 (N_18945,N_18662,N_18657);
or U18946 (N_18946,N_18610,N_18525);
nor U18947 (N_18947,N_18660,N_18608);
xor U18948 (N_18948,N_18540,N_18635);
nor U18949 (N_18949,N_18736,N_18669);
xor U18950 (N_18950,N_18549,N_18665);
or U18951 (N_18951,N_18703,N_18513);
xnor U18952 (N_18952,N_18529,N_18535);
or U18953 (N_18953,N_18741,N_18693);
or U18954 (N_18954,N_18693,N_18556);
nand U18955 (N_18955,N_18703,N_18708);
or U18956 (N_18956,N_18749,N_18686);
nand U18957 (N_18957,N_18626,N_18737);
or U18958 (N_18958,N_18737,N_18533);
nand U18959 (N_18959,N_18712,N_18625);
and U18960 (N_18960,N_18516,N_18590);
nand U18961 (N_18961,N_18536,N_18543);
or U18962 (N_18962,N_18636,N_18521);
xnor U18963 (N_18963,N_18533,N_18595);
xor U18964 (N_18964,N_18681,N_18732);
nor U18965 (N_18965,N_18567,N_18704);
or U18966 (N_18966,N_18692,N_18698);
nor U18967 (N_18967,N_18609,N_18536);
or U18968 (N_18968,N_18690,N_18512);
xnor U18969 (N_18969,N_18737,N_18544);
nand U18970 (N_18970,N_18748,N_18580);
nand U18971 (N_18971,N_18614,N_18638);
and U18972 (N_18972,N_18721,N_18565);
and U18973 (N_18973,N_18706,N_18583);
xor U18974 (N_18974,N_18655,N_18549);
nor U18975 (N_18975,N_18541,N_18691);
and U18976 (N_18976,N_18667,N_18599);
nor U18977 (N_18977,N_18521,N_18610);
nor U18978 (N_18978,N_18733,N_18570);
xnor U18979 (N_18979,N_18528,N_18646);
xnor U18980 (N_18980,N_18713,N_18711);
xnor U18981 (N_18981,N_18721,N_18665);
or U18982 (N_18982,N_18736,N_18610);
or U18983 (N_18983,N_18584,N_18744);
and U18984 (N_18984,N_18501,N_18619);
xnor U18985 (N_18985,N_18626,N_18586);
and U18986 (N_18986,N_18600,N_18721);
or U18987 (N_18987,N_18516,N_18527);
nor U18988 (N_18988,N_18730,N_18503);
nor U18989 (N_18989,N_18512,N_18540);
xor U18990 (N_18990,N_18656,N_18723);
nand U18991 (N_18991,N_18552,N_18536);
or U18992 (N_18992,N_18686,N_18622);
nand U18993 (N_18993,N_18525,N_18591);
nand U18994 (N_18994,N_18716,N_18606);
or U18995 (N_18995,N_18643,N_18651);
and U18996 (N_18996,N_18625,N_18684);
nand U18997 (N_18997,N_18542,N_18655);
xnor U18998 (N_18998,N_18659,N_18592);
xnor U18999 (N_18999,N_18564,N_18713);
nor U19000 (N_19000,N_18758,N_18876);
nor U19001 (N_19001,N_18843,N_18946);
nor U19002 (N_19002,N_18817,N_18846);
nor U19003 (N_19003,N_18844,N_18850);
and U19004 (N_19004,N_18807,N_18877);
nor U19005 (N_19005,N_18774,N_18851);
nor U19006 (N_19006,N_18939,N_18857);
xnor U19007 (N_19007,N_18802,N_18966);
xnor U19008 (N_19008,N_18945,N_18950);
xnor U19009 (N_19009,N_18932,N_18911);
nor U19010 (N_19010,N_18806,N_18975);
nor U19011 (N_19011,N_18860,N_18835);
xor U19012 (N_19012,N_18959,N_18952);
nand U19013 (N_19013,N_18994,N_18971);
xnor U19014 (N_19014,N_18997,N_18920);
nand U19015 (N_19015,N_18987,N_18925);
nand U19016 (N_19016,N_18985,N_18875);
and U19017 (N_19017,N_18951,N_18848);
nand U19018 (N_19018,N_18931,N_18820);
or U19019 (N_19019,N_18893,N_18965);
nand U19020 (N_19020,N_18963,N_18841);
or U19021 (N_19021,N_18888,N_18906);
or U19022 (N_19022,N_18919,N_18929);
nand U19023 (N_19023,N_18755,N_18881);
nor U19024 (N_19024,N_18898,N_18958);
xnor U19025 (N_19025,N_18792,N_18890);
or U19026 (N_19026,N_18883,N_18854);
and U19027 (N_19027,N_18934,N_18779);
and U19028 (N_19028,N_18790,N_18778);
xor U19029 (N_19029,N_18954,N_18927);
nand U19030 (N_19030,N_18940,N_18878);
nor U19031 (N_19031,N_18796,N_18885);
nor U19032 (N_19032,N_18900,N_18801);
xnor U19033 (N_19033,N_18957,N_18988);
and U19034 (N_19034,N_18765,N_18834);
xnor U19035 (N_19035,N_18791,N_18989);
and U19036 (N_19036,N_18836,N_18809);
nor U19037 (N_19037,N_18813,N_18889);
nor U19038 (N_19038,N_18808,N_18759);
nand U19039 (N_19039,N_18936,N_18770);
or U19040 (N_19040,N_18849,N_18899);
or U19041 (N_19041,N_18840,N_18903);
xor U19042 (N_19042,N_18897,N_18865);
and U19043 (N_19043,N_18795,N_18753);
nand U19044 (N_19044,N_18798,N_18956);
xor U19045 (N_19045,N_18980,N_18953);
and U19046 (N_19046,N_18861,N_18831);
and U19047 (N_19047,N_18884,N_18803);
and U19048 (N_19048,N_18826,N_18923);
and U19049 (N_19049,N_18999,N_18754);
and U19050 (N_19050,N_18990,N_18855);
or U19051 (N_19051,N_18852,N_18823);
nor U19052 (N_19052,N_18913,N_18891);
xor U19053 (N_19053,N_18799,N_18873);
xor U19054 (N_19054,N_18812,N_18926);
xnor U19055 (N_19055,N_18894,N_18805);
xor U19056 (N_19056,N_18974,N_18967);
and U19057 (N_19057,N_18781,N_18783);
xnor U19058 (N_19058,N_18948,N_18794);
nor U19059 (N_19059,N_18751,N_18979);
or U19060 (N_19060,N_18968,N_18986);
and U19061 (N_19061,N_18976,N_18858);
xnor U19062 (N_19062,N_18752,N_18845);
nor U19063 (N_19063,N_18814,N_18775);
or U19064 (N_19064,N_18864,N_18872);
and U19065 (N_19065,N_18962,N_18978);
and U19066 (N_19066,N_18960,N_18905);
nand U19067 (N_19067,N_18941,N_18930);
or U19068 (N_19068,N_18830,N_18868);
nor U19069 (N_19069,N_18970,N_18879);
and U19070 (N_19070,N_18943,N_18837);
nand U19071 (N_19071,N_18800,N_18769);
nand U19072 (N_19072,N_18995,N_18811);
nand U19073 (N_19073,N_18763,N_18964);
and U19074 (N_19074,N_18856,N_18859);
nand U19075 (N_19075,N_18869,N_18816);
nand U19076 (N_19076,N_18822,N_18829);
and U19077 (N_19077,N_18993,N_18762);
nor U19078 (N_19078,N_18821,N_18828);
and U19079 (N_19079,N_18910,N_18933);
and U19080 (N_19080,N_18916,N_18904);
nand U19081 (N_19081,N_18760,N_18922);
nor U19082 (N_19082,N_18764,N_18902);
or U19083 (N_19083,N_18847,N_18915);
and U19084 (N_19084,N_18977,N_18757);
or U19085 (N_19085,N_18886,N_18880);
or U19086 (N_19086,N_18983,N_18928);
and U19087 (N_19087,N_18782,N_18810);
nor U19088 (N_19088,N_18773,N_18797);
and U19089 (N_19089,N_18908,N_18766);
nand U19090 (N_19090,N_18921,N_18818);
or U19091 (N_19091,N_18961,N_18761);
nor U19092 (N_19092,N_18909,N_18955);
nor U19093 (N_19093,N_18870,N_18942);
and U19094 (N_19094,N_18787,N_18871);
xor U19095 (N_19095,N_18969,N_18804);
xnor U19096 (N_19096,N_18887,N_18949);
and U19097 (N_19097,N_18882,N_18917);
xor U19098 (N_19098,N_18768,N_18895);
and U19099 (N_19099,N_18780,N_18756);
or U19100 (N_19100,N_18815,N_18833);
nor U19101 (N_19101,N_18984,N_18901);
nand U19102 (N_19102,N_18944,N_18838);
or U19103 (N_19103,N_18785,N_18784);
xor U19104 (N_19104,N_18853,N_18982);
nand U19105 (N_19105,N_18750,N_18827);
and U19106 (N_19106,N_18947,N_18772);
and U19107 (N_19107,N_18789,N_18867);
nor U19108 (N_19108,N_18825,N_18937);
or U19109 (N_19109,N_18767,N_18863);
and U19110 (N_19110,N_18862,N_18912);
or U19111 (N_19111,N_18924,N_18998);
or U19112 (N_19112,N_18992,N_18777);
or U19113 (N_19113,N_18776,N_18793);
and U19114 (N_19114,N_18938,N_18981);
xor U19115 (N_19115,N_18996,N_18839);
xor U19116 (N_19116,N_18991,N_18907);
nand U19117 (N_19117,N_18771,N_18788);
and U19118 (N_19118,N_18842,N_18819);
or U19119 (N_19119,N_18914,N_18874);
or U19120 (N_19120,N_18935,N_18896);
and U19121 (N_19121,N_18892,N_18786);
or U19122 (N_19122,N_18866,N_18972);
nand U19123 (N_19123,N_18832,N_18973);
xor U19124 (N_19124,N_18824,N_18918);
nand U19125 (N_19125,N_18985,N_18902);
xor U19126 (N_19126,N_18758,N_18978);
nand U19127 (N_19127,N_18838,N_18915);
nor U19128 (N_19128,N_18842,N_18808);
xnor U19129 (N_19129,N_18876,N_18763);
or U19130 (N_19130,N_18935,N_18817);
xor U19131 (N_19131,N_18946,N_18955);
xor U19132 (N_19132,N_18767,N_18904);
nor U19133 (N_19133,N_18870,N_18966);
nor U19134 (N_19134,N_18832,N_18865);
or U19135 (N_19135,N_18994,N_18801);
and U19136 (N_19136,N_18882,N_18870);
or U19137 (N_19137,N_18993,N_18922);
xor U19138 (N_19138,N_18906,N_18804);
nand U19139 (N_19139,N_18802,N_18946);
xor U19140 (N_19140,N_18867,N_18878);
nor U19141 (N_19141,N_18856,N_18793);
and U19142 (N_19142,N_18969,N_18752);
or U19143 (N_19143,N_18792,N_18959);
and U19144 (N_19144,N_18847,N_18914);
or U19145 (N_19145,N_18930,N_18916);
and U19146 (N_19146,N_18920,N_18815);
or U19147 (N_19147,N_18946,N_18855);
nor U19148 (N_19148,N_18779,N_18962);
nand U19149 (N_19149,N_18767,N_18750);
and U19150 (N_19150,N_18937,N_18768);
and U19151 (N_19151,N_18906,N_18786);
nor U19152 (N_19152,N_18921,N_18987);
or U19153 (N_19153,N_18969,N_18992);
nor U19154 (N_19154,N_18813,N_18921);
nor U19155 (N_19155,N_18938,N_18869);
and U19156 (N_19156,N_18948,N_18885);
or U19157 (N_19157,N_18846,N_18993);
or U19158 (N_19158,N_18913,N_18766);
nor U19159 (N_19159,N_18912,N_18908);
and U19160 (N_19160,N_18988,N_18764);
or U19161 (N_19161,N_18919,N_18836);
xnor U19162 (N_19162,N_18814,N_18835);
nand U19163 (N_19163,N_18880,N_18965);
or U19164 (N_19164,N_18836,N_18911);
nor U19165 (N_19165,N_18796,N_18870);
and U19166 (N_19166,N_18928,N_18788);
xor U19167 (N_19167,N_18818,N_18983);
and U19168 (N_19168,N_18750,N_18831);
or U19169 (N_19169,N_18946,N_18993);
nand U19170 (N_19170,N_18805,N_18754);
nand U19171 (N_19171,N_18950,N_18884);
xor U19172 (N_19172,N_18902,N_18757);
or U19173 (N_19173,N_18915,N_18874);
nor U19174 (N_19174,N_18925,N_18833);
and U19175 (N_19175,N_18755,N_18915);
or U19176 (N_19176,N_18918,N_18934);
or U19177 (N_19177,N_18920,N_18756);
nand U19178 (N_19178,N_18983,N_18934);
and U19179 (N_19179,N_18813,N_18808);
xnor U19180 (N_19180,N_18907,N_18926);
nor U19181 (N_19181,N_18769,N_18831);
nand U19182 (N_19182,N_18933,N_18836);
xor U19183 (N_19183,N_18862,N_18996);
and U19184 (N_19184,N_18932,N_18899);
xor U19185 (N_19185,N_18939,N_18914);
and U19186 (N_19186,N_18840,N_18888);
xor U19187 (N_19187,N_18825,N_18952);
nand U19188 (N_19188,N_18952,N_18809);
or U19189 (N_19189,N_18773,N_18972);
and U19190 (N_19190,N_18789,N_18877);
xnor U19191 (N_19191,N_18867,N_18922);
or U19192 (N_19192,N_18833,N_18882);
nand U19193 (N_19193,N_18778,N_18851);
xor U19194 (N_19194,N_18859,N_18948);
xor U19195 (N_19195,N_18812,N_18984);
nor U19196 (N_19196,N_18961,N_18841);
xnor U19197 (N_19197,N_18776,N_18959);
nand U19198 (N_19198,N_18882,N_18869);
xor U19199 (N_19199,N_18937,N_18787);
nand U19200 (N_19200,N_18898,N_18870);
nor U19201 (N_19201,N_18985,N_18895);
nor U19202 (N_19202,N_18923,N_18949);
xnor U19203 (N_19203,N_18962,N_18906);
and U19204 (N_19204,N_18968,N_18852);
nand U19205 (N_19205,N_18784,N_18815);
nor U19206 (N_19206,N_18776,N_18831);
nor U19207 (N_19207,N_18967,N_18954);
nand U19208 (N_19208,N_18848,N_18833);
or U19209 (N_19209,N_18890,N_18835);
xor U19210 (N_19210,N_18880,N_18852);
nor U19211 (N_19211,N_18767,N_18940);
nor U19212 (N_19212,N_18906,N_18865);
nand U19213 (N_19213,N_18848,N_18924);
or U19214 (N_19214,N_18815,N_18782);
nand U19215 (N_19215,N_18924,N_18864);
nand U19216 (N_19216,N_18812,N_18819);
or U19217 (N_19217,N_18849,N_18991);
nand U19218 (N_19218,N_18835,N_18759);
or U19219 (N_19219,N_18805,N_18927);
xnor U19220 (N_19220,N_18803,N_18906);
xor U19221 (N_19221,N_18983,N_18861);
xnor U19222 (N_19222,N_18792,N_18858);
and U19223 (N_19223,N_18899,N_18769);
xor U19224 (N_19224,N_18927,N_18840);
nor U19225 (N_19225,N_18939,N_18762);
or U19226 (N_19226,N_18972,N_18858);
and U19227 (N_19227,N_18993,N_18967);
nand U19228 (N_19228,N_18773,N_18805);
or U19229 (N_19229,N_18797,N_18834);
nand U19230 (N_19230,N_18910,N_18770);
or U19231 (N_19231,N_18842,N_18886);
xnor U19232 (N_19232,N_18934,N_18870);
or U19233 (N_19233,N_18943,N_18872);
and U19234 (N_19234,N_18909,N_18996);
nand U19235 (N_19235,N_18764,N_18771);
nor U19236 (N_19236,N_18908,N_18881);
nand U19237 (N_19237,N_18933,N_18783);
nor U19238 (N_19238,N_18940,N_18967);
and U19239 (N_19239,N_18840,N_18941);
or U19240 (N_19240,N_18991,N_18940);
and U19241 (N_19241,N_18798,N_18782);
nor U19242 (N_19242,N_18939,N_18783);
nand U19243 (N_19243,N_18905,N_18823);
xor U19244 (N_19244,N_18811,N_18924);
or U19245 (N_19245,N_18782,N_18917);
xor U19246 (N_19246,N_18797,N_18838);
and U19247 (N_19247,N_18756,N_18951);
nand U19248 (N_19248,N_18775,N_18915);
and U19249 (N_19249,N_18934,N_18944);
nand U19250 (N_19250,N_19242,N_19065);
and U19251 (N_19251,N_19039,N_19161);
nand U19252 (N_19252,N_19213,N_19071);
and U19253 (N_19253,N_19063,N_19077);
nor U19254 (N_19254,N_19171,N_19235);
xnor U19255 (N_19255,N_19234,N_19222);
xnor U19256 (N_19256,N_19047,N_19055);
or U19257 (N_19257,N_19126,N_19033);
xor U19258 (N_19258,N_19231,N_19069);
nand U19259 (N_19259,N_19109,N_19100);
or U19260 (N_19260,N_19167,N_19113);
nor U19261 (N_19261,N_19059,N_19087);
or U19262 (N_19262,N_19203,N_19229);
nor U19263 (N_19263,N_19225,N_19134);
nor U19264 (N_19264,N_19074,N_19156);
xor U19265 (N_19265,N_19004,N_19137);
and U19266 (N_19266,N_19147,N_19185);
nor U19267 (N_19267,N_19014,N_19226);
and U19268 (N_19268,N_19221,N_19043);
or U19269 (N_19269,N_19017,N_19067);
nand U19270 (N_19270,N_19085,N_19159);
or U19271 (N_19271,N_19052,N_19114);
and U19272 (N_19272,N_19209,N_19204);
nor U19273 (N_19273,N_19243,N_19150);
xnor U19274 (N_19274,N_19062,N_19000);
or U19275 (N_19275,N_19086,N_19018);
or U19276 (N_19276,N_19034,N_19178);
nor U19277 (N_19277,N_19236,N_19093);
or U19278 (N_19278,N_19123,N_19041);
and U19279 (N_19279,N_19102,N_19198);
and U19280 (N_19280,N_19073,N_19125);
nor U19281 (N_19281,N_19241,N_19206);
nor U19282 (N_19282,N_19180,N_19082);
xor U19283 (N_19283,N_19094,N_19054);
or U19284 (N_19284,N_19163,N_19110);
nor U19285 (N_19285,N_19160,N_19248);
and U19286 (N_19286,N_19030,N_19058);
or U19287 (N_19287,N_19090,N_19037);
nand U19288 (N_19288,N_19057,N_19227);
nor U19289 (N_19289,N_19189,N_19076);
or U19290 (N_19290,N_19157,N_19146);
and U19291 (N_19291,N_19068,N_19002);
or U19292 (N_19292,N_19128,N_19220);
and U19293 (N_19293,N_19215,N_19207);
or U19294 (N_19294,N_19119,N_19194);
or U19295 (N_19295,N_19045,N_19066);
xor U19296 (N_19296,N_19122,N_19029);
or U19297 (N_19297,N_19024,N_19210);
xnor U19298 (N_19298,N_19032,N_19035);
or U19299 (N_19299,N_19195,N_19028);
nand U19300 (N_19300,N_19211,N_19244);
or U19301 (N_19301,N_19188,N_19232);
nand U19302 (N_19302,N_19246,N_19208);
or U19303 (N_19303,N_19112,N_19048);
xnor U19304 (N_19304,N_19120,N_19136);
or U19305 (N_19305,N_19214,N_19140);
nor U19306 (N_19306,N_19240,N_19031);
and U19307 (N_19307,N_19239,N_19182);
or U19308 (N_19308,N_19199,N_19154);
nand U19309 (N_19309,N_19133,N_19139);
or U19310 (N_19310,N_19165,N_19061);
xnor U19311 (N_19311,N_19238,N_19155);
nor U19312 (N_19312,N_19135,N_19174);
nand U19313 (N_19313,N_19092,N_19224);
xor U19314 (N_19314,N_19015,N_19044);
and U19315 (N_19315,N_19084,N_19183);
and U19316 (N_19316,N_19172,N_19022);
and U19317 (N_19317,N_19237,N_19078);
nor U19318 (N_19318,N_19151,N_19149);
or U19319 (N_19319,N_19091,N_19027);
xor U19320 (N_19320,N_19008,N_19103);
and U19321 (N_19321,N_19104,N_19212);
nand U19322 (N_19322,N_19141,N_19184);
nand U19323 (N_19323,N_19095,N_19176);
and U19324 (N_19324,N_19181,N_19101);
nor U19325 (N_19325,N_19132,N_19191);
xnor U19326 (N_19326,N_19205,N_19042);
and U19327 (N_19327,N_19096,N_19193);
xor U19328 (N_19328,N_19168,N_19072);
nor U19329 (N_19329,N_19023,N_19124);
nand U19330 (N_19330,N_19010,N_19144);
and U19331 (N_19331,N_19088,N_19127);
xnor U19332 (N_19332,N_19164,N_19046);
nor U19333 (N_19333,N_19005,N_19006);
and U19334 (N_19334,N_19097,N_19064);
or U19335 (N_19335,N_19169,N_19099);
or U19336 (N_19336,N_19173,N_19200);
nand U19337 (N_19337,N_19179,N_19056);
and U19338 (N_19338,N_19158,N_19186);
nor U19339 (N_19339,N_19051,N_19129);
xnor U19340 (N_19340,N_19011,N_19075);
or U19341 (N_19341,N_19040,N_19049);
xnor U19342 (N_19342,N_19007,N_19247);
nor U19343 (N_19343,N_19009,N_19217);
nand U19344 (N_19344,N_19013,N_19121);
and U19345 (N_19345,N_19107,N_19079);
xnor U19346 (N_19346,N_19148,N_19142);
or U19347 (N_19347,N_19116,N_19245);
xnor U19348 (N_19348,N_19001,N_19152);
nor U19349 (N_19349,N_19138,N_19021);
xnor U19350 (N_19350,N_19190,N_19233);
or U19351 (N_19351,N_19228,N_19016);
nor U19352 (N_19352,N_19131,N_19130);
nor U19353 (N_19353,N_19105,N_19166);
and U19354 (N_19354,N_19050,N_19162);
nand U19355 (N_19355,N_19080,N_19098);
nor U19356 (N_19356,N_19216,N_19223);
nand U19357 (N_19357,N_19115,N_19038);
xor U19358 (N_19358,N_19019,N_19025);
or U19359 (N_19359,N_19143,N_19053);
xnor U19360 (N_19360,N_19145,N_19196);
xnor U19361 (N_19361,N_19197,N_19036);
nand U19362 (N_19362,N_19153,N_19117);
or U19363 (N_19363,N_19170,N_19249);
xnor U19364 (N_19364,N_19106,N_19089);
xor U19365 (N_19365,N_19020,N_19012);
xor U19366 (N_19366,N_19230,N_19175);
nand U19367 (N_19367,N_19202,N_19081);
nand U19368 (N_19368,N_19118,N_19111);
nor U19369 (N_19369,N_19192,N_19060);
or U19370 (N_19370,N_19219,N_19083);
nor U19371 (N_19371,N_19201,N_19026);
nor U19372 (N_19372,N_19187,N_19177);
nand U19373 (N_19373,N_19218,N_19070);
or U19374 (N_19374,N_19003,N_19108);
nor U19375 (N_19375,N_19176,N_19200);
and U19376 (N_19376,N_19221,N_19233);
nand U19377 (N_19377,N_19083,N_19072);
nor U19378 (N_19378,N_19249,N_19143);
xor U19379 (N_19379,N_19024,N_19113);
nor U19380 (N_19380,N_19179,N_19082);
xor U19381 (N_19381,N_19070,N_19169);
and U19382 (N_19382,N_19217,N_19121);
nand U19383 (N_19383,N_19121,N_19027);
xnor U19384 (N_19384,N_19166,N_19058);
or U19385 (N_19385,N_19195,N_19213);
or U19386 (N_19386,N_19000,N_19018);
nand U19387 (N_19387,N_19030,N_19214);
or U19388 (N_19388,N_19031,N_19177);
or U19389 (N_19389,N_19149,N_19240);
and U19390 (N_19390,N_19074,N_19147);
nor U19391 (N_19391,N_19117,N_19072);
nor U19392 (N_19392,N_19144,N_19121);
or U19393 (N_19393,N_19083,N_19158);
nor U19394 (N_19394,N_19172,N_19108);
or U19395 (N_19395,N_19035,N_19172);
nand U19396 (N_19396,N_19085,N_19221);
nor U19397 (N_19397,N_19051,N_19081);
xnor U19398 (N_19398,N_19077,N_19085);
or U19399 (N_19399,N_19005,N_19009);
nand U19400 (N_19400,N_19223,N_19049);
and U19401 (N_19401,N_19110,N_19087);
nand U19402 (N_19402,N_19222,N_19157);
nor U19403 (N_19403,N_19006,N_19243);
or U19404 (N_19404,N_19062,N_19144);
nand U19405 (N_19405,N_19192,N_19059);
xnor U19406 (N_19406,N_19044,N_19220);
xor U19407 (N_19407,N_19190,N_19195);
and U19408 (N_19408,N_19153,N_19091);
nand U19409 (N_19409,N_19055,N_19042);
and U19410 (N_19410,N_19157,N_19006);
nand U19411 (N_19411,N_19138,N_19052);
nor U19412 (N_19412,N_19069,N_19000);
nand U19413 (N_19413,N_19168,N_19243);
or U19414 (N_19414,N_19101,N_19025);
nand U19415 (N_19415,N_19190,N_19177);
or U19416 (N_19416,N_19125,N_19128);
nand U19417 (N_19417,N_19101,N_19034);
nor U19418 (N_19418,N_19184,N_19209);
and U19419 (N_19419,N_19136,N_19245);
or U19420 (N_19420,N_19162,N_19017);
nand U19421 (N_19421,N_19210,N_19058);
nand U19422 (N_19422,N_19132,N_19217);
or U19423 (N_19423,N_19224,N_19161);
and U19424 (N_19424,N_19007,N_19109);
and U19425 (N_19425,N_19238,N_19131);
or U19426 (N_19426,N_19051,N_19171);
nor U19427 (N_19427,N_19032,N_19165);
xor U19428 (N_19428,N_19102,N_19046);
and U19429 (N_19429,N_19112,N_19045);
or U19430 (N_19430,N_19069,N_19152);
xnor U19431 (N_19431,N_19235,N_19020);
nand U19432 (N_19432,N_19124,N_19110);
or U19433 (N_19433,N_19152,N_19137);
nor U19434 (N_19434,N_19227,N_19006);
or U19435 (N_19435,N_19197,N_19075);
nor U19436 (N_19436,N_19216,N_19209);
nand U19437 (N_19437,N_19083,N_19060);
nor U19438 (N_19438,N_19181,N_19054);
and U19439 (N_19439,N_19041,N_19146);
nor U19440 (N_19440,N_19025,N_19112);
xnor U19441 (N_19441,N_19193,N_19077);
xnor U19442 (N_19442,N_19173,N_19202);
nor U19443 (N_19443,N_19246,N_19153);
nand U19444 (N_19444,N_19166,N_19022);
nand U19445 (N_19445,N_19234,N_19121);
nand U19446 (N_19446,N_19203,N_19002);
nor U19447 (N_19447,N_19159,N_19022);
nor U19448 (N_19448,N_19075,N_19088);
nand U19449 (N_19449,N_19108,N_19228);
nor U19450 (N_19450,N_19138,N_19227);
xnor U19451 (N_19451,N_19062,N_19045);
nor U19452 (N_19452,N_19243,N_19225);
or U19453 (N_19453,N_19150,N_19164);
and U19454 (N_19454,N_19045,N_19124);
or U19455 (N_19455,N_19059,N_19014);
xor U19456 (N_19456,N_19060,N_19010);
and U19457 (N_19457,N_19087,N_19082);
nor U19458 (N_19458,N_19238,N_19150);
xnor U19459 (N_19459,N_19090,N_19102);
nor U19460 (N_19460,N_19185,N_19016);
xor U19461 (N_19461,N_19232,N_19234);
and U19462 (N_19462,N_19108,N_19135);
and U19463 (N_19463,N_19027,N_19048);
and U19464 (N_19464,N_19245,N_19048);
xor U19465 (N_19465,N_19022,N_19100);
and U19466 (N_19466,N_19142,N_19077);
nand U19467 (N_19467,N_19129,N_19183);
and U19468 (N_19468,N_19184,N_19051);
nor U19469 (N_19469,N_19239,N_19046);
and U19470 (N_19470,N_19046,N_19165);
or U19471 (N_19471,N_19239,N_19131);
nand U19472 (N_19472,N_19182,N_19202);
xor U19473 (N_19473,N_19138,N_19190);
nand U19474 (N_19474,N_19229,N_19228);
and U19475 (N_19475,N_19163,N_19085);
xor U19476 (N_19476,N_19017,N_19146);
or U19477 (N_19477,N_19168,N_19164);
xnor U19478 (N_19478,N_19191,N_19008);
nor U19479 (N_19479,N_19218,N_19140);
nand U19480 (N_19480,N_19127,N_19115);
or U19481 (N_19481,N_19235,N_19024);
nand U19482 (N_19482,N_19213,N_19074);
nand U19483 (N_19483,N_19043,N_19105);
and U19484 (N_19484,N_19191,N_19183);
nor U19485 (N_19485,N_19224,N_19145);
nor U19486 (N_19486,N_19087,N_19079);
xnor U19487 (N_19487,N_19112,N_19058);
nor U19488 (N_19488,N_19122,N_19047);
nand U19489 (N_19489,N_19042,N_19032);
xor U19490 (N_19490,N_19054,N_19000);
and U19491 (N_19491,N_19077,N_19044);
and U19492 (N_19492,N_19112,N_19071);
nor U19493 (N_19493,N_19173,N_19118);
or U19494 (N_19494,N_19006,N_19178);
nand U19495 (N_19495,N_19091,N_19140);
nand U19496 (N_19496,N_19081,N_19168);
xor U19497 (N_19497,N_19094,N_19088);
nor U19498 (N_19498,N_19141,N_19118);
nand U19499 (N_19499,N_19176,N_19083);
nand U19500 (N_19500,N_19316,N_19306);
and U19501 (N_19501,N_19479,N_19486);
nand U19502 (N_19502,N_19391,N_19473);
xnor U19503 (N_19503,N_19299,N_19385);
and U19504 (N_19504,N_19492,N_19453);
nand U19505 (N_19505,N_19363,N_19365);
nand U19506 (N_19506,N_19433,N_19389);
nor U19507 (N_19507,N_19472,N_19328);
or U19508 (N_19508,N_19258,N_19387);
or U19509 (N_19509,N_19330,N_19415);
or U19510 (N_19510,N_19458,N_19418);
or U19511 (N_19511,N_19264,N_19375);
nor U19512 (N_19512,N_19430,N_19283);
nand U19513 (N_19513,N_19441,N_19411);
nor U19514 (N_19514,N_19301,N_19340);
xor U19515 (N_19515,N_19321,N_19424);
nand U19516 (N_19516,N_19317,N_19344);
nor U19517 (N_19517,N_19262,N_19488);
xor U19518 (N_19518,N_19390,N_19445);
nor U19519 (N_19519,N_19276,N_19295);
or U19520 (N_19520,N_19482,N_19428);
xnor U19521 (N_19521,N_19468,N_19280);
nand U19522 (N_19522,N_19480,N_19393);
xnor U19523 (N_19523,N_19290,N_19416);
nor U19524 (N_19524,N_19379,N_19487);
nor U19525 (N_19525,N_19271,N_19279);
nor U19526 (N_19526,N_19454,N_19267);
nor U19527 (N_19527,N_19339,N_19254);
nand U19528 (N_19528,N_19308,N_19382);
nand U19529 (N_19529,N_19310,N_19263);
xor U19530 (N_19530,N_19449,N_19348);
xor U19531 (N_19531,N_19498,N_19384);
xnor U19532 (N_19532,N_19327,N_19476);
and U19533 (N_19533,N_19253,N_19402);
or U19534 (N_19534,N_19332,N_19451);
and U19535 (N_19535,N_19426,N_19423);
or U19536 (N_19536,N_19368,N_19297);
nor U19537 (N_19537,N_19336,N_19256);
and U19538 (N_19538,N_19434,N_19437);
nand U19539 (N_19539,N_19350,N_19272);
nand U19540 (N_19540,N_19376,N_19354);
or U19541 (N_19541,N_19431,N_19329);
nor U19542 (N_19542,N_19404,N_19252);
nand U19543 (N_19543,N_19392,N_19410);
or U19544 (N_19544,N_19489,N_19395);
and U19545 (N_19545,N_19323,N_19398);
or U19546 (N_19546,N_19381,N_19491);
or U19547 (N_19547,N_19353,N_19470);
nand U19548 (N_19548,N_19285,N_19464);
nor U19549 (N_19549,N_19360,N_19409);
xor U19550 (N_19550,N_19369,N_19364);
and U19551 (N_19551,N_19361,N_19324);
xnor U19552 (N_19552,N_19477,N_19420);
nor U19553 (N_19553,N_19266,N_19394);
or U19554 (N_19554,N_19335,N_19338);
nor U19555 (N_19555,N_19417,N_19261);
and U19556 (N_19556,N_19461,N_19446);
nand U19557 (N_19557,N_19471,N_19343);
or U19558 (N_19558,N_19463,N_19269);
or U19559 (N_19559,N_19311,N_19282);
xor U19560 (N_19560,N_19366,N_19302);
and U19561 (N_19561,N_19425,N_19495);
and U19562 (N_19562,N_19435,N_19352);
nand U19563 (N_19563,N_19304,N_19377);
xor U19564 (N_19564,N_19483,N_19315);
nor U19565 (N_19565,N_19460,N_19259);
nor U19566 (N_19566,N_19351,N_19403);
or U19567 (N_19567,N_19481,N_19443);
nand U19568 (N_19568,N_19478,N_19313);
xor U19569 (N_19569,N_19422,N_19293);
nand U19570 (N_19570,N_19331,N_19439);
and U19571 (N_19571,N_19493,N_19419);
or U19572 (N_19572,N_19257,N_19292);
nand U19573 (N_19573,N_19341,N_19450);
nand U19574 (N_19574,N_19396,N_19432);
and U19575 (N_19575,N_19260,N_19462);
xnor U19576 (N_19576,N_19337,N_19499);
xnor U19577 (N_19577,N_19345,N_19288);
xnor U19578 (N_19578,N_19320,N_19270);
nand U19579 (N_19579,N_19265,N_19326);
xor U19580 (N_19580,N_19303,N_19277);
xnor U19581 (N_19581,N_19347,N_19342);
nor U19582 (N_19582,N_19444,N_19406);
xnor U19583 (N_19583,N_19494,N_19380);
nor U19584 (N_19584,N_19325,N_19319);
or U19585 (N_19585,N_19485,N_19378);
xor U19586 (N_19586,N_19452,N_19372);
or U19587 (N_19587,N_19250,N_19408);
xor U19588 (N_19588,N_19405,N_19436);
xor U19589 (N_19589,N_19287,N_19346);
nor U19590 (N_19590,N_19412,N_19414);
nor U19591 (N_19591,N_19278,N_19309);
or U19592 (N_19592,N_19255,N_19274);
xor U19593 (N_19593,N_19466,N_19318);
or U19594 (N_19594,N_19307,N_19300);
and U19595 (N_19595,N_19251,N_19497);
nor U19596 (N_19596,N_19362,N_19281);
nand U19597 (N_19597,N_19356,N_19355);
xor U19598 (N_19598,N_19291,N_19371);
nand U19599 (N_19599,N_19349,N_19275);
and U19600 (N_19600,N_19490,N_19370);
nor U19601 (N_19601,N_19457,N_19289);
nor U19602 (N_19602,N_19484,N_19438);
and U19603 (N_19603,N_19474,N_19284);
or U19604 (N_19604,N_19427,N_19407);
or U19605 (N_19605,N_19294,N_19400);
or U19606 (N_19606,N_19383,N_19469);
and U19607 (N_19607,N_19440,N_19322);
and U19608 (N_19608,N_19373,N_19312);
nand U19609 (N_19609,N_19268,N_19399);
or U19610 (N_19610,N_19496,N_19388);
or U19611 (N_19611,N_19357,N_19413);
xor U19612 (N_19612,N_19459,N_19298);
or U19613 (N_19613,N_19456,N_19273);
nand U19614 (N_19614,N_19367,N_19467);
nand U19615 (N_19615,N_19447,N_19314);
nand U19616 (N_19616,N_19455,N_19397);
xor U19617 (N_19617,N_19475,N_19286);
and U19618 (N_19618,N_19429,N_19334);
nor U19619 (N_19619,N_19465,N_19448);
xnor U19620 (N_19620,N_19421,N_19359);
and U19621 (N_19621,N_19358,N_19305);
and U19622 (N_19622,N_19442,N_19296);
or U19623 (N_19623,N_19386,N_19333);
nor U19624 (N_19624,N_19401,N_19374);
xor U19625 (N_19625,N_19430,N_19292);
xor U19626 (N_19626,N_19284,N_19394);
and U19627 (N_19627,N_19348,N_19422);
and U19628 (N_19628,N_19490,N_19371);
and U19629 (N_19629,N_19320,N_19407);
nor U19630 (N_19630,N_19276,N_19334);
or U19631 (N_19631,N_19335,N_19385);
and U19632 (N_19632,N_19398,N_19446);
nand U19633 (N_19633,N_19383,N_19410);
or U19634 (N_19634,N_19410,N_19271);
and U19635 (N_19635,N_19429,N_19293);
nor U19636 (N_19636,N_19375,N_19448);
and U19637 (N_19637,N_19359,N_19361);
and U19638 (N_19638,N_19438,N_19411);
and U19639 (N_19639,N_19453,N_19428);
nor U19640 (N_19640,N_19397,N_19404);
xnor U19641 (N_19641,N_19467,N_19341);
nor U19642 (N_19642,N_19323,N_19251);
nand U19643 (N_19643,N_19338,N_19275);
and U19644 (N_19644,N_19276,N_19378);
nand U19645 (N_19645,N_19441,N_19270);
nor U19646 (N_19646,N_19257,N_19416);
and U19647 (N_19647,N_19361,N_19405);
nand U19648 (N_19648,N_19449,N_19483);
nor U19649 (N_19649,N_19315,N_19462);
nand U19650 (N_19650,N_19322,N_19471);
xnor U19651 (N_19651,N_19383,N_19437);
nor U19652 (N_19652,N_19479,N_19388);
nand U19653 (N_19653,N_19380,N_19289);
nor U19654 (N_19654,N_19409,N_19287);
xnor U19655 (N_19655,N_19447,N_19256);
nand U19656 (N_19656,N_19351,N_19325);
and U19657 (N_19657,N_19423,N_19311);
and U19658 (N_19658,N_19362,N_19408);
or U19659 (N_19659,N_19263,N_19322);
nand U19660 (N_19660,N_19418,N_19337);
or U19661 (N_19661,N_19331,N_19270);
nor U19662 (N_19662,N_19483,N_19459);
xor U19663 (N_19663,N_19436,N_19481);
nand U19664 (N_19664,N_19259,N_19368);
or U19665 (N_19665,N_19276,N_19487);
nor U19666 (N_19666,N_19303,N_19352);
nand U19667 (N_19667,N_19428,N_19315);
nand U19668 (N_19668,N_19498,N_19454);
xor U19669 (N_19669,N_19392,N_19290);
nand U19670 (N_19670,N_19295,N_19308);
nor U19671 (N_19671,N_19315,N_19484);
or U19672 (N_19672,N_19343,N_19446);
and U19673 (N_19673,N_19273,N_19495);
xor U19674 (N_19674,N_19427,N_19305);
nand U19675 (N_19675,N_19348,N_19409);
xor U19676 (N_19676,N_19491,N_19300);
xnor U19677 (N_19677,N_19415,N_19440);
and U19678 (N_19678,N_19265,N_19370);
xor U19679 (N_19679,N_19305,N_19396);
nor U19680 (N_19680,N_19365,N_19268);
nor U19681 (N_19681,N_19360,N_19478);
xnor U19682 (N_19682,N_19387,N_19344);
nor U19683 (N_19683,N_19321,N_19280);
or U19684 (N_19684,N_19449,N_19314);
xnor U19685 (N_19685,N_19397,N_19259);
and U19686 (N_19686,N_19407,N_19382);
xnor U19687 (N_19687,N_19421,N_19465);
nand U19688 (N_19688,N_19336,N_19268);
nor U19689 (N_19689,N_19340,N_19376);
or U19690 (N_19690,N_19378,N_19293);
and U19691 (N_19691,N_19478,N_19475);
nand U19692 (N_19692,N_19467,N_19416);
xnor U19693 (N_19693,N_19468,N_19484);
and U19694 (N_19694,N_19331,N_19285);
nand U19695 (N_19695,N_19431,N_19324);
nand U19696 (N_19696,N_19484,N_19409);
nand U19697 (N_19697,N_19256,N_19310);
nor U19698 (N_19698,N_19495,N_19453);
nand U19699 (N_19699,N_19390,N_19299);
nor U19700 (N_19700,N_19470,N_19387);
nor U19701 (N_19701,N_19490,N_19492);
nor U19702 (N_19702,N_19298,N_19334);
nor U19703 (N_19703,N_19293,N_19438);
or U19704 (N_19704,N_19279,N_19358);
or U19705 (N_19705,N_19358,N_19336);
xor U19706 (N_19706,N_19389,N_19411);
or U19707 (N_19707,N_19279,N_19289);
and U19708 (N_19708,N_19300,N_19367);
nand U19709 (N_19709,N_19328,N_19377);
and U19710 (N_19710,N_19471,N_19314);
xor U19711 (N_19711,N_19262,N_19327);
and U19712 (N_19712,N_19325,N_19476);
nor U19713 (N_19713,N_19310,N_19396);
or U19714 (N_19714,N_19300,N_19312);
nor U19715 (N_19715,N_19390,N_19287);
or U19716 (N_19716,N_19483,N_19326);
and U19717 (N_19717,N_19376,N_19327);
and U19718 (N_19718,N_19351,N_19393);
and U19719 (N_19719,N_19340,N_19393);
and U19720 (N_19720,N_19334,N_19296);
and U19721 (N_19721,N_19259,N_19385);
nand U19722 (N_19722,N_19413,N_19409);
nor U19723 (N_19723,N_19353,N_19400);
and U19724 (N_19724,N_19336,N_19425);
nor U19725 (N_19725,N_19469,N_19441);
and U19726 (N_19726,N_19304,N_19484);
xnor U19727 (N_19727,N_19278,N_19372);
and U19728 (N_19728,N_19434,N_19299);
nand U19729 (N_19729,N_19390,N_19408);
or U19730 (N_19730,N_19383,N_19398);
nand U19731 (N_19731,N_19436,N_19466);
or U19732 (N_19732,N_19446,N_19271);
xnor U19733 (N_19733,N_19457,N_19385);
and U19734 (N_19734,N_19429,N_19276);
or U19735 (N_19735,N_19471,N_19281);
xnor U19736 (N_19736,N_19306,N_19383);
and U19737 (N_19737,N_19351,N_19484);
nor U19738 (N_19738,N_19321,N_19320);
and U19739 (N_19739,N_19451,N_19470);
or U19740 (N_19740,N_19290,N_19498);
nor U19741 (N_19741,N_19344,N_19288);
xnor U19742 (N_19742,N_19402,N_19276);
nor U19743 (N_19743,N_19464,N_19327);
xnor U19744 (N_19744,N_19318,N_19372);
xor U19745 (N_19745,N_19271,N_19463);
nand U19746 (N_19746,N_19445,N_19434);
and U19747 (N_19747,N_19429,N_19321);
and U19748 (N_19748,N_19499,N_19268);
or U19749 (N_19749,N_19414,N_19431);
or U19750 (N_19750,N_19710,N_19665);
xnor U19751 (N_19751,N_19656,N_19550);
nor U19752 (N_19752,N_19732,N_19531);
nand U19753 (N_19753,N_19639,N_19622);
xnor U19754 (N_19754,N_19613,N_19611);
or U19755 (N_19755,N_19529,N_19659);
nand U19756 (N_19756,N_19620,N_19609);
and U19757 (N_19757,N_19733,N_19647);
xor U19758 (N_19758,N_19712,N_19553);
and U19759 (N_19759,N_19561,N_19560);
and U19760 (N_19760,N_19558,N_19722);
or U19761 (N_19761,N_19597,N_19500);
xnor U19762 (N_19762,N_19690,N_19688);
nand U19763 (N_19763,N_19593,N_19739);
nor U19764 (N_19764,N_19705,N_19540);
nand U19765 (N_19765,N_19654,N_19687);
or U19766 (N_19766,N_19582,N_19693);
xor U19767 (N_19767,N_19542,N_19651);
and U19768 (N_19768,N_19644,N_19581);
nand U19769 (N_19769,N_19533,N_19695);
nor U19770 (N_19770,N_19745,N_19616);
or U19771 (N_19771,N_19524,N_19747);
or U19772 (N_19772,N_19727,N_19641);
and U19773 (N_19773,N_19668,N_19617);
nand U19774 (N_19774,N_19743,N_19678);
or U19775 (N_19775,N_19569,N_19587);
xnor U19776 (N_19776,N_19508,N_19509);
xor U19777 (N_19777,N_19518,N_19543);
or U19778 (N_19778,N_19674,N_19720);
nand U19779 (N_19779,N_19520,N_19541);
xor U19780 (N_19780,N_19697,N_19663);
nor U19781 (N_19781,N_19538,N_19565);
nand U19782 (N_19782,N_19682,N_19592);
nand U19783 (N_19783,N_19692,N_19517);
nor U19784 (N_19784,N_19744,N_19707);
or U19785 (N_19785,N_19606,N_19555);
nand U19786 (N_19786,N_19547,N_19539);
or U19787 (N_19787,N_19655,N_19584);
xnor U19788 (N_19788,N_19574,N_19546);
nor U19789 (N_19789,N_19586,N_19632);
or U19790 (N_19790,N_19568,N_19719);
xor U19791 (N_19791,N_19610,N_19590);
xnor U19792 (N_19792,N_19715,N_19507);
and U19793 (N_19793,N_19698,N_19579);
or U19794 (N_19794,N_19725,N_19686);
xor U19795 (N_19795,N_19679,N_19563);
and U19796 (N_19796,N_19623,N_19528);
nand U19797 (N_19797,N_19573,N_19706);
nor U19798 (N_19798,N_19511,N_19591);
and U19799 (N_19799,N_19530,N_19677);
xor U19800 (N_19800,N_19699,N_19653);
nand U19801 (N_19801,N_19726,N_19634);
nand U19802 (N_19802,N_19571,N_19648);
nand U19803 (N_19803,N_19570,N_19545);
xnor U19804 (N_19804,N_19567,N_19701);
xnor U19805 (N_19805,N_19681,N_19527);
and U19806 (N_19806,N_19556,N_19522);
xnor U19807 (N_19807,N_19514,N_19512);
and U19808 (N_19808,N_19510,N_19615);
nor U19809 (N_19809,N_19661,N_19501);
nor U19810 (N_19810,N_19640,N_19714);
and U19811 (N_19811,N_19519,N_19502);
and U19812 (N_19812,N_19526,N_19628);
or U19813 (N_19813,N_19723,N_19562);
and U19814 (N_19814,N_19607,N_19557);
nor U19815 (N_19815,N_19704,N_19596);
nand U19816 (N_19816,N_19626,N_19601);
nand U19817 (N_19817,N_19564,N_19643);
xnor U19818 (N_19818,N_19552,N_19595);
nor U19819 (N_19819,N_19740,N_19621);
nand U19820 (N_19820,N_19669,N_19629);
nor U19821 (N_19821,N_19716,N_19516);
nor U19822 (N_19822,N_19741,N_19548);
and U19823 (N_19823,N_19635,N_19625);
and U19824 (N_19824,N_19559,N_19506);
or U19825 (N_19825,N_19746,N_19638);
xor U19826 (N_19826,N_19551,N_19742);
or U19827 (N_19827,N_19604,N_19703);
nand U19828 (N_19828,N_19535,N_19709);
nor U19829 (N_19829,N_19721,N_19652);
and U19830 (N_19830,N_19736,N_19670);
and U19831 (N_19831,N_19585,N_19602);
and U19832 (N_19832,N_19589,N_19702);
or U19833 (N_19833,N_19608,N_19749);
nand U19834 (N_19834,N_19650,N_19680);
and U19835 (N_19835,N_19633,N_19594);
xor U19836 (N_19836,N_19624,N_19667);
nor U19837 (N_19837,N_19708,N_19619);
xor U19838 (N_19838,N_19649,N_19694);
or U19839 (N_19839,N_19711,N_19504);
and U19840 (N_19840,N_19673,N_19738);
nand U19841 (N_19841,N_19566,N_19549);
xor U19842 (N_19842,N_19684,N_19689);
and U19843 (N_19843,N_19642,N_19537);
and U19844 (N_19844,N_19691,N_19513);
and U19845 (N_19845,N_19748,N_19627);
nand U19846 (N_19846,N_19718,N_19713);
nand U19847 (N_19847,N_19731,N_19576);
nand U19848 (N_19848,N_19657,N_19532);
or U19849 (N_19849,N_19660,N_19536);
nand U19850 (N_19850,N_19662,N_19729);
and U19851 (N_19851,N_19588,N_19675);
or U19852 (N_19852,N_19631,N_19618);
nand U19853 (N_19853,N_19683,N_19525);
nand U19854 (N_19854,N_19599,N_19717);
or U19855 (N_19855,N_19583,N_19605);
and U19856 (N_19856,N_19521,N_19666);
nor U19857 (N_19857,N_19672,N_19577);
and U19858 (N_19858,N_19598,N_19734);
xor U19859 (N_19859,N_19696,N_19600);
nor U19860 (N_19860,N_19630,N_19730);
xor U19861 (N_19861,N_19737,N_19735);
nor U19862 (N_19862,N_19636,N_19544);
nand U19863 (N_19863,N_19700,N_19523);
and U19864 (N_19864,N_19515,N_19612);
xnor U19865 (N_19865,N_19554,N_19728);
nand U19866 (N_19866,N_19575,N_19724);
nand U19867 (N_19867,N_19572,N_19614);
and U19868 (N_19868,N_19580,N_19578);
nor U19869 (N_19869,N_19603,N_19658);
nand U19870 (N_19870,N_19637,N_19685);
nor U19871 (N_19871,N_19676,N_19505);
or U19872 (N_19872,N_19671,N_19664);
and U19873 (N_19873,N_19503,N_19646);
nand U19874 (N_19874,N_19534,N_19645);
xor U19875 (N_19875,N_19739,N_19505);
or U19876 (N_19876,N_19730,N_19558);
and U19877 (N_19877,N_19682,N_19547);
nand U19878 (N_19878,N_19569,N_19518);
nor U19879 (N_19879,N_19727,N_19737);
nor U19880 (N_19880,N_19685,N_19635);
and U19881 (N_19881,N_19574,N_19638);
nand U19882 (N_19882,N_19746,N_19711);
or U19883 (N_19883,N_19519,N_19678);
nor U19884 (N_19884,N_19507,N_19641);
and U19885 (N_19885,N_19666,N_19715);
nand U19886 (N_19886,N_19615,N_19722);
or U19887 (N_19887,N_19603,N_19531);
xnor U19888 (N_19888,N_19539,N_19516);
xnor U19889 (N_19889,N_19625,N_19661);
xnor U19890 (N_19890,N_19605,N_19640);
nand U19891 (N_19891,N_19580,N_19501);
or U19892 (N_19892,N_19711,N_19524);
and U19893 (N_19893,N_19584,N_19634);
xnor U19894 (N_19894,N_19576,N_19611);
or U19895 (N_19895,N_19594,N_19679);
or U19896 (N_19896,N_19578,N_19554);
nand U19897 (N_19897,N_19597,N_19670);
xnor U19898 (N_19898,N_19731,N_19563);
xor U19899 (N_19899,N_19590,N_19631);
nand U19900 (N_19900,N_19622,N_19664);
and U19901 (N_19901,N_19720,N_19640);
nand U19902 (N_19902,N_19515,N_19706);
nor U19903 (N_19903,N_19742,N_19624);
nand U19904 (N_19904,N_19733,N_19648);
nor U19905 (N_19905,N_19684,N_19525);
nor U19906 (N_19906,N_19683,N_19508);
or U19907 (N_19907,N_19585,N_19600);
and U19908 (N_19908,N_19612,N_19626);
nor U19909 (N_19909,N_19591,N_19680);
nand U19910 (N_19910,N_19602,N_19510);
xor U19911 (N_19911,N_19540,N_19742);
nor U19912 (N_19912,N_19719,N_19582);
and U19913 (N_19913,N_19529,N_19589);
xor U19914 (N_19914,N_19635,N_19646);
and U19915 (N_19915,N_19712,N_19607);
nor U19916 (N_19916,N_19665,N_19659);
and U19917 (N_19917,N_19628,N_19555);
nand U19918 (N_19918,N_19573,N_19568);
or U19919 (N_19919,N_19657,N_19742);
nor U19920 (N_19920,N_19659,N_19586);
nor U19921 (N_19921,N_19714,N_19557);
xor U19922 (N_19922,N_19715,N_19612);
nor U19923 (N_19923,N_19590,N_19565);
and U19924 (N_19924,N_19567,N_19601);
and U19925 (N_19925,N_19668,N_19746);
xnor U19926 (N_19926,N_19520,N_19649);
or U19927 (N_19927,N_19597,N_19564);
or U19928 (N_19928,N_19520,N_19738);
and U19929 (N_19929,N_19671,N_19642);
or U19930 (N_19930,N_19671,N_19689);
nand U19931 (N_19931,N_19503,N_19628);
or U19932 (N_19932,N_19624,N_19632);
xor U19933 (N_19933,N_19702,N_19719);
nor U19934 (N_19934,N_19693,N_19697);
or U19935 (N_19935,N_19539,N_19546);
and U19936 (N_19936,N_19610,N_19737);
and U19937 (N_19937,N_19680,N_19550);
and U19938 (N_19938,N_19693,N_19631);
nor U19939 (N_19939,N_19738,N_19743);
nor U19940 (N_19940,N_19701,N_19692);
and U19941 (N_19941,N_19505,N_19519);
or U19942 (N_19942,N_19583,N_19607);
xnor U19943 (N_19943,N_19694,N_19652);
or U19944 (N_19944,N_19746,N_19736);
xor U19945 (N_19945,N_19656,N_19674);
xnor U19946 (N_19946,N_19539,N_19667);
nand U19947 (N_19947,N_19518,N_19663);
or U19948 (N_19948,N_19720,N_19530);
nor U19949 (N_19949,N_19562,N_19706);
nand U19950 (N_19950,N_19680,N_19548);
nor U19951 (N_19951,N_19644,N_19584);
or U19952 (N_19952,N_19670,N_19698);
xor U19953 (N_19953,N_19578,N_19730);
xnor U19954 (N_19954,N_19663,N_19593);
and U19955 (N_19955,N_19658,N_19675);
xnor U19956 (N_19956,N_19502,N_19575);
xor U19957 (N_19957,N_19517,N_19578);
or U19958 (N_19958,N_19725,N_19519);
nor U19959 (N_19959,N_19625,N_19720);
xnor U19960 (N_19960,N_19688,N_19661);
or U19961 (N_19961,N_19695,N_19723);
or U19962 (N_19962,N_19622,N_19715);
nor U19963 (N_19963,N_19743,N_19746);
and U19964 (N_19964,N_19525,N_19620);
or U19965 (N_19965,N_19719,N_19684);
nand U19966 (N_19966,N_19574,N_19642);
nand U19967 (N_19967,N_19558,N_19611);
xor U19968 (N_19968,N_19716,N_19673);
nor U19969 (N_19969,N_19688,N_19741);
nand U19970 (N_19970,N_19620,N_19608);
xor U19971 (N_19971,N_19642,N_19594);
nor U19972 (N_19972,N_19578,N_19589);
or U19973 (N_19973,N_19707,N_19655);
xnor U19974 (N_19974,N_19711,N_19678);
and U19975 (N_19975,N_19737,N_19658);
nand U19976 (N_19976,N_19748,N_19601);
nor U19977 (N_19977,N_19614,N_19695);
and U19978 (N_19978,N_19551,N_19602);
nand U19979 (N_19979,N_19662,N_19684);
xor U19980 (N_19980,N_19728,N_19722);
nor U19981 (N_19981,N_19545,N_19546);
or U19982 (N_19982,N_19550,N_19549);
and U19983 (N_19983,N_19675,N_19608);
xnor U19984 (N_19984,N_19627,N_19505);
and U19985 (N_19985,N_19619,N_19608);
and U19986 (N_19986,N_19688,N_19684);
nand U19987 (N_19987,N_19703,N_19559);
nand U19988 (N_19988,N_19720,N_19533);
nand U19989 (N_19989,N_19619,N_19618);
and U19990 (N_19990,N_19670,N_19561);
and U19991 (N_19991,N_19742,N_19533);
nor U19992 (N_19992,N_19702,N_19536);
nand U19993 (N_19993,N_19500,N_19630);
xor U19994 (N_19994,N_19599,N_19697);
and U19995 (N_19995,N_19534,N_19574);
or U19996 (N_19996,N_19644,N_19608);
nand U19997 (N_19997,N_19645,N_19748);
or U19998 (N_19998,N_19615,N_19653);
and U19999 (N_19999,N_19658,N_19520);
or U20000 (N_20000,N_19910,N_19946);
and U20001 (N_20001,N_19953,N_19782);
nand U20002 (N_20002,N_19951,N_19901);
xor U20003 (N_20003,N_19942,N_19772);
xnor U20004 (N_20004,N_19920,N_19918);
and U20005 (N_20005,N_19776,N_19751);
or U20006 (N_20006,N_19753,N_19868);
xor U20007 (N_20007,N_19988,N_19971);
nor U20008 (N_20008,N_19974,N_19855);
xor U20009 (N_20009,N_19997,N_19986);
xnor U20010 (N_20010,N_19876,N_19956);
nand U20011 (N_20011,N_19797,N_19885);
and U20012 (N_20012,N_19921,N_19898);
xnor U20013 (N_20013,N_19784,N_19763);
xor U20014 (N_20014,N_19820,N_19798);
and U20015 (N_20015,N_19807,N_19819);
xor U20016 (N_20016,N_19982,N_19762);
nand U20017 (N_20017,N_19856,N_19915);
or U20018 (N_20018,N_19939,N_19896);
or U20019 (N_20019,N_19874,N_19968);
nor U20020 (N_20020,N_19756,N_19919);
nand U20021 (N_20021,N_19927,N_19786);
or U20022 (N_20022,N_19995,N_19809);
or U20023 (N_20023,N_19794,N_19799);
nand U20024 (N_20024,N_19859,N_19966);
nor U20025 (N_20025,N_19835,N_19860);
nand U20026 (N_20026,N_19865,N_19911);
nor U20027 (N_20027,N_19792,N_19960);
xnor U20028 (N_20028,N_19948,N_19831);
nand U20029 (N_20029,N_19949,N_19895);
xor U20030 (N_20030,N_19830,N_19889);
xnor U20031 (N_20031,N_19916,N_19976);
xnor U20032 (N_20032,N_19992,N_19793);
and U20033 (N_20033,N_19768,N_19985);
or U20034 (N_20034,N_19935,N_19870);
nor U20035 (N_20035,N_19937,N_19929);
nor U20036 (N_20036,N_19850,N_19778);
nor U20037 (N_20037,N_19817,N_19765);
xor U20038 (N_20038,N_19975,N_19959);
nor U20039 (N_20039,N_19965,N_19833);
and U20040 (N_20040,N_19893,N_19914);
nor U20041 (N_20041,N_19752,N_19963);
nor U20042 (N_20042,N_19900,N_19908);
xnor U20043 (N_20043,N_19866,N_19806);
xnor U20044 (N_20044,N_19987,N_19924);
and U20045 (N_20045,N_19892,N_19769);
and U20046 (N_20046,N_19888,N_19801);
or U20047 (N_20047,N_19872,N_19891);
and U20048 (N_20048,N_19750,N_19867);
xnor U20049 (N_20049,N_19770,N_19862);
nor U20050 (N_20050,N_19869,N_19774);
and U20051 (N_20051,N_19757,N_19854);
and U20052 (N_20052,N_19979,N_19955);
nor U20053 (N_20053,N_19931,N_19962);
or U20054 (N_20054,N_19899,N_19790);
nand U20055 (N_20055,N_19954,N_19771);
nor U20056 (N_20056,N_19863,N_19878);
xor U20057 (N_20057,N_19947,N_19759);
or U20058 (N_20058,N_19787,N_19805);
and U20059 (N_20059,N_19941,N_19844);
and U20060 (N_20060,N_19904,N_19936);
or U20061 (N_20061,N_19788,N_19902);
xnor U20062 (N_20062,N_19907,N_19764);
and U20063 (N_20063,N_19812,N_19883);
xor U20064 (N_20064,N_19897,N_19922);
nand U20065 (N_20065,N_19810,N_19823);
xnor U20066 (N_20066,N_19950,N_19849);
nor U20067 (N_20067,N_19932,N_19933);
and U20068 (N_20068,N_19884,N_19803);
or U20069 (N_20069,N_19852,N_19754);
nor U20070 (N_20070,N_19943,N_19843);
nor U20071 (N_20071,N_19795,N_19917);
nand U20072 (N_20072,N_19926,N_19800);
xor U20073 (N_20073,N_19930,N_19773);
or U20074 (N_20074,N_19813,N_19821);
or U20075 (N_20075,N_19845,N_19758);
nor U20076 (N_20076,N_19964,N_19822);
xor U20077 (N_20077,N_19994,N_19816);
nand U20078 (N_20078,N_19938,N_19814);
nor U20079 (N_20079,N_19837,N_19829);
xnor U20080 (N_20080,N_19970,N_19909);
nand U20081 (N_20081,N_19973,N_19815);
xnor U20082 (N_20082,N_19846,N_19825);
xor U20083 (N_20083,N_19832,N_19905);
nor U20084 (N_20084,N_19875,N_19818);
xor U20085 (N_20085,N_19796,N_19811);
or U20086 (N_20086,N_19828,N_19989);
nor U20087 (N_20087,N_19839,N_19779);
nor U20088 (N_20088,N_19977,N_19802);
xor U20089 (N_20089,N_19777,N_19840);
xnor U20090 (N_20090,N_19780,N_19957);
nor U20091 (N_20091,N_19967,N_19804);
or U20092 (N_20092,N_19767,N_19836);
and U20093 (N_20093,N_19827,N_19912);
and U20094 (N_20094,N_19894,N_19789);
xnor U20095 (N_20095,N_19934,N_19785);
xor U20096 (N_20096,N_19838,N_19991);
nand U20097 (N_20097,N_19945,N_19961);
xor U20098 (N_20098,N_19873,N_19858);
xor U20099 (N_20099,N_19990,N_19940);
or U20100 (N_20100,N_19928,N_19944);
nand U20101 (N_20101,N_19996,N_19906);
and U20102 (N_20102,N_19766,N_19978);
nor U20103 (N_20103,N_19903,N_19882);
and U20104 (N_20104,N_19984,N_19877);
and U20105 (N_20105,N_19972,N_19923);
nand U20106 (N_20106,N_19983,N_19755);
nand U20107 (N_20107,N_19881,N_19969);
nor U20108 (N_20108,N_19880,N_19781);
or U20109 (N_20109,N_19841,N_19853);
xor U20110 (N_20110,N_19993,N_19775);
nand U20111 (N_20111,N_19886,N_19760);
nand U20112 (N_20112,N_19887,N_19980);
nand U20113 (N_20113,N_19999,N_19871);
xor U20114 (N_20114,N_19834,N_19958);
and U20115 (N_20115,N_19826,N_19879);
xor U20116 (N_20116,N_19981,N_19808);
nand U20117 (N_20117,N_19861,N_19848);
or U20118 (N_20118,N_19864,N_19761);
and U20119 (N_20119,N_19998,N_19913);
or U20120 (N_20120,N_19857,N_19925);
and U20121 (N_20121,N_19890,N_19847);
nand U20122 (N_20122,N_19791,N_19842);
nand U20123 (N_20123,N_19952,N_19783);
xnor U20124 (N_20124,N_19824,N_19851);
nand U20125 (N_20125,N_19808,N_19876);
or U20126 (N_20126,N_19979,N_19915);
nor U20127 (N_20127,N_19761,N_19959);
nor U20128 (N_20128,N_19990,N_19839);
nor U20129 (N_20129,N_19805,N_19982);
and U20130 (N_20130,N_19874,N_19985);
nor U20131 (N_20131,N_19958,N_19838);
nor U20132 (N_20132,N_19875,N_19956);
or U20133 (N_20133,N_19983,N_19861);
or U20134 (N_20134,N_19915,N_19872);
nand U20135 (N_20135,N_19998,N_19895);
nor U20136 (N_20136,N_19967,N_19968);
nor U20137 (N_20137,N_19819,N_19814);
nor U20138 (N_20138,N_19918,N_19963);
xor U20139 (N_20139,N_19794,N_19783);
nor U20140 (N_20140,N_19896,N_19816);
nor U20141 (N_20141,N_19937,N_19838);
and U20142 (N_20142,N_19958,N_19770);
and U20143 (N_20143,N_19903,N_19928);
and U20144 (N_20144,N_19828,N_19926);
or U20145 (N_20145,N_19950,N_19798);
or U20146 (N_20146,N_19865,N_19791);
nor U20147 (N_20147,N_19982,N_19782);
nand U20148 (N_20148,N_19972,N_19964);
nand U20149 (N_20149,N_19913,N_19981);
nand U20150 (N_20150,N_19800,N_19948);
and U20151 (N_20151,N_19813,N_19898);
nor U20152 (N_20152,N_19983,N_19790);
xnor U20153 (N_20153,N_19858,N_19915);
nand U20154 (N_20154,N_19771,N_19832);
xnor U20155 (N_20155,N_19831,N_19921);
and U20156 (N_20156,N_19987,N_19871);
or U20157 (N_20157,N_19861,N_19934);
or U20158 (N_20158,N_19805,N_19925);
and U20159 (N_20159,N_19866,N_19776);
and U20160 (N_20160,N_19843,N_19967);
nor U20161 (N_20161,N_19793,N_19781);
or U20162 (N_20162,N_19834,N_19897);
and U20163 (N_20163,N_19986,N_19964);
or U20164 (N_20164,N_19792,N_19788);
and U20165 (N_20165,N_19834,N_19823);
or U20166 (N_20166,N_19794,N_19931);
and U20167 (N_20167,N_19780,N_19799);
and U20168 (N_20168,N_19879,N_19988);
xor U20169 (N_20169,N_19811,N_19877);
nor U20170 (N_20170,N_19941,N_19957);
nand U20171 (N_20171,N_19893,N_19909);
or U20172 (N_20172,N_19984,N_19958);
nand U20173 (N_20173,N_19832,N_19995);
nand U20174 (N_20174,N_19873,N_19886);
or U20175 (N_20175,N_19940,N_19977);
nand U20176 (N_20176,N_19983,N_19854);
and U20177 (N_20177,N_19776,N_19790);
xor U20178 (N_20178,N_19816,N_19938);
nand U20179 (N_20179,N_19829,N_19853);
nor U20180 (N_20180,N_19848,N_19850);
nand U20181 (N_20181,N_19793,N_19797);
nor U20182 (N_20182,N_19893,N_19864);
xnor U20183 (N_20183,N_19850,N_19810);
nand U20184 (N_20184,N_19969,N_19901);
nor U20185 (N_20185,N_19938,N_19986);
nand U20186 (N_20186,N_19763,N_19975);
xor U20187 (N_20187,N_19807,N_19861);
and U20188 (N_20188,N_19840,N_19829);
nor U20189 (N_20189,N_19875,N_19946);
xor U20190 (N_20190,N_19855,N_19750);
nor U20191 (N_20191,N_19934,N_19873);
and U20192 (N_20192,N_19960,N_19922);
nand U20193 (N_20193,N_19766,N_19861);
or U20194 (N_20194,N_19921,N_19758);
and U20195 (N_20195,N_19957,N_19820);
nor U20196 (N_20196,N_19778,N_19799);
xor U20197 (N_20197,N_19968,N_19917);
or U20198 (N_20198,N_19957,N_19811);
xor U20199 (N_20199,N_19952,N_19962);
or U20200 (N_20200,N_19882,N_19956);
nand U20201 (N_20201,N_19960,N_19994);
nand U20202 (N_20202,N_19775,N_19958);
nor U20203 (N_20203,N_19916,N_19769);
nand U20204 (N_20204,N_19957,N_19911);
nor U20205 (N_20205,N_19962,N_19763);
nor U20206 (N_20206,N_19991,N_19872);
nor U20207 (N_20207,N_19794,N_19997);
nor U20208 (N_20208,N_19909,N_19758);
xor U20209 (N_20209,N_19825,N_19969);
nor U20210 (N_20210,N_19828,N_19767);
nor U20211 (N_20211,N_19988,N_19872);
nand U20212 (N_20212,N_19830,N_19805);
nor U20213 (N_20213,N_19908,N_19752);
xor U20214 (N_20214,N_19852,N_19944);
and U20215 (N_20215,N_19787,N_19937);
nand U20216 (N_20216,N_19914,N_19836);
xnor U20217 (N_20217,N_19907,N_19825);
and U20218 (N_20218,N_19951,N_19787);
nand U20219 (N_20219,N_19785,N_19956);
xnor U20220 (N_20220,N_19895,N_19855);
xor U20221 (N_20221,N_19939,N_19836);
xnor U20222 (N_20222,N_19840,N_19894);
xor U20223 (N_20223,N_19962,N_19904);
nand U20224 (N_20224,N_19953,N_19907);
nor U20225 (N_20225,N_19783,N_19863);
and U20226 (N_20226,N_19942,N_19965);
nor U20227 (N_20227,N_19993,N_19776);
and U20228 (N_20228,N_19782,N_19969);
nor U20229 (N_20229,N_19851,N_19947);
nor U20230 (N_20230,N_19956,N_19816);
nor U20231 (N_20231,N_19819,N_19804);
xnor U20232 (N_20232,N_19772,N_19886);
xor U20233 (N_20233,N_19763,N_19843);
or U20234 (N_20234,N_19760,N_19808);
nor U20235 (N_20235,N_19938,N_19889);
nand U20236 (N_20236,N_19812,N_19898);
xor U20237 (N_20237,N_19916,N_19911);
and U20238 (N_20238,N_19872,N_19936);
xor U20239 (N_20239,N_19883,N_19979);
and U20240 (N_20240,N_19835,N_19911);
xnor U20241 (N_20241,N_19824,N_19911);
nand U20242 (N_20242,N_19883,N_19835);
or U20243 (N_20243,N_19893,N_19940);
nor U20244 (N_20244,N_19911,N_19904);
and U20245 (N_20245,N_19883,N_19818);
nor U20246 (N_20246,N_19995,N_19906);
nor U20247 (N_20247,N_19925,N_19882);
nor U20248 (N_20248,N_19951,N_19805);
or U20249 (N_20249,N_19834,N_19843);
or U20250 (N_20250,N_20054,N_20080);
xnor U20251 (N_20251,N_20189,N_20225);
xnor U20252 (N_20252,N_20118,N_20223);
nor U20253 (N_20253,N_20240,N_20127);
nor U20254 (N_20254,N_20132,N_20072);
nor U20255 (N_20255,N_20006,N_20136);
xnor U20256 (N_20256,N_20156,N_20044);
or U20257 (N_20257,N_20096,N_20163);
nand U20258 (N_20258,N_20191,N_20074);
and U20259 (N_20259,N_20018,N_20177);
nor U20260 (N_20260,N_20023,N_20190);
xnor U20261 (N_20261,N_20192,N_20017);
nor U20262 (N_20262,N_20233,N_20198);
and U20263 (N_20263,N_20232,N_20085);
or U20264 (N_20264,N_20236,N_20048);
or U20265 (N_20265,N_20068,N_20115);
nand U20266 (N_20266,N_20143,N_20094);
or U20267 (N_20267,N_20126,N_20152);
nand U20268 (N_20268,N_20078,N_20123);
nand U20269 (N_20269,N_20102,N_20100);
nor U20270 (N_20270,N_20183,N_20065);
or U20271 (N_20271,N_20105,N_20134);
and U20272 (N_20272,N_20237,N_20180);
or U20273 (N_20273,N_20151,N_20057);
xnor U20274 (N_20274,N_20184,N_20154);
or U20275 (N_20275,N_20182,N_20224);
and U20276 (N_20276,N_20167,N_20093);
nand U20277 (N_20277,N_20090,N_20222);
xor U20278 (N_20278,N_20187,N_20249);
nand U20279 (N_20279,N_20168,N_20142);
nor U20280 (N_20280,N_20076,N_20112);
xnor U20281 (N_20281,N_20086,N_20051);
and U20282 (N_20282,N_20034,N_20084);
and U20283 (N_20283,N_20011,N_20208);
xor U20284 (N_20284,N_20111,N_20002);
xor U20285 (N_20285,N_20211,N_20235);
nand U20286 (N_20286,N_20049,N_20073);
or U20287 (N_20287,N_20212,N_20238);
xnor U20288 (N_20288,N_20241,N_20037);
xor U20289 (N_20289,N_20228,N_20114);
and U20290 (N_20290,N_20159,N_20164);
nand U20291 (N_20291,N_20138,N_20032);
and U20292 (N_20292,N_20234,N_20201);
and U20293 (N_20293,N_20013,N_20063);
or U20294 (N_20294,N_20128,N_20082);
or U20295 (N_20295,N_20216,N_20244);
and U20296 (N_20296,N_20066,N_20178);
or U20297 (N_20297,N_20103,N_20033);
nor U20298 (N_20298,N_20088,N_20108);
nor U20299 (N_20299,N_20052,N_20195);
or U20300 (N_20300,N_20171,N_20021);
nor U20301 (N_20301,N_20055,N_20141);
or U20302 (N_20302,N_20121,N_20247);
and U20303 (N_20303,N_20144,N_20149);
nor U20304 (N_20304,N_20014,N_20019);
nor U20305 (N_20305,N_20220,N_20071);
nand U20306 (N_20306,N_20194,N_20101);
nor U20307 (N_20307,N_20147,N_20119);
and U20308 (N_20308,N_20010,N_20125);
xor U20309 (N_20309,N_20122,N_20165);
nor U20310 (N_20310,N_20004,N_20039);
nor U20311 (N_20311,N_20209,N_20137);
or U20312 (N_20312,N_20210,N_20131);
or U20313 (N_20313,N_20193,N_20031);
nor U20314 (N_20314,N_20218,N_20040);
xnor U20315 (N_20315,N_20060,N_20020);
nor U20316 (N_20316,N_20116,N_20160);
or U20317 (N_20317,N_20075,N_20045);
and U20318 (N_20318,N_20161,N_20000);
and U20319 (N_20319,N_20242,N_20214);
or U20320 (N_20320,N_20181,N_20081);
or U20321 (N_20321,N_20083,N_20230);
nor U20322 (N_20322,N_20202,N_20092);
xnor U20323 (N_20323,N_20203,N_20206);
nor U20324 (N_20324,N_20221,N_20227);
nand U20325 (N_20325,N_20009,N_20117);
or U20326 (N_20326,N_20246,N_20248);
nand U20327 (N_20327,N_20162,N_20124);
or U20328 (N_20328,N_20153,N_20174);
xor U20329 (N_20329,N_20135,N_20204);
nor U20330 (N_20330,N_20215,N_20155);
nand U20331 (N_20331,N_20070,N_20058);
nor U20332 (N_20332,N_20219,N_20012);
nand U20333 (N_20333,N_20139,N_20028);
xnor U20334 (N_20334,N_20179,N_20091);
or U20335 (N_20335,N_20196,N_20133);
nand U20336 (N_20336,N_20150,N_20003);
xor U20337 (N_20337,N_20038,N_20186);
or U20338 (N_20338,N_20166,N_20226);
and U20339 (N_20339,N_20169,N_20113);
xnor U20340 (N_20340,N_20175,N_20176);
or U20341 (N_20341,N_20024,N_20005);
and U20342 (N_20342,N_20107,N_20173);
nand U20343 (N_20343,N_20036,N_20061);
nand U20344 (N_20344,N_20095,N_20030);
xnor U20345 (N_20345,N_20087,N_20199);
nor U20346 (N_20346,N_20059,N_20170);
or U20347 (N_20347,N_20213,N_20110);
xor U20348 (N_20348,N_20229,N_20062);
and U20349 (N_20349,N_20231,N_20245);
or U20350 (N_20350,N_20043,N_20200);
nor U20351 (N_20351,N_20007,N_20148);
nand U20352 (N_20352,N_20064,N_20146);
and U20353 (N_20353,N_20129,N_20205);
and U20354 (N_20354,N_20207,N_20077);
nand U20355 (N_20355,N_20140,N_20053);
or U20356 (N_20356,N_20022,N_20098);
or U20357 (N_20357,N_20188,N_20050);
nand U20358 (N_20358,N_20041,N_20217);
or U20359 (N_20359,N_20026,N_20015);
nor U20360 (N_20360,N_20158,N_20239);
nor U20361 (N_20361,N_20197,N_20069);
nor U20362 (N_20362,N_20097,N_20016);
nor U20363 (N_20363,N_20172,N_20008);
nor U20364 (N_20364,N_20046,N_20145);
nor U20365 (N_20365,N_20157,N_20001);
xnor U20366 (N_20366,N_20035,N_20243);
and U20367 (N_20367,N_20025,N_20042);
nor U20368 (N_20368,N_20106,N_20047);
xnor U20369 (N_20369,N_20099,N_20067);
or U20370 (N_20370,N_20056,N_20029);
and U20371 (N_20371,N_20079,N_20089);
xor U20372 (N_20372,N_20130,N_20109);
and U20373 (N_20373,N_20185,N_20120);
nor U20374 (N_20374,N_20027,N_20104);
nand U20375 (N_20375,N_20000,N_20167);
nor U20376 (N_20376,N_20087,N_20084);
or U20377 (N_20377,N_20131,N_20018);
or U20378 (N_20378,N_20236,N_20223);
and U20379 (N_20379,N_20127,N_20139);
or U20380 (N_20380,N_20232,N_20172);
xnor U20381 (N_20381,N_20141,N_20023);
nand U20382 (N_20382,N_20245,N_20000);
or U20383 (N_20383,N_20193,N_20021);
and U20384 (N_20384,N_20234,N_20143);
and U20385 (N_20385,N_20147,N_20108);
nor U20386 (N_20386,N_20205,N_20092);
nand U20387 (N_20387,N_20155,N_20009);
or U20388 (N_20388,N_20166,N_20113);
xor U20389 (N_20389,N_20153,N_20188);
nand U20390 (N_20390,N_20072,N_20189);
xnor U20391 (N_20391,N_20023,N_20085);
nand U20392 (N_20392,N_20166,N_20053);
xnor U20393 (N_20393,N_20019,N_20189);
or U20394 (N_20394,N_20167,N_20015);
nor U20395 (N_20395,N_20200,N_20233);
and U20396 (N_20396,N_20029,N_20197);
and U20397 (N_20397,N_20090,N_20168);
nor U20398 (N_20398,N_20190,N_20223);
xor U20399 (N_20399,N_20083,N_20032);
and U20400 (N_20400,N_20097,N_20012);
xnor U20401 (N_20401,N_20011,N_20239);
nand U20402 (N_20402,N_20105,N_20049);
nor U20403 (N_20403,N_20016,N_20156);
nand U20404 (N_20404,N_20142,N_20123);
xor U20405 (N_20405,N_20116,N_20123);
nand U20406 (N_20406,N_20191,N_20221);
nand U20407 (N_20407,N_20125,N_20128);
and U20408 (N_20408,N_20159,N_20193);
xor U20409 (N_20409,N_20029,N_20173);
nand U20410 (N_20410,N_20022,N_20032);
and U20411 (N_20411,N_20008,N_20062);
nand U20412 (N_20412,N_20126,N_20041);
or U20413 (N_20413,N_20146,N_20148);
nor U20414 (N_20414,N_20063,N_20229);
nand U20415 (N_20415,N_20144,N_20168);
and U20416 (N_20416,N_20101,N_20185);
nor U20417 (N_20417,N_20155,N_20219);
or U20418 (N_20418,N_20151,N_20031);
or U20419 (N_20419,N_20179,N_20065);
xor U20420 (N_20420,N_20222,N_20081);
and U20421 (N_20421,N_20055,N_20163);
or U20422 (N_20422,N_20173,N_20121);
or U20423 (N_20423,N_20190,N_20157);
nand U20424 (N_20424,N_20248,N_20163);
nand U20425 (N_20425,N_20007,N_20100);
and U20426 (N_20426,N_20140,N_20006);
xnor U20427 (N_20427,N_20141,N_20241);
nor U20428 (N_20428,N_20139,N_20060);
and U20429 (N_20429,N_20190,N_20109);
and U20430 (N_20430,N_20069,N_20218);
and U20431 (N_20431,N_20166,N_20051);
or U20432 (N_20432,N_20005,N_20082);
nand U20433 (N_20433,N_20188,N_20045);
and U20434 (N_20434,N_20022,N_20024);
nor U20435 (N_20435,N_20211,N_20099);
nor U20436 (N_20436,N_20204,N_20178);
or U20437 (N_20437,N_20182,N_20069);
xnor U20438 (N_20438,N_20169,N_20055);
nor U20439 (N_20439,N_20026,N_20208);
xor U20440 (N_20440,N_20153,N_20223);
nand U20441 (N_20441,N_20197,N_20195);
nor U20442 (N_20442,N_20181,N_20248);
nand U20443 (N_20443,N_20182,N_20053);
and U20444 (N_20444,N_20173,N_20082);
xor U20445 (N_20445,N_20143,N_20100);
nor U20446 (N_20446,N_20038,N_20002);
nor U20447 (N_20447,N_20094,N_20133);
nand U20448 (N_20448,N_20049,N_20084);
nor U20449 (N_20449,N_20045,N_20094);
or U20450 (N_20450,N_20014,N_20087);
or U20451 (N_20451,N_20183,N_20071);
and U20452 (N_20452,N_20157,N_20002);
xor U20453 (N_20453,N_20091,N_20075);
nor U20454 (N_20454,N_20178,N_20117);
xor U20455 (N_20455,N_20049,N_20125);
xnor U20456 (N_20456,N_20026,N_20012);
or U20457 (N_20457,N_20206,N_20025);
and U20458 (N_20458,N_20149,N_20030);
or U20459 (N_20459,N_20152,N_20073);
or U20460 (N_20460,N_20218,N_20077);
or U20461 (N_20461,N_20075,N_20227);
nand U20462 (N_20462,N_20171,N_20158);
and U20463 (N_20463,N_20116,N_20119);
and U20464 (N_20464,N_20052,N_20113);
xor U20465 (N_20465,N_20009,N_20151);
or U20466 (N_20466,N_20111,N_20110);
and U20467 (N_20467,N_20097,N_20223);
nor U20468 (N_20468,N_20143,N_20187);
xor U20469 (N_20469,N_20236,N_20138);
or U20470 (N_20470,N_20168,N_20031);
and U20471 (N_20471,N_20074,N_20085);
xor U20472 (N_20472,N_20004,N_20098);
nor U20473 (N_20473,N_20033,N_20154);
and U20474 (N_20474,N_20134,N_20109);
nand U20475 (N_20475,N_20192,N_20095);
xnor U20476 (N_20476,N_20248,N_20187);
xor U20477 (N_20477,N_20144,N_20096);
and U20478 (N_20478,N_20124,N_20029);
xnor U20479 (N_20479,N_20219,N_20218);
nand U20480 (N_20480,N_20154,N_20208);
and U20481 (N_20481,N_20135,N_20101);
and U20482 (N_20482,N_20132,N_20081);
and U20483 (N_20483,N_20170,N_20163);
nand U20484 (N_20484,N_20086,N_20220);
xor U20485 (N_20485,N_20193,N_20180);
nand U20486 (N_20486,N_20172,N_20160);
nand U20487 (N_20487,N_20059,N_20029);
nand U20488 (N_20488,N_20122,N_20034);
and U20489 (N_20489,N_20199,N_20095);
nand U20490 (N_20490,N_20093,N_20132);
xnor U20491 (N_20491,N_20100,N_20192);
nor U20492 (N_20492,N_20109,N_20125);
and U20493 (N_20493,N_20088,N_20146);
or U20494 (N_20494,N_20147,N_20092);
xnor U20495 (N_20495,N_20144,N_20070);
and U20496 (N_20496,N_20088,N_20042);
nor U20497 (N_20497,N_20095,N_20166);
or U20498 (N_20498,N_20001,N_20160);
nand U20499 (N_20499,N_20247,N_20210);
nand U20500 (N_20500,N_20435,N_20283);
xor U20501 (N_20501,N_20358,N_20337);
or U20502 (N_20502,N_20257,N_20412);
or U20503 (N_20503,N_20372,N_20431);
nand U20504 (N_20504,N_20485,N_20270);
xnor U20505 (N_20505,N_20459,N_20310);
nand U20506 (N_20506,N_20286,N_20299);
nand U20507 (N_20507,N_20439,N_20492);
nor U20508 (N_20508,N_20329,N_20254);
nand U20509 (N_20509,N_20292,N_20368);
or U20510 (N_20510,N_20256,N_20405);
xnor U20511 (N_20511,N_20441,N_20496);
nor U20512 (N_20512,N_20415,N_20376);
or U20513 (N_20513,N_20274,N_20339);
xnor U20514 (N_20514,N_20378,N_20456);
nor U20515 (N_20515,N_20262,N_20269);
nor U20516 (N_20516,N_20467,N_20389);
xnor U20517 (N_20517,N_20335,N_20319);
nand U20518 (N_20518,N_20450,N_20290);
and U20519 (N_20519,N_20324,N_20287);
and U20520 (N_20520,N_20325,N_20273);
or U20521 (N_20521,N_20359,N_20394);
nor U20522 (N_20522,N_20499,N_20308);
and U20523 (N_20523,N_20313,N_20336);
xnor U20524 (N_20524,N_20426,N_20333);
nand U20525 (N_20525,N_20408,N_20309);
nand U20526 (N_20526,N_20354,N_20442);
nand U20527 (N_20527,N_20478,N_20425);
nand U20528 (N_20528,N_20327,N_20486);
nand U20529 (N_20529,N_20440,N_20414);
nor U20530 (N_20530,N_20422,N_20464);
or U20531 (N_20531,N_20390,N_20465);
or U20532 (N_20532,N_20413,N_20330);
and U20533 (N_20533,N_20312,N_20480);
xor U20534 (N_20534,N_20409,N_20321);
or U20535 (N_20535,N_20391,N_20475);
nor U20536 (N_20536,N_20481,N_20424);
xnor U20537 (N_20537,N_20331,N_20407);
nand U20538 (N_20538,N_20288,N_20268);
nor U20539 (N_20539,N_20373,N_20362);
nand U20540 (N_20540,N_20356,N_20258);
or U20541 (N_20541,N_20493,N_20393);
nand U20542 (N_20542,N_20430,N_20265);
nor U20543 (N_20543,N_20350,N_20472);
or U20544 (N_20544,N_20474,N_20494);
nand U20545 (N_20545,N_20479,N_20326);
nor U20546 (N_20546,N_20346,N_20498);
nand U20547 (N_20547,N_20317,N_20296);
nand U20548 (N_20548,N_20315,N_20451);
and U20549 (N_20549,N_20427,N_20490);
and U20550 (N_20550,N_20416,N_20434);
or U20551 (N_20551,N_20260,N_20297);
nor U20552 (N_20552,N_20251,N_20374);
and U20553 (N_20553,N_20419,N_20381);
xor U20554 (N_20554,N_20495,N_20322);
nand U20555 (N_20555,N_20455,N_20385);
xor U20556 (N_20556,N_20259,N_20444);
nor U20557 (N_20557,N_20396,N_20436);
nor U20558 (N_20558,N_20355,N_20382);
and U20559 (N_20559,N_20250,N_20402);
or U20560 (N_20560,N_20328,N_20448);
nor U20561 (N_20561,N_20305,N_20369);
xor U20562 (N_20562,N_20300,N_20388);
or U20563 (N_20563,N_20302,N_20418);
or U20564 (N_20564,N_20437,N_20314);
and U20565 (N_20565,N_20417,N_20266);
nor U20566 (N_20566,N_20468,N_20357);
xnor U20567 (N_20567,N_20410,N_20399);
nand U20568 (N_20568,N_20352,N_20483);
or U20569 (N_20569,N_20397,N_20395);
and U20570 (N_20570,N_20349,N_20348);
nand U20571 (N_20571,N_20429,N_20370);
xor U20572 (N_20572,N_20353,N_20401);
or U20573 (N_20573,N_20384,N_20295);
or U20574 (N_20574,N_20311,N_20364);
or U20575 (N_20575,N_20281,N_20360);
or U20576 (N_20576,N_20351,N_20289);
or U20577 (N_20577,N_20361,N_20303);
xor U20578 (N_20578,N_20406,N_20377);
nor U20579 (N_20579,N_20386,N_20363);
and U20580 (N_20580,N_20298,N_20340);
nand U20581 (N_20581,N_20477,N_20301);
or U20582 (N_20582,N_20253,N_20423);
nand U20583 (N_20583,N_20445,N_20271);
xnor U20584 (N_20584,N_20411,N_20497);
xor U20585 (N_20585,N_20291,N_20264);
xor U20586 (N_20586,N_20476,N_20438);
or U20587 (N_20587,N_20279,N_20285);
nor U20588 (N_20588,N_20306,N_20458);
nor U20589 (N_20589,N_20400,N_20371);
nor U20590 (N_20590,N_20383,N_20433);
and U20591 (N_20591,N_20294,N_20462);
nor U20592 (N_20592,N_20420,N_20443);
and U20593 (N_20593,N_20454,N_20267);
nand U20594 (N_20594,N_20275,N_20482);
xnor U20595 (N_20595,N_20380,N_20449);
nor U20596 (N_20596,N_20345,N_20404);
nor U20597 (N_20597,N_20334,N_20466);
nor U20598 (N_20598,N_20323,N_20446);
nand U20599 (N_20599,N_20280,N_20491);
nand U20600 (N_20600,N_20365,N_20471);
and U20601 (N_20601,N_20447,N_20341);
nand U20602 (N_20602,N_20284,N_20282);
nand U20603 (N_20603,N_20367,N_20320);
xor U20604 (N_20604,N_20375,N_20421);
nor U20605 (N_20605,N_20484,N_20488);
and U20606 (N_20606,N_20392,N_20278);
or U20607 (N_20607,N_20343,N_20255);
nand U20608 (N_20608,N_20304,N_20261);
nor U20609 (N_20609,N_20463,N_20428);
nand U20610 (N_20610,N_20460,N_20489);
and U20611 (N_20611,N_20252,N_20316);
and U20612 (N_20612,N_20276,N_20453);
and U20613 (N_20613,N_20379,N_20403);
nand U20614 (N_20614,N_20432,N_20293);
and U20615 (N_20615,N_20338,N_20452);
xor U20616 (N_20616,N_20461,N_20470);
or U20617 (N_20617,N_20277,N_20473);
nand U20618 (N_20618,N_20342,N_20272);
or U20619 (N_20619,N_20387,N_20347);
and U20620 (N_20620,N_20307,N_20344);
nand U20621 (N_20621,N_20487,N_20318);
nand U20622 (N_20622,N_20457,N_20398);
and U20623 (N_20623,N_20332,N_20366);
nor U20624 (N_20624,N_20469,N_20263);
nor U20625 (N_20625,N_20333,N_20267);
xnor U20626 (N_20626,N_20269,N_20487);
nand U20627 (N_20627,N_20434,N_20311);
or U20628 (N_20628,N_20338,N_20482);
nor U20629 (N_20629,N_20268,N_20417);
xnor U20630 (N_20630,N_20253,N_20254);
and U20631 (N_20631,N_20471,N_20366);
nand U20632 (N_20632,N_20380,N_20420);
xnor U20633 (N_20633,N_20409,N_20474);
and U20634 (N_20634,N_20324,N_20438);
nor U20635 (N_20635,N_20318,N_20372);
nor U20636 (N_20636,N_20410,N_20420);
nor U20637 (N_20637,N_20452,N_20285);
xor U20638 (N_20638,N_20285,N_20333);
nor U20639 (N_20639,N_20274,N_20314);
nand U20640 (N_20640,N_20426,N_20303);
nand U20641 (N_20641,N_20334,N_20271);
and U20642 (N_20642,N_20282,N_20373);
or U20643 (N_20643,N_20341,N_20283);
xnor U20644 (N_20644,N_20462,N_20490);
nand U20645 (N_20645,N_20366,N_20306);
and U20646 (N_20646,N_20257,N_20414);
and U20647 (N_20647,N_20279,N_20415);
xnor U20648 (N_20648,N_20292,N_20360);
or U20649 (N_20649,N_20286,N_20359);
nand U20650 (N_20650,N_20289,N_20314);
nand U20651 (N_20651,N_20475,N_20345);
nor U20652 (N_20652,N_20286,N_20450);
and U20653 (N_20653,N_20382,N_20363);
nor U20654 (N_20654,N_20339,N_20467);
nand U20655 (N_20655,N_20269,N_20439);
xor U20656 (N_20656,N_20367,N_20433);
nor U20657 (N_20657,N_20271,N_20280);
nand U20658 (N_20658,N_20412,N_20278);
xnor U20659 (N_20659,N_20351,N_20369);
xor U20660 (N_20660,N_20450,N_20358);
xnor U20661 (N_20661,N_20390,N_20250);
and U20662 (N_20662,N_20421,N_20276);
xnor U20663 (N_20663,N_20487,N_20310);
or U20664 (N_20664,N_20300,N_20390);
and U20665 (N_20665,N_20288,N_20475);
and U20666 (N_20666,N_20436,N_20391);
xnor U20667 (N_20667,N_20483,N_20389);
or U20668 (N_20668,N_20432,N_20386);
xor U20669 (N_20669,N_20408,N_20478);
xor U20670 (N_20670,N_20250,N_20400);
and U20671 (N_20671,N_20450,N_20257);
or U20672 (N_20672,N_20483,N_20361);
nand U20673 (N_20673,N_20261,N_20328);
nor U20674 (N_20674,N_20406,N_20473);
or U20675 (N_20675,N_20481,N_20297);
nand U20676 (N_20676,N_20414,N_20332);
and U20677 (N_20677,N_20273,N_20478);
xor U20678 (N_20678,N_20441,N_20339);
xor U20679 (N_20679,N_20280,N_20355);
and U20680 (N_20680,N_20298,N_20474);
and U20681 (N_20681,N_20274,N_20342);
xor U20682 (N_20682,N_20298,N_20251);
or U20683 (N_20683,N_20331,N_20486);
or U20684 (N_20684,N_20391,N_20292);
nor U20685 (N_20685,N_20262,N_20312);
nand U20686 (N_20686,N_20474,N_20472);
xnor U20687 (N_20687,N_20289,N_20283);
and U20688 (N_20688,N_20429,N_20361);
and U20689 (N_20689,N_20313,N_20474);
or U20690 (N_20690,N_20397,N_20434);
nor U20691 (N_20691,N_20332,N_20322);
xnor U20692 (N_20692,N_20348,N_20311);
nand U20693 (N_20693,N_20487,N_20452);
nand U20694 (N_20694,N_20453,N_20384);
xnor U20695 (N_20695,N_20318,N_20350);
nand U20696 (N_20696,N_20385,N_20336);
nand U20697 (N_20697,N_20359,N_20448);
and U20698 (N_20698,N_20342,N_20456);
xnor U20699 (N_20699,N_20471,N_20459);
nor U20700 (N_20700,N_20485,N_20454);
nor U20701 (N_20701,N_20416,N_20459);
and U20702 (N_20702,N_20314,N_20284);
or U20703 (N_20703,N_20295,N_20367);
nand U20704 (N_20704,N_20275,N_20343);
nand U20705 (N_20705,N_20405,N_20400);
nor U20706 (N_20706,N_20488,N_20368);
xnor U20707 (N_20707,N_20463,N_20308);
and U20708 (N_20708,N_20468,N_20297);
xnor U20709 (N_20709,N_20383,N_20265);
nor U20710 (N_20710,N_20307,N_20276);
nand U20711 (N_20711,N_20480,N_20332);
or U20712 (N_20712,N_20386,N_20444);
nand U20713 (N_20713,N_20437,N_20477);
nand U20714 (N_20714,N_20362,N_20383);
nor U20715 (N_20715,N_20349,N_20369);
nand U20716 (N_20716,N_20283,N_20377);
nand U20717 (N_20717,N_20468,N_20395);
xnor U20718 (N_20718,N_20451,N_20489);
nor U20719 (N_20719,N_20370,N_20492);
nor U20720 (N_20720,N_20340,N_20457);
and U20721 (N_20721,N_20345,N_20368);
and U20722 (N_20722,N_20458,N_20307);
or U20723 (N_20723,N_20297,N_20368);
nor U20724 (N_20724,N_20350,N_20477);
and U20725 (N_20725,N_20353,N_20481);
or U20726 (N_20726,N_20350,N_20288);
and U20727 (N_20727,N_20382,N_20468);
or U20728 (N_20728,N_20437,N_20255);
nor U20729 (N_20729,N_20459,N_20373);
or U20730 (N_20730,N_20251,N_20315);
xnor U20731 (N_20731,N_20315,N_20279);
xnor U20732 (N_20732,N_20357,N_20424);
nor U20733 (N_20733,N_20253,N_20437);
or U20734 (N_20734,N_20420,N_20482);
nand U20735 (N_20735,N_20306,N_20475);
nand U20736 (N_20736,N_20318,N_20391);
xnor U20737 (N_20737,N_20327,N_20315);
nand U20738 (N_20738,N_20394,N_20492);
xnor U20739 (N_20739,N_20373,N_20315);
nor U20740 (N_20740,N_20472,N_20338);
xor U20741 (N_20741,N_20295,N_20403);
and U20742 (N_20742,N_20415,N_20455);
nor U20743 (N_20743,N_20444,N_20495);
or U20744 (N_20744,N_20447,N_20400);
xor U20745 (N_20745,N_20488,N_20303);
xnor U20746 (N_20746,N_20377,N_20427);
and U20747 (N_20747,N_20281,N_20459);
nand U20748 (N_20748,N_20272,N_20459);
nand U20749 (N_20749,N_20470,N_20474);
or U20750 (N_20750,N_20747,N_20694);
and U20751 (N_20751,N_20558,N_20611);
nor U20752 (N_20752,N_20743,N_20681);
or U20753 (N_20753,N_20588,N_20744);
nor U20754 (N_20754,N_20587,N_20567);
nor U20755 (N_20755,N_20622,N_20596);
and U20756 (N_20756,N_20742,N_20583);
xor U20757 (N_20757,N_20668,N_20568);
nor U20758 (N_20758,N_20693,N_20663);
and U20759 (N_20759,N_20739,N_20706);
nand U20760 (N_20760,N_20581,N_20711);
xnor U20761 (N_20761,N_20686,N_20606);
nor U20762 (N_20762,N_20505,N_20627);
nand U20763 (N_20763,N_20605,N_20514);
nand U20764 (N_20764,N_20647,N_20705);
xor U20765 (N_20765,N_20502,N_20708);
xnor U20766 (N_20766,N_20552,N_20507);
and U20767 (N_20767,N_20734,N_20538);
nor U20768 (N_20768,N_20547,N_20632);
nor U20769 (N_20769,N_20549,N_20580);
nand U20770 (N_20770,N_20698,N_20709);
or U20771 (N_20771,N_20511,N_20500);
nor U20772 (N_20772,N_20621,N_20566);
nand U20773 (N_20773,N_20603,N_20579);
xnor U20774 (N_20774,N_20569,N_20738);
nand U20775 (N_20775,N_20731,N_20717);
and U20776 (N_20776,N_20737,N_20703);
and U20777 (N_20777,N_20509,N_20609);
and U20778 (N_20778,N_20534,N_20729);
xnor U20779 (N_20779,N_20608,N_20696);
xnor U20780 (N_20780,N_20689,N_20501);
or U20781 (N_20781,N_20562,N_20630);
or U20782 (N_20782,N_20537,N_20667);
nand U20783 (N_20783,N_20676,N_20715);
and U20784 (N_20784,N_20528,N_20617);
and U20785 (N_20785,N_20659,N_20642);
nor U20786 (N_20786,N_20559,N_20556);
xnor U20787 (N_20787,N_20504,N_20526);
nor U20788 (N_20788,N_20530,N_20732);
nand U20789 (N_20789,N_20524,N_20575);
xor U20790 (N_20790,N_20513,N_20506);
or U20791 (N_20791,N_20574,N_20688);
or U20792 (N_20792,N_20702,N_20720);
xnor U20793 (N_20793,N_20607,N_20662);
or U20794 (N_20794,N_20554,N_20683);
xor U20795 (N_20795,N_20675,N_20651);
nand U20796 (N_20796,N_20664,N_20741);
and U20797 (N_20797,N_20631,N_20582);
xor U20798 (N_20798,N_20672,N_20590);
nor U20799 (N_20799,N_20724,N_20529);
or U20800 (N_20800,N_20640,N_20520);
xnor U20801 (N_20801,N_20730,N_20727);
or U20802 (N_20802,N_20592,N_20684);
nor U20803 (N_20803,N_20707,N_20602);
nor U20804 (N_20804,N_20654,N_20718);
nor U20805 (N_20805,N_20548,N_20601);
nand U20806 (N_20806,N_20637,N_20523);
or U20807 (N_20807,N_20619,N_20628);
xnor U20808 (N_20808,N_20650,N_20540);
or U20809 (N_20809,N_20570,N_20682);
xor U20810 (N_20810,N_20623,N_20551);
nand U20811 (N_20811,N_20531,N_20599);
and U20812 (N_20812,N_20745,N_20550);
nand U20813 (N_20813,N_20578,N_20669);
nor U20814 (N_20814,N_20656,N_20598);
or U20815 (N_20815,N_20740,N_20518);
nor U20816 (N_20816,N_20604,N_20503);
or U20817 (N_20817,N_20677,N_20721);
and U20818 (N_20818,N_20673,N_20577);
or U20819 (N_20819,N_20585,N_20643);
or U20820 (N_20820,N_20618,N_20616);
nand U20821 (N_20821,N_20629,N_20645);
nand U20822 (N_20822,N_20726,N_20541);
nor U20823 (N_20823,N_20660,N_20553);
nand U20824 (N_20824,N_20508,N_20639);
and U20825 (N_20825,N_20612,N_20670);
nand U20826 (N_20826,N_20536,N_20722);
or U20827 (N_20827,N_20725,N_20591);
and U20828 (N_20828,N_20748,N_20648);
nand U20829 (N_20829,N_20657,N_20594);
nor U20830 (N_20830,N_20658,N_20680);
or U20831 (N_20831,N_20512,N_20649);
nor U20832 (N_20832,N_20701,N_20564);
and U20833 (N_20833,N_20653,N_20589);
and U20834 (N_20834,N_20521,N_20713);
nand U20835 (N_20835,N_20576,N_20555);
nand U20836 (N_20836,N_20561,N_20638);
nor U20837 (N_20837,N_20544,N_20700);
nor U20838 (N_20838,N_20565,N_20735);
or U20839 (N_20839,N_20665,N_20644);
nand U20840 (N_20840,N_20515,N_20620);
nor U20841 (N_20841,N_20749,N_20595);
or U20842 (N_20842,N_20516,N_20539);
nand U20843 (N_20843,N_20733,N_20615);
nand U20844 (N_20844,N_20692,N_20557);
xor U20845 (N_20845,N_20572,N_20626);
and U20846 (N_20846,N_20691,N_20646);
xor U20847 (N_20847,N_20600,N_20679);
nor U20848 (N_20848,N_20535,N_20690);
and U20849 (N_20849,N_20712,N_20614);
or U20850 (N_20850,N_20573,N_20723);
and U20851 (N_20851,N_20695,N_20685);
xor U20852 (N_20852,N_20635,N_20678);
and U20853 (N_20853,N_20610,N_20527);
xnor U20854 (N_20854,N_20641,N_20625);
or U20855 (N_20855,N_20736,N_20699);
nand U20856 (N_20856,N_20545,N_20728);
xnor U20857 (N_20857,N_20655,N_20517);
and U20858 (N_20858,N_20746,N_20714);
nand U20859 (N_20859,N_20519,N_20697);
xnor U20860 (N_20860,N_20652,N_20563);
nor U20861 (N_20861,N_20674,N_20584);
xnor U20862 (N_20862,N_20710,N_20586);
or U20863 (N_20863,N_20634,N_20522);
nor U20864 (N_20864,N_20666,N_20533);
nand U20865 (N_20865,N_20510,N_20532);
nand U20866 (N_20866,N_20704,N_20593);
and U20867 (N_20867,N_20525,N_20543);
xor U20868 (N_20868,N_20716,N_20633);
and U20869 (N_20869,N_20687,N_20597);
and U20870 (N_20870,N_20546,N_20613);
nand U20871 (N_20871,N_20571,N_20542);
xnor U20872 (N_20872,N_20624,N_20560);
nor U20873 (N_20873,N_20719,N_20671);
nand U20874 (N_20874,N_20661,N_20636);
and U20875 (N_20875,N_20584,N_20714);
or U20876 (N_20876,N_20702,N_20738);
xnor U20877 (N_20877,N_20574,N_20585);
xor U20878 (N_20878,N_20609,N_20648);
xnor U20879 (N_20879,N_20589,N_20687);
nor U20880 (N_20880,N_20603,N_20500);
xnor U20881 (N_20881,N_20565,N_20614);
xnor U20882 (N_20882,N_20662,N_20734);
or U20883 (N_20883,N_20703,N_20701);
xor U20884 (N_20884,N_20743,N_20717);
and U20885 (N_20885,N_20592,N_20717);
nand U20886 (N_20886,N_20603,N_20614);
nand U20887 (N_20887,N_20610,N_20670);
or U20888 (N_20888,N_20511,N_20682);
xnor U20889 (N_20889,N_20665,N_20651);
xor U20890 (N_20890,N_20536,N_20729);
nor U20891 (N_20891,N_20584,N_20747);
nor U20892 (N_20892,N_20669,N_20541);
and U20893 (N_20893,N_20535,N_20521);
xor U20894 (N_20894,N_20524,N_20503);
nor U20895 (N_20895,N_20504,N_20609);
and U20896 (N_20896,N_20606,N_20523);
or U20897 (N_20897,N_20530,N_20665);
nor U20898 (N_20898,N_20506,N_20658);
and U20899 (N_20899,N_20714,N_20748);
nand U20900 (N_20900,N_20580,N_20507);
nand U20901 (N_20901,N_20603,N_20664);
nor U20902 (N_20902,N_20640,N_20589);
nor U20903 (N_20903,N_20508,N_20670);
xor U20904 (N_20904,N_20670,N_20521);
nand U20905 (N_20905,N_20626,N_20558);
nand U20906 (N_20906,N_20515,N_20638);
or U20907 (N_20907,N_20658,N_20718);
or U20908 (N_20908,N_20672,N_20697);
or U20909 (N_20909,N_20563,N_20684);
and U20910 (N_20910,N_20602,N_20646);
and U20911 (N_20911,N_20688,N_20703);
and U20912 (N_20912,N_20748,N_20659);
and U20913 (N_20913,N_20704,N_20588);
nor U20914 (N_20914,N_20746,N_20690);
and U20915 (N_20915,N_20598,N_20501);
or U20916 (N_20916,N_20618,N_20637);
nand U20917 (N_20917,N_20675,N_20687);
nor U20918 (N_20918,N_20680,N_20544);
or U20919 (N_20919,N_20572,N_20524);
xnor U20920 (N_20920,N_20721,N_20644);
xnor U20921 (N_20921,N_20676,N_20625);
nand U20922 (N_20922,N_20553,N_20749);
or U20923 (N_20923,N_20503,N_20638);
or U20924 (N_20924,N_20529,N_20524);
and U20925 (N_20925,N_20570,N_20556);
or U20926 (N_20926,N_20637,N_20679);
nor U20927 (N_20927,N_20557,N_20701);
xnor U20928 (N_20928,N_20570,N_20574);
nand U20929 (N_20929,N_20558,N_20620);
or U20930 (N_20930,N_20747,N_20660);
xor U20931 (N_20931,N_20716,N_20551);
or U20932 (N_20932,N_20720,N_20512);
and U20933 (N_20933,N_20685,N_20681);
nand U20934 (N_20934,N_20544,N_20747);
nand U20935 (N_20935,N_20675,N_20560);
xnor U20936 (N_20936,N_20562,N_20511);
nor U20937 (N_20937,N_20503,N_20679);
nor U20938 (N_20938,N_20554,N_20541);
nand U20939 (N_20939,N_20665,N_20743);
nor U20940 (N_20940,N_20557,N_20702);
nor U20941 (N_20941,N_20641,N_20601);
or U20942 (N_20942,N_20679,N_20673);
xnor U20943 (N_20943,N_20510,N_20538);
nand U20944 (N_20944,N_20685,N_20715);
and U20945 (N_20945,N_20745,N_20532);
nand U20946 (N_20946,N_20589,N_20520);
nand U20947 (N_20947,N_20686,N_20722);
xnor U20948 (N_20948,N_20644,N_20575);
nor U20949 (N_20949,N_20688,N_20738);
nor U20950 (N_20950,N_20714,N_20631);
nand U20951 (N_20951,N_20669,N_20519);
or U20952 (N_20952,N_20514,N_20714);
and U20953 (N_20953,N_20731,N_20679);
nand U20954 (N_20954,N_20508,N_20658);
xnor U20955 (N_20955,N_20668,N_20681);
nor U20956 (N_20956,N_20647,N_20662);
nor U20957 (N_20957,N_20511,N_20698);
nand U20958 (N_20958,N_20528,N_20635);
or U20959 (N_20959,N_20574,N_20609);
and U20960 (N_20960,N_20608,N_20500);
and U20961 (N_20961,N_20540,N_20504);
nand U20962 (N_20962,N_20739,N_20681);
or U20963 (N_20963,N_20613,N_20743);
nor U20964 (N_20964,N_20561,N_20715);
or U20965 (N_20965,N_20568,N_20516);
or U20966 (N_20966,N_20727,N_20560);
nor U20967 (N_20967,N_20653,N_20654);
nor U20968 (N_20968,N_20744,N_20688);
nor U20969 (N_20969,N_20507,N_20690);
or U20970 (N_20970,N_20527,N_20673);
xnor U20971 (N_20971,N_20560,N_20518);
or U20972 (N_20972,N_20593,N_20684);
xnor U20973 (N_20973,N_20695,N_20705);
xnor U20974 (N_20974,N_20725,N_20559);
xor U20975 (N_20975,N_20668,N_20505);
or U20976 (N_20976,N_20728,N_20568);
nor U20977 (N_20977,N_20641,N_20619);
and U20978 (N_20978,N_20672,N_20748);
xnor U20979 (N_20979,N_20723,N_20724);
xor U20980 (N_20980,N_20560,N_20660);
nor U20981 (N_20981,N_20536,N_20614);
or U20982 (N_20982,N_20545,N_20551);
and U20983 (N_20983,N_20733,N_20546);
or U20984 (N_20984,N_20601,N_20733);
and U20985 (N_20985,N_20575,N_20627);
nand U20986 (N_20986,N_20728,N_20622);
xnor U20987 (N_20987,N_20541,N_20637);
nand U20988 (N_20988,N_20569,N_20712);
nand U20989 (N_20989,N_20623,N_20662);
nor U20990 (N_20990,N_20645,N_20595);
nor U20991 (N_20991,N_20695,N_20591);
nor U20992 (N_20992,N_20510,N_20523);
and U20993 (N_20993,N_20631,N_20735);
nor U20994 (N_20994,N_20713,N_20592);
and U20995 (N_20995,N_20592,N_20664);
xor U20996 (N_20996,N_20511,N_20639);
and U20997 (N_20997,N_20699,N_20535);
nand U20998 (N_20998,N_20527,N_20603);
nand U20999 (N_20999,N_20583,N_20518);
xor U21000 (N_21000,N_20953,N_20938);
nand U21001 (N_21001,N_20885,N_20910);
nor U21002 (N_21002,N_20882,N_20987);
and U21003 (N_21003,N_20941,N_20828);
xnor U21004 (N_21004,N_20848,N_20928);
nand U21005 (N_21005,N_20994,N_20875);
xnor U21006 (N_21006,N_20929,N_20786);
and U21007 (N_21007,N_20763,N_20858);
nand U21008 (N_21008,N_20922,N_20901);
and U21009 (N_21009,N_20954,N_20881);
nand U21010 (N_21010,N_20880,N_20797);
or U21011 (N_21011,N_20785,N_20972);
xor U21012 (N_21012,N_20908,N_20787);
nor U21013 (N_21013,N_20969,N_20865);
and U21014 (N_21014,N_20988,N_20822);
xor U21015 (N_21015,N_20951,N_20896);
nand U21016 (N_21016,N_20860,N_20892);
and U21017 (N_21017,N_20996,N_20809);
xor U21018 (N_21018,N_20773,N_20830);
nor U21019 (N_21019,N_20889,N_20779);
nand U21020 (N_21020,N_20991,N_20980);
xnor U21021 (N_21021,N_20837,N_20873);
nand U21022 (N_21022,N_20754,N_20981);
nand U21023 (N_21023,N_20757,N_20820);
or U21024 (N_21024,N_20920,N_20758);
or U21025 (N_21025,N_20755,N_20950);
nor U21026 (N_21026,N_20817,N_20884);
nand U21027 (N_21027,N_20766,N_20772);
or U21028 (N_21028,N_20958,N_20791);
and U21029 (N_21029,N_20923,N_20944);
nor U21030 (N_21030,N_20845,N_20843);
nor U21031 (N_21031,N_20831,N_20833);
nand U21032 (N_21032,N_20915,N_20924);
xnor U21033 (N_21033,N_20871,N_20826);
xor U21034 (N_21034,N_20811,N_20841);
xor U21035 (N_21035,N_20771,N_20899);
and U21036 (N_21036,N_20824,N_20936);
and U21037 (N_21037,N_20907,N_20770);
and U21038 (N_21038,N_20767,N_20973);
xnor U21039 (N_21039,N_20796,N_20983);
xnor U21040 (N_21040,N_20835,N_20840);
nor U21041 (N_21041,N_20753,N_20864);
nand U21042 (N_21042,N_20957,N_20829);
or U21043 (N_21043,N_20946,N_20813);
and U21044 (N_21044,N_20781,N_20808);
or U21045 (N_21045,N_20792,N_20879);
nor U21046 (N_21046,N_20890,N_20959);
nor U21047 (N_21047,N_20782,N_20912);
xor U21048 (N_21048,N_20863,N_20765);
xor U21049 (N_21049,N_20876,N_20776);
nor U21050 (N_21050,N_20818,N_20934);
xnor U21051 (N_21051,N_20764,N_20964);
or U21052 (N_21052,N_20806,N_20992);
nand U21053 (N_21053,N_20900,N_20793);
nor U21054 (N_21054,N_20943,N_20778);
xnor U21055 (N_21055,N_20842,N_20931);
and U21056 (N_21056,N_20825,N_20971);
or U21057 (N_21057,N_20846,N_20985);
nand U21058 (N_21058,N_20962,N_20760);
or U21059 (N_21059,N_20861,N_20878);
xnor U21060 (N_21060,N_20968,N_20850);
xor U21061 (N_21061,N_20844,N_20775);
and U21062 (N_21062,N_20997,N_20891);
nor U21063 (N_21063,N_20932,N_20898);
nor U21064 (N_21064,N_20952,N_20872);
and U21065 (N_21065,N_20868,N_20989);
nand U21066 (N_21066,N_20795,N_20945);
nor U21067 (N_21067,N_20832,N_20759);
nand U21068 (N_21068,N_20963,N_20966);
and U21069 (N_21069,N_20895,N_20993);
xor U21070 (N_21070,N_20851,N_20799);
and U21071 (N_21071,N_20852,N_20904);
and U21072 (N_21072,N_20762,N_20783);
nor U21073 (N_21073,N_20965,N_20769);
nor U21074 (N_21074,N_20918,N_20977);
xnor U21075 (N_21075,N_20866,N_20933);
nor U21076 (N_21076,N_20947,N_20916);
nand U21077 (N_21077,N_20784,N_20902);
nor U21078 (N_21078,N_20930,N_20810);
xor U21079 (N_21079,N_20780,N_20986);
nand U21080 (N_21080,N_20893,N_20847);
nor U21081 (N_21081,N_20883,N_20798);
nand U21082 (N_21082,N_20870,N_20927);
nor U21083 (N_21083,N_20926,N_20949);
nor U21084 (N_21084,N_20752,N_20836);
and U21085 (N_21085,N_20854,N_20849);
nor U21086 (N_21086,N_20812,N_20976);
nor U21087 (N_21087,N_20823,N_20834);
xnor U21088 (N_21088,N_20979,N_20940);
or U21089 (N_21089,N_20905,N_20935);
or U21090 (N_21090,N_20990,N_20982);
nor U21091 (N_21091,N_20995,N_20956);
nor U21092 (N_21092,N_20894,N_20961);
or U21093 (N_21093,N_20867,N_20942);
nand U21094 (N_21094,N_20768,N_20859);
or U21095 (N_21095,N_20777,N_20974);
xnor U21096 (N_21096,N_20827,N_20853);
nand U21097 (N_21097,N_20802,N_20917);
or U21098 (N_21098,N_20805,N_20801);
or U21099 (N_21099,N_20998,N_20948);
or U21100 (N_21100,N_20906,N_20761);
nor U21101 (N_21101,N_20970,N_20803);
and U21102 (N_21102,N_20999,N_20939);
and U21103 (N_21103,N_20921,N_20978);
nand U21104 (N_21104,N_20789,N_20960);
and U21105 (N_21105,N_20794,N_20975);
xnor U21106 (N_21106,N_20815,N_20819);
or U21107 (N_21107,N_20814,N_20937);
nor U21108 (N_21108,N_20807,N_20857);
and U21109 (N_21109,N_20821,N_20984);
nor U21110 (N_21110,N_20790,N_20911);
nand U21111 (N_21111,N_20909,N_20751);
and U21112 (N_21112,N_20897,N_20955);
nor U21113 (N_21113,N_20750,N_20887);
nor U21114 (N_21114,N_20839,N_20838);
nand U21115 (N_21115,N_20869,N_20967);
nor U21116 (N_21116,N_20804,N_20919);
or U21117 (N_21117,N_20914,N_20913);
or U21118 (N_21118,N_20886,N_20774);
or U21119 (N_21119,N_20903,N_20877);
xor U21120 (N_21120,N_20862,N_20925);
xor U21121 (N_21121,N_20788,N_20874);
nor U21122 (N_21122,N_20888,N_20756);
and U21123 (N_21123,N_20855,N_20800);
nand U21124 (N_21124,N_20816,N_20856);
xor U21125 (N_21125,N_20969,N_20931);
nor U21126 (N_21126,N_20992,N_20811);
and U21127 (N_21127,N_20980,N_20916);
nor U21128 (N_21128,N_20923,N_20832);
nor U21129 (N_21129,N_20970,N_20861);
nor U21130 (N_21130,N_20830,N_20785);
or U21131 (N_21131,N_20934,N_20932);
or U21132 (N_21132,N_20808,N_20881);
and U21133 (N_21133,N_20872,N_20923);
and U21134 (N_21134,N_20945,N_20937);
nand U21135 (N_21135,N_20848,N_20901);
nor U21136 (N_21136,N_20932,N_20963);
xor U21137 (N_21137,N_20859,N_20964);
nand U21138 (N_21138,N_20773,N_20797);
nor U21139 (N_21139,N_20779,N_20991);
xnor U21140 (N_21140,N_20755,N_20871);
nand U21141 (N_21141,N_20811,N_20898);
xor U21142 (N_21142,N_20958,N_20821);
or U21143 (N_21143,N_20998,N_20767);
or U21144 (N_21144,N_20859,N_20755);
and U21145 (N_21145,N_20957,N_20841);
or U21146 (N_21146,N_20900,N_20790);
nor U21147 (N_21147,N_20835,N_20811);
and U21148 (N_21148,N_20927,N_20799);
nor U21149 (N_21149,N_20943,N_20802);
and U21150 (N_21150,N_20833,N_20752);
or U21151 (N_21151,N_20914,N_20953);
nor U21152 (N_21152,N_20777,N_20754);
or U21153 (N_21153,N_20960,N_20902);
nor U21154 (N_21154,N_20828,N_20910);
nand U21155 (N_21155,N_20873,N_20882);
and U21156 (N_21156,N_20854,N_20936);
or U21157 (N_21157,N_20798,N_20860);
nand U21158 (N_21158,N_20775,N_20897);
or U21159 (N_21159,N_20989,N_20924);
nand U21160 (N_21160,N_20997,N_20912);
nand U21161 (N_21161,N_20951,N_20940);
or U21162 (N_21162,N_20756,N_20957);
and U21163 (N_21163,N_20776,N_20994);
or U21164 (N_21164,N_20963,N_20797);
nor U21165 (N_21165,N_20829,N_20906);
xnor U21166 (N_21166,N_20826,N_20800);
or U21167 (N_21167,N_20987,N_20926);
or U21168 (N_21168,N_20909,N_20897);
nand U21169 (N_21169,N_20956,N_20953);
xor U21170 (N_21170,N_20959,N_20972);
nand U21171 (N_21171,N_20873,N_20751);
nor U21172 (N_21172,N_20999,N_20894);
nand U21173 (N_21173,N_20831,N_20859);
nand U21174 (N_21174,N_20928,N_20911);
and U21175 (N_21175,N_20918,N_20929);
nand U21176 (N_21176,N_20972,N_20843);
nor U21177 (N_21177,N_20915,N_20916);
or U21178 (N_21178,N_20832,N_20883);
nor U21179 (N_21179,N_20862,N_20784);
and U21180 (N_21180,N_20788,N_20984);
and U21181 (N_21181,N_20818,N_20956);
and U21182 (N_21182,N_20892,N_20950);
xnor U21183 (N_21183,N_20857,N_20875);
and U21184 (N_21184,N_20936,N_20993);
and U21185 (N_21185,N_20803,N_20991);
nand U21186 (N_21186,N_20922,N_20818);
nor U21187 (N_21187,N_20945,N_20877);
and U21188 (N_21188,N_20974,N_20907);
xnor U21189 (N_21189,N_20917,N_20766);
nand U21190 (N_21190,N_20834,N_20887);
nor U21191 (N_21191,N_20841,N_20999);
and U21192 (N_21192,N_20785,N_20834);
and U21193 (N_21193,N_20880,N_20803);
and U21194 (N_21194,N_20888,N_20835);
and U21195 (N_21195,N_20926,N_20924);
nand U21196 (N_21196,N_20873,N_20970);
or U21197 (N_21197,N_20941,N_20800);
or U21198 (N_21198,N_20856,N_20810);
nand U21199 (N_21199,N_20937,N_20991);
nand U21200 (N_21200,N_20893,N_20866);
or U21201 (N_21201,N_20806,N_20805);
nor U21202 (N_21202,N_20934,N_20889);
nor U21203 (N_21203,N_20967,N_20758);
xnor U21204 (N_21204,N_20962,N_20865);
and U21205 (N_21205,N_20900,N_20794);
and U21206 (N_21206,N_20871,N_20932);
or U21207 (N_21207,N_20844,N_20947);
nor U21208 (N_21208,N_20812,N_20783);
and U21209 (N_21209,N_20904,N_20806);
nor U21210 (N_21210,N_20992,N_20773);
nand U21211 (N_21211,N_20887,N_20993);
and U21212 (N_21212,N_20869,N_20751);
nor U21213 (N_21213,N_20874,N_20824);
or U21214 (N_21214,N_20752,N_20827);
and U21215 (N_21215,N_20754,N_20928);
nor U21216 (N_21216,N_20922,N_20911);
nand U21217 (N_21217,N_20833,N_20750);
nand U21218 (N_21218,N_20828,N_20848);
nand U21219 (N_21219,N_20815,N_20784);
nand U21220 (N_21220,N_20904,N_20837);
xnor U21221 (N_21221,N_20832,N_20970);
nand U21222 (N_21222,N_20961,N_20757);
xor U21223 (N_21223,N_20827,N_20814);
nor U21224 (N_21224,N_20866,N_20991);
or U21225 (N_21225,N_20957,N_20959);
nor U21226 (N_21226,N_20842,N_20782);
or U21227 (N_21227,N_20920,N_20785);
nand U21228 (N_21228,N_20911,N_20854);
nand U21229 (N_21229,N_20854,N_20890);
and U21230 (N_21230,N_20887,N_20818);
and U21231 (N_21231,N_20931,N_20763);
xor U21232 (N_21232,N_20998,N_20786);
or U21233 (N_21233,N_20840,N_20925);
nor U21234 (N_21234,N_20964,N_20790);
and U21235 (N_21235,N_20902,N_20779);
nand U21236 (N_21236,N_20854,N_20879);
or U21237 (N_21237,N_20880,N_20817);
and U21238 (N_21238,N_20812,N_20915);
xor U21239 (N_21239,N_20968,N_20908);
or U21240 (N_21240,N_20871,N_20867);
nand U21241 (N_21241,N_20961,N_20753);
and U21242 (N_21242,N_20984,N_20826);
and U21243 (N_21243,N_20824,N_20999);
or U21244 (N_21244,N_20964,N_20804);
or U21245 (N_21245,N_20855,N_20834);
nor U21246 (N_21246,N_20903,N_20944);
xor U21247 (N_21247,N_20968,N_20953);
or U21248 (N_21248,N_20815,N_20804);
nand U21249 (N_21249,N_20828,N_20817);
or U21250 (N_21250,N_21248,N_21244);
or U21251 (N_21251,N_21167,N_21118);
or U21252 (N_21252,N_21245,N_21038);
nand U21253 (N_21253,N_21015,N_21126);
nand U21254 (N_21254,N_21107,N_21215);
xnor U21255 (N_21255,N_21055,N_21064);
or U21256 (N_21256,N_21026,N_21174);
nand U21257 (N_21257,N_21058,N_21071);
nor U21258 (N_21258,N_21082,N_21124);
nor U21259 (N_21259,N_21079,N_21182);
or U21260 (N_21260,N_21194,N_21022);
and U21261 (N_21261,N_21185,N_21001);
and U21262 (N_21262,N_21208,N_21122);
and U21263 (N_21263,N_21009,N_21191);
nand U21264 (N_21264,N_21155,N_21128);
or U21265 (N_21265,N_21057,N_21175);
or U21266 (N_21266,N_21065,N_21223);
nor U21267 (N_21267,N_21203,N_21123);
nor U21268 (N_21268,N_21031,N_21229);
nand U21269 (N_21269,N_21137,N_21041);
nor U21270 (N_21270,N_21192,N_21100);
nor U21271 (N_21271,N_21220,N_21161);
nand U21272 (N_21272,N_21042,N_21154);
or U21273 (N_21273,N_21177,N_21050);
and U21274 (N_21274,N_21000,N_21091);
nand U21275 (N_21275,N_21246,N_21039);
nand U21276 (N_21276,N_21097,N_21078);
nand U21277 (N_21277,N_21088,N_21213);
xnor U21278 (N_21278,N_21206,N_21146);
xor U21279 (N_21279,N_21074,N_21149);
nand U21280 (N_21280,N_21049,N_21111);
and U21281 (N_21281,N_21209,N_21008);
nor U21282 (N_21282,N_21136,N_21061);
or U21283 (N_21283,N_21013,N_21232);
nor U21284 (N_21284,N_21035,N_21093);
nand U21285 (N_21285,N_21186,N_21235);
xor U21286 (N_21286,N_21181,N_21187);
and U21287 (N_21287,N_21032,N_21135);
and U21288 (N_21288,N_21212,N_21153);
nor U21289 (N_21289,N_21142,N_21076);
or U21290 (N_21290,N_21120,N_21140);
nor U21291 (N_21291,N_21138,N_21019);
xnor U21292 (N_21292,N_21133,N_21047);
xor U21293 (N_21293,N_21021,N_21075);
xor U21294 (N_21294,N_21024,N_21114);
and U21295 (N_21295,N_21188,N_21085);
and U21296 (N_21296,N_21169,N_21166);
nor U21297 (N_21297,N_21150,N_21033);
and U21298 (N_21298,N_21204,N_21106);
nor U21299 (N_21299,N_21034,N_21094);
nand U21300 (N_21300,N_21109,N_21130);
xor U21301 (N_21301,N_21226,N_21077);
and U21302 (N_21302,N_21131,N_21016);
or U21303 (N_21303,N_21051,N_21083);
or U21304 (N_21304,N_21028,N_21004);
and U21305 (N_21305,N_21060,N_21224);
or U21306 (N_21306,N_21179,N_21184);
and U21307 (N_21307,N_21110,N_21171);
and U21308 (N_21308,N_21214,N_21062);
nor U21309 (N_21309,N_21147,N_21233);
nand U21310 (N_21310,N_21143,N_21198);
xnor U21311 (N_21311,N_21127,N_21070);
or U21312 (N_21312,N_21092,N_21098);
nor U21313 (N_21313,N_21073,N_21003);
xnor U21314 (N_21314,N_21164,N_21096);
nor U21315 (N_21315,N_21219,N_21129);
or U21316 (N_21316,N_21247,N_21027);
nor U21317 (N_21317,N_21230,N_21172);
xor U21318 (N_21318,N_21242,N_21053);
nor U21319 (N_21319,N_21228,N_21225);
nor U21320 (N_21320,N_21210,N_21002);
or U21321 (N_21321,N_21211,N_21040);
nor U21322 (N_21322,N_21103,N_21072);
xor U21323 (N_21323,N_21159,N_21020);
xor U21324 (N_21324,N_21087,N_21236);
and U21325 (N_21325,N_21139,N_21134);
or U21326 (N_21326,N_21056,N_21066);
or U21327 (N_21327,N_21160,N_21165);
and U21328 (N_21328,N_21157,N_21014);
nor U21329 (N_21329,N_21018,N_21005);
or U21330 (N_21330,N_21141,N_21036);
nand U21331 (N_21331,N_21037,N_21086);
xor U21332 (N_21332,N_21156,N_21237);
and U21333 (N_21333,N_21168,N_21116);
and U21334 (N_21334,N_21195,N_21202);
nand U21335 (N_21335,N_21059,N_21231);
xnor U21336 (N_21336,N_21006,N_21189);
nand U21337 (N_21337,N_21069,N_21145);
and U21338 (N_21338,N_21102,N_21081);
nand U21339 (N_21339,N_21112,N_21068);
or U21340 (N_21340,N_21207,N_21201);
or U21341 (N_21341,N_21176,N_21241);
nor U21342 (N_21342,N_21044,N_21234);
and U21343 (N_21343,N_21029,N_21151);
and U21344 (N_21344,N_21067,N_21063);
and U21345 (N_21345,N_21043,N_21115);
and U21346 (N_21346,N_21183,N_21054);
nor U21347 (N_21347,N_21023,N_21239);
and U21348 (N_21348,N_21012,N_21010);
nor U21349 (N_21349,N_21105,N_21217);
or U21350 (N_21350,N_21190,N_21095);
or U21351 (N_21351,N_21025,N_21243);
or U21352 (N_21352,N_21148,N_21099);
and U21353 (N_21353,N_21080,N_21117);
nor U21354 (N_21354,N_21249,N_21197);
xnor U21355 (N_21355,N_21200,N_21125);
or U21356 (N_21356,N_21144,N_21178);
nand U21357 (N_21357,N_21007,N_21238);
xor U21358 (N_21358,N_21170,N_21101);
xnor U21359 (N_21359,N_21104,N_21152);
nor U21360 (N_21360,N_21132,N_21216);
nand U21361 (N_21361,N_21108,N_21048);
or U21362 (N_21362,N_21196,N_21121);
nand U21363 (N_21363,N_21199,N_21218);
xor U21364 (N_21364,N_21180,N_21119);
or U21365 (N_21365,N_21017,N_21162);
or U21366 (N_21366,N_21030,N_21158);
nor U21367 (N_21367,N_21090,N_21227);
nand U21368 (N_21368,N_21173,N_21193);
and U21369 (N_21369,N_21221,N_21163);
nor U21370 (N_21370,N_21011,N_21113);
nor U21371 (N_21371,N_21240,N_21052);
or U21372 (N_21372,N_21084,N_21089);
and U21373 (N_21373,N_21045,N_21205);
nand U21374 (N_21374,N_21046,N_21222);
and U21375 (N_21375,N_21215,N_21223);
or U21376 (N_21376,N_21046,N_21184);
xor U21377 (N_21377,N_21222,N_21148);
or U21378 (N_21378,N_21007,N_21165);
or U21379 (N_21379,N_21143,N_21035);
xor U21380 (N_21380,N_21113,N_21049);
nor U21381 (N_21381,N_21209,N_21061);
or U21382 (N_21382,N_21181,N_21020);
nand U21383 (N_21383,N_21059,N_21195);
or U21384 (N_21384,N_21110,N_21026);
nor U21385 (N_21385,N_21211,N_21002);
nand U21386 (N_21386,N_21151,N_21243);
nand U21387 (N_21387,N_21224,N_21125);
xor U21388 (N_21388,N_21203,N_21042);
or U21389 (N_21389,N_21014,N_21057);
nor U21390 (N_21390,N_21051,N_21158);
and U21391 (N_21391,N_21155,N_21145);
and U21392 (N_21392,N_21119,N_21200);
nand U21393 (N_21393,N_21203,N_21160);
nand U21394 (N_21394,N_21106,N_21020);
nand U21395 (N_21395,N_21041,N_21104);
nand U21396 (N_21396,N_21180,N_21212);
nand U21397 (N_21397,N_21028,N_21177);
nor U21398 (N_21398,N_21028,N_21175);
nor U21399 (N_21399,N_21120,N_21135);
nor U21400 (N_21400,N_21065,N_21224);
nor U21401 (N_21401,N_21243,N_21146);
and U21402 (N_21402,N_21026,N_21213);
or U21403 (N_21403,N_21161,N_21077);
and U21404 (N_21404,N_21129,N_21075);
nand U21405 (N_21405,N_21099,N_21062);
nand U21406 (N_21406,N_21208,N_21165);
nor U21407 (N_21407,N_21070,N_21105);
nand U21408 (N_21408,N_21101,N_21208);
and U21409 (N_21409,N_21183,N_21079);
and U21410 (N_21410,N_21235,N_21225);
nor U21411 (N_21411,N_21236,N_21028);
nor U21412 (N_21412,N_21083,N_21205);
nand U21413 (N_21413,N_21229,N_21074);
nor U21414 (N_21414,N_21152,N_21243);
or U21415 (N_21415,N_21057,N_21199);
nor U21416 (N_21416,N_21033,N_21218);
xor U21417 (N_21417,N_21004,N_21037);
xor U21418 (N_21418,N_21243,N_21042);
and U21419 (N_21419,N_21236,N_21062);
and U21420 (N_21420,N_21195,N_21178);
nand U21421 (N_21421,N_21002,N_21094);
nor U21422 (N_21422,N_21190,N_21012);
nand U21423 (N_21423,N_21137,N_21142);
or U21424 (N_21424,N_21237,N_21136);
or U21425 (N_21425,N_21049,N_21169);
or U21426 (N_21426,N_21146,N_21175);
xnor U21427 (N_21427,N_21189,N_21190);
and U21428 (N_21428,N_21146,N_21093);
or U21429 (N_21429,N_21151,N_21124);
nand U21430 (N_21430,N_21004,N_21136);
and U21431 (N_21431,N_21113,N_21233);
or U21432 (N_21432,N_21116,N_21086);
nand U21433 (N_21433,N_21158,N_21050);
nor U21434 (N_21434,N_21164,N_21186);
nand U21435 (N_21435,N_21230,N_21247);
nand U21436 (N_21436,N_21205,N_21175);
nor U21437 (N_21437,N_21107,N_21165);
xnor U21438 (N_21438,N_21184,N_21052);
nor U21439 (N_21439,N_21159,N_21177);
nor U21440 (N_21440,N_21040,N_21018);
xor U21441 (N_21441,N_21152,N_21196);
nor U21442 (N_21442,N_21244,N_21163);
or U21443 (N_21443,N_21103,N_21119);
nor U21444 (N_21444,N_21018,N_21065);
xor U21445 (N_21445,N_21209,N_21023);
or U21446 (N_21446,N_21073,N_21167);
and U21447 (N_21447,N_21001,N_21117);
nor U21448 (N_21448,N_21237,N_21204);
nor U21449 (N_21449,N_21213,N_21182);
xnor U21450 (N_21450,N_21081,N_21238);
or U21451 (N_21451,N_21233,N_21093);
and U21452 (N_21452,N_21046,N_21025);
xnor U21453 (N_21453,N_21220,N_21132);
xnor U21454 (N_21454,N_21243,N_21214);
xnor U21455 (N_21455,N_21105,N_21165);
or U21456 (N_21456,N_21048,N_21191);
or U21457 (N_21457,N_21213,N_21076);
nor U21458 (N_21458,N_21155,N_21232);
xor U21459 (N_21459,N_21048,N_21058);
or U21460 (N_21460,N_21065,N_21010);
xor U21461 (N_21461,N_21238,N_21195);
or U21462 (N_21462,N_21131,N_21045);
nand U21463 (N_21463,N_21237,N_21038);
and U21464 (N_21464,N_21166,N_21154);
or U21465 (N_21465,N_21225,N_21058);
nand U21466 (N_21466,N_21073,N_21117);
and U21467 (N_21467,N_21224,N_21184);
and U21468 (N_21468,N_21005,N_21009);
or U21469 (N_21469,N_21214,N_21161);
xnor U21470 (N_21470,N_21026,N_21002);
or U21471 (N_21471,N_21210,N_21070);
and U21472 (N_21472,N_21203,N_21105);
xor U21473 (N_21473,N_21016,N_21171);
and U21474 (N_21474,N_21031,N_21222);
and U21475 (N_21475,N_21194,N_21068);
or U21476 (N_21476,N_21006,N_21023);
nor U21477 (N_21477,N_21114,N_21217);
nor U21478 (N_21478,N_21194,N_21058);
nor U21479 (N_21479,N_21124,N_21065);
and U21480 (N_21480,N_21102,N_21041);
or U21481 (N_21481,N_21247,N_21081);
nand U21482 (N_21482,N_21132,N_21016);
nand U21483 (N_21483,N_21003,N_21001);
xor U21484 (N_21484,N_21081,N_21243);
and U21485 (N_21485,N_21051,N_21142);
nand U21486 (N_21486,N_21034,N_21074);
or U21487 (N_21487,N_21101,N_21138);
and U21488 (N_21488,N_21031,N_21243);
or U21489 (N_21489,N_21206,N_21126);
and U21490 (N_21490,N_21195,N_21181);
or U21491 (N_21491,N_21137,N_21052);
xnor U21492 (N_21492,N_21231,N_21093);
xnor U21493 (N_21493,N_21096,N_21062);
xor U21494 (N_21494,N_21017,N_21097);
nor U21495 (N_21495,N_21189,N_21210);
nor U21496 (N_21496,N_21011,N_21135);
nand U21497 (N_21497,N_21063,N_21218);
xnor U21498 (N_21498,N_21011,N_21062);
xnor U21499 (N_21499,N_21166,N_21149);
and U21500 (N_21500,N_21304,N_21390);
and U21501 (N_21501,N_21379,N_21311);
xnor U21502 (N_21502,N_21387,N_21294);
xor U21503 (N_21503,N_21307,N_21347);
nor U21504 (N_21504,N_21456,N_21290);
or U21505 (N_21505,N_21406,N_21269);
or U21506 (N_21506,N_21392,N_21339);
and U21507 (N_21507,N_21498,N_21431);
and U21508 (N_21508,N_21413,N_21358);
nor U21509 (N_21509,N_21354,N_21409);
xnor U21510 (N_21510,N_21486,N_21322);
nand U21511 (N_21511,N_21285,N_21432);
nand U21512 (N_21512,N_21493,N_21384);
nand U21513 (N_21513,N_21483,N_21455);
xor U21514 (N_21514,N_21378,N_21286);
and U21515 (N_21515,N_21489,N_21436);
nand U21516 (N_21516,N_21444,N_21316);
nand U21517 (N_21517,N_21359,N_21385);
and U21518 (N_21518,N_21492,N_21266);
and U21519 (N_21519,N_21407,N_21345);
xnor U21520 (N_21520,N_21424,N_21302);
or U21521 (N_21521,N_21441,N_21484);
xor U21522 (N_21522,N_21458,N_21496);
xnor U21523 (N_21523,N_21270,N_21418);
nand U21524 (N_21524,N_21466,N_21461);
xor U21525 (N_21525,N_21487,N_21405);
nand U21526 (N_21526,N_21494,N_21279);
or U21527 (N_21527,N_21342,N_21250);
nand U21528 (N_21528,N_21317,N_21420);
nand U21529 (N_21529,N_21370,N_21454);
and U21530 (N_21530,N_21457,N_21333);
or U21531 (N_21531,N_21388,N_21336);
xnor U21532 (N_21532,N_21439,N_21491);
xnor U21533 (N_21533,N_21337,N_21459);
nor U21534 (N_21534,N_21373,N_21481);
and U21535 (N_21535,N_21429,N_21395);
and U21536 (N_21536,N_21295,N_21319);
nand U21537 (N_21537,N_21453,N_21371);
xor U21538 (N_21538,N_21450,N_21306);
nor U21539 (N_21539,N_21289,N_21356);
and U21540 (N_21540,N_21293,N_21334);
nand U21541 (N_21541,N_21391,N_21326);
nor U21542 (N_21542,N_21472,N_21414);
and U21543 (N_21543,N_21366,N_21433);
nor U21544 (N_21544,N_21460,N_21473);
xnor U21545 (N_21545,N_21437,N_21301);
nor U21546 (N_21546,N_21434,N_21416);
xor U21547 (N_21547,N_21386,N_21321);
xnor U21548 (N_21548,N_21251,N_21365);
nor U21549 (N_21549,N_21495,N_21393);
and U21550 (N_21550,N_21445,N_21362);
or U21551 (N_21551,N_21330,N_21258);
and U21552 (N_21552,N_21309,N_21482);
or U21553 (N_21553,N_21363,N_21297);
and U21554 (N_21554,N_21464,N_21257);
xnor U21555 (N_21555,N_21288,N_21446);
or U21556 (N_21556,N_21467,N_21476);
xor U21557 (N_21557,N_21318,N_21299);
nor U21558 (N_21558,N_21300,N_21320);
nor U21559 (N_21559,N_21314,N_21374);
xnor U21560 (N_21560,N_21485,N_21353);
nand U21561 (N_21561,N_21471,N_21283);
nand U21562 (N_21562,N_21335,N_21463);
nand U21563 (N_21563,N_21327,N_21348);
nor U21564 (N_21564,N_21351,N_21470);
nor U21565 (N_21565,N_21389,N_21435);
nor U21566 (N_21566,N_21282,N_21465);
nand U21567 (N_21567,N_21462,N_21346);
or U21568 (N_21568,N_21369,N_21253);
xnor U21569 (N_21569,N_21367,N_21377);
or U21570 (N_21570,N_21260,N_21276);
or U21571 (N_21571,N_21397,N_21394);
nor U21572 (N_21572,N_21448,N_21343);
and U21573 (N_21573,N_21400,N_21344);
nor U21574 (N_21574,N_21252,N_21408);
nand U21575 (N_21575,N_21273,N_21428);
or U21576 (N_21576,N_21468,N_21259);
and U21577 (N_21577,N_21313,N_21488);
nor U21578 (N_21578,N_21310,N_21490);
nor U21579 (N_21579,N_21263,N_21469);
or U21580 (N_21580,N_21399,N_21368);
and U21581 (N_21581,N_21262,N_21277);
or U21582 (N_21582,N_21372,N_21425);
nand U21583 (N_21583,N_21328,N_21324);
nand U21584 (N_21584,N_21338,N_21254);
nand U21585 (N_21585,N_21323,N_21264);
and U21586 (N_21586,N_21275,N_21291);
and U21587 (N_21587,N_21325,N_21440);
nor U21588 (N_21588,N_21315,N_21402);
and U21589 (N_21589,N_21298,N_21380);
and U21590 (N_21590,N_21438,N_21340);
xor U21591 (N_21591,N_21331,N_21422);
or U21592 (N_21592,N_21376,N_21447);
and U21593 (N_21593,N_21364,N_21443);
nand U21594 (N_21594,N_21267,N_21261);
xor U21595 (N_21595,N_21474,N_21398);
nand U21596 (N_21596,N_21401,N_21360);
or U21597 (N_21597,N_21478,N_21427);
nand U21598 (N_21598,N_21423,N_21442);
nor U21599 (N_21599,N_21375,N_21396);
or U21600 (N_21600,N_21271,N_21265);
xor U21601 (N_21601,N_21421,N_21357);
nor U21602 (N_21602,N_21349,N_21452);
nor U21603 (N_21603,N_21287,N_21278);
and U21604 (N_21604,N_21341,N_21382);
nor U21605 (N_21605,N_21499,N_21305);
and U21606 (N_21606,N_21352,N_21403);
or U21607 (N_21607,N_21417,N_21479);
nor U21608 (N_21608,N_21255,N_21274);
and U21609 (N_21609,N_21280,N_21451);
nor U21610 (N_21610,N_21350,N_21449);
xor U21611 (N_21611,N_21268,N_21480);
and U21612 (N_21612,N_21381,N_21419);
nand U21613 (N_21613,N_21292,N_21475);
nor U21614 (N_21614,N_21256,N_21361);
xor U21615 (N_21615,N_21303,N_21415);
or U21616 (N_21616,N_21497,N_21411);
and U21617 (N_21617,N_21332,N_21281);
xnor U21618 (N_21618,N_21355,N_21430);
nor U21619 (N_21619,N_21477,N_21426);
nand U21620 (N_21620,N_21284,N_21312);
nand U21621 (N_21621,N_21412,N_21272);
or U21622 (N_21622,N_21329,N_21383);
and U21623 (N_21623,N_21410,N_21308);
xor U21624 (N_21624,N_21296,N_21404);
or U21625 (N_21625,N_21468,N_21499);
or U21626 (N_21626,N_21444,N_21483);
and U21627 (N_21627,N_21270,N_21395);
nor U21628 (N_21628,N_21307,N_21345);
and U21629 (N_21629,N_21353,N_21254);
or U21630 (N_21630,N_21260,N_21401);
xnor U21631 (N_21631,N_21383,N_21394);
nand U21632 (N_21632,N_21434,N_21384);
nor U21633 (N_21633,N_21380,N_21454);
nor U21634 (N_21634,N_21294,N_21465);
and U21635 (N_21635,N_21418,N_21469);
or U21636 (N_21636,N_21478,N_21324);
and U21637 (N_21637,N_21452,N_21475);
and U21638 (N_21638,N_21317,N_21363);
nor U21639 (N_21639,N_21461,N_21286);
or U21640 (N_21640,N_21352,N_21436);
and U21641 (N_21641,N_21309,N_21483);
nand U21642 (N_21642,N_21416,N_21339);
xnor U21643 (N_21643,N_21494,N_21280);
and U21644 (N_21644,N_21389,N_21437);
xor U21645 (N_21645,N_21263,N_21290);
xor U21646 (N_21646,N_21441,N_21455);
nor U21647 (N_21647,N_21291,N_21268);
nor U21648 (N_21648,N_21317,N_21290);
nand U21649 (N_21649,N_21450,N_21354);
or U21650 (N_21650,N_21443,N_21397);
xor U21651 (N_21651,N_21340,N_21418);
xor U21652 (N_21652,N_21286,N_21366);
xor U21653 (N_21653,N_21288,N_21427);
nand U21654 (N_21654,N_21274,N_21457);
nor U21655 (N_21655,N_21285,N_21428);
nor U21656 (N_21656,N_21350,N_21288);
nand U21657 (N_21657,N_21430,N_21482);
and U21658 (N_21658,N_21475,N_21379);
xor U21659 (N_21659,N_21455,N_21352);
or U21660 (N_21660,N_21327,N_21388);
nor U21661 (N_21661,N_21471,N_21470);
or U21662 (N_21662,N_21268,N_21450);
xor U21663 (N_21663,N_21314,N_21467);
xor U21664 (N_21664,N_21288,N_21399);
nor U21665 (N_21665,N_21299,N_21315);
or U21666 (N_21666,N_21398,N_21323);
and U21667 (N_21667,N_21318,N_21341);
xnor U21668 (N_21668,N_21319,N_21276);
or U21669 (N_21669,N_21316,N_21383);
nand U21670 (N_21670,N_21455,N_21300);
nand U21671 (N_21671,N_21253,N_21378);
nand U21672 (N_21672,N_21345,N_21439);
nand U21673 (N_21673,N_21401,N_21299);
or U21674 (N_21674,N_21269,N_21263);
nor U21675 (N_21675,N_21384,N_21476);
xnor U21676 (N_21676,N_21495,N_21452);
and U21677 (N_21677,N_21276,N_21346);
xnor U21678 (N_21678,N_21368,N_21441);
or U21679 (N_21679,N_21498,N_21451);
nor U21680 (N_21680,N_21314,N_21280);
or U21681 (N_21681,N_21393,N_21311);
or U21682 (N_21682,N_21293,N_21376);
nand U21683 (N_21683,N_21283,N_21285);
or U21684 (N_21684,N_21413,N_21435);
and U21685 (N_21685,N_21496,N_21305);
nor U21686 (N_21686,N_21253,N_21485);
and U21687 (N_21687,N_21258,N_21349);
or U21688 (N_21688,N_21391,N_21320);
xor U21689 (N_21689,N_21416,N_21281);
xor U21690 (N_21690,N_21432,N_21392);
nor U21691 (N_21691,N_21475,N_21280);
nand U21692 (N_21692,N_21367,N_21360);
nand U21693 (N_21693,N_21490,N_21442);
xnor U21694 (N_21694,N_21380,N_21355);
nand U21695 (N_21695,N_21305,N_21382);
and U21696 (N_21696,N_21367,N_21428);
or U21697 (N_21697,N_21342,N_21356);
xnor U21698 (N_21698,N_21300,N_21362);
nand U21699 (N_21699,N_21453,N_21367);
xor U21700 (N_21700,N_21353,N_21337);
nand U21701 (N_21701,N_21479,N_21305);
and U21702 (N_21702,N_21394,N_21409);
nand U21703 (N_21703,N_21309,N_21459);
nand U21704 (N_21704,N_21325,N_21359);
or U21705 (N_21705,N_21433,N_21365);
nor U21706 (N_21706,N_21459,N_21495);
and U21707 (N_21707,N_21367,N_21459);
or U21708 (N_21708,N_21291,N_21401);
and U21709 (N_21709,N_21404,N_21376);
or U21710 (N_21710,N_21351,N_21287);
and U21711 (N_21711,N_21461,N_21474);
and U21712 (N_21712,N_21349,N_21305);
nand U21713 (N_21713,N_21361,N_21441);
nand U21714 (N_21714,N_21461,N_21349);
or U21715 (N_21715,N_21377,N_21267);
and U21716 (N_21716,N_21473,N_21407);
xor U21717 (N_21717,N_21385,N_21255);
xor U21718 (N_21718,N_21452,N_21369);
nand U21719 (N_21719,N_21371,N_21447);
and U21720 (N_21720,N_21449,N_21252);
or U21721 (N_21721,N_21487,N_21477);
or U21722 (N_21722,N_21469,N_21448);
xnor U21723 (N_21723,N_21329,N_21389);
xnor U21724 (N_21724,N_21274,N_21488);
nor U21725 (N_21725,N_21385,N_21401);
xor U21726 (N_21726,N_21423,N_21497);
and U21727 (N_21727,N_21340,N_21400);
and U21728 (N_21728,N_21472,N_21300);
or U21729 (N_21729,N_21487,N_21352);
nor U21730 (N_21730,N_21330,N_21341);
and U21731 (N_21731,N_21336,N_21366);
or U21732 (N_21732,N_21458,N_21310);
and U21733 (N_21733,N_21459,N_21385);
xnor U21734 (N_21734,N_21490,N_21254);
xor U21735 (N_21735,N_21308,N_21253);
and U21736 (N_21736,N_21410,N_21469);
nor U21737 (N_21737,N_21316,N_21321);
xnor U21738 (N_21738,N_21443,N_21427);
nand U21739 (N_21739,N_21443,N_21496);
or U21740 (N_21740,N_21277,N_21467);
and U21741 (N_21741,N_21327,N_21413);
or U21742 (N_21742,N_21402,N_21449);
nand U21743 (N_21743,N_21468,N_21329);
and U21744 (N_21744,N_21260,N_21442);
or U21745 (N_21745,N_21374,N_21382);
nor U21746 (N_21746,N_21296,N_21349);
nor U21747 (N_21747,N_21470,N_21266);
and U21748 (N_21748,N_21388,N_21469);
nand U21749 (N_21749,N_21332,N_21355);
or U21750 (N_21750,N_21647,N_21745);
nor U21751 (N_21751,N_21725,N_21685);
nor U21752 (N_21752,N_21518,N_21541);
nand U21753 (N_21753,N_21503,N_21597);
xnor U21754 (N_21754,N_21687,N_21568);
and U21755 (N_21755,N_21580,N_21555);
nor U21756 (N_21756,N_21623,N_21509);
and U21757 (N_21757,N_21632,N_21746);
xor U21758 (N_21758,N_21524,N_21735);
or U21759 (N_21759,N_21537,N_21507);
nand U21760 (N_21760,N_21646,N_21566);
and U21761 (N_21761,N_21604,N_21523);
nor U21762 (N_21762,N_21726,N_21668);
xnor U21763 (N_21763,N_21689,N_21563);
nor U21764 (N_21764,N_21630,N_21591);
nor U21765 (N_21765,N_21651,N_21637);
xor U21766 (N_21766,N_21716,N_21641);
or U21767 (N_21767,N_21528,N_21636);
or U21768 (N_21768,N_21655,N_21542);
nand U21769 (N_21769,N_21512,N_21624);
nand U21770 (N_21770,N_21607,N_21686);
and U21771 (N_21771,N_21748,N_21645);
or U21772 (N_21772,N_21663,N_21556);
nand U21773 (N_21773,N_21625,N_21565);
or U21774 (N_21774,N_21699,N_21627);
nor U21775 (N_21775,N_21742,N_21703);
and U21776 (N_21776,N_21712,N_21511);
nor U21777 (N_21777,N_21619,N_21538);
and U21778 (N_21778,N_21514,N_21659);
nor U21779 (N_21779,N_21679,N_21690);
or U21780 (N_21780,N_21544,N_21718);
nand U21781 (N_21781,N_21720,N_21631);
or U21782 (N_21782,N_21510,N_21691);
nor U21783 (N_21783,N_21589,N_21711);
nor U21784 (N_21784,N_21586,N_21705);
and U21785 (N_21785,N_21732,N_21525);
nor U21786 (N_21786,N_21724,N_21635);
nor U21787 (N_21787,N_21561,N_21656);
or U21788 (N_21788,N_21572,N_21682);
xor U21789 (N_21789,N_21694,N_21684);
or U21790 (N_21790,N_21529,N_21738);
or U21791 (N_21791,N_21504,N_21642);
and U21792 (N_21792,N_21536,N_21683);
xnor U21793 (N_21793,N_21747,N_21674);
xnor U21794 (N_21794,N_21606,N_21662);
and U21795 (N_21795,N_21734,N_21578);
or U21796 (N_21796,N_21693,N_21643);
nor U21797 (N_21797,N_21658,N_21706);
and U21798 (N_21798,N_21526,N_21558);
and U21799 (N_21799,N_21672,N_21573);
nor U21800 (N_21800,N_21723,N_21605);
nand U21801 (N_21801,N_21553,N_21700);
nand U21802 (N_21802,N_21600,N_21554);
or U21803 (N_21803,N_21519,N_21733);
or U21804 (N_21804,N_21516,N_21571);
nand U21805 (N_21805,N_21736,N_21505);
or U21806 (N_21806,N_21696,N_21522);
or U21807 (N_21807,N_21740,N_21574);
or U21808 (N_21808,N_21613,N_21598);
or U21809 (N_21809,N_21570,N_21649);
nor U21810 (N_21810,N_21681,N_21665);
nor U21811 (N_21811,N_21737,N_21534);
nand U21812 (N_21812,N_21585,N_21640);
and U21813 (N_21813,N_21587,N_21673);
nand U21814 (N_21814,N_21626,N_21533);
and U21815 (N_21815,N_21500,N_21654);
nand U21816 (N_21816,N_21715,N_21633);
nand U21817 (N_21817,N_21702,N_21618);
or U21818 (N_21818,N_21515,N_21729);
nand U21819 (N_21819,N_21588,N_21582);
or U21820 (N_21820,N_21678,N_21648);
or U21821 (N_21821,N_21548,N_21546);
and U21822 (N_21822,N_21677,N_21728);
nor U21823 (N_21823,N_21730,N_21695);
nand U21824 (N_21824,N_21727,N_21698);
xor U21825 (N_21825,N_21670,N_21562);
nor U21826 (N_21826,N_21506,N_21743);
nor U21827 (N_21827,N_21549,N_21594);
or U21828 (N_21828,N_21545,N_21601);
xnor U21829 (N_21829,N_21629,N_21527);
xnor U21830 (N_21830,N_21575,N_21559);
xnor U21831 (N_21831,N_21620,N_21731);
xnor U21832 (N_21832,N_21661,N_21638);
or U21833 (N_21833,N_21657,N_21688);
or U21834 (N_21834,N_21628,N_21653);
and U21835 (N_21835,N_21671,N_21584);
nor U21836 (N_21836,N_21701,N_21521);
or U21837 (N_21837,N_21719,N_21721);
nor U21838 (N_21838,N_21547,N_21577);
nor U21839 (N_21839,N_21741,N_21581);
and U21840 (N_21840,N_21707,N_21722);
nor U21841 (N_21841,N_21540,N_21713);
or U21842 (N_21842,N_21520,N_21660);
xor U21843 (N_21843,N_21602,N_21644);
nand U21844 (N_21844,N_21650,N_21517);
and U21845 (N_21845,N_21708,N_21615);
xor U21846 (N_21846,N_21676,N_21513);
or U21847 (N_21847,N_21608,N_21739);
nand U21848 (N_21848,N_21579,N_21609);
and U21849 (N_21849,N_21557,N_21614);
nand U21850 (N_21850,N_21622,N_21508);
xnor U21851 (N_21851,N_21610,N_21564);
nor U21852 (N_21852,N_21697,N_21704);
xnor U21853 (N_21853,N_21539,N_21596);
nor U21854 (N_21854,N_21590,N_21560);
and U21855 (N_21855,N_21501,N_21675);
and U21856 (N_21856,N_21744,N_21531);
and U21857 (N_21857,N_21535,N_21612);
or U21858 (N_21858,N_21593,N_21569);
and U21859 (N_21859,N_21599,N_21709);
nand U21860 (N_21860,N_21714,N_21576);
or U21861 (N_21861,N_21692,N_21639);
or U21862 (N_21862,N_21667,N_21749);
xor U21863 (N_21863,N_21551,N_21680);
nor U21864 (N_21864,N_21611,N_21543);
nor U21865 (N_21865,N_21592,N_21669);
or U21866 (N_21866,N_21616,N_21532);
nand U21867 (N_21867,N_21603,N_21617);
and U21868 (N_21868,N_21666,N_21664);
nor U21869 (N_21869,N_21552,N_21595);
nand U21870 (N_21870,N_21550,N_21634);
xnor U21871 (N_21871,N_21652,N_21717);
xnor U21872 (N_21872,N_21567,N_21583);
nor U21873 (N_21873,N_21530,N_21710);
nand U21874 (N_21874,N_21621,N_21502);
xnor U21875 (N_21875,N_21524,N_21542);
xnor U21876 (N_21876,N_21591,N_21582);
and U21877 (N_21877,N_21572,N_21652);
nand U21878 (N_21878,N_21500,N_21717);
xor U21879 (N_21879,N_21555,N_21558);
and U21880 (N_21880,N_21685,N_21691);
and U21881 (N_21881,N_21727,N_21537);
or U21882 (N_21882,N_21546,N_21714);
or U21883 (N_21883,N_21624,N_21517);
and U21884 (N_21884,N_21567,N_21599);
and U21885 (N_21885,N_21593,N_21607);
and U21886 (N_21886,N_21667,N_21717);
xor U21887 (N_21887,N_21703,N_21537);
and U21888 (N_21888,N_21513,N_21612);
nor U21889 (N_21889,N_21512,N_21597);
xnor U21890 (N_21890,N_21535,N_21714);
nand U21891 (N_21891,N_21600,N_21602);
and U21892 (N_21892,N_21734,N_21645);
or U21893 (N_21893,N_21554,N_21716);
or U21894 (N_21894,N_21615,N_21631);
nor U21895 (N_21895,N_21634,N_21553);
or U21896 (N_21896,N_21614,N_21654);
or U21897 (N_21897,N_21660,N_21548);
or U21898 (N_21898,N_21534,N_21560);
xor U21899 (N_21899,N_21737,N_21572);
or U21900 (N_21900,N_21538,N_21573);
or U21901 (N_21901,N_21703,N_21712);
and U21902 (N_21902,N_21526,N_21681);
and U21903 (N_21903,N_21677,N_21710);
and U21904 (N_21904,N_21724,N_21649);
xnor U21905 (N_21905,N_21655,N_21723);
nor U21906 (N_21906,N_21741,N_21533);
or U21907 (N_21907,N_21592,N_21615);
nand U21908 (N_21908,N_21590,N_21654);
or U21909 (N_21909,N_21564,N_21633);
or U21910 (N_21910,N_21604,N_21583);
or U21911 (N_21911,N_21605,N_21526);
nand U21912 (N_21912,N_21720,N_21661);
nand U21913 (N_21913,N_21700,N_21555);
or U21914 (N_21914,N_21599,N_21671);
xor U21915 (N_21915,N_21579,N_21575);
nand U21916 (N_21916,N_21567,N_21655);
nand U21917 (N_21917,N_21694,N_21653);
xor U21918 (N_21918,N_21501,N_21600);
xor U21919 (N_21919,N_21658,N_21716);
nor U21920 (N_21920,N_21532,N_21560);
nand U21921 (N_21921,N_21644,N_21615);
xnor U21922 (N_21922,N_21660,N_21565);
nand U21923 (N_21923,N_21670,N_21667);
xor U21924 (N_21924,N_21511,N_21587);
or U21925 (N_21925,N_21511,N_21698);
nand U21926 (N_21926,N_21738,N_21573);
and U21927 (N_21927,N_21622,N_21674);
xnor U21928 (N_21928,N_21729,N_21723);
nor U21929 (N_21929,N_21672,N_21663);
nor U21930 (N_21930,N_21599,N_21614);
nand U21931 (N_21931,N_21553,N_21612);
and U21932 (N_21932,N_21689,N_21541);
nand U21933 (N_21933,N_21676,N_21514);
nand U21934 (N_21934,N_21536,N_21622);
nand U21935 (N_21935,N_21679,N_21562);
nand U21936 (N_21936,N_21502,N_21513);
nand U21937 (N_21937,N_21736,N_21580);
or U21938 (N_21938,N_21500,N_21691);
nand U21939 (N_21939,N_21661,N_21657);
and U21940 (N_21940,N_21584,N_21507);
nand U21941 (N_21941,N_21543,N_21507);
xor U21942 (N_21942,N_21745,N_21636);
nand U21943 (N_21943,N_21731,N_21635);
nand U21944 (N_21944,N_21655,N_21603);
and U21945 (N_21945,N_21570,N_21635);
nand U21946 (N_21946,N_21533,N_21615);
and U21947 (N_21947,N_21551,N_21567);
nand U21948 (N_21948,N_21605,N_21721);
nor U21949 (N_21949,N_21556,N_21532);
or U21950 (N_21950,N_21579,N_21726);
and U21951 (N_21951,N_21506,N_21691);
xor U21952 (N_21952,N_21713,N_21550);
nor U21953 (N_21953,N_21554,N_21664);
nor U21954 (N_21954,N_21725,N_21591);
nand U21955 (N_21955,N_21711,N_21688);
and U21956 (N_21956,N_21589,N_21527);
and U21957 (N_21957,N_21634,N_21577);
or U21958 (N_21958,N_21529,N_21574);
xnor U21959 (N_21959,N_21518,N_21644);
or U21960 (N_21960,N_21566,N_21632);
xnor U21961 (N_21961,N_21636,N_21525);
nand U21962 (N_21962,N_21563,N_21646);
nand U21963 (N_21963,N_21695,N_21734);
and U21964 (N_21964,N_21589,N_21561);
nand U21965 (N_21965,N_21665,N_21565);
nor U21966 (N_21966,N_21525,N_21600);
xnor U21967 (N_21967,N_21556,N_21660);
or U21968 (N_21968,N_21593,N_21682);
and U21969 (N_21969,N_21706,N_21692);
and U21970 (N_21970,N_21614,N_21644);
xor U21971 (N_21971,N_21676,N_21593);
nor U21972 (N_21972,N_21563,N_21505);
or U21973 (N_21973,N_21525,N_21697);
and U21974 (N_21974,N_21679,N_21693);
xor U21975 (N_21975,N_21522,N_21741);
and U21976 (N_21976,N_21541,N_21620);
xor U21977 (N_21977,N_21741,N_21528);
nand U21978 (N_21978,N_21559,N_21692);
nand U21979 (N_21979,N_21573,N_21582);
xor U21980 (N_21980,N_21709,N_21560);
or U21981 (N_21981,N_21710,N_21570);
nand U21982 (N_21982,N_21618,N_21595);
nand U21983 (N_21983,N_21728,N_21695);
nor U21984 (N_21984,N_21740,N_21663);
and U21985 (N_21985,N_21651,N_21631);
nor U21986 (N_21986,N_21700,N_21552);
and U21987 (N_21987,N_21664,N_21691);
xnor U21988 (N_21988,N_21658,N_21518);
and U21989 (N_21989,N_21675,N_21523);
xnor U21990 (N_21990,N_21599,N_21714);
nor U21991 (N_21991,N_21697,N_21688);
nand U21992 (N_21992,N_21608,N_21614);
and U21993 (N_21993,N_21728,N_21731);
nand U21994 (N_21994,N_21709,N_21544);
nor U21995 (N_21995,N_21650,N_21672);
or U21996 (N_21996,N_21558,N_21568);
xor U21997 (N_21997,N_21717,N_21560);
and U21998 (N_21998,N_21590,N_21656);
xor U21999 (N_21999,N_21689,N_21592);
or U22000 (N_22000,N_21910,N_21780);
xnor U22001 (N_22001,N_21944,N_21924);
and U22002 (N_22002,N_21804,N_21820);
or U22003 (N_22003,N_21818,N_21759);
and U22004 (N_22004,N_21807,N_21872);
nor U22005 (N_22005,N_21840,N_21869);
and U22006 (N_22006,N_21873,N_21826);
xnor U22007 (N_22007,N_21880,N_21993);
or U22008 (N_22008,N_21850,N_21837);
nor U22009 (N_22009,N_21957,N_21927);
and U22010 (N_22010,N_21801,N_21981);
nor U22011 (N_22011,N_21829,N_21802);
nand U22012 (N_22012,N_21964,N_21750);
nand U22013 (N_22013,N_21943,N_21755);
or U22014 (N_22014,N_21805,N_21968);
and U22015 (N_22015,N_21799,N_21923);
nand U22016 (N_22016,N_21997,N_21996);
nor U22017 (N_22017,N_21941,N_21970);
xnor U22018 (N_22018,N_21868,N_21791);
nand U22019 (N_22019,N_21983,N_21835);
or U22020 (N_22020,N_21914,N_21764);
or U22021 (N_22021,N_21839,N_21925);
and U22022 (N_22022,N_21935,N_21803);
and U22023 (N_22023,N_21976,N_21768);
and U22024 (N_22024,N_21870,N_21784);
and U22025 (N_22025,N_21902,N_21949);
nor U22026 (N_22026,N_21999,N_21861);
xor U22027 (N_22027,N_21948,N_21953);
or U22028 (N_22028,N_21917,N_21849);
nand U22029 (N_22029,N_21796,N_21830);
nand U22030 (N_22030,N_21875,N_21906);
nor U22031 (N_22031,N_21758,N_21920);
nand U22032 (N_22032,N_21794,N_21913);
nor U22033 (N_22033,N_21915,N_21978);
nand U22034 (N_22034,N_21911,N_21961);
or U22035 (N_22035,N_21973,N_21940);
xnor U22036 (N_22036,N_21952,N_21825);
or U22037 (N_22037,N_21832,N_21761);
or U22038 (N_22038,N_21756,N_21762);
xnor U22039 (N_22039,N_21980,N_21918);
or U22040 (N_22040,N_21772,N_21956);
or U22041 (N_22041,N_21921,N_21937);
and U22042 (N_22042,N_21778,N_21848);
and U22043 (N_22043,N_21785,N_21857);
nor U22044 (N_22044,N_21786,N_21821);
xor U22045 (N_22045,N_21753,N_21995);
xnor U22046 (N_22046,N_21955,N_21890);
or U22047 (N_22047,N_21950,N_21893);
or U22048 (N_22048,N_21960,N_21774);
nor U22049 (N_22049,N_21843,N_21962);
or U22050 (N_22050,N_21754,N_21858);
xnor U22051 (N_22051,N_21757,N_21974);
nand U22052 (N_22052,N_21831,N_21930);
xor U22053 (N_22053,N_21847,N_21846);
or U22054 (N_22054,N_21884,N_21777);
nor U22055 (N_22055,N_21966,N_21787);
nor U22056 (N_22056,N_21933,N_21752);
nand U22057 (N_22057,N_21951,N_21864);
and U22058 (N_22058,N_21885,N_21853);
nand U22059 (N_22059,N_21977,N_21958);
and U22060 (N_22060,N_21767,N_21998);
nor U22061 (N_22061,N_21987,N_21844);
and U22062 (N_22062,N_21815,N_21919);
xnor U22063 (N_22063,N_21892,N_21789);
xnor U22064 (N_22064,N_21845,N_21770);
nor U22065 (N_22065,N_21990,N_21899);
xnor U22066 (N_22066,N_21771,N_21975);
xor U22067 (N_22067,N_21889,N_21866);
xnor U22068 (N_22068,N_21905,N_21903);
and U22069 (N_22069,N_21938,N_21841);
xnor U22070 (N_22070,N_21908,N_21793);
xor U22071 (N_22071,N_21863,N_21916);
xnor U22072 (N_22072,N_21854,N_21922);
or U22073 (N_22073,N_21898,N_21912);
or U22074 (N_22074,N_21945,N_21816);
xor U22075 (N_22075,N_21878,N_21986);
nand U22076 (N_22076,N_21751,N_21862);
nand U22077 (N_22077,N_21800,N_21891);
or U22078 (N_22078,N_21817,N_21763);
nand U22079 (N_22079,N_21814,N_21871);
nor U22080 (N_22080,N_21874,N_21808);
nand U22081 (N_22081,N_21887,N_21855);
nand U22082 (N_22082,N_21879,N_21946);
and U22083 (N_22083,N_21901,N_21809);
nand U22084 (N_22084,N_21982,N_21969);
and U22085 (N_22085,N_21783,N_21994);
xor U22086 (N_22086,N_21888,N_21904);
or U22087 (N_22087,N_21876,N_21954);
nor U22088 (N_22088,N_21907,N_21828);
and U22089 (N_22089,N_21965,N_21932);
xnor U22090 (N_22090,N_21824,N_21811);
nor U22091 (N_22091,N_21896,N_21991);
or U22092 (N_22092,N_21838,N_21909);
and U22093 (N_22093,N_21867,N_21959);
and U22094 (N_22094,N_21782,N_21775);
xor U22095 (N_22095,N_21963,N_21779);
xor U22096 (N_22096,N_21886,N_21860);
nand U22097 (N_22097,N_21842,N_21947);
xnor U22098 (N_22098,N_21926,N_21971);
or U22099 (N_22099,N_21967,N_21931);
and U22100 (N_22100,N_21834,N_21984);
nor U22101 (N_22101,N_21900,N_21788);
nand U22102 (N_22102,N_21765,N_21836);
or U22103 (N_22103,N_21942,N_21851);
nand U22104 (N_22104,N_21792,N_21822);
xor U22105 (N_22105,N_21883,N_21856);
or U22106 (N_22106,N_21810,N_21939);
xor U22107 (N_22107,N_21895,N_21766);
nand U22108 (N_22108,N_21806,N_21979);
nand U22109 (N_22109,N_21776,N_21769);
nand U22110 (N_22110,N_21833,N_21773);
nand U22111 (N_22111,N_21819,N_21936);
xor U22112 (N_22112,N_21985,N_21760);
or U22113 (N_22113,N_21798,N_21781);
or U22114 (N_22114,N_21882,N_21812);
and U22115 (N_22115,N_21934,N_21897);
and U22116 (N_22116,N_21827,N_21988);
nand U22117 (N_22117,N_21797,N_21852);
and U22118 (N_22118,N_21790,N_21972);
and U22119 (N_22119,N_21813,N_21823);
xor U22120 (N_22120,N_21795,N_21989);
xor U22121 (N_22121,N_21877,N_21992);
and U22122 (N_22122,N_21865,N_21859);
nor U22123 (N_22123,N_21928,N_21894);
nand U22124 (N_22124,N_21881,N_21929);
and U22125 (N_22125,N_21873,N_21776);
xor U22126 (N_22126,N_21802,N_21995);
xor U22127 (N_22127,N_21924,N_21970);
or U22128 (N_22128,N_21763,N_21951);
nor U22129 (N_22129,N_21914,N_21918);
or U22130 (N_22130,N_21917,N_21876);
and U22131 (N_22131,N_21844,N_21809);
nand U22132 (N_22132,N_21981,N_21933);
and U22133 (N_22133,N_21993,N_21868);
nor U22134 (N_22134,N_21751,N_21852);
or U22135 (N_22135,N_21938,N_21845);
xnor U22136 (N_22136,N_21776,N_21846);
xnor U22137 (N_22137,N_21947,N_21770);
or U22138 (N_22138,N_21816,N_21869);
nand U22139 (N_22139,N_21821,N_21764);
and U22140 (N_22140,N_21799,N_21891);
or U22141 (N_22141,N_21773,N_21835);
xor U22142 (N_22142,N_21808,N_21930);
or U22143 (N_22143,N_21773,N_21969);
and U22144 (N_22144,N_21983,N_21898);
and U22145 (N_22145,N_21931,N_21982);
nand U22146 (N_22146,N_21785,N_21803);
or U22147 (N_22147,N_21902,N_21808);
or U22148 (N_22148,N_21927,N_21971);
or U22149 (N_22149,N_21781,N_21939);
and U22150 (N_22150,N_21974,N_21835);
xnor U22151 (N_22151,N_21751,N_21830);
nor U22152 (N_22152,N_21852,N_21942);
xnor U22153 (N_22153,N_21948,N_21913);
or U22154 (N_22154,N_21869,N_21836);
nand U22155 (N_22155,N_21982,N_21759);
nand U22156 (N_22156,N_21973,N_21789);
and U22157 (N_22157,N_21845,N_21826);
or U22158 (N_22158,N_21755,N_21855);
xor U22159 (N_22159,N_21921,N_21777);
nand U22160 (N_22160,N_21982,N_21868);
xnor U22161 (N_22161,N_21812,N_21821);
xnor U22162 (N_22162,N_21851,N_21971);
and U22163 (N_22163,N_21892,N_21906);
or U22164 (N_22164,N_21804,N_21874);
nand U22165 (N_22165,N_21953,N_21989);
xnor U22166 (N_22166,N_21985,N_21814);
and U22167 (N_22167,N_21968,N_21822);
or U22168 (N_22168,N_21881,N_21810);
nand U22169 (N_22169,N_21839,N_21805);
and U22170 (N_22170,N_21911,N_21950);
and U22171 (N_22171,N_21942,N_21932);
nand U22172 (N_22172,N_21771,N_21848);
and U22173 (N_22173,N_21966,N_21937);
and U22174 (N_22174,N_21872,N_21831);
or U22175 (N_22175,N_21969,N_21915);
and U22176 (N_22176,N_21873,N_21760);
nand U22177 (N_22177,N_21954,N_21780);
nand U22178 (N_22178,N_21903,N_21931);
or U22179 (N_22179,N_21766,N_21757);
nand U22180 (N_22180,N_21762,N_21873);
xnor U22181 (N_22181,N_21930,N_21980);
nand U22182 (N_22182,N_21998,N_21964);
and U22183 (N_22183,N_21866,N_21921);
nand U22184 (N_22184,N_21876,N_21932);
xnor U22185 (N_22185,N_21890,N_21772);
nor U22186 (N_22186,N_21867,N_21914);
xnor U22187 (N_22187,N_21772,N_21925);
or U22188 (N_22188,N_21996,N_21823);
nor U22189 (N_22189,N_21865,N_21897);
and U22190 (N_22190,N_21874,N_21841);
nand U22191 (N_22191,N_21821,N_21755);
or U22192 (N_22192,N_21862,N_21758);
nor U22193 (N_22193,N_21869,N_21901);
nor U22194 (N_22194,N_21772,N_21833);
xnor U22195 (N_22195,N_21770,N_21922);
nand U22196 (N_22196,N_21974,N_21776);
or U22197 (N_22197,N_21934,N_21863);
xor U22198 (N_22198,N_21871,N_21953);
or U22199 (N_22199,N_21925,N_21903);
or U22200 (N_22200,N_21773,N_21923);
xor U22201 (N_22201,N_21915,N_21846);
and U22202 (N_22202,N_21965,N_21948);
xor U22203 (N_22203,N_21765,N_21989);
nand U22204 (N_22204,N_21970,N_21905);
and U22205 (N_22205,N_21901,N_21885);
and U22206 (N_22206,N_21760,N_21859);
and U22207 (N_22207,N_21771,N_21834);
nand U22208 (N_22208,N_21848,N_21776);
and U22209 (N_22209,N_21756,N_21936);
or U22210 (N_22210,N_21881,N_21839);
and U22211 (N_22211,N_21830,N_21801);
nor U22212 (N_22212,N_21909,N_21921);
nor U22213 (N_22213,N_21894,N_21883);
and U22214 (N_22214,N_21910,N_21973);
or U22215 (N_22215,N_21906,N_21784);
nor U22216 (N_22216,N_21803,N_21847);
xnor U22217 (N_22217,N_21981,N_21923);
nor U22218 (N_22218,N_21843,N_21766);
and U22219 (N_22219,N_21975,N_21902);
nand U22220 (N_22220,N_21760,N_21836);
xor U22221 (N_22221,N_21989,N_21778);
or U22222 (N_22222,N_21865,N_21835);
xor U22223 (N_22223,N_21875,N_21973);
nor U22224 (N_22224,N_21764,N_21753);
and U22225 (N_22225,N_21903,N_21855);
or U22226 (N_22226,N_21956,N_21901);
nand U22227 (N_22227,N_21868,N_21884);
nand U22228 (N_22228,N_21977,N_21823);
or U22229 (N_22229,N_21967,N_21906);
or U22230 (N_22230,N_21798,N_21896);
and U22231 (N_22231,N_21767,N_21781);
or U22232 (N_22232,N_21875,N_21760);
xnor U22233 (N_22233,N_21880,N_21904);
or U22234 (N_22234,N_21990,N_21808);
nand U22235 (N_22235,N_21934,N_21762);
nand U22236 (N_22236,N_21793,N_21969);
and U22237 (N_22237,N_21767,N_21870);
or U22238 (N_22238,N_21979,N_21788);
xnor U22239 (N_22239,N_21791,N_21975);
xnor U22240 (N_22240,N_21847,N_21804);
nor U22241 (N_22241,N_21987,N_21865);
and U22242 (N_22242,N_21968,N_21760);
xnor U22243 (N_22243,N_21910,N_21766);
nor U22244 (N_22244,N_21879,N_21923);
nand U22245 (N_22245,N_21755,N_21976);
xnor U22246 (N_22246,N_21949,N_21953);
or U22247 (N_22247,N_21878,N_21808);
or U22248 (N_22248,N_21859,N_21976);
or U22249 (N_22249,N_21971,N_21916);
or U22250 (N_22250,N_22228,N_22229);
nand U22251 (N_22251,N_22111,N_22224);
and U22252 (N_22252,N_22012,N_22219);
xor U22253 (N_22253,N_22011,N_22089);
xor U22254 (N_22254,N_22069,N_22146);
nor U22255 (N_22255,N_22106,N_22031);
xnor U22256 (N_22256,N_22183,N_22223);
nor U22257 (N_22257,N_22195,N_22241);
or U22258 (N_22258,N_22201,N_22074);
nand U22259 (N_22259,N_22249,N_22129);
nor U22260 (N_22260,N_22084,N_22088);
nand U22261 (N_22261,N_22016,N_22049);
nor U22262 (N_22262,N_22046,N_22076);
or U22263 (N_22263,N_22007,N_22145);
or U22264 (N_22264,N_22123,N_22110);
xor U22265 (N_22265,N_22169,N_22151);
nor U22266 (N_22266,N_22214,N_22130);
nand U22267 (N_22267,N_22018,N_22198);
or U22268 (N_22268,N_22148,N_22064);
nor U22269 (N_22269,N_22230,N_22149);
or U22270 (N_22270,N_22248,N_22003);
or U22271 (N_22271,N_22209,N_22190);
xnor U22272 (N_22272,N_22188,N_22085);
or U22273 (N_22273,N_22070,N_22143);
or U22274 (N_22274,N_22171,N_22033);
or U22275 (N_22275,N_22039,N_22023);
and U22276 (N_22276,N_22166,N_22178);
or U22277 (N_22277,N_22222,N_22164);
nor U22278 (N_22278,N_22212,N_22179);
nor U22279 (N_22279,N_22014,N_22105);
nor U22280 (N_22280,N_22004,N_22058);
nand U22281 (N_22281,N_22155,N_22133);
xor U22282 (N_22282,N_22002,N_22211);
nor U22283 (N_22283,N_22109,N_22138);
nand U22284 (N_22284,N_22062,N_22194);
or U22285 (N_22285,N_22090,N_22135);
nor U22286 (N_22286,N_22218,N_22035);
or U22287 (N_22287,N_22186,N_22025);
nor U22288 (N_22288,N_22047,N_22187);
and U22289 (N_22289,N_22142,N_22118);
nor U22290 (N_22290,N_22041,N_22108);
nor U22291 (N_22291,N_22100,N_22122);
xnor U22292 (N_22292,N_22125,N_22052);
or U22293 (N_22293,N_22097,N_22066);
or U22294 (N_22294,N_22128,N_22013);
or U22295 (N_22295,N_22227,N_22192);
and U22296 (N_22296,N_22063,N_22020);
xnor U22297 (N_22297,N_22235,N_22030);
or U22298 (N_22298,N_22029,N_22068);
nor U22299 (N_22299,N_22156,N_22231);
nor U22300 (N_22300,N_22044,N_22082);
nor U22301 (N_22301,N_22057,N_22104);
xnor U22302 (N_22302,N_22072,N_22115);
and U22303 (N_22303,N_22036,N_22180);
and U22304 (N_22304,N_22134,N_22000);
nand U22305 (N_22305,N_22061,N_22019);
and U22306 (N_22306,N_22139,N_22026);
nor U22307 (N_22307,N_22197,N_22060);
nor U22308 (N_22308,N_22159,N_22199);
nor U22309 (N_22309,N_22017,N_22073);
and U22310 (N_22310,N_22167,N_22079);
nand U22311 (N_22311,N_22099,N_22213);
nand U22312 (N_22312,N_22120,N_22216);
nor U22313 (N_22313,N_22181,N_22132);
or U22314 (N_22314,N_22038,N_22098);
nor U22315 (N_22315,N_22027,N_22127);
or U22316 (N_22316,N_22050,N_22095);
nand U22317 (N_22317,N_22237,N_22246);
xor U22318 (N_22318,N_22021,N_22131);
nor U22319 (N_22319,N_22045,N_22147);
nand U22320 (N_22320,N_22206,N_22144);
or U22321 (N_22321,N_22236,N_22006);
nor U22322 (N_22322,N_22185,N_22140);
or U22323 (N_22323,N_22232,N_22163);
or U22324 (N_22324,N_22210,N_22081);
nand U22325 (N_22325,N_22056,N_22240);
nand U22326 (N_22326,N_22177,N_22165);
and U22327 (N_22327,N_22078,N_22215);
and U22328 (N_22328,N_22225,N_22153);
nand U22329 (N_22329,N_22009,N_22043);
and U22330 (N_22330,N_22154,N_22170);
and U22331 (N_22331,N_22032,N_22042);
or U22332 (N_22332,N_22168,N_22244);
or U22333 (N_22333,N_22234,N_22126);
nor U22334 (N_22334,N_22028,N_22051);
and U22335 (N_22335,N_22184,N_22182);
or U22336 (N_22336,N_22161,N_22055);
or U22337 (N_22337,N_22096,N_22034);
nor U22338 (N_22338,N_22217,N_22191);
nor U22339 (N_22339,N_22087,N_22233);
xor U22340 (N_22340,N_22117,N_22238);
xor U22341 (N_22341,N_22173,N_22102);
xnor U22342 (N_22342,N_22220,N_22008);
nand U22343 (N_22343,N_22086,N_22136);
xor U22344 (N_22344,N_22152,N_22037);
xor U22345 (N_22345,N_22243,N_22137);
nor U22346 (N_22346,N_22162,N_22107);
xnor U22347 (N_22347,N_22205,N_22114);
xor U22348 (N_22348,N_22158,N_22176);
or U22349 (N_22349,N_22077,N_22121);
nor U22350 (N_22350,N_22015,N_22174);
xnor U22351 (N_22351,N_22101,N_22172);
nor U22352 (N_22352,N_22080,N_22160);
nor U22353 (N_22353,N_22150,N_22094);
or U22354 (N_22354,N_22059,N_22048);
xnor U22355 (N_22355,N_22221,N_22053);
nand U22356 (N_22356,N_22207,N_22091);
or U22357 (N_22357,N_22247,N_22001);
nand U22358 (N_22358,N_22203,N_22065);
xnor U22359 (N_22359,N_22092,N_22196);
or U22360 (N_22360,N_22239,N_22189);
nor U22361 (N_22361,N_22141,N_22226);
and U22362 (N_22362,N_22175,N_22093);
xnor U22363 (N_22363,N_22202,N_22113);
nor U22364 (N_22364,N_22005,N_22024);
xor U22365 (N_22365,N_22067,N_22075);
nand U22366 (N_22366,N_22157,N_22124);
or U22367 (N_22367,N_22054,N_22208);
nand U22368 (N_22368,N_22083,N_22116);
and U22369 (N_22369,N_22103,N_22200);
and U22370 (N_22370,N_22119,N_22022);
or U22371 (N_22371,N_22242,N_22071);
xor U22372 (N_22372,N_22010,N_22040);
nand U22373 (N_22373,N_22245,N_22193);
xnor U22374 (N_22374,N_22204,N_22112);
nor U22375 (N_22375,N_22178,N_22050);
or U22376 (N_22376,N_22192,N_22167);
nor U22377 (N_22377,N_22246,N_22050);
and U22378 (N_22378,N_22171,N_22191);
or U22379 (N_22379,N_22065,N_22011);
and U22380 (N_22380,N_22221,N_22040);
and U22381 (N_22381,N_22148,N_22013);
and U22382 (N_22382,N_22077,N_22081);
and U22383 (N_22383,N_22187,N_22128);
nand U22384 (N_22384,N_22175,N_22010);
nor U22385 (N_22385,N_22193,N_22000);
nor U22386 (N_22386,N_22143,N_22227);
or U22387 (N_22387,N_22139,N_22186);
xnor U22388 (N_22388,N_22133,N_22008);
xnor U22389 (N_22389,N_22177,N_22145);
nor U22390 (N_22390,N_22110,N_22199);
nand U22391 (N_22391,N_22122,N_22079);
nand U22392 (N_22392,N_22061,N_22185);
nor U22393 (N_22393,N_22224,N_22225);
nor U22394 (N_22394,N_22012,N_22115);
nor U22395 (N_22395,N_22132,N_22058);
or U22396 (N_22396,N_22053,N_22190);
nand U22397 (N_22397,N_22242,N_22185);
nand U22398 (N_22398,N_22161,N_22050);
nand U22399 (N_22399,N_22028,N_22040);
nor U22400 (N_22400,N_22188,N_22183);
and U22401 (N_22401,N_22145,N_22242);
xor U22402 (N_22402,N_22158,N_22127);
nor U22403 (N_22403,N_22120,N_22036);
nand U22404 (N_22404,N_22109,N_22211);
nand U22405 (N_22405,N_22232,N_22075);
and U22406 (N_22406,N_22139,N_22218);
or U22407 (N_22407,N_22147,N_22231);
nor U22408 (N_22408,N_22239,N_22064);
xor U22409 (N_22409,N_22059,N_22087);
or U22410 (N_22410,N_22243,N_22065);
or U22411 (N_22411,N_22155,N_22026);
xnor U22412 (N_22412,N_22088,N_22196);
xnor U22413 (N_22413,N_22080,N_22123);
or U22414 (N_22414,N_22167,N_22088);
xnor U22415 (N_22415,N_22159,N_22226);
nand U22416 (N_22416,N_22153,N_22197);
nand U22417 (N_22417,N_22140,N_22000);
or U22418 (N_22418,N_22008,N_22004);
or U22419 (N_22419,N_22057,N_22247);
and U22420 (N_22420,N_22018,N_22151);
nor U22421 (N_22421,N_22228,N_22191);
and U22422 (N_22422,N_22012,N_22122);
xnor U22423 (N_22423,N_22204,N_22106);
nand U22424 (N_22424,N_22147,N_22126);
nand U22425 (N_22425,N_22092,N_22225);
nand U22426 (N_22426,N_22069,N_22169);
xnor U22427 (N_22427,N_22031,N_22058);
and U22428 (N_22428,N_22242,N_22234);
and U22429 (N_22429,N_22092,N_22203);
and U22430 (N_22430,N_22174,N_22061);
xnor U22431 (N_22431,N_22167,N_22076);
and U22432 (N_22432,N_22171,N_22153);
nor U22433 (N_22433,N_22063,N_22090);
nand U22434 (N_22434,N_22043,N_22218);
nor U22435 (N_22435,N_22119,N_22067);
xnor U22436 (N_22436,N_22234,N_22082);
and U22437 (N_22437,N_22233,N_22010);
and U22438 (N_22438,N_22207,N_22027);
and U22439 (N_22439,N_22061,N_22156);
nand U22440 (N_22440,N_22156,N_22203);
and U22441 (N_22441,N_22039,N_22133);
nand U22442 (N_22442,N_22241,N_22116);
or U22443 (N_22443,N_22219,N_22141);
xnor U22444 (N_22444,N_22201,N_22005);
nor U22445 (N_22445,N_22234,N_22190);
and U22446 (N_22446,N_22006,N_22178);
or U22447 (N_22447,N_22041,N_22027);
nor U22448 (N_22448,N_22205,N_22162);
xor U22449 (N_22449,N_22148,N_22238);
or U22450 (N_22450,N_22200,N_22113);
and U22451 (N_22451,N_22093,N_22220);
or U22452 (N_22452,N_22109,N_22208);
or U22453 (N_22453,N_22209,N_22041);
or U22454 (N_22454,N_22166,N_22157);
nand U22455 (N_22455,N_22230,N_22093);
nand U22456 (N_22456,N_22080,N_22147);
xor U22457 (N_22457,N_22225,N_22082);
xnor U22458 (N_22458,N_22071,N_22094);
or U22459 (N_22459,N_22056,N_22120);
nor U22460 (N_22460,N_22034,N_22208);
or U22461 (N_22461,N_22166,N_22043);
and U22462 (N_22462,N_22194,N_22000);
nor U22463 (N_22463,N_22032,N_22020);
or U22464 (N_22464,N_22217,N_22160);
nand U22465 (N_22465,N_22244,N_22068);
nor U22466 (N_22466,N_22227,N_22061);
xor U22467 (N_22467,N_22142,N_22219);
nand U22468 (N_22468,N_22224,N_22119);
nor U22469 (N_22469,N_22217,N_22248);
nor U22470 (N_22470,N_22103,N_22184);
xnor U22471 (N_22471,N_22173,N_22001);
xor U22472 (N_22472,N_22167,N_22224);
xor U22473 (N_22473,N_22164,N_22211);
nand U22474 (N_22474,N_22003,N_22229);
and U22475 (N_22475,N_22080,N_22007);
nand U22476 (N_22476,N_22050,N_22075);
nor U22477 (N_22477,N_22017,N_22164);
nand U22478 (N_22478,N_22175,N_22191);
nand U22479 (N_22479,N_22067,N_22080);
nor U22480 (N_22480,N_22004,N_22221);
or U22481 (N_22481,N_22080,N_22201);
and U22482 (N_22482,N_22182,N_22025);
or U22483 (N_22483,N_22166,N_22134);
xor U22484 (N_22484,N_22121,N_22081);
or U22485 (N_22485,N_22025,N_22055);
and U22486 (N_22486,N_22023,N_22056);
and U22487 (N_22487,N_22095,N_22245);
nor U22488 (N_22488,N_22072,N_22031);
nand U22489 (N_22489,N_22188,N_22028);
nand U22490 (N_22490,N_22060,N_22175);
or U22491 (N_22491,N_22168,N_22158);
or U22492 (N_22492,N_22156,N_22143);
nand U22493 (N_22493,N_22124,N_22035);
or U22494 (N_22494,N_22189,N_22207);
and U22495 (N_22495,N_22018,N_22245);
nor U22496 (N_22496,N_22094,N_22197);
xor U22497 (N_22497,N_22112,N_22051);
nand U22498 (N_22498,N_22120,N_22163);
or U22499 (N_22499,N_22123,N_22169);
xor U22500 (N_22500,N_22312,N_22363);
nor U22501 (N_22501,N_22497,N_22292);
nand U22502 (N_22502,N_22260,N_22337);
and U22503 (N_22503,N_22380,N_22448);
and U22504 (N_22504,N_22279,N_22254);
nand U22505 (N_22505,N_22457,N_22320);
nand U22506 (N_22506,N_22371,N_22397);
or U22507 (N_22507,N_22314,N_22496);
nor U22508 (N_22508,N_22435,N_22444);
nor U22509 (N_22509,N_22338,N_22470);
xor U22510 (N_22510,N_22465,N_22437);
nor U22511 (N_22511,N_22381,N_22491);
nand U22512 (N_22512,N_22340,N_22336);
and U22513 (N_22513,N_22353,N_22460);
nor U22514 (N_22514,N_22446,N_22481);
nor U22515 (N_22515,N_22480,N_22390);
and U22516 (N_22516,N_22451,N_22351);
xnor U22517 (N_22517,N_22373,N_22447);
nand U22518 (N_22518,N_22303,N_22492);
nand U22519 (N_22519,N_22328,N_22360);
nand U22520 (N_22520,N_22331,N_22479);
xnor U22521 (N_22521,N_22384,N_22277);
nor U22522 (N_22522,N_22493,N_22294);
nor U22523 (N_22523,N_22472,N_22450);
nor U22524 (N_22524,N_22458,N_22339);
nand U22525 (N_22525,N_22443,N_22302);
and U22526 (N_22526,N_22290,N_22454);
and U22527 (N_22527,N_22396,N_22282);
nor U22528 (N_22528,N_22421,N_22250);
xor U22529 (N_22529,N_22318,N_22357);
nor U22530 (N_22530,N_22256,N_22386);
and U22531 (N_22531,N_22334,N_22436);
and U22532 (N_22532,N_22317,N_22273);
xor U22533 (N_22533,N_22494,N_22335);
xor U22534 (N_22534,N_22410,N_22274);
or U22535 (N_22535,N_22284,N_22482);
or U22536 (N_22536,N_22316,N_22322);
nor U22537 (N_22537,N_22356,N_22286);
xor U22538 (N_22538,N_22442,N_22392);
and U22539 (N_22539,N_22252,N_22375);
nand U22540 (N_22540,N_22389,N_22283);
or U22541 (N_22541,N_22441,N_22306);
and U22542 (N_22542,N_22321,N_22427);
nand U22543 (N_22543,N_22330,N_22367);
nor U22544 (N_22544,N_22404,N_22364);
xnor U22545 (N_22545,N_22478,N_22341);
and U22546 (N_22546,N_22269,N_22378);
or U22547 (N_22547,N_22295,N_22313);
nor U22548 (N_22548,N_22434,N_22382);
and U22549 (N_22549,N_22453,N_22455);
or U22550 (N_22550,N_22326,N_22432);
and U22551 (N_22551,N_22297,N_22253);
xor U22552 (N_22552,N_22325,N_22296);
nand U22553 (N_22553,N_22474,N_22307);
and U22554 (N_22554,N_22411,N_22275);
xnor U22555 (N_22555,N_22301,N_22405);
nand U22556 (N_22556,N_22468,N_22426);
nand U22557 (N_22557,N_22452,N_22299);
or U22558 (N_22558,N_22323,N_22399);
nand U22559 (N_22559,N_22311,N_22489);
or U22560 (N_22560,N_22430,N_22477);
or U22561 (N_22561,N_22305,N_22343);
nand U22562 (N_22562,N_22422,N_22308);
or U22563 (N_22563,N_22475,N_22464);
xor U22564 (N_22564,N_22369,N_22476);
or U22565 (N_22565,N_22355,N_22419);
and U22566 (N_22566,N_22485,N_22300);
nor U22567 (N_22567,N_22406,N_22488);
nor U22568 (N_22568,N_22361,N_22459);
nor U22569 (N_22569,N_22346,N_22319);
nor U22570 (N_22570,N_22387,N_22264);
nor U22571 (N_22571,N_22445,N_22379);
xor U22572 (N_22572,N_22262,N_22349);
and U22573 (N_22573,N_22267,N_22259);
xnor U22574 (N_22574,N_22281,N_22394);
and U22575 (N_22575,N_22354,N_22398);
and U22576 (N_22576,N_22388,N_22439);
and U22577 (N_22577,N_22347,N_22414);
and U22578 (N_22578,N_22377,N_22462);
nor U22579 (N_22579,N_22418,N_22383);
nand U22580 (N_22580,N_22350,N_22374);
nand U22581 (N_22581,N_22272,N_22431);
xor U22582 (N_22582,N_22467,N_22304);
and U22583 (N_22583,N_22490,N_22288);
and U22584 (N_22584,N_22393,N_22420);
or U22585 (N_22585,N_22401,N_22263);
nand U22586 (N_22586,N_22428,N_22310);
or U22587 (N_22587,N_22348,N_22332);
nand U22588 (N_22588,N_22329,N_22495);
xnor U22589 (N_22589,N_22425,N_22287);
nor U22590 (N_22590,N_22473,N_22449);
and U22591 (N_22591,N_22423,N_22469);
and U22592 (N_22592,N_22293,N_22483);
and U22593 (N_22593,N_22342,N_22461);
xnor U22594 (N_22594,N_22424,N_22324);
xor U22595 (N_22595,N_22433,N_22266);
xor U22596 (N_22596,N_22278,N_22285);
nand U22597 (N_22597,N_22370,N_22368);
and U22598 (N_22598,N_22289,N_22413);
and U22599 (N_22599,N_22408,N_22471);
and U22600 (N_22600,N_22395,N_22499);
and U22601 (N_22601,N_22352,N_22280);
nand U22602 (N_22602,N_22417,N_22359);
and U22603 (N_22603,N_22271,N_22484);
nand U22604 (N_22604,N_22416,N_22372);
or U22605 (N_22605,N_22440,N_22315);
or U22606 (N_22606,N_22255,N_22400);
and U22607 (N_22607,N_22276,N_22463);
and U22608 (N_22608,N_22366,N_22402);
xor U22609 (N_22609,N_22265,N_22415);
or U22610 (N_22610,N_22327,N_22407);
xnor U22611 (N_22611,N_22466,N_22251);
xor U22612 (N_22612,N_22456,N_22412);
and U22613 (N_22613,N_22486,N_22291);
xor U22614 (N_22614,N_22391,N_22362);
and U22615 (N_22615,N_22358,N_22498);
nand U22616 (N_22616,N_22385,N_22298);
or U22617 (N_22617,N_22268,N_22257);
nor U22618 (N_22618,N_22429,N_22365);
nand U22619 (N_22619,N_22261,N_22487);
or U22620 (N_22620,N_22376,N_22270);
and U22621 (N_22621,N_22344,N_22409);
and U22622 (N_22622,N_22403,N_22333);
nand U22623 (N_22623,N_22309,N_22438);
nand U22624 (N_22624,N_22258,N_22345);
and U22625 (N_22625,N_22297,N_22497);
xnor U22626 (N_22626,N_22359,N_22262);
and U22627 (N_22627,N_22405,N_22311);
xnor U22628 (N_22628,N_22395,N_22453);
xor U22629 (N_22629,N_22437,N_22336);
nor U22630 (N_22630,N_22348,N_22499);
or U22631 (N_22631,N_22272,N_22462);
nand U22632 (N_22632,N_22424,N_22360);
nor U22633 (N_22633,N_22301,N_22285);
xor U22634 (N_22634,N_22442,N_22277);
xor U22635 (N_22635,N_22298,N_22299);
xnor U22636 (N_22636,N_22374,N_22346);
nand U22637 (N_22637,N_22418,N_22414);
nand U22638 (N_22638,N_22252,N_22433);
nand U22639 (N_22639,N_22251,N_22484);
nor U22640 (N_22640,N_22425,N_22420);
or U22641 (N_22641,N_22330,N_22491);
nand U22642 (N_22642,N_22342,N_22331);
nor U22643 (N_22643,N_22375,N_22381);
and U22644 (N_22644,N_22253,N_22324);
xnor U22645 (N_22645,N_22412,N_22292);
nor U22646 (N_22646,N_22437,N_22312);
nand U22647 (N_22647,N_22348,N_22441);
and U22648 (N_22648,N_22332,N_22450);
nand U22649 (N_22649,N_22460,N_22427);
nand U22650 (N_22650,N_22425,N_22380);
and U22651 (N_22651,N_22372,N_22389);
or U22652 (N_22652,N_22471,N_22356);
or U22653 (N_22653,N_22278,N_22308);
xnor U22654 (N_22654,N_22443,N_22345);
nor U22655 (N_22655,N_22283,N_22345);
and U22656 (N_22656,N_22352,N_22369);
xnor U22657 (N_22657,N_22325,N_22302);
xnor U22658 (N_22658,N_22416,N_22355);
and U22659 (N_22659,N_22319,N_22266);
nor U22660 (N_22660,N_22329,N_22487);
xor U22661 (N_22661,N_22287,N_22305);
nor U22662 (N_22662,N_22395,N_22416);
nand U22663 (N_22663,N_22331,N_22445);
xnor U22664 (N_22664,N_22479,N_22472);
nand U22665 (N_22665,N_22264,N_22478);
and U22666 (N_22666,N_22259,N_22461);
xnor U22667 (N_22667,N_22272,N_22252);
or U22668 (N_22668,N_22293,N_22414);
nand U22669 (N_22669,N_22445,N_22465);
and U22670 (N_22670,N_22417,N_22464);
nor U22671 (N_22671,N_22316,N_22278);
nor U22672 (N_22672,N_22313,N_22391);
or U22673 (N_22673,N_22374,N_22464);
or U22674 (N_22674,N_22398,N_22428);
or U22675 (N_22675,N_22408,N_22484);
nor U22676 (N_22676,N_22306,N_22290);
nand U22677 (N_22677,N_22255,N_22495);
or U22678 (N_22678,N_22490,N_22381);
nor U22679 (N_22679,N_22331,N_22471);
nand U22680 (N_22680,N_22492,N_22250);
nand U22681 (N_22681,N_22337,N_22302);
nor U22682 (N_22682,N_22466,N_22340);
or U22683 (N_22683,N_22271,N_22409);
xnor U22684 (N_22684,N_22423,N_22305);
nand U22685 (N_22685,N_22393,N_22284);
or U22686 (N_22686,N_22348,N_22284);
or U22687 (N_22687,N_22321,N_22328);
or U22688 (N_22688,N_22459,N_22468);
nor U22689 (N_22689,N_22299,N_22407);
nand U22690 (N_22690,N_22329,N_22403);
and U22691 (N_22691,N_22381,N_22447);
nor U22692 (N_22692,N_22362,N_22430);
and U22693 (N_22693,N_22459,N_22397);
or U22694 (N_22694,N_22400,N_22288);
xor U22695 (N_22695,N_22391,N_22488);
or U22696 (N_22696,N_22489,N_22280);
and U22697 (N_22697,N_22282,N_22444);
nor U22698 (N_22698,N_22468,N_22327);
or U22699 (N_22699,N_22319,N_22328);
or U22700 (N_22700,N_22280,N_22426);
or U22701 (N_22701,N_22263,N_22370);
nand U22702 (N_22702,N_22419,N_22279);
nor U22703 (N_22703,N_22342,N_22270);
or U22704 (N_22704,N_22321,N_22266);
or U22705 (N_22705,N_22358,N_22270);
nor U22706 (N_22706,N_22351,N_22423);
nor U22707 (N_22707,N_22322,N_22430);
nor U22708 (N_22708,N_22463,N_22364);
and U22709 (N_22709,N_22297,N_22471);
and U22710 (N_22710,N_22266,N_22459);
nor U22711 (N_22711,N_22395,N_22463);
nor U22712 (N_22712,N_22306,N_22303);
or U22713 (N_22713,N_22485,N_22438);
xnor U22714 (N_22714,N_22303,N_22429);
nor U22715 (N_22715,N_22278,N_22464);
nand U22716 (N_22716,N_22453,N_22353);
xnor U22717 (N_22717,N_22358,N_22323);
xnor U22718 (N_22718,N_22450,N_22308);
nor U22719 (N_22719,N_22337,N_22410);
xnor U22720 (N_22720,N_22369,N_22370);
xor U22721 (N_22721,N_22304,N_22365);
nor U22722 (N_22722,N_22350,N_22259);
nor U22723 (N_22723,N_22461,N_22356);
xnor U22724 (N_22724,N_22383,N_22279);
nor U22725 (N_22725,N_22342,N_22478);
nand U22726 (N_22726,N_22341,N_22303);
xor U22727 (N_22727,N_22372,N_22456);
xnor U22728 (N_22728,N_22328,N_22266);
or U22729 (N_22729,N_22366,N_22265);
nor U22730 (N_22730,N_22414,N_22482);
nor U22731 (N_22731,N_22349,N_22345);
or U22732 (N_22732,N_22317,N_22254);
xnor U22733 (N_22733,N_22434,N_22409);
nand U22734 (N_22734,N_22265,N_22289);
nand U22735 (N_22735,N_22346,N_22315);
nor U22736 (N_22736,N_22379,N_22469);
or U22737 (N_22737,N_22442,N_22319);
and U22738 (N_22738,N_22368,N_22475);
nor U22739 (N_22739,N_22251,N_22452);
and U22740 (N_22740,N_22282,N_22492);
nor U22741 (N_22741,N_22351,N_22475);
nor U22742 (N_22742,N_22436,N_22401);
xnor U22743 (N_22743,N_22468,N_22257);
nand U22744 (N_22744,N_22372,N_22497);
nor U22745 (N_22745,N_22418,N_22327);
nand U22746 (N_22746,N_22388,N_22339);
nor U22747 (N_22747,N_22330,N_22373);
and U22748 (N_22748,N_22441,N_22486);
xnor U22749 (N_22749,N_22354,N_22360);
nand U22750 (N_22750,N_22657,N_22747);
or U22751 (N_22751,N_22652,N_22689);
nand U22752 (N_22752,N_22733,N_22697);
nor U22753 (N_22753,N_22625,N_22643);
nand U22754 (N_22754,N_22541,N_22580);
nor U22755 (N_22755,N_22513,N_22512);
nor U22756 (N_22756,N_22590,N_22639);
nand U22757 (N_22757,N_22714,N_22609);
or U22758 (N_22758,N_22572,N_22504);
and U22759 (N_22759,N_22524,N_22745);
or U22760 (N_22760,N_22596,N_22662);
or U22761 (N_22761,N_22537,N_22718);
and U22762 (N_22762,N_22730,N_22505);
and U22763 (N_22763,N_22583,N_22653);
xnor U22764 (N_22764,N_22561,N_22707);
nor U22765 (N_22765,N_22660,N_22691);
or U22766 (N_22766,N_22615,N_22749);
or U22767 (N_22767,N_22716,N_22654);
and U22768 (N_22768,N_22503,N_22741);
nor U22769 (N_22769,N_22594,N_22558);
xnor U22770 (N_22770,N_22532,N_22634);
or U22771 (N_22771,N_22669,N_22578);
or U22772 (N_22772,N_22575,N_22713);
or U22773 (N_22773,N_22507,N_22678);
nor U22774 (N_22774,N_22563,N_22599);
nor U22775 (N_22775,N_22570,N_22728);
and U22776 (N_22776,N_22619,N_22616);
nand U22777 (N_22777,N_22637,N_22506);
nand U22778 (N_22778,N_22602,N_22564);
nor U22779 (N_22779,N_22527,N_22726);
and U22780 (N_22780,N_22631,N_22723);
nand U22781 (N_22781,N_22618,N_22635);
nor U22782 (N_22782,N_22722,N_22579);
and U22783 (N_22783,N_22548,N_22724);
xnor U22784 (N_22784,N_22549,N_22708);
nor U22785 (N_22785,N_22673,N_22606);
and U22786 (N_22786,N_22626,N_22569);
or U22787 (N_22787,N_22629,N_22687);
and U22788 (N_22788,N_22556,N_22638);
and U22789 (N_22789,N_22529,N_22547);
nor U22790 (N_22790,N_22738,N_22603);
or U22791 (N_22791,N_22735,N_22627);
nand U22792 (N_22792,N_22675,N_22628);
xnor U22793 (N_22793,N_22717,N_22676);
xnor U22794 (N_22794,N_22645,N_22582);
xor U22795 (N_22795,N_22699,N_22706);
nor U22796 (N_22796,N_22608,N_22511);
nor U22797 (N_22797,N_22665,N_22624);
or U22798 (N_22798,N_22592,N_22641);
nand U22799 (N_22799,N_22559,N_22555);
nor U22800 (N_22800,N_22604,N_22661);
and U22801 (N_22801,N_22539,N_22659);
nor U22802 (N_22802,N_22646,N_22690);
and U22803 (N_22803,N_22528,N_22593);
and U22804 (N_22804,N_22632,N_22721);
or U22805 (N_22805,N_22671,N_22742);
nor U22806 (N_22806,N_22636,N_22514);
and U22807 (N_22807,N_22702,N_22553);
or U22808 (N_22808,N_22701,N_22725);
xor U22809 (N_22809,N_22623,N_22536);
nand U22810 (N_22810,N_22720,N_22703);
nor U22811 (N_22811,N_22670,N_22746);
or U22812 (N_22812,N_22740,N_22612);
nand U22813 (N_22813,N_22577,N_22538);
or U22814 (N_22814,N_22666,N_22520);
nor U22815 (N_22815,N_22573,N_22607);
or U22816 (N_22816,N_22732,N_22620);
nor U22817 (N_22817,N_22617,N_22684);
xor U22818 (N_22818,N_22682,N_22587);
nand U22819 (N_22819,N_22557,N_22674);
nand U22820 (N_22820,N_22552,N_22719);
nor U22821 (N_22821,N_22656,N_22551);
and U22822 (N_22822,N_22748,N_22501);
or U22823 (N_22823,N_22651,N_22508);
xnor U22824 (N_22824,N_22543,N_22737);
nand U22825 (N_22825,N_22568,N_22509);
xor U22826 (N_22826,N_22709,N_22531);
xnor U22827 (N_22827,N_22712,N_22704);
nor U22828 (N_22828,N_22743,N_22633);
nand U22829 (N_22829,N_22586,N_22605);
nand U22830 (N_22830,N_22640,N_22694);
and U22831 (N_22831,N_22550,N_22515);
or U22832 (N_22832,N_22610,N_22685);
xor U22833 (N_22833,N_22650,N_22522);
nor U22834 (N_22834,N_22710,N_22664);
or U22835 (N_22835,N_22681,N_22734);
nor U22836 (N_22836,N_22560,N_22648);
or U22837 (N_22837,N_22526,N_22688);
xnor U22838 (N_22838,N_22518,N_22516);
nand U22839 (N_22839,N_22567,N_22545);
nor U22840 (N_22840,N_22686,N_22683);
or U22841 (N_22841,N_22614,N_22601);
xor U22842 (N_22842,N_22736,N_22581);
nand U22843 (N_22843,N_22525,N_22621);
xnor U22844 (N_22844,N_22544,N_22655);
nand U22845 (N_22845,N_22546,N_22693);
nand U22846 (N_22846,N_22554,N_22680);
or U22847 (N_22847,N_22521,N_22565);
or U22848 (N_22848,N_22695,N_22588);
xor U22849 (N_22849,N_22647,N_22562);
xnor U22850 (N_22850,N_22744,N_22540);
or U22851 (N_22851,N_22672,N_22510);
nor U22852 (N_22852,N_22658,N_22591);
nand U22853 (N_22853,N_22502,N_22649);
and U22854 (N_22854,N_22585,N_22715);
and U22855 (N_22855,N_22642,N_22668);
or U22856 (N_22856,N_22571,N_22534);
nand U22857 (N_22857,N_22667,N_22519);
and U22858 (N_22858,N_22576,N_22622);
and U22859 (N_22859,N_22533,N_22523);
or U22860 (N_22860,N_22698,N_22679);
and U22861 (N_22861,N_22727,N_22705);
and U22862 (N_22862,N_22500,N_22597);
or U22863 (N_22863,N_22542,N_22692);
xor U22864 (N_22864,N_22644,N_22739);
nor U22865 (N_22865,N_22595,N_22696);
nor U22866 (N_22866,N_22535,N_22517);
nand U22867 (N_22867,N_22711,N_22731);
nand U22868 (N_22868,N_22700,N_22589);
xnor U22869 (N_22869,N_22574,N_22663);
nand U22870 (N_22870,N_22729,N_22530);
nand U22871 (N_22871,N_22598,N_22584);
nand U22872 (N_22872,N_22611,N_22566);
and U22873 (N_22873,N_22677,N_22630);
nand U22874 (N_22874,N_22600,N_22613);
xor U22875 (N_22875,N_22649,N_22744);
nor U22876 (N_22876,N_22730,N_22609);
nor U22877 (N_22877,N_22527,N_22575);
or U22878 (N_22878,N_22523,N_22728);
xnor U22879 (N_22879,N_22680,N_22694);
nand U22880 (N_22880,N_22659,N_22607);
xor U22881 (N_22881,N_22626,N_22689);
or U22882 (N_22882,N_22736,N_22626);
or U22883 (N_22883,N_22643,N_22507);
nand U22884 (N_22884,N_22664,N_22639);
nor U22885 (N_22885,N_22707,N_22722);
or U22886 (N_22886,N_22546,N_22663);
nand U22887 (N_22887,N_22596,N_22503);
nor U22888 (N_22888,N_22543,N_22703);
and U22889 (N_22889,N_22743,N_22685);
nand U22890 (N_22890,N_22725,N_22569);
nand U22891 (N_22891,N_22729,N_22705);
xnor U22892 (N_22892,N_22662,N_22723);
nand U22893 (N_22893,N_22687,N_22737);
nand U22894 (N_22894,N_22640,N_22643);
or U22895 (N_22895,N_22612,N_22540);
and U22896 (N_22896,N_22524,N_22579);
xnor U22897 (N_22897,N_22509,N_22538);
nor U22898 (N_22898,N_22614,N_22646);
nand U22899 (N_22899,N_22523,N_22575);
and U22900 (N_22900,N_22699,N_22516);
nor U22901 (N_22901,N_22670,N_22615);
nand U22902 (N_22902,N_22531,N_22717);
or U22903 (N_22903,N_22685,N_22519);
xnor U22904 (N_22904,N_22531,N_22540);
nand U22905 (N_22905,N_22735,N_22531);
nor U22906 (N_22906,N_22630,N_22653);
nor U22907 (N_22907,N_22570,N_22735);
or U22908 (N_22908,N_22565,N_22513);
nor U22909 (N_22909,N_22693,N_22615);
or U22910 (N_22910,N_22558,N_22541);
and U22911 (N_22911,N_22568,N_22651);
nor U22912 (N_22912,N_22729,N_22698);
or U22913 (N_22913,N_22596,N_22682);
and U22914 (N_22914,N_22666,N_22522);
nor U22915 (N_22915,N_22614,N_22597);
nand U22916 (N_22916,N_22500,N_22691);
and U22917 (N_22917,N_22505,N_22561);
and U22918 (N_22918,N_22610,N_22618);
xor U22919 (N_22919,N_22563,N_22573);
or U22920 (N_22920,N_22504,N_22554);
or U22921 (N_22921,N_22690,N_22737);
xnor U22922 (N_22922,N_22518,N_22687);
nand U22923 (N_22923,N_22670,N_22629);
or U22924 (N_22924,N_22511,N_22583);
or U22925 (N_22925,N_22686,N_22645);
or U22926 (N_22926,N_22510,N_22612);
nand U22927 (N_22927,N_22744,N_22742);
nand U22928 (N_22928,N_22703,N_22592);
nand U22929 (N_22929,N_22650,N_22557);
or U22930 (N_22930,N_22697,N_22522);
and U22931 (N_22931,N_22726,N_22560);
nor U22932 (N_22932,N_22542,N_22543);
nor U22933 (N_22933,N_22527,N_22664);
and U22934 (N_22934,N_22656,N_22561);
nor U22935 (N_22935,N_22558,N_22725);
or U22936 (N_22936,N_22622,N_22665);
or U22937 (N_22937,N_22613,N_22586);
xnor U22938 (N_22938,N_22527,N_22641);
and U22939 (N_22939,N_22540,N_22524);
xnor U22940 (N_22940,N_22558,N_22703);
or U22941 (N_22941,N_22549,N_22647);
or U22942 (N_22942,N_22562,N_22681);
nand U22943 (N_22943,N_22525,N_22660);
xor U22944 (N_22944,N_22628,N_22533);
xnor U22945 (N_22945,N_22591,N_22549);
nor U22946 (N_22946,N_22620,N_22626);
xnor U22947 (N_22947,N_22572,N_22644);
and U22948 (N_22948,N_22709,N_22581);
xor U22949 (N_22949,N_22628,N_22738);
nor U22950 (N_22950,N_22541,N_22505);
or U22951 (N_22951,N_22549,N_22667);
nand U22952 (N_22952,N_22723,N_22524);
and U22953 (N_22953,N_22586,N_22501);
and U22954 (N_22954,N_22639,N_22573);
nand U22955 (N_22955,N_22572,N_22554);
nor U22956 (N_22956,N_22595,N_22712);
xnor U22957 (N_22957,N_22633,N_22732);
or U22958 (N_22958,N_22500,N_22506);
or U22959 (N_22959,N_22560,N_22505);
or U22960 (N_22960,N_22501,N_22729);
nand U22961 (N_22961,N_22661,N_22648);
or U22962 (N_22962,N_22700,N_22618);
or U22963 (N_22963,N_22671,N_22622);
nand U22964 (N_22964,N_22525,N_22640);
or U22965 (N_22965,N_22744,N_22580);
or U22966 (N_22966,N_22587,N_22716);
or U22967 (N_22967,N_22514,N_22516);
or U22968 (N_22968,N_22624,N_22563);
and U22969 (N_22969,N_22586,N_22654);
nand U22970 (N_22970,N_22532,N_22690);
xor U22971 (N_22971,N_22671,N_22737);
or U22972 (N_22972,N_22649,N_22543);
or U22973 (N_22973,N_22524,N_22638);
and U22974 (N_22974,N_22585,N_22744);
or U22975 (N_22975,N_22536,N_22649);
nand U22976 (N_22976,N_22540,N_22599);
and U22977 (N_22977,N_22702,N_22716);
xnor U22978 (N_22978,N_22627,N_22684);
and U22979 (N_22979,N_22716,N_22527);
nand U22980 (N_22980,N_22638,N_22722);
and U22981 (N_22981,N_22696,N_22673);
nor U22982 (N_22982,N_22500,N_22509);
nand U22983 (N_22983,N_22530,N_22715);
and U22984 (N_22984,N_22594,N_22662);
and U22985 (N_22985,N_22745,N_22526);
nand U22986 (N_22986,N_22633,N_22648);
and U22987 (N_22987,N_22565,N_22652);
nor U22988 (N_22988,N_22747,N_22543);
xor U22989 (N_22989,N_22703,N_22674);
or U22990 (N_22990,N_22548,N_22521);
nor U22991 (N_22991,N_22593,N_22537);
and U22992 (N_22992,N_22649,N_22581);
and U22993 (N_22993,N_22573,N_22637);
xnor U22994 (N_22994,N_22615,N_22518);
nand U22995 (N_22995,N_22574,N_22595);
and U22996 (N_22996,N_22645,N_22733);
and U22997 (N_22997,N_22720,N_22592);
nand U22998 (N_22998,N_22704,N_22500);
or U22999 (N_22999,N_22680,N_22608);
and U23000 (N_23000,N_22915,N_22952);
xnor U23001 (N_23001,N_22795,N_22808);
xnor U23002 (N_23002,N_22826,N_22939);
and U23003 (N_23003,N_22773,N_22931);
and U23004 (N_23004,N_22870,N_22832);
nor U23005 (N_23005,N_22886,N_22871);
xnor U23006 (N_23006,N_22760,N_22917);
nor U23007 (N_23007,N_22891,N_22847);
xnor U23008 (N_23008,N_22788,N_22932);
or U23009 (N_23009,N_22767,N_22950);
and U23010 (N_23010,N_22850,N_22991);
nor U23011 (N_23011,N_22887,N_22805);
nand U23012 (N_23012,N_22980,N_22763);
or U23013 (N_23013,N_22992,N_22879);
nor U23014 (N_23014,N_22813,N_22923);
xnor U23015 (N_23015,N_22962,N_22946);
nand U23016 (N_23016,N_22971,N_22831);
or U23017 (N_23017,N_22890,N_22762);
nor U23018 (N_23018,N_22970,N_22920);
xor U23019 (N_23019,N_22827,N_22967);
nor U23020 (N_23020,N_22810,N_22951);
or U23021 (N_23021,N_22872,N_22841);
nand U23022 (N_23022,N_22776,N_22799);
xnor U23023 (N_23023,N_22884,N_22855);
and U23024 (N_23024,N_22780,N_22995);
and U23025 (N_23025,N_22926,N_22944);
and U23026 (N_23026,N_22755,N_22792);
or U23027 (N_23027,N_22924,N_22934);
or U23028 (N_23028,N_22817,N_22938);
or U23029 (N_23029,N_22921,N_22968);
and U23030 (N_23030,N_22818,N_22948);
xnor U23031 (N_23031,N_22791,N_22843);
xnor U23032 (N_23032,N_22957,N_22930);
xnor U23033 (N_23033,N_22947,N_22966);
xor U23034 (N_23034,N_22894,N_22833);
nor U23035 (N_23035,N_22774,N_22965);
xor U23036 (N_23036,N_22954,N_22861);
nor U23037 (N_23037,N_22949,N_22985);
nor U23038 (N_23038,N_22880,N_22840);
nor U23039 (N_23039,N_22860,N_22765);
and U23040 (N_23040,N_22943,N_22769);
or U23041 (N_23041,N_22918,N_22972);
nand U23042 (N_23042,N_22961,N_22825);
nand U23043 (N_23043,N_22858,N_22775);
xnor U23044 (N_23044,N_22936,N_22854);
nand U23045 (N_23045,N_22901,N_22974);
nor U23046 (N_23046,N_22777,N_22781);
xor U23047 (N_23047,N_22839,N_22803);
nor U23048 (N_23048,N_22888,N_22784);
nor U23049 (N_23049,N_22996,N_22830);
nand U23050 (N_23050,N_22778,N_22794);
nand U23051 (N_23051,N_22779,N_22916);
or U23052 (N_23052,N_22896,N_22989);
nor U23053 (N_23053,N_22909,N_22868);
or U23054 (N_23054,N_22874,N_22809);
or U23055 (N_23055,N_22821,N_22897);
or U23056 (N_23056,N_22983,N_22925);
nand U23057 (N_23057,N_22849,N_22940);
nand U23058 (N_23058,N_22990,N_22796);
nor U23059 (N_23059,N_22802,N_22856);
nand U23060 (N_23060,N_22790,N_22812);
xor U23061 (N_23061,N_22999,N_22927);
nand U23062 (N_23062,N_22878,N_22804);
nand U23063 (N_23063,N_22756,N_22875);
nand U23064 (N_23064,N_22751,N_22829);
xnor U23065 (N_23065,N_22753,N_22933);
or U23066 (N_23066,N_22899,N_22876);
and U23067 (N_23067,N_22913,N_22862);
and U23068 (N_23068,N_22864,N_22761);
or U23069 (N_23069,N_22787,N_22772);
nor U23070 (N_23070,N_22977,N_22998);
and U23071 (N_23071,N_22953,N_22837);
and U23072 (N_23072,N_22786,N_22906);
xnor U23073 (N_23073,N_22877,N_22922);
nand U23074 (N_23074,N_22902,N_22835);
xnor U23075 (N_23075,N_22789,N_22758);
xor U23076 (N_23076,N_22801,N_22942);
nor U23077 (N_23077,N_22973,N_22834);
nor U23078 (N_23078,N_22898,N_22811);
nor U23079 (N_23079,N_22853,N_22848);
and U23080 (N_23080,N_22929,N_22873);
and U23081 (N_23081,N_22820,N_22846);
or U23082 (N_23082,N_22987,N_22911);
nand U23083 (N_23083,N_22807,N_22838);
and U23084 (N_23084,N_22759,N_22928);
and U23085 (N_23085,N_22766,N_22867);
xor U23086 (N_23086,N_22941,N_22997);
nand U23087 (N_23087,N_22978,N_22851);
nor U23088 (N_23088,N_22979,N_22919);
nor U23089 (N_23089,N_22893,N_22785);
nor U23090 (N_23090,N_22800,N_22816);
and U23091 (N_23091,N_22844,N_22866);
xnor U23092 (N_23092,N_22845,N_22988);
nand U23093 (N_23093,N_22836,N_22863);
or U23094 (N_23094,N_22806,N_22828);
or U23095 (N_23095,N_22892,N_22793);
or U23096 (N_23096,N_22994,N_22963);
xor U23097 (N_23097,N_22814,N_22815);
nand U23098 (N_23098,N_22959,N_22937);
nand U23099 (N_23099,N_22955,N_22859);
or U23100 (N_23100,N_22907,N_22895);
xnor U23101 (N_23101,N_22905,N_22976);
nor U23102 (N_23102,N_22768,N_22914);
xor U23103 (N_23103,N_22783,N_22900);
nor U23104 (N_23104,N_22869,N_22982);
nand U23105 (N_23105,N_22935,N_22945);
and U23106 (N_23106,N_22822,N_22986);
nand U23107 (N_23107,N_22764,N_22797);
nor U23108 (N_23108,N_22883,N_22984);
nand U23109 (N_23109,N_22752,N_22958);
and U23110 (N_23110,N_22969,N_22750);
nor U23111 (N_23111,N_22885,N_22754);
or U23112 (N_23112,N_22842,N_22889);
nand U23113 (N_23113,N_22912,N_22824);
xnor U23114 (N_23114,N_22975,N_22882);
or U23115 (N_23115,N_22865,N_22903);
or U23116 (N_23116,N_22910,N_22993);
or U23117 (N_23117,N_22819,N_22881);
or U23118 (N_23118,N_22904,N_22981);
or U23119 (N_23119,N_22857,N_22782);
nor U23120 (N_23120,N_22798,N_22823);
or U23121 (N_23121,N_22852,N_22757);
nand U23122 (N_23122,N_22960,N_22964);
or U23123 (N_23123,N_22771,N_22956);
nor U23124 (N_23124,N_22770,N_22908);
xnor U23125 (N_23125,N_22931,N_22781);
and U23126 (N_23126,N_22940,N_22958);
xnor U23127 (N_23127,N_22960,N_22847);
xor U23128 (N_23128,N_22778,N_22875);
or U23129 (N_23129,N_22993,N_22780);
nor U23130 (N_23130,N_22836,N_22961);
xnor U23131 (N_23131,N_22956,N_22975);
or U23132 (N_23132,N_22889,N_22969);
xor U23133 (N_23133,N_22929,N_22977);
and U23134 (N_23134,N_22840,N_22917);
nand U23135 (N_23135,N_22818,N_22956);
xnor U23136 (N_23136,N_22799,N_22885);
nor U23137 (N_23137,N_22967,N_22985);
or U23138 (N_23138,N_22784,N_22766);
nor U23139 (N_23139,N_22909,N_22889);
nand U23140 (N_23140,N_22932,N_22901);
and U23141 (N_23141,N_22830,N_22962);
nor U23142 (N_23142,N_22897,N_22980);
nor U23143 (N_23143,N_22949,N_22752);
nor U23144 (N_23144,N_22934,N_22761);
nor U23145 (N_23145,N_22839,N_22771);
xnor U23146 (N_23146,N_22927,N_22896);
or U23147 (N_23147,N_22760,N_22938);
or U23148 (N_23148,N_22920,N_22830);
and U23149 (N_23149,N_22992,N_22822);
and U23150 (N_23150,N_22768,N_22869);
nand U23151 (N_23151,N_22998,N_22814);
xor U23152 (N_23152,N_22780,N_22880);
or U23153 (N_23153,N_22906,N_22953);
nor U23154 (N_23154,N_22872,N_22947);
or U23155 (N_23155,N_22970,N_22895);
and U23156 (N_23156,N_22970,N_22922);
nor U23157 (N_23157,N_22816,N_22756);
nand U23158 (N_23158,N_22831,N_22854);
and U23159 (N_23159,N_22821,N_22781);
xnor U23160 (N_23160,N_22824,N_22935);
nand U23161 (N_23161,N_22831,N_22816);
xnor U23162 (N_23162,N_22781,N_22921);
xor U23163 (N_23163,N_22851,N_22761);
and U23164 (N_23164,N_22813,N_22920);
nor U23165 (N_23165,N_22944,N_22827);
or U23166 (N_23166,N_22952,N_22837);
nor U23167 (N_23167,N_22759,N_22774);
or U23168 (N_23168,N_22997,N_22965);
or U23169 (N_23169,N_22753,N_22983);
and U23170 (N_23170,N_22978,N_22920);
nor U23171 (N_23171,N_22942,N_22832);
or U23172 (N_23172,N_22787,N_22884);
xor U23173 (N_23173,N_22973,N_22774);
or U23174 (N_23174,N_22771,N_22762);
and U23175 (N_23175,N_22802,N_22930);
xnor U23176 (N_23176,N_22868,N_22887);
or U23177 (N_23177,N_22918,N_22964);
and U23178 (N_23178,N_22826,N_22866);
nand U23179 (N_23179,N_22805,N_22976);
or U23180 (N_23180,N_22858,N_22878);
nor U23181 (N_23181,N_22765,N_22750);
nor U23182 (N_23182,N_22835,N_22782);
or U23183 (N_23183,N_22762,N_22984);
or U23184 (N_23184,N_22885,N_22761);
xnor U23185 (N_23185,N_22836,N_22822);
and U23186 (N_23186,N_22847,N_22844);
or U23187 (N_23187,N_22756,N_22846);
or U23188 (N_23188,N_22962,N_22764);
nand U23189 (N_23189,N_22852,N_22823);
or U23190 (N_23190,N_22768,N_22973);
or U23191 (N_23191,N_22866,N_22815);
or U23192 (N_23192,N_22806,N_22750);
or U23193 (N_23193,N_22755,N_22878);
and U23194 (N_23194,N_22776,N_22949);
or U23195 (N_23195,N_22817,N_22932);
or U23196 (N_23196,N_22952,N_22765);
and U23197 (N_23197,N_22921,N_22758);
nor U23198 (N_23198,N_22845,N_22815);
nor U23199 (N_23199,N_22998,N_22871);
nand U23200 (N_23200,N_22811,N_22885);
or U23201 (N_23201,N_22988,N_22933);
or U23202 (N_23202,N_22962,N_22819);
or U23203 (N_23203,N_22930,N_22806);
and U23204 (N_23204,N_22988,N_22782);
xnor U23205 (N_23205,N_22873,N_22835);
or U23206 (N_23206,N_22962,N_22767);
xor U23207 (N_23207,N_22810,N_22891);
xnor U23208 (N_23208,N_22950,N_22790);
or U23209 (N_23209,N_22752,N_22959);
xor U23210 (N_23210,N_22971,N_22927);
xnor U23211 (N_23211,N_22847,N_22985);
and U23212 (N_23212,N_22781,N_22895);
and U23213 (N_23213,N_22877,N_22869);
and U23214 (N_23214,N_22759,N_22857);
and U23215 (N_23215,N_22768,N_22812);
nor U23216 (N_23216,N_22902,N_22890);
nand U23217 (N_23217,N_22949,N_22777);
nand U23218 (N_23218,N_22984,N_22957);
nand U23219 (N_23219,N_22967,N_22932);
xnor U23220 (N_23220,N_22908,N_22854);
or U23221 (N_23221,N_22842,N_22776);
nand U23222 (N_23222,N_22819,N_22998);
nor U23223 (N_23223,N_22885,N_22919);
nor U23224 (N_23224,N_22858,N_22993);
or U23225 (N_23225,N_22879,N_22761);
nor U23226 (N_23226,N_22996,N_22808);
or U23227 (N_23227,N_22784,N_22894);
nand U23228 (N_23228,N_22909,N_22765);
or U23229 (N_23229,N_22909,N_22824);
nand U23230 (N_23230,N_22991,N_22842);
and U23231 (N_23231,N_22984,N_22889);
and U23232 (N_23232,N_22811,N_22810);
nand U23233 (N_23233,N_22880,N_22864);
nand U23234 (N_23234,N_22758,N_22876);
nand U23235 (N_23235,N_22798,N_22861);
xor U23236 (N_23236,N_22936,N_22776);
nor U23237 (N_23237,N_22863,N_22933);
nand U23238 (N_23238,N_22878,N_22883);
and U23239 (N_23239,N_22875,N_22813);
xor U23240 (N_23240,N_22807,N_22902);
and U23241 (N_23241,N_22922,N_22779);
nand U23242 (N_23242,N_22957,N_22805);
nor U23243 (N_23243,N_22976,N_22875);
xnor U23244 (N_23244,N_22972,N_22815);
xor U23245 (N_23245,N_22909,N_22785);
nor U23246 (N_23246,N_22842,N_22879);
nand U23247 (N_23247,N_22801,N_22777);
xnor U23248 (N_23248,N_22995,N_22809);
xor U23249 (N_23249,N_22861,N_22887);
nand U23250 (N_23250,N_23003,N_23052);
nor U23251 (N_23251,N_23097,N_23195);
xor U23252 (N_23252,N_23226,N_23146);
and U23253 (N_23253,N_23228,N_23090);
and U23254 (N_23254,N_23044,N_23137);
xnor U23255 (N_23255,N_23075,N_23011);
or U23256 (N_23256,N_23229,N_23192);
or U23257 (N_23257,N_23008,N_23110);
and U23258 (N_23258,N_23194,N_23236);
or U23259 (N_23259,N_23221,N_23161);
nand U23260 (N_23260,N_23019,N_23061);
or U23261 (N_23261,N_23000,N_23207);
nor U23262 (N_23262,N_23069,N_23186);
nand U23263 (N_23263,N_23035,N_23010);
and U23264 (N_23264,N_23086,N_23201);
and U23265 (N_23265,N_23203,N_23038);
or U23266 (N_23266,N_23031,N_23135);
nor U23267 (N_23267,N_23223,N_23157);
or U23268 (N_23268,N_23120,N_23138);
nand U23269 (N_23269,N_23119,N_23050);
and U23270 (N_23270,N_23096,N_23141);
nand U23271 (N_23271,N_23217,N_23187);
and U23272 (N_23272,N_23022,N_23104);
and U23273 (N_23273,N_23098,N_23128);
xor U23274 (N_23274,N_23206,N_23015);
or U23275 (N_23275,N_23046,N_23042);
nor U23276 (N_23276,N_23143,N_23188);
nand U23277 (N_23277,N_23125,N_23145);
nor U23278 (N_23278,N_23099,N_23153);
and U23279 (N_23279,N_23248,N_23094);
nor U23280 (N_23280,N_23012,N_23179);
and U23281 (N_23281,N_23001,N_23040);
xor U23282 (N_23282,N_23177,N_23017);
and U23283 (N_23283,N_23156,N_23232);
nand U23284 (N_23284,N_23147,N_23202);
or U23285 (N_23285,N_23112,N_23048);
xnor U23286 (N_23286,N_23133,N_23211);
xnor U23287 (N_23287,N_23111,N_23065);
xor U23288 (N_23288,N_23160,N_23037);
nor U23289 (N_23289,N_23173,N_23164);
nor U23290 (N_23290,N_23126,N_23130);
xnor U23291 (N_23291,N_23100,N_23136);
nor U23292 (N_23292,N_23200,N_23049);
xnor U23293 (N_23293,N_23047,N_23242);
or U23294 (N_23294,N_23152,N_23208);
and U23295 (N_23295,N_23107,N_23004);
nor U23296 (N_23296,N_23005,N_23106);
nor U23297 (N_23297,N_23243,N_23244);
xor U23298 (N_23298,N_23002,N_23155);
or U23299 (N_23299,N_23091,N_23029);
xor U23300 (N_23300,N_23085,N_23093);
xnor U23301 (N_23301,N_23116,N_23034);
and U23302 (N_23302,N_23180,N_23131);
nor U23303 (N_23303,N_23123,N_23174);
nor U23304 (N_23304,N_23247,N_23073);
or U23305 (N_23305,N_23246,N_23058);
or U23306 (N_23306,N_23193,N_23101);
nor U23307 (N_23307,N_23081,N_23064);
nand U23308 (N_23308,N_23235,N_23088);
xnor U23309 (N_23309,N_23055,N_23082);
or U23310 (N_23310,N_23190,N_23020);
nand U23311 (N_23311,N_23166,N_23139);
xor U23312 (N_23312,N_23227,N_23181);
and U23313 (N_23313,N_23033,N_23039);
nand U23314 (N_23314,N_23027,N_23014);
or U23315 (N_23315,N_23071,N_23144);
xnor U23316 (N_23316,N_23108,N_23197);
or U23317 (N_23317,N_23218,N_23238);
xor U23318 (N_23318,N_23067,N_23025);
xor U23319 (N_23319,N_23198,N_23230);
or U23320 (N_23320,N_23016,N_23079);
xor U23321 (N_23321,N_23148,N_23239);
nor U23322 (N_23322,N_23054,N_23165);
or U23323 (N_23323,N_23007,N_23095);
and U23324 (N_23324,N_23185,N_23234);
nand U23325 (N_23325,N_23041,N_23026);
nor U23326 (N_23326,N_23162,N_23122);
nand U23327 (N_23327,N_23220,N_23013);
nand U23328 (N_23328,N_23068,N_23129);
xnor U23329 (N_23329,N_23140,N_23056);
xor U23330 (N_23330,N_23171,N_23105);
and U23331 (N_23331,N_23237,N_23184);
or U23332 (N_23332,N_23231,N_23053);
nand U23333 (N_23333,N_23113,N_23212);
xor U23334 (N_23334,N_23225,N_23009);
nand U23335 (N_23335,N_23233,N_23083);
xnor U23336 (N_23336,N_23151,N_23024);
or U23337 (N_23337,N_23084,N_23109);
or U23338 (N_23338,N_23150,N_23163);
or U23339 (N_23339,N_23209,N_23018);
and U23340 (N_23340,N_23224,N_23149);
or U23341 (N_23341,N_23021,N_23032);
or U23342 (N_23342,N_23216,N_23219);
nand U23343 (N_23343,N_23240,N_23172);
xor U23344 (N_23344,N_23103,N_23063);
xor U23345 (N_23345,N_23030,N_23182);
nor U23346 (N_23346,N_23070,N_23045);
or U23347 (N_23347,N_23154,N_23170);
nor U23348 (N_23348,N_23196,N_23213);
xor U23349 (N_23349,N_23089,N_23215);
nand U23350 (N_23350,N_23072,N_23178);
xnor U23351 (N_23351,N_23167,N_23124);
and U23352 (N_23352,N_23051,N_23210);
or U23353 (N_23353,N_23074,N_23214);
nand U23354 (N_23354,N_23205,N_23183);
nor U23355 (N_23355,N_23092,N_23204);
xor U23356 (N_23356,N_23059,N_23132);
and U23357 (N_23357,N_23115,N_23169);
nor U23358 (N_23358,N_23057,N_23102);
nand U23359 (N_23359,N_23006,N_23158);
and U23360 (N_23360,N_23134,N_23077);
or U23361 (N_23361,N_23114,N_23176);
or U23362 (N_23362,N_23043,N_23028);
nand U23363 (N_23363,N_23121,N_23060);
and U23364 (N_23364,N_23159,N_23062);
nor U23365 (N_23365,N_23023,N_23222);
xnor U23366 (N_23366,N_23142,N_23118);
xnor U23367 (N_23367,N_23078,N_23249);
nand U23368 (N_23368,N_23076,N_23036);
or U23369 (N_23369,N_23199,N_23087);
or U23370 (N_23370,N_23117,N_23191);
and U23371 (N_23371,N_23080,N_23245);
nand U23372 (N_23372,N_23168,N_23066);
nor U23373 (N_23373,N_23241,N_23127);
nand U23374 (N_23374,N_23189,N_23175);
nor U23375 (N_23375,N_23063,N_23178);
nand U23376 (N_23376,N_23207,N_23220);
and U23377 (N_23377,N_23045,N_23241);
xor U23378 (N_23378,N_23108,N_23047);
or U23379 (N_23379,N_23035,N_23102);
and U23380 (N_23380,N_23120,N_23104);
or U23381 (N_23381,N_23164,N_23036);
or U23382 (N_23382,N_23222,N_23129);
nor U23383 (N_23383,N_23096,N_23234);
nor U23384 (N_23384,N_23182,N_23157);
nor U23385 (N_23385,N_23201,N_23178);
nor U23386 (N_23386,N_23095,N_23149);
and U23387 (N_23387,N_23136,N_23150);
nor U23388 (N_23388,N_23042,N_23075);
nand U23389 (N_23389,N_23221,N_23078);
xor U23390 (N_23390,N_23225,N_23149);
xnor U23391 (N_23391,N_23061,N_23198);
and U23392 (N_23392,N_23175,N_23114);
and U23393 (N_23393,N_23104,N_23149);
nand U23394 (N_23394,N_23070,N_23193);
xor U23395 (N_23395,N_23007,N_23004);
nor U23396 (N_23396,N_23067,N_23057);
xor U23397 (N_23397,N_23017,N_23167);
nor U23398 (N_23398,N_23072,N_23059);
nand U23399 (N_23399,N_23184,N_23177);
nor U23400 (N_23400,N_23095,N_23111);
and U23401 (N_23401,N_23124,N_23047);
and U23402 (N_23402,N_23214,N_23035);
or U23403 (N_23403,N_23075,N_23023);
nand U23404 (N_23404,N_23149,N_23106);
or U23405 (N_23405,N_23171,N_23131);
nor U23406 (N_23406,N_23016,N_23145);
and U23407 (N_23407,N_23023,N_23063);
xnor U23408 (N_23408,N_23036,N_23050);
xor U23409 (N_23409,N_23147,N_23120);
nand U23410 (N_23410,N_23219,N_23017);
or U23411 (N_23411,N_23047,N_23153);
xnor U23412 (N_23412,N_23217,N_23113);
nor U23413 (N_23413,N_23154,N_23113);
and U23414 (N_23414,N_23007,N_23181);
nor U23415 (N_23415,N_23178,N_23227);
and U23416 (N_23416,N_23222,N_23175);
and U23417 (N_23417,N_23126,N_23230);
and U23418 (N_23418,N_23038,N_23041);
xor U23419 (N_23419,N_23225,N_23037);
nand U23420 (N_23420,N_23109,N_23194);
xnor U23421 (N_23421,N_23099,N_23199);
nand U23422 (N_23422,N_23172,N_23023);
nor U23423 (N_23423,N_23023,N_23168);
nor U23424 (N_23424,N_23168,N_23045);
and U23425 (N_23425,N_23041,N_23115);
xnor U23426 (N_23426,N_23109,N_23006);
nor U23427 (N_23427,N_23203,N_23243);
xnor U23428 (N_23428,N_23238,N_23215);
xor U23429 (N_23429,N_23080,N_23061);
nor U23430 (N_23430,N_23228,N_23117);
or U23431 (N_23431,N_23039,N_23096);
and U23432 (N_23432,N_23238,N_23235);
nand U23433 (N_23433,N_23046,N_23066);
nand U23434 (N_23434,N_23048,N_23178);
and U23435 (N_23435,N_23000,N_23008);
and U23436 (N_23436,N_23216,N_23103);
or U23437 (N_23437,N_23200,N_23167);
and U23438 (N_23438,N_23009,N_23083);
nor U23439 (N_23439,N_23044,N_23182);
nor U23440 (N_23440,N_23006,N_23140);
or U23441 (N_23441,N_23190,N_23195);
nor U23442 (N_23442,N_23177,N_23092);
or U23443 (N_23443,N_23028,N_23215);
or U23444 (N_23444,N_23126,N_23128);
xnor U23445 (N_23445,N_23122,N_23000);
nor U23446 (N_23446,N_23002,N_23089);
nand U23447 (N_23447,N_23021,N_23087);
xnor U23448 (N_23448,N_23145,N_23206);
or U23449 (N_23449,N_23174,N_23206);
nand U23450 (N_23450,N_23117,N_23070);
or U23451 (N_23451,N_23235,N_23111);
xor U23452 (N_23452,N_23179,N_23010);
xnor U23453 (N_23453,N_23207,N_23010);
nand U23454 (N_23454,N_23095,N_23242);
xor U23455 (N_23455,N_23199,N_23114);
or U23456 (N_23456,N_23218,N_23249);
xor U23457 (N_23457,N_23168,N_23221);
or U23458 (N_23458,N_23048,N_23062);
or U23459 (N_23459,N_23185,N_23208);
or U23460 (N_23460,N_23151,N_23119);
and U23461 (N_23461,N_23079,N_23221);
or U23462 (N_23462,N_23173,N_23155);
nand U23463 (N_23463,N_23089,N_23061);
and U23464 (N_23464,N_23015,N_23081);
and U23465 (N_23465,N_23161,N_23110);
or U23466 (N_23466,N_23170,N_23196);
nor U23467 (N_23467,N_23154,N_23108);
and U23468 (N_23468,N_23105,N_23116);
or U23469 (N_23469,N_23079,N_23119);
nor U23470 (N_23470,N_23010,N_23204);
nand U23471 (N_23471,N_23051,N_23216);
or U23472 (N_23472,N_23231,N_23164);
nor U23473 (N_23473,N_23232,N_23238);
or U23474 (N_23474,N_23176,N_23036);
nand U23475 (N_23475,N_23249,N_23017);
and U23476 (N_23476,N_23015,N_23207);
xnor U23477 (N_23477,N_23122,N_23221);
and U23478 (N_23478,N_23086,N_23227);
nand U23479 (N_23479,N_23138,N_23217);
nand U23480 (N_23480,N_23161,N_23214);
xor U23481 (N_23481,N_23053,N_23221);
or U23482 (N_23482,N_23032,N_23072);
nand U23483 (N_23483,N_23011,N_23154);
or U23484 (N_23484,N_23135,N_23245);
or U23485 (N_23485,N_23111,N_23155);
nand U23486 (N_23486,N_23078,N_23145);
and U23487 (N_23487,N_23246,N_23182);
xor U23488 (N_23488,N_23016,N_23163);
nand U23489 (N_23489,N_23186,N_23112);
or U23490 (N_23490,N_23199,N_23195);
nand U23491 (N_23491,N_23010,N_23090);
and U23492 (N_23492,N_23019,N_23180);
or U23493 (N_23493,N_23159,N_23232);
nor U23494 (N_23494,N_23216,N_23111);
nand U23495 (N_23495,N_23209,N_23004);
and U23496 (N_23496,N_23166,N_23101);
or U23497 (N_23497,N_23239,N_23091);
nand U23498 (N_23498,N_23064,N_23068);
xnor U23499 (N_23499,N_23070,N_23224);
xor U23500 (N_23500,N_23477,N_23280);
or U23501 (N_23501,N_23398,N_23297);
nor U23502 (N_23502,N_23293,N_23429);
or U23503 (N_23503,N_23495,N_23288);
and U23504 (N_23504,N_23370,N_23255);
nand U23505 (N_23505,N_23354,N_23257);
nand U23506 (N_23506,N_23302,N_23410);
or U23507 (N_23507,N_23324,N_23285);
nand U23508 (N_23508,N_23436,N_23405);
nand U23509 (N_23509,N_23435,N_23490);
and U23510 (N_23510,N_23449,N_23369);
xnor U23511 (N_23511,N_23376,N_23278);
and U23512 (N_23512,N_23282,N_23378);
nor U23513 (N_23513,N_23296,N_23326);
nand U23514 (N_23514,N_23385,N_23301);
xor U23515 (N_23515,N_23344,N_23273);
nor U23516 (N_23516,N_23319,N_23414);
or U23517 (N_23517,N_23315,N_23345);
nand U23518 (N_23518,N_23412,N_23377);
nor U23519 (N_23519,N_23409,N_23483);
or U23520 (N_23520,N_23390,N_23379);
nand U23521 (N_23521,N_23389,N_23443);
nor U23522 (N_23522,N_23349,N_23305);
xor U23523 (N_23523,N_23439,N_23467);
or U23524 (N_23524,N_23375,N_23416);
xnor U23525 (N_23525,N_23430,N_23364);
xnor U23526 (N_23526,N_23265,N_23358);
nor U23527 (N_23527,N_23459,N_23386);
or U23528 (N_23528,N_23441,N_23460);
xnor U23529 (N_23529,N_23454,N_23362);
nor U23530 (N_23530,N_23457,N_23406);
or U23531 (N_23531,N_23417,N_23252);
and U23532 (N_23532,N_23472,N_23339);
nand U23533 (N_23533,N_23408,N_23317);
or U23534 (N_23534,N_23404,N_23481);
xor U23535 (N_23535,N_23261,N_23337);
nand U23536 (N_23536,N_23411,N_23399);
xnor U23537 (N_23537,N_23450,N_23298);
and U23538 (N_23538,N_23340,N_23311);
and U23539 (N_23539,N_23401,N_23456);
nor U23540 (N_23540,N_23251,N_23347);
or U23541 (N_23541,N_23445,N_23437);
xnor U23542 (N_23542,N_23356,N_23478);
nor U23543 (N_23543,N_23383,N_23394);
nand U23544 (N_23544,N_23299,N_23473);
and U23545 (N_23545,N_23476,N_23290);
or U23546 (N_23546,N_23359,N_23446);
nor U23547 (N_23547,N_23455,N_23479);
nand U23548 (N_23548,N_23309,N_23426);
nand U23549 (N_23549,N_23253,N_23323);
or U23550 (N_23550,N_23421,N_23488);
and U23551 (N_23551,N_23492,N_23361);
nand U23552 (N_23552,N_23307,N_23402);
or U23553 (N_23553,N_23447,N_23461);
and U23554 (N_23554,N_23300,N_23366);
xnor U23555 (N_23555,N_23275,N_23338);
nor U23556 (N_23556,N_23440,N_23420);
nor U23557 (N_23557,N_23276,N_23465);
or U23558 (N_23558,N_23335,N_23462);
nand U23559 (N_23559,N_23332,N_23487);
xor U23560 (N_23560,N_23343,N_23453);
or U23561 (N_23561,N_23346,N_23499);
or U23562 (N_23562,N_23427,N_23392);
nand U23563 (N_23563,N_23391,N_23452);
and U23564 (N_23564,N_23413,N_23432);
xor U23565 (N_23565,N_23480,N_23388);
xor U23566 (N_23566,N_23496,N_23303);
xor U23567 (N_23567,N_23365,N_23341);
and U23568 (N_23568,N_23397,N_23268);
nor U23569 (N_23569,N_23433,N_23415);
nand U23570 (N_23570,N_23372,N_23403);
nand U23571 (N_23571,N_23491,N_23292);
or U23572 (N_23572,N_23277,N_23428);
nor U23573 (N_23573,N_23310,N_23470);
nor U23574 (N_23574,N_23281,N_23313);
or U23575 (N_23575,N_23424,N_23423);
xor U23576 (N_23576,N_23497,N_23466);
or U23577 (N_23577,N_23387,N_23484);
nand U23578 (N_23578,N_23295,N_23474);
and U23579 (N_23579,N_23327,N_23486);
nor U23580 (N_23580,N_23380,N_23384);
xnor U23581 (N_23581,N_23352,N_23498);
nor U23582 (N_23582,N_23316,N_23489);
nand U23583 (N_23583,N_23314,N_23422);
xor U23584 (N_23584,N_23270,N_23494);
and U23585 (N_23585,N_23328,N_23431);
and U23586 (N_23586,N_23312,N_23438);
or U23587 (N_23587,N_23286,N_23350);
nor U23588 (N_23588,N_23262,N_23321);
and U23589 (N_23589,N_23272,N_23329);
nor U23590 (N_23590,N_23419,N_23373);
and U23591 (N_23591,N_23266,N_23400);
and U23592 (N_23592,N_23331,N_23464);
nand U23593 (N_23593,N_23260,N_23434);
and U23594 (N_23594,N_23374,N_23291);
xor U23595 (N_23595,N_23425,N_23367);
xor U23596 (N_23596,N_23318,N_23469);
nor U23597 (N_23597,N_23418,N_23284);
xor U23598 (N_23598,N_23287,N_23289);
or U23599 (N_23599,N_23250,N_23382);
nand U23600 (N_23600,N_23444,N_23368);
xor U23601 (N_23601,N_23334,N_23306);
nand U23602 (N_23602,N_23485,N_23283);
and U23603 (N_23603,N_23320,N_23355);
nand U23604 (N_23604,N_23294,N_23442);
xnor U23605 (N_23605,N_23395,N_23468);
nand U23606 (N_23606,N_23463,N_23493);
or U23607 (N_23607,N_23256,N_23325);
nand U23608 (N_23608,N_23348,N_23482);
xnor U23609 (N_23609,N_23304,N_23396);
xnor U23610 (N_23610,N_23360,N_23357);
or U23611 (N_23611,N_23342,N_23471);
or U23612 (N_23612,N_23259,N_23254);
nor U23613 (N_23613,N_23271,N_23322);
nand U23614 (N_23614,N_23407,N_23333);
or U23615 (N_23615,N_23475,N_23274);
nor U23616 (N_23616,N_23363,N_23308);
nand U23617 (N_23617,N_23351,N_23353);
xor U23618 (N_23618,N_23267,N_23458);
and U23619 (N_23619,N_23279,N_23393);
or U23620 (N_23620,N_23448,N_23269);
xor U23621 (N_23621,N_23336,N_23264);
nor U23622 (N_23622,N_23330,N_23381);
or U23623 (N_23623,N_23263,N_23451);
and U23624 (N_23624,N_23371,N_23258);
xnor U23625 (N_23625,N_23296,N_23392);
or U23626 (N_23626,N_23482,N_23365);
xnor U23627 (N_23627,N_23415,N_23295);
xor U23628 (N_23628,N_23482,N_23418);
and U23629 (N_23629,N_23392,N_23354);
nor U23630 (N_23630,N_23250,N_23271);
and U23631 (N_23631,N_23453,N_23281);
nand U23632 (N_23632,N_23455,N_23317);
nand U23633 (N_23633,N_23273,N_23271);
and U23634 (N_23634,N_23272,N_23311);
xnor U23635 (N_23635,N_23396,N_23405);
or U23636 (N_23636,N_23427,N_23432);
or U23637 (N_23637,N_23304,N_23309);
nor U23638 (N_23638,N_23369,N_23280);
nand U23639 (N_23639,N_23463,N_23383);
and U23640 (N_23640,N_23356,N_23456);
nor U23641 (N_23641,N_23333,N_23278);
or U23642 (N_23642,N_23315,N_23353);
nor U23643 (N_23643,N_23356,N_23435);
nand U23644 (N_23644,N_23377,N_23462);
or U23645 (N_23645,N_23381,N_23410);
xor U23646 (N_23646,N_23350,N_23344);
or U23647 (N_23647,N_23296,N_23387);
nand U23648 (N_23648,N_23354,N_23316);
nor U23649 (N_23649,N_23427,N_23363);
xnor U23650 (N_23650,N_23443,N_23405);
or U23651 (N_23651,N_23359,N_23323);
nand U23652 (N_23652,N_23444,N_23324);
nor U23653 (N_23653,N_23435,N_23434);
or U23654 (N_23654,N_23334,N_23321);
nor U23655 (N_23655,N_23264,N_23293);
xor U23656 (N_23656,N_23350,N_23366);
xnor U23657 (N_23657,N_23435,N_23424);
nor U23658 (N_23658,N_23256,N_23483);
nand U23659 (N_23659,N_23268,N_23464);
or U23660 (N_23660,N_23438,N_23464);
nor U23661 (N_23661,N_23369,N_23400);
or U23662 (N_23662,N_23459,N_23290);
nor U23663 (N_23663,N_23308,N_23361);
or U23664 (N_23664,N_23441,N_23254);
and U23665 (N_23665,N_23401,N_23300);
and U23666 (N_23666,N_23308,N_23323);
nand U23667 (N_23667,N_23455,N_23260);
xnor U23668 (N_23668,N_23322,N_23309);
xor U23669 (N_23669,N_23274,N_23467);
and U23670 (N_23670,N_23432,N_23479);
nor U23671 (N_23671,N_23333,N_23363);
or U23672 (N_23672,N_23412,N_23475);
xnor U23673 (N_23673,N_23302,N_23420);
and U23674 (N_23674,N_23364,N_23380);
nor U23675 (N_23675,N_23261,N_23406);
nand U23676 (N_23676,N_23337,N_23359);
nand U23677 (N_23677,N_23483,N_23378);
or U23678 (N_23678,N_23270,N_23484);
xor U23679 (N_23679,N_23393,N_23400);
and U23680 (N_23680,N_23272,N_23381);
xor U23681 (N_23681,N_23284,N_23374);
or U23682 (N_23682,N_23413,N_23404);
and U23683 (N_23683,N_23265,N_23469);
nor U23684 (N_23684,N_23438,N_23413);
nor U23685 (N_23685,N_23465,N_23342);
nand U23686 (N_23686,N_23367,N_23487);
nand U23687 (N_23687,N_23331,N_23394);
nand U23688 (N_23688,N_23454,N_23343);
xnor U23689 (N_23689,N_23326,N_23308);
xnor U23690 (N_23690,N_23471,N_23481);
and U23691 (N_23691,N_23466,N_23387);
nand U23692 (N_23692,N_23388,N_23467);
nand U23693 (N_23693,N_23359,N_23466);
or U23694 (N_23694,N_23390,N_23450);
nor U23695 (N_23695,N_23480,N_23390);
or U23696 (N_23696,N_23353,N_23336);
and U23697 (N_23697,N_23376,N_23439);
or U23698 (N_23698,N_23404,N_23290);
or U23699 (N_23699,N_23486,N_23299);
nor U23700 (N_23700,N_23343,N_23251);
xnor U23701 (N_23701,N_23491,N_23474);
nor U23702 (N_23702,N_23429,N_23406);
or U23703 (N_23703,N_23483,N_23305);
and U23704 (N_23704,N_23418,N_23433);
or U23705 (N_23705,N_23494,N_23309);
and U23706 (N_23706,N_23352,N_23325);
and U23707 (N_23707,N_23355,N_23362);
nand U23708 (N_23708,N_23370,N_23279);
nor U23709 (N_23709,N_23367,N_23324);
and U23710 (N_23710,N_23407,N_23324);
and U23711 (N_23711,N_23422,N_23446);
xnor U23712 (N_23712,N_23335,N_23378);
nand U23713 (N_23713,N_23473,N_23271);
nand U23714 (N_23714,N_23276,N_23476);
nor U23715 (N_23715,N_23416,N_23272);
xor U23716 (N_23716,N_23432,N_23426);
nand U23717 (N_23717,N_23341,N_23405);
or U23718 (N_23718,N_23400,N_23306);
nand U23719 (N_23719,N_23392,N_23326);
or U23720 (N_23720,N_23454,N_23364);
nor U23721 (N_23721,N_23402,N_23462);
or U23722 (N_23722,N_23276,N_23376);
and U23723 (N_23723,N_23258,N_23292);
xnor U23724 (N_23724,N_23355,N_23368);
nor U23725 (N_23725,N_23394,N_23361);
xor U23726 (N_23726,N_23256,N_23369);
or U23727 (N_23727,N_23402,N_23459);
and U23728 (N_23728,N_23331,N_23398);
nor U23729 (N_23729,N_23373,N_23484);
nor U23730 (N_23730,N_23369,N_23322);
and U23731 (N_23731,N_23311,N_23287);
and U23732 (N_23732,N_23359,N_23347);
xor U23733 (N_23733,N_23455,N_23463);
nor U23734 (N_23734,N_23355,N_23273);
and U23735 (N_23735,N_23353,N_23347);
nor U23736 (N_23736,N_23474,N_23471);
and U23737 (N_23737,N_23266,N_23425);
or U23738 (N_23738,N_23255,N_23306);
and U23739 (N_23739,N_23417,N_23283);
xnor U23740 (N_23740,N_23366,N_23463);
or U23741 (N_23741,N_23375,N_23261);
or U23742 (N_23742,N_23285,N_23424);
nor U23743 (N_23743,N_23496,N_23417);
and U23744 (N_23744,N_23289,N_23256);
xnor U23745 (N_23745,N_23455,N_23322);
nor U23746 (N_23746,N_23374,N_23336);
xor U23747 (N_23747,N_23388,N_23440);
xor U23748 (N_23748,N_23328,N_23372);
xor U23749 (N_23749,N_23348,N_23414);
nor U23750 (N_23750,N_23651,N_23673);
or U23751 (N_23751,N_23510,N_23664);
nand U23752 (N_23752,N_23554,N_23720);
xor U23753 (N_23753,N_23736,N_23520);
xor U23754 (N_23754,N_23623,N_23712);
nor U23755 (N_23755,N_23693,N_23529);
xor U23756 (N_23756,N_23618,N_23647);
and U23757 (N_23757,N_23732,N_23573);
nor U23758 (N_23758,N_23551,N_23578);
xnor U23759 (N_23759,N_23587,N_23582);
and U23760 (N_23760,N_23719,N_23624);
or U23761 (N_23761,N_23540,N_23718);
nor U23762 (N_23762,N_23592,N_23731);
nor U23763 (N_23763,N_23735,N_23509);
nor U23764 (N_23764,N_23571,N_23629);
nand U23765 (N_23765,N_23748,N_23583);
xnor U23766 (N_23766,N_23628,N_23594);
nor U23767 (N_23767,N_23641,N_23709);
nand U23768 (N_23768,N_23612,N_23625);
and U23769 (N_23769,N_23585,N_23595);
nand U23770 (N_23770,N_23560,N_23686);
and U23771 (N_23771,N_23671,N_23574);
nand U23772 (N_23772,N_23599,N_23521);
xor U23773 (N_23773,N_23701,N_23621);
nor U23774 (N_23774,N_23645,N_23603);
or U23775 (N_23775,N_23743,N_23698);
nand U23776 (N_23776,N_23607,N_23739);
or U23777 (N_23777,N_23593,N_23507);
and U23778 (N_23778,N_23663,N_23503);
xnor U23779 (N_23779,N_23675,N_23626);
and U23780 (N_23780,N_23702,N_23659);
xnor U23781 (N_23781,N_23695,N_23579);
and U23782 (N_23782,N_23559,N_23531);
or U23783 (N_23783,N_23516,N_23734);
nor U23784 (N_23784,N_23564,N_23611);
nand U23785 (N_23785,N_23569,N_23737);
or U23786 (N_23786,N_23655,N_23729);
nor U23787 (N_23787,N_23536,N_23696);
nand U23788 (N_23788,N_23544,N_23676);
or U23789 (N_23789,N_23660,N_23606);
nand U23790 (N_23790,N_23617,N_23613);
nor U23791 (N_23791,N_23545,N_23648);
or U23792 (N_23792,N_23692,N_23657);
nor U23793 (N_23793,N_23513,N_23504);
and U23794 (N_23794,N_23590,N_23668);
nand U23795 (N_23795,N_23656,N_23515);
nand U23796 (N_23796,N_23672,N_23561);
nor U23797 (N_23797,N_23608,N_23689);
and U23798 (N_23798,N_23650,N_23598);
nand U23799 (N_23799,N_23669,N_23519);
xor U23800 (N_23800,N_23722,N_23688);
and U23801 (N_23801,N_23694,N_23563);
nor U23802 (N_23802,N_23570,N_23703);
nand U23803 (N_23803,N_23550,N_23566);
nand U23804 (N_23804,N_23553,N_23605);
xor U23805 (N_23805,N_23716,N_23575);
nand U23806 (N_23806,N_23644,N_23588);
nand U23807 (N_23807,N_23584,N_23638);
nor U23808 (N_23808,N_23522,N_23725);
and U23809 (N_23809,N_23512,N_23745);
xnor U23810 (N_23810,N_23746,N_23508);
or U23811 (N_23811,N_23642,N_23741);
xor U23812 (N_23812,N_23691,N_23630);
nand U23813 (N_23813,N_23622,N_23597);
nand U23814 (N_23814,N_23604,N_23620);
nand U23815 (N_23815,N_23639,N_23723);
or U23816 (N_23816,N_23674,N_23744);
xor U23817 (N_23817,N_23601,N_23524);
xnor U23818 (N_23818,N_23511,N_23680);
and U23819 (N_23819,N_23614,N_23533);
nand U23820 (N_23820,N_23635,N_23730);
and U23821 (N_23821,N_23661,N_23558);
nor U23822 (N_23822,N_23517,N_23690);
nand U23823 (N_23823,N_23742,N_23538);
xnor U23824 (N_23824,N_23546,N_23677);
nor U23825 (N_23825,N_23683,N_23681);
nor U23826 (N_23826,N_23525,N_23537);
or U23827 (N_23827,N_23665,N_23514);
nor U23828 (N_23828,N_23717,N_23609);
or U23829 (N_23829,N_23637,N_23679);
xnor U23830 (N_23830,N_23527,N_23619);
xnor U23831 (N_23831,N_23615,N_23643);
or U23832 (N_23832,N_23653,N_23632);
nor U23833 (N_23833,N_23526,N_23721);
nand U23834 (N_23834,N_23640,N_23633);
nand U23835 (N_23835,N_23646,N_23636);
nor U23836 (N_23836,N_23714,N_23562);
nor U23837 (N_23837,N_23726,N_23530);
nand U23838 (N_23838,N_23580,N_23528);
or U23839 (N_23839,N_23749,N_23576);
and U23840 (N_23840,N_23581,N_23596);
and U23841 (N_23841,N_23577,N_23543);
and U23842 (N_23842,N_23710,N_23740);
xor U23843 (N_23843,N_23685,N_23658);
or U23844 (N_23844,N_23502,N_23738);
xor U23845 (N_23845,N_23523,N_23670);
nand U23846 (N_23846,N_23715,N_23547);
and U23847 (N_23847,N_23631,N_23567);
or U23848 (N_23848,N_23541,N_23724);
nor U23849 (N_23849,N_23542,N_23532);
nand U23850 (N_23850,N_23662,N_23500);
and U23851 (N_23851,N_23616,N_23534);
and U23852 (N_23852,N_23568,N_23687);
nor U23853 (N_23853,N_23649,N_23682);
nand U23854 (N_23854,N_23555,N_23535);
xnor U23855 (N_23855,N_23652,N_23602);
or U23856 (N_23856,N_23667,N_23700);
nor U23857 (N_23857,N_23600,N_23556);
or U23858 (N_23858,N_23549,N_23678);
nor U23859 (N_23859,N_23707,N_23684);
xnor U23860 (N_23860,N_23747,N_23589);
and U23861 (N_23861,N_23666,N_23539);
nand U23862 (N_23862,N_23711,N_23506);
nor U23863 (N_23863,N_23610,N_23697);
or U23864 (N_23864,N_23505,N_23586);
xnor U23865 (N_23865,N_23728,N_23565);
xor U23866 (N_23866,N_23733,N_23548);
nand U23867 (N_23867,N_23727,N_23704);
nand U23868 (N_23868,N_23552,N_23699);
nor U23869 (N_23869,N_23654,N_23706);
and U23870 (N_23870,N_23518,N_23708);
xor U23871 (N_23871,N_23591,N_23634);
or U23872 (N_23872,N_23713,N_23627);
or U23873 (N_23873,N_23572,N_23501);
xnor U23874 (N_23874,N_23557,N_23705);
nor U23875 (N_23875,N_23530,N_23602);
xor U23876 (N_23876,N_23569,N_23661);
and U23877 (N_23877,N_23741,N_23610);
or U23878 (N_23878,N_23533,N_23674);
or U23879 (N_23879,N_23649,N_23623);
and U23880 (N_23880,N_23745,N_23508);
nand U23881 (N_23881,N_23701,N_23727);
nor U23882 (N_23882,N_23555,N_23616);
nor U23883 (N_23883,N_23728,N_23746);
and U23884 (N_23884,N_23560,N_23676);
and U23885 (N_23885,N_23700,N_23672);
nor U23886 (N_23886,N_23552,N_23613);
nor U23887 (N_23887,N_23513,N_23557);
and U23888 (N_23888,N_23645,N_23665);
xnor U23889 (N_23889,N_23561,N_23708);
nor U23890 (N_23890,N_23738,N_23653);
and U23891 (N_23891,N_23692,N_23530);
nand U23892 (N_23892,N_23662,N_23507);
nand U23893 (N_23893,N_23531,N_23691);
xor U23894 (N_23894,N_23575,N_23618);
xor U23895 (N_23895,N_23673,N_23542);
nand U23896 (N_23896,N_23728,N_23711);
or U23897 (N_23897,N_23557,N_23689);
or U23898 (N_23898,N_23546,N_23562);
xnor U23899 (N_23899,N_23642,N_23656);
and U23900 (N_23900,N_23673,N_23520);
xnor U23901 (N_23901,N_23687,N_23585);
nor U23902 (N_23902,N_23508,N_23574);
or U23903 (N_23903,N_23558,N_23744);
nand U23904 (N_23904,N_23568,N_23645);
xnor U23905 (N_23905,N_23645,N_23535);
nand U23906 (N_23906,N_23648,N_23516);
nand U23907 (N_23907,N_23553,N_23635);
and U23908 (N_23908,N_23537,N_23633);
or U23909 (N_23909,N_23500,N_23602);
xor U23910 (N_23910,N_23638,N_23535);
nand U23911 (N_23911,N_23712,N_23658);
nor U23912 (N_23912,N_23558,N_23536);
nand U23913 (N_23913,N_23691,N_23524);
and U23914 (N_23914,N_23744,N_23711);
xor U23915 (N_23915,N_23579,N_23660);
or U23916 (N_23916,N_23647,N_23742);
or U23917 (N_23917,N_23623,N_23526);
nand U23918 (N_23918,N_23514,N_23634);
xor U23919 (N_23919,N_23580,N_23723);
and U23920 (N_23920,N_23628,N_23607);
or U23921 (N_23921,N_23551,N_23584);
or U23922 (N_23922,N_23734,N_23619);
nor U23923 (N_23923,N_23572,N_23556);
nand U23924 (N_23924,N_23632,N_23565);
nor U23925 (N_23925,N_23685,N_23538);
nand U23926 (N_23926,N_23545,N_23746);
or U23927 (N_23927,N_23553,N_23501);
nor U23928 (N_23928,N_23714,N_23624);
nand U23929 (N_23929,N_23592,N_23692);
and U23930 (N_23930,N_23601,N_23712);
nand U23931 (N_23931,N_23607,N_23510);
and U23932 (N_23932,N_23563,N_23661);
xor U23933 (N_23933,N_23645,N_23705);
and U23934 (N_23934,N_23600,N_23673);
nand U23935 (N_23935,N_23544,N_23696);
and U23936 (N_23936,N_23704,N_23588);
nand U23937 (N_23937,N_23681,N_23570);
nor U23938 (N_23938,N_23716,N_23551);
nand U23939 (N_23939,N_23578,N_23575);
or U23940 (N_23940,N_23729,N_23649);
and U23941 (N_23941,N_23691,N_23654);
nand U23942 (N_23942,N_23632,N_23735);
or U23943 (N_23943,N_23709,N_23535);
xor U23944 (N_23944,N_23734,N_23636);
and U23945 (N_23945,N_23608,N_23592);
and U23946 (N_23946,N_23727,N_23604);
nor U23947 (N_23947,N_23517,N_23651);
nor U23948 (N_23948,N_23538,N_23635);
or U23949 (N_23949,N_23666,N_23660);
and U23950 (N_23950,N_23559,N_23684);
nor U23951 (N_23951,N_23690,N_23571);
nor U23952 (N_23952,N_23747,N_23504);
nand U23953 (N_23953,N_23514,N_23692);
or U23954 (N_23954,N_23735,N_23650);
xor U23955 (N_23955,N_23600,N_23646);
nor U23956 (N_23956,N_23546,N_23540);
or U23957 (N_23957,N_23651,N_23505);
nand U23958 (N_23958,N_23523,N_23537);
and U23959 (N_23959,N_23547,N_23738);
nand U23960 (N_23960,N_23588,N_23592);
xor U23961 (N_23961,N_23533,N_23682);
xor U23962 (N_23962,N_23686,N_23666);
and U23963 (N_23963,N_23567,N_23503);
or U23964 (N_23964,N_23744,N_23670);
nand U23965 (N_23965,N_23562,N_23746);
xor U23966 (N_23966,N_23739,N_23710);
xnor U23967 (N_23967,N_23661,N_23722);
nor U23968 (N_23968,N_23542,N_23740);
nand U23969 (N_23969,N_23667,N_23707);
xor U23970 (N_23970,N_23550,N_23602);
and U23971 (N_23971,N_23697,N_23628);
nand U23972 (N_23972,N_23529,N_23502);
nor U23973 (N_23973,N_23504,N_23515);
xor U23974 (N_23974,N_23650,N_23571);
nand U23975 (N_23975,N_23631,N_23747);
or U23976 (N_23976,N_23749,N_23541);
or U23977 (N_23977,N_23743,N_23568);
nor U23978 (N_23978,N_23581,N_23683);
or U23979 (N_23979,N_23695,N_23614);
xnor U23980 (N_23980,N_23747,N_23742);
xnor U23981 (N_23981,N_23653,N_23663);
nor U23982 (N_23982,N_23620,N_23741);
nor U23983 (N_23983,N_23657,N_23506);
nor U23984 (N_23984,N_23590,N_23637);
nand U23985 (N_23985,N_23729,N_23546);
and U23986 (N_23986,N_23595,N_23668);
or U23987 (N_23987,N_23516,N_23728);
nand U23988 (N_23988,N_23710,N_23656);
and U23989 (N_23989,N_23699,N_23707);
nor U23990 (N_23990,N_23653,N_23731);
and U23991 (N_23991,N_23568,N_23624);
or U23992 (N_23992,N_23739,N_23566);
and U23993 (N_23993,N_23635,N_23527);
and U23994 (N_23994,N_23546,N_23675);
nand U23995 (N_23995,N_23609,N_23531);
nor U23996 (N_23996,N_23634,N_23719);
and U23997 (N_23997,N_23642,N_23541);
nor U23998 (N_23998,N_23711,N_23646);
xnor U23999 (N_23999,N_23600,N_23518);
xnor U24000 (N_24000,N_23991,N_23761);
xnor U24001 (N_24001,N_23835,N_23911);
nor U24002 (N_24002,N_23984,N_23905);
or U24003 (N_24003,N_23955,N_23958);
nand U24004 (N_24004,N_23816,N_23933);
xnor U24005 (N_24005,N_23777,N_23756);
or U24006 (N_24006,N_23819,N_23899);
nand U24007 (N_24007,N_23996,N_23898);
and U24008 (N_24008,N_23919,N_23827);
or U24009 (N_24009,N_23948,N_23815);
nor U24010 (N_24010,N_23963,N_23811);
nor U24011 (N_24011,N_23823,N_23800);
nor U24012 (N_24012,N_23754,N_23786);
xor U24013 (N_24013,N_23821,N_23913);
or U24014 (N_24014,N_23975,N_23771);
nor U24015 (N_24015,N_23829,N_23844);
and U24016 (N_24016,N_23953,N_23998);
nand U24017 (N_24017,N_23792,N_23950);
and U24018 (N_24018,N_23971,N_23988);
nand U24019 (N_24019,N_23863,N_23876);
and U24020 (N_24020,N_23799,N_23967);
or U24021 (N_24021,N_23832,N_23989);
nor U24022 (N_24022,N_23782,N_23865);
nor U24023 (N_24023,N_23893,N_23891);
xnor U24024 (N_24024,N_23968,N_23951);
xnor U24025 (N_24025,N_23766,N_23838);
nor U24026 (N_24026,N_23872,N_23980);
and U24027 (N_24027,N_23793,N_23780);
or U24028 (N_24028,N_23914,N_23791);
xor U24029 (N_24029,N_23803,N_23887);
xnor U24030 (N_24030,N_23855,N_23824);
and U24031 (N_24031,N_23931,N_23957);
nand U24032 (N_24032,N_23755,N_23941);
nand U24033 (N_24033,N_23882,N_23928);
xor U24034 (N_24034,N_23814,N_23836);
xor U24035 (N_24035,N_23994,N_23770);
xor U24036 (N_24036,N_23779,N_23869);
nand U24037 (N_24037,N_23973,N_23859);
xnor U24038 (N_24038,N_23896,N_23825);
and U24039 (N_24039,N_23888,N_23810);
or U24040 (N_24040,N_23813,N_23778);
nor U24041 (N_24041,N_23912,N_23759);
nand U24042 (N_24042,N_23993,N_23828);
or U24043 (N_24043,N_23812,N_23972);
or U24044 (N_24044,N_23842,N_23806);
xor U24045 (N_24045,N_23760,N_23808);
nand U24046 (N_24046,N_23880,N_23797);
nand U24047 (N_24047,N_23879,N_23979);
nand U24048 (N_24048,N_23839,N_23868);
or U24049 (N_24049,N_23921,N_23944);
or U24050 (N_24050,N_23978,N_23752);
nand U24051 (N_24051,N_23932,N_23907);
xor U24052 (N_24052,N_23866,N_23751);
nor U24053 (N_24053,N_23787,N_23852);
nor U24054 (N_24054,N_23794,N_23917);
nor U24055 (N_24055,N_23774,N_23795);
or U24056 (N_24056,N_23938,N_23940);
nand U24057 (N_24057,N_23764,N_23909);
xnor U24058 (N_24058,N_23897,N_23850);
nor U24059 (N_24059,N_23822,N_23943);
and U24060 (N_24060,N_23769,N_23790);
nand U24061 (N_24061,N_23809,N_23892);
nand U24062 (N_24062,N_23826,N_23930);
or U24063 (N_24063,N_23960,N_23925);
xor U24064 (N_24064,N_23853,N_23776);
or U24065 (N_24065,N_23935,N_23884);
xor U24066 (N_24066,N_23981,N_23956);
nor U24067 (N_24067,N_23757,N_23871);
xnor U24068 (N_24068,N_23762,N_23966);
or U24069 (N_24069,N_23934,N_23758);
nand U24070 (N_24070,N_23999,N_23773);
and U24071 (N_24071,N_23901,N_23954);
xor U24072 (N_24072,N_23937,N_23987);
xor U24073 (N_24073,N_23969,N_23847);
xor U24074 (N_24074,N_23986,N_23923);
or U24075 (N_24075,N_23936,N_23830);
nand U24076 (N_24076,N_23873,N_23801);
or U24077 (N_24077,N_23962,N_23854);
or U24078 (N_24078,N_23772,N_23906);
or U24079 (N_24079,N_23817,N_23789);
nor U24080 (N_24080,N_23878,N_23807);
or U24081 (N_24081,N_23886,N_23894);
or U24082 (N_24082,N_23964,N_23851);
nand U24083 (N_24083,N_23946,N_23983);
nand U24084 (N_24084,N_23804,N_23834);
xnor U24085 (N_24085,N_23920,N_23856);
or U24086 (N_24086,N_23805,N_23915);
nor U24087 (N_24087,N_23942,N_23970);
and U24088 (N_24088,N_23885,N_23831);
or U24089 (N_24089,N_23883,N_23939);
xnor U24090 (N_24090,N_23837,N_23961);
nor U24091 (N_24091,N_23867,N_23904);
and U24092 (N_24092,N_23916,N_23900);
or U24093 (N_24093,N_23848,N_23802);
and U24094 (N_24094,N_23902,N_23875);
and U24095 (N_24095,N_23908,N_23788);
and U24096 (N_24096,N_23889,N_23768);
nand U24097 (N_24097,N_23895,N_23995);
nand U24098 (N_24098,N_23820,N_23997);
xor U24099 (N_24099,N_23862,N_23903);
and U24100 (N_24100,N_23924,N_23796);
and U24101 (N_24101,N_23949,N_23929);
nor U24102 (N_24102,N_23841,N_23861);
nand U24103 (N_24103,N_23977,N_23785);
nor U24104 (N_24104,N_23767,N_23874);
nand U24105 (N_24105,N_23976,N_23910);
nand U24106 (N_24106,N_23982,N_23840);
and U24107 (N_24107,N_23974,N_23945);
and U24108 (N_24108,N_23753,N_23927);
nor U24109 (N_24109,N_23833,N_23858);
nand U24110 (N_24110,N_23843,N_23922);
and U24111 (N_24111,N_23959,N_23952);
xnor U24112 (N_24112,N_23881,N_23947);
or U24113 (N_24113,N_23890,N_23845);
or U24114 (N_24114,N_23781,N_23783);
nor U24115 (N_24115,N_23992,N_23763);
or U24116 (N_24116,N_23965,N_23926);
xnor U24117 (N_24117,N_23849,N_23798);
nand U24118 (N_24118,N_23864,N_23990);
nor U24119 (N_24119,N_23846,N_23860);
and U24120 (N_24120,N_23775,N_23750);
xnor U24121 (N_24121,N_23918,N_23818);
or U24122 (N_24122,N_23877,N_23985);
nand U24123 (N_24123,N_23765,N_23857);
or U24124 (N_24124,N_23784,N_23870);
or U24125 (N_24125,N_23979,N_23962);
xnor U24126 (N_24126,N_23914,N_23979);
xor U24127 (N_24127,N_23758,N_23846);
or U24128 (N_24128,N_23964,N_23814);
nand U24129 (N_24129,N_23835,N_23931);
or U24130 (N_24130,N_23821,N_23861);
nand U24131 (N_24131,N_23879,N_23926);
and U24132 (N_24132,N_23998,N_23795);
and U24133 (N_24133,N_23883,N_23904);
xnor U24134 (N_24134,N_23954,N_23775);
and U24135 (N_24135,N_23840,N_23919);
xor U24136 (N_24136,N_23870,N_23843);
nor U24137 (N_24137,N_23811,N_23912);
xor U24138 (N_24138,N_23848,N_23878);
and U24139 (N_24139,N_23965,N_23861);
nor U24140 (N_24140,N_23862,N_23986);
xor U24141 (N_24141,N_23893,N_23833);
and U24142 (N_24142,N_23948,N_23930);
nor U24143 (N_24143,N_23885,N_23960);
nand U24144 (N_24144,N_23886,N_23837);
and U24145 (N_24145,N_23808,N_23803);
or U24146 (N_24146,N_23879,N_23934);
xor U24147 (N_24147,N_23878,N_23950);
nand U24148 (N_24148,N_23791,N_23906);
nand U24149 (N_24149,N_23949,N_23773);
nor U24150 (N_24150,N_23927,N_23883);
nor U24151 (N_24151,N_23960,N_23758);
nor U24152 (N_24152,N_23967,N_23981);
xnor U24153 (N_24153,N_23828,N_23907);
xor U24154 (N_24154,N_23781,N_23923);
xor U24155 (N_24155,N_23948,N_23789);
and U24156 (N_24156,N_23763,N_23995);
nor U24157 (N_24157,N_23961,N_23885);
or U24158 (N_24158,N_23840,N_23996);
nand U24159 (N_24159,N_23780,N_23796);
nand U24160 (N_24160,N_23773,N_23864);
nand U24161 (N_24161,N_23775,N_23764);
nand U24162 (N_24162,N_23850,N_23915);
nor U24163 (N_24163,N_23807,N_23870);
nor U24164 (N_24164,N_23771,N_23799);
and U24165 (N_24165,N_23885,N_23841);
or U24166 (N_24166,N_23949,N_23999);
or U24167 (N_24167,N_23811,N_23819);
xnor U24168 (N_24168,N_23828,N_23836);
nand U24169 (N_24169,N_23831,N_23994);
nand U24170 (N_24170,N_23940,N_23772);
nor U24171 (N_24171,N_23820,N_23870);
and U24172 (N_24172,N_23753,N_23834);
xnor U24173 (N_24173,N_23814,N_23825);
or U24174 (N_24174,N_23760,N_23867);
or U24175 (N_24175,N_23909,N_23888);
or U24176 (N_24176,N_23875,N_23897);
nand U24177 (N_24177,N_23776,N_23944);
or U24178 (N_24178,N_23919,N_23881);
nor U24179 (N_24179,N_23975,N_23887);
or U24180 (N_24180,N_23966,N_23977);
nand U24181 (N_24181,N_23820,N_23764);
xor U24182 (N_24182,N_23925,N_23785);
and U24183 (N_24183,N_23992,N_23816);
nand U24184 (N_24184,N_23864,N_23948);
xor U24185 (N_24185,N_23841,N_23938);
xnor U24186 (N_24186,N_23756,N_23998);
nand U24187 (N_24187,N_23899,N_23982);
nand U24188 (N_24188,N_23828,N_23751);
xnor U24189 (N_24189,N_23844,N_23810);
nor U24190 (N_24190,N_23974,N_23810);
or U24191 (N_24191,N_23803,N_23962);
nand U24192 (N_24192,N_23861,N_23801);
nand U24193 (N_24193,N_23900,N_23788);
nor U24194 (N_24194,N_23868,N_23829);
nand U24195 (N_24195,N_23903,N_23933);
and U24196 (N_24196,N_23980,N_23763);
nand U24197 (N_24197,N_23936,N_23946);
or U24198 (N_24198,N_23902,N_23819);
xnor U24199 (N_24199,N_23920,N_23898);
and U24200 (N_24200,N_23913,N_23908);
nand U24201 (N_24201,N_23896,N_23833);
xor U24202 (N_24202,N_23893,N_23804);
xnor U24203 (N_24203,N_23884,N_23826);
xnor U24204 (N_24204,N_23833,N_23956);
and U24205 (N_24205,N_23896,N_23767);
or U24206 (N_24206,N_23985,N_23781);
or U24207 (N_24207,N_23820,N_23834);
xor U24208 (N_24208,N_23841,N_23770);
nand U24209 (N_24209,N_23981,N_23969);
xor U24210 (N_24210,N_23845,N_23911);
xor U24211 (N_24211,N_23766,N_23912);
nor U24212 (N_24212,N_23961,N_23946);
or U24213 (N_24213,N_23772,N_23818);
or U24214 (N_24214,N_23936,N_23758);
nand U24215 (N_24215,N_23757,N_23754);
or U24216 (N_24216,N_23926,N_23813);
and U24217 (N_24217,N_23825,N_23885);
nor U24218 (N_24218,N_23838,N_23920);
and U24219 (N_24219,N_23971,N_23775);
and U24220 (N_24220,N_23875,N_23809);
nor U24221 (N_24221,N_23823,N_23805);
and U24222 (N_24222,N_23829,N_23892);
xnor U24223 (N_24223,N_23885,N_23824);
nor U24224 (N_24224,N_23809,N_23798);
or U24225 (N_24225,N_23772,N_23830);
and U24226 (N_24226,N_23786,N_23825);
nor U24227 (N_24227,N_23958,N_23950);
and U24228 (N_24228,N_23862,N_23904);
and U24229 (N_24229,N_23999,N_23945);
or U24230 (N_24230,N_23765,N_23892);
or U24231 (N_24231,N_23826,N_23870);
nand U24232 (N_24232,N_23771,N_23896);
or U24233 (N_24233,N_23757,N_23891);
or U24234 (N_24234,N_23982,N_23873);
and U24235 (N_24235,N_23823,N_23813);
or U24236 (N_24236,N_23793,N_23998);
and U24237 (N_24237,N_23899,N_23956);
xor U24238 (N_24238,N_23775,N_23889);
and U24239 (N_24239,N_23811,N_23844);
and U24240 (N_24240,N_23792,N_23819);
and U24241 (N_24241,N_23768,N_23984);
nor U24242 (N_24242,N_23922,N_23758);
nor U24243 (N_24243,N_23770,N_23765);
or U24244 (N_24244,N_23949,N_23878);
nor U24245 (N_24245,N_23756,N_23792);
or U24246 (N_24246,N_23947,N_23938);
or U24247 (N_24247,N_23767,N_23964);
nand U24248 (N_24248,N_23894,N_23827);
and U24249 (N_24249,N_23926,N_23793);
nand U24250 (N_24250,N_24069,N_24094);
nand U24251 (N_24251,N_24001,N_24196);
nand U24252 (N_24252,N_24118,N_24065);
nand U24253 (N_24253,N_24029,N_24004);
or U24254 (N_24254,N_24114,N_24047);
and U24255 (N_24255,N_24015,N_24005);
or U24256 (N_24256,N_24055,N_24040);
nand U24257 (N_24257,N_24107,N_24221);
nor U24258 (N_24258,N_24081,N_24038);
and U24259 (N_24259,N_24009,N_24162);
nand U24260 (N_24260,N_24100,N_24138);
nand U24261 (N_24261,N_24084,N_24195);
nand U24262 (N_24262,N_24068,N_24191);
nor U24263 (N_24263,N_24048,N_24067);
or U24264 (N_24264,N_24145,N_24152);
or U24265 (N_24265,N_24211,N_24245);
nand U24266 (N_24266,N_24165,N_24166);
or U24267 (N_24267,N_24051,N_24089);
nor U24268 (N_24268,N_24173,N_24183);
and U24269 (N_24269,N_24144,N_24192);
nor U24270 (N_24270,N_24151,N_24200);
nor U24271 (N_24271,N_24185,N_24000);
xor U24272 (N_24272,N_24031,N_24225);
xnor U24273 (N_24273,N_24063,N_24128);
nor U24274 (N_24274,N_24207,N_24135);
xnor U24275 (N_24275,N_24073,N_24208);
or U24276 (N_24276,N_24109,N_24229);
xor U24277 (N_24277,N_24216,N_24056);
xnor U24278 (N_24278,N_24086,N_24214);
nand U24279 (N_24279,N_24101,N_24045);
nand U24280 (N_24280,N_24062,N_24235);
xnor U24281 (N_24281,N_24198,N_24240);
xor U24282 (N_24282,N_24012,N_24156);
nor U24283 (N_24283,N_24044,N_24078);
nand U24284 (N_24284,N_24110,N_24137);
nand U24285 (N_24285,N_24028,N_24233);
nor U24286 (N_24286,N_24231,N_24034);
and U24287 (N_24287,N_24075,N_24142);
nor U24288 (N_24288,N_24121,N_24146);
and U24289 (N_24289,N_24061,N_24008);
and U24290 (N_24290,N_24213,N_24210);
or U24291 (N_24291,N_24037,N_24134);
nand U24292 (N_24292,N_24096,N_24017);
and U24293 (N_24293,N_24125,N_24158);
and U24294 (N_24294,N_24083,N_24120);
nor U24295 (N_24295,N_24176,N_24030);
xor U24296 (N_24296,N_24197,N_24126);
nor U24297 (N_24297,N_24088,N_24180);
or U24298 (N_24298,N_24018,N_24164);
or U24299 (N_24299,N_24204,N_24168);
or U24300 (N_24300,N_24172,N_24133);
xnor U24301 (N_24301,N_24169,N_24190);
nand U24302 (N_24302,N_24112,N_24021);
or U24303 (N_24303,N_24102,N_24220);
nor U24304 (N_24304,N_24182,N_24087);
nand U24305 (N_24305,N_24074,N_24085);
xnor U24306 (N_24306,N_24022,N_24226);
or U24307 (N_24307,N_24111,N_24239);
and U24308 (N_24308,N_24052,N_24103);
xnor U24309 (N_24309,N_24219,N_24064);
nor U24310 (N_24310,N_24049,N_24193);
xnor U24311 (N_24311,N_24035,N_24202);
nand U24312 (N_24312,N_24227,N_24179);
nand U24313 (N_24313,N_24006,N_24071);
xor U24314 (N_24314,N_24247,N_24119);
and U24315 (N_24315,N_24080,N_24141);
nand U24316 (N_24316,N_24242,N_24025);
xor U24317 (N_24317,N_24236,N_24186);
xnor U24318 (N_24318,N_24076,N_24150);
nand U24319 (N_24319,N_24178,N_24091);
xnor U24320 (N_24320,N_24127,N_24149);
or U24321 (N_24321,N_24093,N_24123);
and U24322 (N_24322,N_24050,N_24222);
or U24323 (N_24323,N_24209,N_24011);
nand U24324 (N_24324,N_24206,N_24113);
or U24325 (N_24325,N_24181,N_24013);
nor U24326 (N_24326,N_24010,N_24224);
and U24327 (N_24327,N_24058,N_24212);
nor U24328 (N_24328,N_24019,N_24187);
nor U24329 (N_24329,N_24249,N_24147);
nor U24330 (N_24330,N_24136,N_24124);
nor U24331 (N_24331,N_24131,N_24027);
xor U24332 (N_24332,N_24203,N_24023);
nor U24333 (N_24333,N_24170,N_24041);
nor U24334 (N_24334,N_24189,N_24230);
and U24335 (N_24335,N_24108,N_24097);
xor U24336 (N_24336,N_24014,N_24139);
nand U24337 (N_24337,N_24057,N_24223);
and U24338 (N_24338,N_24153,N_24199);
nor U24339 (N_24339,N_24082,N_24092);
nand U24340 (N_24340,N_24159,N_24218);
and U24341 (N_24341,N_24154,N_24248);
and U24342 (N_24342,N_24188,N_24116);
xnor U24343 (N_24343,N_24059,N_24043);
xor U24344 (N_24344,N_24140,N_24237);
nand U24345 (N_24345,N_24175,N_24234);
nor U24346 (N_24346,N_24115,N_24066);
and U24347 (N_24347,N_24167,N_24184);
nand U24348 (N_24348,N_24143,N_24130);
nor U24349 (N_24349,N_24042,N_24106);
xnor U24350 (N_24350,N_24228,N_24217);
and U24351 (N_24351,N_24243,N_24174);
xnor U24352 (N_24352,N_24077,N_24104);
and U24353 (N_24353,N_24046,N_24155);
xor U24354 (N_24354,N_24238,N_24244);
nand U24355 (N_24355,N_24194,N_24007);
and U24356 (N_24356,N_24160,N_24079);
nand U24357 (N_24357,N_24036,N_24129);
xnor U24358 (N_24358,N_24163,N_24072);
nor U24359 (N_24359,N_24132,N_24098);
and U24360 (N_24360,N_24033,N_24117);
or U24361 (N_24361,N_24032,N_24157);
nor U24362 (N_24362,N_24020,N_24024);
nor U24363 (N_24363,N_24201,N_24241);
nand U24364 (N_24364,N_24090,N_24105);
nand U24365 (N_24365,N_24026,N_24002);
nor U24366 (N_24366,N_24122,N_24177);
and U24367 (N_24367,N_24054,N_24003);
nand U24368 (N_24368,N_24099,N_24095);
nand U24369 (N_24369,N_24161,N_24171);
nand U24370 (N_24370,N_24039,N_24246);
and U24371 (N_24371,N_24053,N_24205);
or U24372 (N_24372,N_24016,N_24232);
and U24373 (N_24373,N_24060,N_24148);
and U24374 (N_24374,N_24070,N_24215);
and U24375 (N_24375,N_24052,N_24070);
xnor U24376 (N_24376,N_24091,N_24097);
nor U24377 (N_24377,N_24005,N_24078);
and U24378 (N_24378,N_24008,N_24203);
xnor U24379 (N_24379,N_24181,N_24093);
nor U24380 (N_24380,N_24008,N_24152);
and U24381 (N_24381,N_24183,N_24032);
or U24382 (N_24382,N_24130,N_24121);
xnor U24383 (N_24383,N_24232,N_24203);
nand U24384 (N_24384,N_24200,N_24041);
or U24385 (N_24385,N_24182,N_24212);
nor U24386 (N_24386,N_24023,N_24013);
and U24387 (N_24387,N_24157,N_24164);
xnor U24388 (N_24388,N_24106,N_24069);
nor U24389 (N_24389,N_24048,N_24215);
nand U24390 (N_24390,N_24097,N_24198);
or U24391 (N_24391,N_24125,N_24197);
xor U24392 (N_24392,N_24164,N_24118);
and U24393 (N_24393,N_24160,N_24238);
and U24394 (N_24394,N_24131,N_24188);
or U24395 (N_24395,N_24121,N_24074);
and U24396 (N_24396,N_24015,N_24164);
xnor U24397 (N_24397,N_24002,N_24153);
xor U24398 (N_24398,N_24034,N_24184);
nor U24399 (N_24399,N_24148,N_24230);
or U24400 (N_24400,N_24143,N_24200);
nor U24401 (N_24401,N_24016,N_24076);
xnor U24402 (N_24402,N_24226,N_24186);
or U24403 (N_24403,N_24046,N_24022);
nor U24404 (N_24404,N_24061,N_24185);
nand U24405 (N_24405,N_24059,N_24237);
nor U24406 (N_24406,N_24190,N_24029);
xor U24407 (N_24407,N_24150,N_24185);
xor U24408 (N_24408,N_24177,N_24087);
and U24409 (N_24409,N_24090,N_24115);
and U24410 (N_24410,N_24157,N_24178);
xnor U24411 (N_24411,N_24035,N_24044);
nor U24412 (N_24412,N_24218,N_24148);
nand U24413 (N_24413,N_24167,N_24247);
and U24414 (N_24414,N_24150,N_24024);
nor U24415 (N_24415,N_24163,N_24120);
xor U24416 (N_24416,N_24190,N_24104);
and U24417 (N_24417,N_24162,N_24146);
xor U24418 (N_24418,N_24025,N_24057);
and U24419 (N_24419,N_24138,N_24131);
xor U24420 (N_24420,N_24065,N_24087);
or U24421 (N_24421,N_24151,N_24035);
and U24422 (N_24422,N_24062,N_24195);
and U24423 (N_24423,N_24033,N_24229);
xor U24424 (N_24424,N_24189,N_24103);
and U24425 (N_24425,N_24038,N_24192);
xnor U24426 (N_24426,N_24194,N_24060);
xnor U24427 (N_24427,N_24092,N_24192);
nor U24428 (N_24428,N_24162,N_24014);
nor U24429 (N_24429,N_24237,N_24040);
nand U24430 (N_24430,N_24110,N_24045);
or U24431 (N_24431,N_24177,N_24207);
and U24432 (N_24432,N_24044,N_24002);
nor U24433 (N_24433,N_24132,N_24111);
xor U24434 (N_24434,N_24239,N_24196);
and U24435 (N_24435,N_24131,N_24082);
and U24436 (N_24436,N_24236,N_24224);
or U24437 (N_24437,N_24131,N_24137);
xnor U24438 (N_24438,N_24184,N_24074);
and U24439 (N_24439,N_24048,N_24210);
or U24440 (N_24440,N_24242,N_24101);
and U24441 (N_24441,N_24035,N_24166);
nand U24442 (N_24442,N_24108,N_24060);
nor U24443 (N_24443,N_24049,N_24228);
nand U24444 (N_24444,N_24196,N_24172);
and U24445 (N_24445,N_24048,N_24046);
nand U24446 (N_24446,N_24161,N_24229);
and U24447 (N_24447,N_24165,N_24070);
nor U24448 (N_24448,N_24227,N_24115);
and U24449 (N_24449,N_24118,N_24009);
nand U24450 (N_24450,N_24104,N_24129);
and U24451 (N_24451,N_24183,N_24003);
or U24452 (N_24452,N_24208,N_24236);
or U24453 (N_24453,N_24040,N_24203);
nor U24454 (N_24454,N_24097,N_24137);
xor U24455 (N_24455,N_24089,N_24017);
and U24456 (N_24456,N_24154,N_24052);
and U24457 (N_24457,N_24219,N_24198);
and U24458 (N_24458,N_24111,N_24192);
nand U24459 (N_24459,N_24102,N_24180);
or U24460 (N_24460,N_24170,N_24113);
xnor U24461 (N_24461,N_24217,N_24063);
xnor U24462 (N_24462,N_24001,N_24232);
or U24463 (N_24463,N_24207,N_24068);
and U24464 (N_24464,N_24188,N_24004);
xor U24465 (N_24465,N_24070,N_24118);
or U24466 (N_24466,N_24064,N_24043);
nand U24467 (N_24467,N_24000,N_24238);
nor U24468 (N_24468,N_24011,N_24056);
nor U24469 (N_24469,N_24103,N_24055);
xor U24470 (N_24470,N_24063,N_24228);
nand U24471 (N_24471,N_24081,N_24129);
and U24472 (N_24472,N_24117,N_24147);
nor U24473 (N_24473,N_24039,N_24048);
nor U24474 (N_24474,N_24236,N_24180);
nor U24475 (N_24475,N_24049,N_24100);
and U24476 (N_24476,N_24235,N_24241);
or U24477 (N_24477,N_24136,N_24192);
xnor U24478 (N_24478,N_24034,N_24022);
xnor U24479 (N_24479,N_24088,N_24162);
xnor U24480 (N_24480,N_24198,N_24145);
xnor U24481 (N_24481,N_24135,N_24122);
and U24482 (N_24482,N_24182,N_24232);
and U24483 (N_24483,N_24243,N_24192);
and U24484 (N_24484,N_24142,N_24194);
and U24485 (N_24485,N_24128,N_24238);
nor U24486 (N_24486,N_24193,N_24064);
nand U24487 (N_24487,N_24244,N_24199);
or U24488 (N_24488,N_24031,N_24174);
xnor U24489 (N_24489,N_24075,N_24221);
and U24490 (N_24490,N_24221,N_24141);
nor U24491 (N_24491,N_24233,N_24228);
xor U24492 (N_24492,N_24121,N_24132);
xor U24493 (N_24493,N_24133,N_24046);
or U24494 (N_24494,N_24023,N_24162);
xnor U24495 (N_24495,N_24017,N_24170);
nand U24496 (N_24496,N_24134,N_24072);
nor U24497 (N_24497,N_24192,N_24082);
and U24498 (N_24498,N_24045,N_24135);
and U24499 (N_24499,N_24011,N_24092);
nor U24500 (N_24500,N_24492,N_24331);
and U24501 (N_24501,N_24474,N_24396);
xnor U24502 (N_24502,N_24340,N_24329);
nor U24503 (N_24503,N_24481,N_24393);
or U24504 (N_24504,N_24425,N_24464);
or U24505 (N_24505,N_24364,N_24388);
and U24506 (N_24506,N_24321,N_24433);
and U24507 (N_24507,N_24450,N_24440);
nor U24508 (N_24508,N_24298,N_24273);
and U24509 (N_24509,N_24315,N_24429);
and U24510 (N_24510,N_24477,N_24437);
or U24511 (N_24511,N_24270,N_24407);
or U24512 (N_24512,N_24356,N_24443);
nand U24513 (N_24513,N_24381,N_24318);
xor U24514 (N_24514,N_24498,N_24430);
nor U24515 (N_24515,N_24304,N_24328);
or U24516 (N_24516,N_24322,N_24269);
xnor U24517 (N_24517,N_24264,N_24416);
and U24518 (N_24518,N_24278,N_24451);
or U24519 (N_24519,N_24365,N_24403);
and U24520 (N_24520,N_24449,N_24341);
and U24521 (N_24521,N_24327,N_24380);
nand U24522 (N_24522,N_24293,N_24376);
xor U24523 (N_24523,N_24342,N_24374);
and U24524 (N_24524,N_24409,N_24350);
nand U24525 (N_24525,N_24476,N_24307);
xor U24526 (N_24526,N_24339,N_24463);
or U24527 (N_24527,N_24317,N_24326);
xnor U24528 (N_24528,N_24370,N_24490);
and U24529 (N_24529,N_24466,N_24306);
nand U24530 (N_24530,N_24284,N_24468);
nor U24531 (N_24531,N_24420,N_24457);
and U24532 (N_24532,N_24442,N_24296);
nand U24533 (N_24533,N_24413,N_24387);
nor U24534 (N_24534,N_24358,N_24294);
nand U24535 (N_24535,N_24461,N_24299);
nand U24536 (N_24536,N_24343,N_24495);
or U24537 (N_24537,N_24265,N_24372);
nand U24538 (N_24538,N_24333,N_24336);
xor U24539 (N_24539,N_24494,N_24484);
or U24540 (N_24540,N_24319,N_24362);
xor U24541 (N_24541,N_24368,N_24489);
xnor U24542 (N_24542,N_24311,N_24282);
or U24543 (N_24543,N_24330,N_24470);
nor U24544 (N_24544,N_24262,N_24371);
xnor U24545 (N_24545,N_24472,N_24422);
and U24546 (N_24546,N_24428,N_24438);
nand U24547 (N_24547,N_24346,N_24354);
nand U24548 (N_24548,N_24455,N_24395);
and U24549 (N_24549,N_24272,N_24274);
nand U24550 (N_24550,N_24255,N_24454);
or U24551 (N_24551,N_24259,N_24250);
or U24552 (N_24552,N_24447,N_24493);
nor U24553 (N_24553,N_24335,N_24448);
nor U24554 (N_24554,N_24369,N_24267);
nor U24555 (N_24555,N_24431,N_24404);
nor U24556 (N_24556,N_24302,N_24479);
and U24557 (N_24557,N_24486,N_24436);
or U24558 (N_24558,N_24414,N_24383);
nand U24559 (N_24559,N_24456,N_24256);
xor U24560 (N_24560,N_24263,N_24410);
nand U24561 (N_24561,N_24465,N_24287);
xnor U24562 (N_24562,N_24444,N_24497);
nand U24563 (N_24563,N_24300,N_24399);
or U24564 (N_24564,N_24295,N_24441);
nand U24565 (N_24565,N_24459,N_24355);
xor U24566 (N_24566,N_24347,N_24288);
nor U24567 (N_24567,N_24320,N_24310);
and U24568 (N_24568,N_24367,N_24412);
and U24569 (N_24569,N_24392,N_24427);
xnor U24570 (N_24570,N_24480,N_24338);
nor U24571 (N_24571,N_24312,N_24289);
xor U24572 (N_24572,N_24475,N_24488);
xor U24573 (N_24573,N_24446,N_24453);
xor U24574 (N_24574,N_24401,N_24268);
and U24575 (N_24575,N_24275,N_24276);
or U24576 (N_24576,N_24290,N_24258);
or U24577 (N_24577,N_24394,N_24345);
or U24578 (N_24578,N_24499,N_24277);
xor U24579 (N_24579,N_24485,N_24373);
xnor U24580 (N_24580,N_24309,N_24389);
nor U24581 (N_24581,N_24297,N_24363);
nand U24582 (N_24582,N_24419,N_24421);
xnor U24583 (N_24583,N_24266,N_24406);
and U24584 (N_24584,N_24254,N_24286);
or U24585 (N_24585,N_24400,N_24252);
nor U24586 (N_24586,N_24467,N_24473);
or U24587 (N_24587,N_24432,N_24397);
nand U24588 (N_24588,N_24426,N_24348);
nand U24589 (N_24589,N_24332,N_24439);
nand U24590 (N_24590,N_24487,N_24496);
nand U24591 (N_24591,N_24271,N_24375);
and U24592 (N_24592,N_24382,N_24353);
and U24593 (N_24593,N_24385,N_24280);
nor U24594 (N_24594,N_24361,N_24261);
xnor U24595 (N_24595,N_24316,N_24305);
and U24596 (N_24596,N_24313,N_24251);
nor U24597 (N_24597,N_24351,N_24491);
nand U24598 (N_24598,N_24417,N_24458);
nor U24599 (N_24599,N_24323,N_24279);
nor U24600 (N_24600,N_24462,N_24405);
xnor U24601 (N_24601,N_24359,N_24281);
nand U24602 (N_24602,N_24324,N_24391);
nor U24603 (N_24603,N_24291,N_24483);
nor U24604 (N_24604,N_24384,N_24435);
or U24605 (N_24605,N_24292,N_24352);
nand U24606 (N_24606,N_24415,N_24360);
and U24607 (N_24607,N_24349,N_24357);
nand U24608 (N_24608,N_24478,N_24257);
nor U24609 (N_24609,N_24253,N_24452);
and U24610 (N_24610,N_24379,N_24283);
and U24611 (N_24611,N_24334,N_24398);
xnor U24612 (N_24612,N_24301,N_24325);
nor U24613 (N_24613,N_24471,N_24434);
xor U24614 (N_24614,N_24285,N_24337);
nor U24615 (N_24615,N_24411,N_24424);
nand U24616 (N_24616,N_24482,N_24402);
and U24617 (N_24617,N_24314,N_24366);
or U24618 (N_24618,N_24460,N_24423);
and U24619 (N_24619,N_24445,N_24386);
and U24620 (N_24620,N_24344,N_24408);
and U24621 (N_24621,N_24260,N_24390);
nor U24622 (N_24622,N_24378,N_24308);
nor U24623 (N_24623,N_24469,N_24377);
and U24624 (N_24624,N_24303,N_24418);
or U24625 (N_24625,N_24312,N_24376);
and U24626 (N_24626,N_24347,N_24403);
and U24627 (N_24627,N_24465,N_24379);
xnor U24628 (N_24628,N_24495,N_24375);
nor U24629 (N_24629,N_24254,N_24464);
and U24630 (N_24630,N_24384,N_24351);
nor U24631 (N_24631,N_24462,N_24365);
and U24632 (N_24632,N_24374,N_24416);
and U24633 (N_24633,N_24444,N_24488);
xnor U24634 (N_24634,N_24481,N_24468);
nor U24635 (N_24635,N_24273,N_24388);
xor U24636 (N_24636,N_24442,N_24485);
nor U24637 (N_24637,N_24432,N_24339);
and U24638 (N_24638,N_24347,N_24339);
nor U24639 (N_24639,N_24291,N_24273);
or U24640 (N_24640,N_24378,N_24417);
nand U24641 (N_24641,N_24254,N_24351);
nor U24642 (N_24642,N_24386,N_24429);
and U24643 (N_24643,N_24298,N_24463);
and U24644 (N_24644,N_24341,N_24274);
xnor U24645 (N_24645,N_24400,N_24365);
and U24646 (N_24646,N_24342,N_24257);
xor U24647 (N_24647,N_24362,N_24267);
nor U24648 (N_24648,N_24403,N_24435);
xor U24649 (N_24649,N_24428,N_24463);
nand U24650 (N_24650,N_24382,N_24402);
xor U24651 (N_24651,N_24435,N_24278);
and U24652 (N_24652,N_24258,N_24319);
nor U24653 (N_24653,N_24481,N_24381);
or U24654 (N_24654,N_24433,N_24431);
nand U24655 (N_24655,N_24435,N_24378);
nor U24656 (N_24656,N_24285,N_24473);
xor U24657 (N_24657,N_24436,N_24399);
and U24658 (N_24658,N_24316,N_24476);
and U24659 (N_24659,N_24252,N_24450);
nor U24660 (N_24660,N_24292,N_24337);
and U24661 (N_24661,N_24474,N_24261);
or U24662 (N_24662,N_24285,N_24344);
and U24663 (N_24663,N_24472,N_24331);
nor U24664 (N_24664,N_24268,N_24330);
and U24665 (N_24665,N_24428,N_24267);
nor U24666 (N_24666,N_24367,N_24327);
or U24667 (N_24667,N_24461,N_24473);
or U24668 (N_24668,N_24443,N_24271);
and U24669 (N_24669,N_24332,N_24266);
nand U24670 (N_24670,N_24305,N_24310);
and U24671 (N_24671,N_24265,N_24432);
xnor U24672 (N_24672,N_24370,N_24493);
nand U24673 (N_24673,N_24397,N_24403);
xor U24674 (N_24674,N_24272,N_24469);
xnor U24675 (N_24675,N_24335,N_24372);
or U24676 (N_24676,N_24496,N_24334);
and U24677 (N_24677,N_24322,N_24286);
xnor U24678 (N_24678,N_24354,N_24254);
nor U24679 (N_24679,N_24458,N_24436);
nand U24680 (N_24680,N_24310,N_24484);
xor U24681 (N_24681,N_24476,N_24422);
nand U24682 (N_24682,N_24266,N_24419);
xnor U24683 (N_24683,N_24434,N_24314);
and U24684 (N_24684,N_24273,N_24272);
or U24685 (N_24685,N_24265,N_24252);
xor U24686 (N_24686,N_24358,N_24366);
and U24687 (N_24687,N_24371,N_24420);
nor U24688 (N_24688,N_24308,N_24352);
xnor U24689 (N_24689,N_24369,N_24381);
and U24690 (N_24690,N_24339,N_24359);
and U24691 (N_24691,N_24298,N_24488);
nand U24692 (N_24692,N_24478,N_24450);
nand U24693 (N_24693,N_24485,N_24371);
and U24694 (N_24694,N_24446,N_24283);
or U24695 (N_24695,N_24255,N_24469);
nand U24696 (N_24696,N_24250,N_24298);
or U24697 (N_24697,N_24406,N_24370);
or U24698 (N_24698,N_24325,N_24460);
nand U24699 (N_24699,N_24360,N_24303);
or U24700 (N_24700,N_24394,N_24365);
xor U24701 (N_24701,N_24361,N_24448);
nor U24702 (N_24702,N_24384,N_24310);
xor U24703 (N_24703,N_24479,N_24383);
nand U24704 (N_24704,N_24365,N_24259);
and U24705 (N_24705,N_24359,N_24463);
nand U24706 (N_24706,N_24331,N_24272);
nor U24707 (N_24707,N_24314,N_24431);
nor U24708 (N_24708,N_24297,N_24369);
nor U24709 (N_24709,N_24314,N_24497);
nor U24710 (N_24710,N_24253,N_24398);
and U24711 (N_24711,N_24348,N_24382);
nor U24712 (N_24712,N_24266,N_24463);
nand U24713 (N_24713,N_24388,N_24494);
xor U24714 (N_24714,N_24291,N_24338);
or U24715 (N_24715,N_24333,N_24427);
xor U24716 (N_24716,N_24487,N_24271);
nor U24717 (N_24717,N_24285,N_24407);
nor U24718 (N_24718,N_24311,N_24484);
nor U24719 (N_24719,N_24259,N_24474);
nor U24720 (N_24720,N_24339,N_24454);
nand U24721 (N_24721,N_24453,N_24371);
xor U24722 (N_24722,N_24289,N_24407);
nor U24723 (N_24723,N_24485,N_24364);
nor U24724 (N_24724,N_24422,N_24371);
xor U24725 (N_24725,N_24393,N_24267);
nand U24726 (N_24726,N_24465,N_24398);
and U24727 (N_24727,N_24313,N_24270);
nor U24728 (N_24728,N_24397,N_24477);
or U24729 (N_24729,N_24351,N_24411);
nand U24730 (N_24730,N_24261,N_24420);
or U24731 (N_24731,N_24360,N_24344);
xnor U24732 (N_24732,N_24398,N_24391);
and U24733 (N_24733,N_24377,N_24429);
nor U24734 (N_24734,N_24281,N_24256);
xor U24735 (N_24735,N_24298,N_24448);
nor U24736 (N_24736,N_24498,N_24432);
and U24737 (N_24737,N_24251,N_24312);
nand U24738 (N_24738,N_24436,N_24332);
nand U24739 (N_24739,N_24268,N_24381);
nor U24740 (N_24740,N_24300,N_24408);
nand U24741 (N_24741,N_24424,N_24455);
nand U24742 (N_24742,N_24427,N_24314);
nor U24743 (N_24743,N_24305,N_24412);
nand U24744 (N_24744,N_24476,N_24392);
nand U24745 (N_24745,N_24389,N_24316);
nand U24746 (N_24746,N_24387,N_24439);
nor U24747 (N_24747,N_24280,N_24390);
nand U24748 (N_24748,N_24324,N_24298);
or U24749 (N_24749,N_24316,N_24339);
nand U24750 (N_24750,N_24569,N_24650);
nor U24751 (N_24751,N_24661,N_24584);
or U24752 (N_24752,N_24625,N_24746);
nand U24753 (N_24753,N_24713,N_24624);
nor U24754 (N_24754,N_24622,N_24575);
or U24755 (N_24755,N_24508,N_24518);
xor U24756 (N_24756,N_24691,N_24731);
xor U24757 (N_24757,N_24599,N_24593);
nand U24758 (N_24758,N_24534,N_24557);
nor U24759 (N_24759,N_24727,N_24596);
nor U24760 (N_24760,N_24503,N_24700);
or U24761 (N_24761,N_24717,N_24615);
and U24762 (N_24762,N_24737,N_24607);
and U24763 (N_24763,N_24715,N_24634);
xor U24764 (N_24764,N_24679,N_24571);
and U24765 (N_24765,N_24511,N_24649);
and U24766 (N_24766,N_24576,N_24629);
nor U24767 (N_24767,N_24683,N_24682);
xnor U24768 (N_24768,N_24574,N_24704);
or U24769 (N_24769,N_24739,N_24603);
and U24770 (N_24770,N_24560,N_24709);
nor U24771 (N_24771,N_24577,N_24586);
nor U24772 (N_24772,N_24510,N_24501);
nor U24773 (N_24773,N_24564,N_24667);
or U24774 (N_24774,N_24686,N_24705);
and U24775 (N_24775,N_24516,N_24669);
nor U24776 (N_24776,N_24609,N_24589);
or U24777 (N_24777,N_24743,N_24675);
and U24778 (N_24778,N_24707,N_24633);
xor U24779 (N_24779,N_24627,N_24726);
nor U24780 (N_24780,N_24600,N_24712);
nand U24781 (N_24781,N_24733,N_24736);
or U24782 (N_24782,N_24610,N_24690);
nor U24783 (N_24783,N_24671,N_24546);
or U24784 (N_24784,N_24708,N_24528);
and U24785 (N_24785,N_24630,N_24590);
nand U24786 (N_24786,N_24677,N_24541);
nand U24787 (N_24787,N_24660,N_24504);
or U24788 (N_24788,N_24740,N_24538);
and U24789 (N_24789,N_24532,N_24515);
xor U24790 (N_24790,N_24621,N_24573);
or U24791 (N_24791,N_24529,N_24558);
xor U24792 (N_24792,N_24565,N_24628);
nor U24793 (N_24793,N_24655,N_24555);
or U24794 (N_24794,N_24698,N_24735);
nand U24795 (N_24795,N_24587,N_24666);
nor U24796 (N_24796,N_24618,N_24559);
nand U24797 (N_24797,N_24520,N_24725);
xnor U24798 (N_24798,N_24676,N_24659);
nand U24799 (N_24799,N_24517,N_24719);
xnor U24800 (N_24800,N_24581,N_24547);
and U24801 (N_24801,N_24536,N_24722);
xnor U24802 (N_24802,N_24554,N_24572);
xor U24803 (N_24803,N_24638,N_24505);
or U24804 (N_24804,N_24601,N_24647);
or U24805 (N_24805,N_24662,N_24728);
nand U24806 (N_24806,N_24553,N_24668);
nand U24807 (N_24807,N_24670,N_24548);
xnor U24808 (N_24808,N_24651,N_24524);
nor U24809 (N_24809,N_24730,N_24641);
nor U24810 (N_24810,N_24513,N_24561);
nand U24811 (N_24811,N_24544,N_24500);
nand U24812 (N_24812,N_24531,N_24645);
nand U24813 (N_24813,N_24533,N_24642);
nand U24814 (N_24814,N_24566,N_24718);
nand U24815 (N_24815,N_24741,N_24535);
and U24816 (N_24816,N_24522,N_24540);
nand U24817 (N_24817,N_24527,N_24545);
xor U24818 (N_24818,N_24692,N_24711);
nand U24819 (N_24819,N_24543,N_24693);
and U24820 (N_24820,N_24694,N_24563);
nor U24821 (N_24821,N_24732,N_24525);
xor U24822 (N_24822,N_24594,N_24606);
nand U24823 (N_24823,N_24644,N_24588);
xor U24824 (N_24824,N_24714,N_24654);
or U24825 (N_24825,N_24724,N_24568);
xnor U24826 (N_24826,N_24506,N_24602);
xnor U24827 (N_24827,N_24604,N_24672);
nand U24828 (N_24828,N_24749,N_24597);
xor U24829 (N_24829,N_24616,N_24665);
xnor U24830 (N_24830,N_24612,N_24640);
xnor U24831 (N_24831,N_24585,N_24579);
nand U24832 (N_24832,N_24721,N_24570);
nand U24833 (N_24833,N_24514,N_24637);
and U24834 (N_24834,N_24738,N_24747);
nor U24835 (N_24835,N_24542,N_24562);
and U24836 (N_24836,N_24652,N_24552);
and U24837 (N_24837,N_24699,N_24507);
and U24838 (N_24838,N_24697,N_24688);
nand U24839 (N_24839,N_24748,N_24678);
xor U24840 (N_24840,N_24656,N_24530);
nand U24841 (N_24841,N_24556,N_24617);
or U24842 (N_24842,N_24583,N_24681);
nor U24843 (N_24843,N_24674,N_24643);
nand U24844 (N_24844,N_24580,N_24592);
or U24845 (N_24845,N_24742,N_24684);
nor U24846 (N_24846,N_24663,N_24745);
xnor U24847 (N_24847,N_24502,N_24595);
or U24848 (N_24848,N_24729,N_24526);
or U24849 (N_24849,N_24598,N_24710);
xnor U24850 (N_24850,N_24673,N_24523);
xnor U24851 (N_24851,N_24689,N_24605);
and U24852 (N_24852,N_24695,N_24664);
nand U24853 (N_24853,N_24626,N_24578);
or U24854 (N_24854,N_24608,N_24567);
nor U24855 (N_24855,N_24539,N_24720);
xnor U24856 (N_24856,N_24680,N_24653);
and U24857 (N_24857,N_24685,N_24620);
nand U24858 (N_24858,N_24723,N_24582);
nand U24859 (N_24859,N_24639,N_24744);
nand U24860 (N_24860,N_24519,N_24551);
nand U24861 (N_24861,N_24614,N_24635);
xnor U24862 (N_24862,N_24716,N_24537);
or U24863 (N_24863,N_24687,N_24702);
xnor U24864 (N_24864,N_24701,N_24512);
xor U24865 (N_24865,N_24613,N_24550);
xor U24866 (N_24866,N_24657,N_24658);
nand U24867 (N_24867,N_24696,N_24636);
nor U24868 (N_24868,N_24632,N_24648);
and U24869 (N_24869,N_24646,N_24631);
nand U24870 (N_24870,N_24509,N_24521);
nand U24871 (N_24871,N_24549,N_24623);
xor U24872 (N_24872,N_24706,N_24734);
xor U24873 (N_24873,N_24591,N_24703);
and U24874 (N_24874,N_24611,N_24619);
xnor U24875 (N_24875,N_24636,N_24545);
xor U24876 (N_24876,N_24714,N_24629);
nor U24877 (N_24877,N_24505,N_24603);
nor U24878 (N_24878,N_24584,N_24511);
xor U24879 (N_24879,N_24580,N_24546);
nand U24880 (N_24880,N_24500,N_24707);
nor U24881 (N_24881,N_24680,N_24502);
and U24882 (N_24882,N_24643,N_24657);
and U24883 (N_24883,N_24548,N_24659);
xor U24884 (N_24884,N_24618,N_24587);
xor U24885 (N_24885,N_24712,N_24576);
nor U24886 (N_24886,N_24584,N_24739);
nand U24887 (N_24887,N_24571,N_24578);
or U24888 (N_24888,N_24550,N_24523);
xor U24889 (N_24889,N_24615,N_24671);
nand U24890 (N_24890,N_24538,N_24603);
nand U24891 (N_24891,N_24592,N_24533);
nor U24892 (N_24892,N_24520,N_24698);
and U24893 (N_24893,N_24579,N_24619);
or U24894 (N_24894,N_24607,N_24571);
and U24895 (N_24895,N_24506,N_24642);
or U24896 (N_24896,N_24559,N_24534);
nor U24897 (N_24897,N_24595,N_24505);
nand U24898 (N_24898,N_24618,N_24534);
nand U24899 (N_24899,N_24523,N_24563);
nor U24900 (N_24900,N_24575,N_24574);
nor U24901 (N_24901,N_24586,N_24622);
and U24902 (N_24902,N_24601,N_24595);
xnor U24903 (N_24903,N_24598,N_24621);
and U24904 (N_24904,N_24691,N_24742);
nand U24905 (N_24905,N_24676,N_24596);
xnor U24906 (N_24906,N_24562,N_24707);
nand U24907 (N_24907,N_24584,N_24557);
nand U24908 (N_24908,N_24517,N_24710);
nand U24909 (N_24909,N_24519,N_24504);
xnor U24910 (N_24910,N_24542,N_24506);
nor U24911 (N_24911,N_24651,N_24538);
nor U24912 (N_24912,N_24592,N_24666);
or U24913 (N_24913,N_24748,N_24676);
xnor U24914 (N_24914,N_24563,N_24592);
nand U24915 (N_24915,N_24618,N_24740);
or U24916 (N_24916,N_24580,N_24560);
or U24917 (N_24917,N_24736,N_24676);
nor U24918 (N_24918,N_24654,N_24531);
and U24919 (N_24919,N_24575,N_24519);
or U24920 (N_24920,N_24710,N_24749);
nand U24921 (N_24921,N_24691,N_24530);
or U24922 (N_24922,N_24628,N_24652);
or U24923 (N_24923,N_24735,N_24742);
xor U24924 (N_24924,N_24548,N_24706);
and U24925 (N_24925,N_24684,N_24540);
nand U24926 (N_24926,N_24681,N_24508);
xor U24927 (N_24927,N_24739,N_24672);
nor U24928 (N_24928,N_24566,N_24625);
nand U24929 (N_24929,N_24564,N_24526);
xnor U24930 (N_24930,N_24544,N_24636);
nor U24931 (N_24931,N_24639,N_24501);
xnor U24932 (N_24932,N_24642,N_24680);
nor U24933 (N_24933,N_24506,N_24739);
and U24934 (N_24934,N_24676,N_24544);
or U24935 (N_24935,N_24727,N_24614);
and U24936 (N_24936,N_24565,N_24594);
nand U24937 (N_24937,N_24630,N_24691);
nor U24938 (N_24938,N_24728,N_24732);
and U24939 (N_24939,N_24526,N_24565);
and U24940 (N_24940,N_24566,N_24517);
and U24941 (N_24941,N_24521,N_24652);
nor U24942 (N_24942,N_24611,N_24629);
xor U24943 (N_24943,N_24607,N_24731);
xnor U24944 (N_24944,N_24520,N_24579);
and U24945 (N_24945,N_24510,N_24734);
or U24946 (N_24946,N_24587,N_24704);
xor U24947 (N_24947,N_24640,N_24624);
or U24948 (N_24948,N_24625,N_24691);
or U24949 (N_24949,N_24709,N_24666);
nand U24950 (N_24950,N_24566,N_24564);
and U24951 (N_24951,N_24686,N_24668);
and U24952 (N_24952,N_24563,N_24588);
nand U24953 (N_24953,N_24573,N_24544);
or U24954 (N_24954,N_24682,N_24665);
xnor U24955 (N_24955,N_24585,N_24741);
and U24956 (N_24956,N_24620,N_24547);
nor U24957 (N_24957,N_24654,N_24709);
nand U24958 (N_24958,N_24533,N_24644);
nor U24959 (N_24959,N_24693,N_24659);
or U24960 (N_24960,N_24592,N_24650);
xnor U24961 (N_24961,N_24689,N_24557);
and U24962 (N_24962,N_24651,N_24530);
nand U24963 (N_24963,N_24500,N_24656);
nand U24964 (N_24964,N_24575,N_24681);
and U24965 (N_24965,N_24604,N_24725);
nand U24966 (N_24966,N_24526,N_24530);
xnor U24967 (N_24967,N_24638,N_24566);
or U24968 (N_24968,N_24667,N_24632);
xor U24969 (N_24969,N_24541,N_24676);
or U24970 (N_24970,N_24744,N_24630);
nor U24971 (N_24971,N_24684,N_24586);
or U24972 (N_24972,N_24558,N_24564);
xnor U24973 (N_24973,N_24735,N_24503);
nor U24974 (N_24974,N_24615,N_24590);
and U24975 (N_24975,N_24653,N_24676);
nand U24976 (N_24976,N_24631,N_24648);
xor U24977 (N_24977,N_24585,N_24713);
xor U24978 (N_24978,N_24588,N_24682);
nand U24979 (N_24979,N_24726,N_24530);
and U24980 (N_24980,N_24678,N_24742);
and U24981 (N_24981,N_24690,N_24564);
and U24982 (N_24982,N_24734,N_24727);
nand U24983 (N_24983,N_24664,N_24715);
xor U24984 (N_24984,N_24657,N_24688);
xnor U24985 (N_24985,N_24719,N_24731);
or U24986 (N_24986,N_24646,N_24644);
nand U24987 (N_24987,N_24630,N_24595);
nor U24988 (N_24988,N_24711,N_24613);
or U24989 (N_24989,N_24500,N_24547);
xor U24990 (N_24990,N_24516,N_24629);
nor U24991 (N_24991,N_24570,N_24513);
and U24992 (N_24992,N_24519,N_24749);
nor U24993 (N_24993,N_24575,N_24620);
nor U24994 (N_24994,N_24690,N_24693);
or U24995 (N_24995,N_24560,N_24620);
or U24996 (N_24996,N_24652,N_24712);
or U24997 (N_24997,N_24726,N_24581);
nor U24998 (N_24998,N_24539,N_24523);
xnor U24999 (N_24999,N_24591,N_24655);
nand U25000 (N_25000,N_24970,N_24818);
and U25001 (N_25001,N_24964,N_24941);
nor U25002 (N_25002,N_24794,N_24935);
or U25003 (N_25003,N_24979,N_24785);
and U25004 (N_25004,N_24823,N_24922);
nand U25005 (N_25005,N_24909,N_24861);
and U25006 (N_25006,N_24760,N_24907);
or U25007 (N_25007,N_24837,N_24776);
or U25008 (N_25008,N_24839,N_24750);
and U25009 (N_25009,N_24865,N_24921);
or U25010 (N_25010,N_24813,N_24955);
or U25011 (N_25011,N_24761,N_24913);
nor U25012 (N_25012,N_24905,N_24984);
or U25013 (N_25013,N_24965,N_24753);
nand U25014 (N_25014,N_24953,N_24906);
nor U25015 (N_25015,N_24755,N_24876);
or U25016 (N_25016,N_24810,N_24781);
xnor U25017 (N_25017,N_24769,N_24994);
xor U25018 (N_25018,N_24793,N_24784);
nand U25019 (N_25019,N_24757,N_24936);
or U25020 (N_25020,N_24844,N_24801);
nor U25021 (N_25021,N_24947,N_24908);
nand U25022 (N_25022,N_24968,N_24973);
and U25023 (N_25023,N_24963,N_24887);
nor U25024 (N_25024,N_24828,N_24991);
or U25025 (N_25025,N_24983,N_24789);
xnor U25026 (N_25026,N_24838,N_24903);
xnor U25027 (N_25027,N_24816,N_24949);
nor U25028 (N_25028,N_24848,N_24943);
nor U25029 (N_25029,N_24795,N_24897);
and U25030 (N_25030,N_24914,N_24869);
nor U25031 (N_25031,N_24901,N_24763);
or U25032 (N_25032,N_24956,N_24788);
nor U25033 (N_25033,N_24851,N_24778);
nor U25034 (N_25034,N_24923,N_24998);
xor U25035 (N_25035,N_24927,N_24835);
or U25036 (N_25036,N_24791,N_24957);
nand U25037 (N_25037,N_24827,N_24990);
and U25038 (N_25038,N_24751,N_24768);
nor U25039 (N_25039,N_24918,N_24890);
xnor U25040 (N_25040,N_24958,N_24898);
nand U25041 (N_25041,N_24992,N_24834);
and U25042 (N_25042,N_24815,N_24933);
and U25043 (N_25043,N_24948,N_24875);
xnor U25044 (N_25044,N_24989,N_24797);
xnor U25045 (N_25045,N_24812,N_24931);
or U25046 (N_25046,N_24987,N_24764);
nand U25047 (N_25047,N_24995,N_24997);
nor U25048 (N_25048,N_24783,N_24952);
nor U25049 (N_25049,N_24855,N_24773);
nor U25050 (N_25050,N_24765,N_24819);
nor U25051 (N_25051,N_24891,N_24762);
nor U25052 (N_25052,N_24961,N_24900);
nor U25053 (N_25053,N_24808,N_24976);
or U25054 (N_25054,N_24888,N_24960);
or U25055 (N_25055,N_24841,N_24904);
nor U25056 (N_25056,N_24836,N_24988);
nand U25057 (N_25057,N_24800,N_24902);
xor U25058 (N_25058,N_24854,N_24975);
xnor U25059 (N_25059,N_24951,N_24950);
or U25060 (N_25060,N_24895,N_24849);
and U25061 (N_25061,N_24892,N_24805);
xnor U25062 (N_25062,N_24868,N_24862);
nor U25063 (N_25063,N_24972,N_24822);
and U25064 (N_25064,N_24986,N_24889);
and U25065 (N_25065,N_24938,N_24833);
nand U25066 (N_25066,N_24878,N_24982);
and U25067 (N_25067,N_24824,N_24802);
nor U25068 (N_25068,N_24792,N_24872);
nor U25069 (N_25069,N_24756,N_24917);
nor U25070 (N_25070,N_24974,N_24859);
xnor U25071 (N_25071,N_24896,N_24787);
or U25072 (N_25072,N_24911,N_24856);
or U25073 (N_25073,N_24847,N_24884);
or U25074 (N_25074,N_24937,N_24934);
xor U25075 (N_25075,N_24771,N_24831);
xnor U25076 (N_25076,N_24846,N_24967);
nor U25077 (N_25077,N_24799,N_24981);
and U25078 (N_25078,N_24843,N_24814);
xnor U25079 (N_25079,N_24877,N_24996);
and U25080 (N_25080,N_24883,N_24870);
nor U25081 (N_25081,N_24910,N_24920);
and U25082 (N_25082,N_24752,N_24821);
nand U25083 (N_25083,N_24806,N_24894);
nand U25084 (N_25084,N_24929,N_24980);
and U25085 (N_25085,N_24873,N_24852);
xor U25086 (N_25086,N_24863,N_24871);
and U25087 (N_25087,N_24754,N_24829);
xnor U25088 (N_25088,N_24932,N_24817);
and U25089 (N_25089,N_24912,N_24993);
or U25090 (N_25090,N_24779,N_24850);
nand U25091 (N_25091,N_24767,N_24966);
nor U25092 (N_25092,N_24886,N_24971);
xnor U25093 (N_25093,N_24928,N_24759);
and U25094 (N_25094,N_24962,N_24926);
and U25095 (N_25095,N_24925,N_24939);
nand U25096 (N_25096,N_24924,N_24945);
or U25097 (N_25097,N_24845,N_24782);
xnor U25098 (N_25098,N_24803,N_24766);
nor U25099 (N_25099,N_24780,N_24879);
xor U25100 (N_25100,N_24853,N_24899);
nand U25101 (N_25101,N_24880,N_24864);
nand U25102 (N_25102,N_24866,N_24774);
xor U25103 (N_25103,N_24882,N_24916);
xnor U25104 (N_25104,N_24820,N_24915);
and U25105 (N_25105,N_24867,N_24944);
and U25106 (N_25106,N_24969,N_24985);
nor U25107 (N_25107,N_24842,N_24798);
and U25108 (N_25108,N_24858,N_24840);
xnor U25109 (N_25109,N_24999,N_24860);
nor U25110 (N_25110,N_24881,N_24946);
nand U25111 (N_25111,N_24942,N_24857);
nor U25112 (N_25112,N_24811,N_24978);
xor U25113 (N_25113,N_24977,N_24809);
xnor U25114 (N_25114,N_24826,N_24954);
or U25115 (N_25115,N_24832,N_24830);
xor U25116 (N_25116,N_24874,N_24885);
or U25117 (N_25117,N_24959,N_24770);
nand U25118 (N_25118,N_24796,N_24786);
or U25119 (N_25119,N_24804,N_24930);
and U25120 (N_25120,N_24893,N_24825);
and U25121 (N_25121,N_24772,N_24807);
and U25122 (N_25122,N_24758,N_24777);
or U25123 (N_25123,N_24919,N_24790);
or U25124 (N_25124,N_24940,N_24775);
xor U25125 (N_25125,N_24769,N_24962);
and U25126 (N_25126,N_24761,N_24777);
xor U25127 (N_25127,N_24800,N_24973);
nand U25128 (N_25128,N_24793,N_24907);
or U25129 (N_25129,N_24965,N_24783);
nor U25130 (N_25130,N_24967,N_24940);
xor U25131 (N_25131,N_24780,N_24984);
xnor U25132 (N_25132,N_24992,N_24753);
or U25133 (N_25133,N_24992,N_24962);
and U25134 (N_25134,N_24865,N_24773);
xor U25135 (N_25135,N_24792,N_24958);
nor U25136 (N_25136,N_24904,N_24942);
nand U25137 (N_25137,N_24934,N_24988);
and U25138 (N_25138,N_24920,N_24761);
or U25139 (N_25139,N_24754,N_24889);
nor U25140 (N_25140,N_24771,N_24952);
or U25141 (N_25141,N_24833,N_24767);
nor U25142 (N_25142,N_24791,N_24757);
xnor U25143 (N_25143,N_24973,N_24908);
or U25144 (N_25144,N_24808,N_24892);
and U25145 (N_25145,N_24841,N_24786);
or U25146 (N_25146,N_24818,N_24762);
and U25147 (N_25147,N_24782,N_24946);
xor U25148 (N_25148,N_24774,N_24857);
or U25149 (N_25149,N_24974,N_24798);
nor U25150 (N_25150,N_24939,N_24933);
or U25151 (N_25151,N_24765,N_24822);
xor U25152 (N_25152,N_24988,N_24879);
nand U25153 (N_25153,N_24991,N_24942);
nand U25154 (N_25154,N_24906,N_24911);
or U25155 (N_25155,N_24875,N_24770);
nor U25156 (N_25156,N_24837,N_24866);
or U25157 (N_25157,N_24773,N_24878);
or U25158 (N_25158,N_24776,N_24998);
and U25159 (N_25159,N_24821,N_24796);
or U25160 (N_25160,N_24934,N_24805);
xor U25161 (N_25161,N_24759,N_24815);
xnor U25162 (N_25162,N_24767,N_24801);
and U25163 (N_25163,N_24784,N_24785);
or U25164 (N_25164,N_24931,N_24996);
nand U25165 (N_25165,N_24852,N_24847);
xnor U25166 (N_25166,N_24990,N_24899);
nor U25167 (N_25167,N_24800,N_24944);
and U25168 (N_25168,N_24926,N_24864);
or U25169 (N_25169,N_24880,N_24842);
xor U25170 (N_25170,N_24965,N_24816);
nand U25171 (N_25171,N_24943,N_24936);
nand U25172 (N_25172,N_24911,N_24886);
and U25173 (N_25173,N_24986,N_24821);
and U25174 (N_25174,N_24870,N_24925);
nand U25175 (N_25175,N_24751,N_24802);
or U25176 (N_25176,N_24826,N_24809);
and U25177 (N_25177,N_24911,N_24757);
nor U25178 (N_25178,N_24757,N_24905);
or U25179 (N_25179,N_24877,N_24780);
or U25180 (N_25180,N_24759,N_24863);
or U25181 (N_25181,N_24760,N_24838);
or U25182 (N_25182,N_24861,N_24803);
nand U25183 (N_25183,N_24765,N_24953);
and U25184 (N_25184,N_24812,N_24789);
or U25185 (N_25185,N_24950,N_24807);
or U25186 (N_25186,N_24810,N_24971);
and U25187 (N_25187,N_24755,N_24810);
xnor U25188 (N_25188,N_24916,N_24788);
nor U25189 (N_25189,N_24930,N_24921);
and U25190 (N_25190,N_24912,N_24961);
and U25191 (N_25191,N_24934,N_24770);
nand U25192 (N_25192,N_24813,N_24963);
xor U25193 (N_25193,N_24917,N_24845);
nand U25194 (N_25194,N_24878,N_24993);
xnor U25195 (N_25195,N_24770,N_24943);
nand U25196 (N_25196,N_24836,N_24835);
nand U25197 (N_25197,N_24778,N_24876);
or U25198 (N_25198,N_24969,N_24759);
nand U25199 (N_25199,N_24974,N_24831);
or U25200 (N_25200,N_24791,N_24805);
nor U25201 (N_25201,N_24825,N_24923);
xnor U25202 (N_25202,N_24980,N_24839);
nor U25203 (N_25203,N_24811,N_24767);
nor U25204 (N_25204,N_24904,N_24969);
nor U25205 (N_25205,N_24834,N_24845);
or U25206 (N_25206,N_24890,N_24855);
nand U25207 (N_25207,N_24806,N_24805);
xnor U25208 (N_25208,N_24909,N_24864);
and U25209 (N_25209,N_24775,N_24788);
nor U25210 (N_25210,N_24977,N_24956);
nor U25211 (N_25211,N_24948,N_24972);
or U25212 (N_25212,N_24947,N_24994);
and U25213 (N_25213,N_24864,N_24873);
nor U25214 (N_25214,N_24756,N_24758);
or U25215 (N_25215,N_24833,N_24963);
xnor U25216 (N_25216,N_24894,N_24825);
or U25217 (N_25217,N_24811,N_24982);
nand U25218 (N_25218,N_24967,N_24939);
nand U25219 (N_25219,N_24987,N_24772);
and U25220 (N_25220,N_24927,N_24841);
xnor U25221 (N_25221,N_24778,N_24939);
or U25222 (N_25222,N_24819,N_24864);
xnor U25223 (N_25223,N_24768,N_24774);
nor U25224 (N_25224,N_24831,N_24890);
nand U25225 (N_25225,N_24851,N_24987);
and U25226 (N_25226,N_24948,N_24757);
nand U25227 (N_25227,N_24849,N_24788);
nand U25228 (N_25228,N_24977,N_24778);
or U25229 (N_25229,N_24963,N_24869);
nand U25230 (N_25230,N_24817,N_24768);
xnor U25231 (N_25231,N_24841,N_24824);
or U25232 (N_25232,N_24966,N_24780);
or U25233 (N_25233,N_24918,N_24779);
nor U25234 (N_25234,N_24870,N_24926);
xor U25235 (N_25235,N_24947,N_24998);
and U25236 (N_25236,N_24896,N_24883);
xnor U25237 (N_25237,N_24759,N_24853);
nor U25238 (N_25238,N_24929,N_24939);
nor U25239 (N_25239,N_24853,N_24994);
or U25240 (N_25240,N_24852,N_24911);
nand U25241 (N_25241,N_24841,N_24772);
nor U25242 (N_25242,N_24982,N_24977);
and U25243 (N_25243,N_24907,N_24984);
and U25244 (N_25244,N_24897,N_24831);
nor U25245 (N_25245,N_24848,N_24959);
and U25246 (N_25246,N_24753,N_24782);
and U25247 (N_25247,N_24990,N_24786);
and U25248 (N_25248,N_24756,N_24945);
and U25249 (N_25249,N_24853,N_24928);
nor U25250 (N_25250,N_25242,N_25146);
or U25251 (N_25251,N_25214,N_25231);
and U25252 (N_25252,N_25190,N_25246);
xnor U25253 (N_25253,N_25021,N_25067);
xnor U25254 (N_25254,N_25001,N_25085);
and U25255 (N_25255,N_25159,N_25210);
xnor U25256 (N_25256,N_25203,N_25197);
and U25257 (N_25257,N_25007,N_25032);
and U25258 (N_25258,N_25241,N_25225);
nand U25259 (N_25259,N_25013,N_25048);
and U25260 (N_25260,N_25020,N_25071);
and U25261 (N_25261,N_25229,N_25059);
nor U25262 (N_25262,N_25206,N_25155);
xnor U25263 (N_25263,N_25076,N_25248);
or U25264 (N_25264,N_25158,N_25161);
nor U25265 (N_25265,N_25200,N_25141);
or U25266 (N_25266,N_25245,N_25130);
xor U25267 (N_25267,N_25050,N_25038);
nand U25268 (N_25268,N_25019,N_25029);
nand U25269 (N_25269,N_25204,N_25091);
xor U25270 (N_25270,N_25243,N_25008);
nor U25271 (N_25271,N_25072,N_25213);
nand U25272 (N_25272,N_25082,N_25142);
and U25273 (N_25273,N_25124,N_25187);
nor U25274 (N_25274,N_25057,N_25069);
and U25275 (N_25275,N_25235,N_25230);
nor U25276 (N_25276,N_25080,N_25053);
xnor U25277 (N_25277,N_25166,N_25096);
xnor U25278 (N_25278,N_25111,N_25128);
nand U25279 (N_25279,N_25120,N_25063);
or U25280 (N_25280,N_25079,N_25175);
or U25281 (N_25281,N_25193,N_25133);
or U25282 (N_25282,N_25216,N_25217);
xor U25283 (N_25283,N_25132,N_25127);
xor U25284 (N_25284,N_25129,N_25202);
and U25285 (N_25285,N_25030,N_25148);
xor U25286 (N_25286,N_25165,N_25043);
xnor U25287 (N_25287,N_25188,N_25164);
nand U25288 (N_25288,N_25102,N_25075);
or U25289 (N_25289,N_25045,N_25136);
xor U25290 (N_25290,N_25073,N_25035);
and U25291 (N_25291,N_25056,N_25211);
xor U25292 (N_25292,N_25212,N_25171);
nand U25293 (N_25293,N_25249,N_25150);
nand U25294 (N_25294,N_25002,N_25219);
and U25295 (N_25295,N_25110,N_25232);
and U25296 (N_25296,N_25153,N_25240);
xor U25297 (N_25297,N_25147,N_25228);
nand U25298 (N_25298,N_25121,N_25108);
nand U25299 (N_25299,N_25060,N_25103);
nor U25300 (N_25300,N_25037,N_25157);
or U25301 (N_25301,N_25194,N_25015);
xor U25302 (N_25302,N_25047,N_25104);
and U25303 (N_25303,N_25083,N_25006);
nand U25304 (N_25304,N_25170,N_25086);
nor U25305 (N_25305,N_25198,N_25113);
or U25306 (N_25306,N_25179,N_25138);
nor U25307 (N_25307,N_25135,N_25185);
nand U25308 (N_25308,N_25003,N_25034);
nand U25309 (N_25309,N_25101,N_25109);
nor U25310 (N_25310,N_25052,N_25156);
and U25311 (N_25311,N_25036,N_25041);
xor U25312 (N_25312,N_25100,N_25094);
or U25313 (N_25313,N_25236,N_25118);
nor U25314 (N_25314,N_25105,N_25227);
nand U25315 (N_25315,N_25220,N_25183);
xor U25316 (N_25316,N_25040,N_25062);
or U25317 (N_25317,N_25010,N_25224);
and U25318 (N_25318,N_25152,N_25107);
nor U25319 (N_25319,N_25201,N_25051);
and U25320 (N_25320,N_25122,N_25181);
or U25321 (N_25321,N_25095,N_25065);
and U25322 (N_25322,N_25221,N_25115);
xor U25323 (N_25323,N_25024,N_25064);
nand U25324 (N_25324,N_25119,N_25125);
nor U25325 (N_25325,N_25023,N_25077);
xnor U25326 (N_25326,N_25191,N_25112);
nor U25327 (N_25327,N_25247,N_25018);
xnor U25328 (N_25328,N_25144,N_25182);
and U25329 (N_25329,N_25011,N_25149);
or U25330 (N_25330,N_25234,N_25172);
xnor U25331 (N_25331,N_25233,N_25205);
nand U25332 (N_25332,N_25180,N_25087);
nor U25333 (N_25333,N_25131,N_25151);
xor U25334 (N_25334,N_25134,N_25222);
or U25335 (N_25335,N_25044,N_25028);
nor U25336 (N_25336,N_25017,N_25061);
xor U25337 (N_25337,N_25026,N_25046);
xor U25338 (N_25338,N_25081,N_25137);
nand U25339 (N_25339,N_25088,N_25049);
or U25340 (N_25340,N_25055,N_25000);
nor U25341 (N_25341,N_25022,N_25189);
and U25342 (N_25342,N_25114,N_25177);
xnor U25343 (N_25343,N_25173,N_25099);
xor U25344 (N_25344,N_25117,N_25012);
or U25345 (N_25345,N_25116,N_25218);
or U25346 (N_25346,N_25106,N_25009);
xor U25347 (N_25347,N_25042,N_25160);
nor U25348 (N_25348,N_25192,N_25014);
nand U25349 (N_25349,N_25186,N_25097);
or U25350 (N_25350,N_25162,N_25168);
or U25351 (N_25351,N_25176,N_25199);
or U25352 (N_25352,N_25215,N_25143);
nor U25353 (N_25353,N_25004,N_25207);
nand U25354 (N_25354,N_25163,N_25223);
nor U25355 (N_25355,N_25174,N_25237);
xor U25356 (N_25356,N_25178,N_25184);
nand U25357 (N_25357,N_25005,N_25239);
or U25358 (N_25358,N_25169,N_25016);
or U25359 (N_25359,N_25238,N_25070);
and U25360 (N_25360,N_25068,N_25031);
or U25361 (N_25361,N_25084,N_25033);
and U25362 (N_25362,N_25123,N_25090);
or U25363 (N_25363,N_25139,N_25208);
and U25364 (N_25364,N_25078,N_25093);
nand U25365 (N_25365,N_25226,N_25092);
nor U25366 (N_25366,N_25195,N_25209);
nand U25367 (N_25367,N_25126,N_25167);
nand U25368 (N_25368,N_25058,N_25098);
nor U25369 (N_25369,N_25054,N_25039);
nor U25370 (N_25370,N_25025,N_25066);
nand U25371 (N_25371,N_25089,N_25027);
and U25372 (N_25372,N_25244,N_25154);
or U25373 (N_25373,N_25074,N_25145);
or U25374 (N_25374,N_25140,N_25196);
nand U25375 (N_25375,N_25164,N_25122);
and U25376 (N_25376,N_25019,N_25008);
xor U25377 (N_25377,N_25158,N_25136);
nor U25378 (N_25378,N_25003,N_25234);
or U25379 (N_25379,N_25148,N_25073);
nand U25380 (N_25380,N_25159,N_25226);
nand U25381 (N_25381,N_25140,N_25032);
xor U25382 (N_25382,N_25229,N_25188);
nand U25383 (N_25383,N_25138,N_25170);
nor U25384 (N_25384,N_25082,N_25061);
and U25385 (N_25385,N_25165,N_25092);
nor U25386 (N_25386,N_25098,N_25038);
nand U25387 (N_25387,N_25101,N_25087);
or U25388 (N_25388,N_25083,N_25136);
nor U25389 (N_25389,N_25095,N_25164);
xnor U25390 (N_25390,N_25113,N_25117);
nor U25391 (N_25391,N_25174,N_25090);
nand U25392 (N_25392,N_25223,N_25114);
nor U25393 (N_25393,N_25055,N_25128);
nor U25394 (N_25394,N_25156,N_25048);
and U25395 (N_25395,N_25087,N_25107);
and U25396 (N_25396,N_25214,N_25216);
or U25397 (N_25397,N_25022,N_25049);
nand U25398 (N_25398,N_25025,N_25101);
and U25399 (N_25399,N_25048,N_25114);
xor U25400 (N_25400,N_25167,N_25151);
or U25401 (N_25401,N_25094,N_25214);
nor U25402 (N_25402,N_25134,N_25128);
xor U25403 (N_25403,N_25099,N_25032);
or U25404 (N_25404,N_25174,N_25100);
and U25405 (N_25405,N_25180,N_25154);
xor U25406 (N_25406,N_25188,N_25011);
nand U25407 (N_25407,N_25029,N_25240);
or U25408 (N_25408,N_25069,N_25174);
or U25409 (N_25409,N_25178,N_25112);
or U25410 (N_25410,N_25077,N_25231);
and U25411 (N_25411,N_25065,N_25076);
and U25412 (N_25412,N_25223,N_25237);
nor U25413 (N_25413,N_25017,N_25122);
nand U25414 (N_25414,N_25097,N_25239);
or U25415 (N_25415,N_25100,N_25014);
or U25416 (N_25416,N_25153,N_25055);
and U25417 (N_25417,N_25182,N_25071);
and U25418 (N_25418,N_25021,N_25194);
or U25419 (N_25419,N_25004,N_25218);
xor U25420 (N_25420,N_25209,N_25219);
nand U25421 (N_25421,N_25024,N_25145);
nor U25422 (N_25422,N_25241,N_25093);
xnor U25423 (N_25423,N_25015,N_25232);
nand U25424 (N_25424,N_25104,N_25221);
xor U25425 (N_25425,N_25180,N_25016);
nand U25426 (N_25426,N_25135,N_25174);
or U25427 (N_25427,N_25069,N_25098);
nor U25428 (N_25428,N_25128,N_25196);
nand U25429 (N_25429,N_25028,N_25199);
nand U25430 (N_25430,N_25078,N_25233);
or U25431 (N_25431,N_25206,N_25102);
or U25432 (N_25432,N_25218,N_25042);
nand U25433 (N_25433,N_25232,N_25133);
or U25434 (N_25434,N_25030,N_25037);
nor U25435 (N_25435,N_25245,N_25022);
xnor U25436 (N_25436,N_25118,N_25171);
xor U25437 (N_25437,N_25062,N_25013);
nor U25438 (N_25438,N_25244,N_25109);
xor U25439 (N_25439,N_25159,N_25069);
nand U25440 (N_25440,N_25130,N_25186);
or U25441 (N_25441,N_25071,N_25120);
nor U25442 (N_25442,N_25045,N_25200);
nor U25443 (N_25443,N_25071,N_25010);
nor U25444 (N_25444,N_25069,N_25108);
nor U25445 (N_25445,N_25158,N_25064);
xnor U25446 (N_25446,N_25044,N_25067);
or U25447 (N_25447,N_25183,N_25240);
nand U25448 (N_25448,N_25038,N_25056);
xnor U25449 (N_25449,N_25145,N_25131);
xnor U25450 (N_25450,N_25212,N_25221);
xor U25451 (N_25451,N_25079,N_25129);
or U25452 (N_25452,N_25218,N_25214);
nor U25453 (N_25453,N_25027,N_25203);
xnor U25454 (N_25454,N_25122,N_25087);
nand U25455 (N_25455,N_25008,N_25038);
and U25456 (N_25456,N_25113,N_25022);
or U25457 (N_25457,N_25207,N_25213);
nand U25458 (N_25458,N_25129,N_25112);
and U25459 (N_25459,N_25111,N_25223);
xnor U25460 (N_25460,N_25046,N_25183);
or U25461 (N_25461,N_25101,N_25094);
xnor U25462 (N_25462,N_25115,N_25025);
xor U25463 (N_25463,N_25143,N_25079);
nand U25464 (N_25464,N_25176,N_25008);
and U25465 (N_25465,N_25116,N_25029);
nor U25466 (N_25466,N_25154,N_25050);
xnor U25467 (N_25467,N_25023,N_25159);
nor U25468 (N_25468,N_25005,N_25211);
or U25469 (N_25469,N_25082,N_25116);
nand U25470 (N_25470,N_25057,N_25090);
or U25471 (N_25471,N_25228,N_25175);
or U25472 (N_25472,N_25186,N_25129);
and U25473 (N_25473,N_25182,N_25243);
xor U25474 (N_25474,N_25041,N_25127);
and U25475 (N_25475,N_25060,N_25223);
nor U25476 (N_25476,N_25029,N_25054);
nand U25477 (N_25477,N_25243,N_25133);
nor U25478 (N_25478,N_25030,N_25112);
nor U25479 (N_25479,N_25143,N_25149);
nor U25480 (N_25480,N_25227,N_25213);
or U25481 (N_25481,N_25056,N_25104);
or U25482 (N_25482,N_25006,N_25203);
or U25483 (N_25483,N_25056,N_25231);
or U25484 (N_25484,N_25210,N_25230);
and U25485 (N_25485,N_25189,N_25234);
or U25486 (N_25486,N_25008,N_25076);
or U25487 (N_25487,N_25194,N_25216);
or U25488 (N_25488,N_25213,N_25218);
or U25489 (N_25489,N_25066,N_25161);
and U25490 (N_25490,N_25021,N_25125);
nand U25491 (N_25491,N_25105,N_25221);
and U25492 (N_25492,N_25063,N_25138);
and U25493 (N_25493,N_25065,N_25167);
or U25494 (N_25494,N_25222,N_25057);
or U25495 (N_25495,N_25158,N_25017);
or U25496 (N_25496,N_25091,N_25047);
and U25497 (N_25497,N_25017,N_25115);
nand U25498 (N_25498,N_25093,N_25198);
xor U25499 (N_25499,N_25025,N_25207);
nand U25500 (N_25500,N_25475,N_25446);
nor U25501 (N_25501,N_25495,N_25402);
xor U25502 (N_25502,N_25297,N_25442);
and U25503 (N_25503,N_25307,N_25400);
xor U25504 (N_25504,N_25372,N_25310);
nor U25505 (N_25505,N_25412,N_25330);
or U25506 (N_25506,N_25251,N_25258);
nand U25507 (N_25507,N_25303,N_25261);
or U25508 (N_25508,N_25295,N_25314);
nor U25509 (N_25509,N_25476,N_25282);
and U25510 (N_25510,N_25368,N_25255);
nor U25511 (N_25511,N_25459,N_25425);
xnor U25512 (N_25512,N_25386,N_25396);
or U25513 (N_25513,N_25418,N_25379);
and U25514 (N_25514,N_25270,N_25283);
nand U25515 (N_25515,N_25322,N_25268);
and U25516 (N_25516,N_25433,N_25408);
nand U25517 (N_25517,N_25486,N_25325);
nand U25518 (N_25518,N_25407,N_25491);
nor U25519 (N_25519,N_25394,N_25416);
nor U25520 (N_25520,N_25273,N_25329);
nand U25521 (N_25521,N_25356,N_25403);
xnor U25522 (N_25522,N_25361,N_25305);
nor U25523 (N_25523,N_25263,N_25485);
nand U25524 (N_25524,N_25431,N_25462);
nand U25525 (N_25525,N_25346,N_25358);
xor U25526 (N_25526,N_25466,N_25465);
nor U25527 (N_25527,N_25373,N_25450);
nand U25528 (N_25528,N_25279,N_25284);
and U25529 (N_25529,N_25463,N_25404);
or U25530 (N_25530,N_25470,N_25254);
nor U25531 (N_25531,N_25440,N_25441);
xor U25532 (N_25532,N_25331,N_25429);
xnor U25533 (N_25533,N_25388,N_25472);
or U25534 (N_25534,N_25357,N_25336);
or U25535 (N_25535,N_25377,N_25341);
nor U25536 (N_25536,N_25308,N_25264);
nor U25537 (N_25537,N_25409,N_25274);
xnor U25538 (N_25538,N_25318,N_25490);
or U25539 (N_25539,N_25474,N_25387);
nor U25540 (N_25540,N_25483,N_25411);
xor U25541 (N_25541,N_25252,N_25464);
nand U25542 (N_25542,N_25487,N_25398);
nor U25543 (N_25543,N_25309,N_25278);
nor U25544 (N_25544,N_25275,N_25458);
and U25545 (N_25545,N_25337,N_25413);
and U25546 (N_25546,N_25276,N_25311);
nand U25547 (N_25547,N_25468,N_25299);
and U25548 (N_25548,N_25363,N_25488);
and U25549 (N_25549,N_25383,N_25324);
or U25550 (N_25550,N_25456,N_25347);
xnor U25551 (N_25551,N_25477,N_25420);
nand U25552 (N_25552,N_25259,N_25328);
or U25553 (N_25553,N_25371,N_25417);
nand U25554 (N_25554,N_25312,N_25489);
and U25555 (N_25555,N_25344,N_25339);
and U25556 (N_25556,N_25269,N_25382);
nor U25557 (N_25557,N_25348,N_25423);
or U25558 (N_25558,N_25447,N_25340);
and U25559 (N_25559,N_25424,N_25378);
xor U25560 (N_25560,N_25391,N_25497);
nand U25561 (N_25561,N_25281,N_25267);
and U25562 (N_25562,N_25345,N_25498);
or U25563 (N_25563,N_25479,N_25380);
xor U25564 (N_25564,N_25395,N_25410);
and U25565 (N_25565,N_25426,N_25460);
nor U25566 (N_25566,N_25453,N_25292);
nor U25567 (N_25567,N_25353,N_25384);
or U25568 (N_25568,N_25438,N_25291);
or U25569 (N_25569,N_25494,N_25250);
xnor U25570 (N_25570,N_25427,N_25392);
or U25571 (N_25571,N_25422,N_25484);
and U25572 (N_25572,N_25385,N_25351);
nand U25573 (N_25573,N_25436,N_25370);
nand U25574 (N_25574,N_25350,N_25493);
xnor U25575 (N_25575,N_25323,N_25482);
and U25576 (N_25576,N_25319,N_25301);
xnor U25577 (N_25577,N_25359,N_25272);
xnor U25578 (N_25578,N_25454,N_25300);
nor U25579 (N_25579,N_25471,N_25320);
xnor U25580 (N_25580,N_25256,N_25428);
and U25581 (N_25581,N_25302,N_25381);
xnor U25582 (N_25582,N_25327,N_25257);
nand U25583 (N_25583,N_25445,N_25432);
xnor U25584 (N_25584,N_25289,N_25451);
nand U25585 (N_25585,N_25316,N_25306);
xnor U25586 (N_25586,N_25389,N_25304);
or U25587 (N_25587,N_25375,N_25362);
or U25588 (N_25588,N_25321,N_25260);
and U25589 (N_25589,N_25430,N_25277);
nand U25590 (N_25590,N_25461,N_25286);
or U25591 (N_25591,N_25435,N_25390);
and U25592 (N_25592,N_25467,N_25285);
or U25593 (N_25593,N_25326,N_25335);
nor U25594 (N_25594,N_25365,N_25448);
nor U25595 (N_25595,N_25354,N_25294);
xor U25596 (N_25596,N_25290,N_25452);
nand U25597 (N_25597,N_25415,N_25393);
nor U25598 (N_25598,N_25366,N_25332);
or U25599 (N_25599,N_25280,N_25457);
xnor U25600 (N_25600,N_25499,N_25313);
or U25601 (N_25601,N_25360,N_25414);
nand U25602 (N_25602,N_25315,N_25317);
and U25603 (N_25603,N_25293,N_25342);
and U25604 (N_25604,N_25338,N_25405);
and U25605 (N_25605,N_25298,N_25455);
and U25606 (N_25606,N_25364,N_25406);
nor U25607 (N_25607,N_25481,N_25469);
nand U25608 (N_25608,N_25492,N_25271);
nand U25609 (N_25609,N_25421,N_25296);
nor U25610 (N_25610,N_25266,N_25253);
nor U25611 (N_25611,N_25355,N_25262);
and U25612 (N_25612,N_25434,N_25288);
or U25613 (N_25613,N_25349,N_25343);
or U25614 (N_25614,N_25478,N_25437);
nand U25615 (N_25615,N_25374,N_25333);
and U25616 (N_25616,N_25399,N_25439);
and U25617 (N_25617,N_25376,N_25352);
nand U25618 (N_25618,N_25419,N_25444);
nor U25619 (N_25619,N_25369,N_25367);
and U25620 (N_25620,N_25480,N_25473);
or U25621 (N_25621,N_25334,N_25401);
and U25622 (N_25622,N_25443,N_25265);
xor U25623 (N_25623,N_25496,N_25449);
nand U25624 (N_25624,N_25287,N_25397);
nand U25625 (N_25625,N_25369,N_25274);
or U25626 (N_25626,N_25431,N_25281);
or U25627 (N_25627,N_25412,N_25474);
nor U25628 (N_25628,N_25417,N_25294);
nor U25629 (N_25629,N_25360,N_25373);
nor U25630 (N_25630,N_25393,N_25383);
or U25631 (N_25631,N_25415,N_25269);
nor U25632 (N_25632,N_25381,N_25477);
nor U25633 (N_25633,N_25266,N_25389);
nand U25634 (N_25634,N_25281,N_25454);
and U25635 (N_25635,N_25466,N_25339);
nand U25636 (N_25636,N_25387,N_25426);
or U25637 (N_25637,N_25255,N_25423);
or U25638 (N_25638,N_25328,N_25343);
nand U25639 (N_25639,N_25393,N_25307);
nand U25640 (N_25640,N_25259,N_25429);
or U25641 (N_25641,N_25375,N_25409);
nor U25642 (N_25642,N_25420,N_25375);
and U25643 (N_25643,N_25405,N_25310);
nand U25644 (N_25644,N_25338,N_25382);
xnor U25645 (N_25645,N_25394,N_25303);
xnor U25646 (N_25646,N_25461,N_25329);
or U25647 (N_25647,N_25358,N_25427);
nor U25648 (N_25648,N_25352,N_25414);
nor U25649 (N_25649,N_25483,N_25415);
or U25650 (N_25650,N_25472,N_25491);
or U25651 (N_25651,N_25378,N_25472);
and U25652 (N_25652,N_25432,N_25277);
nor U25653 (N_25653,N_25324,N_25417);
xor U25654 (N_25654,N_25435,N_25450);
or U25655 (N_25655,N_25295,N_25307);
xor U25656 (N_25656,N_25417,N_25471);
and U25657 (N_25657,N_25260,N_25416);
xnor U25658 (N_25658,N_25495,N_25356);
nor U25659 (N_25659,N_25462,N_25284);
or U25660 (N_25660,N_25465,N_25350);
nor U25661 (N_25661,N_25275,N_25353);
nand U25662 (N_25662,N_25361,N_25358);
nor U25663 (N_25663,N_25389,N_25467);
nand U25664 (N_25664,N_25442,N_25281);
nor U25665 (N_25665,N_25421,N_25291);
xnor U25666 (N_25666,N_25331,N_25435);
or U25667 (N_25667,N_25453,N_25278);
nand U25668 (N_25668,N_25299,N_25375);
nor U25669 (N_25669,N_25399,N_25278);
xor U25670 (N_25670,N_25354,N_25299);
xnor U25671 (N_25671,N_25496,N_25413);
nand U25672 (N_25672,N_25459,N_25444);
or U25673 (N_25673,N_25492,N_25497);
and U25674 (N_25674,N_25493,N_25473);
xnor U25675 (N_25675,N_25361,N_25299);
nor U25676 (N_25676,N_25388,N_25377);
nor U25677 (N_25677,N_25463,N_25356);
nand U25678 (N_25678,N_25340,N_25364);
or U25679 (N_25679,N_25390,N_25496);
or U25680 (N_25680,N_25312,N_25385);
nand U25681 (N_25681,N_25398,N_25367);
and U25682 (N_25682,N_25485,N_25298);
xnor U25683 (N_25683,N_25272,N_25279);
and U25684 (N_25684,N_25314,N_25381);
and U25685 (N_25685,N_25470,N_25431);
nor U25686 (N_25686,N_25493,N_25381);
xnor U25687 (N_25687,N_25275,N_25428);
or U25688 (N_25688,N_25453,N_25341);
and U25689 (N_25689,N_25406,N_25361);
or U25690 (N_25690,N_25269,N_25385);
nand U25691 (N_25691,N_25328,N_25383);
nand U25692 (N_25692,N_25442,N_25319);
xnor U25693 (N_25693,N_25338,N_25330);
nand U25694 (N_25694,N_25449,N_25326);
xor U25695 (N_25695,N_25400,N_25488);
or U25696 (N_25696,N_25421,N_25344);
nor U25697 (N_25697,N_25375,N_25380);
and U25698 (N_25698,N_25393,N_25378);
and U25699 (N_25699,N_25495,N_25264);
nor U25700 (N_25700,N_25401,N_25490);
nand U25701 (N_25701,N_25397,N_25418);
and U25702 (N_25702,N_25346,N_25403);
xor U25703 (N_25703,N_25396,N_25493);
nand U25704 (N_25704,N_25265,N_25426);
nand U25705 (N_25705,N_25282,N_25396);
nor U25706 (N_25706,N_25408,N_25266);
xnor U25707 (N_25707,N_25430,N_25491);
nand U25708 (N_25708,N_25258,N_25313);
or U25709 (N_25709,N_25468,N_25359);
or U25710 (N_25710,N_25448,N_25441);
xnor U25711 (N_25711,N_25333,N_25419);
and U25712 (N_25712,N_25434,N_25486);
xnor U25713 (N_25713,N_25341,N_25270);
xnor U25714 (N_25714,N_25461,N_25300);
and U25715 (N_25715,N_25371,N_25483);
or U25716 (N_25716,N_25433,N_25282);
and U25717 (N_25717,N_25394,N_25364);
xnor U25718 (N_25718,N_25388,N_25286);
xnor U25719 (N_25719,N_25286,N_25483);
xnor U25720 (N_25720,N_25380,N_25372);
xnor U25721 (N_25721,N_25318,N_25474);
xnor U25722 (N_25722,N_25370,N_25472);
and U25723 (N_25723,N_25499,N_25333);
xor U25724 (N_25724,N_25324,N_25398);
nor U25725 (N_25725,N_25478,N_25341);
or U25726 (N_25726,N_25357,N_25344);
xor U25727 (N_25727,N_25428,N_25271);
xor U25728 (N_25728,N_25342,N_25319);
and U25729 (N_25729,N_25385,N_25401);
nor U25730 (N_25730,N_25341,N_25431);
or U25731 (N_25731,N_25404,N_25420);
nand U25732 (N_25732,N_25481,N_25420);
and U25733 (N_25733,N_25295,N_25434);
nand U25734 (N_25734,N_25303,N_25430);
nor U25735 (N_25735,N_25486,N_25373);
xnor U25736 (N_25736,N_25319,N_25484);
and U25737 (N_25737,N_25488,N_25466);
nor U25738 (N_25738,N_25481,N_25376);
nand U25739 (N_25739,N_25255,N_25339);
or U25740 (N_25740,N_25361,N_25382);
and U25741 (N_25741,N_25492,N_25454);
or U25742 (N_25742,N_25402,N_25261);
nor U25743 (N_25743,N_25332,N_25458);
nor U25744 (N_25744,N_25451,N_25290);
or U25745 (N_25745,N_25334,N_25473);
nand U25746 (N_25746,N_25445,N_25276);
and U25747 (N_25747,N_25406,N_25268);
or U25748 (N_25748,N_25451,N_25416);
nor U25749 (N_25749,N_25334,N_25278);
nand U25750 (N_25750,N_25505,N_25537);
and U25751 (N_25751,N_25529,N_25541);
xnor U25752 (N_25752,N_25508,N_25694);
or U25753 (N_25753,N_25695,N_25673);
nor U25754 (N_25754,N_25503,N_25641);
nor U25755 (N_25755,N_25717,N_25548);
xor U25756 (N_25756,N_25604,N_25701);
nand U25757 (N_25757,N_25561,N_25709);
or U25758 (N_25758,N_25611,N_25521);
nand U25759 (N_25759,N_25674,N_25570);
and U25760 (N_25760,N_25699,N_25589);
nor U25761 (N_25761,N_25680,N_25605);
xor U25762 (N_25762,N_25707,N_25724);
and U25763 (N_25763,N_25645,N_25740);
or U25764 (N_25764,N_25524,N_25650);
and U25765 (N_25765,N_25635,N_25655);
nand U25766 (N_25766,N_25644,N_25585);
or U25767 (N_25767,N_25735,N_25553);
nand U25768 (N_25768,N_25716,N_25666);
nand U25769 (N_25769,N_25579,N_25690);
nand U25770 (N_25770,N_25612,N_25582);
nor U25771 (N_25771,N_25702,N_25522);
or U25772 (N_25772,N_25517,N_25533);
nor U25773 (N_25773,N_25504,N_25621);
xor U25774 (N_25774,N_25500,N_25606);
nor U25775 (N_25775,N_25581,N_25693);
xor U25776 (N_25776,N_25659,N_25719);
xor U25777 (N_25777,N_25728,N_25652);
nand U25778 (N_25778,N_25691,N_25737);
nand U25779 (N_25779,N_25603,N_25557);
and U25780 (N_25780,N_25647,N_25668);
xnor U25781 (N_25781,N_25577,N_25704);
xor U25782 (N_25782,N_25554,N_25639);
or U25783 (N_25783,N_25664,N_25506);
nor U25784 (N_25784,N_25660,N_25653);
nor U25785 (N_25785,N_25591,N_25683);
nand U25786 (N_25786,N_25566,N_25525);
or U25787 (N_25787,N_25528,N_25592);
and U25788 (N_25788,N_25721,N_25527);
nor U25789 (N_25789,N_25720,N_25625);
xnor U25790 (N_25790,N_25600,N_25501);
or U25791 (N_25791,N_25595,N_25609);
or U25792 (N_25792,N_25675,N_25531);
xnor U25793 (N_25793,N_25552,N_25538);
and U25794 (N_25794,N_25615,N_25572);
nand U25795 (N_25795,N_25733,N_25697);
nor U25796 (N_25796,N_25738,N_25640);
nand U25797 (N_25797,N_25692,N_25616);
or U25798 (N_25798,N_25520,N_25620);
nand U25799 (N_25799,N_25715,N_25516);
and U25800 (N_25800,N_25739,N_25565);
xor U25801 (N_25801,N_25560,N_25703);
xnor U25802 (N_25802,N_25624,N_25725);
and U25803 (N_25803,N_25722,N_25672);
or U25804 (N_25804,N_25613,N_25599);
and U25805 (N_25805,N_25656,N_25632);
and U25806 (N_25806,N_25670,N_25558);
nor U25807 (N_25807,N_25545,N_25597);
nor U25808 (N_25808,N_25593,N_25628);
or U25809 (N_25809,N_25530,N_25634);
or U25810 (N_25810,N_25731,N_25630);
and U25811 (N_25811,N_25534,N_25661);
or U25812 (N_25812,N_25590,N_25736);
nand U25813 (N_25813,N_25682,N_25550);
nand U25814 (N_25814,N_25578,N_25532);
nand U25815 (N_25815,N_25514,N_25663);
xnor U25816 (N_25816,N_25676,N_25688);
xnor U25817 (N_25817,N_25681,N_25567);
and U25818 (N_25818,N_25633,N_25610);
xor U25819 (N_25819,N_25562,N_25619);
and U25820 (N_25820,N_25658,N_25511);
and U25821 (N_25821,N_25583,N_25741);
nand U25822 (N_25822,N_25622,N_25623);
or U25823 (N_25823,N_25555,N_25689);
nand U25824 (N_25824,N_25539,N_25526);
and U25825 (N_25825,N_25564,N_25596);
xnor U25826 (N_25826,N_25549,N_25677);
nor U25827 (N_25827,N_25636,N_25732);
and U25828 (N_25828,N_25546,N_25536);
or U25829 (N_25829,N_25711,N_25726);
or U25830 (N_25830,N_25598,N_25512);
xor U25831 (N_25831,N_25573,N_25643);
nand U25832 (N_25832,N_25638,N_25618);
and U25833 (N_25833,N_25543,N_25629);
nand U25834 (N_25834,N_25513,N_25678);
nor U25835 (N_25835,N_25669,N_25617);
and U25836 (N_25836,N_25747,N_25712);
or U25837 (N_25837,N_25729,N_25580);
nand U25838 (N_25838,N_25746,N_25742);
or U25839 (N_25839,N_25667,N_25687);
or U25840 (N_25840,N_25713,N_25705);
xor U25841 (N_25841,N_25587,N_25714);
and U25842 (N_25842,N_25535,N_25540);
nand U25843 (N_25843,N_25651,N_25519);
and U25844 (N_25844,N_25745,N_25556);
and U25845 (N_25845,N_25684,N_25730);
nand U25846 (N_25846,N_25542,N_25734);
and U25847 (N_25847,N_25696,N_25627);
xor U25848 (N_25848,N_25509,N_25642);
or U25849 (N_25849,N_25649,N_25748);
nand U25850 (N_25850,N_25601,N_25665);
or U25851 (N_25851,N_25662,N_25727);
and U25852 (N_25852,N_25700,N_25698);
and U25853 (N_25853,N_25551,N_25631);
nor U25854 (N_25854,N_25547,N_25614);
or U25855 (N_25855,N_25584,N_25654);
or U25856 (N_25856,N_25607,N_25657);
nor U25857 (N_25857,N_25744,N_25706);
and U25858 (N_25858,N_25594,N_25749);
nor U25859 (N_25859,N_25626,N_25569);
xor U25860 (N_25860,N_25571,N_25568);
or U25861 (N_25861,N_25576,N_25718);
and U25862 (N_25862,N_25708,N_25671);
nor U25863 (N_25863,N_25586,N_25646);
or U25864 (N_25864,N_25563,N_25575);
nand U25865 (N_25865,N_25523,N_25723);
nor U25866 (N_25866,N_25588,N_25574);
xor U25867 (N_25867,N_25559,N_25502);
nor U25868 (N_25868,N_25602,N_25648);
or U25869 (N_25869,N_25679,N_25518);
or U25870 (N_25870,N_25686,N_25710);
xnor U25871 (N_25871,N_25507,N_25510);
or U25872 (N_25872,N_25544,N_25685);
xnor U25873 (N_25873,N_25637,N_25743);
or U25874 (N_25874,N_25515,N_25608);
or U25875 (N_25875,N_25526,N_25715);
or U25876 (N_25876,N_25744,N_25631);
nor U25877 (N_25877,N_25686,N_25677);
and U25878 (N_25878,N_25718,N_25742);
or U25879 (N_25879,N_25683,N_25749);
nand U25880 (N_25880,N_25610,N_25584);
nand U25881 (N_25881,N_25506,N_25719);
and U25882 (N_25882,N_25590,N_25698);
xnor U25883 (N_25883,N_25659,N_25514);
xnor U25884 (N_25884,N_25546,N_25738);
nand U25885 (N_25885,N_25547,N_25656);
and U25886 (N_25886,N_25546,N_25717);
nor U25887 (N_25887,N_25668,N_25571);
nand U25888 (N_25888,N_25718,N_25674);
nand U25889 (N_25889,N_25702,N_25747);
or U25890 (N_25890,N_25546,N_25662);
xor U25891 (N_25891,N_25615,N_25728);
nand U25892 (N_25892,N_25569,N_25708);
nor U25893 (N_25893,N_25704,N_25681);
xor U25894 (N_25894,N_25732,N_25554);
xnor U25895 (N_25895,N_25550,N_25647);
and U25896 (N_25896,N_25629,N_25514);
nand U25897 (N_25897,N_25506,N_25689);
nand U25898 (N_25898,N_25657,N_25595);
nor U25899 (N_25899,N_25665,N_25538);
and U25900 (N_25900,N_25571,N_25700);
nor U25901 (N_25901,N_25595,N_25729);
and U25902 (N_25902,N_25573,N_25610);
and U25903 (N_25903,N_25559,N_25670);
nor U25904 (N_25904,N_25727,N_25733);
nand U25905 (N_25905,N_25595,N_25724);
nor U25906 (N_25906,N_25520,N_25661);
nand U25907 (N_25907,N_25730,N_25559);
or U25908 (N_25908,N_25708,N_25523);
nor U25909 (N_25909,N_25685,N_25648);
nor U25910 (N_25910,N_25734,N_25544);
and U25911 (N_25911,N_25524,N_25516);
nor U25912 (N_25912,N_25684,N_25548);
nand U25913 (N_25913,N_25542,N_25602);
and U25914 (N_25914,N_25730,N_25617);
or U25915 (N_25915,N_25664,N_25605);
and U25916 (N_25916,N_25597,N_25746);
xor U25917 (N_25917,N_25685,N_25747);
and U25918 (N_25918,N_25532,N_25527);
and U25919 (N_25919,N_25628,N_25696);
or U25920 (N_25920,N_25643,N_25569);
or U25921 (N_25921,N_25653,N_25608);
or U25922 (N_25922,N_25533,N_25572);
and U25923 (N_25923,N_25718,N_25685);
and U25924 (N_25924,N_25644,N_25676);
and U25925 (N_25925,N_25684,N_25572);
nand U25926 (N_25926,N_25630,N_25553);
or U25927 (N_25927,N_25632,N_25648);
nor U25928 (N_25928,N_25743,N_25739);
or U25929 (N_25929,N_25692,N_25519);
xor U25930 (N_25930,N_25718,N_25729);
nor U25931 (N_25931,N_25536,N_25621);
and U25932 (N_25932,N_25506,N_25726);
or U25933 (N_25933,N_25501,N_25555);
and U25934 (N_25934,N_25648,N_25574);
or U25935 (N_25935,N_25686,N_25518);
or U25936 (N_25936,N_25587,N_25569);
xnor U25937 (N_25937,N_25708,N_25652);
nor U25938 (N_25938,N_25739,N_25569);
nand U25939 (N_25939,N_25565,N_25547);
or U25940 (N_25940,N_25726,N_25649);
or U25941 (N_25941,N_25608,N_25607);
nor U25942 (N_25942,N_25524,N_25534);
xnor U25943 (N_25943,N_25504,N_25736);
nor U25944 (N_25944,N_25520,N_25729);
nand U25945 (N_25945,N_25527,N_25645);
and U25946 (N_25946,N_25640,N_25728);
nand U25947 (N_25947,N_25507,N_25733);
xor U25948 (N_25948,N_25502,N_25654);
nor U25949 (N_25949,N_25600,N_25569);
nor U25950 (N_25950,N_25629,N_25721);
or U25951 (N_25951,N_25724,N_25682);
and U25952 (N_25952,N_25548,N_25685);
nand U25953 (N_25953,N_25724,N_25744);
nor U25954 (N_25954,N_25595,N_25649);
nand U25955 (N_25955,N_25713,N_25638);
nor U25956 (N_25956,N_25681,N_25719);
nor U25957 (N_25957,N_25683,N_25723);
nand U25958 (N_25958,N_25710,N_25547);
or U25959 (N_25959,N_25569,N_25623);
xor U25960 (N_25960,N_25601,N_25700);
and U25961 (N_25961,N_25632,N_25691);
or U25962 (N_25962,N_25646,N_25685);
or U25963 (N_25963,N_25597,N_25670);
nor U25964 (N_25964,N_25669,N_25641);
xnor U25965 (N_25965,N_25617,N_25539);
nand U25966 (N_25966,N_25749,N_25613);
xor U25967 (N_25967,N_25518,N_25517);
or U25968 (N_25968,N_25568,N_25548);
and U25969 (N_25969,N_25512,N_25631);
and U25970 (N_25970,N_25545,N_25538);
or U25971 (N_25971,N_25629,N_25679);
nand U25972 (N_25972,N_25696,N_25618);
xnor U25973 (N_25973,N_25565,N_25629);
nor U25974 (N_25974,N_25549,N_25723);
nor U25975 (N_25975,N_25659,N_25600);
nor U25976 (N_25976,N_25603,N_25713);
nand U25977 (N_25977,N_25644,N_25607);
nor U25978 (N_25978,N_25696,N_25625);
nand U25979 (N_25979,N_25686,N_25688);
or U25980 (N_25980,N_25652,N_25562);
nand U25981 (N_25981,N_25541,N_25717);
nand U25982 (N_25982,N_25502,N_25703);
nand U25983 (N_25983,N_25574,N_25631);
xnor U25984 (N_25984,N_25557,N_25571);
xnor U25985 (N_25985,N_25615,N_25588);
nand U25986 (N_25986,N_25548,N_25620);
or U25987 (N_25987,N_25669,N_25632);
nor U25988 (N_25988,N_25651,N_25509);
nor U25989 (N_25989,N_25687,N_25602);
and U25990 (N_25990,N_25628,N_25658);
and U25991 (N_25991,N_25720,N_25510);
and U25992 (N_25992,N_25664,N_25683);
nand U25993 (N_25993,N_25590,N_25641);
xnor U25994 (N_25994,N_25537,N_25560);
nand U25995 (N_25995,N_25583,N_25627);
xor U25996 (N_25996,N_25643,N_25720);
or U25997 (N_25997,N_25550,N_25697);
nor U25998 (N_25998,N_25611,N_25642);
or U25999 (N_25999,N_25660,N_25517);
and U26000 (N_26000,N_25860,N_25811);
or U26001 (N_26001,N_25907,N_25863);
xnor U26002 (N_26002,N_25776,N_25973);
and U26003 (N_26003,N_25932,N_25981);
nor U26004 (N_26004,N_25906,N_25754);
nor U26005 (N_26005,N_25824,N_25814);
and U26006 (N_26006,N_25812,N_25923);
nand U26007 (N_26007,N_25966,N_25866);
nor U26008 (N_26008,N_25825,N_25831);
nor U26009 (N_26009,N_25997,N_25757);
or U26010 (N_26010,N_25947,N_25765);
xor U26011 (N_26011,N_25818,N_25928);
nor U26012 (N_26012,N_25835,N_25959);
and U26013 (N_26013,N_25964,N_25762);
xnor U26014 (N_26014,N_25832,N_25977);
nor U26015 (N_26015,N_25940,N_25882);
nor U26016 (N_26016,N_25950,N_25927);
xor U26017 (N_26017,N_25802,N_25942);
or U26018 (N_26018,N_25750,N_25853);
xnor U26019 (N_26019,N_25925,N_25893);
nor U26020 (N_26020,N_25770,N_25931);
or U26021 (N_26021,N_25953,N_25944);
nor U26022 (N_26022,N_25808,N_25985);
or U26023 (N_26023,N_25828,N_25979);
xnor U26024 (N_26024,N_25783,N_25993);
nand U26025 (N_26025,N_25924,N_25852);
and U26026 (N_26026,N_25892,N_25817);
xnor U26027 (N_26027,N_25975,N_25803);
or U26028 (N_26028,N_25798,N_25943);
xor U26029 (N_26029,N_25937,N_25779);
or U26030 (N_26030,N_25810,N_25992);
and U26031 (N_26031,N_25954,N_25991);
nor U26032 (N_26032,N_25797,N_25826);
nor U26033 (N_26033,N_25848,N_25902);
and U26034 (N_26034,N_25837,N_25864);
xnor U26035 (N_26035,N_25965,N_25949);
and U26036 (N_26036,N_25969,N_25995);
nand U26037 (N_26037,N_25794,N_25809);
nor U26038 (N_26038,N_25951,N_25891);
and U26039 (N_26039,N_25912,N_25793);
and U26040 (N_26040,N_25865,N_25871);
nor U26041 (N_26041,N_25933,N_25854);
or U26042 (N_26042,N_25820,N_25861);
and U26043 (N_26043,N_25926,N_25792);
nor U26044 (N_26044,N_25915,N_25956);
nand U26045 (N_26045,N_25968,N_25876);
nand U26046 (N_26046,N_25800,N_25782);
nor U26047 (N_26047,N_25796,N_25843);
and U26048 (N_26048,N_25872,N_25880);
xor U26049 (N_26049,N_25938,N_25886);
nand U26050 (N_26050,N_25913,N_25807);
xor U26051 (N_26051,N_25787,N_25763);
or U26052 (N_26052,N_25986,N_25978);
nand U26053 (N_26053,N_25983,N_25767);
or U26054 (N_26054,N_25948,N_25996);
nor U26055 (N_26055,N_25850,N_25778);
or U26056 (N_26056,N_25781,N_25859);
or U26057 (N_26057,N_25957,N_25879);
and U26058 (N_26058,N_25920,N_25955);
and U26059 (N_26059,N_25791,N_25855);
xor U26060 (N_26060,N_25990,N_25771);
or U26061 (N_26061,N_25769,N_25936);
nand U26062 (N_26062,N_25856,N_25958);
and U26063 (N_26063,N_25921,N_25918);
nor U26064 (N_26064,N_25772,N_25945);
and U26065 (N_26065,N_25858,N_25834);
nand U26066 (N_26066,N_25795,N_25841);
and U26067 (N_26067,N_25887,N_25784);
or U26068 (N_26068,N_25967,N_25786);
or U26069 (N_26069,N_25897,N_25759);
xnor U26070 (N_26070,N_25819,N_25890);
nand U26071 (N_26071,N_25885,N_25846);
and U26072 (N_26072,N_25804,N_25823);
xnor U26073 (N_26073,N_25851,N_25868);
nor U26074 (N_26074,N_25889,N_25976);
and U26075 (N_26075,N_25799,N_25941);
xor U26076 (N_26076,N_25972,N_25939);
xnor U26077 (N_26077,N_25994,N_25908);
nor U26078 (N_26078,N_25884,N_25929);
nand U26079 (N_26079,N_25758,N_25960);
or U26080 (N_26080,N_25919,N_25903);
xnor U26081 (N_26081,N_25962,N_25790);
or U26082 (N_26082,N_25873,N_25999);
nor U26083 (N_26083,N_25988,N_25768);
nor U26084 (N_26084,N_25830,N_25833);
or U26085 (N_26085,N_25961,N_25789);
nor U26086 (N_26086,N_25899,N_25829);
nor U26087 (N_26087,N_25755,N_25914);
and U26088 (N_26088,N_25806,N_25774);
nand U26089 (N_26089,N_25836,N_25756);
nand U26090 (N_26090,N_25984,N_25922);
and U26091 (N_26091,N_25935,N_25916);
or U26092 (N_26092,N_25847,N_25875);
nor U26093 (N_26093,N_25844,N_25930);
nand U26094 (N_26094,N_25840,N_25822);
nand U26095 (N_26095,N_25971,N_25894);
and U26096 (N_26096,N_25963,N_25813);
nor U26097 (N_26097,N_25785,N_25917);
or U26098 (N_26098,N_25815,N_25900);
and U26099 (N_26099,N_25821,N_25801);
xor U26100 (N_26100,N_25895,N_25760);
xor U26101 (N_26101,N_25869,N_25827);
or U26102 (N_26102,N_25909,N_25896);
or U26103 (N_26103,N_25934,N_25881);
and U26104 (N_26104,N_25857,N_25970);
nand U26105 (N_26105,N_25761,N_25842);
and U26106 (N_26106,N_25878,N_25862);
and U26107 (N_26107,N_25870,N_25982);
or U26108 (N_26108,N_25877,N_25780);
nor U26109 (N_26109,N_25816,N_25946);
or U26110 (N_26110,N_25838,N_25751);
nor U26111 (N_26111,N_25905,N_25901);
nor U26112 (N_26112,N_25753,N_25775);
xor U26113 (N_26113,N_25898,N_25998);
nand U26114 (N_26114,N_25952,N_25874);
nor U26115 (N_26115,N_25974,N_25911);
or U26116 (N_26116,N_25910,N_25764);
nand U26117 (N_26117,N_25773,N_25867);
nand U26118 (N_26118,N_25904,N_25788);
and U26119 (N_26119,N_25980,N_25989);
nor U26120 (N_26120,N_25987,N_25888);
nor U26121 (N_26121,N_25752,N_25845);
nand U26122 (N_26122,N_25839,N_25766);
and U26123 (N_26123,N_25883,N_25777);
and U26124 (N_26124,N_25849,N_25805);
xnor U26125 (N_26125,N_25940,N_25879);
nand U26126 (N_26126,N_25862,N_25963);
xnor U26127 (N_26127,N_25848,N_25939);
or U26128 (N_26128,N_25771,N_25891);
or U26129 (N_26129,N_25984,N_25997);
and U26130 (N_26130,N_25928,N_25760);
or U26131 (N_26131,N_25880,N_25984);
nand U26132 (N_26132,N_25797,N_25994);
nor U26133 (N_26133,N_25853,N_25926);
xnor U26134 (N_26134,N_25773,N_25817);
nor U26135 (N_26135,N_25808,N_25772);
and U26136 (N_26136,N_25764,N_25861);
and U26137 (N_26137,N_25881,N_25776);
xor U26138 (N_26138,N_25755,N_25779);
or U26139 (N_26139,N_25924,N_25937);
xnor U26140 (N_26140,N_25910,N_25775);
nor U26141 (N_26141,N_25828,N_25919);
xor U26142 (N_26142,N_25776,N_25824);
nor U26143 (N_26143,N_25757,N_25799);
nor U26144 (N_26144,N_25791,N_25899);
or U26145 (N_26145,N_25890,N_25849);
nor U26146 (N_26146,N_25912,N_25892);
and U26147 (N_26147,N_25766,N_25812);
or U26148 (N_26148,N_25937,N_25878);
and U26149 (N_26149,N_25800,N_25989);
xnor U26150 (N_26150,N_25955,N_25998);
or U26151 (N_26151,N_25825,N_25868);
xnor U26152 (N_26152,N_25858,N_25888);
and U26153 (N_26153,N_25829,N_25905);
xor U26154 (N_26154,N_25965,N_25824);
or U26155 (N_26155,N_25937,N_25831);
nand U26156 (N_26156,N_25966,N_25976);
or U26157 (N_26157,N_25830,N_25828);
and U26158 (N_26158,N_25780,N_25899);
nand U26159 (N_26159,N_25844,N_25789);
xnor U26160 (N_26160,N_25855,N_25991);
and U26161 (N_26161,N_25902,N_25785);
and U26162 (N_26162,N_25837,N_25804);
nand U26163 (N_26163,N_25936,N_25765);
xnor U26164 (N_26164,N_25764,N_25884);
and U26165 (N_26165,N_25759,N_25770);
nand U26166 (N_26166,N_25829,N_25893);
or U26167 (N_26167,N_25873,N_25757);
and U26168 (N_26168,N_25887,N_25948);
or U26169 (N_26169,N_25994,N_25861);
nand U26170 (N_26170,N_25804,N_25938);
and U26171 (N_26171,N_25923,N_25988);
nand U26172 (N_26172,N_25839,N_25997);
and U26173 (N_26173,N_25878,N_25764);
xor U26174 (N_26174,N_25964,N_25878);
nor U26175 (N_26175,N_25785,N_25998);
nor U26176 (N_26176,N_25909,N_25844);
nor U26177 (N_26177,N_25833,N_25882);
nor U26178 (N_26178,N_25925,N_25815);
or U26179 (N_26179,N_25816,N_25942);
or U26180 (N_26180,N_25966,N_25810);
nand U26181 (N_26181,N_25982,N_25797);
or U26182 (N_26182,N_25781,N_25912);
or U26183 (N_26183,N_25956,N_25884);
nor U26184 (N_26184,N_25943,N_25783);
or U26185 (N_26185,N_25822,N_25982);
xnor U26186 (N_26186,N_25901,N_25823);
or U26187 (N_26187,N_25883,N_25807);
and U26188 (N_26188,N_25948,N_25816);
nand U26189 (N_26189,N_25920,N_25887);
or U26190 (N_26190,N_25897,N_25905);
nand U26191 (N_26191,N_25783,N_25799);
nand U26192 (N_26192,N_25870,N_25926);
xor U26193 (N_26193,N_25947,N_25987);
nor U26194 (N_26194,N_25925,N_25845);
xor U26195 (N_26195,N_25989,N_25792);
xor U26196 (N_26196,N_25860,N_25912);
or U26197 (N_26197,N_25924,N_25896);
xor U26198 (N_26198,N_25831,N_25992);
nor U26199 (N_26199,N_25825,N_25986);
nor U26200 (N_26200,N_25831,N_25921);
or U26201 (N_26201,N_25963,N_25933);
nor U26202 (N_26202,N_25819,N_25913);
nand U26203 (N_26203,N_25988,N_25897);
nand U26204 (N_26204,N_25959,N_25978);
nor U26205 (N_26205,N_25918,N_25795);
nand U26206 (N_26206,N_25844,N_25767);
nor U26207 (N_26207,N_25932,N_25826);
and U26208 (N_26208,N_25963,N_25971);
nor U26209 (N_26209,N_25970,N_25965);
nor U26210 (N_26210,N_25758,N_25927);
nor U26211 (N_26211,N_25905,N_25808);
nor U26212 (N_26212,N_25783,N_25776);
and U26213 (N_26213,N_25940,N_25878);
nand U26214 (N_26214,N_25974,N_25930);
or U26215 (N_26215,N_25804,N_25831);
or U26216 (N_26216,N_25795,N_25804);
and U26217 (N_26217,N_25807,N_25977);
or U26218 (N_26218,N_25842,N_25844);
and U26219 (N_26219,N_25842,N_25798);
nand U26220 (N_26220,N_25866,N_25881);
nand U26221 (N_26221,N_25769,N_25864);
and U26222 (N_26222,N_25757,N_25897);
xnor U26223 (N_26223,N_25845,N_25874);
and U26224 (N_26224,N_25799,N_25865);
nand U26225 (N_26225,N_25961,N_25873);
and U26226 (N_26226,N_25993,N_25801);
or U26227 (N_26227,N_25961,N_25819);
or U26228 (N_26228,N_25925,N_25896);
xor U26229 (N_26229,N_25995,N_25863);
nand U26230 (N_26230,N_25777,N_25898);
xor U26231 (N_26231,N_25756,N_25989);
nor U26232 (N_26232,N_25994,N_25925);
xnor U26233 (N_26233,N_25791,N_25926);
xnor U26234 (N_26234,N_25975,N_25778);
and U26235 (N_26235,N_25826,N_25929);
nor U26236 (N_26236,N_25994,N_25844);
nor U26237 (N_26237,N_25911,N_25922);
xnor U26238 (N_26238,N_25923,N_25871);
nand U26239 (N_26239,N_25914,N_25912);
xnor U26240 (N_26240,N_25951,N_25795);
nand U26241 (N_26241,N_25919,N_25772);
nand U26242 (N_26242,N_25987,N_25999);
and U26243 (N_26243,N_25980,N_25941);
xnor U26244 (N_26244,N_25987,N_25819);
and U26245 (N_26245,N_25898,N_25807);
or U26246 (N_26246,N_25751,N_25972);
nand U26247 (N_26247,N_25877,N_25931);
xnor U26248 (N_26248,N_25776,N_25997);
nor U26249 (N_26249,N_25995,N_25948);
and U26250 (N_26250,N_26123,N_26017);
xnor U26251 (N_26251,N_26182,N_26047);
or U26252 (N_26252,N_26005,N_26074);
xor U26253 (N_26253,N_26231,N_26156);
nand U26254 (N_26254,N_26011,N_26245);
nor U26255 (N_26255,N_26181,N_26093);
and U26256 (N_26256,N_26111,N_26016);
nand U26257 (N_26257,N_26203,N_26185);
and U26258 (N_26258,N_26078,N_26157);
nor U26259 (N_26259,N_26110,N_26080);
nand U26260 (N_26260,N_26205,N_26006);
nand U26261 (N_26261,N_26153,N_26147);
xnor U26262 (N_26262,N_26090,N_26115);
xnor U26263 (N_26263,N_26081,N_26099);
nor U26264 (N_26264,N_26152,N_26237);
nor U26265 (N_26265,N_26071,N_26077);
nand U26266 (N_26266,N_26024,N_26184);
or U26267 (N_26267,N_26201,N_26218);
nand U26268 (N_26268,N_26094,N_26113);
and U26269 (N_26269,N_26112,N_26163);
nand U26270 (N_26270,N_26073,N_26079);
xor U26271 (N_26271,N_26229,N_26188);
or U26272 (N_26272,N_26215,N_26100);
nand U26273 (N_26273,N_26134,N_26054);
and U26274 (N_26274,N_26133,N_26155);
nand U26275 (N_26275,N_26014,N_26030);
and U26276 (N_26276,N_26043,N_26198);
and U26277 (N_26277,N_26150,N_26171);
and U26278 (N_26278,N_26132,N_26227);
or U26279 (N_26279,N_26128,N_26086);
nand U26280 (N_26280,N_26041,N_26050);
nand U26281 (N_26281,N_26087,N_26162);
xnor U26282 (N_26282,N_26022,N_26160);
and U26283 (N_26283,N_26221,N_26052);
and U26284 (N_26284,N_26097,N_26235);
nor U26285 (N_26285,N_26217,N_26173);
xor U26286 (N_26286,N_26039,N_26108);
nand U26287 (N_26287,N_26020,N_26142);
xor U26288 (N_26288,N_26202,N_26121);
xnor U26289 (N_26289,N_26025,N_26139);
nand U26290 (N_26290,N_26122,N_26089);
and U26291 (N_26291,N_26028,N_26242);
nand U26292 (N_26292,N_26161,N_26058);
and U26293 (N_26293,N_26238,N_26145);
or U26294 (N_26294,N_26210,N_26199);
nand U26295 (N_26295,N_26166,N_26040);
nand U26296 (N_26296,N_26053,N_26228);
and U26297 (N_26297,N_26083,N_26234);
nand U26298 (N_26298,N_26158,N_26044);
xnor U26299 (N_26299,N_26082,N_26193);
nor U26300 (N_26300,N_26008,N_26037);
nor U26301 (N_26301,N_26032,N_26051);
nand U26302 (N_26302,N_26149,N_26222);
nor U26303 (N_26303,N_26187,N_26179);
xor U26304 (N_26304,N_26243,N_26114);
or U26305 (N_26305,N_26164,N_26033);
or U26306 (N_26306,N_26061,N_26177);
and U26307 (N_26307,N_26224,N_26137);
nor U26308 (N_26308,N_26140,N_26023);
or U26309 (N_26309,N_26176,N_26118);
or U26310 (N_26310,N_26214,N_26236);
or U26311 (N_26311,N_26021,N_26013);
xnor U26312 (N_26312,N_26106,N_26146);
nor U26313 (N_26313,N_26064,N_26127);
or U26314 (N_26314,N_26246,N_26190);
and U26315 (N_26315,N_26216,N_26026);
xnor U26316 (N_26316,N_26069,N_26247);
and U26317 (N_26317,N_26129,N_26038);
or U26318 (N_26318,N_26117,N_26101);
or U26319 (N_26319,N_26104,N_26151);
or U26320 (N_26320,N_26131,N_26105);
and U26321 (N_26321,N_26056,N_26000);
or U26322 (N_26322,N_26042,N_26170);
xor U26323 (N_26323,N_26211,N_26136);
and U26324 (N_26324,N_26027,N_26143);
and U26325 (N_26325,N_26168,N_26249);
xor U26326 (N_26326,N_26065,N_26055);
nor U26327 (N_26327,N_26195,N_26148);
and U26328 (N_26328,N_26219,N_26057);
and U26329 (N_26329,N_26107,N_26075);
nand U26330 (N_26330,N_26046,N_26049);
or U26331 (N_26331,N_26126,N_26141);
xor U26332 (N_26332,N_26169,N_26240);
or U26333 (N_26333,N_26091,N_26220);
or U26334 (N_26334,N_26098,N_26072);
nor U26335 (N_26335,N_26095,N_26204);
or U26336 (N_26336,N_26223,N_26036);
xor U26337 (N_26337,N_26230,N_26189);
xnor U26338 (N_26338,N_26062,N_26186);
and U26339 (N_26339,N_26096,N_26088);
nor U26340 (N_26340,N_26120,N_26174);
xor U26341 (N_26341,N_26029,N_26208);
nand U26342 (N_26342,N_26125,N_26226);
or U26343 (N_26343,N_26070,N_26019);
and U26344 (N_26344,N_26035,N_26084);
nand U26345 (N_26345,N_26172,N_26241);
nor U26346 (N_26346,N_26233,N_26119);
or U26347 (N_26347,N_26196,N_26109);
and U26348 (N_26348,N_26175,N_26085);
and U26349 (N_26349,N_26031,N_26213);
or U26350 (N_26350,N_26165,N_26209);
nor U26351 (N_26351,N_26138,N_26180);
and U26352 (N_26352,N_26015,N_26154);
nand U26353 (N_26353,N_26192,N_26178);
or U26354 (N_26354,N_26018,N_26194);
nor U26355 (N_26355,N_26059,N_26124);
and U26356 (N_26356,N_26092,N_26004);
or U26357 (N_26357,N_26068,N_26144);
and U26358 (N_26358,N_26191,N_26001);
or U26359 (N_26359,N_26045,N_26010);
and U26360 (N_26360,N_26063,N_26248);
and U26361 (N_26361,N_26225,N_26012);
and U26362 (N_26362,N_26197,N_26007);
and U26363 (N_26363,N_26066,N_26102);
or U26364 (N_26364,N_26076,N_26135);
and U26365 (N_26365,N_26183,N_26167);
nand U26366 (N_26366,N_26116,N_26207);
and U26367 (N_26367,N_26212,N_26206);
nand U26368 (N_26368,N_26002,N_26034);
nand U26369 (N_26369,N_26009,N_26048);
or U26370 (N_26370,N_26103,N_26239);
and U26371 (N_26371,N_26130,N_26060);
and U26372 (N_26372,N_26200,N_26003);
nand U26373 (N_26373,N_26067,N_26244);
nand U26374 (N_26374,N_26159,N_26232);
or U26375 (N_26375,N_26119,N_26176);
nor U26376 (N_26376,N_26029,N_26238);
and U26377 (N_26377,N_26127,N_26025);
and U26378 (N_26378,N_26013,N_26151);
nor U26379 (N_26379,N_26239,N_26078);
xor U26380 (N_26380,N_26185,N_26111);
nand U26381 (N_26381,N_26024,N_26035);
or U26382 (N_26382,N_26018,N_26140);
xor U26383 (N_26383,N_26060,N_26178);
and U26384 (N_26384,N_26190,N_26004);
or U26385 (N_26385,N_26084,N_26162);
and U26386 (N_26386,N_26059,N_26127);
and U26387 (N_26387,N_26033,N_26195);
nor U26388 (N_26388,N_26077,N_26115);
nor U26389 (N_26389,N_26194,N_26175);
xor U26390 (N_26390,N_26159,N_26248);
and U26391 (N_26391,N_26205,N_26084);
and U26392 (N_26392,N_26217,N_26157);
xor U26393 (N_26393,N_26245,N_26068);
nand U26394 (N_26394,N_26226,N_26014);
and U26395 (N_26395,N_26017,N_26205);
and U26396 (N_26396,N_26040,N_26004);
or U26397 (N_26397,N_26147,N_26108);
xnor U26398 (N_26398,N_26142,N_26238);
nand U26399 (N_26399,N_26140,N_26064);
nor U26400 (N_26400,N_26022,N_26005);
or U26401 (N_26401,N_26208,N_26055);
xnor U26402 (N_26402,N_26161,N_26033);
nand U26403 (N_26403,N_26006,N_26187);
xnor U26404 (N_26404,N_26151,N_26135);
and U26405 (N_26405,N_26246,N_26067);
nor U26406 (N_26406,N_26138,N_26136);
or U26407 (N_26407,N_26231,N_26144);
and U26408 (N_26408,N_26182,N_26246);
xnor U26409 (N_26409,N_26135,N_26206);
and U26410 (N_26410,N_26026,N_26047);
xor U26411 (N_26411,N_26069,N_26090);
nand U26412 (N_26412,N_26236,N_26171);
xor U26413 (N_26413,N_26147,N_26112);
and U26414 (N_26414,N_26198,N_26210);
nand U26415 (N_26415,N_26143,N_26242);
or U26416 (N_26416,N_26191,N_26079);
or U26417 (N_26417,N_26005,N_26057);
nor U26418 (N_26418,N_26132,N_26142);
or U26419 (N_26419,N_26008,N_26138);
and U26420 (N_26420,N_26102,N_26165);
and U26421 (N_26421,N_26025,N_26102);
nor U26422 (N_26422,N_26119,N_26091);
xor U26423 (N_26423,N_26234,N_26014);
nand U26424 (N_26424,N_26103,N_26152);
nor U26425 (N_26425,N_26089,N_26076);
and U26426 (N_26426,N_26222,N_26026);
xor U26427 (N_26427,N_26145,N_26038);
nor U26428 (N_26428,N_26043,N_26016);
and U26429 (N_26429,N_26126,N_26166);
nor U26430 (N_26430,N_26197,N_26111);
xnor U26431 (N_26431,N_26227,N_26146);
xor U26432 (N_26432,N_26089,N_26092);
and U26433 (N_26433,N_26047,N_26121);
or U26434 (N_26434,N_26169,N_26090);
or U26435 (N_26435,N_26112,N_26118);
and U26436 (N_26436,N_26051,N_26247);
nor U26437 (N_26437,N_26027,N_26072);
and U26438 (N_26438,N_26144,N_26223);
or U26439 (N_26439,N_26194,N_26100);
or U26440 (N_26440,N_26239,N_26159);
nand U26441 (N_26441,N_26110,N_26243);
xor U26442 (N_26442,N_26185,N_26047);
and U26443 (N_26443,N_26122,N_26125);
or U26444 (N_26444,N_26164,N_26179);
nand U26445 (N_26445,N_26102,N_26236);
xor U26446 (N_26446,N_26213,N_26051);
nand U26447 (N_26447,N_26125,N_26166);
or U26448 (N_26448,N_26186,N_26235);
nor U26449 (N_26449,N_26043,N_26138);
and U26450 (N_26450,N_26045,N_26144);
xnor U26451 (N_26451,N_26129,N_26212);
nand U26452 (N_26452,N_26133,N_26169);
nor U26453 (N_26453,N_26180,N_26164);
nor U26454 (N_26454,N_26143,N_26114);
nand U26455 (N_26455,N_26105,N_26064);
nand U26456 (N_26456,N_26206,N_26055);
and U26457 (N_26457,N_26081,N_26085);
nand U26458 (N_26458,N_26172,N_26127);
or U26459 (N_26459,N_26059,N_26175);
or U26460 (N_26460,N_26112,N_26151);
nor U26461 (N_26461,N_26024,N_26178);
and U26462 (N_26462,N_26119,N_26074);
and U26463 (N_26463,N_26061,N_26046);
nor U26464 (N_26464,N_26018,N_26231);
xnor U26465 (N_26465,N_26007,N_26097);
xnor U26466 (N_26466,N_26111,N_26191);
xor U26467 (N_26467,N_26166,N_26123);
or U26468 (N_26468,N_26056,N_26109);
and U26469 (N_26469,N_26227,N_26222);
and U26470 (N_26470,N_26101,N_26205);
and U26471 (N_26471,N_26003,N_26070);
and U26472 (N_26472,N_26088,N_26030);
or U26473 (N_26473,N_26108,N_26047);
or U26474 (N_26474,N_26107,N_26047);
or U26475 (N_26475,N_26215,N_26005);
nand U26476 (N_26476,N_26174,N_26230);
or U26477 (N_26477,N_26184,N_26245);
nand U26478 (N_26478,N_26217,N_26008);
or U26479 (N_26479,N_26184,N_26237);
and U26480 (N_26480,N_26012,N_26141);
xor U26481 (N_26481,N_26038,N_26139);
or U26482 (N_26482,N_26185,N_26085);
and U26483 (N_26483,N_26020,N_26184);
and U26484 (N_26484,N_26032,N_26072);
or U26485 (N_26485,N_26219,N_26047);
nor U26486 (N_26486,N_26155,N_26223);
or U26487 (N_26487,N_26048,N_26223);
nand U26488 (N_26488,N_26125,N_26238);
xnor U26489 (N_26489,N_26111,N_26109);
and U26490 (N_26490,N_26150,N_26177);
nand U26491 (N_26491,N_26245,N_26242);
or U26492 (N_26492,N_26087,N_26190);
xnor U26493 (N_26493,N_26062,N_26214);
or U26494 (N_26494,N_26214,N_26096);
xnor U26495 (N_26495,N_26116,N_26148);
nor U26496 (N_26496,N_26065,N_26197);
or U26497 (N_26497,N_26069,N_26122);
and U26498 (N_26498,N_26162,N_26156);
or U26499 (N_26499,N_26078,N_26012);
nor U26500 (N_26500,N_26298,N_26282);
and U26501 (N_26501,N_26380,N_26400);
and U26502 (N_26502,N_26334,N_26269);
or U26503 (N_26503,N_26396,N_26439);
xnor U26504 (N_26504,N_26381,N_26317);
nand U26505 (N_26505,N_26295,N_26277);
or U26506 (N_26506,N_26411,N_26426);
and U26507 (N_26507,N_26284,N_26356);
xor U26508 (N_26508,N_26253,N_26430);
or U26509 (N_26509,N_26499,N_26441);
nor U26510 (N_26510,N_26329,N_26261);
nand U26511 (N_26511,N_26364,N_26325);
xor U26512 (N_26512,N_26466,N_26442);
and U26513 (N_26513,N_26434,N_26348);
nand U26514 (N_26514,N_26266,N_26273);
xnor U26515 (N_26515,N_26283,N_26330);
nor U26516 (N_26516,N_26459,N_26285);
and U26517 (N_26517,N_26491,N_26300);
and U26518 (N_26518,N_26332,N_26395);
nand U26519 (N_26519,N_26357,N_26346);
nor U26520 (N_26520,N_26389,N_26262);
nand U26521 (N_26521,N_26449,N_26256);
or U26522 (N_26522,N_26342,N_26265);
or U26523 (N_26523,N_26331,N_26319);
nand U26524 (N_26524,N_26456,N_26454);
nand U26525 (N_26525,N_26264,N_26323);
nor U26526 (N_26526,N_26363,N_26316);
and U26527 (N_26527,N_26394,N_26350);
nor U26528 (N_26528,N_26289,N_26406);
xnor U26529 (N_26529,N_26290,N_26294);
xor U26530 (N_26530,N_26451,N_26421);
nand U26531 (N_26531,N_26481,N_26445);
nor U26532 (N_26532,N_26494,N_26255);
and U26533 (N_26533,N_26271,N_26372);
or U26534 (N_26534,N_26401,N_26448);
nand U26535 (N_26535,N_26383,N_26384);
nor U26536 (N_26536,N_26299,N_26305);
nand U26537 (N_26537,N_26413,N_26464);
or U26538 (N_26538,N_26309,N_26361);
nand U26539 (N_26539,N_26333,N_26418);
xor U26540 (N_26540,N_26475,N_26352);
and U26541 (N_26541,N_26374,N_26388);
nor U26542 (N_26542,N_26292,N_26447);
nand U26543 (N_26543,N_26251,N_26274);
nor U26544 (N_26544,N_26444,N_26485);
and U26545 (N_26545,N_26250,N_26286);
or U26546 (N_26546,N_26428,N_26386);
and U26547 (N_26547,N_26267,N_26423);
and U26548 (N_26548,N_26301,N_26482);
xor U26549 (N_26549,N_26484,N_26358);
nand U26550 (N_26550,N_26417,N_26322);
nand U26551 (N_26551,N_26368,N_26341);
or U26552 (N_26552,N_26359,N_26349);
and U26553 (N_26553,N_26498,N_26486);
nor U26554 (N_26554,N_26420,N_26462);
nand U26555 (N_26555,N_26488,N_26260);
nand U26556 (N_26556,N_26327,N_26478);
xor U26557 (N_26557,N_26414,N_26258);
nor U26558 (N_26558,N_26391,N_26387);
or U26559 (N_26559,N_26297,N_26446);
nand U26560 (N_26560,N_26440,N_26252);
xor U26561 (N_26561,N_26336,N_26375);
and U26562 (N_26562,N_26480,N_26365);
xor U26563 (N_26563,N_26457,N_26473);
nor U26564 (N_26564,N_26433,N_26438);
nor U26565 (N_26565,N_26477,N_26355);
and U26566 (N_26566,N_26497,N_26405);
nand U26567 (N_26567,N_26338,N_26276);
nand U26568 (N_26568,N_26288,N_26468);
and U26569 (N_26569,N_26326,N_26416);
and U26570 (N_26570,N_26399,N_26419);
and U26571 (N_26571,N_26313,N_26410);
nand U26572 (N_26572,N_26376,N_26487);
xor U26573 (N_26573,N_26312,N_26443);
nand U26574 (N_26574,N_26489,N_26270);
nand U26575 (N_26575,N_26436,N_26351);
nor U26576 (N_26576,N_26345,N_26321);
nand U26577 (N_26577,N_26470,N_26422);
or U26578 (N_26578,N_26385,N_26474);
or U26579 (N_26579,N_26303,N_26369);
nand U26580 (N_26580,N_26450,N_26463);
xnor U26581 (N_26581,N_26461,N_26254);
nor U26582 (N_26582,N_26268,N_26408);
or U26583 (N_26583,N_26307,N_26296);
xor U26584 (N_26584,N_26409,N_26427);
or U26585 (N_26585,N_26437,N_26490);
nand U26586 (N_26586,N_26278,N_26458);
or U26587 (N_26587,N_26367,N_26318);
nor U26588 (N_26588,N_26471,N_26467);
nor U26589 (N_26589,N_26320,N_26393);
nor U26590 (N_26590,N_26306,N_26453);
nor U26591 (N_26591,N_26347,N_26378);
and U26592 (N_26592,N_26460,N_26435);
nand U26593 (N_26593,N_26302,N_26407);
xor U26594 (N_26594,N_26455,N_26452);
nor U26595 (N_26595,N_26310,N_26263);
or U26596 (N_26596,N_26280,N_26415);
xor U26597 (N_26597,N_26343,N_26382);
nand U26598 (N_26598,N_26371,N_26315);
or U26599 (N_26599,N_26311,N_26404);
and U26600 (N_26600,N_26259,N_26370);
and U26601 (N_26601,N_26314,N_26353);
and U26602 (N_26602,N_26291,N_26287);
xnor U26603 (N_26603,N_26360,N_26379);
nor U26604 (N_26604,N_26412,N_26469);
or U26605 (N_26605,N_26425,N_26373);
xor U26606 (N_26606,N_26304,N_26493);
and U26607 (N_26607,N_26337,N_26279);
nor U26608 (N_26608,N_26403,N_26472);
nor U26609 (N_26609,N_26272,N_26366);
nand U26610 (N_26610,N_26308,N_26495);
or U26611 (N_26611,N_26492,N_26340);
xor U26612 (N_26612,N_26362,N_26424);
nand U26613 (N_26613,N_26432,N_26275);
nand U26614 (N_26614,N_26398,N_26431);
or U26615 (N_26615,N_26281,N_26339);
nand U26616 (N_26616,N_26257,N_26465);
nand U26617 (N_26617,N_26496,N_26328);
nand U26618 (N_26618,N_26397,N_26479);
nand U26619 (N_26619,N_26354,N_26377);
and U26620 (N_26620,N_26483,N_26344);
nand U26621 (N_26621,N_26324,N_26293);
xor U26622 (N_26622,N_26476,N_26429);
nand U26623 (N_26623,N_26402,N_26335);
nand U26624 (N_26624,N_26392,N_26390);
and U26625 (N_26625,N_26485,N_26489);
and U26626 (N_26626,N_26446,N_26309);
or U26627 (N_26627,N_26371,N_26487);
xnor U26628 (N_26628,N_26307,N_26409);
nor U26629 (N_26629,N_26261,N_26432);
and U26630 (N_26630,N_26474,N_26483);
or U26631 (N_26631,N_26424,N_26315);
nor U26632 (N_26632,N_26424,N_26370);
nor U26633 (N_26633,N_26320,N_26356);
and U26634 (N_26634,N_26421,N_26317);
or U26635 (N_26635,N_26264,N_26374);
and U26636 (N_26636,N_26359,N_26472);
xor U26637 (N_26637,N_26449,N_26451);
nor U26638 (N_26638,N_26405,N_26266);
or U26639 (N_26639,N_26424,N_26298);
xor U26640 (N_26640,N_26300,N_26257);
nand U26641 (N_26641,N_26495,N_26315);
nand U26642 (N_26642,N_26312,N_26437);
nor U26643 (N_26643,N_26310,N_26290);
or U26644 (N_26644,N_26432,N_26357);
xor U26645 (N_26645,N_26474,N_26452);
xor U26646 (N_26646,N_26286,N_26422);
or U26647 (N_26647,N_26473,N_26490);
and U26648 (N_26648,N_26492,N_26475);
or U26649 (N_26649,N_26390,N_26326);
or U26650 (N_26650,N_26283,N_26455);
nor U26651 (N_26651,N_26409,N_26480);
xnor U26652 (N_26652,N_26394,N_26377);
or U26653 (N_26653,N_26360,N_26385);
nor U26654 (N_26654,N_26368,N_26268);
and U26655 (N_26655,N_26285,N_26359);
and U26656 (N_26656,N_26455,N_26409);
or U26657 (N_26657,N_26285,N_26484);
nor U26658 (N_26658,N_26374,N_26301);
nor U26659 (N_26659,N_26375,N_26391);
xnor U26660 (N_26660,N_26492,N_26294);
and U26661 (N_26661,N_26374,N_26338);
or U26662 (N_26662,N_26422,N_26257);
nor U26663 (N_26663,N_26282,N_26289);
nor U26664 (N_26664,N_26490,N_26277);
nor U26665 (N_26665,N_26463,N_26340);
nand U26666 (N_26666,N_26486,N_26372);
xnor U26667 (N_26667,N_26397,N_26460);
nand U26668 (N_26668,N_26290,N_26412);
and U26669 (N_26669,N_26415,N_26412);
and U26670 (N_26670,N_26324,N_26476);
nor U26671 (N_26671,N_26345,N_26354);
and U26672 (N_26672,N_26430,N_26318);
nor U26673 (N_26673,N_26448,N_26459);
nand U26674 (N_26674,N_26337,N_26304);
and U26675 (N_26675,N_26359,N_26445);
or U26676 (N_26676,N_26447,N_26253);
and U26677 (N_26677,N_26372,N_26324);
nand U26678 (N_26678,N_26446,N_26486);
or U26679 (N_26679,N_26493,N_26366);
or U26680 (N_26680,N_26291,N_26370);
or U26681 (N_26681,N_26428,N_26451);
or U26682 (N_26682,N_26497,N_26359);
nand U26683 (N_26683,N_26312,N_26460);
and U26684 (N_26684,N_26464,N_26446);
xor U26685 (N_26685,N_26330,N_26490);
xor U26686 (N_26686,N_26461,N_26306);
or U26687 (N_26687,N_26289,N_26364);
nand U26688 (N_26688,N_26327,N_26331);
nor U26689 (N_26689,N_26286,N_26334);
xor U26690 (N_26690,N_26394,N_26318);
and U26691 (N_26691,N_26416,N_26367);
nand U26692 (N_26692,N_26309,N_26396);
and U26693 (N_26693,N_26382,N_26324);
nand U26694 (N_26694,N_26262,N_26430);
xor U26695 (N_26695,N_26348,N_26472);
nand U26696 (N_26696,N_26395,N_26264);
nor U26697 (N_26697,N_26301,N_26381);
or U26698 (N_26698,N_26345,N_26438);
and U26699 (N_26699,N_26438,N_26382);
or U26700 (N_26700,N_26441,N_26329);
xnor U26701 (N_26701,N_26358,N_26377);
and U26702 (N_26702,N_26371,N_26337);
and U26703 (N_26703,N_26402,N_26495);
nand U26704 (N_26704,N_26417,N_26426);
nor U26705 (N_26705,N_26349,N_26348);
nor U26706 (N_26706,N_26306,N_26376);
or U26707 (N_26707,N_26460,N_26420);
nor U26708 (N_26708,N_26338,N_26304);
xor U26709 (N_26709,N_26436,N_26362);
or U26710 (N_26710,N_26387,N_26471);
or U26711 (N_26711,N_26333,N_26420);
or U26712 (N_26712,N_26289,N_26376);
and U26713 (N_26713,N_26333,N_26351);
and U26714 (N_26714,N_26313,N_26335);
nand U26715 (N_26715,N_26355,N_26499);
nor U26716 (N_26716,N_26439,N_26268);
nor U26717 (N_26717,N_26337,N_26372);
nor U26718 (N_26718,N_26290,N_26433);
or U26719 (N_26719,N_26350,N_26271);
nor U26720 (N_26720,N_26380,N_26251);
xor U26721 (N_26721,N_26399,N_26380);
xor U26722 (N_26722,N_26416,N_26420);
or U26723 (N_26723,N_26444,N_26467);
or U26724 (N_26724,N_26368,N_26313);
xnor U26725 (N_26725,N_26338,N_26328);
xor U26726 (N_26726,N_26264,N_26414);
xnor U26727 (N_26727,N_26310,N_26304);
nor U26728 (N_26728,N_26418,N_26293);
and U26729 (N_26729,N_26266,N_26395);
and U26730 (N_26730,N_26324,N_26276);
nor U26731 (N_26731,N_26412,N_26423);
and U26732 (N_26732,N_26460,N_26469);
nor U26733 (N_26733,N_26401,N_26354);
nor U26734 (N_26734,N_26279,N_26467);
nand U26735 (N_26735,N_26433,N_26454);
nand U26736 (N_26736,N_26293,N_26450);
or U26737 (N_26737,N_26382,N_26490);
xor U26738 (N_26738,N_26424,N_26263);
nand U26739 (N_26739,N_26301,N_26268);
or U26740 (N_26740,N_26393,N_26472);
xnor U26741 (N_26741,N_26257,N_26402);
and U26742 (N_26742,N_26320,N_26251);
nor U26743 (N_26743,N_26359,N_26298);
xnor U26744 (N_26744,N_26342,N_26390);
or U26745 (N_26745,N_26254,N_26370);
xor U26746 (N_26746,N_26339,N_26318);
nor U26747 (N_26747,N_26250,N_26264);
or U26748 (N_26748,N_26347,N_26256);
and U26749 (N_26749,N_26272,N_26459);
or U26750 (N_26750,N_26620,N_26735);
or U26751 (N_26751,N_26542,N_26636);
and U26752 (N_26752,N_26531,N_26611);
or U26753 (N_26753,N_26548,N_26603);
or U26754 (N_26754,N_26514,N_26709);
and U26755 (N_26755,N_26509,N_26608);
nor U26756 (N_26756,N_26556,N_26551);
xnor U26757 (N_26757,N_26692,N_26663);
or U26758 (N_26758,N_26552,N_26665);
nor U26759 (N_26759,N_26713,N_26572);
or U26760 (N_26760,N_26736,N_26725);
nand U26761 (N_26761,N_26749,N_26539);
xnor U26762 (N_26762,N_26724,N_26529);
nand U26763 (N_26763,N_26717,N_26716);
nor U26764 (N_26764,N_26567,N_26530);
and U26765 (N_26765,N_26670,N_26673);
nor U26766 (N_26766,N_26693,N_26597);
xnor U26767 (N_26767,N_26525,N_26671);
or U26768 (N_26768,N_26591,N_26545);
and U26769 (N_26769,N_26642,N_26721);
or U26770 (N_26770,N_26643,N_26558);
nand U26771 (N_26771,N_26685,N_26571);
and U26772 (N_26772,N_26655,N_26568);
nor U26773 (N_26773,N_26657,N_26607);
or U26774 (N_26774,N_26557,N_26700);
or U26775 (N_26775,N_26689,N_26619);
or U26776 (N_26776,N_26744,N_26522);
nor U26777 (N_26777,N_26511,N_26645);
xnor U26778 (N_26778,N_26742,N_26659);
nand U26779 (N_26779,N_26638,N_26690);
nand U26780 (N_26780,N_26669,N_26602);
xnor U26781 (N_26781,N_26708,N_26565);
nor U26782 (N_26782,N_26569,N_26695);
or U26783 (N_26783,N_26500,N_26507);
or U26784 (N_26784,N_26686,N_26622);
xor U26785 (N_26785,N_26628,N_26730);
or U26786 (N_26786,N_26618,N_26649);
nor U26787 (N_26787,N_26560,N_26647);
or U26788 (N_26788,N_26653,N_26694);
xnor U26789 (N_26789,N_26743,N_26578);
xor U26790 (N_26790,N_26594,N_26727);
and U26791 (N_26791,N_26621,N_26632);
nand U26792 (N_26792,N_26555,N_26606);
or U26793 (N_26793,N_26661,N_26634);
nand U26794 (N_26794,N_26595,N_26515);
xor U26795 (N_26795,N_26523,N_26596);
nand U26796 (N_26796,N_26626,N_26588);
xor U26797 (N_26797,N_26748,N_26741);
nor U26798 (N_26798,N_26575,N_26520);
or U26799 (N_26799,N_26706,N_26587);
xnor U26800 (N_26800,N_26677,N_26691);
xor U26801 (N_26801,N_26605,N_26697);
nand U26802 (N_26802,N_26650,N_26526);
nor U26803 (N_26803,N_26581,N_26517);
and U26804 (N_26804,N_26633,N_26512);
or U26805 (N_26805,N_26674,N_26651);
or U26806 (N_26806,N_26711,N_26519);
nor U26807 (N_26807,N_26687,N_26723);
nand U26808 (N_26808,N_26561,N_26734);
xnor U26809 (N_26809,N_26590,N_26579);
or U26810 (N_26810,N_26506,N_26583);
and U26811 (N_26811,N_26624,N_26654);
nor U26812 (N_26812,N_26662,N_26646);
or U26813 (N_26813,N_26728,N_26553);
xnor U26814 (N_26814,N_26704,N_26580);
nor U26815 (N_26815,N_26683,N_26546);
xor U26816 (N_26816,N_26714,N_26699);
nor U26817 (N_26817,N_26648,N_26532);
xnor U26818 (N_26818,N_26635,N_26524);
nor U26819 (N_26819,N_26574,N_26640);
or U26820 (N_26820,N_26696,N_26745);
and U26821 (N_26821,N_26533,N_26527);
nand U26822 (N_26822,N_26504,N_26541);
and U26823 (N_26823,N_26678,N_26747);
nor U26824 (N_26824,N_26737,N_26613);
and U26825 (N_26825,N_26722,N_26682);
or U26826 (N_26826,N_26508,N_26564);
nand U26827 (N_26827,N_26710,N_26672);
and U26828 (N_26828,N_26688,N_26652);
nand U26829 (N_26829,N_26679,N_26535);
and U26830 (N_26830,N_26536,N_26598);
or U26831 (N_26831,N_26528,N_26701);
xnor U26832 (N_26832,N_26586,N_26601);
or U26833 (N_26833,N_26680,N_26614);
nand U26834 (N_26834,N_26715,N_26510);
nand U26835 (N_26835,N_26582,N_26549);
and U26836 (N_26836,N_26641,N_26610);
or U26837 (N_26837,N_26609,N_26739);
and U26838 (N_26838,N_26627,N_26738);
xor U26839 (N_26839,N_26538,N_26676);
nand U26840 (N_26840,N_26600,N_26726);
nand U26841 (N_26841,N_26599,N_26684);
or U26842 (N_26842,N_26639,N_26720);
or U26843 (N_26843,N_26570,N_26534);
nor U26844 (N_26844,N_26703,N_26584);
or U26845 (N_26845,N_26681,N_26668);
and U26846 (N_26846,N_26516,N_26537);
nor U26847 (N_26847,N_26698,N_26563);
xnor U26848 (N_26848,N_26656,N_26733);
and U26849 (N_26849,N_26585,N_26589);
nand U26850 (N_26850,N_26707,N_26719);
xor U26851 (N_26851,N_26740,N_26518);
and U26852 (N_26852,N_26615,N_26631);
or U26853 (N_26853,N_26521,N_26540);
and U26854 (N_26854,N_26667,N_26718);
and U26855 (N_26855,N_26625,N_26612);
nor U26856 (N_26856,N_26513,N_26550);
or U26857 (N_26857,N_26731,N_26576);
and U26858 (N_26858,N_26562,N_26629);
nand U26859 (N_26859,N_26577,N_26617);
nor U26860 (N_26860,N_26746,N_26623);
and U26861 (N_26861,N_26503,N_26566);
or U26862 (N_26862,N_26675,N_26547);
nor U26863 (N_26863,N_26616,N_26604);
and U26864 (N_26864,N_26573,N_26554);
and U26865 (N_26865,N_26712,N_26664);
and U26866 (N_26866,N_26637,N_26592);
nor U26867 (N_26867,N_26544,N_26630);
xor U26868 (N_26868,N_26644,N_26658);
nor U26869 (N_26869,N_26501,N_26732);
and U26870 (N_26870,N_26729,N_26702);
nor U26871 (N_26871,N_26543,N_26660);
nand U26872 (N_26872,N_26559,N_26502);
nand U26873 (N_26873,N_26593,N_26705);
or U26874 (N_26874,N_26666,N_26505);
or U26875 (N_26875,N_26681,N_26708);
nor U26876 (N_26876,N_26579,N_26571);
nor U26877 (N_26877,N_26619,N_26602);
and U26878 (N_26878,N_26682,N_26564);
and U26879 (N_26879,N_26722,N_26572);
nor U26880 (N_26880,N_26723,N_26508);
and U26881 (N_26881,N_26550,N_26644);
and U26882 (N_26882,N_26557,N_26744);
and U26883 (N_26883,N_26746,N_26677);
nor U26884 (N_26884,N_26605,N_26591);
and U26885 (N_26885,N_26644,N_26535);
and U26886 (N_26886,N_26639,N_26604);
nand U26887 (N_26887,N_26611,N_26602);
nor U26888 (N_26888,N_26524,N_26590);
nand U26889 (N_26889,N_26706,N_26636);
xor U26890 (N_26890,N_26541,N_26538);
nand U26891 (N_26891,N_26736,N_26629);
xnor U26892 (N_26892,N_26501,N_26543);
or U26893 (N_26893,N_26698,N_26726);
nand U26894 (N_26894,N_26568,N_26691);
nor U26895 (N_26895,N_26734,N_26565);
nand U26896 (N_26896,N_26687,N_26528);
nor U26897 (N_26897,N_26651,N_26654);
and U26898 (N_26898,N_26743,N_26611);
and U26899 (N_26899,N_26686,N_26525);
and U26900 (N_26900,N_26636,N_26658);
xnor U26901 (N_26901,N_26710,N_26647);
nor U26902 (N_26902,N_26549,N_26722);
nor U26903 (N_26903,N_26699,N_26534);
nor U26904 (N_26904,N_26739,N_26554);
nor U26905 (N_26905,N_26605,N_26532);
nor U26906 (N_26906,N_26744,N_26578);
xor U26907 (N_26907,N_26719,N_26685);
and U26908 (N_26908,N_26520,N_26634);
nor U26909 (N_26909,N_26696,N_26624);
or U26910 (N_26910,N_26652,N_26631);
and U26911 (N_26911,N_26564,N_26662);
nand U26912 (N_26912,N_26530,N_26667);
nand U26913 (N_26913,N_26553,N_26648);
nand U26914 (N_26914,N_26611,N_26711);
and U26915 (N_26915,N_26578,N_26559);
and U26916 (N_26916,N_26687,N_26571);
or U26917 (N_26917,N_26634,N_26742);
nand U26918 (N_26918,N_26519,N_26609);
xor U26919 (N_26919,N_26688,N_26649);
nand U26920 (N_26920,N_26582,N_26643);
xor U26921 (N_26921,N_26583,N_26712);
nand U26922 (N_26922,N_26718,N_26513);
nor U26923 (N_26923,N_26715,N_26702);
or U26924 (N_26924,N_26567,N_26700);
nand U26925 (N_26925,N_26651,N_26681);
and U26926 (N_26926,N_26712,N_26711);
xor U26927 (N_26927,N_26551,N_26555);
nor U26928 (N_26928,N_26745,N_26579);
nor U26929 (N_26929,N_26628,N_26652);
xor U26930 (N_26930,N_26560,N_26726);
xnor U26931 (N_26931,N_26524,N_26563);
nand U26932 (N_26932,N_26685,N_26512);
nor U26933 (N_26933,N_26530,N_26614);
xor U26934 (N_26934,N_26583,N_26606);
or U26935 (N_26935,N_26615,N_26681);
xnor U26936 (N_26936,N_26644,N_26595);
nand U26937 (N_26937,N_26533,N_26607);
nand U26938 (N_26938,N_26539,N_26737);
nor U26939 (N_26939,N_26551,N_26534);
nor U26940 (N_26940,N_26525,N_26514);
nand U26941 (N_26941,N_26516,N_26661);
nand U26942 (N_26942,N_26593,N_26719);
and U26943 (N_26943,N_26720,N_26611);
nand U26944 (N_26944,N_26667,N_26725);
nor U26945 (N_26945,N_26596,N_26641);
xnor U26946 (N_26946,N_26615,N_26745);
and U26947 (N_26947,N_26545,N_26609);
nor U26948 (N_26948,N_26612,N_26723);
and U26949 (N_26949,N_26615,N_26722);
nand U26950 (N_26950,N_26580,N_26746);
nor U26951 (N_26951,N_26589,N_26563);
nor U26952 (N_26952,N_26533,N_26736);
xor U26953 (N_26953,N_26698,N_26637);
or U26954 (N_26954,N_26666,N_26508);
xnor U26955 (N_26955,N_26615,N_26691);
xnor U26956 (N_26956,N_26731,N_26658);
or U26957 (N_26957,N_26608,N_26596);
and U26958 (N_26958,N_26698,N_26677);
xnor U26959 (N_26959,N_26648,N_26558);
xnor U26960 (N_26960,N_26513,N_26519);
xnor U26961 (N_26961,N_26737,N_26599);
nor U26962 (N_26962,N_26667,N_26560);
or U26963 (N_26963,N_26678,N_26657);
or U26964 (N_26964,N_26510,N_26523);
or U26965 (N_26965,N_26601,N_26554);
xnor U26966 (N_26966,N_26661,N_26537);
xnor U26967 (N_26967,N_26514,N_26673);
xor U26968 (N_26968,N_26593,N_26585);
nor U26969 (N_26969,N_26539,N_26500);
nand U26970 (N_26970,N_26563,N_26611);
nand U26971 (N_26971,N_26590,N_26588);
nor U26972 (N_26972,N_26574,N_26521);
or U26973 (N_26973,N_26724,N_26547);
nand U26974 (N_26974,N_26676,N_26554);
or U26975 (N_26975,N_26703,N_26647);
nor U26976 (N_26976,N_26565,N_26560);
nand U26977 (N_26977,N_26726,N_26561);
or U26978 (N_26978,N_26565,N_26648);
xor U26979 (N_26979,N_26569,N_26518);
or U26980 (N_26980,N_26551,N_26546);
nand U26981 (N_26981,N_26506,N_26637);
nor U26982 (N_26982,N_26725,N_26555);
nand U26983 (N_26983,N_26624,N_26636);
and U26984 (N_26984,N_26726,N_26741);
or U26985 (N_26985,N_26707,N_26702);
nor U26986 (N_26986,N_26610,N_26523);
or U26987 (N_26987,N_26540,N_26594);
nand U26988 (N_26988,N_26693,N_26711);
nand U26989 (N_26989,N_26709,N_26693);
nor U26990 (N_26990,N_26716,N_26747);
xor U26991 (N_26991,N_26716,N_26625);
and U26992 (N_26992,N_26554,N_26742);
xor U26993 (N_26993,N_26546,N_26581);
or U26994 (N_26994,N_26530,N_26630);
and U26995 (N_26995,N_26512,N_26653);
xnor U26996 (N_26996,N_26531,N_26640);
or U26997 (N_26997,N_26620,N_26714);
nand U26998 (N_26998,N_26503,N_26555);
nor U26999 (N_26999,N_26630,N_26710);
or U27000 (N_27000,N_26757,N_26917);
xor U27001 (N_27001,N_26891,N_26921);
xor U27002 (N_27002,N_26907,N_26844);
nand U27003 (N_27003,N_26770,N_26780);
xnor U27004 (N_27004,N_26975,N_26803);
nor U27005 (N_27005,N_26877,N_26806);
nand U27006 (N_27006,N_26768,N_26839);
or U27007 (N_27007,N_26793,N_26832);
nand U27008 (N_27008,N_26911,N_26883);
and U27009 (N_27009,N_26868,N_26794);
and U27010 (N_27010,N_26807,N_26769);
xnor U27011 (N_27011,N_26760,N_26960);
xnor U27012 (N_27012,N_26761,N_26808);
nand U27013 (N_27013,N_26901,N_26848);
nor U27014 (N_27014,N_26783,N_26938);
xor U27015 (N_27015,N_26804,N_26967);
or U27016 (N_27016,N_26976,N_26942);
and U27017 (N_27017,N_26995,N_26983);
xnor U27018 (N_27018,N_26772,N_26950);
xnor U27019 (N_27019,N_26999,N_26801);
xnor U27020 (N_27020,N_26961,N_26885);
xnor U27021 (N_27021,N_26771,N_26862);
and U27022 (N_27022,N_26948,N_26859);
nor U27023 (N_27023,N_26860,N_26871);
nand U27024 (N_27024,N_26810,N_26852);
and U27025 (N_27025,N_26905,N_26799);
xnor U27026 (N_27026,N_26865,N_26841);
nor U27027 (N_27027,N_26896,N_26893);
nor U27028 (N_27028,N_26923,N_26812);
or U27029 (N_27029,N_26889,N_26902);
and U27030 (N_27030,N_26984,N_26945);
xor U27031 (N_27031,N_26930,N_26755);
and U27032 (N_27032,N_26888,N_26826);
or U27033 (N_27033,N_26816,N_26867);
and U27034 (N_27034,N_26864,N_26829);
nor U27035 (N_27035,N_26777,N_26773);
nor U27036 (N_27036,N_26998,N_26973);
nand U27037 (N_27037,N_26964,N_26925);
and U27038 (N_27038,N_26785,N_26842);
and U27039 (N_27039,N_26838,N_26971);
and U27040 (N_27040,N_26963,N_26791);
and U27041 (N_27041,N_26924,N_26845);
and U27042 (N_27042,N_26787,N_26957);
nand U27043 (N_27043,N_26929,N_26764);
and U27044 (N_27044,N_26820,N_26750);
nor U27045 (N_27045,N_26792,N_26951);
xor U27046 (N_27046,N_26979,N_26846);
or U27047 (N_27047,N_26805,N_26993);
xnor U27048 (N_27048,N_26878,N_26899);
nor U27049 (N_27049,N_26751,N_26756);
and U27050 (N_27050,N_26782,N_26814);
nor U27051 (N_27051,N_26759,N_26775);
xnor U27052 (N_27052,N_26953,N_26762);
nand U27053 (N_27053,N_26818,N_26895);
or U27054 (N_27054,N_26861,N_26926);
xnor U27055 (N_27055,N_26904,N_26890);
nor U27056 (N_27056,N_26974,N_26752);
and U27057 (N_27057,N_26855,N_26943);
xor U27058 (N_27058,N_26910,N_26798);
xor U27059 (N_27059,N_26856,N_26858);
xnor U27060 (N_27060,N_26851,N_26830);
xor U27061 (N_27061,N_26790,N_26797);
nand U27062 (N_27062,N_26931,N_26834);
xnor U27063 (N_27063,N_26956,N_26965);
nand U27064 (N_27064,N_26968,N_26898);
nor U27065 (N_27065,N_26928,N_26815);
nor U27066 (N_27066,N_26962,N_26766);
xnor U27067 (N_27067,N_26994,N_26966);
and U27068 (N_27068,N_26900,N_26970);
and U27069 (N_27069,N_26914,N_26837);
and U27070 (N_27070,N_26939,N_26997);
or U27071 (N_27071,N_26795,N_26935);
and U27072 (N_27072,N_26934,N_26919);
xnor U27073 (N_27073,N_26932,N_26875);
nor U27074 (N_27074,N_26915,N_26854);
or U27075 (N_27075,N_26765,N_26982);
and U27076 (N_27076,N_26828,N_26958);
nand U27077 (N_27077,N_26922,N_26882);
nand U27078 (N_27078,N_26788,N_26827);
or U27079 (N_27079,N_26909,N_26884);
and U27080 (N_27080,N_26753,N_26823);
xnor U27081 (N_27081,N_26809,N_26949);
nand U27082 (N_27082,N_26774,N_26903);
nor U27083 (N_27083,N_26936,N_26811);
nand U27084 (N_27084,N_26990,N_26813);
xnor U27085 (N_27085,N_26879,N_26824);
and U27086 (N_27086,N_26822,N_26776);
or U27087 (N_27087,N_26941,N_26853);
xnor U27088 (N_27088,N_26933,N_26996);
nand U27089 (N_27089,N_26987,N_26916);
nand U27090 (N_27090,N_26954,N_26763);
or U27091 (N_27091,N_26959,N_26985);
nor U27092 (N_27092,N_26946,N_26988);
or U27093 (N_27093,N_26972,N_26947);
or U27094 (N_27094,N_26863,N_26789);
xor U27095 (N_27095,N_26836,N_26937);
and U27096 (N_27096,N_26840,N_26952);
nand U27097 (N_27097,N_26991,N_26989);
or U27098 (N_27098,N_26870,N_26778);
nor U27099 (N_27099,N_26955,N_26986);
nand U27100 (N_27100,N_26779,N_26850);
and U27101 (N_27101,N_26940,N_26873);
nand U27102 (N_27102,N_26874,N_26819);
and U27103 (N_27103,N_26857,N_26912);
xnor U27104 (N_27104,N_26847,N_26886);
nand U27105 (N_27105,N_26849,N_26908);
nor U27106 (N_27106,N_26918,N_26833);
xor U27107 (N_27107,N_26978,N_26906);
nor U27108 (N_27108,N_26872,N_26866);
nor U27109 (N_27109,N_26781,N_26887);
xor U27110 (N_27110,N_26980,N_26977);
or U27111 (N_27111,N_26981,N_26843);
xor U27112 (N_27112,N_26831,N_26920);
xnor U27113 (N_27113,N_26927,N_26784);
or U27114 (N_27114,N_26897,N_26821);
nand U27115 (N_27115,N_26892,N_26786);
or U27116 (N_27116,N_26880,N_26796);
xnor U27117 (N_27117,N_26894,N_26992);
xor U27118 (N_27118,N_26758,N_26825);
nor U27119 (N_27119,N_26802,N_26913);
and U27120 (N_27120,N_26767,N_26800);
xor U27121 (N_27121,N_26944,N_26835);
or U27122 (N_27122,N_26754,N_26876);
nor U27123 (N_27123,N_26969,N_26869);
xnor U27124 (N_27124,N_26817,N_26881);
nand U27125 (N_27125,N_26877,N_26929);
xor U27126 (N_27126,N_26999,N_26975);
or U27127 (N_27127,N_26970,N_26981);
nor U27128 (N_27128,N_26787,N_26856);
nand U27129 (N_27129,N_26821,N_26942);
or U27130 (N_27130,N_26990,N_26804);
and U27131 (N_27131,N_26863,N_26922);
nand U27132 (N_27132,N_26870,N_26925);
or U27133 (N_27133,N_26962,N_26927);
or U27134 (N_27134,N_26877,N_26780);
xor U27135 (N_27135,N_26763,N_26951);
nand U27136 (N_27136,N_26795,N_26869);
xor U27137 (N_27137,N_26834,N_26797);
nor U27138 (N_27138,N_26991,N_26810);
or U27139 (N_27139,N_26950,N_26764);
nor U27140 (N_27140,N_26979,N_26910);
nor U27141 (N_27141,N_26819,N_26810);
nor U27142 (N_27142,N_26939,N_26863);
nor U27143 (N_27143,N_26869,N_26889);
or U27144 (N_27144,N_26818,N_26772);
nand U27145 (N_27145,N_26832,N_26939);
xor U27146 (N_27146,N_26905,N_26817);
nand U27147 (N_27147,N_26869,N_26784);
nand U27148 (N_27148,N_26845,N_26843);
nand U27149 (N_27149,N_26798,N_26822);
or U27150 (N_27150,N_26830,N_26799);
xnor U27151 (N_27151,N_26953,N_26997);
and U27152 (N_27152,N_26901,N_26816);
nand U27153 (N_27153,N_26888,N_26922);
and U27154 (N_27154,N_26790,N_26998);
xor U27155 (N_27155,N_26763,N_26931);
nand U27156 (N_27156,N_26809,N_26972);
nor U27157 (N_27157,N_26969,N_26948);
xnor U27158 (N_27158,N_26866,N_26907);
xor U27159 (N_27159,N_26992,N_26872);
and U27160 (N_27160,N_26879,N_26769);
xnor U27161 (N_27161,N_26892,N_26873);
nand U27162 (N_27162,N_26778,N_26803);
xor U27163 (N_27163,N_26751,N_26936);
or U27164 (N_27164,N_26776,N_26950);
nor U27165 (N_27165,N_26854,N_26949);
or U27166 (N_27166,N_26867,N_26932);
or U27167 (N_27167,N_26751,N_26833);
xor U27168 (N_27168,N_26912,N_26881);
nand U27169 (N_27169,N_26937,N_26953);
xor U27170 (N_27170,N_26960,N_26979);
or U27171 (N_27171,N_26974,N_26838);
and U27172 (N_27172,N_26855,N_26874);
or U27173 (N_27173,N_26769,N_26824);
and U27174 (N_27174,N_26922,N_26971);
xnor U27175 (N_27175,N_26962,N_26930);
nor U27176 (N_27176,N_26902,N_26804);
and U27177 (N_27177,N_26773,N_26914);
xnor U27178 (N_27178,N_26815,N_26905);
and U27179 (N_27179,N_26912,N_26886);
and U27180 (N_27180,N_26777,N_26834);
nor U27181 (N_27181,N_26916,N_26891);
and U27182 (N_27182,N_26857,N_26939);
and U27183 (N_27183,N_26837,N_26900);
nor U27184 (N_27184,N_26978,N_26920);
nand U27185 (N_27185,N_26806,N_26957);
nor U27186 (N_27186,N_26888,N_26795);
nand U27187 (N_27187,N_26867,N_26902);
xnor U27188 (N_27188,N_26816,N_26872);
xor U27189 (N_27189,N_26857,N_26867);
nor U27190 (N_27190,N_26891,N_26922);
nand U27191 (N_27191,N_26751,N_26968);
nor U27192 (N_27192,N_26974,N_26910);
nand U27193 (N_27193,N_26864,N_26839);
nand U27194 (N_27194,N_26802,N_26804);
nor U27195 (N_27195,N_26818,N_26790);
xor U27196 (N_27196,N_26784,N_26917);
or U27197 (N_27197,N_26824,N_26821);
nand U27198 (N_27198,N_26793,N_26896);
nand U27199 (N_27199,N_26752,N_26758);
nor U27200 (N_27200,N_26842,N_26998);
xor U27201 (N_27201,N_26754,N_26921);
xnor U27202 (N_27202,N_26848,N_26890);
xor U27203 (N_27203,N_26841,N_26815);
xor U27204 (N_27204,N_26975,N_26771);
xor U27205 (N_27205,N_26808,N_26753);
nor U27206 (N_27206,N_26915,N_26998);
or U27207 (N_27207,N_26846,N_26869);
and U27208 (N_27208,N_26880,N_26884);
or U27209 (N_27209,N_26989,N_26848);
or U27210 (N_27210,N_26981,N_26973);
or U27211 (N_27211,N_26752,N_26951);
xnor U27212 (N_27212,N_26939,N_26970);
nand U27213 (N_27213,N_26768,N_26874);
xnor U27214 (N_27214,N_26885,N_26953);
nor U27215 (N_27215,N_26802,N_26758);
nand U27216 (N_27216,N_26922,N_26761);
nor U27217 (N_27217,N_26836,N_26898);
xor U27218 (N_27218,N_26793,N_26996);
or U27219 (N_27219,N_26825,N_26808);
and U27220 (N_27220,N_26947,N_26858);
nand U27221 (N_27221,N_26768,N_26903);
and U27222 (N_27222,N_26869,N_26817);
xor U27223 (N_27223,N_26915,N_26796);
xnor U27224 (N_27224,N_26781,N_26842);
and U27225 (N_27225,N_26993,N_26875);
and U27226 (N_27226,N_26933,N_26892);
and U27227 (N_27227,N_26755,N_26995);
nor U27228 (N_27228,N_26976,N_26977);
nor U27229 (N_27229,N_26848,N_26828);
and U27230 (N_27230,N_26774,N_26932);
or U27231 (N_27231,N_26907,N_26860);
and U27232 (N_27232,N_26897,N_26967);
and U27233 (N_27233,N_26955,N_26880);
and U27234 (N_27234,N_26909,N_26836);
and U27235 (N_27235,N_26852,N_26936);
nor U27236 (N_27236,N_26886,N_26998);
or U27237 (N_27237,N_26958,N_26769);
or U27238 (N_27238,N_26918,N_26926);
nand U27239 (N_27239,N_26966,N_26946);
and U27240 (N_27240,N_26967,N_26793);
xor U27241 (N_27241,N_26911,N_26870);
and U27242 (N_27242,N_26946,N_26775);
or U27243 (N_27243,N_26754,N_26928);
nand U27244 (N_27244,N_26801,N_26873);
xnor U27245 (N_27245,N_26760,N_26833);
nor U27246 (N_27246,N_26983,N_26981);
or U27247 (N_27247,N_26832,N_26812);
or U27248 (N_27248,N_26889,N_26823);
xnor U27249 (N_27249,N_26857,N_26866);
nand U27250 (N_27250,N_27030,N_27226);
nor U27251 (N_27251,N_27077,N_27122);
nand U27252 (N_27252,N_27163,N_27181);
nand U27253 (N_27253,N_27191,N_27115);
nand U27254 (N_27254,N_27141,N_27009);
xor U27255 (N_27255,N_27154,N_27137);
xor U27256 (N_27256,N_27006,N_27056);
xnor U27257 (N_27257,N_27231,N_27209);
and U27258 (N_27258,N_27085,N_27153);
nand U27259 (N_27259,N_27108,N_27066);
nor U27260 (N_27260,N_27214,N_27213);
and U27261 (N_27261,N_27035,N_27167);
and U27262 (N_27262,N_27051,N_27184);
and U27263 (N_27263,N_27227,N_27235);
and U27264 (N_27264,N_27215,N_27211);
nor U27265 (N_27265,N_27240,N_27183);
and U27266 (N_27266,N_27058,N_27133);
xor U27267 (N_27267,N_27216,N_27152);
xor U27268 (N_27268,N_27146,N_27223);
nand U27269 (N_27269,N_27179,N_27245);
nand U27270 (N_27270,N_27020,N_27221);
nand U27271 (N_27271,N_27145,N_27096);
nor U27272 (N_27272,N_27068,N_27074);
nor U27273 (N_27273,N_27094,N_27149);
or U27274 (N_27274,N_27033,N_27039);
xnor U27275 (N_27275,N_27176,N_27186);
nand U27276 (N_27276,N_27243,N_27125);
xor U27277 (N_27277,N_27185,N_27090);
nor U27278 (N_27278,N_27091,N_27158);
and U27279 (N_27279,N_27002,N_27169);
and U27280 (N_27280,N_27099,N_27175);
or U27281 (N_27281,N_27073,N_27109);
nand U27282 (N_27282,N_27246,N_27082);
nor U27283 (N_27283,N_27098,N_27029);
nor U27284 (N_27284,N_27123,N_27248);
xnor U27285 (N_27285,N_27148,N_27088);
nor U27286 (N_27286,N_27062,N_27120);
nand U27287 (N_27287,N_27071,N_27132);
nor U27288 (N_27288,N_27160,N_27220);
nor U27289 (N_27289,N_27157,N_27206);
nand U27290 (N_27290,N_27081,N_27072);
nand U27291 (N_27291,N_27017,N_27093);
and U27292 (N_27292,N_27144,N_27041);
nand U27293 (N_27293,N_27016,N_27238);
nor U27294 (N_27294,N_27076,N_27044);
nor U27295 (N_27295,N_27104,N_27201);
nand U27296 (N_27296,N_27219,N_27050);
or U27297 (N_27297,N_27013,N_27124);
xor U27298 (N_27298,N_27142,N_27057);
nor U27299 (N_27299,N_27128,N_27178);
and U27300 (N_27300,N_27003,N_27027);
and U27301 (N_27301,N_27233,N_27203);
xnor U27302 (N_27302,N_27180,N_27249);
xor U27303 (N_27303,N_27040,N_27063);
or U27304 (N_27304,N_27037,N_27022);
nand U27305 (N_27305,N_27095,N_27065);
xor U27306 (N_27306,N_27048,N_27159);
nand U27307 (N_27307,N_27112,N_27196);
nor U27308 (N_27308,N_27192,N_27034);
nand U27309 (N_27309,N_27155,N_27084);
nand U27310 (N_27310,N_27079,N_27000);
xnor U27311 (N_27311,N_27031,N_27047);
nand U27312 (N_27312,N_27078,N_27224);
xor U27313 (N_27313,N_27199,N_27054);
nand U27314 (N_27314,N_27126,N_27151);
xor U27315 (N_27315,N_27173,N_27014);
nor U27316 (N_27316,N_27113,N_27028);
or U27317 (N_27317,N_27023,N_27207);
xor U27318 (N_27318,N_27218,N_27182);
nand U27319 (N_27319,N_27060,N_27001);
or U27320 (N_27320,N_27092,N_27036);
nor U27321 (N_27321,N_27134,N_27139);
nor U27322 (N_27322,N_27188,N_27102);
nor U27323 (N_27323,N_27162,N_27189);
xor U27324 (N_27324,N_27121,N_27046);
and U27325 (N_27325,N_27138,N_27097);
or U27326 (N_27326,N_27222,N_27239);
nand U27327 (N_27327,N_27205,N_27170);
xnor U27328 (N_27328,N_27210,N_27197);
and U27329 (N_27329,N_27165,N_27150);
nor U27330 (N_27330,N_27015,N_27193);
or U27331 (N_27331,N_27005,N_27067);
nor U27332 (N_27332,N_27200,N_27212);
xnor U27333 (N_27333,N_27007,N_27042);
and U27334 (N_27334,N_27055,N_27194);
xnor U27335 (N_27335,N_27131,N_27127);
nand U27336 (N_27336,N_27004,N_27118);
or U27337 (N_27337,N_27008,N_27143);
xor U27338 (N_27338,N_27026,N_27236);
xnor U27339 (N_27339,N_27049,N_27043);
and U27340 (N_27340,N_27110,N_27204);
and U27341 (N_27341,N_27129,N_27107);
xnor U27342 (N_27342,N_27166,N_27147);
nand U27343 (N_27343,N_27038,N_27080);
nand U27344 (N_27344,N_27117,N_27247);
and U27345 (N_27345,N_27053,N_27244);
xor U27346 (N_27346,N_27171,N_27089);
nand U27347 (N_27347,N_27208,N_27100);
and U27348 (N_27348,N_27241,N_27119);
nand U27349 (N_27349,N_27135,N_27086);
xor U27350 (N_27350,N_27052,N_27045);
and U27351 (N_27351,N_27234,N_27237);
or U27352 (N_27352,N_27161,N_27156);
nor U27353 (N_27353,N_27024,N_27242);
nor U27354 (N_27354,N_27164,N_27103);
xor U27355 (N_27355,N_27021,N_27232);
nand U27356 (N_27356,N_27069,N_27019);
nand U27357 (N_27357,N_27064,N_27101);
or U27358 (N_27358,N_27136,N_27114);
xor U27359 (N_27359,N_27075,N_27202);
and U27360 (N_27360,N_27140,N_27011);
nand U27361 (N_27361,N_27187,N_27174);
nor U27362 (N_27362,N_27198,N_27195);
nand U27363 (N_27363,N_27025,N_27083);
xnor U27364 (N_27364,N_27032,N_27106);
and U27365 (N_27365,N_27230,N_27217);
nand U27366 (N_27366,N_27229,N_27012);
or U27367 (N_27367,N_27228,N_27225);
xor U27368 (N_27368,N_27105,N_27172);
nor U27369 (N_27369,N_27061,N_27116);
nor U27370 (N_27370,N_27111,N_27010);
and U27371 (N_27371,N_27177,N_27087);
and U27372 (N_27372,N_27168,N_27130);
nand U27373 (N_27373,N_27018,N_27190);
or U27374 (N_27374,N_27059,N_27070);
and U27375 (N_27375,N_27090,N_27188);
nor U27376 (N_27376,N_27171,N_27023);
nor U27377 (N_27377,N_27068,N_27090);
and U27378 (N_27378,N_27170,N_27194);
or U27379 (N_27379,N_27022,N_27098);
and U27380 (N_27380,N_27139,N_27172);
nor U27381 (N_27381,N_27244,N_27007);
nand U27382 (N_27382,N_27051,N_27143);
nor U27383 (N_27383,N_27234,N_27053);
xnor U27384 (N_27384,N_27190,N_27179);
and U27385 (N_27385,N_27001,N_27164);
or U27386 (N_27386,N_27097,N_27142);
xnor U27387 (N_27387,N_27123,N_27163);
nand U27388 (N_27388,N_27222,N_27136);
or U27389 (N_27389,N_27234,N_27137);
nand U27390 (N_27390,N_27151,N_27088);
or U27391 (N_27391,N_27184,N_27082);
nor U27392 (N_27392,N_27226,N_27108);
or U27393 (N_27393,N_27000,N_27128);
nand U27394 (N_27394,N_27196,N_27043);
and U27395 (N_27395,N_27098,N_27074);
nand U27396 (N_27396,N_27028,N_27178);
nor U27397 (N_27397,N_27211,N_27069);
or U27398 (N_27398,N_27199,N_27148);
and U27399 (N_27399,N_27054,N_27102);
xnor U27400 (N_27400,N_27120,N_27194);
nand U27401 (N_27401,N_27159,N_27165);
xnor U27402 (N_27402,N_27190,N_27181);
xnor U27403 (N_27403,N_27221,N_27164);
xor U27404 (N_27404,N_27038,N_27002);
and U27405 (N_27405,N_27000,N_27097);
nor U27406 (N_27406,N_27221,N_27153);
xor U27407 (N_27407,N_27221,N_27158);
nor U27408 (N_27408,N_27075,N_27050);
and U27409 (N_27409,N_27090,N_27057);
and U27410 (N_27410,N_27034,N_27093);
nor U27411 (N_27411,N_27169,N_27072);
nor U27412 (N_27412,N_27228,N_27047);
or U27413 (N_27413,N_27073,N_27072);
or U27414 (N_27414,N_27139,N_27065);
xnor U27415 (N_27415,N_27150,N_27191);
nor U27416 (N_27416,N_27238,N_27219);
xnor U27417 (N_27417,N_27030,N_27019);
or U27418 (N_27418,N_27078,N_27120);
xor U27419 (N_27419,N_27089,N_27081);
or U27420 (N_27420,N_27244,N_27083);
nand U27421 (N_27421,N_27019,N_27242);
or U27422 (N_27422,N_27068,N_27183);
or U27423 (N_27423,N_27204,N_27082);
nor U27424 (N_27424,N_27239,N_27089);
or U27425 (N_27425,N_27239,N_27067);
nand U27426 (N_27426,N_27104,N_27040);
or U27427 (N_27427,N_27006,N_27080);
xor U27428 (N_27428,N_27020,N_27161);
nor U27429 (N_27429,N_27049,N_27225);
nand U27430 (N_27430,N_27100,N_27107);
and U27431 (N_27431,N_27200,N_27202);
or U27432 (N_27432,N_27080,N_27081);
nand U27433 (N_27433,N_27092,N_27156);
xor U27434 (N_27434,N_27001,N_27208);
and U27435 (N_27435,N_27155,N_27175);
nand U27436 (N_27436,N_27060,N_27036);
xor U27437 (N_27437,N_27101,N_27151);
xor U27438 (N_27438,N_27144,N_27197);
or U27439 (N_27439,N_27150,N_27233);
nor U27440 (N_27440,N_27060,N_27019);
nand U27441 (N_27441,N_27048,N_27201);
nand U27442 (N_27442,N_27094,N_27181);
xor U27443 (N_27443,N_27223,N_27000);
nand U27444 (N_27444,N_27242,N_27087);
or U27445 (N_27445,N_27061,N_27071);
and U27446 (N_27446,N_27102,N_27036);
and U27447 (N_27447,N_27198,N_27007);
xnor U27448 (N_27448,N_27233,N_27174);
or U27449 (N_27449,N_27002,N_27029);
nand U27450 (N_27450,N_27165,N_27155);
and U27451 (N_27451,N_27010,N_27175);
nand U27452 (N_27452,N_27179,N_27210);
nand U27453 (N_27453,N_27018,N_27158);
xnor U27454 (N_27454,N_27120,N_27060);
nand U27455 (N_27455,N_27014,N_27198);
nand U27456 (N_27456,N_27003,N_27245);
nor U27457 (N_27457,N_27090,N_27184);
xnor U27458 (N_27458,N_27026,N_27021);
nand U27459 (N_27459,N_27099,N_27095);
or U27460 (N_27460,N_27028,N_27153);
nor U27461 (N_27461,N_27046,N_27129);
nand U27462 (N_27462,N_27181,N_27238);
and U27463 (N_27463,N_27003,N_27214);
or U27464 (N_27464,N_27188,N_27089);
xnor U27465 (N_27465,N_27178,N_27159);
nor U27466 (N_27466,N_27109,N_27094);
and U27467 (N_27467,N_27020,N_27151);
or U27468 (N_27468,N_27230,N_27005);
nand U27469 (N_27469,N_27054,N_27211);
or U27470 (N_27470,N_27047,N_27009);
xor U27471 (N_27471,N_27117,N_27139);
xnor U27472 (N_27472,N_27247,N_27078);
nor U27473 (N_27473,N_27104,N_27231);
nor U27474 (N_27474,N_27177,N_27007);
nor U27475 (N_27475,N_27068,N_27173);
and U27476 (N_27476,N_27204,N_27069);
or U27477 (N_27477,N_27137,N_27178);
nand U27478 (N_27478,N_27194,N_27053);
and U27479 (N_27479,N_27118,N_27134);
nand U27480 (N_27480,N_27190,N_27111);
nor U27481 (N_27481,N_27104,N_27147);
nand U27482 (N_27482,N_27003,N_27084);
nand U27483 (N_27483,N_27230,N_27090);
xnor U27484 (N_27484,N_27108,N_27010);
or U27485 (N_27485,N_27038,N_27011);
nor U27486 (N_27486,N_27023,N_27066);
or U27487 (N_27487,N_27189,N_27169);
and U27488 (N_27488,N_27168,N_27132);
nand U27489 (N_27489,N_27164,N_27076);
or U27490 (N_27490,N_27078,N_27081);
nor U27491 (N_27491,N_27132,N_27081);
xor U27492 (N_27492,N_27246,N_27212);
nor U27493 (N_27493,N_27130,N_27041);
nor U27494 (N_27494,N_27157,N_27174);
and U27495 (N_27495,N_27126,N_27214);
xor U27496 (N_27496,N_27240,N_27050);
nor U27497 (N_27497,N_27091,N_27075);
xnor U27498 (N_27498,N_27145,N_27121);
nand U27499 (N_27499,N_27089,N_27199);
nand U27500 (N_27500,N_27379,N_27426);
or U27501 (N_27501,N_27497,N_27381);
nand U27502 (N_27502,N_27465,N_27344);
and U27503 (N_27503,N_27419,N_27258);
or U27504 (N_27504,N_27361,N_27444);
xor U27505 (N_27505,N_27469,N_27438);
xor U27506 (N_27506,N_27386,N_27380);
xor U27507 (N_27507,N_27481,N_27406);
nand U27508 (N_27508,N_27459,N_27272);
and U27509 (N_27509,N_27388,N_27410);
nand U27510 (N_27510,N_27395,N_27353);
nand U27511 (N_27511,N_27378,N_27394);
nand U27512 (N_27512,N_27478,N_27273);
or U27513 (N_27513,N_27446,N_27259);
xnor U27514 (N_27514,N_27298,N_27311);
or U27515 (N_27515,N_27295,N_27261);
or U27516 (N_27516,N_27254,N_27448);
nor U27517 (N_27517,N_27329,N_27474);
or U27518 (N_27518,N_27418,N_27431);
nor U27519 (N_27519,N_27270,N_27342);
or U27520 (N_27520,N_27323,N_27284);
xnor U27521 (N_27521,N_27376,N_27333);
nor U27522 (N_27522,N_27411,N_27360);
nand U27523 (N_27523,N_27305,N_27286);
nand U27524 (N_27524,N_27451,N_27463);
xor U27525 (N_27525,N_27391,N_27327);
and U27526 (N_27526,N_27276,N_27464);
nand U27527 (N_27527,N_27348,N_27439);
or U27528 (N_27528,N_27309,N_27257);
nand U27529 (N_27529,N_27456,N_27413);
nand U27530 (N_27530,N_27495,N_27351);
or U27531 (N_27531,N_27384,N_27428);
or U27532 (N_27532,N_27499,N_27310);
xor U27533 (N_27533,N_27279,N_27308);
and U27534 (N_27534,N_27458,N_27441);
or U27535 (N_27535,N_27408,N_27319);
nand U27536 (N_27536,N_27472,N_27390);
or U27537 (N_27537,N_27337,N_27407);
nor U27538 (N_27538,N_27397,N_27462);
and U27539 (N_27539,N_27267,N_27409);
or U27540 (N_27540,N_27252,N_27250);
nor U27541 (N_27541,N_27306,N_27285);
nor U27542 (N_27542,N_27335,N_27322);
nand U27543 (N_27543,N_27328,N_27371);
or U27544 (N_27544,N_27287,N_27265);
xor U27545 (N_27545,N_27320,N_27313);
nand U27546 (N_27546,N_27350,N_27432);
xor U27547 (N_27547,N_27483,N_27400);
xor U27548 (N_27548,N_27479,N_27368);
nor U27549 (N_27549,N_27430,N_27263);
and U27550 (N_27550,N_27314,N_27420);
xor U27551 (N_27551,N_27324,N_27355);
or U27552 (N_27552,N_27294,N_27429);
nand U27553 (N_27553,N_27253,N_27480);
or U27554 (N_27554,N_27365,N_27484);
nor U27555 (N_27555,N_27424,N_27281);
xnor U27556 (N_27556,N_27364,N_27433);
nor U27557 (N_27557,N_27452,N_27399);
and U27558 (N_27558,N_27427,N_27437);
nor U27559 (N_27559,N_27346,N_27312);
or U27560 (N_27560,N_27280,N_27435);
xnor U27561 (N_27561,N_27345,N_27491);
or U27562 (N_27562,N_27343,N_27334);
or U27563 (N_27563,N_27369,N_27292);
or U27564 (N_27564,N_27414,N_27260);
and U27565 (N_27565,N_27385,N_27477);
nor U27566 (N_27566,N_27422,N_27423);
or U27567 (N_27567,N_27339,N_27401);
and U27568 (N_27568,N_27326,N_27358);
xnor U27569 (N_27569,N_27296,N_27289);
nand U27570 (N_27570,N_27347,N_27442);
and U27571 (N_27571,N_27340,N_27268);
and U27572 (N_27572,N_27449,N_27332);
nand U27573 (N_27573,N_27301,N_27293);
and U27574 (N_27574,N_27354,N_27398);
nor U27575 (N_27575,N_27275,N_27375);
and U27576 (N_27576,N_27317,N_27269);
xor U27577 (N_27577,N_27330,N_27392);
and U27578 (N_27578,N_27450,N_27473);
or U27579 (N_27579,N_27352,N_27417);
nand U27580 (N_27580,N_27496,N_27377);
and U27581 (N_27581,N_27366,N_27291);
nor U27582 (N_27582,N_27487,N_27443);
nand U27583 (N_27583,N_27297,N_27359);
and U27584 (N_27584,N_27468,N_27304);
xnor U27585 (N_27585,N_27362,N_27485);
xor U27586 (N_27586,N_27382,N_27374);
xor U27587 (N_27587,N_27445,N_27288);
or U27588 (N_27588,N_27393,N_27436);
xnor U27589 (N_27589,N_27300,N_27338);
nor U27590 (N_27590,N_27266,N_27356);
nand U27591 (N_27591,N_27434,N_27492);
and U27592 (N_27592,N_27299,N_27383);
nand U27593 (N_27593,N_27475,N_27396);
xor U27594 (N_27594,N_27494,N_27262);
and U27595 (N_27595,N_27331,N_27486);
or U27596 (N_27596,N_27303,N_27461);
and U27597 (N_27597,N_27470,N_27453);
or U27598 (N_27598,N_27373,N_27302);
or U27599 (N_27599,N_27325,N_27460);
and U27600 (N_27600,N_27307,N_27349);
nand U27601 (N_27601,N_27488,N_27290);
or U27602 (N_27602,N_27370,N_27278);
nor U27603 (N_27603,N_27387,N_27283);
or U27604 (N_27604,N_27403,N_27415);
or U27605 (N_27605,N_27467,N_27389);
nor U27606 (N_27606,N_27336,N_27471);
and U27607 (N_27607,N_27363,N_27341);
xnor U27608 (N_27608,N_27455,N_27440);
nand U27609 (N_27609,N_27318,N_27476);
nor U27610 (N_27610,N_27490,N_27277);
or U27611 (N_27611,N_27447,N_27498);
nor U27612 (N_27612,N_27404,N_27274);
or U27613 (N_27613,N_27405,N_27315);
xor U27614 (N_27614,N_27316,N_27255);
nor U27615 (N_27615,N_27321,N_27251);
nor U27616 (N_27616,N_27264,N_27493);
nand U27617 (N_27617,N_27357,N_27425);
or U27618 (N_27618,N_27256,N_27416);
and U27619 (N_27619,N_27457,N_27372);
xnor U27620 (N_27620,N_27482,N_27412);
nand U27621 (N_27621,N_27489,N_27282);
nor U27622 (N_27622,N_27402,N_27271);
nand U27623 (N_27623,N_27466,N_27421);
and U27624 (N_27624,N_27367,N_27454);
and U27625 (N_27625,N_27446,N_27491);
or U27626 (N_27626,N_27275,N_27468);
xnor U27627 (N_27627,N_27304,N_27321);
xnor U27628 (N_27628,N_27473,N_27485);
nor U27629 (N_27629,N_27389,N_27336);
xnor U27630 (N_27630,N_27468,N_27349);
and U27631 (N_27631,N_27395,N_27437);
or U27632 (N_27632,N_27270,N_27356);
or U27633 (N_27633,N_27444,N_27476);
xor U27634 (N_27634,N_27420,N_27320);
xor U27635 (N_27635,N_27403,N_27417);
or U27636 (N_27636,N_27262,N_27258);
and U27637 (N_27637,N_27387,N_27408);
or U27638 (N_27638,N_27454,N_27336);
xor U27639 (N_27639,N_27357,N_27460);
or U27640 (N_27640,N_27414,N_27453);
nand U27641 (N_27641,N_27374,N_27355);
nand U27642 (N_27642,N_27399,N_27454);
xor U27643 (N_27643,N_27363,N_27420);
nand U27644 (N_27644,N_27462,N_27428);
nand U27645 (N_27645,N_27478,N_27262);
nor U27646 (N_27646,N_27427,N_27302);
nor U27647 (N_27647,N_27309,N_27382);
nor U27648 (N_27648,N_27396,N_27412);
nor U27649 (N_27649,N_27336,N_27441);
or U27650 (N_27650,N_27445,N_27371);
nor U27651 (N_27651,N_27317,N_27371);
or U27652 (N_27652,N_27337,N_27410);
nand U27653 (N_27653,N_27346,N_27382);
nor U27654 (N_27654,N_27325,N_27359);
xor U27655 (N_27655,N_27442,N_27483);
xnor U27656 (N_27656,N_27309,N_27285);
or U27657 (N_27657,N_27385,N_27379);
nor U27658 (N_27658,N_27262,N_27379);
or U27659 (N_27659,N_27377,N_27286);
or U27660 (N_27660,N_27365,N_27382);
nor U27661 (N_27661,N_27475,N_27439);
nor U27662 (N_27662,N_27258,N_27430);
nand U27663 (N_27663,N_27296,N_27306);
nor U27664 (N_27664,N_27319,N_27460);
nor U27665 (N_27665,N_27480,N_27401);
nor U27666 (N_27666,N_27290,N_27256);
and U27667 (N_27667,N_27349,N_27300);
and U27668 (N_27668,N_27350,N_27482);
xnor U27669 (N_27669,N_27266,N_27456);
nor U27670 (N_27670,N_27305,N_27463);
nand U27671 (N_27671,N_27263,N_27311);
xnor U27672 (N_27672,N_27393,N_27423);
xnor U27673 (N_27673,N_27254,N_27369);
and U27674 (N_27674,N_27472,N_27348);
xor U27675 (N_27675,N_27346,N_27335);
nor U27676 (N_27676,N_27375,N_27364);
nor U27677 (N_27677,N_27250,N_27292);
or U27678 (N_27678,N_27489,N_27465);
xnor U27679 (N_27679,N_27496,N_27341);
xor U27680 (N_27680,N_27484,N_27428);
nor U27681 (N_27681,N_27359,N_27328);
or U27682 (N_27682,N_27469,N_27367);
and U27683 (N_27683,N_27285,N_27261);
nand U27684 (N_27684,N_27445,N_27410);
nand U27685 (N_27685,N_27368,N_27401);
xnor U27686 (N_27686,N_27325,N_27444);
or U27687 (N_27687,N_27287,N_27303);
nand U27688 (N_27688,N_27425,N_27306);
xnor U27689 (N_27689,N_27298,N_27475);
xor U27690 (N_27690,N_27318,N_27265);
nand U27691 (N_27691,N_27397,N_27343);
nor U27692 (N_27692,N_27404,N_27379);
nand U27693 (N_27693,N_27328,N_27257);
xnor U27694 (N_27694,N_27320,N_27370);
nor U27695 (N_27695,N_27251,N_27315);
nand U27696 (N_27696,N_27435,N_27424);
and U27697 (N_27697,N_27292,N_27450);
xor U27698 (N_27698,N_27424,N_27264);
or U27699 (N_27699,N_27447,N_27366);
nor U27700 (N_27700,N_27279,N_27254);
nand U27701 (N_27701,N_27291,N_27262);
nand U27702 (N_27702,N_27350,N_27260);
xnor U27703 (N_27703,N_27389,N_27408);
or U27704 (N_27704,N_27498,N_27395);
xnor U27705 (N_27705,N_27323,N_27421);
and U27706 (N_27706,N_27287,N_27467);
and U27707 (N_27707,N_27361,N_27405);
xnor U27708 (N_27708,N_27450,N_27325);
nor U27709 (N_27709,N_27473,N_27498);
nor U27710 (N_27710,N_27476,N_27415);
nand U27711 (N_27711,N_27275,N_27358);
or U27712 (N_27712,N_27481,N_27464);
xnor U27713 (N_27713,N_27483,N_27333);
and U27714 (N_27714,N_27382,N_27277);
nand U27715 (N_27715,N_27412,N_27418);
and U27716 (N_27716,N_27473,N_27263);
nor U27717 (N_27717,N_27362,N_27447);
nand U27718 (N_27718,N_27251,N_27481);
xnor U27719 (N_27719,N_27450,N_27381);
xnor U27720 (N_27720,N_27292,N_27322);
and U27721 (N_27721,N_27476,N_27252);
nand U27722 (N_27722,N_27343,N_27429);
or U27723 (N_27723,N_27448,N_27426);
and U27724 (N_27724,N_27328,N_27430);
and U27725 (N_27725,N_27393,N_27348);
nor U27726 (N_27726,N_27413,N_27375);
and U27727 (N_27727,N_27367,N_27349);
and U27728 (N_27728,N_27273,N_27267);
or U27729 (N_27729,N_27462,N_27437);
or U27730 (N_27730,N_27417,N_27289);
and U27731 (N_27731,N_27413,N_27497);
xor U27732 (N_27732,N_27381,N_27278);
or U27733 (N_27733,N_27364,N_27478);
nor U27734 (N_27734,N_27263,N_27326);
xor U27735 (N_27735,N_27481,N_27441);
nand U27736 (N_27736,N_27452,N_27392);
or U27737 (N_27737,N_27418,N_27320);
nor U27738 (N_27738,N_27415,N_27401);
and U27739 (N_27739,N_27415,N_27285);
and U27740 (N_27740,N_27298,N_27376);
nor U27741 (N_27741,N_27468,N_27431);
xor U27742 (N_27742,N_27341,N_27284);
or U27743 (N_27743,N_27328,N_27275);
and U27744 (N_27744,N_27279,N_27446);
and U27745 (N_27745,N_27391,N_27305);
nor U27746 (N_27746,N_27442,N_27473);
and U27747 (N_27747,N_27302,N_27457);
and U27748 (N_27748,N_27382,N_27304);
or U27749 (N_27749,N_27379,N_27346);
nor U27750 (N_27750,N_27555,N_27743);
or U27751 (N_27751,N_27615,N_27505);
nor U27752 (N_27752,N_27731,N_27507);
nor U27753 (N_27753,N_27727,N_27626);
nand U27754 (N_27754,N_27700,N_27670);
or U27755 (N_27755,N_27646,N_27519);
nand U27756 (N_27756,N_27728,N_27694);
nor U27757 (N_27757,N_27531,N_27748);
nor U27758 (N_27758,N_27545,N_27581);
nand U27759 (N_27759,N_27656,N_27625);
xnor U27760 (N_27760,N_27638,N_27510);
nor U27761 (N_27761,N_27516,N_27683);
nor U27762 (N_27762,N_27650,N_27739);
or U27763 (N_27763,N_27730,N_27508);
or U27764 (N_27764,N_27639,N_27629);
nand U27765 (N_27765,N_27592,N_27597);
and U27766 (N_27766,N_27643,N_27648);
nor U27767 (N_27767,N_27518,N_27610);
nand U27768 (N_27768,N_27537,N_27575);
xnor U27769 (N_27769,N_27533,N_27618);
xor U27770 (N_27770,N_27630,N_27641);
or U27771 (N_27771,N_27582,N_27675);
xor U27772 (N_27772,N_27556,N_27691);
nand U27773 (N_27773,N_27671,N_27652);
and U27774 (N_27774,N_27554,N_27568);
or U27775 (N_27775,N_27529,N_27723);
nand U27776 (N_27776,N_27546,N_27596);
xor U27777 (N_27777,N_27547,N_27594);
or U27778 (N_27778,N_27621,N_27635);
or U27779 (N_27779,N_27721,N_27669);
nand U27780 (N_27780,N_27521,N_27611);
xnor U27781 (N_27781,N_27720,N_27603);
xnor U27782 (N_27782,N_27551,N_27530);
nor U27783 (N_27783,N_27747,N_27679);
or U27784 (N_27784,N_27542,N_27526);
and U27785 (N_27785,N_27714,N_27502);
and U27786 (N_27786,N_27578,N_27732);
and U27787 (N_27787,N_27711,N_27632);
nand U27788 (N_27788,N_27569,N_27572);
xor U27789 (N_27789,N_27738,N_27657);
nand U27790 (N_27790,N_27525,N_27698);
and U27791 (N_27791,N_27701,N_27544);
and U27792 (N_27792,N_27590,N_27702);
and U27793 (N_27793,N_27746,N_27736);
xor U27794 (N_27794,N_27609,N_27565);
nor U27795 (N_27795,N_27685,N_27665);
nor U27796 (N_27796,N_27563,N_27623);
xor U27797 (N_27797,N_27580,N_27552);
nor U27798 (N_27798,N_27735,N_27674);
nand U27799 (N_27799,N_27586,N_27567);
and U27800 (N_27800,N_27570,N_27587);
and U27801 (N_27801,N_27644,N_27617);
or U27802 (N_27802,N_27523,N_27734);
nand U27803 (N_27803,N_27566,N_27719);
nor U27804 (N_27804,N_27699,N_27733);
and U27805 (N_27805,N_27664,N_27584);
or U27806 (N_27806,N_27655,N_27673);
and U27807 (N_27807,N_27686,N_27672);
nor U27808 (N_27808,N_27651,N_27718);
or U27809 (N_27809,N_27593,N_27560);
nor U27810 (N_27810,N_27501,N_27642);
xnor U27811 (N_27811,N_27515,N_27614);
xnor U27812 (N_27812,N_27684,N_27631);
nand U27813 (N_27813,N_27509,N_27576);
nand U27814 (N_27814,N_27729,N_27599);
or U27815 (N_27815,N_27653,N_27662);
xnor U27816 (N_27816,N_27659,N_27500);
and U27817 (N_27817,N_27561,N_27640);
xor U27818 (N_27818,N_27558,N_27588);
and U27819 (N_27819,N_27663,N_27620);
nand U27820 (N_27820,N_27658,N_27715);
or U27821 (N_27821,N_27713,N_27506);
xnor U27822 (N_27822,N_27619,N_27532);
nor U27823 (N_27823,N_27503,N_27744);
and U27824 (N_27824,N_27712,N_27645);
xor U27825 (N_27825,N_27682,N_27608);
xnor U27826 (N_27826,N_27628,N_27716);
xnor U27827 (N_27827,N_27583,N_27520);
xnor U27828 (N_27828,N_27710,N_27602);
nand U27829 (N_27829,N_27697,N_27688);
or U27830 (N_27830,N_27517,N_27541);
nand U27831 (N_27831,N_27540,N_27722);
nand U27832 (N_27832,N_27564,N_27573);
and U27833 (N_27833,N_27690,N_27591);
or U27834 (N_27834,N_27585,N_27601);
xnor U27835 (N_27835,N_27559,N_27707);
and U27836 (N_27836,N_27613,N_27536);
xnor U27837 (N_27837,N_27616,N_27528);
xnor U27838 (N_27838,N_27637,N_27579);
nor U27839 (N_27839,N_27562,N_27557);
nand U27840 (N_27840,N_27737,N_27577);
or U27841 (N_27841,N_27512,N_27681);
and U27842 (N_27842,N_27548,N_27677);
xor U27843 (N_27843,N_27538,N_27705);
and U27844 (N_27844,N_27667,N_27535);
nor U27845 (N_27845,N_27647,N_27513);
xor U27846 (N_27846,N_27696,N_27726);
nand U27847 (N_27847,N_27724,N_27676);
and U27848 (N_27848,N_27571,N_27742);
xor U27849 (N_27849,N_27745,N_27511);
nor U27850 (N_27850,N_27600,N_27704);
xor U27851 (N_27851,N_27607,N_27689);
nor U27852 (N_27852,N_27514,N_27649);
and U27853 (N_27853,N_27539,N_27589);
and U27854 (N_27854,N_27695,N_27543);
nor U27855 (N_27855,N_27678,N_27749);
and U27856 (N_27856,N_27522,N_27574);
or U27857 (N_27857,N_27654,N_27666);
and U27858 (N_27858,N_27660,N_27741);
nor U27859 (N_27859,N_27687,N_27680);
xor U27860 (N_27860,N_27598,N_27668);
xor U27861 (N_27861,N_27636,N_27622);
nor U27862 (N_27862,N_27604,N_27706);
or U27863 (N_27863,N_27703,N_27549);
nand U27864 (N_27864,N_27627,N_27504);
or U27865 (N_27865,N_27605,N_27553);
and U27866 (N_27866,N_27725,N_27534);
and U27867 (N_27867,N_27524,N_27740);
nor U27868 (N_27868,N_27661,N_27692);
and U27869 (N_27869,N_27624,N_27709);
xnor U27870 (N_27870,N_27595,N_27634);
and U27871 (N_27871,N_27606,N_27717);
or U27872 (N_27872,N_27633,N_27708);
or U27873 (N_27873,N_27550,N_27527);
and U27874 (N_27874,N_27693,N_27612);
nand U27875 (N_27875,N_27612,N_27621);
or U27876 (N_27876,N_27653,N_27634);
and U27877 (N_27877,N_27603,N_27606);
xor U27878 (N_27878,N_27642,N_27553);
and U27879 (N_27879,N_27677,N_27602);
and U27880 (N_27880,N_27684,N_27653);
xor U27881 (N_27881,N_27747,N_27654);
xor U27882 (N_27882,N_27596,N_27698);
and U27883 (N_27883,N_27545,N_27518);
nand U27884 (N_27884,N_27625,N_27592);
xnor U27885 (N_27885,N_27637,N_27680);
xor U27886 (N_27886,N_27506,N_27517);
nand U27887 (N_27887,N_27698,N_27567);
xor U27888 (N_27888,N_27612,N_27601);
and U27889 (N_27889,N_27504,N_27713);
nand U27890 (N_27890,N_27525,N_27535);
and U27891 (N_27891,N_27719,N_27707);
xor U27892 (N_27892,N_27542,N_27681);
or U27893 (N_27893,N_27640,N_27702);
and U27894 (N_27894,N_27748,N_27686);
and U27895 (N_27895,N_27674,N_27628);
nor U27896 (N_27896,N_27688,N_27617);
nor U27897 (N_27897,N_27515,N_27619);
or U27898 (N_27898,N_27500,N_27559);
or U27899 (N_27899,N_27716,N_27671);
nor U27900 (N_27900,N_27695,N_27562);
or U27901 (N_27901,N_27613,N_27680);
xnor U27902 (N_27902,N_27629,N_27748);
nor U27903 (N_27903,N_27707,N_27677);
and U27904 (N_27904,N_27554,N_27503);
nor U27905 (N_27905,N_27532,N_27656);
and U27906 (N_27906,N_27634,N_27622);
and U27907 (N_27907,N_27721,N_27741);
and U27908 (N_27908,N_27683,N_27655);
nand U27909 (N_27909,N_27641,N_27616);
nor U27910 (N_27910,N_27733,N_27628);
or U27911 (N_27911,N_27571,N_27633);
nand U27912 (N_27912,N_27732,N_27575);
and U27913 (N_27913,N_27608,N_27743);
and U27914 (N_27914,N_27567,N_27509);
nand U27915 (N_27915,N_27691,N_27673);
xor U27916 (N_27916,N_27671,N_27656);
or U27917 (N_27917,N_27535,N_27512);
or U27918 (N_27918,N_27558,N_27601);
and U27919 (N_27919,N_27748,N_27666);
xor U27920 (N_27920,N_27590,N_27746);
or U27921 (N_27921,N_27728,N_27652);
nand U27922 (N_27922,N_27719,N_27745);
and U27923 (N_27923,N_27512,N_27589);
nand U27924 (N_27924,N_27522,N_27539);
nor U27925 (N_27925,N_27674,N_27640);
xnor U27926 (N_27926,N_27748,N_27506);
xor U27927 (N_27927,N_27563,N_27685);
or U27928 (N_27928,N_27714,N_27501);
xor U27929 (N_27929,N_27583,N_27579);
or U27930 (N_27930,N_27584,N_27504);
nand U27931 (N_27931,N_27661,N_27594);
xnor U27932 (N_27932,N_27555,N_27585);
and U27933 (N_27933,N_27691,N_27694);
or U27934 (N_27934,N_27730,N_27542);
and U27935 (N_27935,N_27566,N_27588);
nor U27936 (N_27936,N_27502,N_27737);
nor U27937 (N_27937,N_27729,N_27601);
xnor U27938 (N_27938,N_27512,N_27504);
nor U27939 (N_27939,N_27746,N_27518);
xnor U27940 (N_27940,N_27620,N_27740);
nand U27941 (N_27941,N_27702,N_27611);
or U27942 (N_27942,N_27706,N_27522);
xnor U27943 (N_27943,N_27715,N_27575);
xnor U27944 (N_27944,N_27655,N_27525);
and U27945 (N_27945,N_27500,N_27605);
nor U27946 (N_27946,N_27722,N_27666);
xnor U27947 (N_27947,N_27517,N_27663);
nand U27948 (N_27948,N_27640,N_27649);
and U27949 (N_27949,N_27575,N_27620);
and U27950 (N_27950,N_27556,N_27531);
nand U27951 (N_27951,N_27691,N_27619);
and U27952 (N_27952,N_27682,N_27746);
and U27953 (N_27953,N_27556,N_27745);
nor U27954 (N_27954,N_27553,N_27634);
and U27955 (N_27955,N_27682,N_27662);
or U27956 (N_27956,N_27600,N_27739);
nor U27957 (N_27957,N_27652,N_27680);
xor U27958 (N_27958,N_27729,N_27695);
and U27959 (N_27959,N_27542,N_27622);
nor U27960 (N_27960,N_27518,N_27573);
xor U27961 (N_27961,N_27586,N_27528);
nor U27962 (N_27962,N_27657,N_27501);
or U27963 (N_27963,N_27688,N_27730);
or U27964 (N_27964,N_27690,N_27703);
xor U27965 (N_27965,N_27646,N_27625);
xor U27966 (N_27966,N_27539,N_27676);
xor U27967 (N_27967,N_27697,N_27648);
or U27968 (N_27968,N_27683,N_27502);
xnor U27969 (N_27969,N_27728,N_27703);
or U27970 (N_27970,N_27524,N_27748);
or U27971 (N_27971,N_27718,N_27557);
or U27972 (N_27972,N_27622,N_27556);
and U27973 (N_27973,N_27645,N_27594);
nand U27974 (N_27974,N_27658,N_27627);
xor U27975 (N_27975,N_27565,N_27707);
or U27976 (N_27976,N_27733,N_27706);
or U27977 (N_27977,N_27603,N_27698);
or U27978 (N_27978,N_27716,N_27516);
xnor U27979 (N_27979,N_27694,N_27714);
nor U27980 (N_27980,N_27654,N_27737);
nand U27981 (N_27981,N_27616,N_27620);
xor U27982 (N_27982,N_27550,N_27706);
nand U27983 (N_27983,N_27729,N_27528);
and U27984 (N_27984,N_27738,N_27685);
nor U27985 (N_27985,N_27661,N_27664);
and U27986 (N_27986,N_27547,N_27622);
and U27987 (N_27987,N_27670,N_27676);
or U27988 (N_27988,N_27732,N_27664);
or U27989 (N_27989,N_27507,N_27553);
or U27990 (N_27990,N_27724,N_27533);
or U27991 (N_27991,N_27692,N_27567);
and U27992 (N_27992,N_27607,N_27604);
or U27993 (N_27993,N_27512,N_27713);
nor U27994 (N_27994,N_27625,N_27684);
nor U27995 (N_27995,N_27696,N_27697);
and U27996 (N_27996,N_27744,N_27708);
xor U27997 (N_27997,N_27548,N_27595);
nor U27998 (N_27998,N_27733,N_27615);
nand U27999 (N_27999,N_27525,N_27508);
and U28000 (N_28000,N_27908,N_27833);
and U28001 (N_28001,N_27941,N_27946);
and U28002 (N_28002,N_27846,N_27944);
nand U28003 (N_28003,N_27774,N_27884);
or U28004 (N_28004,N_27843,N_27834);
nand U28005 (N_28005,N_27878,N_27874);
xor U28006 (N_28006,N_27877,N_27916);
nand U28007 (N_28007,N_27760,N_27807);
nor U28008 (N_28008,N_27893,N_27872);
xnor U28009 (N_28009,N_27912,N_27771);
xor U28010 (N_28010,N_27921,N_27915);
nand U28011 (N_28011,N_27759,N_27993);
xnor U28012 (N_28012,N_27920,N_27959);
nand U28013 (N_28013,N_27974,N_27952);
or U28014 (N_28014,N_27802,N_27769);
nor U28015 (N_28015,N_27987,N_27927);
and U28016 (N_28016,N_27899,N_27831);
and U28017 (N_28017,N_27910,N_27785);
nand U28018 (N_28018,N_27782,N_27888);
or U28019 (N_28019,N_27783,N_27863);
or U28020 (N_28020,N_27776,N_27875);
and U28021 (N_28021,N_27837,N_27985);
xnor U28022 (N_28022,N_27918,N_27906);
and U28023 (N_28023,N_27857,N_27964);
xor U28024 (N_28024,N_27886,N_27935);
xnor U28025 (N_28025,N_27975,N_27994);
or U28026 (N_28026,N_27767,N_27779);
or U28027 (N_28027,N_27758,N_27813);
and U28028 (N_28028,N_27913,N_27992);
or U28029 (N_28029,N_27945,N_27977);
xor U28030 (N_28030,N_27953,N_27887);
xnor U28031 (N_28031,N_27838,N_27812);
nor U28032 (N_28032,N_27811,N_27864);
or U28033 (N_28033,N_27961,N_27972);
and U28034 (N_28034,N_27907,N_27911);
nor U28035 (N_28035,N_27784,N_27998);
xor U28036 (N_28036,N_27789,N_27896);
nor U28037 (N_28037,N_27967,N_27809);
xor U28038 (N_28038,N_27826,N_27989);
nand U28039 (N_28039,N_27932,N_27971);
and U28040 (N_28040,N_27850,N_27873);
or U28041 (N_28041,N_27750,N_27866);
and U28042 (N_28042,N_27969,N_27777);
nor U28043 (N_28043,N_27781,N_27855);
nor U28044 (N_28044,N_27995,N_27889);
xor U28045 (N_28045,N_27894,N_27824);
nor U28046 (N_28046,N_27938,N_27775);
nor U28047 (N_28047,N_27757,N_27876);
nor U28048 (N_28048,N_27954,N_27835);
nor U28049 (N_28049,N_27870,N_27885);
and U28050 (N_28050,N_27847,N_27751);
nor U28051 (N_28051,N_27981,N_27839);
or U28052 (N_28052,N_27796,N_27902);
nand U28053 (N_28053,N_27780,N_27792);
nor U28054 (N_28054,N_27900,N_27936);
xnor U28055 (N_28055,N_27787,N_27799);
nand U28056 (N_28056,N_27763,N_27949);
and U28057 (N_28057,N_27815,N_27845);
nand U28058 (N_28058,N_27805,N_27940);
and U28059 (N_28059,N_27798,N_27970);
or U28060 (N_28060,N_27860,N_27820);
nor U28061 (N_28061,N_27895,N_27923);
xor U28062 (N_28062,N_27755,N_27773);
or U28063 (N_28063,N_27897,N_27862);
nand U28064 (N_28064,N_27853,N_27948);
nand U28065 (N_28065,N_27823,N_27973);
nand U28066 (N_28066,N_27890,N_27778);
and U28067 (N_28067,N_27841,N_27849);
nand U28068 (N_28068,N_27898,N_27976);
and U28069 (N_28069,N_27880,N_27955);
and U28070 (N_28070,N_27762,N_27858);
nor U28071 (N_28071,N_27934,N_27868);
nor U28072 (N_28072,N_27914,N_27978);
or U28073 (N_28073,N_27871,N_27883);
and U28074 (N_28074,N_27904,N_27930);
nor U28075 (N_28075,N_27806,N_27905);
or U28076 (N_28076,N_27800,N_27752);
and U28077 (N_28077,N_27957,N_27814);
xnor U28078 (N_28078,N_27892,N_27988);
nor U28079 (N_28079,N_27869,N_27919);
and U28080 (N_28080,N_27786,N_27772);
or U28081 (N_28081,N_27943,N_27803);
and U28082 (N_28082,N_27965,N_27817);
or U28083 (N_28083,N_27810,N_27801);
nand U28084 (N_28084,N_27951,N_27765);
nand U28085 (N_28085,N_27818,N_27939);
xnor U28086 (N_28086,N_27891,N_27832);
nor U28087 (N_28087,N_27984,N_27881);
and U28088 (N_28088,N_27848,N_27980);
nor U28089 (N_28089,N_27983,N_27753);
and U28090 (N_28090,N_27942,N_27958);
or U28091 (N_28091,N_27804,N_27851);
xnor U28092 (N_28092,N_27861,N_27962);
nand U28093 (N_28093,N_27822,N_27859);
xnor U28094 (N_28094,N_27950,N_27986);
nand U28095 (N_28095,N_27790,N_27795);
nor U28096 (N_28096,N_27829,N_27917);
nor U28097 (N_28097,N_27909,N_27996);
and U28098 (N_28098,N_27768,N_27856);
nor U28099 (N_28099,N_27793,N_27836);
nor U28100 (N_28100,N_27852,N_27922);
xor U28101 (N_28101,N_27766,N_27937);
nor U28102 (N_28102,N_27791,N_27867);
or U28103 (N_28103,N_27854,N_27788);
xnor U28104 (N_28104,N_27821,N_27956);
nor U28105 (N_28105,N_27928,N_27991);
and U28106 (N_28106,N_27840,N_27999);
nor U28107 (N_28107,N_27960,N_27865);
nor U28108 (N_28108,N_27901,N_27797);
and U28109 (N_28109,N_27816,N_27844);
xor U28110 (N_28110,N_27842,N_27770);
nor U28111 (N_28111,N_27968,N_27879);
nand U28112 (N_28112,N_27828,N_27990);
and U28113 (N_28113,N_27979,N_27947);
and U28114 (N_28114,N_27756,N_27933);
nand U28115 (N_28115,N_27761,N_27929);
or U28116 (N_28116,N_27794,N_27966);
xor U28117 (N_28117,N_27830,N_27754);
nand U28118 (N_28118,N_27925,N_27825);
or U28119 (N_28119,N_27808,N_27882);
nor U28120 (N_28120,N_27931,N_27819);
nor U28121 (N_28121,N_27926,N_27764);
nor U28122 (N_28122,N_27924,N_27827);
and U28123 (N_28123,N_27997,N_27903);
or U28124 (N_28124,N_27963,N_27982);
xnor U28125 (N_28125,N_27791,N_27876);
nor U28126 (N_28126,N_27946,N_27763);
or U28127 (N_28127,N_27990,N_27842);
and U28128 (N_28128,N_27920,N_27869);
xnor U28129 (N_28129,N_27872,N_27868);
xor U28130 (N_28130,N_27801,N_27975);
nand U28131 (N_28131,N_27848,N_27982);
nor U28132 (N_28132,N_27887,N_27807);
nand U28133 (N_28133,N_27832,N_27875);
or U28134 (N_28134,N_27807,N_27842);
nand U28135 (N_28135,N_27846,N_27766);
and U28136 (N_28136,N_27854,N_27752);
or U28137 (N_28137,N_27832,N_27955);
and U28138 (N_28138,N_27888,N_27957);
nor U28139 (N_28139,N_27942,N_27865);
nor U28140 (N_28140,N_27806,N_27814);
nor U28141 (N_28141,N_27980,N_27912);
or U28142 (N_28142,N_27809,N_27916);
xor U28143 (N_28143,N_27883,N_27939);
and U28144 (N_28144,N_27882,N_27858);
and U28145 (N_28145,N_27952,N_27939);
xor U28146 (N_28146,N_27929,N_27908);
and U28147 (N_28147,N_27802,N_27945);
and U28148 (N_28148,N_27996,N_27851);
nor U28149 (N_28149,N_27779,N_27837);
or U28150 (N_28150,N_27909,N_27858);
nand U28151 (N_28151,N_27762,N_27889);
nand U28152 (N_28152,N_27846,N_27824);
and U28153 (N_28153,N_27908,N_27912);
and U28154 (N_28154,N_27895,N_27930);
or U28155 (N_28155,N_27871,N_27823);
nor U28156 (N_28156,N_27972,N_27862);
nand U28157 (N_28157,N_27891,N_27971);
and U28158 (N_28158,N_27777,N_27796);
nand U28159 (N_28159,N_27882,N_27985);
xor U28160 (N_28160,N_27989,N_27972);
nor U28161 (N_28161,N_27753,N_27784);
nor U28162 (N_28162,N_27890,N_27845);
or U28163 (N_28163,N_27813,N_27963);
xor U28164 (N_28164,N_27856,N_27953);
and U28165 (N_28165,N_27758,N_27868);
nand U28166 (N_28166,N_27899,N_27872);
xor U28167 (N_28167,N_27839,N_27898);
xnor U28168 (N_28168,N_27809,N_27910);
nand U28169 (N_28169,N_27812,N_27882);
xnor U28170 (N_28170,N_27941,N_27914);
nand U28171 (N_28171,N_27900,N_27985);
nand U28172 (N_28172,N_27893,N_27987);
and U28173 (N_28173,N_27790,N_27912);
xnor U28174 (N_28174,N_27954,N_27949);
nor U28175 (N_28175,N_27883,N_27866);
xnor U28176 (N_28176,N_27856,N_27964);
and U28177 (N_28177,N_27827,N_27769);
and U28178 (N_28178,N_27893,N_27935);
xor U28179 (N_28179,N_27970,N_27850);
or U28180 (N_28180,N_27871,N_27894);
or U28181 (N_28181,N_27895,N_27776);
nand U28182 (N_28182,N_27756,N_27786);
nand U28183 (N_28183,N_27849,N_27988);
or U28184 (N_28184,N_27870,N_27774);
xor U28185 (N_28185,N_27784,N_27942);
and U28186 (N_28186,N_27945,N_27832);
and U28187 (N_28187,N_27835,N_27809);
nor U28188 (N_28188,N_27878,N_27792);
or U28189 (N_28189,N_27913,N_27841);
or U28190 (N_28190,N_27754,N_27838);
and U28191 (N_28191,N_27834,N_27969);
xnor U28192 (N_28192,N_27893,N_27879);
xnor U28193 (N_28193,N_27776,N_27750);
or U28194 (N_28194,N_27853,N_27777);
and U28195 (N_28195,N_27995,N_27763);
xnor U28196 (N_28196,N_27781,N_27801);
and U28197 (N_28197,N_27969,N_27862);
xnor U28198 (N_28198,N_27866,N_27820);
nor U28199 (N_28199,N_27980,N_27903);
and U28200 (N_28200,N_27986,N_27785);
and U28201 (N_28201,N_27917,N_27925);
xor U28202 (N_28202,N_27914,N_27784);
nor U28203 (N_28203,N_27775,N_27807);
nor U28204 (N_28204,N_27755,N_27870);
and U28205 (N_28205,N_27907,N_27904);
xnor U28206 (N_28206,N_27880,N_27913);
and U28207 (N_28207,N_27841,N_27811);
xnor U28208 (N_28208,N_27964,N_27956);
xnor U28209 (N_28209,N_27945,N_27987);
nor U28210 (N_28210,N_27887,N_27942);
nand U28211 (N_28211,N_27927,N_27770);
nand U28212 (N_28212,N_27930,N_27753);
or U28213 (N_28213,N_27997,N_27821);
xnor U28214 (N_28214,N_27812,N_27750);
nand U28215 (N_28215,N_27822,N_27758);
nand U28216 (N_28216,N_27811,N_27819);
nor U28217 (N_28217,N_27912,N_27902);
nand U28218 (N_28218,N_27947,N_27901);
xor U28219 (N_28219,N_27769,N_27897);
or U28220 (N_28220,N_27971,N_27984);
xor U28221 (N_28221,N_27762,N_27771);
nand U28222 (N_28222,N_27986,N_27764);
xor U28223 (N_28223,N_27835,N_27932);
or U28224 (N_28224,N_27912,N_27964);
and U28225 (N_28225,N_27921,N_27987);
or U28226 (N_28226,N_27953,N_27892);
xor U28227 (N_28227,N_27988,N_27960);
and U28228 (N_28228,N_27827,N_27851);
or U28229 (N_28229,N_27987,N_27907);
xnor U28230 (N_28230,N_27962,N_27786);
xnor U28231 (N_28231,N_27777,N_27752);
xor U28232 (N_28232,N_27769,N_27839);
nand U28233 (N_28233,N_27814,N_27883);
nand U28234 (N_28234,N_27928,N_27963);
nor U28235 (N_28235,N_27862,N_27778);
or U28236 (N_28236,N_27951,N_27893);
or U28237 (N_28237,N_27844,N_27808);
xor U28238 (N_28238,N_27756,N_27845);
xnor U28239 (N_28239,N_27910,N_27803);
nor U28240 (N_28240,N_27796,N_27992);
or U28241 (N_28241,N_27915,N_27876);
nand U28242 (N_28242,N_27888,N_27795);
nand U28243 (N_28243,N_27855,N_27861);
xnor U28244 (N_28244,N_27842,N_27929);
nand U28245 (N_28245,N_27906,N_27908);
nor U28246 (N_28246,N_27922,N_27941);
and U28247 (N_28247,N_27785,N_27771);
nand U28248 (N_28248,N_27883,N_27874);
nor U28249 (N_28249,N_27991,N_27923);
and U28250 (N_28250,N_28057,N_28146);
xor U28251 (N_28251,N_28027,N_28088);
and U28252 (N_28252,N_28169,N_28185);
xor U28253 (N_28253,N_28175,N_28229);
xor U28254 (N_28254,N_28133,N_28147);
nand U28255 (N_28255,N_28194,N_28078);
xor U28256 (N_28256,N_28203,N_28040);
and U28257 (N_28257,N_28236,N_28199);
nand U28258 (N_28258,N_28020,N_28011);
and U28259 (N_28259,N_28012,N_28024);
nor U28260 (N_28260,N_28039,N_28149);
xnor U28261 (N_28261,N_28121,N_28184);
and U28262 (N_28262,N_28033,N_28224);
xnor U28263 (N_28263,N_28059,N_28195);
nand U28264 (N_28264,N_28163,N_28161);
nor U28265 (N_28265,N_28207,N_28227);
and U28266 (N_28266,N_28035,N_28122);
xor U28267 (N_28267,N_28116,N_28215);
xor U28268 (N_28268,N_28134,N_28052);
xnor U28269 (N_28269,N_28109,N_28232);
or U28270 (N_28270,N_28148,N_28120);
and U28271 (N_28271,N_28096,N_28031);
and U28272 (N_28272,N_28063,N_28070);
xnor U28273 (N_28273,N_28093,N_28200);
or U28274 (N_28274,N_28102,N_28136);
nand U28275 (N_28275,N_28076,N_28189);
xor U28276 (N_28276,N_28151,N_28142);
or U28277 (N_28277,N_28104,N_28126);
or U28278 (N_28278,N_28029,N_28089);
nand U28279 (N_28279,N_28044,N_28087);
nor U28280 (N_28280,N_28009,N_28036);
and U28281 (N_28281,N_28001,N_28099);
nand U28282 (N_28282,N_28108,N_28066);
xor U28283 (N_28283,N_28005,N_28174);
xnor U28284 (N_28284,N_28113,N_28038);
nand U28285 (N_28285,N_28157,N_28034);
or U28286 (N_28286,N_28019,N_28239);
nor U28287 (N_28287,N_28056,N_28115);
nand U28288 (N_28288,N_28172,N_28166);
or U28289 (N_28289,N_28135,N_28238);
xor U28290 (N_28290,N_28119,N_28190);
nor U28291 (N_28291,N_28138,N_28107);
nor U28292 (N_28292,N_28140,N_28068);
nand U28293 (N_28293,N_28193,N_28128);
or U28294 (N_28294,N_28018,N_28145);
or U28295 (N_28295,N_28055,N_28106);
or U28296 (N_28296,N_28230,N_28085);
and U28297 (N_28297,N_28141,N_28111);
nand U28298 (N_28298,N_28181,N_28216);
nand U28299 (N_28299,N_28051,N_28178);
and U28300 (N_28300,N_28082,N_28065);
nand U28301 (N_28301,N_28205,N_28002);
or U28302 (N_28302,N_28220,N_28118);
and U28303 (N_28303,N_28062,N_28092);
or U28304 (N_28304,N_28127,N_28170);
nand U28305 (N_28305,N_28043,N_28084);
xor U28306 (N_28306,N_28014,N_28124);
or U28307 (N_28307,N_28155,N_28053);
and U28308 (N_28308,N_28162,N_28240);
or U28309 (N_28309,N_28214,N_28192);
nand U28310 (N_28310,N_28110,N_28191);
nor U28311 (N_28311,N_28248,N_28032);
nor U28312 (N_28312,N_28047,N_28112);
or U28313 (N_28313,N_28208,N_28160);
xnor U28314 (N_28314,N_28049,N_28177);
xnor U28315 (N_28315,N_28245,N_28086);
nor U28316 (N_28316,N_28223,N_28152);
or U28317 (N_28317,N_28182,N_28101);
xor U28318 (N_28318,N_28204,N_28218);
nand U28319 (N_28319,N_28064,N_28130);
and U28320 (N_28320,N_28060,N_28016);
or U28321 (N_28321,N_28156,N_28197);
xnor U28322 (N_28322,N_28054,N_28237);
or U28323 (N_28323,N_28188,N_28150);
nor U28324 (N_28324,N_28231,N_28090);
xnor U28325 (N_28325,N_28129,N_28061);
or U28326 (N_28326,N_28132,N_28241);
nor U28327 (N_28327,N_28168,N_28069);
nor U28328 (N_28328,N_28105,N_28021);
xor U28329 (N_28329,N_28023,N_28222);
xor U28330 (N_28330,N_28081,N_28030);
or U28331 (N_28331,N_28212,N_28103);
nor U28332 (N_28332,N_28213,N_28198);
xor U28333 (N_28333,N_28028,N_28117);
xor U28334 (N_28334,N_28221,N_28098);
nand U28335 (N_28335,N_28042,N_28073);
and U28336 (N_28336,N_28226,N_28210);
or U28337 (N_28337,N_28097,N_28167);
or U28338 (N_28338,N_28080,N_28143);
nor U28339 (N_28339,N_28046,N_28094);
nand U28340 (N_28340,N_28144,N_28050);
and U28341 (N_28341,N_28211,N_28074);
and U28342 (N_28342,N_28164,N_28008);
xor U28343 (N_28343,N_28183,N_28077);
and U28344 (N_28344,N_28048,N_28247);
nor U28345 (N_28345,N_28131,N_28010);
nand U28346 (N_28346,N_28246,N_28176);
nor U28347 (N_28347,N_28075,N_28139);
xnor U28348 (N_28348,N_28067,N_28100);
or U28349 (N_28349,N_28006,N_28003);
nand U28350 (N_28350,N_28114,N_28015);
xnor U28351 (N_28351,N_28013,N_28079);
and U28352 (N_28352,N_28196,N_28091);
nand U28353 (N_28353,N_28137,N_28180);
or U28354 (N_28354,N_28233,N_28217);
and U28355 (N_28355,N_28201,N_28000);
nor U28356 (N_28356,N_28154,N_28072);
nor U28357 (N_28357,N_28158,N_28249);
and U28358 (N_28358,N_28045,N_28083);
xor U28359 (N_28359,N_28206,N_28025);
and U28360 (N_28360,N_28007,N_28209);
nor U28361 (N_28361,N_28219,N_28123);
or U28362 (N_28362,N_28125,N_28244);
and U28363 (N_28363,N_28242,N_28234);
and U28364 (N_28364,N_28004,N_28228);
nand U28365 (N_28365,N_28017,N_28026);
xnor U28366 (N_28366,N_28041,N_28202);
nand U28367 (N_28367,N_28243,N_28095);
and U28368 (N_28368,N_28165,N_28022);
nand U28369 (N_28369,N_28187,N_28071);
nand U28370 (N_28370,N_28058,N_28153);
nand U28371 (N_28371,N_28159,N_28173);
nor U28372 (N_28372,N_28225,N_28171);
xnor U28373 (N_28373,N_28037,N_28179);
nor U28374 (N_28374,N_28186,N_28235);
nor U28375 (N_28375,N_28189,N_28060);
or U28376 (N_28376,N_28058,N_28137);
xor U28377 (N_28377,N_28184,N_28053);
or U28378 (N_28378,N_28120,N_28145);
xnor U28379 (N_28379,N_28109,N_28056);
xnor U28380 (N_28380,N_28016,N_28211);
nand U28381 (N_28381,N_28099,N_28167);
nor U28382 (N_28382,N_28112,N_28009);
nor U28383 (N_28383,N_28188,N_28062);
nand U28384 (N_28384,N_28168,N_28210);
xnor U28385 (N_28385,N_28085,N_28059);
or U28386 (N_28386,N_28025,N_28185);
nand U28387 (N_28387,N_28088,N_28072);
xnor U28388 (N_28388,N_28223,N_28126);
and U28389 (N_28389,N_28148,N_28052);
nor U28390 (N_28390,N_28059,N_28094);
and U28391 (N_28391,N_28131,N_28108);
and U28392 (N_28392,N_28247,N_28036);
or U28393 (N_28393,N_28007,N_28139);
nor U28394 (N_28394,N_28010,N_28030);
nor U28395 (N_28395,N_28172,N_28181);
nand U28396 (N_28396,N_28091,N_28133);
nand U28397 (N_28397,N_28200,N_28049);
or U28398 (N_28398,N_28089,N_28098);
or U28399 (N_28399,N_28159,N_28100);
nor U28400 (N_28400,N_28198,N_28224);
or U28401 (N_28401,N_28232,N_28172);
xor U28402 (N_28402,N_28243,N_28055);
nor U28403 (N_28403,N_28079,N_28140);
or U28404 (N_28404,N_28036,N_28225);
nor U28405 (N_28405,N_28104,N_28224);
nor U28406 (N_28406,N_28085,N_28134);
xor U28407 (N_28407,N_28173,N_28022);
nand U28408 (N_28408,N_28039,N_28130);
or U28409 (N_28409,N_28032,N_28104);
xor U28410 (N_28410,N_28141,N_28057);
xor U28411 (N_28411,N_28200,N_28135);
or U28412 (N_28412,N_28032,N_28222);
nor U28413 (N_28413,N_28244,N_28231);
or U28414 (N_28414,N_28161,N_28180);
and U28415 (N_28415,N_28233,N_28231);
and U28416 (N_28416,N_28139,N_28064);
nand U28417 (N_28417,N_28222,N_28219);
nand U28418 (N_28418,N_28019,N_28146);
nand U28419 (N_28419,N_28158,N_28221);
nand U28420 (N_28420,N_28198,N_28080);
nand U28421 (N_28421,N_28247,N_28079);
nand U28422 (N_28422,N_28001,N_28206);
xnor U28423 (N_28423,N_28115,N_28231);
nand U28424 (N_28424,N_28240,N_28001);
and U28425 (N_28425,N_28146,N_28212);
and U28426 (N_28426,N_28053,N_28084);
nor U28427 (N_28427,N_28055,N_28238);
xnor U28428 (N_28428,N_28099,N_28053);
nand U28429 (N_28429,N_28011,N_28031);
nand U28430 (N_28430,N_28182,N_28175);
or U28431 (N_28431,N_28056,N_28142);
xnor U28432 (N_28432,N_28242,N_28239);
or U28433 (N_28433,N_28248,N_28049);
or U28434 (N_28434,N_28102,N_28157);
or U28435 (N_28435,N_28229,N_28231);
nand U28436 (N_28436,N_28084,N_28029);
xnor U28437 (N_28437,N_28039,N_28146);
xnor U28438 (N_28438,N_28236,N_28218);
or U28439 (N_28439,N_28203,N_28051);
nor U28440 (N_28440,N_28190,N_28084);
and U28441 (N_28441,N_28045,N_28129);
or U28442 (N_28442,N_28217,N_28184);
xor U28443 (N_28443,N_28144,N_28136);
nand U28444 (N_28444,N_28001,N_28070);
nand U28445 (N_28445,N_28017,N_28040);
nor U28446 (N_28446,N_28184,N_28173);
nand U28447 (N_28447,N_28085,N_28171);
nand U28448 (N_28448,N_28034,N_28229);
nand U28449 (N_28449,N_28103,N_28241);
or U28450 (N_28450,N_28178,N_28228);
or U28451 (N_28451,N_28141,N_28145);
xor U28452 (N_28452,N_28053,N_28017);
and U28453 (N_28453,N_28155,N_28106);
nor U28454 (N_28454,N_28002,N_28023);
nor U28455 (N_28455,N_28120,N_28192);
nand U28456 (N_28456,N_28230,N_28089);
nor U28457 (N_28457,N_28067,N_28183);
nand U28458 (N_28458,N_28087,N_28050);
nor U28459 (N_28459,N_28047,N_28146);
and U28460 (N_28460,N_28133,N_28218);
nor U28461 (N_28461,N_28034,N_28119);
and U28462 (N_28462,N_28086,N_28088);
nand U28463 (N_28463,N_28112,N_28033);
or U28464 (N_28464,N_28232,N_28040);
xor U28465 (N_28465,N_28079,N_28011);
xor U28466 (N_28466,N_28032,N_28100);
or U28467 (N_28467,N_28172,N_28202);
xnor U28468 (N_28468,N_28149,N_28100);
xor U28469 (N_28469,N_28209,N_28016);
nand U28470 (N_28470,N_28239,N_28108);
nand U28471 (N_28471,N_28229,N_28027);
xnor U28472 (N_28472,N_28084,N_28222);
nand U28473 (N_28473,N_28243,N_28227);
nand U28474 (N_28474,N_28003,N_28196);
nand U28475 (N_28475,N_28126,N_28177);
xor U28476 (N_28476,N_28200,N_28003);
nand U28477 (N_28477,N_28239,N_28204);
xor U28478 (N_28478,N_28244,N_28194);
nor U28479 (N_28479,N_28240,N_28247);
or U28480 (N_28480,N_28016,N_28042);
and U28481 (N_28481,N_28064,N_28124);
nand U28482 (N_28482,N_28191,N_28083);
xor U28483 (N_28483,N_28160,N_28187);
nor U28484 (N_28484,N_28159,N_28116);
xnor U28485 (N_28485,N_28138,N_28246);
and U28486 (N_28486,N_28243,N_28125);
or U28487 (N_28487,N_28132,N_28020);
nor U28488 (N_28488,N_28078,N_28094);
xnor U28489 (N_28489,N_28111,N_28166);
or U28490 (N_28490,N_28109,N_28163);
and U28491 (N_28491,N_28209,N_28136);
nand U28492 (N_28492,N_28213,N_28015);
nor U28493 (N_28493,N_28021,N_28046);
nand U28494 (N_28494,N_28067,N_28231);
and U28495 (N_28495,N_28017,N_28074);
nor U28496 (N_28496,N_28051,N_28092);
nand U28497 (N_28497,N_28215,N_28195);
or U28498 (N_28498,N_28089,N_28010);
xnor U28499 (N_28499,N_28053,N_28204);
or U28500 (N_28500,N_28353,N_28250);
or U28501 (N_28501,N_28399,N_28275);
or U28502 (N_28502,N_28254,N_28436);
nor U28503 (N_28503,N_28478,N_28325);
nand U28504 (N_28504,N_28271,N_28311);
nor U28505 (N_28505,N_28346,N_28387);
xor U28506 (N_28506,N_28265,N_28323);
xor U28507 (N_28507,N_28442,N_28397);
xnor U28508 (N_28508,N_28284,N_28391);
or U28509 (N_28509,N_28261,N_28430);
or U28510 (N_28510,N_28290,N_28260);
or U28511 (N_28511,N_28384,N_28274);
xor U28512 (N_28512,N_28447,N_28339);
nand U28513 (N_28513,N_28465,N_28443);
nor U28514 (N_28514,N_28475,N_28354);
or U28515 (N_28515,N_28350,N_28258);
nand U28516 (N_28516,N_28431,N_28422);
or U28517 (N_28517,N_28267,N_28364);
xor U28518 (N_28518,N_28415,N_28379);
nor U28519 (N_28519,N_28300,N_28445);
nand U28520 (N_28520,N_28288,N_28266);
and U28521 (N_28521,N_28345,N_28488);
nand U28522 (N_28522,N_28427,N_28388);
xnor U28523 (N_28523,N_28419,N_28356);
nand U28524 (N_28524,N_28262,N_28413);
xnor U28525 (N_28525,N_28468,N_28362);
xor U28526 (N_28526,N_28278,N_28259);
nand U28527 (N_28527,N_28307,N_28380);
xor U28528 (N_28528,N_28309,N_28410);
or U28529 (N_28529,N_28474,N_28452);
nor U28530 (N_28530,N_28371,N_28302);
xor U28531 (N_28531,N_28322,N_28480);
xor U28532 (N_28532,N_28414,N_28349);
nor U28533 (N_28533,N_28327,N_28303);
and U28534 (N_28534,N_28470,N_28330);
nand U28535 (N_28535,N_28337,N_28299);
nor U28536 (N_28536,N_28441,N_28272);
and U28537 (N_28537,N_28453,N_28333);
xnor U28538 (N_28538,N_28424,N_28378);
nand U28539 (N_28539,N_28398,N_28412);
and U28540 (N_28540,N_28448,N_28263);
xnor U28541 (N_28541,N_28273,N_28357);
xnor U28542 (N_28542,N_28460,N_28375);
or U28543 (N_28543,N_28440,N_28348);
and U28544 (N_28544,N_28490,N_28476);
and U28545 (N_28545,N_28423,N_28359);
nand U28546 (N_28546,N_28301,N_28368);
nor U28547 (N_28547,N_28434,N_28317);
xnor U28548 (N_28548,N_28276,N_28429);
and U28549 (N_28549,N_28283,N_28432);
and U28550 (N_28550,N_28491,N_28407);
nand U28551 (N_28551,N_28459,N_28462);
or U28552 (N_28552,N_28435,N_28433);
nor U28553 (N_28553,N_28269,N_28361);
and U28554 (N_28554,N_28268,N_28363);
xnor U28555 (N_28555,N_28411,N_28409);
nor U28556 (N_28556,N_28485,N_28285);
and U28557 (N_28557,N_28444,N_28426);
nand U28558 (N_28558,N_28377,N_28467);
nand U28559 (N_28559,N_28331,N_28400);
xor U28560 (N_28560,N_28366,N_28402);
xnor U28561 (N_28561,N_28486,N_28342);
nand U28562 (N_28562,N_28291,N_28373);
and U28563 (N_28563,N_28312,N_28489);
or U28564 (N_28564,N_28336,N_28293);
nand U28565 (N_28565,N_28484,N_28393);
xor U28566 (N_28566,N_28252,N_28449);
and U28567 (N_28567,N_28358,N_28332);
and U28568 (N_28568,N_28334,N_28438);
nor U28569 (N_28569,N_28401,N_28463);
or U28570 (N_28570,N_28324,N_28352);
xor U28571 (N_28571,N_28374,N_28295);
nand U28572 (N_28572,N_28277,N_28256);
nand U28573 (N_28573,N_28439,N_28496);
xor U28574 (N_28574,N_28481,N_28341);
xnor U28575 (N_28575,N_28370,N_28394);
nand U28576 (N_28576,N_28479,N_28417);
and U28577 (N_28577,N_28360,N_28286);
nand U28578 (N_28578,N_28310,N_28347);
or U28579 (N_28579,N_28495,N_28456);
or U28580 (N_28580,N_28280,N_28306);
and U28581 (N_28581,N_28313,N_28482);
or U28582 (N_28582,N_28251,N_28257);
or U28583 (N_28583,N_28458,N_28304);
xor U28584 (N_28584,N_28270,N_28319);
or U28585 (N_28585,N_28297,N_28471);
xor U28586 (N_28586,N_28383,N_28494);
and U28587 (N_28587,N_28326,N_28461);
nor U28588 (N_28588,N_28405,N_28382);
xor U28589 (N_28589,N_28320,N_28403);
and U28590 (N_28590,N_28316,N_28483);
nor U28591 (N_28591,N_28492,N_28425);
nand U28592 (N_28592,N_28365,N_28385);
and U28593 (N_28593,N_28386,N_28446);
nor U28594 (N_28594,N_28454,N_28421);
xor U28595 (N_28595,N_28390,N_28338);
and U28596 (N_28596,N_28308,N_28294);
nand U28597 (N_28597,N_28466,N_28437);
xnor U28598 (N_28598,N_28420,N_28396);
and U28599 (N_28599,N_28329,N_28344);
nand U28600 (N_28600,N_28455,N_28493);
and U28601 (N_28601,N_28497,N_28340);
nand U28602 (N_28602,N_28450,N_28395);
or U28603 (N_28603,N_28318,N_28473);
nand U28604 (N_28604,N_28457,N_28315);
xor U28605 (N_28605,N_28321,N_28499);
and U28606 (N_28606,N_28343,N_28298);
and U28607 (N_28607,N_28351,N_28408);
nand U28608 (N_28608,N_28369,N_28281);
or U28609 (N_28609,N_28328,N_28279);
nand U28610 (N_28610,N_28255,N_28389);
nor U28611 (N_28611,N_28416,N_28253);
or U28612 (N_28612,N_28335,N_28406);
nand U28613 (N_28613,N_28287,N_28381);
or U28614 (N_28614,N_28428,N_28487);
or U28615 (N_28615,N_28367,N_28292);
or U28616 (N_28616,N_28289,N_28451);
and U28617 (N_28617,N_28464,N_28376);
or U28618 (N_28618,N_28469,N_28418);
xor U28619 (N_28619,N_28282,N_28355);
nor U28620 (N_28620,N_28392,N_28472);
and U28621 (N_28621,N_28477,N_28296);
or U28622 (N_28622,N_28372,N_28264);
and U28623 (N_28623,N_28305,N_28314);
nor U28624 (N_28624,N_28404,N_28498);
xnor U28625 (N_28625,N_28485,N_28356);
nand U28626 (N_28626,N_28479,N_28438);
xor U28627 (N_28627,N_28432,N_28429);
nor U28628 (N_28628,N_28309,N_28376);
and U28629 (N_28629,N_28369,N_28378);
nor U28630 (N_28630,N_28399,N_28367);
nand U28631 (N_28631,N_28312,N_28479);
nor U28632 (N_28632,N_28276,N_28479);
xnor U28633 (N_28633,N_28453,N_28271);
nand U28634 (N_28634,N_28439,N_28369);
nor U28635 (N_28635,N_28479,N_28283);
nand U28636 (N_28636,N_28430,N_28401);
nor U28637 (N_28637,N_28311,N_28448);
nor U28638 (N_28638,N_28298,N_28430);
xor U28639 (N_28639,N_28442,N_28432);
xnor U28640 (N_28640,N_28360,N_28425);
nand U28641 (N_28641,N_28453,N_28316);
and U28642 (N_28642,N_28432,N_28268);
nor U28643 (N_28643,N_28275,N_28290);
and U28644 (N_28644,N_28380,N_28443);
nor U28645 (N_28645,N_28474,N_28252);
nor U28646 (N_28646,N_28454,N_28402);
or U28647 (N_28647,N_28449,N_28283);
or U28648 (N_28648,N_28493,N_28437);
xnor U28649 (N_28649,N_28396,N_28414);
nand U28650 (N_28650,N_28262,N_28424);
or U28651 (N_28651,N_28420,N_28294);
nor U28652 (N_28652,N_28317,N_28255);
or U28653 (N_28653,N_28305,N_28401);
xor U28654 (N_28654,N_28440,N_28480);
or U28655 (N_28655,N_28475,N_28338);
nor U28656 (N_28656,N_28477,N_28310);
xor U28657 (N_28657,N_28266,N_28342);
nand U28658 (N_28658,N_28386,N_28255);
nand U28659 (N_28659,N_28410,N_28260);
and U28660 (N_28660,N_28448,N_28431);
and U28661 (N_28661,N_28464,N_28348);
or U28662 (N_28662,N_28351,N_28471);
xnor U28663 (N_28663,N_28260,N_28306);
or U28664 (N_28664,N_28471,N_28446);
nand U28665 (N_28665,N_28337,N_28431);
xor U28666 (N_28666,N_28401,N_28458);
and U28667 (N_28667,N_28277,N_28451);
or U28668 (N_28668,N_28433,N_28327);
xor U28669 (N_28669,N_28465,N_28383);
or U28670 (N_28670,N_28344,N_28313);
and U28671 (N_28671,N_28294,N_28477);
xor U28672 (N_28672,N_28277,N_28340);
xor U28673 (N_28673,N_28379,N_28420);
or U28674 (N_28674,N_28459,N_28465);
nand U28675 (N_28675,N_28383,N_28350);
nor U28676 (N_28676,N_28395,N_28375);
nor U28677 (N_28677,N_28488,N_28351);
and U28678 (N_28678,N_28486,N_28334);
xor U28679 (N_28679,N_28411,N_28371);
xor U28680 (N_28680,N_28423,N_28274);
nor U28681 (N_28681,N_28469,N_28437);
and U28682 (N_28682,N_28479,N_28367);
nand U28683 (N_28683,N_28423,N_28411);
xnor U28684 (N_28684,N_28333,N_28367);
nor U28685 (N_28685,N_28475,N_28305);
or U28686 (N_28686,N_28340,N_28428);
or U28687 (N_28687,N_28487,N_28381);
nand U28688 (N_28688,N_28447,N_28464);
xor U28689 (N_28689,N_28324,N_28498);
xnor U28690 (N_28690,N_28354,N_28301);
xnor U28691 (N_28691,N_28389,N_28397);
nand U28692 (N_28692,N_28257,N_28366);
or U28693 (N_28693,N_28385,N_28348);
nor U28694 (N_28694,N_28253,N_28386);
or U28695 (N_28695,N_28368,N_28430);
xor U28696 (N_28696,N_28274,N_28367);
or U28697 (N_28697,N_28293,N_28265);
xnor U28698 (N_28698,N_28470,N_28447);
xnor U28699 (N_28699,N_28354,N_28482);
or U28700 (N_28700,N_28313,N_28404);
nand U28701 (N_28701,N_28383,N_28436);
nor U28702 (N_28702,N_28402,N_28431);
xor U28703 (N_28703,N_28438,N_28395);
xor U28704 (N_28704,N_28310,N_28460);
and U28705 (N_28705,N_28478,N_28291);
and U28706 (N_28706,N_28370,N_28426);
or U28707 (N_28707,N_28269,N_28330);
xnor U28708 (N_28708,N_28331,N_28399);
and U28709 (N_28709,N_28499,N_28296);
nand U28710 (N_28710,N_28324,N_28358);
and U28711 (N_28711,N_28306,N_28366);
xor U28712 (N_28712,N_28317,N_28475);
nand U28713 (N_28713,N_28498,N_28278);
xnor U28714 (N_28714,N_28334,N_28453);
xnor U28715 (N_28715,N_28337,N_28388);
xnor U28716 (N_28716,N_28380,N_28433);
xnor U28717 (N_28717,N_28476,N_28449);
and U28718 (N_28718,N_28363,N_28478);
or U28719 (N_28719,N_28447,N_28376);
nand U28720 (N_28720,N_28405,N_28261);
nand U28721 (N_28721,N_28477,N_28408);
and U28722 (N_28722,N_28407,N_28333);
xnor U28723 (N_28723,N_28391,N_28497);
nor U28724 (N_28724,N_28299,N_28480);
xnor U28725 (N_28725,N_28482,N_28459);
nor U28726 (N_28726,N_28339,N_28326);
nand U28727 (N_28727,N_28376,N_28302);
nand U28728 (N_28728,N_28491,N_28406);
and U28729 (N_28729,N_28432,N_28352);
or U28730 (N_28730,N_28366,N_28399);
nand U28731 (N_28731,N_28482,N_28389);
nor U28732 (N_28732,N_28266,N_28421);
nor U28733 (N_28733,N_28482,N_28259);
nor U28734 (N_28734,N_28420,N_28382);
and U28735 (N_28735,N_28391,N_28473);
or U28736 (N_28736,N_28399,N_28354);
nor U28737 (N_28737,N_28286,N_28376);
nand U28738 (N_28738,N_28389,N_28463);
nor U28739 (N_28739,N_28462,N_28370);
nor U28740 (N_28740,N_28421,N_28463);
nand U28741 (N_28741,N_28313,N_28254);
or U28742 (N_28742,N_28450,N_28282);
and U28743 (N_28743,N_28304,N_28326);
and U28744 (N_28744,N_28489,N_28377);
nand U28745 (N_28745,N_28379,N_28471);
nor U28746 (N_28746,N_28365,N_28370);
nor U28747 (N_28747,N_28399,N_28384);
and U28748 (N_28748,N_28313,N_28479);
nor U28749 (N_28749,N_28460,N_28455);
nand U28750 (N_28750,N_28533,N_28614);
xor U28751 (N_28751,N_28617,N_28641);
nand U28752 (N_28752,N_28733,N_28718);
and U28753 (N_28753,N_28640,N_28577);
nand U28754 (N_28754,N_28698,N_28535);
and U28755 (N_28755,N_28619,N_28727);
and U28756 (N_28756,N_28507,N_28642);
xnor U28757 (N_28757,N_28512,N_28610);
and U28758 (N_28758,N_28513,N_28748);
nand U28759 (N_28759,N_28508,N_28729);
nor U28760 (N_28760,N_28655,N_28519);
nand U28761 (N_28761,N_28529,N_28570);
xnor U28762 (N_28762,N_28561,N_28633);
nor U28763 (N_28763,N_28602,N_28663);
nor U28764 (N_28764,N_28590,N_28639);
nand U28765 (N_28765,N_28681,N_28580);
nor U28766 (N_28766,N_28726,N_28562);
and U28767 (N_28767,N_28711,N_28611);
nand U28768 (N_28768,N_28690,N_28695);
xor U28769 (N_28769,N_28588,N_28616);
or U28770 (N_28770,N_28716,N_28500);
nor U28771 (N_28771,N_28520,N_28649);
and U28772 (N_28772,N_28702,N_28556);
nor U28773 (N_28773,N_28571,N_28591);
nand U28774 (N_28774,N_28662,N_28630);
nand U28775 (N_28775,N_28675,N_28717);
nand U28776 (N_28776,N_28521,N_28682);
or U28777 (N_28777,N_28618,N_28514);
or U28778 (N_28778,N_28604,N_28502);
or U28779 (N_28779,N_28730,N_28582);
or U28780 (N_28780,N_28539,N_28693);
nor U28781 (N_28781,N_28615,N_28605);
nor U28782 (N_28782,N_28665,N_28537);
nor U28783 (N_28783,N_28623,N_28701);
or U28784 (N_28784,N_28548,N_28731);
or U28785 (N_28785,N_28517,N_28524);
xnor U28786 (N_28786,N_28527,N_28593);
or U28787 (N_28787,N_28549,N_28509);
and U28788 (N_28788,N_28585,N_28708);
nor U28789 (N_28789,N_28565,N_28657);
xnor U28790 (N_28790,N_28558,N_28581);
or U28791 (N_28791,N_28723,N_28686);
nand U28792 (N_28792,N_28559,N_28722);
xor U28793 (N_28793,N_28721,N_28528);
xor U28794 (N_28794,N_28551,N_28575);
or U28795 (N_28795,N_28504,N_28706);
nor U28796 (N_28796,N_28697,N_28530);
nand U28797 (N_28797,N_28555,N_28595);
xor U28798 (N_28798,N_28710,N_28645);
or U28799 (N_28799,N_28647,N_28525);
nor U28800 (N_28800,N_28659,N_28739);
nand U28801 (N_28801,N_28749,N_28676);
nand U28802 (N_28802,N_28724,N_28734);
and U28803 (N_28803,N_28511,N_28713);
or U28804 (N_28804,N_28703,N_28705);
or U28805 (N_28805,N_28691,N_28546);
xor U28806 (N_28806,N_28725,N_28668);
and U28807 (N_28807,N_28720,N_28576);
nor U28808 (N_28808,N_28568,N_28597);
and U28809 (N_28809,N_28531,N_28601);
and U28810 (N_28810,N_28737,N_28685);
nand U28811 (N_28811,N_28715,N_28547);
and U28812 (N_28812,N_28743,N_28628);
or U28813 (N_28813,N_28586,N_28566);
nor U28814 (N_28814,N_28719,N_28596);
or U28815 (N_28815,N_28683,N_28506);
and U28816 (N_28816,N_28741,N_28745);
and U28817 (N_28817,N_28545,N_28684);
and U28818 (N_28818,N_28603,N_28728);
nand U28819 (N_28819,N_28563,N_28678);
xnor U28820 (N_28820,N_28666,N_28510);
nand U28821 (N_28821,N_28608,N_28516);
nor U28822 (N_28822,N_28583,N_28599);
nor U28823 (N_28823,N_28632,N_28573);
or U28824 (N_28824,N_28631,N_28636);
or U28825 (N_28825,N_28694,N_28624);
and U28826 (N_28826,N_28589,N_28552);
nand U28827 (N_28827,N_28541,N_28522);
and U28828 (N_28828,N_28612,N_28526);
nand U28829 (N_28829,N_28592,N_28637);
and U28830 (N_28830,N_28661,N_28664);
nand U28831 (N_28831,N_28532,N_28560);
xnor U28832 (N_28832,N_28704,N_28550);
and U28833 (N_28833,N_28638,N_28621);
xor U28834 (N_28834,N_28584,N_28687);
nand U28835 (N_28835,N_28736,N_28742);
nand U28836 (N_28836,N_28578,N_28680);
nand U28837 (N_28837,N_28712,N_28627);
nor U28838 (N_28838,N_28620,N_28518);
xor U28839 (N_28839,N_28643,N_28609);
or U28840 (N_28840,N_28626,N_28579);
nor U28841 (N_28841,N_28644,N_28653);
and U28842 (N_28842,N_28543,N_28622);
xor U28843 (N_28843,N_28635,N_28746);
xnor U28844 (N_28844,N_28542,N_28672);
xnor U28845 (N_28845,N_28651,N_28667);
xnor U28846 (N_28846,N_28569,N_28646);
and U28847 (N_28847,N_28594,N_28696);
or U28848 (N_28848,N_28732,N_28606);
and U28849 (N_28849,N_28700,N_28654);
or U28850 (N_28850,N_28707,N_28536);
nor U28851 (N_28851,N_28699,N_28544);
and U28852 (N_28852,N_28673,N_28738);
nor U28853 (N_28853,N_28540,N_28650);
or U28854 (N_28854,N_28515,N_28648);
nand U28855 (N_28855,N_28553,N_28677);
nor U28856 (N_28856,N_28658,N_28689);
nor U28857 (N_28857,N_28501,N_28670);
nand U28858 (N_28858,N_28505,N_28598);
or U28859 (N_28859,N_28692,N_28613);
and U28860 (N_28860,N_28747,N_28709);
or U28861 (N_28861,N_28574,N_28744);
xnor U28862 (N_28862,N_28735,N_28572);
and U28863 (N_28863,N_28629,N_28634);
and U28864 (N_28864,N_28587,N_28656);
or U28865 (N_28865,N_28607,N_28714);
and U28866 (N_28866,N_28688,N_28660);
nand U28867 (N_28867,N_28600,N_28523);
or U28868 (N_28868,N_28674,N_28671);
xor U28869 (N_28869,N_28652,N_28557);
and U28870 (N_28870,N_28625,N_28567);
nor U28871 (N_28871,N_28554,N_28503);
xor U28872 (N_28872,N_28669,N_28564);
or U28873 (N_28873,N_28740,N_28538);
nand U28874 (N_28874,N_28679,N_28534);
or U28875 (N_28875,N_28670,N_28657);
or U28876 (N_28876,N_28522,N_28666);
and U28877 (N_28877,N_28739,N_28517);
or U28878 (N_28878,N_28583,N_28680);
and U28879 (N_28879,N_28593,N_28515);
or U28880 (N_28880,N_28553,N_28533);
or U28881 (N_28881,N_28511,N_28541);
nor U28882 (N_28882,N_28691,N_28748);
nor U28883 (N_28883,N_28501,N_28543);
nand U28884 (N_28884,N_28573,N_28699);
or U28885 (N_28885,N_28574,N_28734);
nand U28886 (N_28886,N_28610,N_28746);
nor U28887 (N_28887,N_28591,N_28618);
nand U28888 (N_28888,N_28720,N_28547);
nand U28889 (N_28889,N_28727,N_28725);
or U28890 (N_28890,N_28708,N_28649);
and U28891 (N_28891,N_28590,N_28739);
nand U28892 (N_28892,N_28643,N_28591);
or U28893 (N_28893,N_28585,N_28594);
and U28894 (N_28894,N_28716,N_28591);
xnor U28895 (N_28895,N_28686,N_28567);
or U28896 (N_28896,N_28610,N_28511);
or U28897 (N_28897,N_28545,N_28516);
or U28898 (N_28898,N_28664,N_28731);
nor U28899 (N_28899,N_28668,N_28727);
or U28900 (N_28900,N_28515,N_28641);
nor U28901 (N_28901,N_28568,N_28562);
nand U28902 (N_28902,N_28661,N_28749);
nand U28903 (N_28903,N_28660,N_28610);
and U28904 (N_28904,N_28572,N_28612);
xnor U28905 (N_28905,N_28673,N_28630);
xor U28906 (N_28906,N_28529,N_28563);
or U28907 (N_28907,N_28540,N_28582);
nand U28908 (N_28908,N_28720,N_28549);
nand U28909 (N_28909,N_28622,N_28607);
xnor U28910 (N_28910,N_28650,N_28594);
nor U28911 (N_28911,N_28719,N_28569);
and U28912 (N_28912,N_28676,N_28663);
nand U28913 (N_28913,N_28644,N_28717);
nor U28914 (N_28914,N_28646,N_28632);
or U28915 (N_28915,N_28575,N_28737);
nor U28916 (N_28916,N_28675,N_28601);
xor U28917 (N_28917,N_28527,N_28731);
nand U28918 (N_28918,N_28657,N_28708);
xnor U28919 (N_28919,N_28661,N_28643);
and U28920 (N_28920,N_28613,N_28627);
and U28921 (N_28921,N_28512,N_28593);
xor U28922 (N_28922,N_28594,N_28531);
nand U28923 (N_28923,N_28740,N_28506);
nand U28924 (N_28924,N_28695,N_28548);
nor U28925 (N_28925,N_28570,N_28715);
nor U28926 (N_28926,N_28713,N_28728);
nand U28927 (N_28927,N_28749,N_28702);
and U28928 (N_28928,N_28535,N_28748);
and U28929 (N_28929,N_28632,N_28732);
nor U28930 (N_28930,N_28642,N_28681);
nor U28931 (N_28931,N_28521,N_28731);
nand U28932 (N_28932,N_28571,N_28501);
nand U28933 (N_28933,N_28631,N_28583);
nand U28934 (N_28934,N_28507,N_28737);
and U28935 (N_28935,N_28510,N_28562);
nor U28936 (N_28936,N_28696,N_28727);
or U28937 (N_28937,N_28517,N_28612);
or U28938 (N_28938,N_28666,N_28547);
and U28939 (N_28939,N_28699,N_28734);
and U28940 (N_28940,N_28522,N_28656);
or U28941 (N_28941,N_28702,N_28582);
nand U28942 (N_28942,N_28532,N_28501);
xnor U28943 (N_28943,N_28689,N_28710);
xor U28944 (N_28944,N_28698,N_28647);
xor U28945 (N_28945,N_28611,N_28529);
xor U28946 (N_28946,N_28674,N_28560);
nor U28947 (N_28947,N_28698,N_28560);
nand U28948 (N_28948,N_28597,N_28621);
nor U28949 (N_28949,N_28630,N_28588);
or U28950 (N_28950,N_28602,N_28572);
nand U28951 (N_28951,N_28597,N_28539);
nor U28952 (N_28952,N_28701,N_28721);
and U28953 (N_28953,N_28594,N_28693);
and U28954 (N_28954,N_28670,N_28510);
nor U28955 (N_28955,N_28617,N_28535);
and U28956 (N_28956,N_28521,N_28723);
nor U28957 (N_28957,N_28640,N_28741);
nand U28958 (N_28958,N_28523,N_28529);
xor U28959 (N_28959,N_28558,N_28692);
or U28960 (N_28960,N_28629,N_28657);
or U28961 (N_28961,N_28527,N_28601);
xor U28962 (N_28962,N_28679,N_28734);
nand U28963 (N_28963,N_28641,N_28681);
xnor U28964 (N_28964,N_28670,N_28602);
and U28965 (N_28965,N_28628,N_28629);
nor U28966 (N_28966,N_28679,N_28655);
nand U28967 (N_28967,N_28674,N_28629);
nand U28968 (N_28968,N_28686,N_28542);
nor U28969 (N_28969,N_28642,N_28731);
xor U28970 (N_28970,N_28707,N_28714);
xnor U28971 (N_28971,N_28511,N_28698);
or U28972 (N_28972,N_28659,N_28624);
and U28973 (N_28973,N_28588,N_28596);
xnor U28974 (N_28974,N_28679,N_28730);
nor U28975 (N_28975,N_28522,N_28704);
nor U28976 (N_28976,N_28536,N_28729);
or U28977 (N_28977,N_28611,N_28520);
nand U28978 (N_28978,N_28729,N_28556);
xnor U28979 (N_28979,N_28586,N_28696);
or U28980 (N_28980,N_28638,N_28647);
nand U28981 (N_28981,N_28518,N_28610);
or U28982 (N_28982,N_28694,N_28605);
xor U28983 (N_28983,N_28608,N_28698);
nor U28984 (N_28984,N_28512,N_28540);
nor U28985 (N_28985,N_28626,N_28587);
or U28986 (N_28986,N_28543,N_28646);
and U28987 (N_28987,N_28626,N_28739);
and U28988 (N_28988,N_28606,N_28601);
xor U28989 (N_28989,N_28678,N_28686);
nor U28990 (N_28990,N_28727,N_28726);
xor U28991 (N_28991,N_28571,N_28627);
and U28992 (N_28992,N_28534,N_28559);
xnor U28993 (N_28993,N_28572,N_28627);
and U28994 (N_28994,N_28644,N_28595);
and U28995 (N_28995,N_28581,N_28625);
nor U28996 (N_28996,N_28553,N_28747);
or U28997 (N_28997,N_28692,N_28579);
nor U28998 (N_28998,N_28733,N_28657);
nand U28999 (N_28999,N_28551,N_28543);
or U29000 (N_29000,N_28915,N_28896);
nand U29001 (N_29001,N_28796,N_28939);
nor U29002 (N_29002,N_28867,N_28982);
nor U29003 (N_29003,N_28839,N_28759);
or U29004 (N_29004,N_28996,N_28856);
nand U29005 (N_29005,N_28878,N_28859);
nand U29006 (N_29006,N_28795,N_28751);
xor U29007 (N_29007,N_28928,N_28998);
nand U29008 (N_29008,N_28918,N_28969);
xnor U29009 (N_29009,N_28841,N_28756);
and U29010 (N_29010,N_28934,N_28792);
nand U29011 (N_29011,N_28767,N_28852);
nand U29012 (N_29012,N_28973,N_28970);
and U29013 (N_29013,N_28848,N_28858);
nor U29014 (N_29014,N_28765,N_28819);
and U29015 (N_29015,N_28788,N_28902);
xnor U29016 (N_29016,N_28961,N_28750);
xor U29017 (N_29017,N_28886,N_28964);
nand U29018 (N_29018,N_28962,N_28942);
nand U29019 (N_29019,N_28836,N_28978);
nand U29020 (N_29020,N_28823,N_28757);
and U29021 (N_29021,N_28953,N_28776);
xnor U29022 (N_29022,N_28903,N_28826);
nand U29023 (N_29023,N_28794,N_28763);
and U29024 (N_29024,N_28883,N_28809);
nor U29025 (N_29025,N_28793,N_28875);
xor U29026 (N_29026,N_28943,N_28887);
nor U29027 (N_29027,N_28944,N_28917);
or U29028 (N_29028,N_28881,N_28766);
or U29029 (N_29029,N_28815,N_28864);
xor U29030 (N_29030,N_28929,N_28895);
nand U29031 (N_29031,N_28938,N_28817);
xor U29032 (N_29032,N_28808,N_28912);
nor U29033 (N_29033,N_28968,N_28862);
nor U29034 (N_29034,N_28870,N_28910);
nand U29035 (N_29035,N_28785,N_28778);
nand U29036 (N_29036,N_28958,N_28775);
nor U29037 (N_29037,N_28913,N_28866);
or U29038 (N_29038,N_28777,N_28773);
nand U29039 (N_29039,N_28937,N_28892);
nand U29040 (N_29040,N_28916,N_28879);
nor U29041 (N_29041,N_28835,N_28779);
xor U29042 (N_29042,N_28814,N_28807);
or U29043 (N_29043,N_28921,N_28963);
nand U29044 (N_29044,N_28984,N_28798);
xor U29045 (N_29045,N_28806,N_28832);
or U29046 (N_29046,N_28956,N_28891);
or U29047 (N_29047,N_28803,N_28908);
or U29048 (N_29048,N_28853,N_28829);
nand U29049 (N_29049,N_28760,N_28905);
xor U29050 (N_29050,N_28752,N_28847);
or U29051 (N_29051,N_28999,N_28790);
or U29052 (N_29052,N_28889,N_28898);
xor U29053 (N_29053,N_28936,N_28843);
or U29054 (N_29054,N_28783,N_28799);
xor U29055 (N_29055,N_28805,N_28769);
nand U29056 (N_29056,N_28840,N_28972);
and U29057 (N_29057,N_28827,N_28894);
nand U29058 (N_29058,N_28957,N_28874);
nand U29059 (N_29059,N_28876,N_28945);
xnor U29060 (N_29060,N_28791,N_28824);
or U29061 (N_29061,N_28959,N_28872);
nand U29062 (N_29062,N_28911,N_28940);
or U29063 (N_29063,N_28860,N_28981);
and U29064 (N_29064,N_28993,N_28787);
xor U29065 (N_29065,N_28979,N_28931);
or U29066 (N_29066,N_28927,N_28971);
nand U29067 (N_29067,N_28770,N_28967);
nor U29068 (N_29068,N_28897,N_28988);
and U29069 (N_29069,N_28987,N_28922);
nor U29070 (N_29070,N_28828,N_28965);
and U29071 (N_29071,N_28857,N_28816);
nand U29072 (N_29072,N_28850,N_28997);
or U29073 (N_29073,N_28994,N_28904);
nor U29074 (N_29074,N_28920,N_28755);
and U29075 (N_29075,N_28985,N_28907);
nand U29076 (N_29076,N_28764,N_28820);
xor U29077 (N_29077,N_28849,N_28954);
nand U29078 (N_29078,N_28761,N_28933);
nand U29079 (N_29079,N_28831,N_28797);
and U29080 (N_29080,N_28837,N_28762);
nand U29081 (N_29081,N_28885,N_28990);
or U29082 (N_29082,N_28935,N_28789);
xor U29083 (N_29083,N_28854,N_28974);
and U29084 (N_29084,N_28774,N_28890);
nand U29085 (N_29085,N_28845,N_28949);
nor U29086 (N_29086,N_28865,N_28966);
and U29087 (N_29087,N_28871,N_28782);
nand U29088 (N_29088,N_28926,N_28882);
and U29089 (N_29089,N_28975,N_28880);
xor U29090 (N_29090,N_28977,N_28822);
and U29091 (N_29091,N_28877,N_28952);
nand U29092 (N_29092,N_28893,N_28951);
or U29093 (N_29093,N_28818,N_28801);
nor U29094 (N_29094,N_28950,N_28834);
nor U29095 (N_29095,N_28821,N_28914);
nor U29096 (N_29096,N_28842,N_28989);
xnor U29097 (N_29097,N_28812,N_28986);
and U29098 (N_29098,N_28861,N_28802);
nand U29099 (N_29099,N_28899,N_28909);
or U29100 (N_29100,N_28781,N_28771);
xor U29101 (N_29101,N_28924,N_28955);
and U29102 (N_29102,N_28784,N_28855);
or U29103 (N_29103,N_28780,N_28923);
and U29104 (N_29104,N_28948,N_28932);
and U29105 (N_29105,N_28800,N_28869);
and U29106 (N_29106,N_28992,N_28930);
and U29107 (N_29107,N_28753,N_28754);
nand U29108 (N_29108,N_28830,N_28825);
nand U29109 (N_29109,N_28946,N_28873);
xnor U29110 (N_29110,N_28925,N_28844);
or U29111 (N_29111,N_28863,N_28810);
xor U29112 (N_29112,N_28851,N_28811);
xor U29113 (N_29113,N_28846,N_28884);
nand U29114 (N_29114,N_28868,N_28786);
xnor U29115 (N_29115,N_28838,N_28941);
or U29116 (N_29116,N_28804,N_28991);
nor U29117 (N_29117,N_28901,N_28919);
xor U29118 (N_29118,N_28813,N_28995);
xnor U29119 (N_29119,N_28947,N_28900);
or U29120 (N_29120,N_28833,N_28976);
and U29121 (N_29121,N_28980,N_28983);
or U29122 (N_29122,N_28906,N_28758);
nor U29123 (N_29123,N_28768,N_28888);
or U29124 (N_29124,N_28772,N_28960);
or U29125 (N_29125,N_28977,N_28784);
or U29126 (N_29126,N_28997,N_28756);
and U29127 (N_29127,N_28941,N_28971);
nand U29128 (N_29128,N_28843,N_28777);
xnor U29129 (N_29129,N_28807,N_28751);
xnor U29130 (N_29130,N_28763,N_28856);
xor U29131 (N_29131,N_28860,N_28958);
or U29132 (N_29132,N_28834,N_28880);
nand U29133 (N_29133,N_28972,N_28882);
nor U29134 (N_29134,N_28753,N_28916);
nand U29135 (N_29135,N_28940,N_28967);
and U29136 (N_29136,N_28787,N_28758);
nor U29137 (N_29137,N_28753,N_28806);
or U29138 (N_29138,N_28799,N_28862);
nor U29139 (N_29139,N_28986,N_28875);
and U29140 (N_29140,N_28923,N_28909);
nand U29141 (N_29141,N_28856,N_28903);
and U29142 (N_29142,N_28924,N_28873);
xnor U29143 (N_29143,N_28865,N_28816);
xnor U29144 (N_29144,N_28997,N_28821);
nand U29145 (N_29145,N_28898,N_28904);
or U29146 (N_29146,N_28909,N_28912);
nor U29147 (N_29147,N_28891,N_28973);
and U29148 (N_29148,N_28865,N_28903);
or U29149 (N_29149,N_28782,N_28754);
nand U29150 (N_29150,N_28906,N_28913);
nor U29151 (N_29151,N_28790,N_28990);
xnor U29152 (N_29152,N_28879,N_28789);
and U29153 (N_29153,N_28805,N_28939);
nor U29154 (N_29154,N_28974,N_28941);
nand U29155 (N_29155,N_28861,N_28988);
and U29156 (N_29156,N_28876,N_28903);
and U29157 (N_29157,N_28940,N_28813);
or U29158 (N_29158,N_28808,N_28940);
xor U29159 (N_29159,N_28762,N_28831);
or U29160 (N_29160,N_28780,N_28994);
or U29161 (N_29161,N_28980,N_28998);
and U29162 (N_29162,N_28957,N_28849);
nand U29163 (N_29163,N_28817,N_28891);
xor U29164 (N_29164,N_28863,N_28935);
or U29165 (N_29165,N_28796,N_28944);
or U29166 (N_29166,N_28771,N_28841);
nor U29167 (N_29167,N_28823,N_28903);
nor U29168 (N_29168,N_28848,N_28873);
nor U29169 (N_29169,N_28863,N_28988);
nand U29170 (N_29170,N_28936,N_28890);
nand U29171 (N_29171,N_28981,N_28841);
nor U29172 (N_29172,N_28970,N_28808);
and U29173 (N_29173,N_28991,N_28995);
nand U29174 (N_29174,N_28779,N_28982);
nand U29175 (N_29175,N_28885,N_28919);
nand U29176 (N_29176,N_28830,N_28988);
xnor U29177 (N_29177,N_28883,N_28792);
nand U29178 (N_29178,N_28762,N_28835);
or U29179 (N_29179,N_28985,N_28897);
xnor U29180 (N_29180,N_28927,N_28879);
or U29181 (N_29181,N_28781,N_28812);
xor U29182 (N_29182,N_28782,N_28834);
or U29183 (N_29183,N_28875,N_28949);
and U29184 (N_29184,N_28837,N_28900);
nor U29185 (N_29185,N_28967,N_28911);
or U29186 (N_29186,N_28847,N_28965);
or U29187 (N_29187,N_28976,N_28979);
nand U29188 (N_29188,N_28790,N_28793);
and U29189 (N_29189,N_28862,N_28914);
or U29190 (N_29190,N_28957,N_28833);
xor U29191 (N_29191,N_28962,N_28950);
nor U29192 (N_29192,N_28891,N_28914);
nor U29193 (N_29193,N_28757,N_28820);
nor U29194 (N_29194,N_28895,N_28983);
and U29195 (N_29195,N_28943,N_28871);
nand U29196 (N_29196,N_28980,N_28786);
nand U29197 (N_29197,N_28975,N_28775);
nor U29198 (N_29198,N_28885,N_28957);
xor U29199 (N_29199,N_28938,N_28848);
nor U29200 (N_29200,N_28884,N_28988);
nand U29201 (N_29201,N_28794,N_28888);
nand U29202 (N_29202,N_28906,N_28805);
nand U29203 (N_29203,N_28808,N_28931);
nand U29204 (N_29204,N_28994,N_28963);
and U29205 (N_29205,N_28964,N_28813);
nor U29206 (N_29206,N_28782,N_28965);
nor U29207 (N_29207,N_28910,N_28907);
xor U29208 (N_29208,N_28807,N_28857);
nor U29209 (N_29209,N_28983,N_28884);
or U29210 (N_29210,N_28857,N_28840);
or U29211 (N_29211,N_28938,N_28832);
or U29212 (N_29212,N_28793,N_28768);
or U29213 (N_29213,N_28958,N_28990);
and U29214 (N_29214,N_28883,N_28948);
nor U29215 (N_29215,N_28926,N_28942);
xor U29216 (N_29216,N_28918,N_28876);
and U29217 (N_29217,N_28889,N_28826);
nor U29218 (N_29218,N_28898,N_28982);
nand U29219 (N_29219,N_28887,N_28901);
and U29220 (N_29220,N_28973,N_28968);
or U29221 (N_29221,N_28822,N_28931);
nor U29222 (N_29222,N_28865,N_28886);
xnor U29223 (N_29223,N_28971,N_28852);
xor U29224 (N_29224,N_28917,N_28812);
and U29225 (N_29225,N_28784,N_28900);
or U29226 (N_29226,N_28991,N_28954);
and U29227 (N_29227,N_28910,N_28845);
and U29228 (N_29228,N_28838,N_28768);
or U29229 (N_29229,N_28760,N_28781);
nor U29230 (N_29230,N_28771,N_28955);
nor U29231 (N_29231,N_28767,N_28825);
or U29232 (N_29232,N_28785,N_28961);
nor U29233 (N_29233,N_28760,N_28853);
and U29234 (N_29234,N_28936,N_28993);
xor U29235 (N_29235,N_28900,N_28811);
nor U29236 (N_29236,N_28768,N_28764);
xnor U29237 (N_29237,N_28987,N_28753);
or U29238 (N_29238,N_28951,N_28963);
or U29239 (N_29239,N_28956,N_28950);
and U29240 (N_29240,N_28787,N_28914);
nor U29241 (N_29241,N_28856,N_28761);
nor U29242 (N_29242,N_28786,N_28855);
or U29243 (N_29243,N_28969,N_28810);
nand U29244 (N_29244,N_28841,N_28755);
xor U29245 (N_29245,N_28848,N_28889);
xnor U29246 (N_29246,N_28977,N_28794);
nand U29247 (N_29247,N_28758,N_28947);
or U29248 (N_29248,N_28799,N_28785);
nand U29249 (N_29249,N_28793,N_28905);
nand U29250 (N_29250,N_29244,N_29097);
nor U29251 (N_29251,N_29236,N_29240);
or U29252 (N_29252,N_29031,N_29177);
xor U29253 (N_29253,N_29207,N_29117);
nand U29254 (N_29254,N_29011,N_29182);
xor U29255 (N_29255,N_29110,N_29028);
and U29256 (N_29256,N_29226,N_29176);
xor U29257 (N_29257,N_29037,N_29052);
nor U29258 (N_29258,N_29094,N_29151);
nor U29259 (N_29259,N_29133,N_29090);
or U29260 (N_29260,N_29223,N_29054);
or U29261 (N_29261,N_29169,N_29118);
xnor U29262 (N_29262,N_29022,N_29019);
and U29263 (N_29263,N_29233,N_29068);
nor U29264 (N_29264,N_29100,N_29039);
or U29265 (N_29265,N_29196,N_29087);
or U29266 (N_29266,N_29030,N_29245);
xor U29267 (N_29267,N_29212,N_29101);
nor U29268 (N_29268,N_29173,N_29040);
xor U29269 (N_29269,N_29130,N_29153);
nor U29270 (N_29270,N_29138,N_29201);
or U29271 (N_29271,N_29045,N_29184);
nor U29272 (N_29272,N_29034,N_29145);
or U29273 (N_29273,N_29164,N_29204);
or U29274 (N_29274,N_29246,N_29210);
nor U29275 (N_29275,N_29088,N_29092);
or U29276 (N_29276,N_29242,N_29041);
and U29277 (N_29277,N_29220,N_29044);
xor U29278 (N_29278,N_29005,N_29111);
nand U29279 (N_29279,N_29155,N_29132);
or U29280 (N_29280,N_29183,N_29229);
nor U29281 (N_29281,N_29208,N_29074);
and U29282 (N_29282,N_29163,N_29181);
and U29283 (N_29283,N_29107,N_29228);
and U29284 (N_29284,N_29065,N_29168);
nand U29285 (N_29285,N_29061,N_29070);
xor U29286 (N_29286,N_29033,N_29002);
nand U29287 (N_29287,N_29072,N_29116);
xor U29288 (N_29288,N_29160,N_29016);
xor U29289 (N_29289,N_29053,N_29025);
nor U29290 (N_29290,N_29069,N_29214);
nand U29291 (N_29291,N_29077,N_29066);
and U29292 (N_29292,N_29215,N_29056);
nor U29293 (N_29293,N_29147,N_29239);
nor U29294 (N_29294,N_29199,N_29194);
nor U29295 (N_29295,N_29172,N_29216);
and U29296 (N_29296,N_29222,N_29139);
xnor U29297 (N_29297,N_29067,N_29165);
or U29298 (N_29298,N_29079,N_29095);
xor U29299 (N_29299,N_29142,N_29080);
and U29300 (N_29300,N_29075,N_29178);
nor U29301 (N_29301,N_29119,N_29180);
and U29302 (N_29302,N_29186,N_29064);
or U29303 (N_29303,N_29000,N_29193);
and U29304 (N_29304,N_29235,N_29157);
xnor U29305 (N_29305,N_29108,N_29049);
or U29306 (N_29306,N_29148,N_29021);
xnor U29307 (N_29307,N_29013,N_29035);
xor U29308 (N_29308,N_29237,N_29185);
nand U29309 (N_29309,N_29209,N_29230);
xor U29310 (N_29310,N_29225,N_29241);
xor U29311 (N_29311,N_29202,N_29018);
and U29312 (N_29312,N_29047,N_29006);
nand U29313 (N_29313,N_29113,N_29057);
and U29314 (N_29314,N_29023,N_29140);
xnor U29315 (N_29315,N_29008,N_29048);
nor U29316 (N_29316,N_29096,N_29091);
and U29317 (N_29317,N_29143,N_29050);
xnor U29318 (N_29318,N_29024,N_29027);
nand U29319 (N_29319,N_29082,N_29234);
nor U29320 (N_29320,N_29170,N_29159);
xnor U29321 (N_29321,N_29106,N_29017);
or U29322 (N_29322,N_29156,N_29051);
xor U29323 (N_29323,N_29227,N_29109);
nor U29324 (N_29324,N_29029,N_29224);
or U29325 (N_29325,N_29131,N_29136);
nand U29326 (N_29326,N_29158,N_29063);
nand U29327 (N_29327,N_29007,N_29012);
or U29328 (N_29328,N_29078,N_29003);
or U29329 (N_29329,N_29032,N_29010);
nand U29330 (N_29330,N_29200,N_29055);
xnor U29331 (N_29331,N_29102,N_29152);
xor U29332 (N_29332,N_29043,N_29076);
nor U29333 (N_29333,N_29205,N_29015);
and U29334 (N_29334,N_29127,N_29114);
nand U29335 (N_29335,N_29103,N_29026);
xor U29336 (N_29336,N_29219,N_29203);
nand U29337 (N_29337,N_29206,N_29059);
or U29338 (N_29338,N_29174,N_29238);
nor U29339 (N_29339,N_29104,N_29195);
or U29340 (N_29340,N_29060,N_29062);
nor U29341 (N_29341,N_29073,N_29046);
nor U29342 (N_29342,N_29084,N_29071);
nor U29343 (N_29343,N_29099,N_29122);
or U29344 (N_29344,N_29190,N_29086);
or U29345 (N_29345,N_29081,N_29129);
nor U29346 (N_29346,N_29009,N_29083);
nand U29347 (N_29347,N_29232,N_29105);
nor U29348 (N_29348,N_29243,N_29188);
nor U29349 (N_29349,N_29213,N_29014);
nor U29350 (N_29350,N_29248,N_29218);
nand U29351 (N_29351,N_29141,N_29115);
xnor U29352 (N_29352,N_29217,N_29098);
xor U29353 (N_29353,N_29001,N_29189);
nor U29354 (N_29354,N_29161,N_29038);
nand U29355 (N_29355,N_29144,N_29231);
xnor U29356 (N_29356,N_29126,N_29150);
or U29357 (N_29357,N_29197,N_29162);
nor U29358 (N_29358,N_29249,N_29089);
xnor U29359 (N_29359,N_29042,N_29124);
nand U29360 (N_29360,N_29154,N_29175);
xnor U29361 (N_29361,N_29125,N_29036);
nor U29362 (N_29362,N_29128,N_29192);
xor U29363 (N_29363,N_29179,N_29112);
nand U29364 (N_29364,N_29211,N_29146);
nor U29365 (N_29365,N_29020,N_29191);
and U29366 (N_29366,N_29137,N_29093);
and U29367 (N_29367,N_29149,N_29166);
nand U29368 (N_29368,N_29171,N_29187);
xnor U29369 (N_29369,N_29247,N_29058);
xnor U29370 (N_29370,N_29085,N_29167);
nand U29371 (N_29371,N_29123,N_29134);
nand U29372 (N_29372,N_29121,N_29120);
or U29373 (N_29373,N_29221,N_29004);
nor U29374 (N_29374,N_29135,N_29198);
and U29375 (N_29375,N_29225,N_29228);
nor U29376 (N_29376,N_29067,N_29023);
xor U29377 (N_29377,N_29198,N_29147);
nor U29378 (N_29378,N_29083,N_29015);
xnor U29379 (N_29379,N_29068,N_29122);
nor U29380 (N_29380,N_29244,N_29089);
nor U29381 (N_29381,N_29245,N_29063);
nand U29382 (N_29382,N_29075,N_29240);
nand U29383 (N_29383,N_29056,N_29101);
xor U29384 (N_29384,N_29238,N_29191);
nand U29385 (N_29385,N_29082,N_29076);
and U29386 (N_29386,N_29164,N_29189);
and U29387 (N_29387,N_29064,N_29209);
nor U29388 (N_29388,N_29137,N_29217);
and U29389 (N_29389,N_29156,N_29044);
and U29390 (N_29390,N_29159,N_29024);
nand U29391 (N_29391,N_29186,N_29002);
xnor U29392 (N_29392,N_29218,N_29044);
nand U29393 (N_29393,N_29244,N_29104);
or U29394 (N_29394,N_29134,N_29069);
or U29395 (N_29395,N_29076,N_29027);
and U29396 (N_29396,N_29009,N_29068);
and U29397 (N_29397,N_29030,N_29243);
or U29398 (N_29398,N_29036,N_29200);
or U29399 (N_29399,N_29217,N_29088);
and U29400 (N_29400,N_29066,N_29056);
nor U29401 (N_29401,N_29094,N_29113);
or U29402 (N_29402,N_29053,N_29184);
xor U29403 (N_29403,N_29111,N_29191);
nand U29404 (N_29404,N_29047,N_29150);
or U29405 (N_29405,N_29061,N_29063);
nor U29406 (N_29406,N_29161,N_29245);
and U29407 (N_29407,N_29060,N_29075);
nor U29408 (N_29408,N_29095,N_29017);
and U29409 (N_29409,N_29104,N_29041);
xor U29410 (N_29410,N_29161,N_29210);
nand U29411 (N_29411,N_29223,N_29147);
nor U29412 (N_29412,N_29244,N_29229);
nor U29413 (N_29413,N_29134,N_29074);
nand U29414 (N_29414,N_29045,N_29127);
and U29415 (N_29415,N_29129,N_29136);
nor U29416 (N_29416,N_29206,N_29195);
nand U29417 (N_29417,N_29068,N_29105);
nor U29418 (N_29418,N_29115,N_29214);
and U29419 (N_29419,N_29037,N_29192);
nor U29420 (N_29420,N_29154,N_29161);
nand U29421 (N_29421,N_29218,N_29164);
nor U29422 (N_29422,N_29194,N_29229);
nor U29423 (N_29423,N_29052,N_29115);
nor U29424 (N_29424,N_29222,N_29239);
xor U29425 (N_29425,N_29144,N_29058);
xnor U29426 (N_29426,N_29199,N_29103);
xnor U29427 (N_29427,N_29135,N_29168);
nand U29428 (N_29428,N_29144,N_29174);
and U29429 (N_29429,N_29177,N_29145);
or U29430 (N_29430,N_29052,N_29025);
nor U29431 (N_29431,N_29156,N_29099);
nand U29432 (N_29432,N_29087,N_29185);
or U29433 (N_29433,N_29063,N_29083);
xnor U29434 (N_29434,N_29118,N_29236);
nor U29435 (N_29435,N_29004,N_29186);
xor U29436 (N_29436,N_29072,N_29141);
nand U29437 (N_29437,N_29049,N_29127);
and U29438 (N_29438,N_29201,N_29212);
nor U29439 (N_29439,N_29019,N_29066);
or U29440 (N_29440,N_29076,N_29074);
xnor U29441 (N_29441,N_29207,N_29172);
or U29442 (N_29442,N_29035,N_29016);
nand U29443 (N_29443,N_29123,N_29173);
nand U29444 (N_29444,N_29181,N_29247);
xor U29445 (N_29445,N_29166,N_29046);
and U29446 (N_29446,N_29129,N_29224);
nor U29447 (N_29447,N_29229,N_29037);
and U29448 (N_29448,N_29135,N_29243);
and U29449 (N_29449,N_29160,N_29099);
or U29450 (N_29450,N_29110,N_29107);
xnor U29451 (N_29451,N_29007,N_29116);
nand U29452 (N_29452,N_29167,N_29028);
and U29453 (N_29453,N_29018,N_29021);
and U29454 (N_29454,N_29062,N_29051);
or U29455 (N_29455,N_29206,N_29233);
xor U29456 (N_29456,N_29096,N_29231);
xnor U29457 (N_29457,N_29089,N_29150);
nor U29458 (N_29458,N_29077,N_29117);
nand U29459 (N_29459,N_29009,N_29082);
and U29460 (N_29460,N_29231,N_29047);
or U29461 (N_29461,N_29075,N_29071);
xor U29462 (N_29462,N_29096,N_29018);
or U29463 (N_29463,N_29159,N_29087);
nand U29464 (N_29464,N_29055,N_29117);
xnor U29465 (N_29465,N_29172,N_29058);
and U29466 (N_29466,N_29155,N_29228);
xor U29467 (N_29467,N_29174,N_29212);
xnor U29468 (N_29468,N_29099,N_29163);
and U29469 (N_29469,N_29082,N_29025);
and U29470 (N_29470,N_29076,N_29084);
and U29471 (N_29471,N_29160,N_29168);
nand U29472 (N_29472,N_29029,N_29058);
and U29473 (N_29473,N_29062,N_29031);
nor U29474 (N_29474,N_29224,N_29119);
and U29475 (N_29475,N_29143,N_29167);
nand U29476 (N_29476,N_29212,N_29192);
nor U29477 (N_29477,N_29087,N_29055);
and U29478 (N_29478,N_29127,N_29012);
and U29479 (N_29479,N_29161,N_29023);
nand U29480 (N_29480,N_29126,N_29207);
and U29481 (N_29481,N_29180,N_29208);
nand U29482 (N_29482,N_29149,N_29063);
nor U29483 (N_29483,N_29064,N_29042);
xor U29484 (N_29484,N_29082,N_29072);
xor U29485 (N_29485,N_29032,N_29203);
nand U29486 (N_29486,N_29009,N_29019);
xor U29487 (N_29487,N_29098,N_29068);
nor U29488 (N_29488,N_29012,N_29157);
and U29489 (N_29489,N_29116,N_29046);
or U29490 (N_29490,N_29040,N_29172);
and U29491 (N_29491,N_29117,N_29159);
or U29492 (N_29492,N_29172,N_29123);
or U29493 (N_29493,N_29094,N_29137);
and U29494 (N_29494,N_29003,N_29101);
xor U29495 (N_29495,N_29014,N_29075);
nand U29496 (N_29496,N_29003,N_29229);
nor U29497 (N_29497,N_29135,N_29026);
nor U29498 (N_29498,N_29229,N_29225);
nand U29499 (N_29499,N_29036,N_29029);
and U29500 (N_29500,N_29278,N_29284);
nand U29501 (N_29501,N_29488,N_29341);
nand U29502 (N_29502,N_29308,N_29429);
xor U29503 (N_29503,N_29280,N_29337);
nand U29504 (N_29504,N_29479,N_29371);
xnor U29505 (N_29505,N_29387,N_29362);
or U29506 (N_29506,N_29476,N_29426);
or U29507 (N_29507,N_29309,N_29264);
nor U29508 (N_29508,N_29345,N_29364);
xor U29509 (N_29509,N_29367,N_29305);
and U29510 (N_29510,N_29442,N_29296);
xnor U29511 (N_29511,N_29381,N_29303);
and U29512 (N_29512,N_29409,N_29462);
nand U29513 (N_29513,N_29433,N_29456);
xnor U29514 (N_29514,N_29434,N_29385);
nand U29515 (N_29515,N_29436,N_29487);
and U29516 (N_29516,N_29316,N_29317);
or U29517 (N_29517,N_29457,N_29472);
or U29518 (N_29518,N_29423,N_29389);
nor U29519 (N_29519,N_29422,N_29478);
nand U29520 (N_29520,N_29283,N_29333);
nor U29521 (N_29521,N_29412,N_29377);
and U29522 (N_29522,N_29289,N_29494);
or U29523 (N_29523,N_29304,N_29482);
or U29524 (N_29524,N_29467,N_29461);
and U29525 (N_29525,N_29495,N_29291);
and U29526 (N_29526,N_29307,N_29471);
nand U29527 (N_29527,N_29393,N_29483);
or U29528 (N_29528,N_29411,N_29342);
nor U29529 (N_29529,N_29300,N_29344);
or U29530 (N_29530,N_29297,N_29298);
and U29531 (N_29531,N_29282,N_29383);
or U29532 (N_29532,N_29469,N_29489);
xnor U29533 (N_29533,N_29392,N_29408);
nand U29534 (N_29534,N_29465,N_29491);
nand U29535 (N_29535,N_29336,N_29400);
nor U29536 (N_29536,N_29338,N_29349);
and U29537 (N_29537,N_29359,N_29398);
and U29538 (N_29538,N_29295,N_29390);
and U29539 (N_29539,N_29260,N_29499);
nand U29540 (N_29540,N_29481,N_29424);
nand U29541 (N_29541,N_29454,N_29447);
or U29542 (N_29542,N_29274,N_29375);
or U29543 (N_29543,N_29287,N_29370);
or U29544 (N_29544,N_29458,N_29276);
or U29545 (N_29545,N_29428,N_29437);
nor U29546 (N_29546,N_29379,N_29259);
and U29547 (N_29547,N_29380,N_29443);
and U29548 (N_29548,N_29480,N_29324);
nor U29549 (N_29549,N_29357,N_29313);
nand U29550 (N_29550,N_29281,N_29372);
xor U29551 (N_29551,N_29498,N_29477);
or U29552 (N_29552,N_29360,N_29258);
or U29553 (N_29553,N_29473,N_29493);
and U29554 (N_29554,N_29446,N_29431);
and U29555 (N_29555,N_29358,N_29413);
xor U29556 (N_29556,N_29331,N_29396);
nor U29557 (N_29557,N_29301,N_29374);
nor U29558 (N_29558,N_29451,N_29449);
nand U29559 (N_29559,N_29293,N_29382);
or U29560 (N_29560,N_29311,N_29352);
xnor U29561 (N_29561,N_29463,N_29397);
or U29562 (N_29562,N_29448,N_29438);
or U29563 (N_29563,N_29273,N_29266);
or U29564 (N_29564,N_29460,N_29497);
xnor U29565 (N_29565,N_29421,N_29290);
or U29566 (N_29566,N_29286,N_29302);
nor U29567 (N_29567,N_29319,N_29368);
or U29568 (N_29568,N_29415,N_29418);
and U29569 (N_29569,N_29350,N_29326);
and U29570 (N_29570,N_29470,N_29403);
and U29571 (N_29571,N_29348,N_29275);
nand U29572 (N_29572,N_29486,N_29288);
nand U29573 (N_29573,N_29254,N_29366);
xor U29574 (N_29574,N_29416,N_29420);
xor U29575 (N_29575,N_29262,N_29475);
or U29576 (N_29576,N_29328,N_29419);
xor U29577 (N_29577,N_29277,N_29373);
xor U29578 (N_29578,N_29255,N_29430);
xnor U29579 (N_29579,N_29490,N_29365);
or U29580 (N_29580,N_29312,N_29414);
nand U29581 (N_29581,N_29445,N_29363);
or U29582 (N_29582,N_29261,N_29285);
and U29583 (N_29583,N_29399,N_29452);
nand U29584 (N_29584,N_29492,N_29332);
or U29585 (N_29585,N_29455,N_29339);
nand U29586 (N_29586,N_29356,N_29444);
or U29587 (N_29587,N_29318,N_29484);
nand U29588 (N_29588,N_29417,N_29441);
and U29589 (N_29589,N_29315,N_29388);
nor U29590 (N_29590,N_29405,N_29346);
or U29591 (N_29591,N_29269,N_29395);
xor U29592 (N_29592,N_29485,N_29402);
and U29593 (N_29593,N_29340,N_29321);
or U29594 (N_29594,N_29453,N_29468);
nand U29595 (N_29595,N_29263,N_29253);
xnor U29596 (N_29596,N_29252,N_29268);
or U29597 (N_29597,N_29272,N_29320);
nor U29598 (N_29598,N_29427,N_29386);
nand U29599 (N_29599,N_29323,N_29270);
and U29600 (N_29600,N_29251,N_29292);
nand U29601 (N_29601,N_29322,N_29474);
or U29602 (N_29602,N_29353,N_29355);
xor U29603 (N_29603,N_29410,N_29330);
and U29604 (N_29604,N_29391,N_29351);
or U29605 (N_29605,N_29369,N_29384);
or U29606 (N_29606,N_29378,N_29394);
and U29607 (N_29607,N_29347,N_29354);
nor U29608 (N_29608,N_29325,N_29271);
nor U29609 (N_29609,N_29294,N_29256);
xnor U29610 (N_29610,N_29404,N_29439);
nor U29611 (N_29611,N_29334,N_29466);
nor U29612 (N_29612,N_29361,N_29440);
nor U29613 (N_29613,N_29407,N_29265);
and U29614 (N_29614,N_29327,N_29432);
nand U29615 (N_29615,N_29459,N_29450);
nand U29616 (N_29616,N_29314,N_29376);
xnor U29617 (N_29617,N_29267,N_29435);
nand U29618 (N_29618,N_29464,N_29306);
nand U29619 (N_29619,N_29343,N_29496);
nand U29620 (N_29620,N_29299,N_29335);
xor U29621 (N_29621,N_29257,N_29406);
nand U29622 (N_29622,N_29425,N_29401);
nand U29623 (N_29623,N_29329,N_29250);
and U29624 (N_29624,N_29310,N_29279);
or U29625 (N_29625,N_29309,N_29390);
nor U29626 (N_29626,N_29266,N_29440);
nor U29627 (N_29627,N_29461,N_29459);
xnor U29628 (N_29628,N_29451,N_29496);
and U29629 (N_29629,N_29314,N_29395);
nor U29630 (N_29630,N_29391,N_29284);
nand U29631 (N_29631,N_29283,N_29309);
nand U29632 (N_29632,N_29335,N_29326);
nor U29633 (N_29633,N_29490,N_29317);
or U29634 (N_29634,N_29281,N_29368);
nor U29635 (N_29635,N_29481,N_29313);
xor U29636 (N_29636,N_29438,N_29324);
xor U29637 (N_29637,N_29426,N_29283);
xor U29638 (N_29638,N_29366,N_29272);
or U29639 (N_29639,N_29485,N_29443);
and U29640 (N_29640,N_29359,N_29274);
or U29641 (N_29641,N_29302,N_29461);
and U29642 (N_29642,N_29454,N_29428);
and U29643 (N_29643,N_29402,N_29299);
and U29644 (N_29644,N_29446,N_29387);
xor U29645 (N_29645,N_29365,N_29257);
xor U29646 (N_29646,N_29312,N_29318);
nand U29647 (N_29647,N_29390,N_29330);
nor U29648 (N_29648,N_29316,N_29347);
nor U29649 (N_29649,N_29405,N_29260);
nor U29650 (N_29650,N_29256,N_29419);
or U29651 (N_29651,N_29304,N_29399);
or U29652 (N_29652,N_29437,N_29270);
or U29653 (N_29653,N_29394,N_29400);
or U29654 (N_29654,N_29336,N_29356);
nor U29655 (N_29655,N_29488,N_29428);
xor U29656 (N_29656,N_29307,N_29306);
and U29657 (N_29657,N_29349,N_29276);
or U29658 (N_29658,N_29313,N_29494);
nand U29659 (N_29659,N_29419,N_29284);
nor U29660 (N_29660,N_29348,N_29359);
and U29661 (N_29661,N_29491,N_29444);
nor U29662 (N_29662,N_29371,N_29496);
nor U29663 (N_29663,N_29443,N_29361);
and U29664 (N_29664,N_29305,N_29336);
xor U29665 (N_29665,N_29268,N_29384);
and U29666 (N_29666,N_29385,N_29440);
or U29667 (N_29667,N_29350,N_29494);
nand U29668 (N_29668,N_29386,N_29368);
xnor U29669 (N_29669,N_29453,N_29253);
xor U29670 (N_29670,N_29461,N_29498);
and U29671 (N_29671,N_29349,N_29392);
xor U29672 (N_29672,N_29260,N_29448);
or U29673 (N_29673,N_29417,N_29412);
nand U29674 (N_29674,N_29430,N_29471);
and U29675 (N_29675,N_29419,N_29336);
or U29676 (N_29676,N_29466,N_29483);
xnor U29677 (N_29677,N_29258,N_29330);
or U29678 (N_29678,N_29432,N_29264);
nand U29679 (N_29679,N_29377,N_29499);
and U29680 (N_29680,N_29264,N_29431);
or U29681 (N_29681,N_29408,N_29442);
xnor U29682 (N_29682,N_29417,N_29304);
or U29683 (N_29683,N_29437,N_29465);
nor U29684 (N_29684,N_29286,N_29356);
or U29685 (N_29685,N_29277,N_29348);
nand U29686 (N_29686,N_29419,N_29281);
xnor U29687 (N_29687,N_29306,N_29414);
and U29688 (N_29688,N_29491,N_29493);
nand U29689 (N_29689,N_29336,N_29446);
and U29690 (N_29690,N_29411,N_29493);
nand U29691 (N_29691,N_29360,N_29294);
nor U29692 (N_29692,N_29281,N_29342);
or U29693 (N_29693,N_29471,N_29294);
or U29694 (N_29694,N_29405,N_29341);
nand U29695 (N_29695,N_29429,N_29400);
or U29696 (N_29696,N_29254,N_29305);
and U29697 (N_29697,N_29489,N_29303);
and U29698 (N_29698,N_29407,N_29278);
nand U29699 (N_29699,N_29433,N_29340);
nand U29700 (N_29700,N_29383,N_29392);
xor U29701 (N_29701,N_29398,N_29393);
and U29702 (N_29702,N_29394,N_29365);
nor U29703 (N_29703,N_29286,N_29362);
nand U29704 (N_29704,N_29268,N_29479);
nor U29705 (N_29705,N_29396,N_29295);
nand U29706 (N_29706,N_29484,N_29268);
nand U29707 (N_29707,N_29458,N_29279);
nand U29708 (N_29708,N_29311,N_29443);
nand U29709 (N_29709,N_29459,N_29343);
nor U29710 (N_29710,N_29381,N_29457);
nand U29711 (N_29711,N_29300,N_29454);
and U29712 (N_29712,N_29349,N_29396);
or U29713 (N_29713,N_29286,N_29265);
or U29714 (N_29714,N_29335,N_29290);
nand U29715 (N_29715,N_29349,N_29322);
xor U29716 (N_29716,N_29314,N_29320);
or U29717 (N_29717,N_29477,N_29364);
and U29718 (N_29718,N_29365,N_29266);
xnor U29719 (N_29719,N_29336,N_29494);
nor U29720 (N_29720,N_29468,N_29299);
and U29721 (N_29721,N_29369,N_29375);
and U29722 (N_29722,N_29421,N_29334);
nand U29723 (N_29723,N_29399,N_29264);
and U29724 (N_29724,N_29390,N_29446);
nand U29725 (N_29725,N_29284,N_29480);
nand U29726 (N_29726,N_29391,N_29468);
nand U29727 (N_29727,N_29416,N_29422);
and U29728 (N_29728,N_29292,N_29408);
and U29729 (N_29729,N_29488,N_29251);
nand U29730 (N_29730,N_29344,N_29281);
nand U29731 (N_29731,N_29384,N_29381);
xnor U29732 (N_29732,N_29314,N_29419);
nand U29733 (N_29733,N_29416,N_29308);
nand U29734 (N_29734,N_29325,N_29498);
and U29735 (N_29735,N_29267,N_29465);
xor U29736 (N_29736,N_29266,N_29433);
nor U29737 (N_29737,N_29286,N_29290);
nand U29738 (N_29738,N_29323,N_29400);
nor U29739 (N_29739,N_29326,N_29437);
and U29740 (N_29740,N_29310,N_29345);
xor U29741 (N_29741,N_29400,N_29266);
and U29742 (N_29742,N_29277,N_29473);
nor U29743 (N_29743,N_29304,N_29276);
and U29744 (N_29744,N_29458,N_29355);
and U29745 (N_29745,N_29477,N_29388);
xnor U29746 (N_29746,N_29404,N_29270);
xor U29747 (N_29747,N_29406,N_29355);
nand U29748 (N_29748,N_29469,N_29343);
and U29749 (N_29749,N_29296,N_29266);
and U29750 (N_29750,N_29657,N_29566);
nor U29751 (N_29751,N_29679,N_29713);
xnor U29752 (N_29752,N_29707,N_29702);
nor U29753 (N_29753,N_29692,N_29530);
nor U29754 (N_29754,N_29511,N_29550);
or U29755 (N_29755,N_29584,N_29589);
or U29756 (N_29756,N_29529,N_29690);
nand U29757 (N_29757,N_29672,N_29634);
nor U29758 (N_29758,N_29606,N_29726);
or U29759 (N_29759,N_29581,N_29641);
nor U29760 (N_29760,N_29734,N_29723);
xnor U29761 (N_29761,N_29704,N_29663);
and U29762 (N_29762,N_29653,N_29555);
nand U29763 (N_29763,N_29677,N_29630);
and U29764 (N_29764,N_29515,N_29522);
and U29765 (N_29765,N_29727,N_29595);
nand U29766 (N_29766,N_29614,N_29632);
or U29767 (N_29767,N_29502,N_29536);
or U29768 (N_29768,N_29538,N_29739);
or U29769 (N_29769,N_29691,N_29615);
xnor U29770 (N_29770,N_29675,N_29639);
or U29771 (N_29771,N_29593,N_29527);
and U29772 (N_29772,N_29616,N_29701);
and U29773 (N_29773,N_29721,N_29735);
or U29774 (N_29774,N_29742,N_29728);
nand U29775 (N_29775,N_29700,N_29662);
nor U29776 (N_29776,N_29681,N_29666);
xor U29777 (N_29777,N_29596,N_29668);
or U29778 (N_29778,N_29516,N_29543);
and U29779 (N_29779,N_29580,N_29680);
and U29780 (N_29780,N_29558,N_29508);
nor U29781 (N_29781,N_29695,N_29733);
and U29782 (N_29782,N_29642,N_29740);
nor U29783 (N_29783,N_29711,N_29703);
nor U29784 (N_29784,N_29546,N_29505);
xor U29785 (N_29785,N_29590,N_29658);
or U29786 (N_29786,N_29521,N_29559);
or U29787 (N_29787,N_29732,N_29542);
or U29788 (N_29788,N_29561,N_29591);
or U29789 (N_29789,N_29725,N_29683);
xnor U29790 (N_29790,N_29510,N_29674);
nand U29791 (N_29791,N_29652,N_29665);
and U29792 (N_29792,N_29587,N_29729);
and U29793 (N_29793,N_29548,N_29715);
nand U29794 (N_29794,N_29688,N_29519);
nor U29795 (N_29795,N_29686,N_29537);
nand U29796 (N_29796,N_29601,N_29636);
nor U29797 (N_29797,N_29655,N_29592);
and U29798 (N_29798,N_29717,N_29583);
and U29799 (N_29799,N_29646,N_29608);
nor U29800 (N_29800,N_29556,N_29564);
or U29801 (N_29801,N_29718,N_29746);
nor U29802 (N_29802,N_29749,N_29562);
and U29803 (N_29803,N_29716,N_29607);
nor U29804 (N_29804,N_29597,N_29709);
and U29805 (N_29805,N_29619,N_29504);
nand U29806 (N_29806,N_29673,N_29545);
and U29807 (N_29807,N_29544,N_29647);
nor U29808 (N_29808,N_29605,N_29512);
nor U29809 (N_29809,N_29560,N_29637);
or U29810 (N_29810,N_29533,N_29551);
and U29811 (N_29811,N_29588,N_29617);
nand U29812 (N_29812,N_29626,N_29517);
nand U29813 (N_29813,N_29618,N_29500);
nand U29814 (N_29814,N_29730,N_29513);
and U29815 (N_29815,N_29603,N_29509);
nand U29816 (N_29816,N_29557,N_29549);
or U29817 (N_29817,N_29640,N_29693);
xor U29818 (N_29818,N_29660,N_29643);
nor U29819 (N_29819,N_29578,N_29623);
and U29820 (N_29820,N_29525,N_29722);
and U29821 (N_29821,N_29670,N_29567);
xnor U29822 (N_29822,N_29532,N_29667);
and U29823 (N_29823,N_29661,N_29585);
or U29824 (N_29824,N_29621,N_29633);
xnor U29825 (N_29825,N_29629,N_29696);
nor U29826 (N_29826,N_29547,N_29720);
or U29827 (N_29827,N_29523,N_29609);
or U29828 (N_29828,N_29697,N_29602);
nor U29829 (N_29829,N_29625,N_29599);
xor U29830 (N_29830,N_29503,N_29507);
nand U29831 (N_29831,N_29610,N_29654);
nor U29832 (N_29832,N_29671,N_29676);
or U29833 (N_29833,N_29649,N_29531);
and U29834 (N_29834,N_29689,N_29565);
or U29835 (N_29835,N_29612,N_29737);
or U29836 (N_29836,N_29520,N_29644);
nor U29837 (N_29837,N_29708,N_29645);
nand U29838 (N_29838,N_29540,N_29631);
or U29839 (N_29839,N_29628,N_29594);
or U29840 (N_29840,N_29659,N_29579);
nand U29841 (N_29841,N_29526,N_29620);
xor U29842 (N_29842,N_29600,N_29745);
or U29843 (N_29843,N_29685,N_29698);
nand U29844 (N_29844,N_29748,N_29743);
nor U29845 (N_29845,N_29714,N_29577);
or U29846 (N_29846,N_29534,N_29541);
and U29847 (N_29847,N_29747,N_29741);
nor U29848 (N_29848,N_29712,N_29694);
nor U29849 (N_29849,N_29575,N_29506);
nand U29850 (N_29850,N_29571,N_29611);
xnor U29851 (N_29851,N_29552,N_29651);
nand U29852 (N_29852,N_29604,N_29650);
xnor U29853 (N_29853,N_29572,N_29699);
nand U29854 (N_29854,N_29669,N_29687);
nand U29855 (N_29855,N_29731,N_29514);
nand U29856 (N_29856,N_29744,N_29568);
and U29857 (N_29857,N_29710,N_29656);
and U29858 (N_29858,N_29586,N_29518);
and U29859 (N_29859,N_29535,N_29570);
nor U29860 (N_29860,N_29719,N_29598);
xnor U29861 (N_29861,N_29705,N_29573);
xnor U29862 (N_29862,N_29622,N_29627);
or U29863 (N_29863,N_29706,N_29678);
xnor U29864 (N_29864,N_29664,N_29638);
and U29865 (N_29865,N_29635,N_29528);
nand U29866 (N_29866,N_29736,N_29501);
xnor U29867 (N_29867,N_29524,N_29553);
or U29868 (N_29868,N_29613,N_29738);
xnor U29869 (N_29869,N_29563,N_29582);
or U29870 (N_29870,N_29648,N_29684);
nand U29871 (N_29871,N_29682,N_29539);
xor U29872 (N_29872,N_29724,N_29574);
nand U29873 (N_29873,N_29576,N_29569);
nand U29874 (N_29874,N_29554,N_29624);
or U29875 (N_29875,N_29704,N_29669);
nor U29876 (N_29876,N_29610,N_29565);
nand U29877 (N_29877,N_29728,N_29714);
nand U29878 (N_29878,N_29571,N_29623);
nor U29879 (N_29879,N_29645,N_29733);
xnor U29880 (N_29880,N_29696,N_29522);
and U29881 (N_29881,N_29696,N_29654);
nor U29882 (N_29882,N_29530,N_29573);
and U29883 (N_29883,N_29731,N_29637);
and U29884 (N_29884,N_29709,N_29517);
and U29885 (N_29885,N_29504,N_29509);
nand U29886 (N_29886,N_29517,N_29614);
and U29887 (N_29887,N_29646,N_29664);
or U29888 (N_29888,N_29622,N_29552);
nor U29889 (N_29889,N_29599,N_29701);
and U29890 (N_29890,N_29677,N_29662);
or U29891 (N_29891,N_29705,N_29679);
nor U29892 (N_29892,N_29716,N_29711);
or U29893 (N_29893,N_29629,N_29713);
or U29894 (N_29894,N_29559,N_29535);
xnor U29895 (N_29895,N_29649,N_29538);
or U29896 (N_29896,N_29540,N_29564);
nor U29897 (N_29897,N_29561,N_29743);
and U29898 (N_29898,N_29742,N_29551);
nor U29899 (N_29899,N_29748,N_29699);
nor U29900 (N_29900,N_29566,N_29717);
nor U29901 (N_29901,N_29552,N_29522);
nand U29902 (N_29902,N_29503,N_29551);
nand U29903 (N_29903,N_29597,N_29595);
xnor U29904 (N_29904,N_29629,N_29548);
nand U29905 (N_29905,N_29694,N_29530);
nand U29906 (N_29906,N_29516,N_29650);
nand U29907 (N_29907,N_29714,N_29746);
and U29908 (N_29908,N_29718,N_29713);
nor U29909 (N_29909,N_29507,N_29684);
nand U29910 (N_29910,N_29739,N_29673);
nor U29911 (N_29911,N_29658,N_29572);
and U29912 (N_29912,N_29700,N_29523);
nor U29913 (N_29913,N_29639,N_29627);
nor U29914 (N_29914,N_29552,N_29631);
nand U29915 (N_29915,N_29607,N_29706);
nand U29916 (N_29916,N_29507,N_29607);
nand U29917 (N_29917,N_29697,N_29611);
nor U29918 (N_29918,N_29732,N_29684);
or U29919 (N_29919,N_29513,N_29592);
or U29920 (N_29920,N_29632,N_29606);
xnor U29921 (N_29921,N_29638,N_29651);
and U29922 (N_29922,N_29697,N_29711);
nand U29923 (N_29923,N_29609,N_29505);
and U29924 (N_29924,N_29632,N_29526);
and U29925 (N_29925,N_29504,N_29697);
nor U29926 (N_29926,N_29668,N_29576);
nand U29927 (N_29927,N_29644,N_29592);
and U29928 (N_29928,N_29731,N_29703);
and U29929 (N_29929,N_29686,N_29547);
nand U29930 (N_29930,N_29705,N_29724);
nand U29931 (N_29931,N_29685,N_29635);
and U29932 (N_29932,N_29597,N_29701);
or U29933 (N_29933,N_29649,N_29599);
and U29934 (N_29934,N_29654,N_29588);
nor U29935 (N_29935,N_29604,N_29515);
and U29936 (N_29936,N_29706,N_29649);
xnor U29937 (N_29937,N_29532,N_29617);
or U29938 (N_29938,N_29571,N_29659);
nand U29939 (N_29939,N_29671,N_29702);
and U29940 (N_29940,N_29665,N_29649);
or U29941 (N_29941,N_29725,N_29749);
nor U29942 (N_29942,N_29738,N_29557);
and U29943 (N_29943,N_29684,N_29558);
nor U29944 (N_29944,N_29515,N_29645);
xor U29945 (N_29945,N_29727,N_29665);
and U29946 (N_29946,N_29613,N_29588);
xor U29947 (N_29947,N_29527,N_29574);
and U29948 (N_29948,N_29661,N_29730);
and U29949 (N_29949,N_29521,N_29681);
and U29950 (N_29950,N_29506,N_29503);
or U29951 (N_29951,N_29695,N_29529);
nand U29952 (N_29952,N_29708,N_29715);
nor U29953 (N_29953,N_29586,N_29729);
nand U29954 (N_29954,N_29703,N_29696);
xnor U29955 (N_29955,N_29702,N_29637);
nand U29956 (N_29956,N_29704,N_29749);
or U29957 (N_29957,N_29715,N_29632);
xor U29958 (N_29958,N_29568,N_29607);
or U29959 (N_29959,N_29565,N_29663);
xor U29960 (N_29960,N_29653,N_29661);
and U29961 (N_29961,N_29502,N_29700);
nor U29962 (N_29962,N_29724,N_29681);
xor U29963 (N_29963,N_29594,N_29561);
nor U29964 (N_29964,N_29715,N_29636);
nand U29965 (N_29965,N_29606,N_29683);
nor U29966 (N_29966,N_29567,N_29683);
nor U29967 (N_29967,N_29628,N_29738);
or U29968 (N_29968,N_29576,N_29604);
or U29969 (N_29969,N_29620,N_29668);
nand U29970 (N_29970,N_29572,N_29720);
and U29971 (N_29971,N_29663,N_29712);
xnor U29972 (N_29972,N_29697,N_29724);
nand U29973 (N_29973,N_29575,N_29582);
and U29974 (N_29974,N_29560,N_29593);
and U29975 (N_29975,N_29695,N_29659);
nor U29976 (N_29976,N_29558,N_29650);
and U29977 (N_29977,N_29598,N_29553);
xor U29978 (N_29978,N_29621,N_29729);
or U29979 (N_29979,N_29516,N_29737);
or U29980 (N_29980,N_29577,N_29674);
nand U29981 (N_29981,N_29707,N_29571);
xnor U29982 (N_29982,N_29588,N_29667);
or U29983 (N_29983,N_29651,N_29543);
or U29984 (N_29984,N_29671,N_29746);
and U29985 (N_29985,N_29566,N_29691);
nor U29986 (N_29986,N_29504,N_29669);
xor U29987 (N_29987,N_29513,N_29745);
or U29988 (N_29988,N_29541,N_29590);
or U29989 (N_29989,N_29645,N_29650);
and U29990 (N_29990,N_29640,N_29500);
and U29991 (N_29991,N_29743,N_29626);
and U29992 (N_29992,N_29578,N_29678);
nor U29993 (N_29993,N_29523,N_29701);
nand U29994 (N_29994,N_29505,N_29640);
and U29995 (N_29995,N_29723,N_29731);
nor U29996 (N_29996,N_29576,N_29661);
or U29997 (N_29997,N_29557,N_29548);
xnor U29998 (N_29998,N_29618,N_29713);
and U29999 (N_29999,N_29546,N_29744);
and U30000 (N_30000,N_29866,N_29838);
xnor U30001 (N_30001,N_29917,N_29770);
and U30002 (N_30002,N_29831,N_29983);
xor U30003 (N_30003,N_29799,N_29950);
nor U30004 (N_30004,N_29891,N_29790);
nor U30005 (N_30005,N_29949,N_29852);
and U30006 (N_30006,N_29843,N_29875);
or U30007 (N_30007,N_29992,N_29754);
and U30008 (N_30008,N_29773,N_29892);
nor U30009 (N_30009,N_29925,N_29981);
or U30010 (N_30010,N_29819,N_29780);
xnor U30011 (N_30011,N_29970,N_29832);
nor U30012 (N_30012,N_29807,N_29812);
nand U30013 (N_30013,N_29862,N_29840);
nor U30014 (N_30014,N_29768,N_29873);
and U30015 (N_30015,N_29813,N_29967);
or U30016 (N_30016,N_29936,N_29800);
xnor U30017 (N_30017,N_29935,N_29913);
and U30018 (N_30018,N_29816,N_29869);
xor U30019 (N_30019,N_29764,N_29774);
and U30020 (N_30020,N_29872,N_29955);
and U30021 (N_30021,N_29995,N_29962);
xnor U30022 (N_30022,N_29779,N_29763);
or U30023 (N_30023,N_29814,N_29825);
and U30024 (N_30024,N_29788,N_29841);
and U30025 (N_30025,N_29857,N_29883);
xor U30026 (N_30026,N_29961,N_29853);
nor U30027 (N_30027,N_29829,N_29794);
nand U30028 (N_30028,N_29946,N_29987);
xnor U30029 (N_30029,N_29985,N_29751);
nor U30030 (N_30030,N_29923,N_29797);
xor U30031 (N_30031,N_29926,N_29876);
or U30032 (N_30032,N_29858,N_29885);
nand U30033 (N_30033,N_29954,N_29920);
xnor U30034 (N_30034,N_29821,N_29766);
xnor U30035 (N_30035,N_29999,N_29815);
nor U30036 (N_30036,N_29994,N_29906);
and U30037 (N_30037,N_29809,N_29998);
and U30038 (N_30038,N_29806,N_29752);
nand U30039 (N_30039,N_29842,N_29911);
and U30040 (N_30040,N_29945,N_29834);
or U30041 (N_30041,N_29856,N_29989);
xor U30042 (N_30042,N_29960,N_29966);
nand U30043 (N_30043,N_29976,N_29775);
or U30044 (N_30044,N_29896,N_29828);
xor U30045 (N_30045,N_29868,N_29783);
nor U30046 (N_30046,N_29924,N_29947);
nor U30047 (N_30047,N_29940,N_29756);
xnor U30048 (N_30048,N_29964,N_29824);
and U30049 (N_30049,N_29888,N_29881);
nand U30050 (N_30050,N_29982,N_29755);
xnor U30051 (N_30051,N_29953,N_29895);
nor U30052 (N_30052,N_29776,N_29948);
and U30053 (N_30053,N_29889,N_29943);
nand U30054 (N_30054,N_29811,N_29884);
and U30055 (N_30055,N_29965,N_29851);
xnor U30056 (N_30056,N_29956,N_29870);
or U30057 (N_30057,N_29772,N_29952);
nand U30058 (N_30058,N_29867,N_29951);
or U30059 (N_30059,N_29781,N_29786);
or U30060 (N_30060,N_29898,N_29972);
or U30061 (N_30061,N_29769,N_29904);
xnor U30062 (N_30062,N_29902,N_29863);
nand U30063 (N_30063,N_29930,N_29912);
nor U30064 (N_30064,N_29900,N_29878);
or U30065 (N_30065,N_29918,N_29777);
nand U30066 (N_30066,N_29931,N_29818);
and U30067 (N_30067,N_29791,N_29826);
or U30068 (N_30068,N_29975,N_29803);
nor U30069 (N_30069,N_29905,N_29986);
xnor U30070 (N_30070,N_29845,N_29977);
xor U30071 (N_30071,N_29796,N_29957);
xnor U30072 (N_30072,N_29919,N_29984);
or U30073 (N_30073,N_29785,N_29859);
xnor U30074 (N_30074,N_29890,N_29759);
xnor U30075 (N_30075,N_29808,N_29839);
and U30076 (N_30076,N_29929,N_29901);
nand U30077 (N_30077,N_29894,N_29877);
or U30078 (N_30078,N_29927,N_29810);
nand U30079 (N_30079,N_29789,N_29938);
nor U30080 (N_30080,N_29844,N_29849);
nand U30081 (N_30081,N_29830,N_29990);
nand U30082 (N_30082,N_29805,N_29980);
or U30083 (N_30083,N_29934,N_29916);
xor U30084 (N_30084,N_29823,N_29968);
xor U30085 (N_30085,N_29847,N_29941);
or U30086 (N_30086,N_29991,N_29903);
or U30087 (N_30087,N_29897,N_29793);
nand U30088 (N_30088,N_29871,N_29973);
and U30089 (N_30089,N_29874,N_29928);
nor U30090 (N_30090,N_29758,N_29795);
xnor U30091 (N_30091,N_29865,N_29753);
nand U30092 (N_30092,N_29932,N_29761);
or U30093 (N_30093,N_29864,N_29848);
nor U30094 (N_30094,N_29910,N_29939);
nor U30095 (N_30095,N_29978,N_29996);
and U30096 (N_30096,N_29979,N_29802);
and U30097 (N_30097,N_29778,N_29782);
nor U30098 (N_30098,N_29861,N_29988);
and U30099 (N_30099,N_29854,N_29762);
nor U30100 (N_30100,N_29907,N_29914);
or U30101 (N_30101,N_29909,N_29971);
and U30102 (N_30102,N_29792,N_29969);
and U30103 (N_30103,N_29942,N_29879);
or U30104 (N_30104,N_29750,N_29757);
and U30105 (N_30105,N_29963,N_29921);
and U30106 (N_30106,N_29798,N_29765);
nand U30107 (N_30107,N_29855,N_29837);
or U30108 (N_30108,N_29933,N_29827);
nand U30109 (N_30109,N_29922,N_29959);
and U30110 (N_30110,N_29822,N_29937);
nand U30111 (N_30111,N_29771,N_29801);
xor U30112 (N_30112,N_29997,N_29908);
xor U30113 (N_30113,N_29836,N_29817);
xor U30114 (N_30114,N_29833,N_29787);
nor U30115 (N_30115,N_29760,N_29993);
or U30116 (N_30116,N_29893,N_29899);
nor U30117 (N_30117,N_29880,N_29915);
nand U30118 (N_30118,N_29846,N_29887);
nor U30119 (N_30119,N_29882,N_29820);
nand U30120 (N_30120,N_29886,N_29944);
and U30121 (N_30121,N_29804,N_29850);
and U30122 (N_30122,N_29784,N_29958);
and U30123 (N_30123,N_29974,N_29767);
nand U30124 (N_30124,N_29835,N_29860);
and U30125 (N_30125,N_29838,N_29791);
or U30126 (N_30126,N_29846,N_29907);
or U30127 (N_30127,N_29843,N_29775);
nand U30128 (N_30128,N_29868,N_29821);
and U30129 (N_30129,N_29941,N_29771);
nor U30130 (N_30130,N_29980,N_29896);
xor U30131 (N_30131,N_29915,N_29850);
and U30132 (N_30132,N_29849,N_29881);
nand U30133 (N_30133,N_29795,N_29859);
nand U30134 (N_30134,N_29988,N_29828);
nand U30135 (N_30135,N_29980,N_29802);
nor U30136 (N_30136,N_29923,N_29935);
and U30137 (N_30137,N_29935,N_29770);
nand U30138 (N_30138,N_29844,N_29782);
and U30139 (N_30139,N_29855,N_29890);
or U30140 (N_30140,N_29862,N_29948);
and U30141 (N_30141,N_29753,N_29997);
nor U30142 (N_30142,N_29961,N_29839);
nand U30143 (N_30143,N_29814,N_29750);
and U30144 (N_30144,N_29798,N_29978);
and U30145 (N_30145,N_29980,N_29905);
nand U30146 (N_30146,N_29763,N_29842);
nand U30147 (N_30147,N_29847,N_29758);
and U30148 (N_30148,N_29764,N_29767);
or U30149 (N_30149,N_29987,N_29953);
or U30150 (N_30150,N_29776,N_29848);
xnor U30151 (N_30151,N_29894,N_29977);
nand U30152 (N_30152,N_29895,N_29791);
nor U30153 (N_30153,N_29914,N_29956);
xnor U30154 (N_30154,N_29867,N_29783);
xor U30155 (N_30155,N_29808,N_29966);
nor U30156 (N_30156,N_29988,N_29836);
or U30157 (N_30157,N_29925,N_29938);
xnor U30158 (N_30158,N_29945,N_29920);
and U30159 (N_30159,N_29897,N_29866);
or U30160 (N_30160,N_29991,N_29883);
nand U30161 (N_30161,N_29766,N_29977);
nand U30162 (N_30162,N_29792,N_29927);
xnor U30163 (N_30163,N_29769,N_29812);
xnor U30164 (N_30164,N_29969,N_29835);
xnor U30165 (N_30165,N_29840,N_29777);
or U30166 (N_30166,N_29892,N_29996);
nand U30167 (N_30167,N_29877,N_29988);
nand U30168 (N_30168,N_29810,N_29850);
or U30169 (N_30169,N_29956,N_29852);
xnor U30170 (N_30170,N_29932,N_29842);
nand U30171 (N_30171,N_29927,N_29958);
xor U30172 (N_30172,N_29764,N_29957);
and U30173 (N_30173,N_29780,N_29944);
or U30174 (N_30174,N_29939,N_29771);
nand U30175 (N_30175,N_29933,N_29794);
nor U30176 (N_30176,N_29821,N_29893);
nor U30177 (N_30177,N_29751,N_29939);
and U30178 (N_30178,N_29809,N_29966);
and U30179 (N_30179,N_29945,N_29889);
or U30180 (N_30180,N_29982,N_29816);
and U30181 (N_30181,N_29761,N_29928);
nand U30182 (N_30182,N_29771,N_29940);
nor U30183 (N_30183,N_29892,N_29872);
nand U30184 (N_30184,N_29862,N_29996);
or U30185 (N_30185,N_29800,N_29921);
or U30186 (N_30186,N_29953,N_29954);
nor U30187 (N_30187,N_29767,N_29917);
nand U30188 (N_30188,N_29981,N_29831);
or U30189 (N_30189,N_29987,N_29788);
nor U30190 (N_30190,N_29885,N_29941);
nor U30191 (N_30191,N_29949,N_29874);
nor U30192 (N_30192,N_29822,N_29899);
and U30193 (N_30193,N_29973,N_29832);
and U30194 (N_30194,N_29899,N_29849);
or U30195 (N_30195,N_29853,N_29931);
nand U30196 (N_30196,N_29973,N_29960);
or U30197 (N_30197,N_29998,N_29864);
and U30198 (N_30198,N_29953,N_29923);
and U30199 (N_30199,N_29902,N_29776);
nand U30200 (N_30200,N_29768,N_29964);
and U30201 (N_30201,N_29961,N_29999);
and U30202 (N_30202,N_29842,N_29940);
or U30203 (N_30203,N_29841,N_29879);
xor U30204 (N_30204,N_29993,N_29906);
xor U30205 (N_30205,N_29943,N_29867);
nand U30206 (N_30206,N_29764,N_29917);
nand U30207 (N_30207,N_29777,N_29992);
and U30208 (N_30208,N_29948,N_29789);
and U30209 (N_30209,N_29983,N_29754);
or U30210 (N_30210,N_29982,N_29870);
or U30211 (N_30211,N_29811,N_29969);
nor U30212 (N_30212,N_29806,N_29944);
and U30213 (N_30213,N_29867,N_29821);
xnor U30214 (N_30214,N_29984,N_29960);
xor U30215 (N_30215,N_29990,N_29850);
nor U30216 (N_30216,N_29826,N_29772);
and U30217 (N_30217,N_29815,N_29985);
and U30218 (N_30218,N_29909,N_29876);
and U30219 (N_30219,N_29988,N_29814);
xnor U30220 (N_30220,N_29971,N_29878);
nor U30221 (N_30221,N_29983,N_29905);
or U30222 (N_30222,N_29795,N_29861);
xor U30223 (N_30223,N_29941,N_29958);
and U30224 (N_30224,N_29926,N_29786);
nor U30225 (N_30225,N_29768,N_29972);
nor U30226 (N_30226,N_29825,N_29882);
nand U30227 (N_30227,N_29920,N_29805);
nand U30228 (N_30228,N_29780,N_29784);
or U30229 (N_30229,N_29814,N_29911);
nor U30230 (N_30230,N_29908,N_29922);
nand U30231 (N_30231,N_29889,N_29816);
nor U30232 (N_30232,N_29871,N_29820);
or U30233 (N_30233,N_29768,N_29934);
or U30234 (N_30234,N_29860,N_29995);
and U30235 (N_30235,N_29834,N_29756);
nor U30236 (N_30236,N_29818,N_29800);
nor U30237 (N_30237,N_29792,N_29891);
and U30238 (N_30238,N_29822,N_29974);
or U30239 (N_30239,N_29994,N_29929);
nand U30240 (N_30240,N_29771,N_29832);
or U30241 (N_30241,N_29832,N_29852);
or U30242 (N_30242,N_29833,N_29898);
nand U30243 (N_30243,N_29818,N_29975);
xor U30244 (N_30244,N_29849,N_29839);
and U30245 (N_30245,N_29966,N_29835);
nand U30246 (N_30246,N_29765,N_29838);
and U30247 (N_30247,N_29778,N_29967);
nor U30248 (N_30248,N_29805,N_29867);
or U30249 (N_30249,N_29990,N_29996);
nand U30250 (N_30250,N_30128,N_30241);
or U30251 (N_30251,N_30106,N_30169);
or U30252 (N_30252,N_30129,N_30055);
nor U30253 (N_30253,N_30238,N_30236);
nor U30254 (N_30254,N_30138,N_30047);
or U30255 (N_30255,N_30109,N_30148);
xor U30256 (N_30256,N_30090,N_30030);
nand U30257 (N_30257,N_30020,N_30174);
nand U30258 (N_30258,N_30065,N_30078);
xnor U30259 (N_30259,N_30134,N_30125);
or U30260 (N_30260,N_30146,N_30019);
nand U30261 (N_30261,N_30100,N_30122);
or U30262 (N_30262,N_30203,N_30028);
nand U30263 (N_30263,N_30082,N_30229);
and U30264 (N_30264,N_30080,N_30156);
or U30265 (N_30265,N_30123,N_30194);
nand U30266 (N_30266,N_30231,N_30186);
or U30267 (N_30267,N_30058,N_30097);
or U30268 (N_30268,N_30176,N_30165);
and U30269 (N_30269,N_30230,N_30042);
and U30270 (N_30270,N_30151,N_30101);
or U30271 (N_30271,N_30223,N_30215);
nand U30272 (N_30272,N_30202,N_30222);
and U30273 (N_30273,N_30112,N_30064);
nand U30274 (N_30274,N_30089,N_30029);
nor U30275 (N_30275,N_30168,N_30037);
and U30276 (N_30276,N_30027,N_30031);
and U30277 (N_30277,N_30085,N_30152);
and U30278 (N_30278,N_30017,N_30224);
xor U30279 (N_30279,N_30088,N_30135);
nor U30280 (N_30280,N_30188,N_30095);
xor U30281 (N_30281,N_30225,N_30197);
nor U30282 (N_30282,N_30103,N_30012);
nor U30283 (N_30283,N_30192,N_30150);
or U30284 (N_30284,N_30113,N_30048);
xnor U30285 (N_30285,N_30136,N_30161);
xnor U30286 (N_30286,N_30071,N_30092);
nand U30287 (N_30287,N_30116,N_30121);
nor U30288 (N_30288,N_30118,N_30235);
nor U30289 (N_30289,N_30158,N_30093);
and U30290 (N_30290,N_30084,N_30057);
nor U30291 (N_30291,N_30201,N_30008);
nand U30292 (N_30292,N_30204,N_30043);
or U30293 (N_30293,N_30066,N_30119);
nor U30294 (N_30294,N_30040,N_30033);
nand U30295 (N_30295,N_30175,N_30131);
nand U30296 (N_30296,N_30217,N_30180);
xor U30297 (N_30297,N_30178,N_30007);
xor U30298 (N_30298,N_30233,N_30021);
nor U30299 (N_30299,N_30177,N_30243);
or U30300 (N_30300,N_30210,N_30115);
or U30301 (N_30301,N_30081,N_30034);
nand U30302 (N_30302,N_30004,N_30039);
or U30303 (N_30303,N_30181,N_30237);
and U30304 (N_30304,N_30209,N_30145);
or U30305 (N_30305,N_30214,N_30227);
xor U30306 (N_30306,N_30193,N_30107);
nor U30307 (N_30307,N_30132,N_30036);
and U30308 (N_30308,N_30102,N_30144);
or U30309 (N_30309,N_30137,N_30218);
xnor U30310 (N_30310,N_30014,N_30173);
xnor U30311 (N_30311,N_30157,N_30244);
and U30312 (N_30312,N_30091,N_30025);
nand U30313 (N_30313,N_30035,N_30022);
or U30314 (N_30314,N_30044,N_30130);
nor U30315 (N_30315,N_30154,N_30094);
and U30316 (N_30316,N_30075,N_30163);
nor U30317 (N_30317,N_30069,N_30179);
nor U30318 (N_30318,N_30005,N_30232);
or U30319 (N_30319,N_30024,N_30247);
nand U30320 (N_30320,N_30032,N_30054);
xnor U30321 (N_30321,N_30073,N_30006);
nor U30322 (N_30322,N_30207,N_30001);
nand U30323 (N_30323,N_30205,N_30219);
or U30324 (N_30324,N_30234,N_30052);
or U30325 (N_30325,N_30242,N_30068);
and U30326 (N_30326,N_30041,N_30162);
or U30327 (N_30327,N_30059,N_30086);
xor U30328 (N_30328,N_30167,N_30117);
nor U30329 (N_30329,N_30221,N_30015);
and U30330 (N_30330,N_30184,N_30003);
or U30331 (N_30331,N_30228,N_30002);
nand U30332 (N_30332,N_30142,N_30038);
nor U30333 (N_30333,N_30139,N_30171);
nor U30334 (N_30334,N_30240,N_30198);
nor U30335 (N_30335,N_30147,N_30170);
xnor U30336 (N_30336,N_30124,N_30143);
or U30337 (N_30337,N_30099,N_30083);
nand U30338 (N_30338,N_30016,N_30245);
nand U30339 (N_30339,N_30062,N_30049);
and U30340 (N_30340,N_30190,N_30182);
nand U30341 (N_30341,N_30098,N_30200);
or U30342 (N_30342,N_30216,N_30220);
and U30343 (N_30343,N_30189,N_30000);
xor U30344 (N_30344,N_30056,N_30072);
nor U30345 (N_30345,N_30160,N_30166);
or U30346 (N_30346,N_30013,N_30191);
nand U30347 (N_30347,N_30110,N_30213);
xnor U30348 (N_30348,N_30023,N_30141);
nand U30349 (N_30349,N_30249,N_30239);
or U30350 (N_30350,N_30153,N_30120);
and U30351 (N_30351,N_30104,N_30155);
nor U30352 (N_30352,N_30053,N_30076);
xnor U30353 (N_30353,N_30159,N_30140);
and U30354 (N_30354,N_30070,N_30010);
or U30355 (N_30355,N_30087,N_30195);
or U30356 (N_30356,N_30108,N_30111);
or U30357 (N_30357,N_30067,N_30050);
and U30358 (N_30358,N_30096,N_30060);
or U30359 (N_30359,N_30126,N_30061);
xor U30360 (N_30360,N_30105,N_30208);
nand U30361 (N_30361,N_30009,N_30026);
nand U30362 (N_30362,N_30114,N_30248);
nand U30363 (N_30363,N_30077,N_30212);
or U30364 (N_30364,N_30187,N_30199);
nand U30365 (N_30365,N_30079,N_30183);
or U30366 (N_30366,N_30127,N_30185);
and U30367 (N_30367,N_30172,N_30226);
nor U30368 (N_30368,N_30018,N_30133);
nand U30369 (N_30369,N_30246,N_30164);
or U30370 (N_30370,N_30149,N_30206);
xor U30371 (N_30371,N_30211,N_30063);
nand U30372 (N_30372,N_30045,N_30046);
and U30373 (N_30373,N_30196,N_30051);
or U30374 (N_30374,N_30011,N_30074);
xnor U30375 (N_30375,N_30103,N_30224);
or U30376 (N_30376,N_30228,N_30231);
nor U30377 (N_30377,N_30249,N_30152);
or U30378 (N_30378,N_30132,N_30198);
nand U30379 (N_30379,N_30082,N_30128);
nand U30380 (N_30380,N_30078,N_30050);
and U30381 (N_30381,N_30078,N_30021);
nor U30382 (N_30382,N_30102,N_30219);
and U30383 (N_30383,N_30006,N_30232);
or U30384 (N_30384,N_30196,N_30218);
or U30385 (N_30385,N_30195,N_30019);
nor U30386 (N_30386,N_30112,N_30005);
nand U30387 (N_30387,N_30165,N_30020);
xnor U30388 (N_30388,N_30019,N_30067);
and U30389 (N_30389,N_30128,N_30105);
or U30390 (N_30390,N_30015,N_30008);
nand U30391 (N_30391,N_30178,N_30242);
xor U30392 (N_30392,N_30024,N_30112);
nor U30393 (N_30393,N_30046,N_30193);
and U30394 (N_30394,N_30160,N_30110);
nor U30395 (N_30395,N_30083,N_30169);
and U30396 (N_30396,N_30026,N_30047);
or U30397 (N_30397,N_30067,N_30152);
nor U30398 (N_30398,N_30052,N_30189);
and U30399 (N_30399,N_30152,N_30209);
nand U30400 (N_30400,N_30109,N_30226);
or U30401 (N_30401,N_30017,N_30170);
nand U30402 (N_30402,N_30143,N_30247);
xnor U30403 (N_30403,N_30112,N_30228);
nand U30404 (N_30404,N_30177,N_30013);
nor U30405 (N_30405,N_30071,N_30226);
xnor U30406 (N_30406,N_30168,N_30044);
or U30407 (N_30407,N_30052,N_30113);
xor U30408 (N_30408,N_30243,N_30141);
or U30409 (N_30409,N_30169,N_30097);
or U30410 (N_30410,N_30210,N_30223);
nor U30411 (N_30411,N_30036,N_30042);
xnor U30412 (N_30412,N_30197,N_30105);
and U30413 (N_30413,N_30195,N_30101);
xor U30414 (N_30414,N_30122,N_30043);
and U30415 (N_30415,N_30140,N_30127);
or U30416 (N_30416,N_30009,N_30222);
xnor U30417 (N_30417,N_30236,N_30116);
nor U30418 (N_30418,N_30181,N_30001);
nor U30419 (N_30419,N_30208,N_30038);
nand U30420 (N_30420,N_30172,N_30146);
and U30421 (N_30421,N_30186,N_30028);
and U30422 (N_30422,N_30104,N_30244);
nand U30423 (N_30423,N_30111,N_30002);
nor U30424 (N_30424,N_30112,N_30179);
and U30425 (N_30425,N_30235,N_30116);
and U30426 (N_30426,N_30146,N_30065);
nand U30427 (N_30427,N_30068,N_30041);
and U30428 (N_30428,N_30195,N_30102);
or U30429 (N_30429,N_30088,N_30232);
xor U30430 (N_30430,N_30083,N_30201);
nand U30431 (N_30431,N_30151,N_30055);
and U30432 (N_30432,N_30205,N_30075);
or U30433 (N_30433,N_30207,N_30125);
or U30434 (N_30434,N_30148,N_30237);
or U30435 (N_30435,N_30065,N_30216);
nor U30436 (N_30436,N_30022,N_30237);
nor U30437 (N_30437,N_30223,N_30068);
nor U30438 (N_30438,N_30041,N_30109);
or U30439 (N_30439,N_30072,N_30095);
xnor U30440 (N_30440,N_30201,N_30204);
xnor U30441 (N_30441,N_30105,N_30009);
and U30442 (N_30442,N_30105,N_30050);
or U30443 (N_30443,N_30093,N_30126);
nand U30444 (N_30444,N_30237,N_30037);
nor U30445 (N_30445,N_30090,N_30102);
or U30446 (N_30446,N_30191,N_30040);
and U30447 (N_30447,N_30143,N_30137);
or U30448 (N_30448,N_30082,N_30073);
xor U30449 (N_30449,N_30083,N_30094);
nand U30450 (N_30450,N_30144,N_30186);
or U30451 (N_30451,N_30153,N_30048);
xor U30452 (N_30452,N_30092,N_30057);
xor U30453 (N_30453,N_30180,N_30024);
nor U30454 (N_30454,N_30045,N_30004);
xor U30455 (N_30455,N_30178,N_30183);
and U30456 (N_30456,N_30207,N_30235);
xnor U30457 (N_30457,N_30229,N_30149);
nand U30458 (N_30458,N_30048,N_30011);
nand U30459 (N_30459,N_30180,N_30096);
and U30460 (N_30460,N_30000,N_30233);
nand U30461 (N_30461,N_30132,N_30235);
nand U30462 (N_30462,N_30237,N_30034);
or U30463 (N_30463,N_30085,N_30141);
xor U30464 (N_30464,N_30105,N_30221);
and U30465 (N_30465,N_30227,N_30131);
or U30466 (N_30466,N_30027,N_30109);
and U30467 (N_30467,N_30129,N_30068);
and U30468 (N_30468,N_30120,N_30191);
or U30469 (N_30469,N_30184,N_30015);
and U30470 (N_30470,N_30168,N_30150);
nand U30471 (N_30471,N_30129,N_30099);
nand U30472 (N_30472,N_30114,N_30215);
and U30473 (N_30473,N_30012,N_30238);
nor U30474 (N_30474,N_30154,N_30157);
nor U30475 (N_30475,N_30201,N_30220);
xor U30476 (N_30476,N_30176,N_30084);
xnor U30477 (N_30477,N_30121,N_30013);
xor U30478 (N_30478,N_30117,N_30099);
or U30479 (N_30479,N_30050,N_30107);
nand U30480 (N_30480,N_30059,N_30037);
xor U30481 (N_30481,N_30102,N_30122);
or U30482 (N_30482,N_30126,N_30156);
nor U30483 (N_30483,N_30238,N_30214);
nor U30484 (N_30484,N_30206,N_30037);
nor U30485 (N_30485,N_30240,N_30026);
xnor U30486 (N_30486,N_30133,N_30142);
or U30487 (N_30487,N_30007,N_30008);
nand U30488 (N_30488,N_30134,N_30129);
nor U30489 (N_30489,N_30178,N_30228);
and U30490 (N_30490,N_30161,N_30162);
and U30491 (N_30491,N_30003,N_30241);
and U30492 (N_30492,N_30194,N_30177);
or U30493 (N_30493,N_30179,N_30050);
xnor U30494 (N_30494,N_30027,N_30069);
xnor U30495 (N_30495,N_30042,N_30203);
nand U30496 (N_30496,N_30142,N_30209);
and U30497 (N_30497,N_30156,N_30134);
nor U30498 (N_30498,N_30002,N_30140);
nand U30499 (N_30499,N_30074,N_30077);
xnor U30500 (N_30500,N_30331,N_30262);
nor U30501 (N_30501,N_30329,N_30430);
xor U30502 (N_30502,N_30404,N_30441);
nor U30503 (N_30503,N_30377,N_30333);
or U30504 (N_30504,N_30324,N_30270);
nor U30505 (N_30505,N_30408,N_30350);
xnor U30506 (N_30506,N_30337,N_30474);
nor U30507 (N_30507,N_30315,N_30269);
or U30508 (N_30508,N_30473,N_30436);
nor U30509 (N_30509,N_30462,N_30274);
or U30510 (N_30510,N_30318,N_30424);
and U30511 (N_30511,N_30470,N_30385);
nand U30512 (N_30512,N_30364,N_30412);
xor U30513 (N_30513,N_30493,N_30427);
nand U30514 (N_30514,N_30375,N_30479);
nand U30515 (N_30515,N_30252,N_30456);
xor U30516 (N_30516,N_30384,N_30458);
xor U30517 (N_30517,N_30278,N_30343);
xor U30518 (N_30518,N_30344,N_30486);
nand U30519 (N_30519,N_30332,N_30299);
and U30520 (N_30520,N_30438,N_30292);
or U30521 (N_30521,N_30279,N_30357);
xnor U30522 (N_30522,N_30472,N_30300);
xnor U30523 (N_30523,N_30446,N_30354);
nor U30524 (N_30524,N_30314,N_30319);
and U30525 (N_30525,N_30437,N_30434);
xnor U30526 (N_30526,N_30416,N_30305);
and U30527 (N_30527,N_30448,N_30328);
or U30528 (N_30528,N_30353,N_30256);
and U30529 (N_30529,N_30302,N_30263);
nand U30530 (N_30530,N_30330,N_30449);
xor U30531 (N_30531,N_30457,N_30264);
or U30532 (N_30532,N_30372,N_30445);
xnor U30533 (N_30533,N_30414,N_30310);
nand U30534 (N_30534,N_30466,N_30387);
nand U30535 (N_30535,N_30351,N_30494);
nand U30536 (N_30536,N_30442,N_30499);
nor U30537 (N_30537,N_30272,N_30439);
nor U30538 (N_30538,N_30275,N_30400);
nand U30539 (N_30539,N_30386,N_30482);
or U30540 (N_30540,N_30476,N_30428);
nor U30541 (N_30541,N_30397,N_30451);
xor U30542 (N_30542,N_30268,N_30266);
nor U30543 (N_30543,N_30382,N_30356);
or U30544 (N_30544,N_30379,N_30309);
xnor U30545 (N_30545,N_30260,N_30368);
nor U30546 (N_30546,N_30392,N_30471);
nor U30547 (N_30547,N_30429,N_30413);
nor U30548 (N_30548,N_30398,N_30496);
or U30549 (N_30549,N_30267,N_30423);
or U30550 (N_30550,N_30338,N_30317);
xor U30551 (N_30551,N_30468,N_30421);
nand U30552 (N_30552,N_30396,N_30401);
nand U30553 (N_30553,N_30406,N_30326);
xnor U30554 (N_30554,N_30453,N_30322);
or U30555 (N_30555,N_30461,N_30321);
and U30556 (N_30556,N_30422,N_30383);
nor U30557 (N_30557,N_30261,N_30289);
and U30558 (N_30558,N_30452,N_30459);
or U30559 (N_30559,N_30367,N_30447);
xor U30560 (N_30560,N_30286,N_30417);
and U30561 (N_30561,N_30298,N_30435);
xor U30562 (N_30562,N_30373,N_30498);
and U30563 (N_30563,N_30376,N_30280);
nand U30564 (N_30564,N_30371,N_30355);
nor U30565 (N_30565,N_30454,N_30378);
xor U30566 (N_30566,N_30480,N_30464);
or U30567 (N_30567,N_30399,N_30402);
and U30568 (N_30568,N_30250,N_30380);
nor U30569 (N_30569,N_30358,N_30475);
nor U30570 (N_30570,N_30362,N_30393);
nor U30571 (N_30571,N_30405,N_30258);
and U30572 (N_30572,N_30418,N_30483);
and U30573 (N_30573,N_30293,N_30285);
xor U30574 (N_30574,N_30254,N_30395);
nor U30575 (N_30575,N_30361,N_30259);
xor U30576 (N_30576,N_30455,N_30487);
nand U30577 (N_30577,N_30349,N_30391);
xnor U30578 (N_30578,N_30444,N_30359);
nand U30579 (N_30579,N_30478,N_30463);
or U30580 (N_30580,N_30291,N_30295);
nor U30581 (N_30581,N_30307,N_30410);
nand U30582 (N_30582,N_30335,N_30346);
nand U30583 (N_30583,N_30273,N_30495);
or U30584 (N_30584,N_30497,N_30450);
nand U30585 (N_30585,N_30255,N_30419);
nand U30586 (N_30586,N_30325,N_30374);
nand U30587 (N_30587,N_30323,N_30334);
or U30588 (N_30588,N_30320,N_30342);
nand U30589 (N_30589,N_30488,N_30296);
and U30590 (N_30590,N_30303,N_30431);
or U30591 (N_30591,N_30257,N_30363);
xor U30592 (N_30592,N_30403,N_30366);
or U30593 (N_30593,N_30369,N_30433);
nand U30594 (N_30594,N_30301,N_30460);
nand U30595 (N_30595,N_30284,N_30306);
and U30596 (N_30596,N_30253,N_30415);
nor U30597 (N_30597,N_30304,N_30420);
or U30598 (N_30598,N_30316,N_30282);
and U30599 (N_30599,N_30288,N_30347);
nor U30600 (N_30600,N_30465,N_30389);
or U30601 (N_30601,N_30443,N_30283);
xor U30602 (N_30602,N_30492,N_30481);
nand U30603 (N_30603,N_30271,N_30348);
nor U30604 (N_30604,N_30265,N_30360);
nand U30605 (N_30605,N_30341,N_30440);
nor U30606 (N_30606,N_30425,N_30411);
nor U30607 (N_30607,N_30312,N_30491);
or U30608 (N_30608,N_30340,N_30345);
xor U30609 (N_30609,N_30313,N_30251);
or U30610 (N_30610,N_30477,N_30394);
nor U30611 (N_30611,N_30281,N_30409);
and U30612 (N_30612,N_30365,N_30484);
nor U30613 (N_30613,N_30297,N_30388);
and U30614 (N_30614,N_30336,N_30381);
or U30615 (N_30615,N_30390,N_30339);
and U30616 (N_30616,N_30469,N_30276);
and U30617 (N_30617,N_30290,N_30352);
nor U30618 (N_30618,N_30426,N_30370);
nand U30619 (N_30619,N_30277,N_30467);
xor U30620 (N_30620,N_30407,N_30489);
and U30621 (N_30621,N_30311,N_30294);
and U30622 (N_30622,N_30490,N_30485);
nand U30623 (N_30623,N_30287,N_30432);
and U30624 (N_30624,N_30308,N_30327);
or U30625 (N_30625,N_30486,N_30324);
xor U30626 (N_30626,N_30336,N_30422);
or U30627 (N_30627,N_30364,N_30401);
and U30628 (N_30628,N_30326,N_30342);
nand U30629 (N_30629,N_30496,N_30261);
or U30630 (N_30630,N_30447,N_30490);
nor U30631 (N_30631,N_30478,N_30292);
and U30632 (N_30632,N_30308,N_30426);
nand U30633 (N_30633,N_30452,N_30473);
and U30634 (N_30634,N_30317,N_30409);
or U30635 (N_30635,N_30292,N_30355);
or U30636 (N_30636,N_30294,N_30316);
and U30637 (N_30637,N_30386,N_30490);
or U30638 (N_30638,N_30264,N_30272);
nor U30639 (N_30639,N_30485,N_30468);
xor U30640 (N_30640,N_30427,N_30352);
xnor U30641 (N_30641,N_30487,N_30430);
nor U30642 (N_30642,N_30391,N_30412);
xor U30643 (N_30643,N_30486,N_30294);
and U30644 (N_30644,N_30289,N_30363);
xnor U30645 (N_30645,N_30375,N_30485);
nand U30646 (N_30646,N_30274,N_30298);
or U30647 (N_30647,N_30474,N_30275);
and U30648 (N_30648,N_30483,N_30409);
and U30649 (N_30649,N_30314,N_30320);
nand U30650 (N_30650,N_30381,N_30434);
or U30651 (N_30651,N_30456,N_30309);
nand U30652 (N_30652,N_30296,N_30465);
nand U30653 (N_30653,N_30451,N_30265);
or U30654 (N_30654,N_30380,N_30474);
or U30655 (N_30655,N_30381,N_30382);
and U30656 (N_30656,N_30493,N_30347);
and U30657 (N_30657,N_30439,N_30314);
or U30658 (N_30658,N_30311,N_30319);
or U30659 (N_30659,N_30392,N_30487);
or U30660 (N_30660,N_30386,N_30383);
or U30661 (N_30661,N_30374,N_30420);
nor U30662 (N_30662,N_30251,N_30264);
and U30663 (N_30663,N_30477,N_30388);
or U30664 (N_30664,N_30277,N_30321);
xor U30665 (N_30665,N_30367,N_30269);
nand U30666 (N_30666,N_30366,N_30398);
nand U30667 (N_30667,N_30348,N_30384);
and U30668 (N_30668,N_30375,N_30372);
or U30669 (N_30669,N_30398,N_30263);
nand U30670 (N_30670,N_30280,N_30359);
nor U30671 (N_30671,N_30427,N_30261);
nor U30672 (N_30672,N_30396,N_30402);
nand U30673 (N_30673,N_30332,N_30267);
xnor U30674 (N_30674,N_30341,N_30297);
or U30675 (N_30675,N_30486,N_30340);
nor U30676 (N_30676,N_30415,N_30422);
or U30677 (N_30677,N_30481,N_30424);
nor U30678 (N_30678,N_30404,N_30257);
nand U30679 (N_30679,N_30454,N_30476);
xnor U30680 (N_30680,N_30450,N_30440);
and U30681 (N_30681,N_30405,N_30251);
or U30682 (N_30682,N_30470,N_30253);
or U30683 (N_30683,N_30303,N_30413);
nand U30684 (N_30684,N_30338,N_30495);
and U30685 (N_30685,N_30384,N_30275);
and U30686 (N_30686,N_30269,N_30277);
or U30687 (N_30687,N_30335,N_30363);
nand U30688 (N_30688,N_30294,N_30428);
nor U30689 (N_30689,N_30443,N_30405);
nand U30690 (N_30690,N_30495,N_30305);
nor U30691 (N_30691,N_30420,N_30326);
xnor U30692 (N_30692,N_30329,N_30454);
and U30693 (N_30693,N_30466,N_30369);
or U30694 (N_30694,N_30401,N_30461);
nor U30695 (N_30695,N_30423,N_30364);
nor U30696 (N_30696,N_30265,N_30498);
nand U30697 (N_30697,N_30447,N_30327);
xor U30698 (N_30698,N_30287,N_30433);
and U30699 (N_30699,N_30277,N_30291);
nand U30700 (N_30700,N_30442,N_30374);
nand U30701 (N_30701,N_30477,N_30440);
xor U30702 (N_30702,N_30448,N_30383);
xor U30703 (N_30703,N_30351,N_30419);
and U30704 (N_30704,N_30436,N_30404);
xor U30705 (N_30705,N_30300,N_30378);
nor U30706 (N_30706,N_30455,N_30321);
nor U30707 (N_30707,N_30336,N_30264);
nand U30708 (N_30708,N_30469,N_30474);
nand U30709 (N_30709,N_30273,N_30409);
and U30710 (N_30710,N_30322,N_30446);
or U30711 (N_30711,N_30359,N_30253);
or U30712 (N_30712,N_30447,N_30448);
nor U30713 (N_30713,N_30304,N_30256);
xor U30714 (N_30714,N_30263,N_30305);
xnor U30715 (N_30715,N_30254,N_30333);
or U30716 (N_30716,N_30271,N_30370);
and U30717 (N_30717,N_30363,N_30341);
nand U30718 (N_30718,N_30342,N_30383);
nor U30719 (N_30719,N_30369,N_30479);
xnor U30720 (N_30720,N_30468,N_30313);
xor U30721 (N_30721,N_30417,N_30456);
and U30722 (N_30722,N_30415,N_30328);
or U30723 (N_30723,N_30447,N_30379);
xor U30724 (N_30724,N_30387,N_30454);
nand U30725 (N_30725,N_30473,N_30370);
xnor U30726 (N_30726,N_30372,N_30433);
nand U30727 (N_30727,N_30450,N_30277);
nand U30728 (N_30728,N_30359,N_30369);
nand U30729 (N_30729,N_30487,N_30452);
xor U30730 (N_30730,N_30375,N_30293);
or U30731 (N_30731,N_30358,N_30467);
or U30732 (N_30732,N_30379,N_30347);
nand U30733 (N_30733,N_30420,N_30487);
nor U30734 (N_30734,N_30306,N_30366);
nor U30735 (N_30735,N_30408,N_30268);
nand U30736 (N_30736,N_30385,N_30348);
nor U30737 (N_30737,N_30329,N_30411);
nand U30738 (N_30738,N_30314,N_30353);
xor U30739 (N_30739,N_30402,N_30465);
and U30740 (N_30740,N_30409,N_30383);
xor U30741 (N_30741,N_30365,N_30329);
nand U30742 (N_30742,N_30250,N_30315);
xor U30743 (N_30743,N_30443,N_30369);
nand U30744 (N_30744,N_30291,N_30474);
nand U30745 (N_30745,N_30282,N_30494);
or U30746 (N_30746,N_30357,N_30358);
or U30747 (N_30747,N_30432,N_30342);
and U30748 (N_30748,N_30296,N_30292);
nand U30749 (N_30749,N_30339,N_30268);
nor U30750 (N_30750,N_30550,N_30719);
or U30751 (N_30751,N_30680,N_30722);
or U30752 (N_30752,N_30560,N_30564);
nand U30753 (N_30753,N_30549,N_30583);
nor U30754 (N_30754,N_30594,N_30712);
and U30755 (N_30755,N_30693,N_30612);
nand U30756 (N_30756,N_30642,N_30537);
nand U30757 (N_30757,N_30724,N_30524);
nand U30758 (N_30758,N_30559,N_30701);
or U30759 (N_30759,N_30606,N_30522);
or U30760 (N_30760,N_30726,N_30632);
nor U30761 (N_30761,N_30660,N_30626);
nand U30762 (N_30762,N_30734,N_30519);
and U30763 (N_30763,N_30725,N_30572);
nor U30764 (N_30764,N_30618,N_30707);
nor U30765 (N_30765,N_30562,N_30639);
or U30766 (N_30766,N_30715,N_30615);
nand U30767 (N_30767,N_30716,N_30570);
nor U30768 (N_30768,N_30717,N_30739);
or U30769 (N_30769,N_30706,N_30690);
nand U30770 (N_30770,N_30573,N_30600);
xnor U30771 (N_30771,N_30684,N_30507);
xor U30772 (N_30772,N_30575,N_30585);
nand U30773 (N_30773,N_30675,N_30566);
and U30774 (N_30774,N_30628,N_30595);
nand U30775 (N_30775,N_30687,N_30678);
nand U30776 (N_30776,N_30609,N_30649);
and U30777 (N_30777,N_30699,N_30619);
nand U30778 (N_30778,N_30588,N_30605);
nor U30779 (N_30779,N_30622,N_30544);
and U30780 (N_30780,N_30538,N_30694);
or U30781 (N_30781,N_30708,N_30532);
xnor U30782 (N_30782,N_30679,N_30598);
or U30783 (N_30783,N_30700,N_30651);
xnor U30784 (N_30784,N_30533,N_30714);
and U30785 (N_30785,N_30616,N_30603);
nor U30786 (N_30786,N_30723,N_30508);
nand U30787 (N_30787,N_30516,N_30514);
or U30788 (N_30788,N_30637,N_30521);
or U30789 (N_30789,N_30674,N_30696);
or U30790 (N_30790,N_30703,N_30540);
nor U30791 (N_30791,N_30506,N_30740);
nand U30792 (N_30792,N_30737,N_30556);
or U30793 (N_30793,N_30689,N_30691);
nor U30794 (N_30794,N_30535,N_30744);
or U30795 (N_30795,N_30665,N_30747);
and U30796 (N_30796,N_30713,N_30662);
and U30797 (N_30797,N_30623,N_30681);
nand U30798 (N_30798,N_30643,N_30543);
xnor U30799 (N_30799,N_30647,N_30523);
nand U30800 (N_30800,N_30501,N_30511);
or U30801 (N_30801,N_30614,N_30646);
nor U30802 (N_30802,N_30705,N_30648);
nand U30803 (N_30803,N_30733,N_30650);
or U30804 (N_30804,N_30657,N_30663);
or U30805 (N_30805,N_30576,N_30546);
or U30806 (N_30806,N_30685,N_30654);
and U30807 (N_30807,N_30698,N_30539);
or U30808 (N_30808,N_30688,N_30574);
xnor U30809 (N_30809,N_30569,N_30620);
or U30810 (N_30810,N_30579,N_30526);
and U30811 (N_30811,N_30509,N_30629);
or U30812 (N_30812,N_30520,N_30607);
or U30813 (N_30813,N_30593,N_30563);
or U30814 (N_30814,N_30502,N_30658);
xor U30815 (N_30815,N_30621,N_30721);
and U30816 (N_30816,N_30636,N_30590);
xor U30817 (N_30817,N_30731,N_30518);
xor U30818 (N_30818,N_30624,N_30672);
nand U30819 (N_30819,N_30503,N_30517);
nand U30820 (N_30820,N_30697,N_30673);
nor U30821 (N_30821,N_30627,N_30541);
nand U30822 (N_30822,N_30584,N_30676);
xnor U30823 (N_30823,N_30631,N_30611);
and U30824 (N_30824,N_30510,N_30586);
and U30825 (N_30825,N_30551,N_30710);
xor U30826 (N_30826,N_30525,N_30727);
or U30827 (N_30827,N_30513,N_30592);
or U30828 (N_30828,N_30635,N_30587);
and U30829 (N_30829,N_30531,N_30746);
and U30830 (N_30830,N_30512,N_30601);
xor U30831 (N_30831,N_30547,N_30630);
nand U30832 (N_30832,N_30655,N_30548);
and U30833 (N_30833,N_30641,N_30553);
and U30834 (N_30834,N_30561,N_30656);
and U30835 (N_30835,N_30709,N_30666);
nand U30836 (N_30836,N_30671,N_30597);
nor U30837 (N_30837,N_30500,N_30683);
or U30838 (N_30838,N_30555,N_30711);
nor U30839 (N_30839,N_30677,N_30728);
xor U30840 (N_30840,N_30589,N_30736);
or U30841 (N_30841,N_30745,N_30599);
or U30842 (N_30842,N_30530,N_30552);
and U30843 (N_30843,N_30704,N_30610);
xor U30844 (N_30844,N_30670,N_30743);
nand U30845 (N_30845,N_30617,N_30652);
nor U30846 (N_30846,N_30528,N_30742);
and U30847 (N_30847,N_30633,N_30702);
and U30848 (N_30848,N_30504,N_30568);
xor U30849 (N_30849,N_30730,N_30529);
nor U30850 (N_30850,N_30667,N_30735);
xnor U30851 (N_30851,N_30640,N_30515);
xnor U30852 (N_30852,N_30738,N_30580);
xnor U30853 (N_30853,N_30613,N_30659);
and U30854 (N_30854,N_30686,N_30581);
or U30855 (N_30855,N_30554,N_30602);
xor U30856 (N_30856,N_30720,N_30565);
nor U30857 (N_30857,N_30578,N_30558);
or U30858 (N_30858,N_30692,N_30577);
xor U30859 (N_30859,N_30591,N_30741);
or U30860 (N_30860,N_30527,N_30534);
nor U30861 (N_30861,N_30664,N_30604);
or U30862 (N_30862,N_30729,N_30718);
or U30863 (N_30863,N_30625,N_30661);
nor U30864 (N_30864,N_30582,N_30695);
xor U30865 (N_30865,N_30668,N_30571);
or U30866 (N_30866,N_30638,N_30567);
or U30867 (N_30867,N_30542,N_30682);
nor U30868 (N_30868,N_30545,N_30669);
xnor U30869 (N_30869,N_30596,N_30732);
nand U30870 (N_30870,N_30749,N_30505);
nor U30871 (N_30871,N_30634,N_30557);
xor U30872 (N_30872,N_30645,N_30608);
nand U30873 (N_30873,N_30748,N_30536);
nor U30874 (N_30874,N_30644,N_30653);
or U30875 (N_30875,N_30551,N_30717);
or U30876 (N_30876,N_30633,N_30672);
xor U30877 (N_30877,N_30606,N_30661);
and U30878 (N_30878,N_30615,N_30583);
xnor U30879 (N_30879,N_30711,N_30577);
and U30880 (N_30880,N_30714,N_30736);
or U30881 (N_30881,N_30571,N_30720);
or U30882 (N_30882,N_30641,N_30554);
nor U30883 (N_30883,N_30632,N_30631);
or U30884 (N_30884,N_30576,N_30713);
nor U30885 (N_30885,N_30637,N_30614);
nor U30886 (N_30886,N_30730,N_30656);
and U30887 (N_30887,N_30611,N_30732);
or U30888 (N_30888,N_30682,N_30538);
xnor U30889 (N_30889,N_30531,N_30538);
nor U30890 (N_30890,N_30675,N_30691);
nand U30891 (N_30891,N_30653,N_30663);
nor U30892 (N_30892,N_30628,N_30679);
or U30893 (N_30893,N_30682,N_30504);
and U30894 (N_30894,N_30704,N_30620);
nand U30895 (N_30895,N_30634,N_30516);
nand U30896 (N_30896,N_30739,N_30615);
or U30897 (N_30897,N_30676,N_30720);
and U30898 (N_30898,N_30616,N_30575);
or U30899 (N_30899,N_30578,N_30592);
nor U30900 (N_30900,N_30548,N_30608);
and U30901 (N_30901,N_30657,N_30603);
xnor U30902 (N_30902,N_30504,N_30614);
nand U30903 (N_30903,N_30608,N_30690);
xnor U30904 (N_30904,N_30576,N_30737);
xor U30905 (N_30905,N_30635,N_30507);
and U30906 (N_30906,N_30682,N_30743);
or U30907 (N_30907,N_30547,N_30707);
nor U30908 (N_30908,N_30698,N_30704);
nand U30909 (N_30909,N_30611,N_30557);
nor U30910 (N_30910,N_30546,N_30618);
nor U30911 (N_30911,N_30505,N_30626);
xor U30912 (N_30912,N_30584,N_30517);
nand U30913 (N_30913,N_30572,N_30708);
nor U30914 (N_30914,N_30541,N_30598);
and U30915 (N_30915,N_30748,N_30540);
nand U30916 (N_30916,N_30541,N_30533);
or U30917 (N_30917,N_30583,N_30712);
and U30918 (N_30918,N_30607,N_30699);
and U30919 (N_30919,N_30623,N_30642);
and U30920 (N_30920,N_30631,N_30714);
or U30921 (N_30921,N_30594,N_30657);
or U30922 (N_30922,N_30705,N_30584);
or U30923 (N_30923,N_30665,N_30586);
and U30924 (N_30924,N_30663,N_30595);
nor U30925 (N_30925,N_30604,N_30549);
nand U30926 (N_30926,N_30598,N_30580);
xnor U30927 (N_30927,N_30588,N_30502);
and U30928 (N_30928,N_30737,N_30638);
and U30929 (N_30929,N_30563,N_30727);
or U30930 (N_30930,N_30728,N_30504);
or U30931 (N_30931,N_30601,N_30504);
or U30932 (N_30932,N_30684,N_30565);
nor U30933 (N_30933,N_30601,N_30656);
xor U30934 (N_30934,N_30532,N_30527);
and U30935 (N_30935,N_30563,N_30674);
and U30936 (N_30936,N_30744,N_30585);
and U30937 (N_30937,N_30689,N_30738);
nand U30938 (N_30938,N_30642,N_30538);
xnor U30939 (N_30939,N_30671,N_30699);
nand U30940 (N_30940,N_30621,N_30697);
xor U30941 (N_30941,N_30554,N_30529);
or U30942 (N_30942,N_30689,N_30706);
xor U30943 (N_30943,N_30743,N_30531);
nand U30944 (N_30944,N_30530,N_30540);
and U30945 (N_30945,N_30547,N_30518);
and U30946 (N_30946,N_30607,N_30582);
nand U30947 (N_30947,N_30609,N_30542);
or U30948 (N_30948,N_30709,N_30600);
xnor U30949 (N_30949,N_30717,N_30574);
nand U30950 (N_30950,N_30574,N_30539);
nor U30951 (N_30951,N_30623,N_30545);
or U30952 (N_30952,N_30537,N_30523);
nor U30953 (N_30953,N_30636,N_30721);
xor U30954 (N_30954,N_30516,N_30561);
nor U30955 (N_30955,N_30685,N_30528);
and U30956 (N_30956,N_30638,N_30727);
nand U30957 (N_30957,N_30511,N_30672);
nand U30958 (N_30958,N_30511,N_30545);
or U30959 (N_30959,N_30586,N_30639);
xor U30960 (N_30960,N_30606,N_30623);
or U30961 (N_30961,N_30688,N_30659);
nand U30962 (N_30962,N_30623,N_30512);
or U30963 (N_30963,N_30578,N_30709);
xnor U30964 (N_30964,N_30570,N_30663);
xor U30965 (N_30965,N_30634,N_30616);
xnor U30966 (N_30966,N_30734,N_30644);
nor U30967 (N_30967,N_30510,N_30573);
and U30968 (N_30968,N_30579,N_30730);
nand U30969 (N_30969,N_30672,N_30708);
nand U30970 (N_30970,N_30614,N_30527);
or U30971 (N_30971,N_30544,N_30735);
and U30972 (N_30972,N_30517,N_30654);
xnor U30973 (N_30973,N_30529,N_30557);
nor U30974 (N_30974,N_30695,N_30694);
xnor U30975 (N_30975,N_30559,N_30578);
or U30976 (N_30976,N_30685,N_30709);
and U30977 (N_30977,N_30614,N_30532);
or U30978 (N_30978,N_30551,N_30699);
nand U30979 (N_30979,N_30727,N_30632);
xnor U30980 (N_30980,N_30735,N_30647);
nand U30981 (N_30981,N_30606,N_30711);
nor U30982 (N_30982,N_30606,N_30529);
nor U30983 (N_30983,N_30673,N_30696);
nand U30984 (N_30984,N_30547,N_30597);
or U30985 (N_30985,N_30672,N_30524);
or U30986 (N_30986,N_30650,N_30609);
nand U30987 (N_30987,N_30595,N_30518);
and U30988 (N_30988,N_30699,N_30532);
xor U30989 (N_30989,N_30701,N_30705);
and U30990 (N_30990,N_30649,N_30714);
xor U30991 (N_30991,N_30613,N_30503);
xor U30992 (N_30992,N_30672,N_30599);
xor U30993 (N_30993,N_30651,N_30684);
xor U30994 (N_30994,N_30594,N_30604);
xor U30995 (N_30995,N_30651,N_30742);
nor U30996 (N_30996,N_30648,N_30565);
nand U30997 (N_30997,N_30592,N_30530);
or U30998 (N_30998,N_30715,N_30662);
nand U30999 (N_30999,N_30722,N_30655);
nand U31000 (N_31000,N_30952,N_30759);
and U31001 (N_31001,N_30940,N_30892);
xor U31002 (N_31002,N_30863,N_30920);
nand U31003 (N_31003,N_30933,N_30874);
nand U31004 (N_31004,N_30967,N_30969);
xor U31005 (N_31005,N_30907,N_30924);
or U31006 (N_31006,N_30807,N_30965);
nand U31007 (N_31007,N_30806,N_30912);
and U31008 (N_31008,N_30964,N_30829);
and U31009 (N_31009,N_30886,N_30899);
nand U31010 (N_31010,N_30769,N_30849);
nor U31011 (N_31011,N_30750,N_30783);
nor U31012 (N_31012,N_30900,N_30843);
nand U31013 (N_31013,N_30795,N_30754);
and U31014 (N_31014,N_30794,N_30976);
nor U31015 (N_31015,N_30793,N_30963);
xnor U31016 (N_31016,N_30842,N_30764);
or U31017 (N_31017,N_30796,N_30858);
and U31018 (N_31018,N_30848,N_30936);
or U31019 (N_31019,N_30988,N_30875);
or U31020 (N_31020,N_30786,N_30770);
or U31021 (N_31021,N_30774,N_30763);
and U31022 (N_31022,N_30890,N_30881);
and U31023 (N_31023,N_30766,N_30974);
or U31024 (N_31024,N_30878,N_30817);
and U31025 (N_31025,N_30841,N_30951);
or U31026 (N_31026,N_30827,N_30761);
nor U31027 (N_31027,N_30929,N_30943);
nor U31028 (N_31028,N_30953,N_30950);
or U31029 (N_31029,N_30777,N_30859);
nor U31030 (N_31030,N_30934,N_30828);
nor U31031 (N_31031,N_30882,N_30866);
and U31032 (N_31032,N_30853,N_30855);
and U31033 (N_31033,N_30909,N_30871);
and U31034 (N_31034,N_30998,N_30864);
or U31035 (N_31035,N_30787,N_30992);
nand U31036 (N_31036,N_30895,N_30986);
xor U31037 (N_31037,N_30814,N_30928);
and U31038 (N_31038,N_30993,N_30815);
or U31039 (N_31039,N_30824,N_30847);
nor U31040 (N_31040,N_30941,N_30994);
nand U31041 (N_31041,N_30823,N_30876);
and U31042 (N_31042,N_30756,N_30903);
nor U31043 (N_31043,N_30962,N_30808);
nand U31044 (N_31044,N_30954,N_30984);
nand U31045 (N_31045,N_30898,N_30942);
xor U31046 (N_31046,N_30927,N_30785);
nand U31047 (N_31047,N_30801,N_30836);
nor U31048 (N_31048,N_30802,N_30985);
xor U31049 (N_31049,N_30872,N_30753);
nor U31050 (N_31050,N_30885,N_30956);
or U31051 (N_31051,N_30916,N_30851);
and U31052 (N_31052,N_30865,N_30758);
nand U31053 (N_31053,N_30910,N_30803);
xor U31054 (N_31054,N_30883,N_30911);
nand U31055 (N_31055,N_30922,N_30778);
nor U31056 (N_31056,N_30884,N_30804);
xnor U31057 (N_31057,N_30811,N_30930);
nor U31058 (N_31058,N_30935,N_30854);
and U31059 (N_31059,N_30757,N_30879);
or U31060 (N_31060,N_30995,N_30955);
nor U31061 (N_31061,N_30977,N_30790);
nand U31062 (N_31062,N_30780,N_30887);
xnor U31063 (N_31063,N_30914,N_30945);
and U31064 (N_31064,N_30908,N_30972);
nand U31065 (N_31065,N_30792,N_30773);
or U31066 (N_31066,N_30921,N_30996);
and U31067 (N_31067,N_30968,N_30846);
or U31068 (N_31068,N_30873,N_30791);
and U31069 (N_31069,N_30970,N_30822);
xor U31070 (N_31070,N_30821,N_30771);
xor U31071 (N_31071,N_30939,N_30832);
nand U31072 (N_31072,N_30946,N_30852);
nand U31073 (N_31073,N_30931,N_30856);
nor U31074 (N_31074,N_30833,N_30980);
xor U31075 (N_31075,N_30888,N_30925);
nor U31076 (N_31076,N_30889,N_30966);
nor U31077 (N_31077,N_30752,N_30989);
and U31078 (N_31078,N_30957,N_30971);
and U31079 (N_31079,N_30997,N_30897);
nor U31080 (N_31080,N_30901,N_30902);
or U31081 (N_31081,N_30818,N_30978);
or U31082 (N_31082,N_30835,N_30990);
nor U31083 (N_31083,N_30798,N_30973);
or U31084 (N_31084,N_30772,N_30809);
and U31085 (N_31085,N_30775,N_30938);
nand U31086 (N_31086,N_30776,N_30805);
or U31087 (N_31087,N_30813,N_30755);
and U31088 (N_31088,N_30760,N_30987);
and U31089 (N_31089,N_30944,N_30932);
or U31090 (N_31090,N_30860,N_30812);
nor U31091 (N_31091,N_30923,N_30831);
nor U31092 (N_31092,N_30782,N_30918);
nor U31093 (N_31093,N_30869,N_30784);
nor U31094 (N_31094,N_30819,N_30820);
nor U31095 (N_31095,N_30816,N_30797);
nor U31096 (N_31096,N_30904,N_30975);
xor U31097 (N_31097,N_30868,N_30982);
xnor U31098 (N_31098,N_30983,N_30762);
nand U31099 (N_31099,N_30960,N_30915);
xor U31100 (N_31100,N_30959,N_30880);
and U31101 (N_31101,N_30837,N_30961);
nor U31102 (N_31102,N_30896,N_30857);
or U31103 (N_31103,N_30862,N_30991);
xor U31104 (N_31104,N_30799,N_30926);
nand U31105 (N_31105,N_30893,N_30981);
and U31106 (N_31106,N_30948,N_30894);
xnor U31107 (N_31107,N_30979,N_30891);
nor U31108 (N_31108,N_30937,N_30830);
and U31109 (N_31109,N_30826,N_30839);
nor U31110 (N_31110,N_30949,N_30781);
and U31111 (N_31111,N_30768,N_30906);
nor U31112 (N_31112,N_30861,N_30767);
or U31113 (N_31113,N_30825,N_30840);
or U31114 (N_31114,N_30870,N_30845);
and U31115 (N_31115,N_30913,N_30765);
xnor U31116 (N_31116,N_30958,N_30788);
or U31117 (N_31117,N_30844,N_30867);
xnor U31118 (N_31118,N_30810,N_30947);
nand U31119 (N_31119,N_30751,N_30877);
and U31120 (N_31120,N_30919,N_30850);
xor U31121 (N_31121,N_30779,N_30999);
xnor U31122 (N_31122,N_30917,N_30838);
and U31123 (N_31123,N_30905,N_30789);
and U31124 (N_31124,N_30800,N_30834);
and U31125 (N_31125,N_30900,N_30884);
and U31126 (N_31126,N_30837,N_30827);
nand U31127 (N_31127,N_30883,N_30872);
and U31128 (N_31128,N_30756,N_30967);
nand U31129 (N_31129,N_30976,N_30773);
and U31130 (N_31130,N_30926,N_30911);
nor U31131 (N_31131,N_30769,N_30917);
and U31132 (N_31132,N_30887,N_30809);
nor U31133 (N_31133,N_30911,N_30867);
nand U31134 (N_31134,N_30939,N_30961);
and U31135 (N_31135,N_30969,N_30839);
nand U31136 (N_31136,N_30756,N_30767);
xnor U31137 (N_31137,N_30990,N_30850);
xor U31138 (N_31138,N_30878,N_30920);
and U31139 (N_31139,N_30866,N_30823);
nand U31140 (N_31140,N_30967,N_30948);
nor U31141 (N_31141,N_30761,N_30863);
xnor U31142 (N_31142,N_30773,N_30973);
nand U31143 (N_31143,N_30865,N_30953);
nor U31144 (N_31144,N_30875,N_30945);
nand U31145 (N_31145,N_30755,N_30753);
nand U31146 (N_31146,N_30884,N_30783);
nand U31147 (N_31147,N_30789,N_30764);
nand U31148 (N_31148,N_30873,N_30991);
or U31149 (N_31149,N_30988,N_30786);
nand U31150 (N_31150,N_30959,N_30791);
nand U31151 (N_31151,N_30783,N_30828);
nor U31152 (N_31152,N_30816,N_30940);
xnor U31153 (N_31153,N_30973,N_30971);
and U31154 (N_31154,N_30793,N_30825);
and U31155 (N_31155,N_30920,N_30890);
xnor U31156 (N_31156,N_30855,N_30948);
xor U31157 (N_31157,N_30818,N_30867);
nor U31158 (N_31158,N_30778,N_30808);
xor U31159 (N_31159,N_30852,N_30970);
or U31160 (N_31160,N_30900,N_30759);
or U31161 (N_31161,N_30783,N_30910);
nor U31162 (N_31162,N_30770,N_30818);
or U31163 (N_31163,N_30947,N_30990);
xnor U31164 (N_31164,N_30942,N_30842);
and U31165 (N_31165,N_30935,N_30813);
nand U31166 (N_31166,N_30896,N_30838);
xor U31167 (N_31167,N_30956,N_30905);
and U31168 (N_31168,N_30863,N_30813);
nand U31169 (N_31169,N_30796,N_30812);
xor U31170 (N_31170,N_30931,N_30754);
nand U31171 (N_31171,N_30829,N_30900);
or U31172 (N_31172,N_30786,N_30849);
or U31173 (N_31173,N_30907,N_30912);
xor U31174 (N_31174,N_30896,N_30873);
and U31175 (N_31175,N_30803,N_30940);
and U31176 (N_31176,N_30939,N_30920);
nand U31177 (N_31177,N_30960,N_30896);
xor U31178 (N_31178,N_30850,N_30979);
nand U31179 (N_31179,N_30861,N_30839);
nand U31180 (N_31180,N_30956,N_30841);
or U31181 (N_31181,N_30906,N_30888);
xnor U31182 (N_31182,N_30887,N_30825);
nand U31183 (N_31183,N_30939,N_30855);
and U31184 (N_31184,N_30838,N_30822);
nor U31185 (N_31185,N_30828,N_30793);
or U31186 (N_31186,N_30941,N_30802);
nor U31187 (N_31187,N_30862,N_30893);
nor U31188 (N_31188,N_30955,N_30978);
nand U31189 (N_31189,N_30813,N_30956);
and U31190 (N_31190,N_30825,N_30761);
nor U31191 (N_31191,N_30954,N_30870);
xor U31192 (N_31192,N_30948,N_30752);
or U31193 (N_31193,N_30903,N_30908);
or U31194 (N_31194,N_30843,N_30756);
nor U31195 (N_31195,N_30860,N_30848);
and U31196 (N_31196,N_30980,N_30892);
or U31197 (N_31197,N_30879,N_30851);
nand U31198 (N_31198,N_30931,N_30750);
and U31199 (N_31199,N_30759,N_30854);
or U31200 (N_31200,N_30982,N_30851);
xnor U31201 (N_31201,N_30859,N_30802);
nand U31202 (N_31202,N_30957,N_30849);
and U31203 (N_31203,N_30841,N_30974);
nand U31204 (N_31204,N_30970,N_30922);
nor U31205 (N_31205,N_30772,N_30994);
xnor U31206 (N_31206,N_30875,N_30809);
or U31207 (N_31207,N_30785,N_30753);
nor U31208 (N_31208,N_30809,N_30914);
nand U31209 (N_31209,N_30886,N_30879);
xor U31210 (N_31210,N_30847,N_30878);
nor U31211 (N_31211,N_30793,N_30863);
nor U31212 (N_31212,N_30776,N_30775);
nand U31213 (N_31213,N_30930,N_30976);
nand U31214 (N_31214,N_30951,N_30843);
nand U31215 (N_31215,N_30839,N_30894);
xnor U31216 (N_31216,N_30947,N_30949);
nor U31217 (N_31217,N_30959,N_30799);
nand U31218 (N_31218,N_30982,N_30881);
xor U31219 (N_31219,N_30952,N_30819);
or U31220 (N_31220,N_30987,N_30763);
xnor U31221 (N_31221,N_30825,N_30964);
or U31222 (N_31222,N_30886,N_30763);
nand U31223 (N_31223,N_30992,N_30962);
xnor U31224 (N_31224,N_30971,N_30759);
nor U31225 (N_31225,N_30810,N_30890);
or U31226 (N_31226,N_30835,N_30822);
nand U31227 (N_31227,N_30881,N_30986);
nor U31228 (N_31228,N_30900,N_30919);
nor U31229 (N_31229,N_30928,N_30960);
and U31230 (N_31230,N_30874,N_30949);
and U31231 (N_31231,N_30824,N_30849);
nor U31232 (N_31232,N_30774,N_30917);
or U31233 (N_31233,N_30833,N_30845);
and U31234 (N_31234,N_30942,N_30765);
nor U31235 (N_31235,N_30939,N_30934);
nand U31236 (N_31236,N_30796,N_30932);
xnor U31237 (N_31237,N_30912,N_30909);
nor U31238 (N_31238,N_30970,N_30886);
nand U31239 (N_31239,N_30797,N_30988);
nand U31240 (N_31240,N_30842,N_30848);
xnor U31241 (N_31241,N_30868,N_30897);
nor U31242 (N_31242,N_30774,N_30998);
and U31243 (N_31243,N_30760,N_30863);
or U31244 (N_31244,N_30980,N_30994);
and U31245 (N_31245,N_30969,N_30788);
or U31246 (N_31246,N_30937,N_30834);
and U31247 (N_31247,N_30805,N_30971);
and U31248 (N_31248,N_30911,N_30854);
xor U31249 (N_31249,N_30918,N_30923);
or U31250 (N_31250,N_31157,N_31048);
and U31251 (N_31251,N_31150,N_31137);
and U31252 (N_31252,N_31143,N_31201);
and U31253 (N_31253,N_31067,N_31158);
or U31254 (N_31254,N_31189,N_31068);
or U31255 (N_31255,N_31064,N_31040);
or U31256 (N_31256,N_31090,N_31019);
xnor U31257 (N_31257,N_31088,N_31066);
and U31258 (N_31258,N_31000,N_31050);
nor U31259 (N_31259,N_31245,N_31011);
nand U31260 (N_31260,N_31186,N_31237);
or U31261 (N_31261,N_31145,N_31176);
xor U31262 (N_31262,N_31012,N_31168);
nand U31263 (N_31263,N_31170,N_31192);
or U31264 (N_31264,N_31004,N_31230);
xnor U31265 (N_31265,N_31219,N_31041);
nor U31266 (N_31266,N_31093,N_31075);
nand U31267 (N_31267,N_31156,N_31139);
nor U31268 (N_31268,N_31122,N_31119);
or U31269 (N_31269,N_31118,N_31001);
or U31270 (N_31270,N_31023,N_31130);
or U31271 (N_31271,N_31181,N_31208);
nand U31272 (N_31272,N_31211,N_31206);
nor U31273 (N_31273,N_31077,N_31248);
xnor U31274 (N_31274,N_31106,N_31178);
and U31275 (N_31275,N_31129,N_31190);
nor U31276 (N_31276,N_31007,N_31217);
xnor U31277 (N_31277,N_31022,N_31229);
or U31278 (N_31278,N_31015,N_31243);
nor U31279 (N_31279,N_31202,N_31117);
nor U31280 (N_31280,N_31128,N_31037);
or U31281 (N_31281,N_31153,N_31020);
nor U31282 (N_31282,N_31021,N_31172);
and U31283 (N_31283,N_31095,N_31113);
xor U31284 (N_31284,N_31197,N_31084);
nor U31285 (N_31285,N_31140,N_31127);
or U31286 (N_31286,N_31204,N_31134);
and U31287 (N_31287,N_31205,N_31044);
nor U31288 (N_31288,N_31138,N_31058);
xnor U31289 (N_31289,N_31108,N_31086);
and U31290 (N_31290,N_31141,N_31161);
nand U31291 (N_31291,N_31238,N_31220);
and U31292 (N_31292,N_31036,N_31212);
nand U31293 (N_31293,N_31039,N_31236);
and U31294 (N_31294,N_31191,N_31029);
or U31295 (N_31295,N_31144,N_31227);
or U31296 (N_31296,N_31087,N_31125);
and U31297 (N_31297,N_31203,N_31196);
xnor U31298 (N_31298,N_31160,N_31060);
xor U31299 (N_31299,N_31146,N_31225);
and U31300 (N_31300,N_31026,N_31148);
or U31301 (N_31301,N_31092,N_31193);
nor U31302 (N_31302,N_31226,N_31155);
and U31303 (N_31303,N_31006,N_31057);
or U31304 (N_31304,N_31249,N_31016);
or U31305 (N_31305,N_31235,N_31246);
nor U31306 (N_31306,N_31222,N_31078);
and U31307 (N_31307,N_31213,N_31123);
nor U31308 (N_31308,N_31173,N_31059);
and U31309 (N_31309,N_31080,N_31214);
and U31310 (N_31310,N_31244,N_31098);
and U31311 (N_31311,N_31200,N_31224);
or U31312 (N_31312,N_31194,N_31136);
and U31313 (N_31313,N_31198,N_31107);
nor U31314 (N_31314,N_31232,N_31180);
and U31315 (N_31315,N_31076,N_31010);
nand U31316 (N_31316,N_31069,N_31115);
nand U31317 (N_31317,N_31074,N_31133);
nor U31318 (N_31318,N_31241,N_31215);
nand U31319 (N_31319,N_31152,N_31008);
nand U31320 (N_31320,N_31096,N_31182);
nor U31321 (N_31321,N_31223,N_31177);
xor U31322 (N_31322,N_31174,N_31154);
or U31323 (N_31323,N_31147,N_31165);
nor U31324 (N_31324,N_31065,N_31171);
nand U31325 (N_31325,N_31184,N_31073);
or U31326 (N_31326,N_31116,N_31185);
nand U31327 (N_31327,N_31110,N_31179);
xnor U31328 (N_31328,N_31013,N_31135);
nor U31329 (N_31329,N_31027,N_31091);
nor U31330 (N_31330,N_31089,N_31045);
nor U31331 (N_31331,N_31131,N_31028);
or U31332 (N_31332,N_31104,N_31183);
nor U31333 (N_31333,N_31017,N_31210);
nor U31334 (N_31334,N_31142,N_31187);
and U31335 (N_31335,N_31018,N_31149);
nand U31336 (N_31336,N_31112,N_31126);
nor U31337 (N_31337,N_31053,N_31030);
xor U31338 (N_31338,N_31056,N_31162);
or U31339 (N_31339,N_31070,N_31046);
nand U31340 (N_31340,N_31097,N_31024);
nor U31341 (N_31341,N_31071,N_31207);
or U31342 (N_31342,N_31221,N_31043);
nand U31343 (N_31343,N_31175,N_31188);
xnor U31344 (N_31344,N_31240,N_31099);
nor U31345 (N_31345,N_31083,N_31049);
or U31346 (N_31346,N_31005,N_31072);
or U31347 (N_31347,N_31047,N_31062);
and U31348 (N_31348,N_31082,N_31033);
nor U31349 (N_31349,N_31063,N_31014);
xnor U31350 (N_31350,N_31151,N_31216);
nor U31351 (N_31351,N_31035,N_31034);
nor U31352 (N_31352,N_31163,N_31103);
and U31353 (N_31353,N_31061,N_31231);
xor U31354 (N_31354,N_31124,N_31009);
and U31355 (N_31355,N_31242,N_31218);
xor U31356 (N_31356,N_31101,N_31052);
nand U31357 (N_31357,N_31054,N_31164);
and U31358 (N_31358,N_31239,N_31051);
nand U31359 (N_31359,N_31209,N_31169);
nand U31360 (N_31360,N_31081,N_31132);
nor U31361 (N_31361,N_31032,N_31111);
nand U31362 (N_31362,N_31195,N_31121);
or U31363 (N_31363,N_31003,N_31100);
or U31364 (N_31364,N_31055,N_31042);
and U31365 (N_31365,N_31247,N_31105);
and U31366 (N_31366,N_31233,N_31120);
and U31367 (N_31367,N_31114,N_31038);
nand U31368 (N_31368,N_31002,N_31031);
xor U31369 (N_31369,N_31085,N_31079);
nand U31370 (N_31370,N_31166,N_31094);
and U31371 (N_31371,N_31109,N_31025);
nor U31372 (N_31372,N_31159,N_31167);
nor U31373 (N_31373,N_31234,N_31102);
nor U31374 (N_31374,N_31199,N_31228);
nor U31375 (N_31375,N_31032,N_31075);
xor U31376 (N_31376,N_31136,N_31051);
xnor U31377 (N_31377,N_31225,N_31155);
xor U31378 (N_31378,N_31137,N_31072);
nor U31379 (N_31379,N_31016,N_31065);
and U31380 (N_31380,N_31020,N_31001);
nand U31381 (N_31381,N_31240,N_31074);
nand U31382 (N_31382,N_31236,N_31159);
nand U31383 (N_31383,N_31028,N_31080);
xnor U31384 (N_31384,N_31174,N_31061);
nor U31385 (N_31385,N_31219,N_31050);
and U31386 (N_31386,N_31057,N_31047);
nand U31387 (N_31387,N_31127,N_31121);
or U31388 (N_31388,N_31034,N_31151);
and U31389 (N_31389,N_31144,N_31134);
nand U31390 (N_31390,N_31199,N_31108);
nand U31391 (N_31391,N_31105,N_31132);
xnor U31392 (N_31392,N_31057,N_31078);
nand U31393 (N_31393,N_31246,N_31107);
xor U31394 (N_31394,N_31185,N_31178);
nand U31395 (N_31395,N_31161,N_31035);
and U31396 (N_31396,N_31076,N_31007);
and U31397 (N_31397,N_31233,N_31069);
xnor U31398 (N_31398,N_31228,N_31129);
and U31399 (N_31399,N_31039,N_31001);
nor U31400 (N_31400,N_31009,N_31034);
xor U31401 (N_31401,N_31105,N_31053);
or U31402 (N_31402,N_31031,N_31074);
nand U31403 (N_31403,N_31027,N_31208);
nor U31404 (N_31404,N_31149,N_31178);
and U31405 (N_31405,N_31242,N_31019);
and U31406 (N_31406,N_31020,N_31056);
or U31407 (N_31407,N_31082,N_31136);
or U31408 (N_31408,N_31150,N_31201);
or U31409 (N_31409,N_31110,N_31187);
and U31410 (N_31410,N_31084,N_31070);
nor U31411 (N_31411,N_31055,N_31012);
xor U31412 (N_31412,N_31129,N_31021);
nor U31413 (N_31413,N_31129,N_31145);
nor U31414 (N_31414,N_31001,N_31218);
nand U31415 (N_31415,N_31159,N_31240);
and U31416 (N_31416,N_31143,N_31194);
xor U31417 (N_31417,N_31129,N_31139);
and U31418 (N_31418,N_31010,N_31242);
or U31419 (N_31419,N_31121,N_31060);
xnor U31420 (N_31420,N_31148,N_31133);
and U31421 (N_31421,N_31178,N_31013);
or U31422 (N_31422,N_31109,N_31223);
or U31423 (N_31423,N_31066,N_31187);
nand U31424 (N_31424,N_31151,N_31168);
xnor U31425 (N_31425,N_31121,N_31125);
and U31426 (N_31426,N_31147,N_31193);
and U31427 (N_31427,N_31077,N_31057);
nor U31428 (N_31428,N_31229,N_31223);
xnor U31429 (N_31429,N_31114,N_31087);
nor U31430 (N_31430,N_31076,N_31105);
and U31431 (N_31431,N_31197,N_31085);
or U31432 (N_31432,N_31195,N_31215);
xnor U31433 (N_31433,N_31236,N_31248);
xnor U31434 (N_31434,N_31186,N_31004);
or U31435 (N_31435,N_31082,N_31072);
and U31436 (N_31436,N_31133,N_31031);
or U31437 (N_31437,N_31074,N_31175);
and U31438 (N_31438,N_31064,N_31112);
xnor U31439 (N_31439,N_31012,N_31021);
xor U31440 (N_31440,N_31016,N_31041);
and U31441 (N_31441,N_31225,N_31189);
nor U31442 (N_31442,N_31142,N_31005);
nor U31443 (N_31443,N_31117,N_31227);
or U31444 (N_31444,N_31071,N_31237);
nand U31445 (N_31445,N_31249,N_31167);
xnor U31446 (N_31446,N_31009,N_31102);
nor U31447 (N_31447,N_31185,N_31134);
nand U31448 (N_31448,N_31179,N_31062);
xnor U31449 (N_31449,N_31148,N_31100);
xnor U31450 (N_31450,N_31233,N_31026);
nand U31451 (N_31451,N_31089,N_31225);
or U31452 (N_31452,N_31247,N_31062);
or U31453 (N_31453,N_31202,N_31112);
xor U31454 (N_31454,N_31046,N_31133);
and U31455 (N_31455,N_31050,N_31063);
nor U31456 (N_31456,N_31141,N_31017);
nor U31457 (N_31457,N_31123,N_31187);
or U31458 (N_31458,N_31189,N_31167);
or U31459 (N_31459,N_31200,N_31238);
nand U31460 (N_31460,N_31093,N_31033);
xnor U31461 (N_31461,N_31182,N_31015);
nand U31462 (N_31462,N_31187,N_31058);
or U31463 (N_31463,N_31009,N_31048);
and U31464 (N_31464,N_31114,N_31033);
and U31465 (N_31465,N_31202,N_31010);
or U31466 (N_31466,N_31101,N_31177);
xnor U31467 (N_31467,N_31141,N_31202);
and U31468 (N_31468,N_31146,N_31088);
and U31469 (N_31469,N_31042,N_31041);
nand U31470 (N_31470,N_31068,N_31007);
nor U31471 (N_31471,N_31224,N_31004);
xnor U31472 (N_31472,N_31246,N_31209);
or U31473 (N_31473,N_31152,N_31053);
or U31474 (N_31474,N_31130,N_31022);
nand U31475 (N_31475,N_31142,N_31220);
nand U31476 (N_31476,N_31162,N_31002);
nor U31477 (N_31477,N_31203,N_31084);
nand U31478 (N_31478,N_31087,N_31230);
and U31479 (N_31479,N_31016,N_31006);
and U31480 (N_31480,N_31189,N_31076);
nand U31481 (N_31481,N_31111,N_31098);
nor U31482 (N_31482,N_31049,N_31137);
and U31483 (N_31483,N_31004,N_31009);
nand U31484 (N_31484,N_31207,N_31067);
nand U31485 (N_31485,N_31048,N_31153);
nand U31486 (N_31486,N_31129,N_31134);
or U31487 (N_31487,N_31087,N_31206);
xnor U31488 (N_31488,N_31148,N_31169);
or U31489 (N_31489,N_31207,N_31037);
and U31490 (N_31490,N_31186,N_31239);
and U31491 (N_31491,N_31244,N_31201);
nor U31492 (N_31492,N_31154,N_31055);
and U31493 (N_31493,N_31245,N_31189);
or U31494 (N_31494,N_31217,N_31131);
nand U31495 (N_31495,N_31229,N_31072);
and U31496 (N_31496,N_31186,N_31227);
xor U31497 (N_31497,N_31168,N_31065);
and U31498 (N_31498,N_31228,N_31226);
xnor U31499 (N_31499,N_31058,N_31223);
xnor U31500 (N_31500,N_31298,N_31353);
xnor U31501 (N_31501,N_31466,N_31492);
and U31502 (N_31502,N_31361,N_31380);
nand U31503 (N_31503,N_31384,N_31342);
or U31504 (N_31504,N_31407,N_31397);
xnor U31505 (N_31505,N_31474,N_31475);
or U31506 (N_31506,N_31365,N_31280);
and U31507 (N_31507,N_31458,N_31467);
nand U31508 (N_31508,N_31476,N_31269);
xnor U31509 (N_31509,N_31419,N_31303);
or U31510 (N_31510,N_31430,N_31473);
xor U31511 (N_31511,N_31322,N_31329);
and U31512 (N_31512,N_31477,N_31369);
nand U31513 (N_31513,N_31424,N_31441);
xnor U31514 (N_31514,N_31404,N_31325);
nor U31515 (N_31515,N_31381,N_31488);
nor U31516 (N_31516,N_31320,N_31406);
or U31517 (N_31517,N_31425,N_31330);
nor U31518 (N_31518,N_31388,N_31394);
and U31519 (N_31519,N_31251,N_31375);
xnor U31520 (N_31520,N_31376,N_31429);
and U31521 (N_31521,N_31343,N_31428);
nand U31522 (N_31522,N_31326,N_31440);
and U31523 (N_31523,N_31308,N_31378);
nand U31524 (N_31524,N_31347,N_31294);
nand U31525 (N_31525,N_31287,N_31420);
nor U31526 (N_31526,N_31447,N_31354);
xnor U31527 (N_31527,N_31297,N_31493);
nor U31528 (N_31528,N_31261,N_31254);
nand U31529 (N_31529,N_31334,N_31451);
and U31530 (N_31530,N_31283,N_31484);
nor U31531 (N_31531,N_31323,N_31469);
nand U31532 (N_31532,N_31457,N_31305);
and U31533 (N_31533,N_31485,N_31316);
nor U31534 (N_31534,N_31332,N_31299);
or U31535 (N_31535,N_31363,N_31417);
xnor U31536 (N_31536,N_31266,N_31393);
or U31537 (N_31537,N_31450,N_31437);
xnor U31538 (N_31538,N_31433,N_31482);
nand U31539 (N_31539,N_31495,N_31300);
or U31540 (N_31540,N_31403,N_31253);
xor U31541 (N_31541,N_31321,N_31351);
or U31542 (N_31542,N_31374,N_31324);
and U31543 (N_31543,N_31360,N_31355);
nand U31544 (N_31544,N_31465,N_31333);
or U31545 (N_31545,N_31278,N_31338);
nand U31546 (N_31546,N_31284,N_31263);
xor U31547 (N_31547,N_31344,N_31413);
and U31548 (N_31548,N_31348,N_31383);
and U31549 (N_31549,N_31389,N_31312);
and U31550 (N_31550,N_31277,N_31289);
xor U31551 (N_31551,N_31423,N_31445);
xnor U31552 (N_31552,N_31331,N_31496);
or U31553 (N_31553,N_31267,N_31454);
and U31554 (N_31554,N_31319,N_31398);
nand U31555 (N_31555,N_31391,N_31442);
or U31556 (N_31556,N_31314,N_31415);
and U31557 (N_31557,N_31260,N_31274);
or U31558 (N_31558,N_31282,N_31396);
nor U31559 (N_31559,N_31346,N_31499);
or U31560 (N_31560,N_31257,N_31327);
nand U31561 (N_31561,N_31352,N_31262);
xnor U31562 (N_31562,N_31358,N_31452);
xor U31563 (N_31563,N_31416,N_31498);
xnor U31564 (N_31564,N_31341,N_31273);
nand U31565 (N_31565,N_31411,N_31304);
and U31566 (N_31566,N_31453,N_31478);
or U31567 (N_31567,N_31456,N_31436);
xor U31568 (N_31568,N_31395,N_31311);
xnor U31569 (N_31569,N_31292,N_31318);
and U31570 (N_31570,N_31382,N_31408);
nor U31571 (N_31571,N_31336,N_31368);
and U31572 (N_31572,N_31310,N_31306);
nand U31573 (N_31573,N_31434,N_31276);
or U31574 (N_31574,N_31377,N_31446);
xor U31575 (N_31575,N_31410,N_31497);
and U31576 (N_31576,N_31448,N_31345);
and U31577 (N_31577,N_31443,N_31462);
or U31578 (N_31578,N_31431,N_31255);
and U31579 (N_31579,N_31252,N_31480);
xor U31580 (N_31580,N_31405,N_31399);
or U31581 (N_31581,N_31401,N_31422);
and U31582 (N_31582,N_31302,N_31455);
xor U31583 (N_31583,N_31444,N_31258);
nand U31584 (N_31584,N_31373,N_31421);
or U31585 (N_31585,N_31315,N_31486);
nor U31586 (N_31586,N_31460,N_31432);
nand U31587 (N_31587,N_31349,N_31402);
xor U31588 (N_31588,N_31390,N_31271);
xnor U31589 (N_31589,N_31288,N_31275);
xnor U31590 (N_31590,N_31350,N_31439);
and U31591 (N_31591,N_31412,N_31268);
nor U31592 (N_31592,N_31285,N_31470);
xor U31593 (N_31593,N_31464,N_31372);
and U31594 (N_31594,N_31291,N_31362);
xor U31595 (N_31595,N_31370,N_31264);
xnor U31596 (N_31596,N_31385,N_31392);
or U31597 (N_31597,N_31340,N_31293);
nor U31598 (N_31598,N_31418,N_31317);
xnor U31599 (N_31599,N_31270,N_31296);
nor U31600 (N_31600,N_31427,N_31471);
xnor U31601 (N_31601,N_31364,N_31371);
nand U31602 (N_31602,N_31468,N_31286);
xor U31603 (N_31603,N_31479,N_31463);
or U31604 (N_31604,N_31487,N_31265);
nand U31605 (N_31605,N_31438,N_31309);
nor U31606 (N_31606,N_31281,N_31359);
nand U31607 (N_31607,N_31367,N_31301);
xnor U31608 (N_31608,N_31357,N_31272);
and U31609 (N_31609,N_31313,N_31481);
and U31610 (N_31610,N_31494,N_31426);
and U31611 (N_31611,N_31356,N_31414);
xnor U31612 (N_31612,N_31250,N_31295);
nor U31613 (N_31613,N_31490,N_31256);
and U31614 (N_31614,N_31400,N_31290);
or U31615 (N_31615,N_31279,N_31461);
nand U31616 (N_31616,N_31409,N_31328);
nor U31617 (N_31617,N_31491,N_31459);
and U31618 (N_31618,N_31386,N_31472);
nor U31619 (N_31619,N_31489,N_31335);
and U31620 (N_31620,N_31337,N_31435);
and U31621 (N_31621,N_31339,N_31449);
nor U31622 (N_31622,N_31259,N_31483);
nand U31623 (N_31623,N_31379,N_31387);
nor U31624 (N_31624,N_31307,N_31366);
xor U31625 (N_31625,N_31494,N_31365);
nor U31626 (N_31626,N_31250,N_31394);
nand U31627 (N_31627,N_31414,N_31492);
or U31628 (N_31628,N_31257,N_31416);
nand U31629 (N_31629,N_31371,N_31425);
nand U31630 (N_31630,N_31446,N_31395);
and U31631 (N_31631,N_31428,N_31365);
and U31632 (N_31632,N_31259,N_31461);
and U31633 (N_31633,N_31348,N_31399);
xor U31634 (N_31634,N_31335,N_31394);
or U31635 (N_31635,N_31467,N_31283);
nand U31636 (N_31636,N_31330,N_31386);
xor U31637 (N_31637,N_31269,N_31332);
nand U31638 (N_31638,N_31481,N_31448);
nand U31639 (N_31639,N_31386,N_31426);
xor U31640 (N_31640,N_31362,N_31260);
and U31641 (N_31641,N_31485,N_31393);
or U31642 (N_31642,N_31397,N_31424);
or U31643 (N_31643,N_31486,N_31389);
nand U31644 (N_31644,N_31395,N_31416);
nor U31645 (N_31645,N_31481,N_31452);
nor U31646 (N_31646,N_31458,N_31435);
xor U31647 (N_31647,N_31495,N_31461);
nor U31648 (N_31648,N_31433,N_31446);
xor U31649 (N_31649,N_31314,N_31498);
or U31650 (N_31650,N_31494,N_31446);
nand U31651 (N_31651,N_31453,N_31365);
nand U31652 (N_31652,N_31463,N_31446);
nor U31653 (N_31653,N_31445,N_31304);
or U31654 (N_31654,N_31330,N_31482);
xor U31655 (N_31655,N_31426,N_31401);
xnor U31656 (N_31656,N_31418,N_31446);
xnor U31657 (N_31657,N_31461,N_31362);
nand U31658 (N_31658,N_31467,N_31268);
nand U31659 (N_31659,N_31260,N_31402);
nand U31660 (N_31660,N_31272,N_31462);
or U31661 (N_31661,N_31310,N_31262);
nand U31662 (N_31662,N_31400,N_31356);
nand U31663 (N_31663,N_31364,N_31457);
nand U31664 (N_31664,N_31362,N_31300);
and U31665 (N_31665,N_31407,N_31329);
or U31666 (N_31666,N_31300,N_31485);
nor U31667 (N_31667,N_31255,N_31375);
and U31668 (N_31668,N_31300,N_31316);
nor U31669 (N_31669,N_31458,N_31407);
xnor U31670 (N_31670,N_31277,N_31430);
xnor U31671 (N_31671,N_31427,N_31413);
or U31672 (N_31672,N_31356,N_31399);
nor U31673 (N_31673,N_31417,N_31268);
nor U31674 (N_31674,N_31463,N_31409);
or U31675 (N_31675,N_31264,N_31461);
nor U31676 (N_31676,N_31455,N_31328);
xnor U31677 (N_31677,N_31456,N_31329);
and U31678 (N_31678,N_31255,N_31488);
nand U31679 (N_31679,N_31465,N_31324);
or U31680 (N_31680,N_31452,N_31278);
and U31681 (N_31681,N_31252,N_31492);
nor U31682 (N_31682,N_31391,N_31425);
nand U31683 (N_31683,N_31405,N_31415);
nand U31684 (N_31684,N_31339,N_31311);
nand U31685 (N_31685,N_31351,N_31475);
or U31686 (N_31686,N_31280,N_31254);
xor U31687 (N_31687,N_31264,N_31334);
or U31688 (N_31688,N_31276,N_31347);
nor U31689 (N_31689,N_31277,N_31319);
nor U31690 (N_31690,N_31318,N_31313);
nor U31691 (N_31691,N_31414,N_31377);
nand U31692 (N_31692,N_31319,N_31475);
xnor U31693 (N_31693,N_31326,N_31379);
nor U31694 (N_31694,N_31343,N_31279);
or U31695 (N_31695,N_31486,N_31432);
or U31696 (N_31696,N_31371,N_31337);
nor U31697 (N_31697,N_31470,N_31437);
xor U31698 (N_31698,N_31408,N_31448);
or U31699 (N_31699,N_31379,N_31446);
and U31700 (N_31700,N_31324,N_31318);
and U31701 (N_31701,N_31255,N_31473);
or U31702 (N_31702,N_31374,N_31489);
nor U31703 (N_31703,N_31274,N_31291);
nand U31704 (N_31704,N_31274,N_31417);
or U31705 (N_31705,N_31404,N_31342);
nor U31706 (N_31706,N_31393,N_31343);
or U31707 (N_31707,N_31384,N_31416);
nand U31708 (N_31708,N_31295,N_31438);
xnor U31709 (N_31709,N_31342,N_31316);
or U31710 (N_31710,N_31340,N_31287);
and U31711 (N_31711,N_31368,N_31463);
nor U31712 (N_31712,N_31389,N_31285);
nand U31713 (N_31713,N_31273,N_31261);
nand U31714 (N_31714,N_31315,N_31300);
and U31715 (N_31715,N_31463,N_31378);
or U31716 (N_31716,N_31354,N_31390);
or U31717 (N_31717,N_31375,N_31425);
or U31718 (N_31718,N_31296,N_31475);
nand U31719 (N_31719,N_31356,N_31448);
nand U31720 (N_31720,N_31313,N_31460);
and U31721 (N_31721,N_31376,N_31480);
and U31722 (N_31722,N_31481,N_31261);
nand U31723 (N_31723,N_31457,N_31437);
nor U31724 (N_31724,N_31362,N_31303);
nand U31725 (N_31725,N_31300,N_31404);
nor U31726 (N_31726,N_31256,N_31483);
and U31727 (N_31727,N_31311,N_31259);
xor U31728 (N_31728,N_31330,N_31280);
and U31729 (N_31729,N_31439,N_31411);
nand U31730 (N_31730,N_31321,N_31354);
or U31731 (N_31731,N_31260,N_31475);
and U31732 (N_31732,N_31308,N_31453);
and U31733 (N_31733,N_31364,N_31251);
or U31734 (N_31734,N_31340,N_31397);
nor U31735 (N_31735,N_31357,N_31492);
and U31736 (N_31736,N_31364,N_31293);
and U31737 (N_31737,N_31490,N_31389);
nor U31738 (N_31738,N_31456,N_31280);
nor U31739 (N_31739,N_31449,N_31442);
xnor U31740 (N_31740,N_31372,N_31488);
nand U31741 (N_31741,N_31282,N_31260);
nor U31742 (N_31742,N_31467,N_31400);
nand U31743 (N_31743,N_31349,N_31453);
nand U31744 (N_31744,N_31273,N_31352);
xor U31745 (N_31745,N_31489,N_31433);
xor U31746 (N_31746,N_31414,N_31383);
nor U31747 (N_31747,N_31262,N_31459);
or U31748 (N_31748,N_31306,N_31288);
xor U31749 (N_31749,N_31329,N_31375);
xor U31750 (N_31750,N_31591,N_31575);
or U31751 (N_31751,N_31518,N_31505);
xor U31752 (N_31752,N_31695,N_31698);
xor U31753 (N_31753,N_31665,N_31623);
nand U31754 (N_31754,N_31707,N_31712);
nor U31755 (N_31755,N_31603,N_31585);
xor U31756 (N_31756,N_31721,N_31554);
xnor U31757 (N_31757,N_31602,N_31634);
xor U31758 (N_31758,N_31744,N_31731);
xor U31759 (N_31759,N_31613,N_31599);
and U31760 (N_31760,N_31746,N_31523);
or U31761 (N_31761,N_31558,N_31749);
and U31762 (N_31762,N_31565,N_31573);
nand U31763 (N_31763,N_31525,N_31535);
or U31764 (N_31764,N_31670,N_31552);
xor U31765 (N_31765,N_31600,N_31657);
nand U31766 (N_31766,N_31546,N_31606);
xor U31767 (N_31767,N_31740,N_31519);
xnor U31768 (N_31768,N_31550,N_31640);
nand U31769 (N_31769,N_31693,N_31516);
nor U31770 (N_31770,N_31564,N_31524);
nor U31771 (N_31771,N_31563,N_31651);
nand U31772 (N_31772,N_31675,N_31580);
nor U31773 (N_31773,N_31539,N_31582);
and U31774 (N_31774,N_31714,N_31612);
nand U31775 (N_31775,N_31742,N_31646);
xnor U31776 (N_31776,N_31589,N_31534);
nand U31777 (N_31777,N_31512,N_31619);
nor U31778 (N_31778,N_31687,N_31562);
nand U31779 (N_31779,N_31653,N_31551);
and U31780 (N_31780,N_31709,N_31700);
or U31781 (N_31781,N_31608,N_31584);
nand U31782 (N_31782,N_31655,N_31520);
nor U31783 (N_31783,N_31542,N_31701);
nand U31784 (N_31784,N_31737,N_31574);
nand U31785 (N_31785,N_31622,N_31579);
nor U31786 (N_31786,N_31652,N_31664);
and U31787 (N_31787,N_31681,N_31596);
and U31788 (N_31788,N_31560,N_31691);
or U31789 (N_31789,N_31632,N_31631);
xor U31790 (N_31790,N_31511,N_31702);
nand U31791 (N_31791,N_31654,N_31706);
nand U31792 (N_31792,N_31604,N_31607);
xor U31793 (N_31793,N_31671,N_31504);
nand U31794 (N_31794,N_31548,N_31747);
and U31795 (N_31795,N_31650,N_31645);
or U31796 (N_31796,N_31696,N_31583);
xnor U31797 (N_31797,N_31557,N_31588);
xnor U31798 (N_31798,N_31628,N_31724);
or U31799 (N_31799,N_31643,N_31748);
xnor U31800 (N_31800,N_31649,N_31629);
nor U31801 (N_31801,N_31532,N_31609);
and U31802 (N_31802,N_31630,N_31537);
xor U31803 (N_31803,N_31559,N_31644);
and U31804 (N_31804,N_31533,N_31704);
nor U31805 (N_31805,N_31605,N_31692);
or U31806 (N_31806,N_31528,N_31586);
or U31807 (N_31807,N_31662,N_31745);
nand U31808 (N_31808,N_31581,N_31699);
nand U31809 (N_31809,N_31517,N_31572);
nor U31810 (N_31810,N_31708,N_31728);
nand U31811 (N_31811,N_31647,N_31726);
nand U31812 (N_31812,N_31686,N_31587);
nand U31813 (N_31813,N_31680,N_31509);
or U31814 (N_31814,N_31642,N_31648);
and U31815 (N_31815,N_31732,N_31531);
xor U31816 (N_31816,N_31510,N_31635);
nor U31817 (N_31817,N_31667,N_31641);
nor U31818 (N_31818,N_31624,N_31618);
and U31819 (N_31819,N_31536,N_31636);
or U31820 (N_31820,N_31679,N_31555);
nor U31821 (N_31821,N_31567,N_31719);
xnor U31822 (N_31822,N_31717,N_31727);
or U31823 (N_31823,N_31741,N_31595);
xnor U31824 (N_31824,N_31625,N_31514);
xnor U31825 (N_31825,N_31570,N_31673);
nand U31826 (N_31826,N_31729,N_31601);
nor U31827 (N_31827,N_31716,N_31666);
or U31828 (N_31828,N_31627,N_31522);
nand U31829 (N_31829,N_31538,N_31713);
or U31830 (N_31830,N_31598,N_31569);
nand U31831 (N_31831,N_31690,N_31730);
and U31832 (N_31832,N_31617,N_31529);
or U31833 (N_31833,N_31566,N_31659);
xnor U31834 (N_31834,N_31683,N_31568);
xor U31835 (N_31835,N_31610,N_31658);
nand U31836 (N_31836,N_31725,N_31743);
and U31837 (N_31837,N_31736,N_31685);
or U31838 (N_31838,N_31543,N_31722);
xor U31839 (N_31839,N_31615,N_31526);
xnor U31840 (N_31840,N_31638,N_31739);
nand U31841 (N_31841,N_31500,N_31689);
xor U31842 (N_31842,N_31668,N_31592);
xnor U31843 (N_31843,N_31571,N_31672);
and U31844 (N_31844,N_31656,N_31549);
xor U31845 (N_31845,N_31710,N_31633);
nor U31846 (N_31846,N_31507,N_31614);
xor U31847 (N_31847,N_31547,N_31723);
and U31848 (N_31848,N_31578,N_31711);
and U31849 (N_31849,N_31734,N_31521);
or U31850 (N_31850,N_31501,N_31684);
xor U31851 (N_31851,N_31738,N_31694);
xor U31852 (N_31852,N_31720,N_31576);
and U31853 (N_31853,N_31527,N_31682);
nor U31854 (N_31854,N_31735,N_31513);
xor U31855 (N_31855,N_31688,N_31669);
and U31856 (N_31856,N_31621,N_31597);
or U31857 (N_31857,N_31661,N_31502);
and U31858 (N_31858,N_31611,N_31674);
and U31859 (N_31859,N_31540,N_31541);
and U31860 (N_31860,N_31545,N_31715);
xor U31861 (N_31861,N_31553,N_31637);
nand U31862 (N_31862,N_31590,N_31660);
and U31863 (N_31863,N_31676,N_31626);
and U31864 (N_31864,N_31733,N_31506);
nor U31865 (N_31865,N_31530,N_31703);
nor U31866 (N_31866,N_31561,N_31663);
nand U31867 (N_31867,N_31577,N_31620);
nand U31868 (N_31868,N_31556,N_31678);
or U31869 (N_31869,N_31718,N_31515);
xor U31870 (N_31870,N_31705,N_31639);
nand U31871 (N_31871,N_31593,N_31697);
nor U31872 (N_31872,N_31544,N_31616);
nor U31873 (N_31873,N_31594,N_31503);
or U31874 (N_31874,N_31677,N_31508);
or U31875 (N_31875,N_31584,N_31632);
and U31876 (N_31876,N_31687,N_31691);
and U31877 (N_31877,N_31520,N_31568);
nor U31878 (N_31878,N_31707,N_31559);
nor U31879 (N_31879,N_31618,N_31670);
xor U31880 (N_31880,N_31592,N_31589);
xnor U31881 (N_31881,N_31507,N_31564);
nand U31882 (N_31882,N_31640,N_31649);
nor U31883 (N_31883,N_31503,N_31544);
xor U31884 (N_31884,N_31702,N_31683);
nand U31885 (N_31885,N_31583,N_31646);
and U31886 (N_31886,N_31708,N_31525);
nor U31887 (N_31887,N_31731,N_31517);
xnor U31888 (N_31888,N_31654,N_31704);
and U31889 (N_31889,N_31644,N_31661);
nand U31890 (N_31890,N_31623,N_31595);
nand U31891 (N_31891,N_31539,N_31594);
nor U31892 (N_31892,N_31664,N_31689);
xnor U31893 (N_31893,N_31686,N_31590);
nor U31894 (N_31894,N_31686,N_31617);
or U31895 (N_31895,N_31706,N_31716);
and U31896 (N_31896,N_31670,N_31707);
nor U31897 (N_31897,N_31681,N_31735);
nor U31898 (N_31898,N_31542,N_31737);
and U31899 (N_31899,N_31584,N_31541);
nand U31900 (N_31900,N_31561,N_31524);
nand U31901 (N_31901,N_31697,N_31694);
and U31902 (N_31902,N_31620,N_31576);
and U31903 (N_31903,N_31582,N_31597);
or U31904 (N_31904,N_31510,N_31714);
and U31905 (N_31905,N_31570,N_31737);
xnor U31906 (N_31906,N_31638,N_31717);
xor U31907 (N_31907,N_31633,N_31657);
nor U31908 (N_31908,N_31701,N_31727);
and U31909 (N_31909,N_31715,N_31687);
xor U31910 (N_31910,N_31576,N_31664);
nor U31911 (N_31911,N_31617,N_31642);
nand U31912 (N_31912,N_31690,N_31655);
nor U31913 (N_31913,N_31668,N_31604);
and U31914 (N_31914,N_31688,N_31665);
nand U31915 (N_31915,N_31553,N_31670);
nor U31916 (N_31916,N_31688,N_31541);
xor U31917 (N_31917,N_31733,N_31541);
xor U31918 (N_31918,N_31576,N_31693);
nand U31919 (N_31919,N_31680,N_31609);
nand U31920 (N_31920,N_31543,N_31749);
nor U31921 (N_31921,N_31706,N_31585);
or U31922 (N_31922,N_31530,N_31746);
nor U31923 (N_31923,N_31548,N_31537);
xnor U31924 (N_31924,N_31511,N_31549);
and U31925 (N_31925,N_31704,N_31564);
nor U31926 (N_31926,N_31720,N_31662);
and U31927 (N_31927,N_31654,N_31743);
xor U31928 (N_31928,N_31609,N_31530);
or U31929 (N_31929,N_31524,N_31576);
and U31930 (N_31930,N_31596,N_31621);
nand U31931 (N_31931,N_31691,N_31606);
nor U31932 (N_31932,N_31749,N_31624);
or U31933 (N_31933,N_31511,N_31543);
and U31934 (N_31934,N_31537,N_31532);
nor U31935 (N_31935,N_31650,N_31653);
and U31936 (N_31936,N_31680,N_31731);
nor U31937 (N_31937,N_31671,N_31587);
and U31938 (N_31938,N_31644,N_31741);
xnor U31939 (N_31939,N_31720,N_31625);
and U31940 (N_31940,N_31701,N_31567);
or U31941 (N_31941,N_31652,N_31599);
and U31942 (N_31942,N_31669,N_31525);
and U31943 (N_31943,N_31519,N_31502);
nor U31944 (N_31944,N_31514,N_31582);
or U31945 (N_31945,N_31560,N_31546);
and U31946 (N_31946,N_31645,N_31608);
nor U31947 (N_31947,N_31625,N_31539);
nand U31948 (N_31948,N_31736,N_31728);
xor U31949 (N_31949,N_31737,N_31626);
nand U31950 (N_31950,N_31626,N_31636);
or U31951 (N_31951,N_31705,N_31555);
and U31952 (N_31952,N_31718,N_31726);
xor U31953 (N_31953,N_31720,N_31681);
nand U31954 (N_31954,N_31578,N_31741);
nor U31955 (N_31955,N_31730,N_31514);
or U31956 (N_31956,N_31579,N_31712);
nor U31957 (N_31957,N_31627,N_31609);
nand U31958 (N_31958,N_31719,N_31706);
xnor U31959 (N_31959,N_31737,N_31651);
and U31960 (N_31960,N_31724,N_31546);
and U31961 (N_31961,N_31580,N_31699);
and U31962 (N_31962,N_31617,N_31536);
nor U31963 (N_31963,N_31556,N_31668);
nor U31964 (N_31964,N_31548,N_31570);
and U31965 (N_31965,N_31647,N_31629);
nor U31966 (N_31966,N_31576,N_31705);
xor U31967 (N_31967,N_31713,N_31593);
nand U31968 (N_31968,N_31528,N_31653);
or U31969 (N_31969,N_31500,N_31592);
and U31970 (N_31970,N_31576,N_31535);
xnor U31971 (N_31971,N_31571,N_31546);
nand U31972 (N_31972,N_31575,N_31730);
xnor U31973 (N_31973,N_31697,N_31582);
and U31974 (N_31974,N_31621,N_31613);
or U31975 (N_31975,N_31720,N_31728);
nand U31976 (N_31976,N_31705,N_31744);
nand U31977 (N_31977,N_31699,N_31727);
nand U31978 (N_31978,N_31560,N_31694);
xor U31979 (N_31979,N_31656,N_31677);
or U31980 (N_31980,N_31695,N_31625);
nand U31981 (N_31981,N_31562,N_31538);
nor U31982 (N_31982,N_31648,N_31586);
xnor U31983 (N_31983,N_31508,N_31607);
or U31984 (N_31984,N_31632,N_31503);
and U31985 (N_31985,N_31616,N_31714);
xor U31986 (N_31986,N_31562,N_31581);
and U31987 (N_31987,N_31723,N_31722);
xnor U31988 (N_31988,N_31544,N_31718);
or U31989 (N_31989,N_31715,N_31718);
and U31990 (N_31990,N_31577,N_31536);
xnor U31991 (N_31991,N_31728,N_31688);
xor U31992 (N_31992,N_31623,N_31730);
nand U31993 (N_31993,N_31676,N_31678);
xnor U31994 (N_31994,N_31659,N_31586);
xor U31995 (N_31995,N_31645,N_31603);
nand U31996 (N_31996,N_31671,N_31727);
or U31997 (N_31997,N_31520,N_31608);
or U31998 (N_31998,N_31584,N_31513);
and U31999 (N_31999,N_31659,N_31563);
and U32000 (N_32000,N_31886,N_31995);
xor U32001 (N_32001,N_31892,N_31985);
xor U32002 (N_32002,N_31891,N_31823);
nand U32003 (N_32003,N_31988,N_31820);
nor U32004 (N_32004,N_31797,N_31944);
xnor U32005 (N_32005,N_31909,N_31761);
and U32006 (N_32006,N_31812,N_31830);
or U32007 (N_32007,N_31868,N_31908);
nor U32008 (N_32008,N_31941,N_31772);
nand U32009 (N_32009,N_31914,N_31816);
nand U32010 (N_32010,N_31850,N_31825);
xor U32011 (N_32011,N_31884,N_31976);
nand U32012 (N_32012,N_31873,N_31752);
xnor U32013 (N_32013,N_31800,N_31813);
nand U32014 (N_32014,N_31801,N_31763);
nor U32015 (N_32015,N_31770,N_31915);
and U32016 (N_32016,N_31781,N_31848);
nand U32017 (N_32017,N_31880,N_31836);
xor U32018 (N_32018,N_31981,N_31856);
xnor U32019 (N_32019,N_31968,N_31936);
xor U32020 (N_32020,N_31771,N_31977);
and U32021 (N_32021,N_31997,N_31765);
or U32022 (N_32022,N_31948,N_31955);
and U32023 (N_32023,N_31972,N_31792);
xor U32024 (N_32024,N_31924,N_31827);
and U32025 (N_32025,N_31863,N_31951);
xnor U32026 (N_32026,N_31773,N_31853);
nor U32027 (N_32027,N_31932,N_31804);
nor U32028 (N_32028,N_31893,N_31987);
nand U32029 (N_32029,N_31845,N_31885);
xor U32030 (N_32030,N_31831,N_31808);
nand U32031 (N_32031,N_31938,N_31998);
xor U32032 (N_32032,N_31787,N_31990);
nand U32033 (N_32033,N_31922,N_31837);
nor U32034 (N_32034,N_31978,N_31815);
xnor U32035 (N_32035,N_31961,N_31790);
or U32036 (N_32036,N_31973,N_31878);
xnor U32037 (N_32037,N_31942,N_31777);
or U32038 (N_32038,N_31791,N_31925);
or U32039 (N_32039,N_31965,N_31992);
nand U32040 (N_32040,N_31994,N_31774);
nor U32041 (N_32041,N_31946,N_31835);
nand U32042 (N_32042,N_31959,N_31940);
xnor U32043 (N_32043,N_31905,N_31846);
xor U32044 (N_32044,N_31866,N_31785);
nand U32045 (N_32045,N_31963,N_31962);
or U32046 (N_32046,N_31766,N_31903);
or U32047 (N_32047,N_31964,N_31859);
and U32048 (N_32048,N_31764,N_31969);
xor U32049 (N_32049,N_31960,N_31876);
and U32050 (N_32050,N_31916,N_31796);
nor U32051 (N_32051,N_31755,N_31814);
xnor U32052 (N_32052,N_31887,N_31996);
and U32053 (N_32053,N_31828,N_31867);
nand U32054 (N_32054,N_31810,N_31970);
or U32055 (N_32055,N_31919,N_31906);
nand U32056 (N_32056,N_31953,N_31881);
nor U32057 (N_32057,N_31871,N_31849);
and U32058 (N_32058,N_31933,N_31847);
and U32059 (N_32059,N_31947,N_31930);
and U32060 (N_32060,N_31901,N_31842);
nand U32061 (N_32061,N_31894,N_31890);
and U32062 (N_32062,N_31860,N_31870);
or U32063 (N_32063,N_31883,N_31805);
nor U32064 (N_32064,N_31769,N_31979);
nor U32065 (N_32065,N_31819,N_31935);
and U32066 (N_32066,N_31911,N_31897);
nand U32067 (N_32067,N_31851,N_31754);
and U32068 (N_32068,N_31945,N_31896);
xnor U32069 (N_32069,N_31879,N_31753);
nor U32070 (N_32070,N_31923,N_31966);
and U32071 (N_32071,N_31840,N_31877);
xnor U32072 (N_32072,N_31907,N_31864);
and U32073 (N_32073,N_31928,N_31931);
xnor U32074 (N_32074,N_31875,N_31821);
nand U32075 (N_32075,N_31759,N_31900);
or U32076 (N_32076,N_31934,N_31854);
xor U32077 (N_32077,N_31760,N_31829);
nand U32078 (N_32078,N_31809,N_31844);
and U32079 (N_32079,N_31874,N_31950);
or U32080 (N_32080,N_31902,N_31912);
or U32081 (N_32081,N_31824,N_31986);
or U32082 (N_32082,N_31852,N_31768);
nor U32083 (N_32083,N_31794,N_31982);
nor U32084 (N_32084,N_31855,N_31807);
or U32085 (N_32085,N_31975,N_31802);
nand U32086 (N_32086,N_31958,N_31949);
xnor U32087 (N_32087,N_31782,N_31952);
nand U32088 (N_32088,N_31869,N_31775);
nand U32089 (N_32089,N_31898,N_31889);
or U32090 (N_32090,N_31939,N_31806);
and U32091 (N_32091,N_31917,N_31750);
and U32092 (N_32092,N_31793,N_31882);
or U32093 (N_32093,N_31904,N_31984);
nand U32094 (N_32094,N_31993,N_31920);
nand U32095 (N_32095,N_31872,N_31834);
or U32096 (N_32096,N_31756,N_31957);
xor U32097 (N_32097,N_31913,N_31788);
and U32098 (N_32098,N_31784,N_31817);
nor U32099 (N_32099,N_31778,N_31974);
or U32100 (N_32100,N_31811,N_31991);
nor U32101 (N_32101,N_31971,N_31803);
nor U32102 (N_32102,N_31822,N_31943);
xnor U32103 (N_32103,N_31918,N_31799);
xnor U32104 (N_32104,N_31798,N_31956);
xor U32105 (N_32105,N_31862,N_31789);
and U32106 (N_32106,N_31888,N_31954);
or U32107 (N_32107,N_31865,N_31832);
or U32108 (N_32108,N_31937,N_31818);
nor U32109 (N_32109,N_31762,N_31841);
nand U32110 (N_32110,N_31899,N_31861);
and U32111 (N_32111,N_31910,N_31926);
nand U32112 (N_32112,N_31843,N_31826);
nor U32113 (N_32113,N_31795,N_31980);
and U32114 (N_32114,N_31967,N_31751);
xor U32115 (N_32115,N_31989,N_31767);
or U32116 (N_32116,N_31783,N_31786);
nor U32117 (N_32117,N_31758,N_31776);
nor U32118 (N_32118,N_31780,N_31999);
nand U32119 (N_32119,N_31895,N_31927);
nor U32120 (N_32120,N_31833,N_31858);
xnor U32121 (N_32121,N_31838,N_31857);
nand U32122 (N_32122,N_31757,N_31921);
nand U32123 (N_32123,N_31929,N_31983);
and U32124 (N_32124,N_31779,N_31839);
and U32125 (N_32125,N_31852,N_31969);
xor U32126 (N_32126,N_31806,N_31885);
xnor U32127 (N_32127,N_31765,N_31975);
and U32128 (N_32128,N_31913,N_31976);
xor U32129 (N_32129,N_31775,N_31878);
nand U32130 (N_32130,N_31978,N_31937);
or U32131 (N_32131,N_31942,N_31922);
nand U32132 (N_32132,N_31875,N_31752);
and U32133 (N_32133,N_31924,N_31813);
xor U32134 (N_32134,N_31981,N_31798);
nor U32135 (N_32135,N_31751,N_31860);
and U32136 (N_32136,N_31815,N_31794);
xnor U32137 (N_32137,N_31858,N_31961);
or U32138 (N_32138,N_31757,N_31972);
nor U32139 (N_32139,N_31860,N_31919);
nand U32140 (N_32140,N_31761,N_31778);
and U32141 (N_32141,N_31828,N_31834);
or U32142 (N_32142,N_31805,N_31999);
xor U32143 (N_32143,N_31768,N_31801);
xnor U32144 (N_32144,N_31969,N_31869);
and U32145 (N_32145,N_31871,N_31817);
and U32146 (N_32146,N_31958,N_31758);
nand U32147 (N_32147,N_31911,N_31842);
or U32148 (N_32148,N_31801,N_31853);
nand U32149 (N_32149,N_31930,N_31793);
xnor U32150 (N_32150,N_31881,N_31982);
nand U32151 (N_32151,N_31955,N_31848);
and U32152 (N_32152,N_31989,N_31904);
and U32153 (N_32153,N_31856,N_31905);
or U32154 (N_32154,N_31874,N_31775);
or U32155 (N_32155,N_31904,N_31780);
nor U32156 (N_32156,N_31756,N_31964);
and U32157 (N_32157,N_31921,N_31937);
nor U32158 (N_32158,N_31989,N_31844);
xor U32159 (N_32159,N_31872,N_31795);
nor U32160 (N_32160,N_31859,N_31895);
xor U32161 (N_32161,N_31842,N_31844);
nor U32162 (N_32162,N_31876,N_31852);
or U32163 (N_32163,N_31975,N_31865);
xor U32164 (N_32164,N_31791,N_31919);
or U32165 (N_32165,N_31881,N_31753);
xnor U32166 (N_32166,N_31922,N_31989);
nor U32167 (N_32167,N_31920,N_31759);
xnor U32168 (N_32168,N_31933,N_31755);
xor U32169 (N_32169,N_31814,N_31957);
nand U32170 (N_32170,N_31880,N_31794);
or U32171 (N_32171,N_31756,N_31901);
xnor U32172 (N_32172,N_31791,N_31780);
nor U32173 (N_32173,N_31759,N_31789);
nand U32174 (N_32174,N_31767,N_31808);
nand U32175 (N_32175,N_31974,N_31871);
nor U32176 (N_32176,N_31902,N_31986);
nand U32177 (N_32177,N_31862,N_31810);
nand U32178 (N_32178,N_31853,N_31761);
nor U32179 (N_32179,N_31868,N_31943);
and U32180 (N_32180,N_31773,N_31908);
nor U32181 (N_32181,N_31859,N_31937);
nor U32182 (N_32182,N_31957,N_31760);
and U32183 (N_32183,N_31883,N_31999);
nand U32184 (N_32184,N_31762,N_31986);
xnor U32185 (N_32185,N_31965,N_31894);
or U32186 (N_32186,N_31813,N_31923);
nor U32187 (N_32187,N_31860,N_31760);
xor U32188 (N_32188,N_31807,N_31864);
nand U32189 (N_32189,N_31937,N_31850);
or U32190 (N_32190,N_31925,N_31832);
or U32191 (N_32191,N_31791,N_31838);
nor U32192 (N_32192,N_31985,N_31886);
nor U32193 (N_32193,N_31816,N_31909);
nor U32194 (N_32194,N_31860,N_31974);
nand U32195 (N_32195,N_31864,N_31868);
and U32196 (N_32196,N_31759,N_31889);
xor U32197 (N_32197,N_31840,N_31818);
xnor U32198 (N_32198,N_31939,N_31917);
xor U32199 (N_32199,N_31970,N_31973);
and U32200 (N_32200,N_31898,N_31978);
nand U32201 (N_32201,N_31911,N_31926);
xnor U32202 (N_32202,N_31936,N_31992);
nand U32203 (N_32203,N_31887,N_31879);
and U32204 (N_32204,N_31911,N_31885);
xnor U32205 (N_32205,N_31985,N_31926);
or U32206 (N_32206,N_31790,N_31821);
nor U32207 (N_32207,N_31774,N_31923);
nor U32208 (N_32208,N_31879,N_31848);
or U32209 (N_32209,N_31847,N_31950);
and U32210 (N_32210,N_31890,N_31942);
xor U32211 (N_32211,N_31832,N_31986);
xnor U32212 (N_32212,N_31971,N_31869);
nand U32213 (N_32213,N_31818,N_31867);
xnor U32214 (N_32214,N_31941,N_31924);
nor U32215 (N_32215,N_31893,N_31997);
nor U32216 (N_32216,N_31765,N_31870);
nand U32217 (N_32217,N_31881,N_31927);
nor U32218 (N_32218,N_31757,N_31901);
nor U32219 (N_32219,N_31830,N_31920);
or U32220 (N_32220,N_31919,N_31833);
xnor U32221 (N_32221,N_31874,N_31944);
xor U32222 (N_32222,N_31893,N_31915);
nor U32223 (N_32223,N_31875,N_31816);
nor U32224 (N_32224,N_31771,N_31904);
and U32225 (N_32225,N_31803,N_31917);
xnor U32226 (N_32226,N_31770,N_31992);
or U32227 (N_32227,N_31992,N_31937);
or U32228 (N_32228,N_31966,N_31785);
and U32229 (N_32229,N_31797,N_31750);
or U32230 (N_32230,N_31984,N_31825);
and U32231 (N_32231,N_31974,N_31910);
nor U32232 (N_32232,N_31929,N_31801);
nor U32233 (N_32233,N_31825,N_31979);
and U32234 (N_32234,N_31853,N_31881);
nand U32235 (N_32235,N_31788,N_31930);
nor U32236 (N_32236,N_31999,N_31977);
nand U32237 (N_32237,N_31998,N_31968);
xnor U32238 (N_32238,N_31987,N_31926);
or U32239 (N_32239,N_31933,N_31985);
nand U32240 (N_32240,N_31809,N_31865);
nand U32241 (N_32241,N_31787,N_31923);
or U32242 (N_32242,N_31823,N_31969);
and U32243 (N_32243,N_31820,N_31999);
nor U32244 (N_32244,N_31857,N_31969);
xnor U32245 (N_32245,N_31790,N_31990);
and U32246 (N_32246,N_31757,N_31995);
nor U32247 (N_32247,N_31780,N_31858);
nor U32248 (N_32248,N_31847,N_31887);
nor U32249 (N_32249,N_31835,N_31918);
nor U32250 (N_32250,N_32144,N_32165);
and U32251 (N_32251,N_32094,N_32171);
nand U32252 (N_32252,N_32107,N_32003);
and U32253 (N_32253,N_32093,N_32245);
nor U32254 (N_32254,N_32157,N_32080);
or U32255 (N_32255,N_32132,N_32065);
and U32256 (N_32256,N_32062,N_32191);
xnor U32257 (N_32257,N_32007,N_32148);
nor U32258 (N_32258,N_32208,N_32218);
nor U32259 (N_32259,N_32002,N_32237);
xnor U32260 (N_32260,N_32209,N_32089);
xnor U32261 (N_32261,N_32142,N_32083);
nor U32262 (N_32262,N_32185,N_32225);
xor U32263 (N_32263,N_32044,N_32195);
and U32264 (N_32264,N_32217,N_32096);
nor U32265 (N_32265,N_32121,N_32162);
or U32266 (N_32266,N_32203,N_32126);
or U32267 (N_32267,N_32239,N_32196);
nor U32268 (N_32268,N_32169,N_32134);
and U32269 (N_32269,N_32108,N_32084);
or U32270 (N_32270,N_32075,N_32155);
and U32271 (N_32271,N_32127,N_32056);
nand U32272 (N_32272,N_32248,N_32151);
xor U32273 (N_32273,N_32106,N_32078);
xor U32274 (N_32274,N_32207,N_32175);
nand U32275 (N_32275,N_32043,N_32079);
or U32276 (N_32276,N_32058,N_32051);
or U32277 (N_32277,N_32041,N_32098);
nand U32278 (N_32278,N_32066,N_32205);
and U32279 (N_32279,N_32221,N_32130);
and U32280 (N_32280,N_32071,N_32244);
or U32281 (N_32281,N_32045,N_32211);
nor U32282 (N_32282,N_32095,N_32109);
and U32283 (N_32283,N_32215,N_32116);
nand U32284 (N_32284,N_32183,N_32088);
nand U32285 (N_32285,N_32189,N_32230);
nand U32286 (N_32286,N_32010,N_32133);
and U32287 (N_32287,N_32087,N_32216);
nand U32288 (N_32288,N_32050,N_32223);
nand U32289 (N_32289,N_32009,N_32020);
nand U32290 (N_32290,N_32064,N_32068);
nor U32291 (N_32291,N_32160,N_32081);
and U32292 (N_32292,N_32170,N_32188);
xor U32293 (N_32293,N_32114,N_32105);
nand U32294 (N_32294,N_32000,N_32037);
and U32295 (N_32295,N_32152,N_32057);
nor U32296 (N_32296,N_32053,N_32243);
and U32297 (N_32297,N_32159,N_32115);
nand U32298 (N_32298,N_32186,N_32073);
or U32299 (N_32299,N_32011,N_32032);
nor U32300 (N_32300,N_32219,N_32101);
and U32301 (N_32301,N_32125,N_32097);
or U32302 (N_32302,N_32240,N_32061);
and U32303 (N_32303,N_32118,N_32140);
nor U32304 (N_32304,N_32055,N_32220);
xnor U32305 (N_32305,N_32092,N_32236);
nand U32306 (N_32306,N_32103,N_32222);
or U32307 (N_32307,N_32163,N_32131);
or U32308 (N_32308,N_32076,N_32104);
or U32309 (N_32309,N_32172,N_32113);
xnor U32310 (N_32310,N_32168,N_32201);
xor U32311 (N_32311,N_32138,N_32005);
xor U32312 (N_32312,N_32085,N_32039);
xnor U32313 (N_32313,N_32204,N_32069);
xor U32314 (N_32314,N_32004,N_32102);
nor U32315 (N_32315,N_32174,N_32090);
nor U32316 (N_32316,N_32154,N_32197);
xnor U32317 (N_32317,N_32123,N_32070);
or U32318 (N_32318,N_32137,N_32120);
xor U32319 (N_32319,N_32246,N_32178);
and U32320 (N_32320,N_32141,N_32086);
nand U32321 (N_32321,N_32153,N_32200);
xnor U32322 (N_32322,N_32112,N_32136);
xor U32323 (N_32323,N_32021,N_32206);
xor U32324 (N_32324,N_32117,N_32014);
xnor U32325 (N_32325,N_32158,N_32119);
xnor U32326 (N_32326,N_32166,N_32226);
nand U32327 (N_32327,N_32028,N_32006);
xor U32328 (N_32328,N_32234,N_32035);
or U32329 (N_32329,N_32099,N_32235);
nand U32330 (N_32330,N_32023,N_32143);
and U32331 (N_32331,N_32231,N_32048);
xor U32332 (N_32332,N_32135,N_32022);
xor U32333 (N_32333,N_32012,N_32192);
xnor U32334 (N_32334,N_32124,N_32031);
xor U32335 (N_32335,N_32129,N_32190);
and U32336 (N_32336,N_32173,N_32038);
nand U32337 (N_32337,N_32150,N_32214);
nor U32338 (N_32338,N_32161,N_32074);
nand U32339 (N_32339,N_32180,N_32018);
nand U32340 (N_32340,N_32008,N_32111);
and U32341 (N_32341,N_32001,N_32026);
xor U32342 (N_32342,N_32149,N_32210);
and U32343 (N_32343,N_32242,N_32034);
or U32344 (N_32344,N_32224,N_32040);
nor U32345 (N_32345,N_32077,N_32241);
nand U32346 (N_32346,N_32060,N_32063);
or U32347 (N_32347,N_32030,N_32049);
and U32348 (N_32348,N_32199,N_32091);
xnor U32349 (N_32349,N_32013,N_32042);
nand U32350 (N_32350,N_32233,N_32100);
and U32351 (N_32351,N_32019,N_32025);
or U32352 (N_32352,N_32016,N_32247);
nor U32353 (N_32353,N_32194,N_32128);
nor U32354 (N_32354,N_32229,N_32145);
xor U32355 (N_32355,N_32072,N_32033);
nand U32356 (N_32356,N_32024,N_32213);
or U32357 (N_32357,N_32027,N_32198);
xnor U32358 (N_32358,N_32164,N_32187);
or U32359 (N_32359,N_32036,N_32212);
nor U32360 (N_32360,N_32193,N_32177);
or U32361 (N_32361,N_32015,N_32238);
nand U32362 (N_32362,N_32046,N_32067);
nand U32363 (N_32363,N_32059,N_32146);
xnor U32364 (N_32364,N_32249,N_32122);
or U32365 (N_32365,N_32179,N_32202);
nand U32366 (N_32366,N_32156,N_32047);
xnor U32367 (N_32367,N_32181,N_32017);
nand U32368 (N_32368,N_32082,N_32232);
nand U32369 (N_32369,N_32139,N_32110);
xor U32370 (N_32370,N_32184,N_32054);
nor U32371 (N_32371,N_32176,N_32147);
nand U32372 (N_32372,N_32228,N_32052);
nor U32373 (N_32373,N_32227,N_32167);
xnor U32374 (N_32374,N_32029,N_32182);
nor U32375 (N_32375,N_32076,N_32120);
nand U32376 (N_32376,N_32192,N_32005);
or U32377 (N_32377,N_32014,N_32174);
xor U32378 (N_32378,N_32136,N_32162);
nand U32379 (N_32379,N_32042,N_32219);
nand U32380 (N_32380,N_32236,N_32208);
xor U32381 (N_32381,N_32191,N_32174);
and U32382 (N_32382,N_32038,N_32110);
or U32383 (N_32383,N_32024,N_32183);
nor U32384 (N_32384,N_32193,N_32190);
nand U32385 (N_32385,N_32233,N_32045);
nor U32386 (N_32386,N_32137,N_32052);
nand U32387 (N_32387,N_32007,N_32028);
or U32388 (N_32388,N_32168,N_32077);
nor U32389 (N_32389,N_32047,N_32224);
nand U32390 (N_32390,N_32090,N_32209);
nor U32391 (N_32391,N_32247,N_32178);
or U32392 (N_32392,N_32081,N_32057);
nand U32393 (N_32393,N_32248,N_32218);
nand U32394 (N_32394,N_32192,N_32162);
or U32395 (N_32395,N_32182,N_32214);
or U32396 (N_32396,N_32185,N_32123);
xor U32397 (N_32397,N_32161,N_32117);
nor U32398 (N_32398,N_32114,N_32081);
xnor U32399 (N_32399,N_32136,N_32173);
or U32400 (N_32400,N_32238,N_32152);
nand U32401 (N_32401,N_32040,N_32072);
or U32402 (N_32402,N_32110,N_32123);
nand U32403 (N_32403,N_32248,N_32089);
nor U32404 (N_32404,N_32012,N_32050);
and U32405 (N_32405,N_32201,N_32070);
xor U32406 (N_32406,N_32076,N_32026);
or U32407 (N_32407,N_32025,N_32132);
nand U32408 (N_32408,N_32068,N_32196);
or U32409 (N_32409,N_32234,N_32115);
nand U32410 (N_32410,N_32019,N_32055);
or U32411 (N_32411,N_32233,N_32199);
nor U32412 (N_32412,N_32099,N_32176);
or U32413 (N_32413,N_32139,N_32204);
and U32414 (N_32414,N_32245,N_32084);
xnor U32415 (N_32415,N_32179,N_32033);
nor U32416 (N_32416,N_32155,N_32232);
nor U32417 (N_32417,N_32153,N_32065);
and U32418 (N_32418,N_32100,N_32043);
nor U32419 (N_32419,N_32234,N_32067);
and U32420 (N_32420,N_32115,N_32113);
nor U32421 (N_32421,N_32231,N_32098);
nor U32422 (N_32422,N_32121,N_32025);
and U32423 (N_32423,N_32161,N_32236);
nor U32424 (N_32424,N_32238,N_32045);
xnor U32425 (N_32425,N_32189,N_32208);
nor U32426 (N_32426,N_32014,N_32119);
or U32427 (N_32427,N_32010,N_32061);
nand U32428 (N_32428,N_32148,N_32020);
nor U32429 (N_32429,N_32182,N_32069);
nand U32430 (N_32430,N_32176,N_32245);
nand U32431 (N_32431,N_32002,N_32101);
or U32432 (N_32432,N_32015,N_32044);
xnor U32433 (N_32433,N_32234,N_32038);
or U32434 (N_32434,N_32089,N_32176);
nand U32435 (N_32435,N_32160,N_32061);
nand U32436 (N_32436,N_32182,N_32107);
xor U32437 (N_32437,N_32059,N_32142);
and U32438 (N_32438,N_32063,N_32058);
or U32439 (N_32439,N_32030,N_32039);
nor U32440 (N_32440,N_32130,N_32133);
and U32441 (N_32441,N_32174,N_32140);
or U32442 (N_32442,N_32064,N_32142);
or U32443 (N_32443,N_32054,N_32033);
nand U32444 (N_32444,N_32052,N_32235);
and U32445 (N_32445,N_32105,N_32094);
nand U32446 (N_32446,N_32240,N_32067);
or U32447 (N_32447,N_32211,N_32249);
and U32448 (N_32448,N_32171,N_32141);
and U32449 (N_32449,N_32186,N_32002);
nand U32450 (N_32450,N_32037,N_32188);
or U32451 (N_32451,N_32225,N_32122);
nor U32452 (N_32452,N_32048,N_32062);
or U32453 (N_32453,N_32204,N_32225);
nand U32454 (N_32454,N_32080,N_32158);
nor U32455 (N_32455,N_32240,N_32087);
nor U32456 (N_32456,N_32000,N_32193);
or U32457 (N_32457,N_32065,N_32062);
and U32458 (N_32458,N_32217,N_32011);
nand U32459 (N_32459,N_32223,N_32167);
xor U32460 (N_32460,N_32097,N_32238);
and U32461 (N_32461,N_32240,N_32202);
and U32462 (N_32462,N_32142,N_32046);
nor U32463 (N_32463,N_32042,N_32240);
nand U32464 (N_32464,N_32064,N_32174);
nand U32465 (N_32465,N_32217,N_32221);
and U32466 (N_32466,N_32010,N_32238);
and U32467 (N_32467,N_32068,N_32225);
nor U32468 (N_32468,N_32221,N_32053);
and U32469 (N_32469,N_32017,N_32238);
xor U32470 (N_32470,N_32158,N_32027);
nor U32471 (N_32471,N_32166,N_32045);
or U32472 (N_32472,N_32111,N_32240);
nor U32473 (N_32473,N_32018,N_32240);
or U32474 (N_32474,N_32065,N_32030);
xnor U32475 (N_32475,N_32146,N_32054);
or U32476 (N_32476,N_32097,N_32202);
and U32477 (N_32477,N_32202,N_32123);
nor U32478 (N_32478,N_32152,N_32076);
or U32479 (N_32479,N_32182,N_32225);
nand U32480 (N_32480,N_32239,N_32055);
and U32481 (N_32481,N_32239,N_32195);
and U32482 (N_32482,N_32113,N_32085);
and U32483 (N_32483,N_32146,N_32098);
and U32484 (N_32484,N_32236,N_32186);
nand U32485 (N_32485,N_32075,N_32194);
xor U32486 (N_32486,N_32184,N_32003);
and U32487 (N_32487,N_32062,N_32013);
xnor U32488 (N_32488,N_32108,N_32101);
and U32489 (N_32489,N_32174,N_32221);
xor U32490 (N_32490,N_32241,N_32147);
and U32491 (N_32491,N_32015,N_32223);
nor U32492 (N_32492,N_32026,N_32042);
nor U32493 (N_32493,N_32026,N_32166);
xnor U32494 (N_32494,N_32002,N_32134);
xnor U32495 (N_32495,N_32151,N_32075);
nor U32496 (N_32496,N_32157,N_32223);
and U32497 (N_32497,N_32152,N_32088);
xor U32498 (N_32498,N_32056,N_32130);
nand U32499 (N_32499,N_32062,N_32122);
and U32500 (N_32500,N_32261,N_32339);
or U32501 (N_32501,N_32359,N_32372);
nand U32502 (N_32502,N_32462,N_32376);
nand U32503 (N_32503,N_32387,N_32268);
or U32504 (N_32504,N_32408,N_32377);
nor U32505 (N_32505,N_32320,N_32271);
nor U32506 (N_32506,N_32390,N_32357);
xor U32507 (N_32507,N_32471,N_32447);
nor U32508 (N_32508,N_32440,N_32498);
and U32509 (N_32509,N_32319,N_32276);
xnor U32510 (N_32510,N_32267,N_32413);
nor U32511 (N_32511,N_32383,N_32250);
nand U32512 (N_32512,N_32433,N_32285);
xnor U32513 (N_32513,N_32441,N_32449);
or U32514 (N_32514,N_32463,N_32481);
nor U32515 (N_32515,N_32448,N_32489);
or U32516 (N_32516,N_32274,N_32355);
nand U32517 (N_32517,N_32352,N_32416);
nand U32518 (N_32518,N_32254,N_32337);
nor U32519 (N_32519,N_32304,N_32461);
and U32520 (N_32520,N_32289,N_32346);
nor U32521 (N_32521,N_32443,N_32403);
xor U32522 (N_32522,N_32412,N_32343);
nor U32523 (N_32523,N_32453,N_32389);
nor U32524 (N_32524,N_32392,N_32340);
or U32525 (N_32525,N_32353,N_32341);
nand U32526 (N_32526,N_32253,N_32306);
and U32527 (N_32527,N_32480,N_32310);
and U32528 (N_32528,N_32264,N_32493);
and U32529 (N_32529,N_32325,N_32410);
nand U32530 (N_32530,N_32458,N_32332);
and U32531 (N_32531,N_32475,N_32259);
xnor U32532 (N_32532,N_32331,N_32428);
nor U32533 (N_32533,N_32445,N_32257);
nand U32534 (N_32534,N_32361,N_32314);
xnor U32535 (N_32535,N_32280,N_32400);
or U32536 (N_32536,N_32496,N_32405);
or U32537 (N_32537,N_32411,N_32299);
or U32538 (N_32538,N_32328,N_32307);
xnor U32539 (N_32539,N_32270,N_32393);
or U32540 (N_32540,N_32497,N_32479);
nor U32541 (N_32541,N_32386,N_32266);
and U32542 (N_32542,N_32363,N_32450);
nor U32543 (N_32543,N_32351,N_32309);
xnor U32544 (N_32544,N_32371,N_32382);
and U32545 (N_32545,N_32296,N_32315);
nor U32546 (N_32546,N_32301,N_32467);
or U32547 (N_32547,N_32385,N_32338);
or U32548 (N_32548,N_32415,N_32330);
and U32549 (N_32549,N_32273,N_32362);
nand U32550 (N_32550,N_32396,N_32406);
nand U32551 (N_32551,N_32476,N_32483);
nor U32552 (N_32552,N_32348,N_32425);
and U32553 (N_32553,N_32401,N_32278);
or U32554 (N_32554,N_32418,N_32350);
nor U32555 (N_32555,N_32398,N_32367);
and U32556 (N_32556,N_32327,N_32432);
nand U32557 (N_32557,N_32437,N_32399);
and U32558 (N_32558,N_32300,N_32251);
xor U32559 (N_32559,N_32308,N_32446);
and U32560 (N_32560,N_32414,N_32313);
and U32561 (N_32561,N_32265,N_32349);
nor U32562 (N_32562,N_32460,N_32459);
nand U32563 (N_32563,N_32404,N_32286);
and U32564 (N_32564,N_32358,N_32435);
nand U32565 (N_32565,N_32488,N_32336);
nand U32566 (N_32566,N_32391,N_32490);
xnor U32567 (N_32567,N_32395,N_32269);
nor U32568 (N_32568,N_32487,N_32292);
xor U32569 (N_32569,N_32262,N_32409);
nand U32570 (N_32570,N_32454,N_32263);
and U32571 (N_32571,N_32255,N_32482);
nand U32572 (N_32572,N_32347,N_32438);
or U32573 (N_32573,N_32378,N_32284);
nand U32574 (N_32574,N_32303,N_32470);
nor U32575 (N_32575,N_32258,N_32423);
and U32576 (N_32576,N_32485,N_32431);
xor U32577 (N_32577,N_32442,N_32466);
xnor U32578 (N_32578,N_32464,N_32334);
xnor U32579 (N_32579,N_32290,N_32429);
and U32580 (N_32580,N_32370,N_32472);
or U32581 (N_32581,N_32426,N_32495);
xnor U32582 (N_32582,N_32397,N_32275);
and U32583 (N_32583,N_32407,N_32288);
and U32584 (N_32584,N_32282,N_32379);
nor U32585 (N_32585,N_32468,N_32486);
nor U32586 (N_32586,N_32388,N_32298);
nand U32587 (N_32587,N_32434,N_32421);
nor U32588 (N_32588,N_32333,N_32455);
xor U32589 (N_32589,N_32342,N_32294);
xor U32590 (N_32590,N_32439,N_32402);
nand U32591 (N_32591,N_32305,N_32424);
or U32592 (N_32592,N_32324,N_32365);
and U32593 (N_32593,N_32364,N_32469);
and U32594 (N_32594,N_32419,N_32491);
nand U32595 (N_32595,N_32316,N_32473);
or U32596 (N_32596,N_32368,N_32302);
xnor U32597 (N_32597,N_32456,N_32272);
xor U32598 (N_32598,N_32394,N_32318);
and U32599 (N_32599,N_32279,N_32317);
nand U32600 (N_32600,N_32451,N_32277);
nor U32601 (N_32601,N_32384,N_32452);
nor U32602 (N_32602,N_32256,N_32322);
or U32603 (N_32603,N_32457,N_32260);
nor U32604 (N_32604,N_32380,N_32474);
and U32605 (N_32605,N_32356,N_32492);
xnor U32606 (N_32606,N_32373,N_32297);
nor U32607 (N_32607,N_32354,N_32252);
xnor U32608 (N_32608,N_32311,N_32281);
xnor U32609 (N_32609,N_32369,N_32427);
xor U32610 (N_32610,N_32335,N_32326);
nand U32611 (N_32611,N_32420,N_32312);
or U32612 (N_32612,N_32375,N_32494);
and U32613 (N_32613,N_32381,N_32422);
xnor U32614 (N_32614,N_32323,N_32484);
or U32615 (N_32615,N_32436,N_32329);
or U32616 (N_32616,N_32430,N_32366);
nor U32617 (N_32617,N_32465,N_32295);
nor U32618 (N_32618,N_32477,N_32360);
nor U32619 (N_32619,N_32283,N_32287);
and U32620 (N_32620,N_32321,N_32293);
and U32621 (N_32621,N_32444,N_32417);
or U32622 (N_32622,N_32374,N_32478);
xor U32623 (N_32623,N_32499,N_32344);
nand U32624 (N_32624,N_32345,N_32291);
and U32625 (N_32625,N_32382,N_32428);
xnor U32626 (N_32626,N_32482,N_32374);
or U32627 (N_32627,N_32454,N_32464);
nand U32628 (N_32628,N_32387,N_32254);
nor U32629 (N_32629,N_32498,N_32358);
xor U32630 (N_32630,N_32259,N_32341);
nand U32631 (N_32631,N_32407,N_32419);
xnor U32632 (N_32632,N_32346,N_32424);
nand U32633 (N_32633,N_32441,N_32421);
and U32634 (N_32634,N_32257,N_32389);
xor U32635 (N_32635,N_32422,N_32425);
nor U32636 (N_32636,N_32322,N_32465);
nand U32637 (N_32637,N_32263,N_32316);
nor U32638 (N_32638,N_32481,N_32483);
nand U32639 (N_32639,N_32428,N_32358);
and U32640 (N_32640,N_32347,N_32260);
and U32641 (N_32641,N_32321,N_32271);
and U32642 (N_32642,N_32377,N_32342);
nor U32643 (N_32643,N_32399,N_32278);
or U32644 (N_32644,N_32477,N_32301);
nor U32645 (N_32645,N_32453,N_32498);
nor U32646 (N_32646,N_32260,N_32497);
xor U32647 (N_32647,N_32451,N_32446);
xnor U32648 (N_32648,N_32347,N_32358);
nand U32649 (N_32649,N_32432,N_32424);
nand U32650 (N_32650,N_32356,N_32259);
nand U32651 (N_32651,N_32406,N_32424);
or U32652 (N_32652,N_32361,N_32383);
nor U32653 (N_32653,N_32330,N_32310);
nor U32654 (N_32654,N_32391,N_32298);
or U32655 (N_32655,N_32461,N_32472);
nor U32656 (N_32656,N_32260,N_32375);
and U32657 (N_32657,N_32287,N_32348);
and U32658 (N_32658,N_32258,N_32371);
nor U32659 (N_32659,N_32469,N_32350);
nand U32660 (N_32660,N_32341,N_32456);
or U32661 (N_32661,N_32453,N_32406);
nand U32662 (N_32662,N_32299,N_32466);
or U32663 (N_32663,N_32391,N_32259);
xor U32664 (N_32664,N_32309,N_32334);
nand U32665 (N_32665,N_32477,N_32374);
and U32666 (N_32666,N_32374,N_32368);
or U32667 (N_32667,N_32324,N_32309);
or U32668 (N_32668,N_32444,N_32335);
nand U32669 (N_32669,N_32451,N_32312);
or U32670 (N_32670,N_32489,N_32366);
or U32671 (N_32671,N_32448,N_32326);
and U32672 (N_32672,N_32260,N_32431);
nor U32673 (N_32673,N_32393,N_32254);
nor U32674 (N_32674,N_32420,N_32351);
xor U32675 (N_32675,N_32275,N_32478);
xnor U32676 (N_32676,N_32326,N_32435);
nand U32677 (N_32677,N_32393,N_32427);
xnor U32678 (N_32678,N_32467,N_32323);
and U32679 (N_32679,N_32255,N_32363);
and U32680 (N_32680,N_32458,N_32268);
or U32681 (N_32681,N_32325,N_32402);
or U32682 (N_32682,N_32303,N_32337);
and U32683 (N_32683,N_32454,N_32344);
nand U32684 (N_32684,N_32284,N_32257);
xnor U32685 (N_32685,N_32404,N_32269);
nand U32686 (N_32686,N_32305,N_32288);
or U32687 (N_32687,N_32363,N_32299);
nand U32688 (N_32688,N_32466,N_32377);
xor U32689 (N_32689,N_32382,N_32253);
or U32690 (N_32690,N_32325,N_32446);
and U32691 (N_32691,N_32460,N_32413);
or U32692 (N_32692,N_32358,N_32287);
xor U32693 (N_32693,N_32412,N_32295);
and U32694 (N_32694,N_32313,N_32321);
and U32695 (N_32695,N_32342,N_32284);
and U32696 (N_32696,N_32287,N_32301);
xnor U32697 (N_32697,N_32427,N_32259);
or U32698 (N_32698,N_32275,N_32458);
xnor U32699 (N_32699,N_32328,N_32400);
nor U32700 (N_32700,N_32431,N_32310);
nor U32701 (N_32701,N_32350,N_32343);
xnor U32702 (N_32702,N_32280,N_32318);
nor U32703 (N_32703,N_32308,N_32344);
and U32704 (N_32704,N_32459,N_32383);
xor U32705 (N_32705,N_32301,N_32375);
nand U32706 (N_32706,N_32371,N_32429);
or U32707 (N_32707,N_32280,N_32441);
or U32708 (N_32708,N_32430,N_32344);
xor U32709 (N_32709,N_32253,N_32261);
nor U32710 (N_32710,N_32453,N_32495);
nor U32711 (N_32711,N_32420,N_32334);
and U32712 (N_32712,N_32326,N_32365);
xnor U32713 (N_32713,N_32454,N_32449);
and U32714 (N_32714,N_32304,N_32390);
xor U32715 (N_32715,N_32407,N_32281);
nor U32716 (N_32716,N_32400,N_32257);
nor U32717 (N_32717,N_32402,N_32405);
or U32718 (N_32718,N_32257,N_32278);
nor U32719 (N_32719,N_32355,N_32292);
and U32720 (N_32720,N_32253,N_32344);
xor U32721 (N_32721,N_32447,N_32496);
nor U32722 (N_32722,N_32384,N_32376);
or U32723 (N_32723,N_32257,N_32408);
xnor U32724 (N_32724,N_32258,N_32406);
or U32725 (N_32725,N_32435,N_32476);
nand U32726 (N_32726,N_32361,N_32295);
nor U32727 (N_32727,N_32410,N_32270);
and U32728 (N_32728,N_32327,N_32421);
or U32729 (N_32729,N_32304,N_32404);
nor U32730 (N_32730,N_32478,N_32388);
nand U32731 (N_32731,N_32262,N_32270);
xor U32732 (N_32732,N_32403,N_32337);
nor U32733 (N_32733,N_32271,N_32446);
and U32734 (N_32734,N_32268,N_32321);
xnor U32735 (N_32735,N_32460,N_32252);
xor U32736 (N_32736,N_32439,N_32396);
nand U32737 (N_32737,N_32303,N_32440);
or U32738 (N_32738,N_32476,N_32376);
nand U32739 (N_32739,N_32411,N_32489);
and U32740 (N_32740,N_32323,N_32266);
nor U32741 (N_32741,N_32478,N_32460);
or U32742 (N_32742,N_32272,N_32489);
xor U32743 (N_32743,N_32276,N_32418);
nand U32744 (N_32744,N_32297,N_32262);
and U32745 (N_32745,N_32415,N_32278);
and U32746 (N_32746,N_32411,N_32485);
nand U32747 (N_32747,N_32464,N_32322);
or U32748 (N_32748,N_32391,N_32460);
nor U32749 (N_32749,N_32498,N_32352);
and U32750 (N_32750,N_32619,N_32627);
and U32751 (N_32751,N_32719,N_32628);
or U32752 (N_32752,N_32660,N_32596);
nor U32753 (N_32753,N_32698,N_32583);
nor U32754 (N_32754,N_32564,N_32650);
nand U32755 (N_32755,N_32533,N_32507);
nand U32756 (N_32756,N_32707,N_32638);
xor U32757 (N_32757,N_32633,N_32555);
and U32758 (N_32758,N_32557,N_32662);
nand U32759 (N_32759,N_32513,N_32609);
or U32760 (N_32760,N_32712,N_32735);
nor U32761 (N_32761,N_32641,N_32611);
and U32762 (N_32762,N_32673,N_32636);
xnor U32763 (N_32763,N_32672,N_32692);
or U32764 (N_32764,N_32706,N_32710);
nor U32765 (N_32765,N_32670,N_32589);
xnor U32766 (N_32766,N_32543,N_32567);
nand U32767 (N_32767,N_32695,N_32541);
xnor U32768 (N_32768,N_32529,N_32518);
xnor U32769 (N_32769,N_32514,N_32547);
xor U32770 (N_32770,N_32632,N_32648);
and U32771 (N_32771,N_32720,N_32747);
nor U32772 (N_32772,N_32665,N_32681);
and U32773 (N_32773,N_32524,N_32744);
or U32774 (N_32774,N_32510,N_32739);
xnor U32775 (N_32775,N_32709,N_32714);
nand U32776 (N_32776,N_32553,N_32540);
nor U32777 (N_32777,N_32661,N_32624);
xor U32778 (N_32778,N_32642,N_32565);
nand U32779 (N_32779,N_32504,N_32597);
or U32780 (N_32780,N_32689,N_32519);
nand U32781 (N_32781,N_32625,N_32502);
and U32782 (N_32782,N_32595,N_32621);
xnor U32783 (N_32783,N_32604,N_32708);
nor U32784 (N_32784,N_32570,N_32738);
nor U32785 (N_32785,N_32727,N_32729);
and U32786 (N_32786,N_32560,N_32556);
nor U32787 (N_32787,N_32591,N_32525);
or U32788 (N_32788,N_32684,N_32615);
xor U32789 (N_32789,N_32749,N_32563);
and U32790 (N_32790,N_32551,N_32520);
and U32791 (N_32791,N_32705,N_32617);
or U32792 (N_32792,N_32581,N_32594);
xnor U32793 (N_32793,N_32618,N_32580);
nor U32794 (N_32794,N_32506,N_32701);
nor U32795 (N_32795,N_32603,N_32616);
xnor U32796 (N_32796,N_32716,N_32649);
nand U32797 (N_32797,N_32511,N_32571);
nand U32798 (N_32798,N_32503,N_32659);
and U32799 (N_32799,N_32626,N_32667);
nor U32800 (N_32800,N_32577,N_32645);
xnor U32801 (N_32801,N_32653,N_32568);
nor U32802 (N_32802,N_32635,N_32606);
and U32803 (N_32803,N_32538,N_32713);
nor U32804 (N_32804,N_32679,N_32535);
nor U32805 (N_32805,N_32654,N_32607);
nand U32806 (N_32806,N_32732,N_32702);
nand U32807 (N_32807,N_32746,N_32512);
or U32808 (N_32808,N_32505,N_32664);
nand U32809 (N_32809,N_32523,N_32687);
and U32810 (N_32810,N_32558,N_32554);
xor U32811 (N_32811,N_32620,N_32742);
or U32812 (N_32812,N_32640,N_32584);
or U32813 (N_32813,N_32522,N_32723);
xnor U32814 (N_32814,N_32601,N_32587);
and U32815 (N_32815,N_32599,N_32715);
and U32816 (N_32816,N_32509,N_32526);
xnor U32817 (N_32817,N_32657,N_32717);
and U32818 (N_32818,N_32500,N_32630);
or U32819 (N_32819,N_32697,N_32721);
and U32820 (N_32820,N_32734,N_32546);
nor U32821 (N_32821,N_32562,N_32652);
and U32822 (N_32822,N_32532,N_32600);
or U32823 (N_32823,N_32559,N_32743);
nor U32824 (N_32824,N_32578,N_32688);
or U32825 (N_32825,N_32639,N_32588);
or U32826 (N_32826,N_32544,N_32646);
or U32827 (N_32827,N_32737,N_32542);
or U32828 (N_32828,N_32521,N_32605);
nor U32829 (N_32829,N_32671,N_32678);
nor U32830 (N_32830,N_32548,N_32573);
nor U32831 (N_32831,N_32592,N_32655);
or U32832 (N_32832,N_32730,N_32682);
nor U32833 (N_32833,N_32722,N_32608);
xnor U32834 (N_32834,N_32602,N_32574);
and U32835 (N_32835,N_32718,N_32598);
or U32836 (N_32836,N_32725,N_32516);
nor U32837 (N_32837,N_32666,N_32585);
or U32838 (N_32838,N_32728,N_32731);
xor U32839 (N_32839,N_32508,N_32663);
xnor U32840 (N_32840,N_32569,N_32593);
nor U32841 (N_32841,N_32685,N_32647);
nor U32842 (N_32842,N_32623,N_32700);
nor U32843 (N_32843,N_32745,N_32552);
or U32844 (N_32844,N_32528,N_32634);
xor U32845 (N_32845,N_32531,N_32579);
or U32846 (N_32846,N_32515,N_32545);
nor U32847 (N_32847,N_32674,N_32656);
nor U32848 (N_32848,N_32686,N_32699);
xor U32849 (N_32849,N_32582,N_32675);
nand U32850 (N_32850,N_32677,N_32680);
or U32851 (N_32851,N_32612,N_32631);
xnor U32852 (N_32852,N_32703,N_32586);
and U32853 (N_32853,N_32530,N_32566);
or U32854 (N_32854,N_32614,N_32740);
or U32855 (N_32855,N_32724,N_32549);
xor U32856 (N_32856,N_32683,N_32610);
nor U32857 (N_32857,N_32539,N_32733);
nor U32858 (N_32858,N_32643,N_32613);
nand U32859 (N_32859,N_32590,N_32676);
xnor U32860 (N_32860,N_32576,N_32572);
xnor U32861 (N_32861,N_32694,N_32501);
xor U32862 (N_32862,N_32726,N_32622);
xnor U32863 (N_32863,N_32669,N_32748);
xor U32864 (N_32864,N_32629,N_32534);
nor U32865 (N_32865,N_32690,N_32644);
and U32866 (N_32866,N_32668,N_32711);
xnor U32867 (N_32867,N_32736,N_32537);
nor U32868 (N_32868,N_32696,N_32691);
nand U32869 (N_32869,N_32575,N_32550);
nor U32870 (N_32870,N_32704,N_32536);
and U32871 (N_32871,N_32527,N_32658);
nand U32872 (N_32872,N_32637,N_32693);
nand U32873 (N_32873,N_32651,N_32561);
nor U32874 (N_32874,N_32741,N_32517);
and U32875 (N_32875,N_32643,N_32682);
and U32876 (N_32876,N_32699,N_32647);
and U32877 (N_32877,N_32605,N_32591);
and U32878 (N_32878,N_32629,N_32631);
and U32879 (N_32879,N_32671,N_32689);
nor U32880 (N_32880,N_32502,N_32603);
xnor U32881 (N_32881,N_32651,N_32684);
nand U32882 (N_32882,N_32575,N_32513);
nor U32883 (N_32883,N_32540,N_32708);
nor U32884 (N_32884,N_32520,N_32667);
nor U32885 (N_32885,N_32622,N_32556);
xnor U32886 (N_32886,N_32515,N_32668);
or U32887 (N_32887,N_32580,N_32554);
xnor U32888 (N_32888,N_32542,N_32693);
nand U32889 (N_32889,N_32676,N_32541);
nand U32890 (N_32890,N_32657,N_32663);
xor U32891 (N_32891,N_32534,N_32690);
nand U32892 (N_32892,N_32678,N_32657);
xor U32893 (N_32893,N_32544,N_32627);
and U32894 (N_32894,N_32611,N_32633);
or U32895 (N_32895,N_32534,N_32621);
or U32896 (N_32896,N_32713,N_32501);
nor U32897 (N_32897,N_32544,N_32733);
xor U32898 (N_32898,N_32742,N_32618);
nand U32899 (N_32899,N_32704,N_32719);
nand U32900 (N_32900,N_32710,N_32557);
nand U32901 (N_32901,N_32670,N_32686);
nand U32902 (N_32902,N_32564,N_32691);
or U32903 (N_32903,N_32547,N_32541);
xnor U32904 (N_32904,N_32630,N_32736);
nand U32905 (N_32905,N_32527,N_32533);
nor U32906 (N_32906,N_32660,N_32574);
nor U32907 (N_32907,N_32586,N_32644);
or U32908 (N_32908,N_32602,N_32592);
nand U32909 (N_32909,N_32622,N_32723);
or U32910 (N_32910,N_32627,N_32514);
nand U32911 (N_32911,N_32651,N_32722);
xor U32912 (N_32912,N_32748,N_32567);
nand U32913 (N_32913,N_32547,N_32562);
or U32914 (N_32914,N_32627,N_32748);
or U32915 (N_32915,N_32705,N_32557);
or U32916 (N_32916,N_32607,N_32524);
or U32917 (N_32917,N_32507,N_32689);
or U32918 (N_32918,N_32521,N_32514);
xnor U32919 (N_32919,N_32592,N_32677);
nor U32920 (N_32920,N_32706,N_32504);
or U32921 (N_32921,N_32694,N_32728);
nor U32922 (N_32922,N_32583,N_32620);
nor U32923 (N_32923,N_32741,N_32726);
xnor U32924 (N_32924,N_32726,N_32574);
and U32925 (N_32925,N_32687,N_32509);
nor U32926 (N_32926,N_32702,N_32743);
xnor U32927 (N_32927,N_32696,N_32543);
xor U32928 (N_32928,N_32519,N_32723);
and U32929 (N_32929,N_32614,N_32580);
nand U32930 (N_32930,N_32685,N_32614);
and U32931 (N_32931,N_32595,N_32732);
xnor U32932 (N_32932,N_32634,N_32567);
nor U32933 (N_32933,N_32728,N_32542);
or U32934 (N_32934,N_32671,N_32623);
nor U32935 (N_32935,N_32555,N_32529);
and U32936 (N_32936,N_32626,N_32507);
and U32937 (N_32937,N_32741,N_32572);
xnor U32938 (N_32938,N_32504,N_32694);
and U32939 (N_32939,N_32622,N_32695);
nor U32940 (N_32940,N_32638,N_32591);
nor U32941 (N_32941,N_32563,N_32658);
or U32942 (N_32942,N_32689,N_32570);
xnor U32943 (N_32943,N_32558,N_32649);
xor U32944 (N_32944,N_32660,N_32580);
xor U32945 (N_32945,N_32688,N_32559);
or U32946 (N_32946,N_32721,N_32690);
xnor U32947 (N_32947,N_32578,N_32599);
nor U32948 (N_32948,N_32743,N_32601);
xnor U32949 (N_32949,N_32681,N_32536);
or U32950 (N_32950,N_32519,N_32518);
or U32951 (N_32951,N_32677,N_32707);
nor U32952 (N_32952,N_32668,N_32578);
nor U32953 (N_32953,N_32639,N_32630);
nor U32954 (N_32954,N_32662,N_32565);
nor U32955 (N_32955,N_32576,N_32738);
or U32956 (N_32956,N_32671,N_32747);
nor U32957 (N_32957,N_32515,N_32656);
and U32958 (N_32958,N_32684,N_32623);
and U32959 (N_32959,N_32717,N_32622);
nand U32960 (N_32960,N_32566,N_32684);
nand U32961 (N_32961,N_32549,N_32690);
or U32962 (N_32962,N_32612,N_32683);
nand U32963 (N_32963,N_32723,N_32516);
and U32964 (N_32964,N_32601,N_32507);
nand U32965 (N_32965,N_32547,N_32667);
nand U32966 (N_32966,N_32621,N_32536);
and U32967 (N_32967,N_32516,N_32749);
nor U32968 (N_32968,N_32715,N_32702);
and U32969 (N_32969,N_32554,N_32736);
nor U32970 (N_32970,N_32735,N_32657);
and U32971 (N_32971,N_32735,N_32683);
or U32972 (N_32972,N_32501,N_32512);
and U32973 (N_32973,N_32703,N_32692);
and U32974 (N_32974,N_32622,N_32517);
xnor U32975 (N_32975,N_32586,N_32519);
nor U32976 (N_32976,N_32618,N_32626);
nand U32977 (N_32977,N_32722,N_32692);
xor U32978 (N_32978,N_32736,N_32745);
or U32979 (N_32979,N_32680,N_32576);
xnor U32980 (N_32980,N_32555,N_32660);
nor U32981 (N_32981,N_32745,N_32528);
or U32982 (N_32982,N_32667,N_32540);
nor U32983 (N_32983,N_32568,N_32577);
nand U32984 (N_32984,N_32533,N_32525);
xnor U32985 (N_32985,N_32670,N_32596);
and U32986 (N_32986,N_32708,N_32672);
and U32987 (N_32987,N_32711,N_32667);
xor U32988 (N_32988,N_32671,N_32691);
and U32989 (N_32989,N_32609,N_32603);
nand U32990 (N_32990,N_32609,N_32611);
nand U32991 (N_32991,N_32603,N_32635);
nand U32992 (N_32992,N_32696,N_32657);
and U32993 (N_32993,N_32599,N_32593);
xor U32994 (N_32994,N_32736,N_32602);
nand U32995 (N_32995,N_32715,N_32717);
nand U32996 (N_32996,N_32543,N_32555);
nor U32997 (N_32997,N_32628,N_32583);
or U32998 (N_32998,N_32588,N_32742);
and U32999 (N_32999,N_32710,N_32567);
nor U33000 (N_33000,N_32947,N_32794);
nand U33001 (N_33001,N_32764,N_32894);
xor U33002 (N_33002,N_32851,N_32801);
nor U33003 (N_33003,N_32855,N_32774);
and U33004 (N_33004,N_32974,N_32782);
nand U33005 (N_33005,N_32937,N_32762);
and U33006 (N_33006,N_32791,N_32816);
and U33007 (N_33007,N_32799,N_32893);
or U33008 (N_33008,N_32999,N_32953);
nor U33009 (N_33009,N_32991,N_32892);
xnor U33010 (N_33010,N_32758,N_32926);
or U33011 (N_33011,N_32772,N_32853);
nor U33012 (N_33012,N_32865,N_32787);
nor U33013 (N_33013,N_32860,N_32882);
nor U33014 (N_33014,N_32757,N_32863);
nor U33015 (N_33015,N_32760,N_32890);
or U33016 (N_33016,N_32839,N_32888);
nand U33017 (N_33017,N_32846,N_32884);
or U33018 (N_33018,N_32763,N_32939);
nand U33019 (N_33019,N_32809,N_32807);
nor U33020 (N_33020,N_32908,N_32810);
nor U33021 (N_33021,N_32792,N_32910);
xor U33022 (N_33022,N_32815,N_32964);
nand U33023 (N_33023,N_32978,N_32907);
nand U33024 (N_33024,N_32990,N_32979);
nor U33025 (N_33025,N_32814,N_32784);
xnor U33026 (N_33026,N_32837,N_32822);
nor U33027 (N_33027,N_32820,N_32903);
or U33028 (N_33028,N_32891,N_32971);
nand U33029 (N_33029,N_32995,N_32955);
and U33030 (N_33030,N_32766,N_32925);
and U33031 (N_33031,N_32959,N_32924);
and U33032 (N_33032,N_32927,N_32994);
or U33033 (N_33033,N_32871,N_32946);
and U33034 (N_33034,N_32818,N_32840);
xnor U33035 (N_33035,N_32933,N_32821);
nor U33036 (N_33036,N_32988,N_32786);
xnor U33037 (N_33037,N_32962,N_32977);
nor U33038 (N_33038,N_32886,N_32843);
nand U33039 (N_33039,N_32832,N_32864);
xor U33040 (N_33040,N_32836,N_32795);
nand U33041 (N_33041,N_32875,N_32844);
or U33042 (N_33042,N_32852,N_32993);
nand U33043 (N_33043,N_32986,N_32773);
or U33044 (N_33044,N_32916,N_32896);
or U33045 (N_33045,N_32826,N_32847);
nor U33046 (N_33046,N_32948,N_32951);
and U33047 (N_33047,N_32835,N_32841);
nor U33048 (N_33048,N_32788,N_32833);
and U33049 (N_33049,N_32917,N_32883);
nor U33050 (N_33050,N_32845,N_32831);
nand U33051 (N_33051,N_32755,N_32957);
nor U33052 (N_33052,N_32857,N_32872);
and U33053 (N_33053,N_32806,N_32797);
or U33054 (N_33054,N_32877,N_32779);
and U33055 (N_33055,N_32906,N_32811);
and U33056 (N_33056,N_32767,N_32935);
and U33057 (N_33057,N_32854,N_32889);
or U33058 (N_33058,N_32929,N_32873);
nor U33059 (N_33059,N_32751,N_32842);
and U33060 (N_33060,N_32998,N_32928);
or U33061 (N_33061,N_32954,N_32895);
and U33062 (N_33062,N_32973,N_32808);
or U33063 (N_33063,N_32769,N_32879);
xnor U33064 (N_33064,N_32915,N_32753);
nor U33065 (N_33065,N_32966,N_32805);
xnor U33066 (N_33066,N_32777,N_32756);
nand U33067 (N_33067,N_32980,N_32931);
and U33068 (N_33068,N_32950,N_32898);
nor U33069 (N_33069,N_32752,N_32969);
nor U33070 (N_33070,N_32913,N_32970);
or U33071 (N_33071,N_32941,N_32942);
nand U33072 (N_33072,N_32904,N_32914);
nor U33073 (N_33073,N_32902,N_32824);
xor U33074 (N_33074,N_32900,N_32975);
nand U33075 (N_33075,N_32923,N_32934);
nor U33076 (N_33076,N_32936,N_32972);
nor U33077 (N_33077,N_32861,N_32823);
or U33078 (N_33078,N_32776,N_32858);
or U33079 (N_33079,N_32862,N_32930);
xor U33080 (N_33080,N_32850,N_32870);
or U33081 (N_33081,N_32905,N_32874);
and U33082 (N_33082,N_32897,N_32802);
xor U33083 (N_33083,N_32768,N_32921);
and U33084 (N_33084,N_32952,N_32868);
or U33085 (N_33085,N_32912,N_32922);
nand U33086 (N_33086,N_32789,N_32798);
and U33087 (N_33087,N_32825,N_32943);
and U33088 (N_33088,N_32830,N_32876);
nand U33089 (N_33089,N_32920,N_32911);
nor U33090 (N_33090,N_32958,N_32982);
nor U33091 (N_33091,N_32800,N_32765);
or U33092 (N_33092,N_32828,N_32867);
nand U33093 (N_33093,N_32849,N_32938);
nand U33094 (N_33094,N_32987,N_32940);
nand U33095 (N_33095,N_32856,N_32778);
xor U33096 (N_33096,N_32750,N_32785);
and U33097 (N_33097,N_32881,N_32793);
nor U33098 (N_33098,N_32848,N_32780);
nor U33099 (N_33099,N_32992,N_32869);
nand U33100 (N_33100,N_32996,N_32997);
nand U33101 (N_33101,N_32761,N_32866);
or U33102 (N_33102,N_32887,N_32960);
xnor U33103 (N_33103,N_32963,N_32984);
or U33104 (N_33104,N_32961,N_32919);
nor U33105 (N_33105,N_32918,N_32945);
and U33106 (N_33106,N_32949,N_32944);
xnor U33107 (N_33107,N_32956,N_32796);
nor U33108 (N_33108,N_32965,N_32968);
xnor U33109 (N_33109,N_32838,N_32976);
xor U33110 (N_33110,N_32859,N_32901);
and U33111 (N_33111,N_32909,N_32771);
or U33112 (N_33112,N_32770,N_32878);
nand U33113 (N_33113,N_32817,N_32812);
nor U33114 (N_33114,N_32827,N_32981);
nand U33115 (N_33115,N_32932,N_32781);
nor U33116 (N_33116,N_32880,N_32829);
or U33117 (N_33117,N_32989,N_32819);
nand U33118 (N_33118,N_32885,N_32790);
and U33119 (N_33119,N_32967,N_32813);
and U33120 (N_33120,N_32759,N_32834);
xor U33121 (N_33121,N_32775,N_32754);
and U33122 (N_33122,N_32803,N_32899);
and U33123 (N_33123,N_32804,N_32983);
nand U33124 (N_33124,N_32783,N_32985);
xor U33125 (N_33125,N_32780,N_32966);
xor U33126 (N_33126,N_32820,N_32834);
and U33127 (N_33127,N_32827,N_32799);
nor U33128 (N_33128,N_32996,N_32955);
or U33129 (N_33129,N_32949,N_32960);
nand U33130 (N_33130,N_32915,N_32855);
and U33131 (N_33131,N_32871,N_32933);
or U33132 (N_33132,N_32990,N_32834);
and U33133 (N_33133,N_32914,N_32759);
nor U33134 (N_33134,N_32770,N_32802);
nand U33135 (N_33135,N_32762,N_32848);
or U33136 (N_33136,N_32766,N_32866);
xor U33137 (N_33137,N_32892,N_32913);
nand U33138 (N_33138,N_32912,N_32816);
nand U33139 (N_33139,N_32772,N_32791);
xor U33140 (N_33140,N_32991,N_32923);
and U33141 (N_33141,N_32900,N_32862);
or U33142 (N_33142,N_32844,N_32821);
nand U33143 (N_33143,N_32895,N_32855);
nor U33144 (N_33144,N_32981,N_32898);
xor U33145 (N_33145,N_32856,N_32962);
nand U33146 (N_33146,N_32762,N_32947);
and U33147 (N_33147,N_32919,N_32783);
or U33148 (N_33148,N_32858,N_32924);
and U33149 (N_33149,N_32829,N_32870);
or U33150 (N_33150,N_32924,N_32985);
nand U33151 (N_33151,N_32877,N_32981);
nor U33152 (N_33152,N_32835,N_32946);
xor U33153 (N_33153,N_32804,N_32789);
xnor U33154 (N_33154,N_32833,N_32836);
or U33155 (N_33155,N_32962,N_32769);
xnor U33156 (N_33156,N_32794,N_32964);
nand U33157 (N_33157,N_32803,N_32942);
nor U33158 (N_33158,N_32869,N_32900);
xnor U33159 (N_33159,N_32783,N_32856);
nand U33160 (N_33160,N_32970,N_32781);
or U33161 (N_33161,N_32924,N_32931);
and U33162 (N_33162,N_32853,N_32983);
xor U33163 (N_33163,N_32840,N_32889);
or U33164 (N_33164,N_32868,N_32922);
nor U33165 (N_33165,N_32866,N_32804);
or U33166 (N_33166,N_32757,N_32777);
and U33167 (N_33167,N_32997,N_32773);
xor U33168 (N_33168,N_32858,N_32877);
nand U33169 (N_33169,N_32904,N_32991);
nor U33170 (N_33170,N_32869,N_32921);
or U33171 (N_33171,N_32784,N_32957);
or U33172 (N_33172,N_32921,N_32972);
xnor U33173 (N_33173,N_32807,N_32900);
xor U33174 (N_33174,N_32891,N_32866);
nor U33175 (N_33175,N_32847,N_32893);
xor U33176 (N_33176,N_32969,N_32793);
nand U33177 (N_33177,N_32824,N_32825);
nand U33178 (N_33178,N_32878,N_32774);
xor U33179 (N_33179,N_32803,N_32790);
nand U33180 (N_33180,N_32906,N_32872);
nand U33181 (N_33181,N_32928,N_32847);
or U33182 (N_33182,N_32989,N_32824);
xor U33183 (N_33183,N_32879,N_32905);
nand U33184 (N_33184,N_32891,N_32758);
nand U33185 (N_33185,N_32845,N_32889);
nand U33186 (N_33186,N_32872,N_32864);
nor U33187 (N_33187,N_32979,N_32977);
xor U33188 (N_33188,N_32881,N_32801);
and U33189 (N_33189,N_32791,N_32901);
xor U33190 (N_33190,N_32792,N_32823);
or U33191 (N_33191,N_32778,N_32773);
xnor U33192 (N_33192,N_32996,N_32777);
xor U33193 (N_33193,N_32765,N_32780);
nor U33194 (N_33194,N_32905,N_32930);
xor U33195 (N_33195,N_32835,N_32762);
xnor U33196 (N_33196,N_32923,N_32795);
nor U33197 (N_33197,N_32986,N_32994);
and U33198 (N_33198,N_32892,N_32860);
nand U33199 (N_33199,N_32875,N_32800);
xnor U33200 (N_33200,N_32882,N_32862);
nand U33201 (N_33201,N_32863,N_32974);
or U33202 (N_33202,N_32789,N_32808);
xor U33203 (N_33203,N_32853,N_32867);
nor U33204 (N_33204,N_32792,N_32923);
and U33205 (N_33205,N_32793,N_32855);
xnor U33206 (N_33206,N_32921,N_32848);
nand U33207 (N_33207,N_32911,N_32910);
nor U33208 (N_33208,N_32903,N_32950);
and U33209 (N_33209,N_32914,N_32786);
nor U33210 (N_33210,N_32985,N_32827);
xnor U33211 (N_33211,N_32870,N_32811);
nand U33212 (N_33212,N_32976,N_32963);
nor U33213 (N_33213,N_32762,N_32976);
nand U33214 (N_33214,N_32752,N_32894);
nor U33215 (N_33215,N_32949,N_32834);
xnor U33216 (N_33216,N_32764,N_32848);
nor U33217 (N_33217,N_32863,N_32901);
or U33218 (N_33218,N_32945,N_32787);
xnor U33219 (N_33219,N_32894,N_32994);
nor U33220 (N_33220,N_32928,N_32932);
nand U33221 (N_33221,N_32943,N_32882);
nor U33222 (N_33222,N_32812,N_32940);
xnor U33223 (N_33223,N_32911,N_32907);
nor U33224 (N_33224,N_32896,N_32801);
nand U33225 (N_33225,N_32883,N_32893);
nand U33226 (N_33226,N_32909,N_32920);
xor U33227 (N_33227,N_32917,N_32927);
or U33228 (N_33228,N_32808,N_32778);
xor U33229 (N_33229,N_32825,N_32808);
and U33230 (N_33230,N_32848,N_32985);
xnor U33231 (N_33231,N_32896,N_32934);
and U33232 (N_33232,N_32869,N_32963);
xnor U33233 (N_33233,N_32863,N_32993);
nor U33234 (N_33234,N_32844,N_32796);
xor U33235 (N_33235,N_32918,N_32871);
xor U33236 (N_33236,N_32758,N_32936);
nand U33237 (N_33237,N_32788,N_32880);
or U33238 (N_33238,N_32857,N_32800);
or U33239 (N_33239,N_32926,N_32869);
xor U33240 (N_33240,N_32982,N_32933);
xor U33241 (N_33241,N_32902,N_32876);
xor U33242 (N_33242,N_32865,N_32788);
or U33243 (N_33243,N_32784,N_32992);
nand U33244 (N_33244,N_32935,N_32769);
and U33245 (N_33245,N_32806,N_32962);
and U33246 (N_33246,N_32885,N_32855);
and U33247 (N_33247,N_32917,N_32952);
nor U33248 (N_33248,N_32851,N_32911);
and U33249 (N_33249,N_32764,N_32877);
and U33250 (N_33250,N_33155,N_33134);
nand U33251 (N_33251,N_33200,N_33184);
xnor U33252 (N_33252,N_33076,N_33091);
and U33253 (N_33253,N_33154,N_33085);
or U33254 (N_33254,N_33034,N_33088);
nand U33255 (N_33255,N_33008,N_33003);
nand U33256 (N_33256,N_33232,N_33016);
xor U33257 (N_33257,N_33179,N_33055);
or U33258 (N_33258,N_33137,N_33147);
nor U33259 (N_33259,N_33124,N_33056);
xnor U33260 (N_33260,N_33209,N_33130);
and U33261 (N_33261,N_33082,N_33001);
nand U33262 (N_33262,N_33033,N_33065);
nor U33263 (N_33263,N_33216,N_33060);
and U33264 (N_33264,N_33096,N_33111);
or U33265 (N_33265,N_33139,N_33170);
nor U33266 (N_33266,N_33173,N_33078);
nand U33267 (N_33267,N_33140,N_33119);
and U33268 (N_33268,N_33004,N_33046);
nand U33269 (N_33269,N_33141,N_33198);
and U33270 (N_33270,N_33236,N_33213);
xnor U33271 (N_33271,N_33208,N_33148);
xnor U33272 (N_33272,N_33159,N_33166);
and U33273 (N_33273,N_33183,N_33071);
xnor U33274 (N_33274,N_33158,N_33125);
or U33275 (N_33275,N_33029,N_33019);
nand U33276 (N_33276,N_33066,N_33245);
xnor U33277 (N_33277,N_33222,N_33114);
nand U33278 (N_33278,N_33126,N_33075);
or U33279 (N_33279,N_33070,N_33049);
and U33280 (N_33280,N_33117,N_33084);
and U33281 (N_33281,N_33015,N_33249);
or U33282 (N_33282,N_33052,N_33053);
nor U33283 (N_33283,N_33087,N_33247);
and U33284 (N_33284,N_33248,N_33131);
nor U33285 (N_33285,N_33107,N_33187);
nand U33286 (N_33286,N_33108,N_33039);
and U33287 (N_33287,N_33207,N_33010);
or U33288 (N_33288,N_33058,N_33239);
xor U33289 (N_33289,N_33143,N_33097);
or U33290 (N_33290,N_33113,N_33150);
nor U33291 (N_33291,N_33174,N_33229);
nand U33292 (N_33292,N_33109,N_33040);
xnor U33293 (N_33293,N_33128,N_33189);
and U33294 (N_33294,N_33037,N_33152);
nor U33295 (N_33295,N_33181,N_33226);
xnor U33296 (N_33296,N_33202,N_33009);
or U33297 (N_33297,N_33063,N_33211);
nand U33298 (N_33298,N_33241,N_33156);
or U33299 (N_33299,N_33074,N_33079);
or U33300 (N_33300,N_33233,N_33185);
nand U33301 (N_33301,N_33178,N_33116);
or U33302 (N_33302,N_33215,N_33218);
nand U33303 (N_33303,N_33234,N_33204);
nor U33304 (N_33304,N_33112,N_33212);
nand U33305 (N_33305,N_33243,N_33086);
and U33306 (N_33306,N_33106,N_33038);
or U33307 (N_33307,N_33205,N_33242);
or U33308 (N_33308,N_33099,N_33172);
xor U33309 (N_33309,N_33036,N_33118);
or U33310 (N_33310,N_33035,N_33228);
nor U33311 (N_33311,N_33121,N_33146);
xnor U33312 (N_33312,N_33238,N_33018);
nand U33313 (N_33313,N_33094,N_33157);
nand U33314 (N_33314,N_33031,N_33013);
xor U33315 (N_33315,N_33110,N_33014);
and U33316 (N_33316,N_33197,N_33007);
nand U33317 (N_33317,N_33048,N_33221);
xnor U33318 (N_33318,N_33235,N_33098);
nand U33319 (N_33319,N_33244,N_33102);
or U33320 (N_33320,N_33028,N_33201);
xor U33321 (N_33321,N_33095,N_33044);
and U33322 (N_33322,N_33153,N_33214);
nand U33323 (N_33323,N_33127,N_33051);
nand U33324 (N_33324,N_33026,N_33105);
nor U33325 (N_33325,N_33080,N_33050);
and U33326 (N_33326,N_33047,N_33103);
nor U33327 (N_33327,N_33162,N_33192);
nor U33328 (N_33328,N_33024,N_33145);
nand U33329 (N_33329,N_33230,N_33220);
or U33330 (N_33330,N_33129,N_33240);
nor U33331 (N_33331,N_33133,N_33077);
xnor U33332 (N_33332,N_33149,N_33101);
nand U33333 (N_33333,N_33142,N_33136);
and U33334 (N_33334,N_33135,N_33164);
and U33335 (N_33335,N_33180,N_33025);
xnor U33336 (N_33336,N_33196,N_33092);
nor U33337 (N_33337,N_33203,N_33045);
or U33338 (N_33338,N_33123,N_33195);
nor U33339 (N_33339,N_33072,N_33020);
nand U33340 (N_33340,N_33064,N_33163);
xor U33341 (N_33341,N_33224,N_33081);
or U33342 (N_33342,N_33165,N_33167);
and U33343 (N_33343,N_33011,N_33223);
xor U33344 (N_33344,N_33062,N_33017);
xnor U33345 (N_33345,N_33231,N_33237);
nand U33346 (N_33346,N_33169,N_33093);
and U33347 (N_33347,N_33191,N_33002);
nor U33348 (N_33348,N_33089,N_33000);
nor U33349 (N_33349,N_33030,N_33041);
and U33350 (N_33350,N_33083,N_33182);
nor U33351 (N_33351,N_33246,N_33067);
nand U33352 (N_33352,N_33190,N_33032);
nor U33353 (N_33353,N_33061,N_33069);
xor U33354 (N_33354,N_33073,N_33193);
xor U33355 (N_33355,N_33021,N_33005);
or U33356 (N_33356,N_33219,N_33012);
nor U33357 (N_33357,N_33199,N_33206);
and U33358 (N_33358,N_33138,N_33217);
nand U33359 (N_33359,N_33068,N_33115);
or U33360 (N_33360,N_33054,N_33090);
or U33361 (N_33361,N_33171,N_33104);
or U33362 (N_33362,N_33194,N_33023);
xor U33363 (N_33363,N_33100,N_33120);
and U33364 (N_33364,N_33177,N_33188);
nand U33365 (N_33365,N_33210,N_33168);
and U33366 (N_33366,N_33151,N_33227);
xnor U33367 (N_33367,N_33027,N_33043);
xor U33368 (N_33368,N_33059,N_33042);
nor U33369 (N_33369,N_33225,N_33161);
nand U33370 (N_33370,N_33160,N_33186);
nor U33371 (N_33371,N_33176,N_33057);
or U33372 (N_33372,N_33144,N_33006);
nand U33373 (N_33373,N_33022,N_33175);
nor U33374 (N_33374,N_33132,N_33122);
nor U33375 (N_33375,N_33241,N_33082);
or U33376 (N_33376,N_33196,N_33045);
and U33377 (N_33377,N_33145,N_33160);
nand U33378 (N_33378,N_33034,N_33090);
or U33379 (N_33379,N_33182,N_33077);
xnor U33380 (N_33380,N_33000,N_33020);
nand U33381 (N_33381,N_33076,N_33021);
nor U33382 (N_33382,N_33147,N_33188);
xor U33383 (N_33383,N_33143,N_33196);
nor U33384 (N_33384,N_33187,N_33202);
nand U33385 (N_33385,N_33016,N_33007);
xor U33386 (N_33386,N_33119,N_33044);
nor U33387 (N_33387,N_33204,N_33198);
nor U33388 (N_33388,N_33028,N_33186);
and U33389 (N_33389,N_33245,N_33198);
xor U33390 (N_33390,N_33103,N_33038);
or U33391 (N_33391,N_33020,N_33245);
nor U33392 (N_33392,N_33051,N_33066);
nor U33393 (N_33393,N_33248,N_33155);
xnor U33394 (N_33394,N_33209,N_33190);
and U33395 (N_33395,N_33183,N_33098);
or U33396 (N_33396,N_33177,N_33097);
and U33397 (N_33397,N_33149,N_33233);
nand U33398 (N_33398,N_33159,N_33134);
xnor U33399 (N_33399,N_33210,N_33119);
nand U33400 (N_33400,N_33071,N_33110);
and U33401 (N_33401,N_33048,N_33198);
nand U33402 (N_33402,N_33098,N_33023);
xor U33403 (N_33403,N_33062,N_33107);
xor U33404 (N_33404,N_33162,N_33121);
xnor U33405 (N_33405,N_33229,N_33246);
nand U33406 (N_33406,N_33091,N_33041);
and U33407 (N_33407,N_33223,N_33024);
and U33408 (N_33408,N_33221,N_33232);
nand U33409 (N_33409,N_33196,N_33055);
nand U33410 (N_33410,N_33181,N_33052);
nor U33411 (N_33411,N_33237,N_33011);
nor U33412 (N_33412,N_33101,N_33161);
or U33413 (N_33413,N_33161,N_33073);
xnor U33414 (N_33414,N_33074,N_33008);
xor U33415 (N_33415,N_33228,N_33084);
nand U33416 (N_33416,N_33014,N_33066);
or U33417 (N_33417,N_33163,N_33170);
xor U33418 (N_33418,N_33074,N_33178);
nor U33419 (N_33419,N_33010,N_33233);
or U33420 (N_33420,N_33232,N_33116);
nand U33421 (N_33421,N_33047,N_33163);
and U33422 (N_33422,N_33072,N_33092);
xnor U33423 (N_33423,N_33147,N_33061);
and U33424 (N_33424,N_33048,N_33206);
or U33425 (N_33425,N_33098,N_33198);
and U33426 (N_33426,N_33120,N_33044);
and U33427 (N_33427,N_33079,N_33116);
nand U33428 (N_33428,N_33242,N_33021);
or U33429 (N_33429,N_33135,N_33183);
and U33430 (N_33430,N_33208,N_33224);
nor U33431 (N_33431,N_33092,N_33074);
and U33432 (N_33432,N_33034,N_33187);
or U33433 (N_33433,N_33007,N_33054);
xnor U33434 (N_33434,N_33045,N_33130);
and U33435 (N_33435,N_33183,N_33054);
xnor U33436 (N_33436,N_33121,N_33046);
nand U33437 (N_33437,N_33021,N_33077);
or U33438 (N_33438,N_33068,N_33092);
or U33439 (N_33439,N_33074,N_33135);
and U33440 (N_33440,N_33010,N_33229);
and U33441 (N_33441,N_33121,N_33246);
or U33442 (N_33442,N_33040,N_33042);
and U33443 (N_33443,N_33028,N_33031);
and U33444 (N_33444,N_33100,N_33013);
and U33445 (N_33445,N_33214,N_33145);
nor U33446 (N_33446,N_33208,N_33219);
xnor U33447 (N_33447,N_33029,N_33232);
xnor U33448 (N_33448,N_33083,N_33122);
nand U33449 (N_33449,N_33025,N_33150);
and U33450 (N_33450,N_33210,N_33077);
nor U33451 (N_33451,N_33038,N_33168);
nand U33452 (N_33452,N_33241,N_33181);
nand U33453 (N_33453,N_33193,N_33054);
or U33454 (N_33454,N_33160,N_33205);
and U33455 (N_33455,N_33120,N_33003);
nand U33456 (N_33456,N_33045,N_33153);
and U33457 (N_33457,N_33228,N_33113);
nor U33458 (N_33458,N_33232,N_33239);
nand U33459 (N_33459,N_33094,N_33028);
nand U33460 (N_33460,N_33219,N_33149);
xnor U33461 (N_33461,N_33203,N_33140);
xnor U33462 (N_33462,N_33013,N_33242);
nand U33463 (N_33463,N_33029,N_33075);
xnor U33464 (N_33464,N_33113,N_33062);
and U33465 (N_33465,N_33140,N_33130);
nand U33466 (N_33466,N_33226,N_33003);
nor U33467 (N_33467,N_33180,N_33186);
nor U33468 (N_33468,N_33027,N_33029);
nor U33469 (N_33469,N_33055,N_33059);
nor U33470 (N_33470,N_33221,N_33029);
nand U33471 (N_33471,N_33117,N_33026);
or U33472 (N_33472,N_33177,N_33003);
and U33473 (N_33473,N_33216,N_33113);
or U33474 (N_33474,N_33162,N_33091);
or U33475 (N_33475,N_33214,N_33030);
nand U33476 (N_33476,N_33246,N_33162);
nand U33477 (N_33477,N_33158,N_33130);
nand U33478 (N_33478,N_33162,N_33005);
nor U33479 (N_33479,N_33103,N_33164);
xor U33480 (N_33480,N_33244,N_33153);
or U33481 (N_33481,N_33003,N_33002);
xor U33482 (N_33482,N_33146,N_33044);
nand U33483 (N_33483,N_33018,N_33242);
or U33484 (N_33484,N_33240,N_33125);
xnor U33485 (N_33485,N_33017,N_33154);
nand U33486 (N_33486,N_33157,N_33018);
and U33487 (N_33487,N_33069,N_33225);
or U33488 (N_33488,N_33103,N_33174);
nor U33489 (N_33489,N_33225,N_33207);
or U33490 (N_33490,N_33115,N_33210);
or U33491 (N_33491,N_33078,N_33135);
and U33492 (N_33492,N_33097,N_33167);
nor U33493 (N_33493,N_33080,N_33203);
nor U33494 (N_33494,N_33053,N_33131);
or U33495 (N_33495,N_33212,N_33040);
nand U33496 (N_33496,N_33018,N_33105);
xor U33497 (N_33497,N_33073,N_33107);
or U33498 (N_33498,N_33023,N_33083);
nor U33499 (N_33499,N_33170,N_33192);
or U33500 (N_33500,N_33300,N_33376);
nand U33501 (N_33501,N_33260,N_33261);
xor U33502 (N_33502,N_33262,N_33280);
nand U33503 (N_33503,N_33383,N_33309);
or U33504 (N_33504,N_33380,N_33359);
and U33505 (N_33505,N_33445,N_33282);
nand U33506 (N_33506,N_33346,N_33312);
xor U33507 (N_33507,N_33281,N_33434);
or U33508 (N_33508,N_33394,N_33420);
nand U33509 (N_33509,N_33306,N_33360);
nor U33510 (N_33510,N_33259,N_33453);
nand U33511 (N_33511,N_33494,N_33456);
nand U33512 (N_33512,N_33419,N_33322);
nor U33513 (N_33513,N_33329,N_33374);
nand U33514 (N_33514,N_33484,N_33341);
or U33515 (N_33515,N_33366,N_33271);
nand U33516 (N_33516,N_33303,N_33370);
nor U33517 (N_33517,N_33351,N_33408);
xnor U33518 (N_33518,N_33317,N_33294);
nand U33519 (N_33519,N_33290,N_33468);
nand U33520 (N_33520,N_33490,N_33495);
or U33521 (N_33521,N_33373,N_33343);
nor U33522 (N_33522,N_33263,N_33340);
xor U33523 (N_33523,N_33257,N_33333);
xnor U33524 (N_33524,N_33254,N_33289);
or U33525 (N_33525,N_33472,N_33273);
xnor U33526 (N_33526,N_33344,N_33311);
and U33527 (N_33527,N_33488,N_33279);
xnor U33528 (N_33528,N_33362,N_33414);
nand U33529 (N_33529,N_33301,N_33473);
or U33530 (N_33530,N_33367,N_33403);
and U33531 (N_33531,N_33441,N_33493);
nand U33532 (N_33532,N_33424,N_33497);
nor U33533 (N_33533,N_33267,N_33285);
nor U33534 (N_33534,N_33327,N_33252);
and U33535 (N_33535,N_33391,N_33265);
nor U33536 (N_33536,N_33464,N_33481);
nand U33537 (N_33537,N_33363,N_33286);
or U33538 (N_33538,N_33385,N_33345);
or U33539 (N_33539,N_33466,N_33264);
and U33540 (N_33540,N_33469,N_33347);
nor U33541 (N_33541,N_33392,N_33284);
or U33542 (N_33542,N_33283,N_33378);
nand U33543 (N_33543,N_33353,N_33297);
nor U33544 (N_33544,N_33478,N_33358);
xnor U33545 (N_33545,N_33407,N_33357);
nand U33546 (N_33546,N_33399,N_33298);
nor U33547 (N_33547,N_33452,N_33411);
nor U33548 (N_33548,N_33389,N_33498);
nand U33549 (N_33549,N_33320,N_33471);
nor U33550 (N_33550,N_33477,N_33275);
nor U33551 (N_33551,N_33336,N_33458);
nor U33552 (N_33552,N_33324,N_33272);
or U33553 (N_33553,N_33379,N_33395);
nand U33554 (N_33554,N_33465,N_33323);
xor U33555 (N_33555,N_33486,N_33328);
and U33556 (N_33556,N_33470,N_33483);
or U33557 (N_33557,N_33292,N_33446);
nand U33558 (N_33558,N_33390,N_33430);
and U33559 (N_33559,N_33332,N_33296);
xor U33560 (N_33560,N_33269,N_33369);
and U33561 (N_33561,N_33314,N_33382);
xnor U33562 (N_33562,N_33476,N_33404);
and U33563 (N_33563,N_33426,N_33308);
nand U33564 (N_33564,N_33480,N_33432);
nand U33565 (N_33565,N_33461,N_33428);
or U33566 (N_33566,N_33293,N_33489);
or U33567 (N_33567,N_33406,N_33318);
nor U33568 (N_33568,N_33416,N_33425);
or U33569 (N_33569,N_33496,N_33485);
nor U33570 (N_33570,N_33460,N_33474);
nand U33571 (N_33571,N_33361,N_33413);
or U33572 (N_33572,N_33276,N_33335);
or U33573 (N_33573,N_33393,N_33482);
nand U33574 (N_33574,N_33331,N_33454);
xor U33575 (N_33575,N_33371,N_33352);
or U33576 (N_33576,N_33386,N_33338);
nor U33577 (N_33577,N_33409,N_33295);
or U33578 (N_33578,N_33450,N_33436);
or U33579 (N_33579,N_33348,N_33457);
or U33580 (N_33580,N_33449,N_33487);
xor U33581 (N_33581,N_33277,N_33268);
or U33582 (N_33582,N_33455,N_33440);
or U33583 (N_33583,N_33448,N_33305);
xnor U33584 (N_33584,N_33415,N_33253);
and U33585 (N_33585,N_33326,N_33310);
or U33586 (N_33586,N_33435,N_33319);
nor U33587 (N_33587,N_33372,N_33307);
xnor U33588 (N_33588,N_33429,N_33447);
or U33589 (N_33589,N_33421,N_33339);
and U33590 (N_33590,N_33475,N_33398);
nor U33591 (N_33591,N_33384,N_33401);
nand U33592 (N_33592,N_33459,N_33304);
xnor U33593 (N_33593,N_33479,N_33334);
and U33594 (N_33594,N_33388,N_33377);
nand U33595 (N_33595,N_33356,N_33443);
and U33596 (N_33596,N_33499,N_33274);
or U33597 (N_33597,N_33349,N_33412);
nor U33598 (N_33598,N_33337,N_33270);
xor U33599 (N_33599,N_33330,N_33256);
and U33600 (N_33600,N_33375,N_33278);
nor U33601 (N_33601,N_33410,N_33368);
or U33602 (N_33602,N_33400,N_33402);
and U33603 (N_33603,N_33316,N_33405);
nand U33604 (N_33604,N_33266,N_33437);
or U33605 (N_33605,N_33355,N_33491);
xor U33606 (N_33606,N_33291,N_33433);
nor U33607 (N_33607,N_33463,N_33251);
and U33608 (N_33608,N_33451,N_33427);
and U33609 (N_33609,N_33422,N_33396);
xnor U33610 (N_33610,N_33417,N_33255);
or U33611 (N_33611,N_33439,N_33381);
nor U33612 (N_33612,N_33492,N_33354);
nor U33613 (N_33613,N_33258,N_33313);
or U33614 (N_33614,N_33442,N_33467);
nand U33615 (N_33615,N_33325,N_33250);
xor U33616 (N_33616,N_33365,N_33431);
nand U33617 (N_33617,N_33444,N_33438);
and U33618 (N_33618,N_33302,N_33397);
or U33619 (N_33619,N_33387,N_33364);
nor U33620 (N_33620,N_33423,N_33315);
nand U33621 (N_33621,N_33350,N_33418);
xnor U33622 (N_33622,N_33342,N_33299);
and U33623 (N_33623,N_33321,N_33288);
xnor U33624 (N_33624,N_33287,N_33462);
nand U33625 (N_33625,N_33298,N_33291);
nand U33626 (N_33626,N_33282,N_33342);
nand U33627 (N_33627,N_33324,N_33402);
and U33628 (N_33628,N_33260,N_33481);
nor U33629 (N_33629,N_33282,N_33385);
and U33630 (N_33630,N_33258,N_33341);
nor U33631 (N_33631,N_33330,N_33373);
xor U33632 (N_33632,N_33253,N_33348);
xnor U33633 (N_33633,N_33394,N_33378);
or U33634 (N_33634,N_33270,N_33464);
xor U33635 (N_33635,N_33423,N_33402);
nor U33636 (N_33636,N_33464,N_33449);
nor U33637 (N_33637,N_33292,N_33423);
and U33638 (N_33638,N_33252,N_33354);
xnor U33639 (N_33639,N_33267,N_33385);
xnor U33640 (N_33640,N_33334,N_33461);
and U33641 (N_33641,N_33393,N_33334);
nor U33642 (N_33642,N_33378,N_33324);
nand U33643 (N_33643,N_33302,N_33353);
nor U33644 (N_33644,N_33460,N_33361);
or U33645 (N_33645,N_33359,N_33325);
nand U33646 (N_33646,N_33453,N_33360);
or U33647 (N_33647,N_33334,N_33369);
xor U33648 (N_33648,N_33267,N_33403);
nand U33649 (N_33649,N_33300,N_33344);
nor U33650 (N_33650,N_33369,N_33452);
nand U33651 (N_33651,N_33465,N_33399);
nand U33652 (N_33652,N_33438,N_33455);
or U33653 (N_33653,N_33310,N_33402);
and U33654 (N_33654,N_33357,N_33273);
or U33655 (N_33655,N_33294,N_33445);
nor U33656 (N_33656,N_33318,N_33300);
nor U33657 (N_33657,N_33453,N_33306);
nand U33658 (N_33658,N_33268,N_33477);
nor U33659 (N_33659,N_33347,N_33441);
or U33660 (N_33660,N_33276,N_33410);
nor U33661 (N_33661,N_33277,N_33315);
xnor U33662 (N_33662,N_33371,N_33363);
xnor U33663 (N_33663,N_33415,N_33300);
nand U33664 (N_33664,N_33371,N_33455);
nor U33665 (N_33665,N_33375,N_33350);
or U33666 (N_33666,N_33431,N_33273);
nand U33667 (N_33667,N_33316,N_33273);
nor U33668 (N_33668,N_33447,N_33296);
or U33669 (N_33669,N_33398,N_33322);
nand U33670 (N_33670,N_33250,N_33425);
nand U33671 (N_33671,N_33390,N_33269);
and U33672 (N_33672,N_33444,N_33254);
nor U33673 (N_33673,N_33378,N_33437);
nand U33674 (N_33674,N_33347,N_33404);
xnor U33675 (N_33675,N_33343,N_33416);
nor U33676 (N_33676,N_33277,N_33312);
and U33677 (N_33677,N_33328,N_33262);
xnor U33678 (N_33678,N_33288,N_33299);
xnor U33679 (N_33679,N_33449,N_33436);
and U33680 (N_33680,N_33286,N_33290);
or U33681 (N_33681,N_33290,N_33482);
xor U33682 (N_33682,N_33353,N_33384);
nand U33683 (N_33683,N_33266,N_33391);
and U33684 (N_33684,N_33426,N_33258);
nor U33685 (N_33685,N_33292,N_33330);
or U33686 (N_33686,N_33389,N_33401);
and U33687 (N_33687,N_33292,N_33415);
xnor U33688 (N_33688,N_33302,N_33449);
nand U33689 (N_33689,N_33492,N_33487);
xor U33690 (N_33690,N_33293,N_33317);
nand U33691 (N_33691,N_33262,N_33466);
and U33692 (N_33692,N_33424,N_33293);
xor U33693 (N_33693,N_33322,N_33456);
xnor U33694 (N_33694,N_33399,N_33253);
or U33695 (N_33695,N_33455,N_33475);
nand U33696 (N_33696,N_33251,N_33300);
nand U33697 (N_33697,N_33422,N_33302);
nand U33698 (N_33698,N_33464,N_33445);
xor U33699 (N_33699,N_33373,N_33469);
or U33700 (N_33700,N_33470,N_33480);
xor U33701 (N_33701,N_33324,N_33401);
nor U33702 (N_33702,N_33410,N_33297);
or U33703 (N_33703,N_33448,N_33441);
nor U33704 (N_33704,N_33494,N_33498);
or U33705 (N_33705,N_33496,N_33366);
nand U33706 (N_33706,N_33401,N_33421);
and U33707 (N_33707,N_33412,N_33260);
and U33708 (N_33708,N_33409,N_33348);
xnor U33709 (N_33709,N_33395,N_33384);
nand U33710 (N_33710,N_33424,N_33339);
nand U33711 (N_33711,N_33462,N_33463);
xnor U33712 (N_33712,N_33443,N_33393);
nor U33713 (N_33713,N_33471,N_33394);
and U33714 (N_33714,N_33412,N_33402);
and U33715 (N_33715,N_33365,N_33423);
nand U33716 (N_33716,N_33396,N_33284);
xnor U33717 (N_33717,N_33330,N_33325);
nand U33718 (N_33718,N_33277,N_33389);
and U33719 (N_33719,N_33329,N_33422);
nor U33720 (N_33720,N_33484,N_33280);
or U33721 (N_33721,N_33459,N_33390);
or U33722 (N_33722,N_33352,N_33358);
nor U33723 (N_33723,N_33473,N_33315);
or U33724 (N_33724,N_33464,N_33496);
xnor U33725 (N_33725,N_33406,N_33437);
or U33726 (N_33726,N_33466,N_33281);
or U33727 (N_33727,N_33273,N_33421);
nand U33728 (N_33728,N_33378,N_33493);
or U33729 (N_33729,N_33398,N_33345);
and U33730 (N_33730,N_33379,N_33298);
nand U33731 (N_33731,N_33281,N_33284);
nor U33732 (N_33732,N_33476,N_33462);
nor U33733 (N_33733,N_33330,N_33390);
or U33734 (N_33734,N_33492,N_33457);
nand U33735 (N_33735,N_33442,N_33428);
nor U33736 (N_33736,N_33409,N_33498);
nor U33737 (N_33737,N_33430,N_33410);
nor U33738 (N_33738,N_33333,N_33251);
xor U33739 (N_33739,N_33314,N_33348);
nand U33740 (N_33740,N_33499,N_33296);
and U33741 (N_33741,N_33396,N_33281);
nor U33742 (N_33742,N_33336,N_33262);
xnor U33743 (N_33743,N_33471,N_33262);
nor U33744 (N_33744,N_33410,N_33362);
or U33745 (N_33745,N_33307,N_33450);
nand U33746 (N_33746,N_33413,N_33448);
xor U33747 (N_33747,N_33389,N_33485);
nand U33748 (N_33748,N_33319,N_33444);
nand U33749 (N_33749,N_33496,N_33491);
nor U33750 (N_33750,N_33728,N_33712);
nor U33751 (N_33751,N_33533,N_33564);
xor U33752 (N_33752,N_33686,N_33709);
and U33753 (N_33753,N_33741,N_33676);
nor U33754 (N_33754,N_33550,N_33559);
nand U33755 (N_33755,N_33706,N_33580);
or U33756 (N_33756,N_33745,N_33684);
or U33757 (N_33757,N_33589,N_33690);
or U33758 (N_33758,N_33726,N_33625);
or U33759 (N_33759,N_33658,N_33556);
nor U33760 (N_33760,N_33557,N_33668);
and U33761 (N_33761,N_33567,N_33730);
nand U33762 (N_33762,N_33717,N_33599);
nand U33763 (N_33763,N_33651,N_33724);
nand U33764 (N_33764,N_33694,N_33507);
nor U33765 (N_33765,N_33638,N_33672);
xnor U33766 (N_33766,N_33544,N_33572);
or U33767 (N_33767,N_33523,N_33650);
nor U33768 (N_33768,N_33562,N_33683);
nor U33769 (N_33769,N_33721,N_33525);
and U33770 (N_33770,N_33646,N_33570);
nor U33771 (N_33771,N_33510,N_33629);
and U33772 (N_33772,N_33720,N_33667);
nor U33773 (N_33773,N_33675,N_33665);
or U33774 (N_33774,N_33620,N_33538);
nand U33775 (N_33775,N_33504,N_33532);
xnor U33776 (N_33776,N_33663,N_33633);
and U33777 (N_33777,N_33531,N_33699);
and U33778 (N_33778,N_33627,N_33641);
nor U33779 (N_33779,N_33588,N_33542);
or U33780 (N_33780,N_33613,N_33615);
and U33781 (N_33781,N_33614,N_33734);
nand U33782 (N_33782,N_33673,N_33630);
nand U33783 (N_33783,N_33695,N_33514);
or U33784 (N_33784,N_33568,N_33597);
and U33785 (N_33785,N_33601,N_33592);
or U33786 (N_33786,N_33579,N_33591);
nor U33787 (N_33787,N_33685,N_33689);
nor U33788 (N_33788,N_33600,N_33594);
nor U33789 (N_33789,N_33539,N_33565);
nand U33790 (N_33790,N_33583,N_33590);
or U33791 (N_33791,N_33652,N_33576);
and U33792 (N_33792,N_33598,N_33534);
xnor U33793 (N_33793,N_33698,N_33512);
nor U33794 (N_33794,N_33605,N_33656);
nor U33795 (N_33795,N_33554,N_33528);
xor U33796 (N_33796,N_33513,N_33527);
xor U33797 (N_33797,N_33563,N_33596);
and U33798 (N_33798,N_33716,N_33645);
nand U33799 (N_33799,N_33737,N_33704);
nand U33800 (N_33800,N_33587,N_33648);
and U33801 (N_33801,N_33657,N_33653);
xnor U33802 (N_33802,N_33530,N_33623);
nor U33803 (N_33803,N_33607,N_33549);
or U33804 (N_33804,N_33518,N_33707);
and U33805 (N_33805,N_33671,N_33618);
nand U33806 (N_33806,N_33746,N_33691);
or U33807 (N_33807,N_33541,N_33516);
and U33808 (N_33808,N_33526,N_33509);
or U33809 (N_33809,N_33515,N_33543);
nand U33810 (N_33810,N_33626,N_33740);
and U33811 (N_33811,N_33708,N_33582);
and U33812 (N_33812,N_33616,N_33603);
nor U33813 (N_33813,N_33586,N_33508);
nor U33814 (N_33814,N_33643,N_33631);
or U33815 (N_33815,N_33732,N_33609);
nor U33816 (N_33816,N_33692,N_33678);
nand U33817 (N_33817,N_33622,N_33578);
or U33818 (N_33818,N_33696,N_33608);
nand U33819 (N_33819,N_33624,N_33647);
or U33820 (N_33820,N_33640,N_33529);
nand U33821 (N_33821,N_33661,N_33610);
or U33822 (N_33822,N_33522,N_33577);
and U33823 (N_33823,N_33602,N_33584);
nand U33824 (N_33824,N_33546,N_33574);
nor U33825 (N_33825,N_33738,N_33679);
xor U33826 (N_33826,N_33537,N_33511);
and U33827 (N_33827,N_33634,N_33552);
nor U33828 (N_33828,N_33617,N_33621);
xnor U33829 (N_33829,N_33722,N_33705);
xnor U33830 (N_33830,N_33575,N_33674);
nand U33831 (N_33831,N_33519,N_33748);
xor U33832 (N_33832,N_33566,N_33500);
nand U33833 (N_33833,N_33733,N_33561);
or U33834 (N_33834,N_33560,N_33711);
nor U33835 (N_33835,N_33662,N_33693);
nor U33836 (N_33836,N_33700,N_33535);
nand U33837 (N_33837,N_33612,N_33581);
xor U33838 (N_33838,N_33713,N_33747);
nand U33839 (N_33839,N_33506,N_33619);
and U33840 (N_33840,N_33517,N_33555);
and U33841 (N_33841,N_33731,N_33719);
and U33842 (N_33842,N_33502,N_33670);
nor U33843 (N_33843,N_33736,N_33639);
nand U33844 (N_33844,N_33688,N_33729);
and U33845 (N_33845,N_33505,N_33606);
nand U33846 (N_33846,N_33501,N_33710);
nand U33847 (N_33847,N_33725,N_33585);
or U33848 (N_33848,N_33742,N_33604);
nor U33849 (N_33849,N_33701,N_33545);
nand U33850 (N_33850,N_33636,N_33659);
xnor U33851 (N_33851,N_33735,N_33520);
nand U33852 (N_33852,N_33715,N_33681);
nand U33853 (N_33853,N_33703,N_33655);
nor U33854 (N_33854,N_33743,N_33540);
or U33855 (N_33855,N_33553,N_33573);
xnor U33856 (N_33856,N_33660,N_33524);
and U33857 (N_33857,N_33551,N_33687);
nor U33858 (N_33858,N_33723,N_33521);
nor U33859 (N_33859,N_33503,N_33649);
xnor U33860 (N_33860,N_33727,N_33593);
and U33861 (N_33861,N_33536,N_33664);
or U33862 (N_33862,N_33714,N_33611);
and U33863 (N_33863,N_33680,N_33644);
nand U33864 (N_33864,N_33595,N_33635);
and U33865 (N_33865,N_33628,N_33548);
nor U33866 (N_33866,N_33669,N_33571);
or U33867 (N_33867,N_33682,N_33677);
and U33868 (N_33868,N_33569,N_33642);
xor U33869 (N_33869,N_33697,N_33547);
and U33870 (N_33870,N_33744,N_33702);
nor U33871 (N_33871,N_33739,N_33654);
and U33872 (N_33872,N_33749,N_33558);
nor U33873 (N_33873,N_33718,N_33666);
and U33874 (N_33874,N_33632,N_33637);
xor U33875 (N_33875,N_33514,N_33622);
nor U33876 (N_33876,N_33721,N_33681);
xnor U33877 (N_33877,N_33500,N_33682);
nand U33878 (N_33878,N_33715,N_33700);
nand U33879 (N_33879,N_33609,N_33589);
and U33880 (N_33880,N_33734,N_33626);
or U33881 (N_33881,N_33656,N_33597);
or U33882 (N_33882,N_33687,N_33727);
nand U33883 (N_33883,N_33624,N_33690);
nor U33884 (N_33884,N_33540,N_33533);
xnor U33885 (N_33885,N_33667,N_33563);
nand U33886 (N_33886,N_33720,N_33665);
nand U33887 (N_33887,N_33743,N_33502);
and U33888 (N_33888,N_33669,N_33513);
xor U33889 (N_33889,N_33684,N_33508);
nand U33890 (N_33890,N_33610,N_33730);
nand U33891 (N_33891,N_33571,N_33646);
nor U33892 (N_33892,N_33511,N_33710);
or U33893 (N_33893,N_33732,N_33712);
xor U33894 (N_33894,N_33584,N_33595);
xor U33895 (N_33895,N_33729,N_33692);
nand U33896 (N_33896,N_33682,N_33627);
nor U33897 (N_33897,N_33621,N_33746);
nand U33898 (N_33898,N_33511,N_33674);
nand U33899 (N_33899,N_33657,N_33537);
xnor U33900 (N_33900,N_33626,N_33720);
xor U33901 (N_33901,N_33613,N_33512);
nor U33902 (N_33902,N_33547,N_33699);
or U33903 (N_33903,N_33610,N_33591);
or U33904 (N_33904,N_33533,N_33501);
xnor U33905 (N_33905,N_33641,N_33529);
nor U33906 (N_33906,N_33504,N_33588);
xnor U33907 (N_33907,N_33536,N_33721);
or U33908 (N_33908,N_33611,N_33693);
nand U33909 (N_33909,N_33557,N_33716);
nor U33910 (N_33910,N_33535,N_33682);
xnor U33911 (N_33911,N_33747,N_33607);
and U33912 (N_33912,N_33619,N_33525);
nor U33913 (N_33913,N_33521,N_33537);
nand U33914 (N_33914,N_33693,N_33604);
nand U33915 (N_33915,N_33503,N_33564);
nand U33916 (N_33916,N_33526,N_33670);
xnor U33917 (N_33917,N_33523,N_33676);
nand U33918 (N_33918,N_33650,N_33684);
xnor U33919 (N_33919,N_33545,N_33565);
or U33920 (N_33920,N_33663,N_33660);
xor U33921 (N_33921,N_33670,N_33625);
and U33922 (N_33922,N_33698,N_33642);
and U33923 (N_33923,N_33513,N_33549);
nor U33924 (N_33924,N_33702,N_33529);
or U33925 (N_33925,N_33632,N_33659);
nand U33926 (N_33926,N_33514,N_33568);
or U33927 (N_33927,N_33690,N_33681);
or U33928 (N_33928,N_33551,N_33649);
or U33929 (N_33929,N_33672,N_33648);
nand U33930 (N_33930,N_33536,N_33566);
and U33931 (N_33931,N_33519,N_33520);
and U33932 (N_33932,N_33729,N_33550);
xnor U33933 (N_33933,N_33653,N_33723);
or U33934 (N_33934,N_33519,N_33571);
or U33935 (N_33935,N_33502,N_33681);
and U33936 (N_33936,N_33716,N_33593);
nor U33937 (N_33937,N_33535,N_33627);
and U33938 (N_33938,N_33650,N_33620);
and U33939 (N_33939,N_33645,N_33506);
nor U33940 (N_33940,N_33694,N_33738);
xor U33941 (N_33941,N_33507,N_33571);
xor U33942 (N_33942,N_33717,N_33742);
or U33943 (N_33943,N_33727,N_33530);
nor U33944 (N_33944,N_33586,N_33579);
or U33945 (N_33945,N_33679,N_33703);
nor U33946 (N_33946,N_33526,N_33696);
nor U33947 (N_33947,N_33649,N_33528);
or U33948 (N_33948,N_33510,N_33617);
xnor U33949 (N_33949,N_33619,N_33696);
and U33950 (N_33950,N_33549,N_33505);
xor U33951 (N_33951,N_33549,N_33609);
nand U33952 (N_33952,N_33622,N_33749);
nor U33953 (N_33953,N_33664,N_33508);
and U33954 (N_33954,N_33539,N_33606);
or U33955 (N_33955,N_33719,N_33664);
xnor U33956 (N_33956,N_33619,N_33569);
nor U33957 (N_33957,N_33671,N_33702);
xnor U33958 (N_33958,N_33608,N_33652);
nor U33959 (N_33959,N_33532,N_33513);
and U33960 (N_33960,N_33556,N_33689);
xnor U33961 (N_33961,N_33663,N_33725);
and U33962 (N_33962,N_33719,N_33682);
nor U33963 (N_33963,N_33617,N_33515);
xor U33964 (N_33964,N_33650,N_33691);
and U33965 (N_33965,N_33604,N_33585);
xnor U33966 (N_33966,N_33740,N_33588);
or U33967 (N_33967,N_33710,N_33679);
or U33968 (N_33968,N_33644,N_33598);
xor U33969 (N_33969,N_33745,N_33625);
and U33970 (N_33970,N_33615,N_33582);
or U33971 (N_33971,N_33685,N_33579);
and U33972 (N_33972,N_33664,N_33574);
and U33973 (N_33973,N_33581,N_33673);
nand U33974 (N_33974,N_33654,N_33680);
nand U33975 (N_33975,N_33612,N_33596);
xnor U33976 (N_33976,N_33551,N_33595);
and U33977 (N_33977,N_33533,N_33697);
or U33978 (N_33978,N_33622,N_33746);
and U33979 (N_33979,N_33709,N_33672);
or U33980 (N_33980,N_33667,N_33548);
or U33981 (N_33981,N_33603,N_33685);
nor U33982 (N_33982,N_33705,N_33532);
nor U33983 (N_33983,N_33645,N_33541);
nand U33984 (N_33984,N_33520,N_33727);
or U33985 (N_33985,N_33618,N_33732);
xnor U33986 (N_33986,N_33649,N_33700);
nor U33987 (N_33987,N_33504,N_33745);
nand U33988 (N_33988,N_33507,N_33657);
or U33989 (N_33989,N_33611,N_33699);
and U33990 (N_33990,N_33717,N_33654);
and U33991 (N_33991,N_33627,N_33564);
nor U33992 (N_33992,N_33609,N_33642);
or U33993 (N_33993,N_33644,N_33654);
xor U33994 (N_33994,N_33630,N_33734);
and U33995 (N_33995,N_33645,N_33529);
xor U33996 (N_33996,N_33712,N_33585);
or U33997 (N_33997,N_33672,N_33548);
or U33998 (N_33998,N_33674,N_33671);
xnor U33999 (N_33999,N_33657,N_33530);
and U34000 (N_34000,N_33875,N_33978);
xor U34001 (N_34001,N_33835,N_33874);
nand U34002 (N_34002,N_33940,N_33948);
nand U34003 (N_34003,N_33869,N_33992);
or U34004 (N_34004,N_33920,N_33906);
and U34005 (N_34005,N_33963,N_33901);
nand U34006 (N_34006,N_33919,N_33872);
or U34007 (N_34007,N_33985,N_33921);
nand U34008 (N_34008,N_33810,N_33947);
or U34009 (N_34009,N_33828,N_33776);
xor U34010 (N_34010,N_33945,N_33786);
or U34011 (N_34011,N_33793,N_33896);
xor U34012 (N_34012,N_33783,N_33836);
and U34013 (N_34013,N_33900,N_33885);
and U34014 (N_34014,N_33808,N_33762);
xnor U34015 (N_34015,N_33818,N_33751);
nand U34016 (N_34016,N_33784,N_33974);
nand U34017 (N_34017,N_33863,N_33880);
xor U34018 (N_34018,N_33763,N_33857);
nor U34019 (N_34019,N_33865,N_33870);
nand U34020 (N_34020,N_33792,N_33803);
xnor U34021 (N_34021,N_33981,N_33767);
xnor U34022 (N_34022,N_33971,N_33859);
nand U34023 (N_34023,N_33922,N_33991);
or U34024 (N_34024,N_33843,N_33798);
or U34025 (N_34025,N_33815,N_33902);
xor U34026 (N_34026,N_33976,N_33856);
nand U34027 (N_34027,N_33779,N_33944);
and U34028 (N_34028,N_33753,N_33941);
xnor U34029 (N_34029,N_33952,N_33782);
or U34030 (N_34030,N_33791,N_33802);
nand U34031 (N_34031,N_33908,N_33912);
and U34032 (N_34032,N_33849,N_33967);
nand U34033 (N_34033,N_33889,N_33755);
xor U34034 (N_34034,N_33807,N_33927);
nand U34035 (N_34035,N_33958,N_33822);
nor U34036 (N_34036,N_33853,N_33917);
nand U34037 (N_34037,N_33916,N_33891);
nor U34038 (N_34038,N_33995,N_33794);
or U34039 (N_34039,N_33984,N_33955);
xor U34040 (N_34040,N_33910,N_33797);
nand U34041 (N_34041,N_33928,N_33897);
nor U34042 (N_34042,N_33997,N_33894);
or U34043 (N_34043,N_33813,N_33913);
nand U34044 (N_34044,N_33766,N_33761);
nand U34045 (N_34045,N_33970,N_33867);
or U34046 (N_34046,N_33787,N_33829);
nand U34047 (N_34047,N_33983,N_33760);
or U34048 (N_34048,N_33858,N_33979);
or U34049 (N_34049,N_33914,N_33980);
and U34050 (N_34050,N_33750,N_33960);
nor U34051 (N_34051,N_33977,N_33778);
nor U34052 (N_34052,N_33809,N_33752);
and U34053 (N_34053,N_33769,N_33820);
nand U34054 (N_34054,N_33986,N_33898);
and U34055 (N_34055,N_33883,N_33957);
xor U34056 (N_34056,N_33969,N_33765);
nor U34057 (N_34057,N_33929,N_33774);
nand U34058 (N_34058,N_33972,N_33993);
nor U34059 (N_34059,N_33890,N_33826);
nor U34060 (N_34060,N_33852,N_33909);
nor U34061 (N_34061,N_33956,N_33805);
xor U34062 (N_34062,N_33942,N_33824);
and U34063 (N_34063,N_33934,N_33895);
xor U34064 (N_34064,N_33832,N_33842);
nand U34065 (N_34065,N_33893,N_33790);
or U34066 (N_34066,N_33770,N_33932);
or U34067 (N_34067,N_33848,N_33772);
nand U34068 (N_34068,N_33982,N_33968);
nand U34069 (N_34069,N_33788,N_33907);
nor U34070 (N_34070,N_33823,N_33975);
xor U34071 (N_34071,N_33878,N_33905);
xor U34072 (N_34072,N_33881,N_33887);
nand U34073 (N_34073,N_33888,N_33918);
xnor U34074 (N_34074,N_33768,N_33953);
and U34075 (N_34075,N_33827,N_33882);
nor U34076 (N_34076,N_33817,N_33994);
xnor U34077 (N_34077,N_33904,N_33833);
nor U34078 (N_34078,N_33946,N_33854);
and U34079 (N_34079,N_33844,N_33951);
or U34080 (N_34080,N_33850,N_33996);
nor U34081 (N_34081,N_33915,N_33847);
nand U34082 (N_34082,N_33924,N_33756);
and U34083 (N_34083,N_33931,N_33877);
nand U34084 (N_34084,N_33830,N_33795);
or U34085 (N_34085,N_33937,N_33962);
or U34086 (N_34086,N_33764,N_33899);
nor U34087 (N_34087,N_33930,N_33838);
or U34088 (N_34088,N_33757,N_33841);
nor U34089 (N_34089,N_33845,N_33825);
nor U34090 (N_34090,N_33939,N_33965);
and U34091 (N_34091,N_33886,N_33804);
nand U34092 (N_34092,N_33911,N_33831);
xnor U34093 (N_34093,N_33864,N_33925);
xor U34094 (N_34094,N_33949,N_33785);
nor U34095 (N_34095,N_33879,N_33990);
or U34096 (N_34096,N_33923,N_33855);
xor U34097 (N_34097,N_33780,N_33871);
nand U34098 (N_34098,N_33821,N_33775);
nor U34099 (N_34099,N_33781,N_33846);
nor U34100 (N_34100,N_33777,N_33840);
nor U34101 (N_34101,N_33812,N_33903);
or U34102 (N_34102,N_33961,N_33861);
nor U34103 (N_34103,N_33873,N_33868);
or U34104 (N_34104,N_33999,N_33959);
nor U34105 (N_34105,N_33964,N_33800);
nor U34106 (N_34106,N_33884,N_33876);
nor U34107 (N_34107,N_33839,N_33801);
nor U34108 (N_34108,N_33796,N_33773);
nand U34109 (N_34109,N_33933,N_33866);
and U34110 (N_34110,N_33862,N_33950);
nor U34111 (N_34111,N_33799,N_33754);
or U34112 (N_34112,N_33989,N_33892);
nand U34113 (N_34113,N_33819,N_33811);
nor U34114 (N_34114,N_33771,N_33998);
or U34115 (N_34115,N_33935,N_33954);
or U34116 (N_34116,N_33988,N_33837);
and U34117 (N_34117,N_33759,N_33943);
or U34118 (N_34118,N_33816,N_33834);
xnor U34119 (N_34119,N_33758,N_33936);
xnor U34120 (N_34120,N_33926,N_33851);
and U34121 (N_34121,N_33814,N_33973);
nand U34122 (N_34122,N_33966,N_33789);
nor U34123 (N_34123,N_33806,N_33987);
xor U34124 (N_34124,N_33860,N_33938);
xor U34125 (N_34125,N_33918,N_33778);
nand U34126 (N_34126,N_33878,N_33965);
nor U34127 (N_34127,N_33848,N_33906);
and U34128 (N_34128,N_33781,N_33852);
nor U34129 (N_34129,N_33995,N_33766);
nand U34130 (N_34130,N_33907,N_33881);
or U34131 (N_34131,N_33806,N_33868);
nor U34132 (N_34132,N_33803,N_33856);
nand U34133 (N_34133,N_33952,N_33811);
nor U34134 (N_34134,N_33880,N_33889);
or U34135 (N_34135,N_33897,N_33801);
nor U34136 (N_34136,N_33965,N_33892);
xnor U34137 (N_34137,N_33828,N_33873);
xor U34138 (N_34138,N_33931,N_33752);
nor U34139 (N_34139,N_33821,N_33844);
nor U34140 (N_34140,N_33952,N_33875);
nor U34141 (N_34141,N_33770,N_33760);
xnor U34142 (N_34142,N_33801,N_33774);
or U34143 (N_34143,N_33877,N_33769);
and U34144 (N_34144,N_33881,N_33860);
xnor U34145 (N_34145,N_33936,N_33871);
nor U34146 (N_34146,N_33837,N_33946);
nand U34147 (N_34147,N_33813,N_33780);
nor U34148 (N_34148,N_33863,N_33855);
nor U34149 (N_34149,N_33985,N_33942);
nor U34150 (N_34150,N_33933,N_33924);
or U34151 (N_34151,N_33927,N_33996);
nand U34152 (N_34152,N_33809,N_33886);
xor U34153 (N_34153,N_33878,N_33834);
nand U34154 (N_34154,N_33983,N_33860);
nor U34155 (N_34155,N_33808,N_33943);
nor U34156 (N_34156,N_33829,N_33796);
and U34157 (N_34157,N_33800,N_33819);
nor U34158 (N_34158,N_33958,N_33971);
or U34159 (N_34159,N_33865,N_33810);
and U34160 (N_34160,N_33912,N_33806);
or U34161 (N_34161,N_33991,N_33900);
nor U34162 (N_34162,N_33778,N_33858);
xor U34163 (N_34163,N_33825,N_33961);
or U34164 (N_34164,N_33919,N_33941);
and U34165 (N_34165,N_33999,N_33973);
nand U34166 (N_34166,N_33893,N_33997);
nor U34167 (N_34167,N_33884,N_33787);
nand U34168 (N_34168,N_33929,N_33853);
or U34169 (N_34169,N_33907,N_33955);
nand U34170 (N_34170,N_33862,N_33873);
or U34171 (N_34171,N_33884,N_33983);
and U34172 (N_34172,N_33974,N_33955);
and U34173 (N_34173,N_33756,N_33840);
xnor U34174 (N_34174,N_33936,N_33850);
nor U34175 (N_34175,N_33815,N_33954);
xnor U34176 (N_34176,N_33968,N_33772);
or U34177 (N_34177,N_33878,N_33898);
xnor U34178 (N_34178,N_33768,N_33757);
or U34179 (N_34179,N_33814,N_33844);
nor U34180 (N_34180,N_33980,N_33797);
nand U34181 (N_34181,N_33848,N_33997);
and U34182 (N_34182,N_33799,N_33998);
nand U34183 (N_34183,N_33863,N_33901);
xnor U34184 (N_34184,N_33942,N_33996);
xor U34185 (N_34185,N_33937,N_33853);
xor U34186 (N_34186,N_33998,N_33888);
and U34187 (N_34187,N_33802,N_33765);
nor U34188 (N_34188,N_33828,N_33866);
nand U34189 (N_34189,N_33895,N_33915);
xnor U34190 (N_34190,N_33898,N_33763);
nand U34191 (N_34191,N_33822,N_33906);
or U34192 (N_34192,N_33888,N_33778);
or U34193 (N_34193,N_33823,N_33965);
nand U34194 (N_34194,N_33914,N_33870);
nor U34195 (N_34195,N_33908,N_33886);
nand U34196 (N_34196,N_33817,N_33785);
nor U34197 (N_34197,N_33799,N_33902);
or U34198 (N_34198,N_33753,N_33801);
and U34199 (N_34199,N_33951,N_33794);
and U34200 (N_34200,N_33844,N_33872);
xnor U34201 (N_34201,N_33936,N_33885);
xnor U34202 (N_34202,N_33962,N_33812);
xnor U34203 (N_34203,N_33933,N_33805);
and U34204 (N_34204,N_33963,N_33840);
nor U34205 (N_34205,N_33899,N_33967);
or U34206 (N_34206,N_33878,N_33929);
nor U34207 (N_34207,N_33889,N_33993);
xor U34208 (N_34208,N_33904,N_33925);
nand U34209 (N_34209,N_33970,N_33854);
xnor U34210 (N_34210,N_33752,N_33944);
or U34211 (N_34211,N_33971,N_33986);
xor U34212 (N_34212,N_33750,N_33826);
nor U34213 (N_34213,N_33832,N_33992);
nor U34214 (N_34214,N_33869,N_33854);
or U34215 (N_34215,N_33873,N_33802);
nor U34216 (N_34216,N_33813,N_33996);
xor U34217 (N_34217,N_33865,N_33855);
xor U34218 (N_34218,N_33830,N_33892);
xor U34219 (N_34219,N_33861,N_33830);
or U34220 (N_34220,N_33936,N_33985);
and U34221 (N_34221,N_33898,N_33876);
and U34222 (N_34222,N_33755,N_33946);
xor U34223 (N_34223,N_33758,N_33946);
nor U34224 (N_34224,N_33851,N_33824);
xor U34225 (N_34225,N_33845,N_33832);
and U34226 (N_34226,N_33886,N_33781);
nand U34227 (N_34227,N_33860,N_33852);
or U34228 (N_34228,N_33762,N_33957);
and U34229 (N_34229,N_33755,N_33843);
xor U34230 (N_34230,N_33986,N_33999);
or U34231 (N_34231,N_33948,N_33790);
nand U34232 (N_34232,N_33789,N_33808);
xor U34233 (N_34233,N_33864,N_33758);
nand U34234 (N_34234,N_33900,N_33931);
nand U34235 (N_34235,N_33784,N_33843);
and U34236 (N_34236,N_33815,N_33992);
nand U34237 (N_34237,N_33898,N_33843);
and U34238 (N_34238,N_33871,N_33785);
xnor U34239 (N_34239,N_33919,N_33770);
xnor U34240 (N_34240,N_33987,N_33914);
nand U34241 (N_34241,N_33967,N_33907);
or U34242 (N_34242,N_33874,N_33917);
or U34243 (N_34243,N_33802,N_33936);
nand U34244 (N_34244,N_33882,N_33843);
and U34245 (N_34245,N_33993,N_33948);
xnor U34246 (N_34246,N_33968,N_33800);
and U34247 (N_34247,N_33789,N_33864);
or U34248 (N_34248,N_33859,N_33760);
xnor U34249 (N_34249,N_33976,N_33994);
and U34250 (N_34250,N_34177,N_34046);
and U34251 (N_34251,N_34003,N_34120);
nor U34252 (N_34252,N_34209,N_34065);
and U34253 (N_34253,N_34213,N_34074);
and U34254 (N_34254,N_34128,N_34064);
or U34255 (N_34255,N_34160,N_34108);
xor U34256 (N_34256,N_34114,N_34144);
nand U34257 (N_34257,N_34097,N_34188);
nand U34258 (N_34258,N_34212,N_34035);
nor U34259 (N_34259,N_34230,N_34210);
and U34260 (N_34260,N_34198,N_34155);
nor U34261 (N_34261,N_34235,N_34118);
nor U34262 (N_34262,N_34094,N_34164);
nand U34263 (N_34263,N_34219,N_34163);
and U34264 (N_34264,N_34132,N_34151);
nor U34265 (N_34265,N_34047,N_34113);
nor U34266 (N_34266,N_34220,N_34009);
xor U34267 (N_34267,N_34150,N_34143);
or U34268 (N_34268,N_34023,N_34153);
or U34269 (N_34269,N_34227,N_34195);
xor U34270 (N_34270,N_34244,N_34201);
nor U34271 (N_34271,N_34060,N_34127);
nor U34272 (N_34272,N_34142,N_34246);
and U34273 (N_34273,N_34145,N_34167);
and U34274 (N_34274,N_34225,N_34184);
or U34275 (N_34275,N_34099,N_34166);
nor U34276 (N_34276,N_34083,N_34096);
and U34277 (N_34277,N_34182,N_34134);
or U34278 (N_34278,N_34093,N_34079);
xnor U34279 (N_34279,N_34071,N_34139);
nor U34280 (N_34280,N_34076,N_34051);
nor U34281 (N_34281,N_34122,N_34156);
or U34282 (N_34282,N_34208,N_34125);
or U34283 (N_34283,N_34206,N_34234);
or U34284 (N_34284,N_34205,N_34175);
or U34285 (N_34285,N_34007,N_34039);
and U34286 (N_34286,N_34050,N_34199);
nand U34287 (N_34287,N_34106,N_34131);
or U34288 (N_34288,N_34067,N_34034);
and U34289 (N_34289,N_34077,N_34135);
nand U34290 (N_34290,N_34123,N_34136);
or U34291 (N_34291,N_34087,N_34028);
or U34292 (N_34292,N_34149,N_34006);
nand U34293 (N_34293,N_34124,N_34178);
and U34294 (N_34294,N_34186,N_34174);
or U34295 (N_34295,N_34098,N_34063);
nand U34296 (N_34296,N_34116,N_34168);
nor U34297 (N_34297,N_34044,N_34200);
nand U34298 (N_34298,N_34223,N_34226);
and U34299 (N_34299,N_34172,N_34229);
and U34300 (N_34300,N_34102,N_34045);
nor U34301 (N_34301,N_34085,N_34187);
or U34302 (N_34302,N_34148,N_34197);
and U34303 (N_34303,N_34231,N_34084);
xor U34304 (N_34304,N_34130,N_34126);
nand U34305 (N_34305,N_34075,N_34202);
or U34306 (N_34306,N_34032,N_34239);
xnor U34307 (N_34307,N_34066,N_34068);
or U34308 (N_34308,N_34017,N_34043);
nor U34309 (N_34309,N_34117,N_34176);
and U34310 (N_34310,N_34058,N_34000);
xor U34311 (N_34311,N_34042,N_34241);
or U34312 (N_34312,N_34086,N_34033);
nand U34313 (N_34313,N_34215,N_34104);
nand U34314 (N_34314,N_34004,N_34165);
or U34315 (N_34315,N_34052,N_34110);
and U34316 (N_34316,N_34185,N_34247);
xor U34317 (N_34317,N_34189,N_34192);
nand U34318 (N_34318,N_34237,N_34037);
or U34319 (N_34319,N_34245,N_34211);
nor U34320 (N_34320,N_34129,N_34055);
xnor U34321 (N_34321,N_34101,N_34091);
or U34322 (N_34322,N_34013,N_34062);
nor U34323 (N_34323,N_34181,N_34224);
nor U34324 (N_34324,N_34173,N_34190);
nand U34325 (N_34325,N_34152,N_34012);
nand U34326 (N_34326,N_34089,N_34238);
xor U34327 (N_34327,N_34141,N_34222);
xnor U34328 (N_34328,N_34020,N_34029);
xor U34329 (N_34329,N_34008,N_34217);
nand U34330 (N_34330,N_34090,N_34140);
nand U34331 (N_34331,N_34001,N_34196);
xor U34332 (N_34332,N_34081,N_34053);
xnor U34333 (N_34333,N_34002,N_34169);
and U34334 (N_34334,N_34105,N_34030);
and U34335 (N_34335,N_34137,N_34038);
xor U34336 (N_34336,N_34072,N_34183);
xnor U34337 (N_34337,N_34059,N_34111);
xnor U34338 (N_34338,N_34218,N_34147);
or U34339 (N_34339,N_34049,N_34016);
nand U34340 (N_34340,N_34103,N_34095);
nand U34341 (N_34341,N_34249,N_34041);
nand U34342 (N_34342,N_34203,N_34031);
and U34343 (N_34343,N_34221,N_34080);
nor U34344 (N_34344,N_34048,N_34170);
and U34345 (N_34345,N_34025,N_34232);
or U34346 (N_34346,N_34194,N_34161);
and U34347 (N_34347,N_34216,N_34022);
nand U34348 (N_34348,N_34119,N_34158);
nor U34349 (N_34349,N_34040,N_34191);
and U34350 (N_34350,N_34204,N_34107);
or U34351 (N_34351,N_34024,N_34162);
nand U34352 (N_34352,N_34138,N_34243);
and U34353 (N_34353,N_34027,N_34036);
nor U34354 (N_34354,N_34069,N_34019);
and U34355 (N_34355,N_34248,N_34121);
nand U34356 (N_34356,N_34082,N_34073);
or U34357 (N_34357,N_34015,N_34014);
xor U34358 (N_34358,N_34018,N_34159);
xnor U34359 (N_34359,N_34010,N_34233);
xor U34360 (N_34360,N_34133,N_34061);
and U34361 (N_34361,N_34088,N_34005);
xor U34362 (N_34362,N_34180,N_34109);
or U34363 (N_34363,N_34054,N_34171);
nor U34364 (N_34364,N_34092,N_34207);
nor U34365 (N_34365,N_34236,N_34115);
xnor U34366 (N_34366,N_34078,N_34179);
or U34367 (N_34367,N_34157,N_34070);
nand U34368 (N_34368,N_34240,N_34112);
or U34369 (N_34369,N_34193,N_34100);
and U34370 (N_34370,N_34146,N_34011);
nor U34371 (N_34371,N_34214,N_34154);
nand U34372 (N_34372,N_34056,N_34242);
nand U34373 (N_34373,N_34057,N_34026);
and U34374 (N_34374,N_34021,N_34228);
nand U34375 (N_34375,N_34172,N_34220);
xor U34376 (N_34376,N_34105,N_34045);
xnor U34377 (N_34377,N_34125,N_34127);
nand U34378 (N_34378,N_34134,N_34219);
nand U34379 (N_34379,N_34025,N_34040);
or U34380 (N_34380,N_34092,N_34168);
or U34381 (N_34381,N_34102,N_34233);
nor U34382 (N_34382,N_34004,N_34242);
nor U34383 (N_34383,N_34153,N_34077);
nand U34384 (N_34384,N_34000,N_34192);
nand U34385 (N_34385,N_34138,N_34125);
or U34386 (N_34386,N_34240,N_34017);
xor U34387 (N_34387,N_34044,N_34119);
nor U34388 (N_34388,N_34132,N_34018);
or U34389 (N_34389,N_34060,N_34074);
and U34390 (N_34390,N_34023,N_34092);
nor U34391 (N_34391,N_34183,N_34220);
nand U34392 (N_34392,N_34239,N_34104);
xnor U34393 (N_34393,N_34156,N_34128);
nor U34394 (N_34394,N_34109,N_34132);
or U34395 (N_34395,N_34113,N_34137);
nor U34396 (N_34396,N_34214,N_34061);
nand U34397 (N_34397,N_34199,N_34120);
nor U34398 (N_34398,N_34218,N_34045);
xnor U34399 (N_34399,N_34089,N_34023);
nand U34400 (N_34400,N_34247,N_34170);
nor U34401 (N_34401,N_34132,N_34240);
nor U34402 (N_34402,N_34064,N_34073);
nor U34403 (N_34403,N_34065,N_34070);
nor U34404 (N_34404,N_34227,N_34198);
and U34405 (N_34405,N_34240,N_34001);
or U34406 (N_34406,N_34143,N_34021);
and U34407 (N_34407,N_34050,N_34104);
and U34408 (N_34408,N_34120,N_34158);
nor U34409 (N_34409,N_34017,N_34112);
nor U34410 (N_34410,N_34065,N_34036);
xnor U34411 (N_34411,N_34226,N_34193);
and U34412 (N_34412,N_34211,N_34241);
nand U34413 (N_34413,N_34138,N_34242);
or U34414 (N_34414,N_34144,N_34145);
and U34415 (N_34415,N_34115,N_34179);
nor U34416 (N_34416,N_34236,N_34070);
xnor U34417 (N_34417,N_34085,N_34116);
or U34418 (N_34418,N_34159,N_34183);
nor U34419 (N_34419,N_34087,N_34217);
nand U34420 (N_34420,N_34044,N_34175);
xor U34421 (N_34421,N_34010,N_34012);
xnor U34422 (N_34422,N_34165,N_34153);
xor U34423 (N_34423,N_34105,N_34189);
xnor U34424 (N_34424,N_34135,N_34117);
nand U34425 (N_34425,N_34019,N_34234);
or U34426 (N_34426,N_34002,N_34243);
and U34427 (N_34427,N_34047,N_34152);
nor U34428 (N_34428,N_34204,N_34182);
and U34429 (N_34429,N_34248,N_34215);
and U34430 (N_34430,N_34246,N_34048);
nand U34431 (N_34431,N_34013,N_34129);
nor U34432 (N_34432,N_34241,N_34206);
and U34433 (N_34433,N_34054,N_34072);
xnor U34434 (N_34434,N_34039,N_34024);
or U34435 (N_34435,N_34203,N_34128);
and U34436 (N_34436,N_34122,N_34211);
xor U34437 (N_34437,N_34080,N_34010);
nor U34438 (N_34438,N_34044,N_34137);
and U34439 (N_34439,N_34012,N_34115);
nand U34440 (N_34440,N_34223,N_34033);
nand U34441 (N_34441,N_34031,N_34022);
and U34442 (N_34442,N_34239,N_34078);
nand U34443 (N_34443,N_34136,N_34092);
nand U34444 (N_34444,N_34238,N_34131);
nand U34445 (N_34445,N_34213,N_34192);
xor U34446 (N_34446,N_34078,N_34092);
and U34447 (N_34447,N_34058,N_34239);
or U34448 (N_34448,N_34178,N_34181);
nor U34449 (N_34449,N_34222,N_34026);
xnor U34450 (N_34450,N_34091,N_34204);
or U34451 (N_34451,N_34032,N_34052);
nor U34452 (N_34452,N_34107,N_34231);
or U34453 (N_34453,N_34236,N_34166);
nor U34454 (N_34454,N_34144,N_34167);
nand U34455 (N_34455,N_34169,N_34121);
nor U34456 (N_34456,N_34084,N_34148);
nand U34457 (N_34457,N_34140,N_34091);
nand U34458 (N_34458,N_34031,N_34061);
and U34459 (N_34459,N_34077,N_34152);
nor U34460 (N_34460,N_34151,N_34175);
xor U34461 (N_34461,N_34111,N_34148);
and U34462 (N_34462,N_34170,N_34033);
and U34463 (N_34463,N_34063,N_34020);
nor U34464 (N_34464,N_34213,N_34091);
xnor U34465 (N_34465,N_34169,N_34051);
and U34466 (N_34466,N_34203,N_34092);
nor U34467 (N_34467,N_34147,N_34015);
and U34468 (N_34468,N_34145,N_34081);
nor U34469 (N_34469,N_34009,N_34031);
xnor U34470 (N_34470,N_34004,N_34082);
and U34471 (N_34471,N_34103,N_34062);
xor U34472 (N_34472,N_34095,N_34048);
nor U34473 (N_34473,N_34033,N_34230);
nand U34474 (N_34474,N_34213,N_34212);
nand U34475 (N_34475,N_34073,N_34160);
nand U34476 (N_34476,N_34225,N_34180);
xor U34477 (N_34477,N_34198,N_34043);
xor U34478 (N_34478,N_34205,N_34158);
or U34479 (N_34479,N_34171,N_34206);
xnor U34480 (N_34480,N_34164,N_34122);
nand U34481 (N_34481,N_34044,N_34182);
nand U34482 (N_34482,N_34008,N_34169);
and U34483 (N_34483,N_34182,N_34170);
or U34484 (N_34484,N_34183,N_34226);
xor U34485 (N_34485,N_34212,N_34243);
xnor U34486 (N_34486,N_34234,N_34105);
and U34487 (N_34487,N_34238,N_34181);
nor U34488 (N_34488,N_34125,N_34134);
or U34489 (N_34489,N_34132,N_34220);
or U34490 (N_34490,N_34150,N_34108);
nand U34491 (N_34491,N_34237,N_34061);
and U34492 (N_34492,N_34092,N_34090);
or U34493 (N_34493,N_34161,N_34180);
and U34494 (N_34494,N_34070,N_34000);
nor U34495 (N_34495,N_34026,N_34194);
or U34496 (N_34496,N_34203,N_34115);
nand U34497 (N_34497,N_34068,N_34159);
or U34498 (N_34498,N_34114,N_34042);
or U34499 (N_34499,N_34124,N_34088);
nor U34500 (N_34500,N_34463,N_34293);
nand U34501 (N_34501,N_34400,N_34417);
and U34502 (N_34502,N_34260,N_34345);
or U34503 (N_34503,N_34268,N_34271);
and U34504 (N_34504,N_34428,N_34276);
xor U34505 (N_34505,N_34344,N_34437);
nand U34506 (N_34506,N_34342,N_34378);
and U34507 (N_34507,N_34315,N_34280);
xnor U34508 (N_34508,N_34384,N_34495);
or U34509 (N_34509,N_34311,N_34318);
or U34510 (N_34510,N_34429,N_34256);
nor U34511 (N_34511,N_34422,N_34261);
or U34512 (N_34512,N_34385,N_34478);
or U34513 (N_34513,N_34307,N_34432);
and U34514 (N_34514,N_34264,N_34454);
and U34515 (N_34515,N_34298,N_34372);
and U34516 (N_34516,N_34353,N_34259);
or U34517 (N_34517,N_34450,N_34380);
or U34518 (N_34518,N_34337,N_34425);
nor U34519 (N_34519,N_34263,N_34462);
or U34520 (N_34520,N_34424,N_34395);
nor U34521 (N_34521,N_34414,N_34363);
and U34522 (N_34522,N_34447,N_34274);
nand U34523 (N_34523,N_34273,N_34409);
nand U34524 (N_34524,N_34300,N_34396);
nand U34525 (N_34525,N_34309,N_34381);
and U34526 (N_34526,N_34379,N_34369);
xnor U34527 (N_34527,N_34481,N_34430);
or U34528 (N_34528,N_34418,N_34347);
or U34529 (N_34529,N_34442,N_34270);
nand U34530 (N_34530,N_34404,N_34482);
xnor U34531 (N_34531,N_34492,N_34496);
and U34532 (N_34532,N_34332,N_34446);
xor U34533 (N_34533,N_34489,N_34296);
or U34534 (N_34534,N_34316,N_34460);
nor U34535 (N_34535,N_34288,N_34279);
xnor U34536 (N_34536,N_34451,N_34403);
nor U34537 (N_34537,N_34359,N_34301);
and U34538 (N_34538,N_34408,N_34304);
nor U34539 (N_34539,N_34366,N_34367);
or U34540 (N_34540,N_34299,N_34443);
or U34541 (N_34541,N_34376,N_34453);
nand U34542 (N_34542,N_34470,N_34354);
nand U34543 (N_34543,N_34466,N_34329);
and U34544 (N_34544,N_34471,N_34253);
xnor U34545 (N_34545,N_34459,N_34421);
nor U34546 (N_34546,N_34440,N_34473);
nand U34547 (N_34547,N_34290,N_34281);
or U34548 (N_34548,N_34491,N_34386);
and U34549 (N_34549,N_34358,N_34383);
or U34550 (N_34550,N_34328,N_34339);
and U34551 (N_34551,N_34483,N_34258);
or U34552 (N_34552,N_34297,N_34444);
xor U34553 (N_34553,N_34475,N_34493);
and U34554 (N_34554,N_34278,N_34319);
or U34555 (N_34555,N_34340,N_34349);
nand U34556 (N_34556,N_34449,N_34388);
nor U34557 (N_34557,N_34302,N_34286);
and U34558 (N_34558,N_34357,N_34393);
nor U34559 (N_34559,N_34487,N_34368);
and U34560 (N_34560,N_34387,N_34490);
nand U34561 (N_34561,N_34295,N_34479);
nand U34562 (N_34562,N_34445,N_34448);
and U34563 (N_34563,N_34435,N_34306);
nand U34564 (N_34564,N_34391,N_34294);
or U34565 (N_34565,N_34333,N_34499);
and U34566 (N_34566,N_34269,N_34350);
nand U34567 (N_34567,N_34282,N_34255);
nand U34568 (N_34568,N_34360,N_34485);
xor U34569 (N_34569,N_34374,N_34257);
nand U34570 (N_34570,N_34251,N_34305);
or U34571 (N_34571,N_34474,N_34427);
and U34572 (N_34572,N_34335,N_34484);
or U34573 (N_34573,N_34284,N_34287);
and U34574 (N_34574,N_34252,N_34277);
nor U34575 (N_34575,N_34322,N_34285);
or U34576 (N_34576,N_34262,N_34476);
and U34577 (N_34577,N_34321,N_34406);
or U34578 (N_34578,N_34423,N_34402);
or U34579 (N_34579,N_34494,N_34438);
and U34580 (N_34580,N_34272,N_34331);
and U34581 (N_34581,N_34392,N_34289);
and U34582 (N_34582,N_34283,N_34434);
or U34583 (N_34583,N_34415,N_34313);
xnor U34584 (N_34584,N_34410,N_34413);
nand U34585 (N_34585,N_34426,N_34394);
and U34586 (N_34586,N_34364,N_34433);
xnor U34587 (N_34587,N_34265,N_34497);
xnor U34588 (N_34588,N_34389,N_34412);
or U34589 (N_34589,N_34320,N_34254);
and U34590 (N_34590,N_34275,N_34405);
nor U34591 (N_34591,N_34464,N_34292);
nand U34592 (N_34592,N_34330,N_34373);
nand U34593 (N_34593,N_34441,N_34407);
xor U34594 (N_34594,N_34377,N_34334);
nand U34595 (N_34595,N_34398,N_34390);
xor U34596 (N_34596,N_34362,N_34346);
and U34597 (N_34597,N_34326,N_34488);
nor U34598 (N_34598,N_34314,N_34397);
xnor U34599 (N_34599,N_34267,N_34312);
nor U34600 (N_34600,N_34465,N_34303);
and U34601 (N_34601,N_34310,N_34472);
or U34602 (N_34602,N_34401,N_34480);
or U34603 (N_34603,N_34375,N_34341);
nand U34604 (N_34604,N_34324,N_34457);
or U34605 (N_34605,N_34419,N_34371);
nor U34606 (N_34606,N_34436,N_34308);
nand U34607 (N_34607,N_34250,N_34323);
nand U34608 (N_34608,N_34317,N_34361);
or U34609 (N_34609,N_34431,N_34336);
nand U34610 (N_34610,N_34439,N_34382);
and U34611 (N_34611,N_34351,N_34469);
xnor U34612 (N_34612,N_34356,N_34468);
nor U34613 (N_34613,N_34365,N_34411);
nor U34614 (N_34614,N_34456,N_34467);
or U34615 (N_34615,N_34291,N_34486);
or U34616 (N_34616,N_34370,N_34498);
and U34617 (N_34617,N_34452,N_34348);
xnor U34618 (N_34618,N_34477,N_34338);
nand U34619 (N_34619,N_34343,N_34352);
nor U34620 (N_34620,N_34355,N_34399);
or U34621 (N_34621,N_34455,N_34416);
and U34622 (N_34622,N_34327,N_34266);
and U34623 (N_34623,N_34420,N_34458);
nor U34624 (N_34624,N_34461,N_34325);
or U34625 (N_34625,N_34410,N_34430);
or U34626 (N_34626,N_34461,N_34380);
and U34627 (N_34627,N_34397,N_34377);
nand U34628 (N_34628,N_34289,N_34368);
and U34629 (N_34629,N_34432,N_34352);
xnor U34630 (N_34630,N_34385,N_34395);
nand U34631 (N_34631,N_34256,N_34377);
or U34632 (N_34632,N_34348,N_34298);
nand U34633 (N_34633,N_34498,N_34351);
xnor U34634 (N_34634,N_34475,N_34441);
and U34635 (N_34635,N_34465,N_34262);
xnor U34636 (N_34636,N_34453,N_34257);
or U34637 (N_34637,N_34285,N_34418);
and U34638 (N_34638,N_34468,N_34310);
xnor U34639 (N_34639,N_34251,N_34307);
xor U34640 (N_34640,N_34285,N_34314);
or U34641 (N_34641,N_34479,N_34411);
and U34642 (N_34642,N_34418,N_34466);
nand U34643 (N_34643,N_34281,N_34447);
nand U34644 (N_34644,N_34432,N_34395);
nand U34645 (N_34645,N_34354,N_34366);
and U34646 (N_34646,N_34489,N_34304);
nor U34647 (N_34647,N_34389,N_34285);
or U34648 (N_34648,N_34262,N_34353);
xor U34649 (N_34649,N_34297,N_34299);
nand U34650 (N_34650,N_34397,N_34471);
xnor U34651 (N_34651,N_34295,N_34339);
nand U34652 (N_34652,N_34447,N_34308);
and U34653 (N_34653,N_34459,N_34335);
nand U34654 (N_34654,N_34349,N_34277);
and U34655 (N_34655,N_34267,N_34311);
nand U34656 (N_34656,N_34383,N_34290);
or U34657 (N_34657,N_34476,N_34254);
and U34658 (N_34658,N_34453,N_34342);
xor U34659 (N_34659,N_34358,N_34424);
and U34660 (N_34660,N_34461,N_34454);
nand U34661 (N_34661,N_34327,N_34463);
nand U34662 (N_34662,N_34323,N_34355);
nor U34663 (N_34663,N_34326,N_34484);
xor U34664 (N_34664,N_34440,N_34296);
nand U34665 (N_34665,N_34276,N_34498);
nor U34666 (N_34666,N_34478,N_34458);
or U34667 (N_34667,N_34486,N_34404);
nand U34668 (N_34668,N_34484,N_34377);
and U34669 (N_34669,N_34303,N_34459);
or U34670 (N_34670,N_34395,N_34402);
xnor U34671 (N_34671,N_34316,N_34337);
nand U34672 (N_34672,N_34404,N_34421);
and U34673 (N_34673,N_34448,N_34363);
and U34674 (N_34674,N_34268,N_34286);
or U34675 (N_34675,N_34479,N_34452);
and U34676 (N_34676,N_34435,N_34264);
and U34677 (N_34677,N_34371,N_34306);
nor U34678 (N_34678,N_34392,N_34297);
xor U34679 (N_34679,N_34412,N_34391);
and U34680 (N_34680,N_34470,N_34397);
nor U34681 (N_34681,N_34353,N_34477);
and U34682 (N_34682,N_34341,N_34369);
and U34683 (N_34683,N_34270,N_34481);
nor U34684 (N_34684,N_34384,N_34372);
and U34685 (N_34685,N_34372,N_34253);
or U34686 (N_34686,N_34376,N_34485);
and U34687 (N_34687,N_34421,N_34272);
xor U34688 (N_34688,N_34394,N_34489);
xor U34689 (N_34689,N_34336,N_34453);
nor U34690 (N_34690,N_34384,N_34299);
nand U34691 (N_34691,N_34373,N_34411);
nand U34692 (N_34692,N_34432,N_34365);
nand U34693 (N_34693,N_34266,N_34302);
and U34694 (N_34694,N_34470,N_34284);
nand U34695 (N_34695,N_34364,N_34463);
and U34696 (N_34696,N_34442,N_34388);
nand U34697 (N_34697,N_34287,N_34264);
nor U34698 (N_34698,N_34385,N_34490);
nand U34699 (N_34699,N_34365,N_34293);
xor U34700 (N_34700,N_34455,N_34397);
nor U34701 (N_34701,N_34289,N_34490);
xor U34702 (N_34702,N_34366,N_34421);
and U34703 (N_34703,N_34444,N_34315);
nor U34704 (N_34704,N_34343,N_34384);
xnor U34705 (N_34705,N_34388,N_34447);
and U34706 (N_34706,N_34399,N_34460);
xor U34707 (N_34707,N_34321,N_34405);
xor U34708 (N_34708,N_34493,N_34283);
nand U34709 (N_34709,N_34474,N_34302);
or U34710 (N_34710,N_34466,N_34370);
xor U34711 (N_34711,N_34396,N_34382);
nor U34712 (N_34712,N_34436,N_34362);
xor U34713 (N_34713,N_34330,N_34466);
or U34714 (N_34714,N_34477,N_34322);
and U34715 (N_34715,N_34280,N_34314);
nor U34716 (N_34716,N_34314,N_34490);
or U34717 (N_34717,N_34276,N_34435);
nor U34718 (N_34718,N_34401,N_34386);
and U34719 (N_34719,N_34459,N_34291);
or U34720 (N_34720,N_34400,N_34462);
xnor U34721 (N_34721,N_34355,N_34281);
nor U34722 (N_34722,N_34447,N_34483);
nor U34723 (N_34723,N_34420,N_34435);
or U34724 (N_34724,N_34354,N_34296);
nand U34725 (N_34725,N_34460,N_34309);
nand U34726 (N_34726,N_34456,N_34444);
and U34727 (N_34727,N_34291,N_34398);
nand U34728 (N_34728,N_34498,N_34387);
and U34729 (N_34729,N_34313,N_34421);
nand U34730 (N_34730,N_34375,N_34398);
nand U34731 (N_34731,N_34461,N_34471);
nor U34732 (N_34732,N_34300,N_34290);
nor U34733 (N_34733,N_34355,N_34364);
or U34734 (N_34734,N_34406,N_34444);
xnor U34735 (N_34735,N_34464,N_34462);
nor U34736 (N_34736,N_34444,N_34284);
and U34737 (N_34737,N_34273,N_34329);
nor U34738 (N_34738,N_34355,N_34383);
and U34739 (N_34739,N_34283,N_34260);
and U34740 (N_34740,N_34260,N_34288);
and U34741 (N_34741,N_34402,N_34456);
nor U34742 (N_34742,N_34264,N_34251);
nor U34743 (N_34743,N_34467,N_34258);
nand U34744 (N_34744,N_34343,N_34497);
nor U34745 (N_34745,N_34393,N_34378);
and U34746 (N_34746,N_34393,N_34404);
xnor U34747 (N_34747,N_34435,N_34254);
nor U34748 (N_34748,N_34363,N_34331);
and U34749 (N_34749,N_34393,N_34498);
xor U34750 (N_34750,N_34666,N_34664);
xor U34751 (N_34751,N_34571,N_34705);
nor U34752 (N_34752,N_34513,N_34656);
xnor U34753 (N_34753,N_34601,N_34665);
and U34754 (N_34754,N_34711,N_34519);
nor U34755 (N_34755,N_34611,N_34678);
nand U34756 (N_34756,N_34731,N_34539);
xor U34757 (N_34757,N_34604,N_34594);
or U34758 (N_34758,N_34749,N_34639);
or U34759 (N_34759,N_34680,N_34723);
nand U34760 (N_34760,N_34699,N_34581);
nand U34761 (N_34761,N_34582,N_34536);
or U34762 (N_34762,N_34575,N_34722);
nand U34763 (N_34763,N_34623,N_34561);
nor U34764 (N_34764,N_34620,N_34626);
or U34765 (N_34765,N_34634,N_34578);
nand U34766 (N_34766,N_34650,N_34653);
nand U34767 (N_34767,N_34606,N_34654);
nor U34768 (N_34768,N_34658,N_34500);
nand U34769 (N_34769,N_34533,N_34547);
and U34770 (N_34770,N_34735,N_34717);
nor U34771 (N_34771,N_34707,N_34511);
nand U34772 (N_34772,N_34538,N_34612);
xor U34773 (N_34773,N_34507,N_34599);
or U34774 (N_34774,N_34632,N_34745);
and U34775 (N_34775,N_34649,N_34591);
xor U34776 (N_34776,N_34543,N_34532);
xor U34777 (N_34777,N_34638,N_34588);
nor U34778 (N_34778,N_34747,N_34506);
xnor U34779 (N_34779,N_34583,N_34508);
and U34780 (N_34780,N_34744,N_34563);
nor U34781 (N_34781,N_34695,N_34660);
nor U34782 (N_34782,N_34509,N_34585);
or U34783 (N_34783,N_34577,N_34530);
nor U34784 (N_34784,N_34555,N_34694);
or U34785 (N_34785,N_34633,N_34684);
nor U34786 (N_34786,N_34527,N_34729);
nand U34787 (N_34787,N_34631,N_34554);
and U34788 (N_34788,N_34748,N_34551);
nand U34789 (N_34789,N_34702,N_34685);
nand U34790 (N_34790,N_34687,N_34505);
nor U34791 (N_34791,N_34728,N_34580);
nand U34792 (N_34792,N_34550,N_34710);
or U34793 (N_34793,N_34718,N_34697);
xnor U34794 (N_34794,N_34524,N_34537);
nand U34795 (N_34795,N_34616,N_34515);
and U34796 (N_34796,N_34574,N_34677);
and U34797 (N_34797,N_34609,N_34726);
or U34798 (N_34798,N_34641,N_34683);
or U34799 (N_34799,N_34607,N_34706);
xor U34800 (N_34800,N_34688,N_34739);
nand U34801 (N_34801,N_34682,N_34659);
and U34802 (N_34802,N_34572,N_34640);
xnor U34803 (N_34803,N_34647,N_34504);
and U34804 (N_34804,N_34635,N_34681);
xor U34805 (N_34805,N_34645,N_34686);
nor U34806 (N_34806,N_34624,N_34674);
nand U34807 (N_34807,N_34715,N_34534);
or U34808 (N_34808,N_34627,N_34737);
nor U34809 (N_34809,N_34557,N_34596);
nand U34810 (N_34810,N_34512,N_34546);
or U34811 (N_34811,N_34568,N_34614);
xor U34812 (N_34812,N_34503,N_34522);
or U34813 (N_34813,N_34714,N_34567);
or U34814 (N_34814,N_34712,N_34535);
and U34815 (N_34815,N_34592,N_34556);
xnor U34816 (N_34816,N_34548,N_34738);
xor U34817 (N_34817,N_34733,N_34618);
xor U34818 (N_34818,N_34671,N_34516);
and U34819 (N_34819,N_34720,N_34603);
nand U34820 (N_34820,N_34544,N_34713);
nand U34821 (N_34821,N_34740,N_34570);
and U34822 (N_34822,N_34617,N_34589);
and U34823 (N_34823,N_34502,N_34545);
and U34824 (N_34824,N_34630,N_34520);
nor U34825 (N_34825,N_34540,N_34719);
or U34826 (N_34826,N_34598,N_34562);
nand U34827 (N_34827,N_34689,N_34560);
nor U34828 (N_34828,N_34673,N_34622);
and U34829 (N_34829,N_34619,N_34730);
nand U34830 (N_34830,N_34741,N_34661);
xnor U34831 (N_34831,N_34724,N_34644);
nor U34832 (N_34832,N_34734,N_34595);
xor U34833 (N_34833,N_34700,N_34558);
nand U34834 (N_34834,N_34675,N_34746);
nor U34835 (N_34835,N_34668,N_34629);
or U34836 (N_34836,N_34549,N_34651);
or U34837 (N_34837,N_34663,N_34643);
xnor U34838 (N_34838,N_34667,N_34565);
and U34839 (N_34839,N_34662,N_34669);
and U34840 (N_34840,N_34691,N_34727);
nor U34841 (N_34841,N_34701,N_34721);
xnor U34842 (N_34842,N_34655,N_34742);
or U34843 (N_34843,N_34510,N_34566);
xor U34844 (N_34844,N_34579,N_34648);
nand U34845 (N_34845,N_34608,N_34716);
xor U34846 (N_34846,N_34693,N_34602);
nor U34847 (N_34847,N_34528,N_34698);
or U34848 (N_34848,N_34553,N_34559);
nand U34849 (N_34849,N_34610,N_34708);
nor U34850 (N_34850,N_34696,N_34517);
xor U34851 (N_34851,N_34736,N_34637);
nor U34852 (N_34852,N_34525,N_34672);
nor U34853 (N_34853,N_34732,N_34605);
xnor U34854 (N_34854,N_34514,N_34584);
nand U34855 (N_34855,N_34586,N_34652);
xor U34856 (N_34856,N_34590,N_34690);
and U34857 (N_34857,N_34615,N_34636);
nand U34858 (N_34858,N_34569,N_34704);
xor U34859 (N_34859,N_34518,N_34541);
xnor U34860 (N_34860,N_34521,N_34529);
or U34861 (N_34861,N_34597,N_34621);
nand U34862 (N_34862,N_34709,N_34743);
or U34863 (N_34863,N_34501,N_34628);
or U34864 (N_34864,N_34646,N_34573);
xnor U34865 (N_34865,N_34552,N_34523);
xor U34866 (N_34866,N_34593,N_34676);
xor U34867 (N_34867,N_34657,N_34587);
or U34868 (N_34868,N_34600,N_34725);
nor U34869 (N_34869,N_34679,N_34642);
nor U34870 (N_34870,N_34703,N_34564);
nor U34871 (N_34871,N_34625,N_34613);
nand U34872 (N_34872,N_34692,N_34531);
or U34873 (N_34873,N_34576,N_34542);
xnor U34874 (N_34874,N_34670,N_34526);
or U34875 (N_34875,N_34629,N_34700);
and U34876 (N_34876,N_34703,N_34708);
nand U34877 (N_34877,N_34681,N_34592);
nor U34878 (N_34878,N_34568,N_34684);
nand U34879 (N_34879,N_34570,N_34503);
or U34880 (N_34880,N_34651,N_34735);
xor U34881 (N_34881,N_34565,N_34701);
and U34882 (N_34882,N_34626,N_34511);
nor U34883 (N_34883,N_34602,N_34744);
and U34884 (N_34884,N_34705,N_34724);
nor U34885 (N_34885,N_34531,N_34656);
nor U34886 (N_34886,N_34638,N_34742);
xnor U34887 (N_34887,N_34714,N_34639);
nand U34888 (N_34888,N_34680,N_34562);
or U34889 (N_34889,N_34525,N_34660);
nand U34890 (N_34890,N_34601,N_34644);
nor U34891 (N_34891,N_34696,N_34726);
nand U34892 (N_34892,N_34500,N_34596);
and U34893 (N_34893,N_34710,N_34622);
nand U34894 (N_34894,N_34662,N_34523);
or U34895 (N_34895,N_34597,N_34559);
nand U34896 (N_34896,N_34693,N_34656);
nor U34897 (N_34897,N_34601,N_34742);
and U34898 (N_34898,N_34504,N_34513);
and U34899 (N_34899,N_34561,N_34626);
and U34900 (N_34900,N_34707,N_34528);
or U34901 (N_34901,N_34614,N_34691);
nor U34902 (N_34902,N_34593,N_34614);
or U34903 (N_34903,N_34722,N_34509);
nand U34904 (N_34904,N_34703,N_34697);
or U34905 (N_34905,N_34696,N_34741);
and U34906 (N_34906,N_34597,N_34521);
and U34907 (N_34907,N_34718,N_34705);
nor U34908 (N_34908,N_34644,N_34614);
xnor U34909 (N_34909,N_34581,N_34664);
nor U34910 (N_34910,N_34620,N_34584);
nand U34911 (N_34911,N_34732,N_34648);
nand U34912 (N_34912,N_34596,N_34617);
or U34913 (N_34913,N_34568,N_34600);
and U34914 (N_34914,N_34672,N_34557);
nor U34915 (N_34915,N_34536,N_34624);
and U34916 (N_34916,N_34610,N_34677);
or U34917 (N_34917,N_34549,N_34626);
or U34918 (N_34918,N_34741,N_34557);
nand U34919 (N_34919,N_34505,N_34580);
or U34920 (N_34920,N_34736,N_34669);
and U34921 (N_34921,N_34589,N_34744);
or U34922 (N_34922,N_34731,N_34664);
xor U34923 (N_34923,N_34590,N_34539);
nor U34924 (N_34924,N_34554,N_34569);
or U34925 (N_34925,N_34549,N_34563);
xor U34926 (N_34926,N_34735,N_34670);
or U34927 (N_34927,N_34600,N_34732);
xor U34928 (N_34928,N_34551,N_34529);
nor U34929 (N_34929,N_34693,N_34592);
xor U34930 (N_34930,N_34538,N_34593);
and U34931 (N_34931,N_34643,N_34521);
nor U34932 (N_34932,N_34562,N_34557);
or U34933 (N_34933,N_34549,N_34681);
and U34934 (N_34934,N_34525,N_34675);
nor U34935 (N_34935,N_34670,N_34698);
and U34936 (N_34936,N_34516,N_34661);
xor U34937 (N_34937,N_34654,N_34520);
or U34938 (N_34938,N_34670,N_34618);
or U34939 (N_34939,N_34507,N_34747);
or U34940 (N_34940,N_34688,N_34699);
or U34941 (N_34941,N_34525,N_34530);
or U34942 (N_34942,N_34525,N_34506);
or U34943 (N_34943,N_34616,N_34714);
or U34944 (N_34944,N_34695,N_34519);
and U34945 (N_34945,N_34637,N_34720);
and U34946 (N_34946,N_34648,N_34516);
and U34947 (N_34947,N_34575,N_34661);
nand U34948 (N_34948,N_34567,N_34663);
or U34949 (N_34949,N_34658,N_34593);
nor U34950 (N_34950,N_34687,N_34644);
xor U34951 (N_34951,N_34623,N_34581);
xnor U34952 (N_34952,N_34746,N_34576);
and U34953 (N_34953,N_34634,N_34549);
and U34954 (N_34954,N_34589,N_34514);
nor U34955 (N_34955,N_34526,N_34627);
and U34956 (N_34956,N_34656,N_34588);
nor U34957 (N_34957,N_34645,N_34512);
nand U34958 (N_34958,N_34530,N_34745);
xnor U34959 (N_34959,N_34695,N_34710);
nand U34960 (N_34960,N_34554,N_34728);
and U34961 (N_34961,N_34664,N_34551);
and U34962 (N_34962,N_34708,N_34738);
and U34963 (N_34963,N_34715,N_34512);
and U34964 (N_34964,N_34651,N_34545);
nand U34965 (N_34965,N_34591,N_34575);
xnor U34966 (N_34966,N_34618,N_34589);
nor U34967 (N_34967,N_34719,N_34661);
or U34968 (N_34968,N_34746,N_34522);
and U34969 (N_34969,N_34576,N_34521);
or U34970 (N_34970,N_34579,N_34676);
nor U34971 (N_34971,N_34663,N_34527);
nor U34972 (N_34972,N_34510,N_34586);
or U34973 (N_34973,N_34504,N_34638);
nand U34974 (N_34974,N_34559,N_34598);
and U34975 (N_34975,N_34514,N_34612);
nor U34976 (N_34976,N_34699,N_34658);
or U34977 (N_34977,N_34511,N_34561);
nor U34978 (N_34978,N_34669,N_34609);
xor U34979 (N_34979,N_34516,N_34529);
nand U34980 (N_34980,N_34628,N_34682);
and U34981 (N_34981,N_34542,N_34605);
xnor U34982 (N_34982,N_34642,N_34669);
nand U34983 (N_34983,N_34749,N_34703);
and U34984 (N_34984,N_34737,N_34631);
nand U34985 (N_34985,N_34613,N_34722);
and U34986 (N_34986,N_34648,N_34696);
nor U34987 (N_34987,N_34500,N_34621);
or U34988 (N_34988,N_34520,N_34606);
xor U34989 (N_34989,N_34717,N_34739);
nor U34990 (N_34990,N_34738,N_34652);
nor U34991 (N_34991,N_34621,N_34737);
nor U34992 (N_34992,N_34582,N_34690);
xor U34993 (N_34993,N_34662,N_34712);
and U34994 (N_34994,N_34612,N_34579);
and U34995 (N_34995,N_34724,N_34565);
xor U34996 (N_34996,N_34657,N_34580);
xnor U34997 (N_34997,N_34561,N_34600);
nand U34998 (N_34998,N_34742,N_34526);
and U34999 (N_34999,N_34573,N_34578);
nand U35000 (N_35000,N_34855,N_34793);
nor U35001 (N_35001,N_34851,N_34905);
and U35002 (N_35002,N_34760,N_34956);
nand U35003 (N_35003,N_34824,N_34904);
xor U35004 (N_35004,N_34900,N_34960);
nor U35005 (N_35005,N_34856,N_34970);
nor U35006 (N_35006,N_34854,N_34850);
and U35007 (N_35007,N_34944,N_34898);
xor U35008 (N_35008,N_34769,N_34958);
xnor U35009 (N_35009,N_34835,N_34811);
nand U35010 (N_35010,N_34826,N_34876);
and U35011 (N_35011,N_34801,N_34772);
nand U35012 (N_35012,N_34788,N_34830);
nand U35013 (N_35013,N_34996,N_34800);
xor U35014 (N_35014,N_34833,N_34950);
and U35015 (N_35015,N_34763,N_34984);
xnor U35016 (N_35016,N_34980,N_34959);
nand U35017 (N_35017,N_34778,N_34815);
or U35018 (N_35018,N_34822,N_34864);
xnor U35019 (N_35019,N_34859,N_34818);
nor U35020 (N_35020,N_34852,N_34917);
nand U35021 (N_35021,N_34899,N_34813);
xnor U35022 (N_35022,N_34922,N_34988);
or U35023 (N_35023,N_34911,N_34909);
xor U35024 (N_35024,N_34873,N_34979);
or U35025 (N_35025,N_34957,N_34761);
nor U35026 (N_35026,N_34963,N_34771);
or U35027 (N_35027,N_34969,N_34974);
or U35028 (N_35028,N_34783,N_34762);
nor U35029 (N_35029,N_34947,N_34910);
xor U35030 (N_35030,N_34918,N_34775);
or U35031 (N_35031,N_34878,N_34983);
and U35032 (N_35032,N_34895,N_34903);
nor U35033 (N_35033,N_34759,N_34894);
xor U35034 (N_35034,N_34828,N_34923);
or U35035 (N_35035,N_34782,N_34861);
and U35036 (N_35036,N_34934,N_34990);
and U35037 (N_35037,N_34972,N_34848);
nand U35038 (N_35038,N_34886,N_34884);
xnor U35039 (N_35039,N_34966,N_34953);
nand U35040 (N_35040,N_34827,N_34912);
nand U35041 (N_35041,N_34916,N_34942);
nor U35042 (N_35042,N_34929,N_34949);
nor U35043 (N_35043,N_34755,N_34882);
or U35044 (N_35044,N_34915,N_34844);
or U35045 (N_35045,N_34885,N_34802);
nand U35046 (N_35046,N_34840,N_34932);
xnor U35047 (N_35047,N_34770,N_34773);
nor U35048 (N_35048,N_34794,N_34820);
nor U35049 (N_35049,N_34881,N_34816);
xor U35050 (N_35050,N_34753,N_34943);
xnor U35051 (N_35051,N_34893,N_34868);
nand U35052 (N_35052,N_34857,N_34807);
or U35053 (N_35053,N_34875,N_34921);
xnor U35054 (N_35054,N_34831,N_34757);
nand U35055 (N_35055,N_34751,N_34987);
or U35056 (N_35056,N_34780,N_34926);
nor U35057 (N_35057,N_34823,N_34936);
or U35058 (N_35058,N_34791,N_34964);
and U35059 (N_35059,N_34941,N_34940);
or U35060 (N_35060,N_34986,N_34797);
nor U35061 (N_35061,N_34862,N_34896);
and U35062 (N_35062,N_34999,N_34821);
nor U35063 (N_35063,N_34869,N_34892);
nand U35064 (N_35064,N_34790,N_34832);
and U35065 (N_35065,N_34995,N_34784);
xor U35066 (N_35066,N_34781,N_34786);
or U35067 (N_35067,N_34845,N_34982);
xnor U35068 (N_35068,N_34955,N_34925);
nor U35069 (N_35069,N_34798,N_34973);
xnor U35070 (N_35070,N_34808,N_34937);
nand U35071 (N_35071,N_34887,N_34870);
xnor U35072 (N_35072,N_34817,N_34795);
xor U35073 (N_35073,N_34805,N_34866);
and U35074 (N_35074,N_34906,N_34946);
nor U35075 (N_35075,N_34834,N_34752);
and U35076 (N_35076,N_34927,N_34779);
and U35077 (N_35077,N_34841,N_34931);
or U35078 (N_35078,N_34825,N_34994);
xor U35079 (N_35079,N_34858,N_34992);
and U35080 (N_35080,N_34810,N_34948);
xnor U35081 (N_35081,N_34819,N_34812);
and U35082 (N_35082,N_34928,N_34939);
or U35083 (N_35083,N_34890,N_34765);
nand U35084 (N_35084,N_34938,N_34768);
xor U35085 (N_35085,N_34806,N_34754);
and U35086 (N_35086,N_34907,N_34897);
and U35087 (N_35087,N_34872,N_34766);
nor U35088 (N_35088,N_34993,N_34814);
nor U35089 (N_35089,N_34977,N_34968);
and U35090 (N_35090,N_34976,N_34991);
nor U35091 (N_35091,N_34924,N_34838);
or U35092 (N_35092,N_34774,N_34933);
nand U35093 (N_35093,N_34920,N_34837);
nor U35094 (N_35094,N_34776,N_34961);
or U35095 (N_35095,N_34792,N_34945);
nand U35096 (N_35096,N_34930,N_34750);
xnor U35097 (N_35097,N_34971,N_34997);
or U35098 (N_35098,N_34799,N_34901);
nor U35099 (N_35099,N_34985,N_34981);
or U35100 (N_35100,N_34975,N_34871);
xnor U35101 (N_35101,N_34785,N_34846);
nand U35102 (N_35102,N_34935,N_34954);
or U35103 (N_35103,N_34860,N_34839);
xor U35104 (N_35104,N_34804,N_34847);
or U35105 (N_35105,N_34874,N_34998);
nand U35106 (N_35106,N_34888,N_34758);
or U35107 (N_35107,N_34836,N_34789);
and U35108 (N_35108,N_34889,N_34809);
nand U35109 (N_35109,N_34919,N_34849);
nand U35110 (N_35110,N_34865,N_34880);
nor U35111 (N_35111,N_34803,N_34796);
nand U35112 (N_35112,N_34853,N_34877);
nand U35113 (N_35113,N_34914,N_34843);
or U35114 (N_35114,N_34978,N_34883);
nor U35115 (N_35115,N_34913,N_34891);
xor U35116 (N_35116,N_34756,N_34777);
nor U35117 (N_35117,N_34863,N_34879);
and U35118 (N_35118,N_34787,N_34967);
or U35119 (N_35119,N_34829,N_34767);
nor U35120 (N_35120,N_34764,N_34867);
or U35121 (N_35121,N_34962,N_34952);
or U35122 (N_35122,N_34951,N_34908);
xnor U35123 (N_35123,N_34965,N_34902);
nand U35124 (N_35124,N_34842,N_34989);
and U35125 (N_35125,N_34812,N_34954);
or U35126 (N_35126,N_34840,N_34835);
nand U35127 (N_35127,N_34879,N_34988);
nand U35128 (N_35128,N_34785,N_34760);
nor U35129 (N_35129,N_34793,N_34866);
nand U35130 (N_35130,N_34935,N_34893);
nor U35131 (N_35131,N_34946,N_34968);
and U35132 (N_35132,N_34821,N_34993);
xor U35133 (N_35133,N_34940,N_34763);
xnor U35134 (N_35134,N_34769,N_34984);
nand U35135 (N_35135,N_34809,N_34870);
xnor U35136 (N_35136,N_34762,N_34832);
nand U35137 (N_35137,N_34769,N_34875);
xor U35138 (N_35138,N_34959,N_34810);
nor U35139 (N_35139,N_34796,N_34952);
or U35140 (N_35140,N_34872,N_34891);
or U35141 (N_35141,N_34889,N_34963);
nor U35142 (N_35142,N_34863,N_34990);
nor U35143 (N_35143,N_34780,N_34985);
or U35144 (N_35144,N_34940,N_34849);
and U35145 (N_35145,N_34852,N_34976);
nand U35146 (N_35146,N_34865,N_34981);
or U35147 (N_35147,N_34790,N_34912);
and U35148 (N_35148,N_34802,N_34751);
xnor U35149 (N_35149,N_34950,N_34871);
nor U35150 (N_35150,N_34962,N_34837);
and U35151 (N_35151,N_34906,N_34767);
or U35152 (N_35152,N_34849,N_34841);
and U35153 (N_35153,N_34981,N_34782);
nand U35154 (N_35154,N_34940,N_34790);
nor U35155 (N_35155,N_34958,N_34910);
or U35156 (N_35156,N_34959,N_34752);
and U35157 (N_35157,N_34774,N_34912);
or U35158 (N_35158,N_34870,N_34865);
xor U35159 (N_35159,N_34854,N_34900);
nor U35160 (N_35160,N_34822,N_34890);
nor U35161 (N_35161,N_34813,N_34956);
xnor U35162 (N_35162,N_34756,N_34927);
xnor U35163 (N_35163,N_34832,N_34769);
or U35164 (N_35164,N_34936,N_34956);
nor U35165 (N_35165,N_34931,N_34960);
nand U35166 (N_35166,N_34875,N_34937);
or U35167 (N_35167,N_34871,N_34909);
or U35168 (N_35168,N_34798,N_34914);
xnor U35169 (N_35169,N_34871,N_34832);
xnor U35170 (N_35170,N_34778,N_34944);
nand U35171 (N_35171,N_34985,N_34917);
nand U35172 (N_35172,N_34949,N_34992);
nand U35173 (N_35173,N_34926,N_34865);
xnor U35174 (N_35174,N_34995,N_34807);
or U35175 (N_35175,N_34929,N_34782);
nand U35176 (N_35176,N_34826,N_34855);
or U35177 (N_35177,N_34851,N_34776);
nor U35178 (N_35178,N_34808,N_34959);
and U35179 (N_35179,N_34854,N_34812);
or U35180 (N_35180,N_34820,N_34951);
nand U35181 (N_35181,N_34800,N_34884);
and U35182 (N_35182,N_34996,N_34874);
nand U35183 (N_35183,N_34905,N_34820);
and U35184 (N_35184,N_34904,N_34892);
nor U35185 (N_35185,N_34878,N_34925);
nand U35186 (N_35186,N_34880,N_34820);
or U35187 (N_35187,N_34792,N_34941);
and U35188 (N_35188,N_34941,N_34795);
nor U35189 (N_35189,N_34923,N_34902);
xnor U35190 (N_35190,N_34997,N_34802);
and U35191 (N_35191,N_34851,N_34945);
nor U35192 (N_35192,N_34840,N_34787);
or U35193 (N_35193,N_34858,N_34789);
or U35194 (N_35194,N_34968,N_34910);
or U35195 (N_35195,N_34845,N_34896);
or U35196 (N_35196,N_34892,N_34927);
nand U35197 (N_35197,N_34903,N_34965);
nor U35198 (N_35198,N_34945,N_34938);
nand U35199 (N_35199,N_34886,N_34824);
nand U35200 (N_35200,N_34769,N_34793);
or U35201 (N_35201,N_34955,N_34824);
and U35202 (N_35202,N_34814,N_34927);
and U35203 (N_35203,N_34995,N_34933);
or U35204 (N_35204,N_34783,N_34909);
nand U35205 (N_35205,N_34846,N_34914);
xor U35206 (N_35206,N_34929,N_34993);
nand U35207 (N_35207,N_34849,N_34971);
and U35208 (N_35208,N_34864,N_34902);
and U35209 (N_35209,N_34920,N_34759);
xor U35210 (N_35210,N_34798,N_34931);
xor U35211 (N_35211,N_34793,N_34871);
or U35212 (N_35212,N_34957,N_34804);
xor U35213 (N_35213,N_34826,N_34844);
nor U35214 (N_35214,N_34774,N_34775);
nor U35215 (N_35215,N_34900,N_34987);
or U35216 (N_35216,N_34778,N_34905);
nor U35217 (N_35217,N_34872,N_34969);
nor U35218 (N_35218,N_34800,N_34753);
nand U35219 (N_35219,N_34992,N_34869);
and U35220 (N_35220,N_34998,N_34906);
or U35221 (N_35221,N_34972,N_34880);
and U35222 (N_35222,N_34777,N_34906);
nand U35223 (N_35223,N_34941,N_34878);
nand U35224 (N_35224,N_34938,N_34778);
nor U35225 (N_35225,N_34987,N_34879);
and U35226 (N_35226,N_34792,N_34949);
xnor U35227 (N_35227,N_34954,N_34947);
or U35228 (N_35228,N_34753,N_34759);
and U35229 (N_35229,N_34946,N_34985);
nand U35230 (N_35230,N_34809,N_34880);
xor U35231 (N_35231,N_34815,N_34832);
nor U35232 (N_35232,N_34806,N_34885);
xor U35233 (N_35233,N_34785,N_34823);
nor U35234 (N_35234,N_34917,N_34812);
nand U35235 (N_35235,N_34767,N_34921);
nand U35236 (N_35236,N_34854,N_34861);
or U35237 (N_35237,N_34911,N_34774);
or U35238 (N_35238,N_34949,N_34845);
or U35239 (N_35239,N_34997,N_34963);
or U35240 (N_35240,N_34832,N_34932);
nand U35241 (N_35241,N_34894,N_34996);
and U35242 (N_35242,N_34898,N_34781);
or U35243 (N_35243,N_34921,N_34759);
nand U35244 (N_35244,N_34820,N_34989);
xor U35245 (N_35245,N_34932,N_34907);
nor U35246 (N_35246,N_34934,N_34967);
or U35247 (N_35247,N_34823,N_34857);
or U35248 (N_35248,N_34768,N_34890);
and U35249 (N_35249,N_34995,N_34814);
xnor U35250 (N_35250,N_35082,N_35007);
and U35251 (N_35251,N_35106,N_35225);
and U35252 (N_35252,N_35046,N_35170);
nor U35253 (N_35253,N_35075,N_35044);
or U35254 (N_35254,N_35195,N_35206);
nor U35255 (N_35255,N_35148,N_35053);
and U35256 (N_35256,N_35030,N_35086);
and U35257 (N_35257,N_35192,N_35061);
nor U35258 (N_35258,N_35015,N_35246);
nand U35259 (N_35259,N_35085,N_35240);
or U35260 (N_35260,N_35114,N_35071);
and U35261 (N_35261,N_35076,N_35105);
or U35262 (N_35262,N_35109,N_35167);
and U35263 (N_35263,N_35131,N_35163);
nand U35264 (N_35264,N_35247,N_35023);
or U35265 (N_35265,N_35237,N_35037);
and U35266 (N_35266,N_35222,N_35204);
xnor U35267 (N_35267,N_35201,N_35129);
xor U35268 (N_35268,N_35039,N_35099);
or U35269 (N_35269,N_35056,N_35115);
or U35270 (N_35270,N_35002,N_35124);
xnor U35271 (N_35271,N_35134,N_35233);
or U35272 (N_35272,N_35213,N_35097);
nand U35273 (N_35273,N_35108,N_35009);
and U35274 (N_35274,N_35171,N_35040);
and U35275 (N_35275,N_35162,N_35184);
nand U35276 (N_35276,N_35178,N_35060);
nor U35277 (N_35277,N_35014,N_35197);
xor U35278 (N_35278,N_35054,N_35215);
and U35279 (N_35279,N_35051,N_35140);
and U35280 (N_35280,N_35059,N_35057);
nand U35281 (N_35281,N_35234,N_35083);
and U35282 (N_35282,N_35216,N_35136);
nor U35283 (N_35283,N_35066,N_35187);
and U35284 (N_35284,N_35118,N_35226);
or U35285 (N_35285,N_35239,N_35000);
and U35286 (N_35286,N_35011,N_35149);
or U35287 (N_35287,N_35169,N_35006);
nor U35288 (N_35288,N_35073,N_35160);
xor U35289 (N_35289,N_35021,N_35048);
xor U35290 (N_35290,N_35022,N_35205);
nand U35291 (N_35291,N_35005,N_35123);
or U35292 (N_35292,N_35091,N_35089);
and U35293 (N_35293,N_35209,N_35119);
nor U35294 (N_35294,N_35227,N_35135);
or U35295 (N_35295,N_35094,N_35219);
and U35296 (N_35296,N_35102,N_35095);
nand U35297 (N_35297,N_35043,N_35034);
xnor U35298 (N_35298,N_35045,N_35103);
nor U35299 (N_35299,N_35027,N_35231);
or U35300 (N_35300,N_35036,N_35024);
and U35301 (N_35301,N_35152,N_35088);
nand U35302 (N_35302,N_35138,N_35228);
nand U35303 (N_35303,N_35223,N_35245);
and U35304 (N_35304,N_35230,N_35087);
or U35305 (N_35305,N_35025,N_35132);
nand U35306 (N_35306,N_35202,N_35133);
xnor U35307 (N_35307,N_35067,N_35010);
xor U35308 (N_35308,N_35074,N_35012);
xor U35309 (N_35309,N_35249,N_35093);
or U35310 (N_35310,N_35125,N_35190);
or U35311 (N_35311,N_35026,N_35098);
nor U35312 (N_35312,N_35235,N_35144);
nand U35313 (N_35313,N_35180,N_35236);
and U35314 (N_35314,N_35181,N_35052);
and U35315 (N_35315,N_35092,N_35191);
nand U35316 (N_35316,N_35154,N_35101);
nor U35317 (N_35317,N_35084,N_35153);
nand U35318 (N_35318,N_35156,N_35242);
nand U35319 (N_35319,N_35185,N_35035);
and U35320 (N_35320,N_35165,N_35243);
xor U35321 (N_35321,N_35127,N_35121);
or U35322 (N_35322,N_35017,N_35207);
xor U35323 (N_35323,N_35161,N_35186);
and U35324 (N_35324,N_35173,N_35199);
xnor U35325 (N_35325,N_35116,N_35200);
xnor U35326 (N_35326,N_35218,N_35068);
nand U35327 (N_35327,N_35177,N_35155);
nand U35328 (N_35328,N_35244,N_35077);
or U35329 (N_35329,N_35238,N_35117);
xnor U35330 (N_35330,N_35078,N_35072);
nor U35331 (N_35331,N_35016,N_35220);
xnor U35332 (N_35332,N_35176,N_35122);
nand U35333 (N_35333,N_35164,N_35157);
xnor U35334 (N_35334,N_35189,N_35113);
or U35335 (N_35335,N_35158,N_35179);
nor U35336 (N_35336,N_35018,N_35159);
xnor U35337 (N_35337,N_35062,N_35174);
and U35338 (N_35338,N_35055,N_35110);
nor U35339 (N_35339,N_35100,N_35150);
nor U35340 (N_35340,N_35193,N_35019);
and U35341 (N_35341,N_35065,N_35241);
or U35342 (N_35342,N_35001,N_35188);
and U35343 (N_35343,N_35194,N_35080);
nand U35344 (N_35344,N_35137,N_35013);
and U35345 (N_35345,N_35146,N_35111);
xor U35346 (N_35346,N_35064,N_35151);
nand U35347 (N_35347,N_35031,N_35079);
nand U35348 (N_35348,N_35112,N_35143);
and U35349 (N_35349,N_35248,N_35050);
or U35350 (N_35350,N_35211,N_35120);
and U35351 (N_35351,N_35020,N_35203);
nand U35352 (N_35352,N_35008,N_35032);
xnor U35353 (N_35353,N_35217,N_35081);
nand U35354 (N_35354,N_35063,N_35198);
nand U35355 (N_35355,N_35214,N_35104);
or U35356 (N_35356,N_35130,N_35196);
xnor U35357 (N_35357,N_35172,N_35128);
xor U35358 (N_35358,N_35232,N_35208);
nor U35359 (N_35359,N_35182,N_35126);
or U35360 (N_35360,N_35229,N_35090);
xor U35361 (N_35361,N_35212,N_35042);
xor U35362 (N_35362,N_35139,N_35004);
xor U35363 (N_35363,N_35145,N_35224);
and U35364 (N_35364,N_35107,N_35058);
xor U35365 (N_35365,N_35028,N_35047);
nor U35366 (N_35366,N_35142,N_35141);
nor U35367 (N_35367,N_35003,N_35183);
nor U35368 (N_35368,N_35168,N_35029);
xor U35369 (N_35369,N_35038,N_35069);
nor U35370 (N_35370,N_35041,N_35049);
nand U35371 (N_35371,N_35096,N_35070);
and U35372 (N_35372,N_35147,N_35175);
or U35373 (N_35373,N_35210,N_35166);
and U35374 (N_35374,N_35221,N_35033);
nor U35375 (N_35375,N_35211,N_35128);
nand U35376 (N_35376,N_35211,N_35230);
nor U35377 (N_35377,N_35058,N_35103);
xor U35378 (N_35378,N_35171,N_35152);
and U35379 (N_35379,N_35104,N_35181);
or U35380 (N_35380,N_35092,N_35185);
xnor U35381 (N_35381,N_35085,N_35051);
nor U35382 (N_35382,N_35182,N_35067);
nor U35383 (N_35383,N_35034,N_35219);
and U35384 (N_35384,N_35248,N_35121);
nor U35385 (N_35385,N_35130,N_35110);
nor U35386 (N_35386,N_35236,N_35029);
or U35387 (N_35387,N_35073,N_35167);
nor U35388 (N_35388,N_35062,N_35221);
nand U35389 (N_35389,N_35068,N_35063);
or U35390 (N_35390,N_35101,N_35064);
or U35391 (N_35391,N_35238,N_35094);
nand U35392 (N_35392,N_35162,N_35088);
nand U35393 (N_35393,N_35050,N_35220);
or U35394 (N_35394,N_35219,N_35028);
nor U35395 (N_35395,N_35089,N_35236);
xnor U35396 (N_35396,N_35178,N_35048);
xnor U35397 (N_35397,N_35115,N_35154);
and U35398 (N_35398,N_35245,N_35124);
or U35399 (N_35399,N_35206,N_35130);
nand U35400 (N_35400,N_35058,N_35130);
and U35401 (N_35401,N_35071,N_35038);
nand U35402 (N_35402,N_35226,N_35047);
or U35403 (N_35403,N_35053,N_35095);
xor U35404 (N_35404,N_35059,N_35167);
nor U35405 (N_35405,N_35170,N_35136);
and U35406 (N_35406,N_35066,N_35071);
or U35407 (N_35407,N_35180,N_35116);
and U35408 (N_35408,N_35068,N_35240);
nor U35409 (N_35409,N_35143,N_35220);
nand U35410 (N_35410,N_35111,N_35181);
nand U35411 (N_35411,N_35060,N_35243);
nand U35412 (N_35412,N_35147,N_35218);
nand U35413 (N_35413,N_35143,N_35170);
xor U35414 (N_35414,N_35182,N_35234);
xnor U35415 (N_35415,N_35027,N_35148);
or U35416 (N_35416,N_35232,N_35121);
nor U35417 (N_35417,N_35014,N_35077);
and U35418 (N_35418,N_35182,N_35043);
nor U35419 (N_35419,N_35023,N_35112);
xnor U35420 (N_35420,N_35141,N_35198);
nand U35421 (N_35421,N_35073,N_35157);
nand U35422 (N_35422,N_35205,N_35075);
or U35423 (N_35423,N_35206,N_35000);
nor U35424 (N_35424,N_35108,N_35002);
nand U35425 (N_35425,N_35146,N_35033);
xnor U35426 (N_35426,N_35110,N_35119);
nand U35427 (N_35427,N_35158,N_35045);
nand U35428 (N_35428,N_35097,N_35208);
or U35429 (N_35429,N_35168,N_35004);
nand U35430 (N_35430,N_35033,N_35222);
nand U35431 (N_35431,N_35088,N_35180);
nand U35432 (N_35432,N_35070,N_35246);
nor U35433 (N_35433,N_35210,N_35046);
and U35434 (N_35434,N_35195,N_35201);
or U35435 (N_35435,N_35207,N_35000);
and U35436 (N_35436,N_35099,N_35068);
or U35437 (N_35437,N_35033,N_35171);
nand U35438 (N_35438,N_35044,N_35066);
xnor U35439 (N_35439,N_35171,N_35032);
and U35440 (N_35440,N_35064,N_35004);
nand U35441 (N_35441,N_35214,N_35191);
nor U35442 (N_35442,N_35142,N_35037);
nand U35443 (N_35443,N_35025,N_35123);
or U35444 (N_35444,N_35027,N_35003);
nor U35445 (N_35445,N_35078,N_35001);
nand U35446 (N_35446,N_35052,N_35247);
xor U35447 (N_35447,N_35161,N_35050);
nor U35448 (N_35448,N_35146,N_35082);
and U35449 (N_35449,N_35163,N_35032);
xor U35450 (N_35450,N_35038,N_35180);
nand U35451 (N_35451,N_35230,N_35125);
and U35452 (N_35452,N_35090,N_35153);
nor U35453 (N_35453,N_35030,N_35010);
and U35454 (N_35454,N_35041,N_35220);
xor U35455 (N_35455,N_35071,N_35083);
or U35456 (N_35456,N_35057,N_35064);
and U35457 (N_35457,N_35229,N_35119);
nor U35458 (N_35458,N_35131,N_35029);
nor U35459 (N_35459,N_35061,N_35078);
xnor U35460 (N_35460,N_35003,N_35142);
xor U35461 (N_35461,N_35059,N_35086);
nor U35462 (N_35462,N_35053,N_35062);
nor U35463 (N_35463,N_35142,N_35215);
and U35464 (N_35464,N_35159,N_35007);
nand U35465 (N_35465,N_35069,N_35205);
nand U35466 (N_35466,N_35228,N_35007);
nor U35467 (N_35467,N_35079,N_35025);
nor U35468 (N_35468,N_35075,N_35178);
and U35469 (N_35469,N_35203,N_35161);
or U35470 (N_35470,N_35189,N_35057);
nor U35471 (N_35471,N_35066,N_35137);
xnor U35472 (N_35472,N_35213,N_35038);
and U35473 (N_35473,N_35126,N_35045);
nand U35474 (N_35474,N_35004,N_35117);
nor U35475 (N_35475,N_35207,N_35123);
or U35476 (N_35476,N_35245,N_35156);
and U35477 (N_35477,N_35144,N_35212);
nor U35478 (N_35478,N_35242,N_35106);
nand U35479 (N_35479,N_35158,N_35124);
and U35480 (N_35480,N_35127,N_35168);
nor U35481 (N_35481,N_35118,N_35172);
and U35482 (N_35482,N_35006,N_35142);
nor U35483 (N_35483,N_35190,N_35072);
nand U35484 (N_35484,N_35057,N_35019);
nand U35485 (N_35485,N_35236,N_35121);
and U35486 (N_35486,N_35148,N_35007);
and U35487 (N_35487,N_35083,N_35173);
and U35488 (N_35488,N_35142,N_35117);
or U35489 (N_35489,N_35040,N_35206);
and U35490 (N_35490,N_35076,N_35176);
or U35491 (N_35491,N_35157,N_35138);
or U35492 (N_35492,N_35073,N_35237);
nor U35493 (N_35493,N_35180,N_35190);
or U35494 (N_35494,N_35065,N_35043);
nor U35495 (N_35495,N_35024,N_35142);
and U35496 (N_35496,N_35224,N_35042);
nor U35497 (N_35497,N_35108,N_35238);
nand U35498 (N_35498,N_35180,N_35130);
or U35499 (N_35499,N_35034,N_35090);
nor U35500 (N_35500,N_35370,N_35368);
and U35501 (N_35501,N_35402,N_35284);
and U35502 (N_35502,N_35452,N_35393);
and U35503 (N_35503,N_35351,N_35415);
xnor U35504 (N_35504,N_35425,N_35430);
and U35505 (N_35505,N_35277,N_35285);
and U35506 (N_35506,N_35282,N_35389);
and U35507 (N_35507,N_35434,N_35395);
xor U35508 (N_35508,N_35288,N_35275);
xor U35509 (N_35509,N_35380,N_35323);
nand U35510 (N_35510,N_35459,N_35458);
or U35511 (N_35511,N_35305,N_35291);
xor U35512 (N_35512,N_35441,N_35426);
xnor U35513 (N_35513,N_35475,N_35278);
nand U35514 (N_35514,N_35480,N_35332);
or U35515 (N_35515,N_35442,N_35422);
nor U35516 (N_35516,N_35479,N_35372);
nand U35517 (N_35517,N_35322,N_35270);
and U35518 (N_35518,N_35478,N_35319);
or U35519 (N_35519,N_35465,N_35439);
xnor U35520 (N_35520,N_35431,N_35286);
or U35521 (N_35521,N_35413,N_35261);
or U35522 (N_35522,N_35259,N_35367);
and U35523 (N_35523,N_35271,N_35295);
nand U35524 (N_35524,N_35390,N_35409);
nor U35525 (N_35525,N_35348,N_35418);
or U35526 (N_35526,N_35363,N_35349);
and U35527 (N_35527,N_35398,N_35283);
xnor U35528 (N_35528,N_35341,N_35481);
and U35529 (N_35529,N_35451,N_35336);
and U35530 (N_35530,N_35362,N_35460);
nand U35531 (N_35531,N_35350,N_35345);
and U35532 (N_35532,N_35330,N_35464);
or U35533 (N_35533,N_35400,N_35308);
nand U35534 (N_35534,N_35429,N_35366);
nand U35535 (N_35535,N_35498,N_35469);
xnor U35536 (N_35536,N_35450,N_35326);
nor U35537 (N_35537,N_35416,N_35489);
xor U35538 (N_35538,N_35387,N_35353);
nor U35539 (N_35539,N_35280,N_35455);
xnor U35540 (N_35540,N_35297,N_35281);
nand U35541 (N_35541,N_35411,N_35352);
nand U35542 (N_35542,N_35333,N_35437);
xnor U35543 (N_35543,N_35392,N_35384);
or U35544 (N_35544,N_35378,N_35444);
nand U35545 (N_35545,N_35253,N_35254);
xnor U35546 (N_35546,N_35347,N_35321);
or U35547 (N_35547,N_35410,N_35360);
or U35548 (N_35548,N_35412,N_35406);
and U35549 (N_35549,N_35274,N_35487);
or U35550 (N_35550,N_35421,N_35260);
and U35551 (N_35551,N_35493,N_35334);
nand U35552 (N_35552,N_35289,N_35327);
nand U35553 (N_35553,N_35420,N_35265);
nor U35554 (N_35554,N_35382,N_35462);
nor U35555 (N_35555,N_35267,N_35309);
nor U35556 (N_35556,N_35339,N_35371);
and U35557 (N_35557,N_35302,N_35375);
and U35558 (N_35558,N_35468,N_35456);
xor U35559 (N_35559,N_35419,N_35445);
and U35560 (N_35560,N_35407,N_35258);
nand U35561 (N_35561,N_35293,N_35374);
xor U35562 (N_35562,N_35318,N_35401);
nor U35563 (N_35563,N_35474,N_35262);
xnor U35564 (N_35564,N_35325,N_35391);
xnor U35565 (N_35565,N_35476,N_35461);
nand U35566 (N_35566,N_35383,N_35317);
or U35567 (N_35567,N_35495,N_35306);
nand U35568 (N_35568,N_35359,N_35335);
xor U35569 (N_35569,N_35453,N_35255);
xnor U35570 (N_35570,N_35328,N_35273);
nor U35571 (N_35571,N_35342,N_35446);
nand U35572 (N_35572,N_35377,N_35344);
and U35573 (N_35573,N_35443,N_35449);
and U35574 (N_35574,N_35436,N_35405);
nand U35575 (N_35575,N_35399,N_35435);
nor U35576 (N_35576,N_35263,N_35397);
nor U35577 (N_35577,N_35269,N_35304);
xor U35578 (N_35578,N_35463,N_35264);
and U35579 (N_35579,N_35340,N_35354);
and U35580 (N_35580,N_35329,N_35250);
and U35581 (N_35581,N_35396,N_35364);
nor U35582 (N_35582,N_35355,N_35346);
and U35583 (N_35583,N_35408,N_35386);
or U35584 (N_35584,N_35448,N_35338);
and U35585 (N_35585,N_35484,N_35432);
and U35586 (N_35586,N_35365,N_35482);
or U35587 (N_35587,N_35256,N_35470);
nor U35588 (N_35588,N_35257,N_35454);
and U35589 (N_35589,N_35294,N_35385);
or U35590 (N_35590,N_35314,N_35343);
xnor U35591 (N_35591,N_35485,N_35313);
and U35592 (N_35592,N_35272,N_35361);
or U35593 (N_35593,N_35494,N_35252);
xnor U35594 (N_35594,N_35491,N_35320);
and U35595 (N_35595,N_35486,N_35403);
and U35596 (N_35596,N_35466,N_35497);
nor U35597 (N_35597,N_35279,N_35483);
xor U35598 (N_35598,N_35388,N_35417);
and U35599 (N_35599,N_35251,N_35467);
nand U35600 (N_35600,N_35471,N_35331);
xnor U35601 (N_35601,N_35316,N_35447);
or U35602 (N_35602,N_35490,N_35303);
nand U35603 (N_35603,N_35337,N_35358);
nor U35604 (N_35604,N_35296,N_35496);
or U35605 (N_35605,N_35369,N_35300);
and U35606 (N_35606,N_35299,N_35488);
nand U35607 (N_35607,N_35457,N_35324);
nand U35608 (N_35608,N_35428,N_35427);
nor U35609 (N_35609,N_35473,N_35268);
nor U35610 (N_35610,N_35292,N_35477);
and U35611 (N_35611,N_35440,N_35307);
or U35612 (N_35612,N_35472,N_35276);
and U35613 (N_35613,N_35287,N_35379);
xor U35614 (N_35614,N_35433,N_35356);
nand U35615 (N_35615,N_35301,N_35298);
or U35616 (N_35616,N_35499,N_35357);
nor U35617 (N_35617,N_35381,N_35404);
nand U35618 (N_35618,N_35312,N_35266);
nor U35619 (N_35619,N_35394,N_35315);
nor U35620 (N_35620,N_35492,N_35424);
nand U35621 (N_35621,N_35310,N_35414);
xnor U35622 (N_35622,N_35290,N_35376);
xnor U35623 (N_35623,N_35423,N_35438);
and U35624 (N_35624,N_35373,N_35311);
xor U35625 (N_35625,N_35353,N_35390);
nor U35626 (N_35626,N_35492,N_35433);
nand U35627 (N_35627,N_35440,N_35415);
nor U35628 (N_35628,N_35294,N_35382);
or U35629 (N_35629,N_35349,N_35301);
or U35630 (N_35630,N_35432,N_35332);
xor U35631 (N_35631,N_35394,N_35251);
nand U35632 (N_35632,N_35476,N_35431);
and U35633 (N_35633,N_35471,N_35363);
and U35634 (N_35634,N_35309,N_35483);
and U35635 (N_35635,N_35260,N_35353);
nor U35636 (N_35636,N_35424,N_35289);
nor U35637 (N_35637,N_35301,N_35291);
or U35638 (N_35638,N_35472,N_35479);
or U35639 (N_35639,N_35326,N_35266);
or U35640 (N_35640,N_35328,N_35433);
nand U35641 (N_35641,N_35494,N_35410);
xnor U35642 (N_35642,N_35378,N_35366);
and U35643 (N_35643,N_35334,N_35440);
nand U35644 (N_35644,N_35322,N_35328);
or U35645 (N_35645,N_35463,N_35423);
and U35646 (N_35646,N_35384,N_35436);
xnor U35647 (N_35647,N_35456,N_35366);
or U35648 (N_35648,N_35288,N_35416);
or U35649 (N_35649,N_35350,N_35308);
and U35650 (N_35650,N_35344,N_35342);
and U35651 (N_35651,N_35471,N_35481);
or U35652 (N_35652,N_35354,N_35353);
nand U35653 (N_35653,N_35434,N_35315);
nand U35654 (N_35654,N_35438,N_35294);
nand U35655 (N_35655,N_35367,N_35469);
and U35656 (N_35656,N_35456,N_35264);
nor U35657 (N_35657,N_35468,N_35349);
and U35658 (N_35658,N_35317,N_35423);
xor U35659 (N_35659,N_35426,N_35395);
nor U35660 (N_35660,N_35474,N_35451);
nand U35661 (N_35661,N_35488,N_35410);
and U35662 (N_35662,N_35384,N_35387);
and U35663 (N_35663,N_35291,N_35472);
and U35664 (N_35664,N_35330,N_35451);
xnor U35665 (N_35665,N_35490,N_35428);
xnor U35666 (N_35666,N_35339,N_35350);
and U35667 (N_35667,N_35337,N_35371);
xnor U35668 (N_35668,N_35488,N_35491);
or U35669 (N_35669,N_35438,N_35331);
or U35670 (N_35670,N_35407,N_35423);
or U35671 (N_35671,N_35470,N_35434);
and U35672 (N_35672,N_35311,N_35443);
nand U35673 (N_35673,N_35427,N_35314);
nor U35674 (N_35674,N_35251,N_35384);
nand U35675 (N_35675,N_35343,N_35297);
and U35676 (N_35676,N_35352,N_35288);
nand U35677 (N_35677,N_35326,N_35374);
nor U35678 (N_35678,N_35388,N_35278);
nand U35679 (N_35679,N_35440,N_35330);
nor U35680 (N_35680,N_35424,N_35262);
nor U35681 (N_35681,N_35380,N_35270);
and U35682 (N_35682,N_35383,N_35308);
nand U35683 (N_35683,N_35413,N_35448);
nor U35684 (N_35684,N_35479,N_35389);
nor U35685 (N_35685,N_35377,N_35477);
or U35686 (N_35686,N_35361,N_35383);
and U35687 (N_35687,N_35488,N_35324);
nand U35688 (N_35688,N_35356,N_35460);
and U35689 (N_35689,N_35404,N_35371);
or U35690 (N_35690,N_35370,N_35398);
xnor U35691 (N_35691,N_35287,N_35308);
xor U35692 (N_35692,N_35486,N_35431);
and U35693 (N_35693,N_35275,N_35373);
nor U35694 (N_35694,N_35459,N_35279);
or U35695 (N_35695,N_35389,N_35344);
nand U35696 (N_35696,N_35377,N_35399);
xor U35697 (N_35697,N_35264,N_35285);
xnor U35698 (N_35698,N_35296,N_35321);
nor U35699 (N_35699,N_35311,N_35271);
xnor U35700 (N_35700,N_35294,N_35478);
xor U35701 (N_35701,N_35432,N_35373);
nand U35702 (N_35702,N_35470,N_35490);
and U35703 (N_35703,N_35443,N_35462);
nor U35704 (N_35704,N_35469,N_35441);
nor U35705 (N_35705,N_35314,N_35349);
nand U35706 (N_35706,N_35261,N_35301);
and U35707 (N_35707,N_35351,N_35473);
nor U35708 (N_35708,N_35327,N_35468);
nor U35709 (N_35709,N_35465,N_35406);
xor U35710 (N_35710,N_35384,N_35372);
nor U35711 (N_35711,N_35462,N_35386);
xnor U35712 (N_35712,N_35349,N_35384);
or U35713 (N_35713,N_35307,N_35443);
xnor U35714 (N_35714,N_35488,N_35273);
nand U35715 (N_35715,N_35304,N_35423);
or U35716 (N_35716,N_35423,N_35443);
or U35717 (N_35717,N_35474,N_35435);
nand U35718 (N_35718,N_35259,N_35387);
nor U35719 (N_35719,N_35382,N_35257);
nand U35720 (N_35720,N_35430,N_35283);
or U35721 (N_35721,N_35288,N_35413);
nor U35722 (N_35722,N_35462,N_35275);
or U35723 (N_35723,N_35386,N_35335);
and U35724 (N_35724,N_35450,N_35437);
nor U35725 (N_35725,N_35485,N_35374);
or U35726 (N_35726,N_35419,N_35343);
xnor U35727 (N_35727,N_35495,N_35314);
xnor U35728 (N_35728,N_35331,N_35272);
or U35729 (N_35729,N_35473,N_35449);
nor U35730 (N_35730,N_35300,N_35341);
nor U35731 (N_35731,N_35314,N_35338);
nand U35732 (N_35732,N_35434,N_35421);
or U35733 (N_35733,N_35367,N_35458);
xor U35734 (N_35734,N_35462,N_35266);
xor U35735 (N_35735,N_35433,N_35280);
nor U35736 (N_35736,N_35480,N_35437);
nor U35737 (N_35737,N_35314,N_35479);
xor U35738 (N_35738,N_35490,N_35418);
nand U35739 (N_35739,N_35370,N_35266);
and U35740 (N_35740,N_35444,N_35384);
xor U35741 (N_35741,N_35344,N_35462);
nand U35742 (N_35742,N_35341,N_35434);
nand U35743 (N_35743,N_35433,N_35404);
nor U35744 (N_35744,N_35416,N_35330);
nand U35745 (N_35745,N_35367,N_35286);
or U35746 (N_35746,N_35264,N_35355);
nor U35747 (N_35747,N_35364,N_35288);
and U35748 (N_35748,N_35487,N_35273);
nor U35749 (N_35749,N_35328,N_35250);
and U35750 (N_35750,N_35528,N_35575);
nor U35751 (N_35751,N_35701,N_35716);
or U35752 (N_35752,N_35541,N_35569);
xor U35753 (N_35753,N_35645,N_35508);
and U35754 (N_35754,N_35593,N_35678);
or U35755 (N_35755,N_35551,N_35705);
nor U35756 (N_35756,N_35549,N_35522);
or U35757 (N_35757,N_35666,N_35709);
and U35758 (N_35758,N_35662,N_35746);
nand U35759 (N_35759,N_35553,N_35505);
and U35760 (N_35760,N_35591,N_35511);
nand U35761 (N_35761,N_35675,N_35580);
and U35762 (N_35762,N_35589,N_35558);
or U35763 (N_35763,N_35628,N_35543);
nor U35764 (N_35764,N_35739,N_35620);
xor U35765 (N_35765,N_35597,N_35725);
or U35766 (N_35766,N_35616,N_35512);
xor U35767 (N_35767,N_35563,N_35586);
nor U35768 (N_35768,N_35680,N_35603);
and U35769 (N_35769,N_35587,N_35656);
and U35770 (N_35770,N_35623,N_35719);
and U35771 (N_35771,N_35595,N_35704);
or U35772 (N_35772,N_35609,N_35599);
or U35773 (N_35773,N_35721,N_35674);
nor U35774 (N_35774,N_35652,N_35577);
nand U35775 (N_35775,N_35735,N_35607);
and U35776 (N_35776,N_35622,N_35556);
nor U35777 (N_35777,N_35625,N_35745);
and U35778 (N_35778,N_35687,N_35600);
nand U35779 (N_35779,N_35540,N_35516);
or U35780 (N_35780,N_35657,N_35738);
and U35781 (N_35781,N_35530,N_35631);
nand U35782 (N_35782,N_35510,N_35611);
or U35783 (N_35783,N_35546,N_35677);
or U35784 (N_35784,N_35736,N_35690);
nor U35785 (N_35785,N_35639,N_35732);
nor U35786 (N_35786,N_35727,N_35536);
and U35787 (N_35787,N_35682,N_35728);
nor U35788 (N_35788,N_35706,N_35723);
or U35789 (N_35789,N_35545,N_35720);
xor U35790 (N_35790,N_35604,N_35668);
and U35791 (N_35791,N_35564,N_35646);
or U35792 (N_35792,N_35585,N_35697);
or U35793 (N_35793,N_35681,N_35602);
and U35794 (N_35794,N_35520,N_35529);
and U35795 (N_35795,N_35596,N_35629);
and U35796 (N_35796,N_35747,N_35547);
xor U35797 (N_35797,N_35647,N_35513);
and U35798 (N_35798,N_35658,N_35671);
or U35799 (N_35799,N_35708,N_35743);
nor U35800 (N_35800,N_35581,N_35571);
nand U35801 (N_35801,N_35518,N_35670);
nor U35802 (N_35802,N_35521,N_35523);
xnor U35803 (N_35803,N_35576,N_35637);
xor U35804 (N_35804,N_35660,N_35742);
nor U35805 (N_35805,N_35506,N_35694);
nor U35806 (N_35806,N_35538,N_35578);
nand U35807 (N_35807,N_35626,N_35582);
xnor U35808 (N_35808,N_35726,N_35534);
nand U35809 (N_35809,N_35574,N_35729);
nand U35810 (N_35810,N_35627,N_35684);
xor U35811 (N_35811,N_35612,N_35749);
nor U35812 (N_35812,N_35557,N_35568);
nand U35813 (N_35813,N_35698,N_35696);
nor U35814 (N_35814,N_35524,N_35614);
xor U35815 (N_35815,N_35640,N_35615);
xor U35816 (N_35816,N_35648,N_35651);
or U35817 (N_35817,N_35608,N_35526);
or U35818 (N_35818,N_35592,N_35503);
nor U35819 (N_35819,N_35606,N_35552);
nor U35820 (N_35820,N_35643,N_35744);
and U35821 (N_35821,N_35531,N_35533);
or U35822 (N_35822,N_35559,N_35644);
and U35823 (N_35823,N_35554,N_35693);
xnor U35824 (N_35824,N_35669,N_35686);
and U35825 (N_35825,N_35740,N_35642);
and U35826 (N_35826,N_35741,N_35562);
nand U35827 (N_35827,N_35548,N_35679);
or U35828 (N_35828,N_35689,N_35717);
xnor U35829 (N_35829,N_35565,N_35653);
nand U35830 (N_35830,N_35673,N_35624);
and U35831 (N_35831,N_35509,N_35663);
or U35832 (N_35832,N_35699,N_35667);
and U35833 (N_35833,N_35542,N_35598);
nand U35834 (N_35834,N_35590,N_35504);
xor U35835 (N_35835,N_35573,N_35567);
xnor U35836 (N_35836,N_35733,N_35617);
nand U35837 (N_35837,N_35527,N_35532);
nand U35838 (N_35838,N_35621,N_35692);
nor U35839 (N_35839,N_35664,N_35650);
xor U35840 (N_35840,N_35584,N_35712);
or U35841 (N_35841,N_35594,N_35630);
or U35842 (N_35842,N_35579,N_35714);
or U35843 (N_35843,N_35730,N_35535);
xor U35844 (N_35844,N_35537,N_35702);
nand U35845 (N_35845,N_35649,N_35710);
and U35846 (N_35846,N_35539,N_35501);
or U35847 (N_35847,N_35560,N_35665);
or U35848 (N_35848,N_35588,N_35700);
nand U35849 (N_35849,N_35507,N_35676);
and U35850 (N_35850,N_35661,N_35724);
nand U35851 (N_35851,N_35722,N_35655);
nand U35852 (N_35852,N_35659,N_35517);
nand U35853 (N_35853,N_35634,N_35672);
and U35854 (N_35854,N_35561,N_35515);
nor U35855 (N_35855,N_35550,N_35711);
and U35856 (N_35856,N_35737,N_35618);
nor U35857 (N_35857,N_35500,N_35525);
xnor U35858 (N_35858,N_35683,N_35555);
nand U35859 (N_35859,N_35583,N_35502);
nand U35860 (N_35860,N_35734,N_35748);
nor U35861 (N_35861,N_35641,N_35703);
nor U35862 (N_35862,N_35654,N_35570);
nand U35863 (N_35863,N_35638,N_35605);
nor U35864 (N_35864,N_35613,N_35572);
and U35865 (N_35865,N_35632,N_35718);
or U35866 (N_35866,N_35636,N_35688);
and U35867 (N_35867,N_35691,N_35715);
or U35868 (N_35868,N_35635,N_35731);
and U35869 (N_35869,N_35685,N_35544);
or U35870 (N_35870,N_35619,N_35633);
and U35871 (N_35871,N_35713,N_35695);
nor U35872 (N_35872,N_35514,N_35707);
and U35873 (N_35873,N_35601,N_35610);
xnor U35874 (N_35874,N_35519,N_35566);
and U35875 (N_35875,N_35536,N_35570);
nand U35876 (N_35876,N_35628,N_35729);
and U35877 (N_35877,N_35539,N_35592);
nand U35878 (N_35878,N_35687,N_35514);
and U35879 (N_35879,N_35610,N_35685);
or U35880 (N_35880,N_35535,N_35552);
nor U35881 (N_35881,N_35676,N_35742);
xor U35882 (N_35882,N_35659,N_35670);
nor U35883 (N_35883,N_35739,N_35602);
or U35884 (N_35884,N_35560,N_35579);
nand U35885 (N_35885,N_35685,N_35733);
and U35886 (N_35886,N_35666,N_35653);
nand U35887 (N_35887,N_35677,N_35606);
nand U35888 (N_35888,N_35682,N_35742);
or U35889 (N_35889,N_35733,N_35679);
nand U35890 (N_35890,N_35579,N_35588);
xor U35891 (N_35891,N_35581,N_35725);
or U35892 (N_35892,N_35570,N_35632);
xnor U35893 (N_35893,N_35502,N_35501);
and U35894 (N_35894,N_35610,N_35742);
and U35895 (N_35895,N_35746,N_35522);
xor U35896 (N_35896,N_35629,N_35678);
or U35897 (N_35897,N_35660,N_35726);
or U35898 (N_35898,N_35624,N_35587);
xor U35899 (N_35899,N_35697,N_35514);
or U35900 (N_35900,N_35734,N_35655);
xor U35901 (N_35901,N_35584,N_35514);
and U35902 (N_35902,N_35636,N_35648);
xnor U35903 (N_35903,N_35643,N_35557);
and U35904 (N_35904,N_35700,N_35551);
nand U35905 (N_35905,N_35578,N_35544);
and U35906 (N_35906,N_35631,N_35669);
nand U35907 (N_35907,N_35676,N_35517);
xnor U35908 (N_35908,N_35672,N_35568);
xor U35909 (N_35909,N_35652,N_35521);
or U35910 (N_35910,N_35520,N_35513);
and U35911 (N_35911,N_35696,N_35731);
and U35912 (N_35912,N_35631,N_35711);
xor U35913 (N_35913,N_35748,N_35703);
or U35914 (N_35914,N_35554,N_35709);
nand U35915 (N_35915,N_35508,N_35634);
or U35916 (N_35916,N_35655,N_35747);
nor U35917 (N_35917,N_35582,N_35598);
or U35918 (N_35918,N_35589,N_35538);
and U35919 (N_35919,N_35631,N_35606);
xor U35920 (N_35920,N_35617,N_35543);
xnor U35921 (N_35921,N_35704,N_35549);
and U35922 (N_35922,N_35689,N_35595);
and U35923 (N_35923,N_35543,N_35520);
nand U35924 (N_35924,N_35538,N_35633);
xnor U35925 (N_35925,N_35704,N_35531);
and U35926 (N_35926,N_35636,N_35503);
xor U35927 (N_35927,N_35634,N_35693);
and U35928 (N_35928,N_35719,N_35599);
and U35929 (N_35929,N_35640,N_35599);
or U35930 (N_35930,N_35685,N_35525);
xnor U35931 (N_35931,N_35657,N_35562);
xnor U35932 (N_35932,N_35721,N_35675);
or U35933 (N_35933,N_35514,N_35643);
or U35934 (N_35934,N_35720,N_35690);
nor U35935 (N_35935,N_35572,N_35585);
or U35936 (N_35936,N_35572,N_35664);
and U35937 (N_35937,N_35645,N_35650);
nor U35938 (N_35938,N_35655,N_35719);
and U35939 (N_35939,N_35590,N_35532);
nor U35940 (N_35940,N_35749,N_35576);
nand U35941 (N_35941,N_35513,N_35626);
and U35942 (N_35942,N_35669,N_35723);
and U35943 (N_35943,N_35738,N_35610);
nand U35944 (N_35944,N_35663,N_35709);
xnor U35945 (N_35945,N_35599,N_35519);
nand U35946 (N_35946,N_35642,N_35664);
nand U35947 (N_35947,N_35563,N_35546);
or U35948 (N_35948,N_35614,N_35566);
nor U35949 (N_35949,N_35604,N_35745);
nand U35950 (N_35950,N_35710,N_35650);
and U35951 (N_35951,N_35734,N_35621);
nand U35952 (N_35952,N_35541,N_35509);
nor U35953 (N_35953,N_35604,N_35564);
and U35954 (N_35954,N_35566,N_35629);
nor U35955 (N_35955,N_35631,N_35663);
or U35956 (N_35956,N_35605,N_35716);
nor U35957 (N_35957,N_35679,N_35656);
nor U35958 (N_35958,N_35634,N_35624);
nor U35959 (N_35959,N_35704,N_35637);
nand U35960 (N_35960,N_35665,N_35544);
nor U35961 (N_35961,N_35528,N_35661);
or U35962 (N_35962,N_35654,N_35566);
or U35963 (N_35963,N_35629,N_35557);
and U35964 (N_35964,N_35747,N_35673);
and U35965 (N_35965,N_35668,N_35731);
nand U35966 (N_35966,N_35674,N_35516);
or U35967 (N_35967,N_35704,N_35605);
nor U35968 (N_35968,N_35601,N_35701);
and U35969 (N_35969,N_35608,N_35671);
xor U35970 (N_35970,N_35608,N_35690);
and U35971 (N_35971,N_35651,N_35733);
or U35972 (N_35972,N_35657,N_35670);
or U35973 (N_35973,N_35603,N_35741);
xnor U35974 (N_35974,N_35586,N_35700);
nor U35975 (N_35975,N_35506,N_35571);
xnor U35976 (N_35976,N_35699,N_35703);
nor U35977 (N_35977,N_35711,N_35556);
nand U35978 (N_35978,N_35715,N_35502);
and U35979 (N_35979,N_35627,N_35547);
or U35980 (N_35980,N_35549,N_35626);
and U35981 (N_35981,N_35653,N_35595);
nor U35982 (N_35982,N_35678,N_35690);
nand U35983 (N_35983,N_35701,N_35727);
nand U35984 (N_35984,N_35517,N_35579);
and U35985 (N_35985,N_35726,N_35664);
or U35986 (N_35986,N_35507,N_35504);
and U35987 (N_35987,N_35620,N_35584);
and U35988 (N_35988,N_35671,N_35523);
nand U35989 (N_35989,N_35507,N_35703);
and U35990 (N_35990,N_35621,N_35536);
xnor U35991 (N_35991,N_35569,N_35677);
xor U35992 (N_35992,N_35622,N_35646);
or U35993 (N_35993,N_35731,N_35570);
nand U35994 (N_35994,N_35614,N_35687);
and U35995 (N_35995,N_35732,N_35602);
nand U35996 (N_35996,N_35551,N_35660);
xnor U35997 (N_35997,N_35525,N_35570);
nor U35998 (N_35998,N_35504,N_35693);
nand U35999 (N_35999,N_35633,N_35621);
or U36000 (N_36000,N_35812,N_35860);
nand U36001 (N_36001,N_35964,N_35959);
nand U36002 (N_36002,N_35914,N_35930);
and U36003 (N_36003,N_35985,N_35897);
xnor U36004 (N_36004,N_35990,N_35983);
and U36005 (N_36005,N_35858,N_35942);
nand U36006 (N_36006,N_35881,N_35760);
xnor U36007 (N_36007,N_35789,N_35788);
nor U36008 (N_36008,N_35813,N_35893);
nor U36009 (N_36009,N_35937,N_35989);
xnor U36010 (N_36010,N_35886,N_35764);
or U36011 (N_36011,N_35817,N_35808);
xnor U36012 (N_36012,N_35868,N_35856);
nand U36013 (N_36013,N_35908,N_35899);
or U36014 (N_36014,N_35978,N_35870);
nor U36015 (N_36015,N_35915,N_35963);
nand U36016 (N_36016,N_35782,N_35861);
or U36017 (N_36017,N_35774,N_35962);
nor U36018 (N_36018,N_35887,N_35957);
xor U36019 (N_36019,N_35755,N_35997);
nand U36020 (N_36020,N_35877,N_35982);
xor U36021 (N_36021,N_35876,N_35929);
xor U36022 (N_36022,N_35864,N_35776);
and U36023 (N_36023,N_35979,N_35973);
xnor U36024 (N_36024,N_35980,N_35814);
nand U36025 (N_36025,N_35923,N_35885);
and U36026 (N_36026,N_35777,N_35780);
nand U36027 (N_36027,N_35822,N_35800);
nor U36028 (N_36028,N_35976,N_35775);
and U36029 (N_36029,N_35875,N_35918);
nor U36030 (N_36030,N_35912,N_35878);
nand U36031 (N_36031,N_35867,N_35894);
nor U36032 (N_36032,N_35954,N_35783);
nand U36033 (N_36033,N_35994,N_35836);
xnor U36034 (N_36034,N_35773,N_35905);
and U36035 (N_36035,N_35916,N_35890);
xnor U36036 (N_36036,N_35975,N_35825);
nand U36037 (N_36037,N_35892,N_35940);
and U36038 (N_36038,N_35960,N_35831);
and U36039 (N_36039,N_35901,N_35902);
xnor U36040 (N_36040,N_35966,N_35874);
and U36041 (N_36041,N_35798,N_35819);
nand U36042 (N_36042,N_35784,N_35811);
or U36043 (N_36043,N_35830,N_35810);
nand U36044 (N_36044,N_35913,N_35770);
nand U36045 (N_36045,N_35873,N_35761);
and U36046 (N_36046,N_35993,N_35991);
nor U36047 (N_36047,N_35933,N_35945);
nor U36048 (N_36048,N_35880,N_35907);
and U36049 (N_36049,N_35840,N_35750);
nand U36050 (N_36050,N_35944,N_35824);
nand U36051 (N_36051,N_35906,N_35792);
and U36052 (N_36052,N_35882,N_35790);
nand U36053 (N_36053,N_35818,N_35953);
nor U36054 (N_36054,N_35943,N_35757);
and U36055 (N_36055,N_35932,N_35767);
or U36056 (N_36056,N_35851,N_35846);
nand U36057 (N_36057,N_35816,N_35794);
and U36058 (N_36058,N_35884,N_35986);
or U36059 (N_36059,N_35758,N_35765);
or U36060 (N_36060,N_35947,N_35834);
or U36061 (N_36061,N_35863,N_35772);
nor U36062 (N_36062,N_35859,N_35766);
nand U36063 (N_36063,N_35987,N_35970);
xor U36064 (N_36064,N_35936,N_35807);
or U36065 (N_36065,N_35862,N_35967);
and U36066 (N_36066,N_35852,N_35797);
nor U36067 (N_36067,N_35857,N_35998);
xor U36068 (N_36068,N_35778,N_35823);
and U36069 (N_36069,N_35903,N_35977);
nand U36070 (N_36070,N_35809,N_35839);
and U36071 (N_36071,N_35958,N_35971);
and U36072 (N_36072,N_35802,N_35796);
xor U36073 (N_36073,N_35974,N_35785);
nand U36074 (N_36074,N_35759,N_35879);
nand U36075 (N_36075,N_35951,N_35826);
nand U36076 (N_36076,N_35869,N_35843);
and U36077 (N_36077,N_35753,N_35769);
nand U36078 (N_36078,N_35921,N_35838);
xnor U36079 (N_36079,N_35804,N_35752);
xnor U36080 (N_36080,N_35820,N_35791);
nand U36081 (N_36081,N_35754,N_35756);
or U36082 (N_36082,N_35949,N_35786);
xnor U36083 (N_36083,N_35925,N_35931);
xnor U36084 (N_36084,N_35854,N_35898);
and U36085 (N_36085,N_35848,N_35992);
xnor U36086 (N_36086,N_35946,N_35855);
xor U36087 (N_36087,N_35799,N_35909);
nor U36088 (N_36088,N_35888,N_35941);
nand U36089 (N_36089,N_35803,N_35763);
and U36090 (N_36090,N_35883,N_35935);
and U36091 (N_36091,N_35779,N_35965);
nor U36092 (N_36092,N_35853,N_35806);
or U36093 (N_36093,N_35981,N_35926);
nand U36094 (N_36094,N_35847,N_35844);
nand U36095 (N_36095,N_35845,N_35781);
nor U36096 (N_36096,N_35969,N_35872);
or U36097 (N_36097,N_35850,N_35948);
xnor U36098 (N_36098,N_35793,N_35900);
nor U36099 (N_36099,N_35842,N_35787);
xor U36100 (N_36100,N_35833,N_35972);
and U36101 (N_36101,N_35927,N_35996);
nor U36102 (N_36102,N_35865,N_35896);
nand U36103 (N_36103,N_35762,N_35919);
and U36104 (N_36104,N_35968,N_35827);
and U36105 (N_36105,N_35871,N_35911);
or U36106 (N_36106,N_35832,N_35866);
and U36107 (N_36107,N_35956,N_35828);
and U36108 (N_36108,N_35934,N_35904);
nand U36109 (N_36109,N_35895,N_35961);
nor U36110 (N_36110,N_35917,N_35920);
and U36111 (N_36111,N_35837,N_35999);
or U36112 (N_36112,N_35835,N_35805);
xor U36113 (N_36113,N_35939,N_35952);
nor U36114 (N_36114,N_35821,N_35815);
and U36115 (N_36115,N_35988,N_35938);
or U36116 (N_36116,N_35801,N_35928);
xnor U36117 (N_36117,N_35955,N_35849);
xnor U36118 (N_36118,N_35995,N_35891);
or U36119 (N_36119,N_35922,N_35751);
xor U36120 (N_36120,N_35768,N_35950);
xor U36121 (N_36121,N_35795,N_35841);
nand U36122 (N_36122,N_35829,N_35924);
nand U36123 (N_36123,N_35910,N_35984);
xnor U36124 (N_36124,N_35771,N_35889);
nand U36125 (N_36125,N_35850,N_35997);
xor U36126 (N_36126,N_35857,N_35823);
nor U36127 (N_36127,N_35956,N_35805);
nor U36128 (N_36128,N_35977,N_35821);
or U36129 (N_36129,N_35873,N_35897);
xnor U36130 (N_36130,N_35981,N_35862);
and U36131 (N_36131,N_35854,N_35973);
or U36132 (N_36132,N_35817,N_35958);
or U36133 (N_36133,N_35789,N_35924);
nand U36134 (N_36134,N_35976,N_35926);
nor U36135 (N_36135,N_35923,N_35975);
xnor U36136 (N_36136,N_35788,N_35822);
nand U36137 (N_36137,N_35912,N_35883);
or U36138 (N_36138,N_35966,N_35758);
xnor U36139 (N_36139,N_35800,N_35828);
or U36140 (N_36140,N_35767,N_35770);
or U36141 (N_36141,N_35876,N_35849);
xor U36142 (N_36142,N_35831,N_35822);
or U36143 (N_36143,N_35829,N_35779);
xor U36144 (N_36144,N_35892,N_35894);
nor U36145 (N_36145,N_35809,N_35825);
xor U36146 (N_36146,N_35974,N_35811);
or U36147 (N_36147,N_35942,N_35999);
xor U36148 (N_36148,N_35826,N_35864);
and U36149 (N_36149,N_35966,N_35762);
xnor U36150 (N_36150,N_35861,N_35875);
and U36151 (N_36151,N_35976,N_35764);
or U36152 (N_36152,N_35816,N_35841);
or U36153 (N_36153,N_35774,N_35904);
nand U36154 (N_36154,N_35961,N_35947);
or U36155 (N_36155,N_35900,N_35912);
or U36156 (N_36156,N_35899,N_35951);
and U36157 (N_36157,N_35892,N_35913);
xnor U36158 (N_36158,N_35845,N_35806);
nor U36159 (N_36159,N_35914,N_35808);
or U36160 (N_36160,N_35800,N_35757);
nor U36161 (N_36161,N_35999,N_35753);
or U36162 (N_36162,N_35973,N_35777);
nand U36163 (N_36163,N_35849,N_35971);
nor U36164 (N_36164,N_35839,N_35903);
nor U36165 (N_36165,N_35839,N_35779);
or U36166 (N_36166,N_35935,N_35970);
and U36167 (N_36167,N_35813,N_35891);
xnor U36168 (N_36168,N_35999,N_35862);
xor U36169 (N_36169,N_35776,N_35915);
nor U36170 (N_36170,N_35919,N_35874);
nor U36171 (N_36171,N_35775,N_35859);
nand U36172 (N_36172,N_35906,N_35942);
nor U36173 (N_36173,N_35977,N_35938);
or U36174 (N_36174,N_35757,N_35871);
and U36175 (N_36175,N_35802,N_35989);
nand U36176 (N_36176,N_35789,N_35818);
and U36177 (N_36177,N_35911,N_35931);
xnor U36178 (N_36178,N_35993,N_35869);
and U36179 (N_36179,N_35991,N_35924);
and U36180 (N_36180,N_35851,N_35924);
or U36181 (N_36181,N_35768,N_35903);
nand U36182 (N_36182,N_35982,N_35870);
nor U36183 (N_36183,N_35934,N_35840);
or U36184 (N_36184,N_35876,N_35840);
or U36185 (N_36185,N_35761,N_35817);
nand U36186 (N_36186,N_35795,N_35796);
nand U36187 (N_36187,N_35963,N_35833);
xnor U36188 (N_36188,N_35792,N_35986);
nand U36189 (N_36189,N_35800,N_35935);
nor U36190 (N_36190,N_35844,N_35965);
nand U36191 (N_36191,N_35752,N_35920);
or U36192 (N_36192,N_35977,N_35882);
nand U36193 (N_36193,N_35843,N_35793);
and U36194 (N_36194,N_35875,N_35950);
and U36195 (N_36195,N_35763,N_35965);
nor U36196 (N_36196,N_35919,N_35934);
nand U36197 (N_36197,N_35937,N_35806);
nand U36198 (N_36198,N_35792,N_35993);
nand U36199 (N_36199,N_35796,N_35994);
or U36200 (N_36200,N_35960,N_35917);
or U36201 (N_36201,N_35816,N_35783);
xnor U36202 (N_36202,N_35933,N_35813);
xnor U36203 (N_36203,N_35775,N_35900);
or U36204 (N_36204,N_35768,N_35913);
nor U36205 (N_36205,N_35935,N_35875);
xor U36206 (N_36206,N_35979,N_35919);
xor U36207 (N_36207,N_35906,N_35844);
or U36208 (N_36208,N_35999,N_35922);
nand U36209 (N_36209,N_35902,N_35765);
xor U36210 (N_36210,N_35771,N_35767);
or U36211 (N_36211,N_35886,N_35933);
nor U36212 (N_36212,N_35948,N_35984);
nand U36213 (N_36213,N_35751,N_35847);
nor U36214 (N_36214,N_35849,N_35900);
xor U36215 (N_36215,N_35824,N_35868);
nand U36216 (N_36216,N_35848,N_35882);
or U36217 (N_36217,N_35933,N_35987);
nor U36218 (N_36218,N_35779,N_35943);
nor U36219 (N_36219,N_35914,N_35860);
nor U36220 (N_36220,N_35872,N_35996);
or U36221 (N_36221,N_35910,N_35977);
nor U36222 (N_36222,N_35760,N_35886);
xnor U36223 (N_36223,N_35949,N_35914);
nor U36224 (N_36224,N_35753,N_35838);
nor U36225 (N_36225,N_35926,N_35761);
or U36226 (N_36226,N_35810,N_35944);
nor U36227 (N_36227,N_35989,N_35992);
nor U36228 (N_36228,N_35781,N_35973);
nor U36229 (N_36229,N_35833,N_35836);
and U36230 (N_36230,N_35973,N_35882);
nand U36231 (N_36231,N_35884,N_35788);
or U36232 (N_36232,N_35893,N_35911);
xor U36233 (N_36233,N_35876,N_35785);
or U36234 (N_36234,N_35971,N_35936);
nand U36235 (N_36235,N_35784,N_35891);
and U36236 (N_36236,N_35843,N_35920);
and U36237 (N_36237,N_35810,N_35934);
xor U36238 (N_36238,N_35918,N_35759);
and U36239 (N_36239,N_35759,N_35895);
and U36240 (N_36240,N_35803,N_35873);
and U36241 (N_36241,N_35888,N_35769);
nand U36242 (N_36242,N_35808,N_35916);
xnor U36243 (N_36243,N_35967,N_35888);
nor U36244 (N_36244,N_35994,N_35977);
nor U36245 (N_36245,N_35791,N_35802);
nand U36246 (N_36246,N_35802,N_35974);
and U36247 (N_36247,N_35936,N_35809);
nand U36248 (N_36248,N_35773,N_35911);
nand U36249 (N_36249,N_35839,N_35820);
or U36250 (N_36250,N_36182,N_36047);
and U36251 (N_36251,N_36002,N_36236);
nor U36252 (N_36252,N_36228,N_36204);
and U36253 (N_36253,N_36107,N_36185);
nand U36254 (N_36254,N_36093,N_36230);
or U36255 (N_36255,N_36134,N_36101);
or U36256 (N_36256,N_36037,N_36108);
and U36257 (N_36257,N_36021,N_36009);
xnor U36258 (N_36258,N_36171,N_36102);
or U36259 (N_36259,N_36215,N_36241);
xor U36260 (N_36260,N_36232,N_36062);
and U36261 (N_36261,N_36106,N_36068);
or U36262 (N_36262,N_36012,N_36162);
nand U36263 (N_36263,N_36087,N_36027);
nor U36264 (N_36264,N_36126,N_36054);
and U36265 (N_36265,N_36081,N_36077);
nor U36266 (N_36266,N_36235,N_36195);
nor U36267 (N_36267,N_36223,N_36092);
xor U36268 (N_36268,N_36175,N_36104);
nor U36269 (N_36269,N_36017,N_36247);
and U36270 (N_36270,N_36084,N_36048);
and U36271 (N_36271,N_36217,N_36016);
xor U36272 (N_36272,N_36115,N_36160);
xor U36273 (N_36273,N_36111,N_36187);
nand U36274 (N_36274,N_36177,N_36186);
or U36275 (N_36275,N_36000,N_36089);
and U36276 (N_36276,N_36070,N_36044);
nor U36277 (N_36277,N_36146,N_36008);
xnor U36278 (N_36278,N_36165,N_36095);
nand U36279 (N_36279,N_36032,N_36130);
xor U36280 (N_36280,N_36063,N_36196);
and U36281 (N_36281,N_36082,N_36238);
nand U36282 (N_36282,N_36189,N_36213);
or U36283 (N_36283,N_36031,N_36096);
xor U36284 (N_36284,N_36212,N_36197);
nand U36285 (N_36285,N_36139,N_36100);
or U36286 (N_36286,N_36065,N_36210);
xnor U36287 (N_36287,N_36099,N_36073);
or U36288 (N_36288,N_36148,N_36194);
nor U36289 (N_36289,N_36056,N_36038);
nand U36290 (N_36290,N_36103,N_36136);
and U36291 (N_36291,N_36137,N_36117);
nor U36292 (N_36292,N_36173,N_36124);
nand U36293 (N_36293,N_36046,N_36242);
and U36294 (N_36294,N_36222,N_36119);
nor U36295 (N_36295,N_36132,N_36180);
nand U36296 (N_36296,N_36018,N_36026);
xnor U36297 (N_36297,N_36216,N_36041);
or U36298 (N_36298,N_36151,N_36156);
nor U36299 (N_36299,N_36020,N_36015);
nor U36300 (N_36300,N_36135,N_36067);
and U36301 (N_36301,N_36050,N_36221);
xnor U36302 (N_36302,N_36200,N_36231);
or U36303 (N_36303,N_36239,N_36086);
nor U36304 (N_36304,N_36105,N_36227);
nor U36305 (N_36305,N_36207,N_36198);
or U36306 (N_36306,N_36010,N_36094);
and U36307 (N_36307,N_36209,N_36014);
or U36308 (N_36308,N_36055,N_36188);
and U36309 (N_36309,N_36074,N_36022);
xor U36310 (N_36310,N_36005,N_36006);
nand U36311 (N_36311,N_36249,N_36152);
or U36312 (N_36312,N_36127,N_36208);
xor U36313 (N_36313,N_36097,N_36019);
xor U36314 (N_36314,N_36202,N_36233);
xor U36315 (N_36315,N_36001,N_36150);
or U36316 (N_36316,N_36224,N_36024);
xor U36317 (N_36317,N_36168,N_36237);
xnor U36318 (N_36318,N_36218,N_36121);
nand U36319 (N_36319,N_36199,N_36179);
nor U36320 (N_36320,N_36145,N_36064);
xor U36321 (N_36321,N_36118,N_36140);
xnor U36322 (N_36322,N_36114,N_36120);
and U36323 (N_36323,N_36225,N_36109);
and U36324 (N_36324,N_36061,N_36098);
or U36325 (N_36325,N_36085,N_36040);
nor U36326 (N_36326,N_36122,N_36033);
or U36327 (N_36327,N_36243,N_36161);
or U36328 (N_36328,N_36112,N_36157);
nor U36329 (N_36329,N_36158,N_36244);
nand U36330 (N_36330,N_36003,N_36029);
xnor U36331 (N_36331,N_36190,N_36052);
and U36332 (N_36332,N_36181,N_36051);
nand U36333 (N_36333,N_36049,N_36110);
nor U36334 (N_36334,N_36229,N_36036);
xor U36335 (N_36335,N_36028,N_36240);
or U36336 (N_36336,N_36133,N_36039);
and U36337 (N_36337,N_36206,N_36025);
nor U36338 (N_36338,N_36174,N_36219);
nor U36339 (N_36339,N_36131,N_36201);
and U36340 (N_36340,N_36043,N_36142);
nand U36341 (N_36341,N_36205,N_36203);
nand U36342 (N_36342,N_36220,N_36141);
or U36343 (N_36343,N_36079,N_36149);
or U36344 (N_36344,N_36246,N_36076);
xnor U36345 (N_36345,N_36023,N_36080);
and U36346 (N_36346,N_36013,N_36153);
or U36347 (N_36347,N_36091,N_36167);
and U36348 (N_36348,N_36069,N_36007);
xor U36349 (N_36349,N_36170,N_36172);
or U36350 (N_36350,N_36072,N_36211);
nand U36351 (N_36351,N_36058,N_36113);
xor U36352 (N_36352,N_36083,N_36075);
xnor U36353 (N_36353,N_36169,N_36060);
or U36354 (N_36354,N_36226,N_36045);
nand U36355 (N_36355,N_36214,N_36154);
nor U36356 (N_36356,N_36193,N_36138);
xor U36357 (N_36357,N_36192,N_36143);
xor U36358 (N_36358,N_36166,N_36248);
or U36359 (N_36359,N_36057,N_36159);
or U36360 (N_36360,N_36147,N_36245);
xnor U36361 (N_36361,N_36144,N_36034);
and U36362 (N_36362,N_36155,N_36129);
nor U36363 (N_36363,N_36176,N_36004);
or U36364 (N_36364,N_36088,N_36163);
nor U36365 (N_36365,N_36090,N_36234);
nand U36366 (N_36366,N_36164,N_36128);
or U36367 (N_36367,N_36066,N_36071);
and U36368 (N_36368,N_36123,N_36030);
and U36369 (N_36369,N_36125,N_36059);
xor U36370 (N_36370,N_36042,N_36183);
xor U36371 (N_36371,N_36011,N_36178);
nor U36372 (N_36372,N_36053,N_36078);
nand U36373 (N_36373,N_36035,N_36191);
nand U36374 (N_36374,N_36116,N_36184);
or U36375 (N_36375,N_36188,N_36071);
xnor U36376 (N_36376,N_36161,N_36201);
xnor U36377 (N_36377,N_36107,N_36146);
or U36378 (N_36378,N_36014,N_36004);
nand U36379 (N_36379,N_36152,N_36207);
or U36380 (N_36380,N_36119,N_36233);
and U36381 (N_36381,N_36101,N_36200);
nor U36382 (N_36382,N_36059,N_36055);
or U36383 (N_36383,N_36138,N_36022);
or U36384 (N_36384,N_36041,N_36085);
or U36385 (N_36385,N_36059,N_36229);
and U36386 (N_36386,N_36229,N_36066);
or U36387 (N_36387,N_36121,N_36124);
nand U36388 (N_36388,N_36188,N_36048);
or U36389 (N_36389,N_36172,N_36052);
nor U36390 (N_36390,N_36208,N_36222);
xnor U36391 (N_36391,N_36240,N_36093);
and U36392 (N_36392,N_36063,N_36066);
nor U36393 (N_36393,N_36147,N_36221);
nand U36394 (N_36394,N_36245,N_36198);
and U36395 (N_36395,N_36231,N_36220);
nor U36396 (N_36396,N_36196,N_36171);
and U36397 (N_36397,N_36083,N_36187);
xnor U36398 (N_36398,N_36224,N_36118);
nand U36399 (N_36399,N_36214,N_36003);
nor U36400 (N_36400,N_36170,N_36049);
or U36401 (N_36401,N_36100,N_36206);
nand U36402 (N_36402,N_36047,N_36037);
or U36403 (N_36403,N_36056,N_36084);
or U36404 (N_36404,N_36169,N_36195);
nand U36405 (N_36405,N_36035,N_36025);
nor U36406 (N_36406,N_36115,N_36201);
nor U36407 (N_36407,N_36092,N_36120);
or U36408 (N_36408,N_36242,N_36040);
xnor U36409 (N_36409,N_36205,N_36160);
nand U36410 (N_36410,N_36026,N_36136);
xor U36411 (N_36411,N_36071,N_36054);
nor U36412 (N_36412,N_36020,N_36042);
nand U36413 (N_36413,N_36039,N_36120);
or U36414 (N_36414,N_36123,N_36147);
nand U36415 (N_36415,N_36048,N_36016);
or U36416 (N_36416,N_36108,N_36009);
or U36417 (N_36417,N_36212,N_36112);
nand U36418 (N_36418,N_36142,N_36151);
and U36419 (N_36419,N_36184,N_36087);
or U36420 (N_36420,N_36184,N_36206);
xor U36421 (N_36421,N_36029,N_36141);
or U36422 (N_36422,N_36175,N_36050);
nor U36423 (N_36423,N_36147,N_36064);
xnor U36424 (N_36424,N_36010,N_36151);
nand U36425 (N_36425,N_36183,N_36242);
nand U36426 (N_36426,N_36019,N_36111);
xnor U36427 (N_36427,N_36152,N_36051);
nor U36428 (N_36428,N_36096,N_36090);
and U36429 (N_36429,N_36193,N_36100);
nor U36430 (N_36430,N_36089,N_36097);
xnor U36431 (N_36431,N_36165,N_36061);
or U36432 (N_36432,N_36164,N_36000);
xor U36433 (N_36433,N_36130,N_36139);
nor U36434 (N_36434,N_36169,N_36061);
and U36435 (N_36435,N_36010,N_36058);
nand U36436 (N_36436,N_36011,N_36002);
nor U36437 (N_36437,N_36181,N_36091);
nand U36438 (N_36438,N_36196,N_36248);
xor U36439 (N_36439,N_36108,N_36093);
nor U36440 (N_36440,N_36132,N_36036);
or U36441 (N_36441,N_36036,N_36021);
or U36442 (N_36442,N_36091,N_36204);
and U36443 (N_36443,N_36217,N_36148);
and U36444 (N_36444,N_36173,N_36190);
or U36445 (N_36445,N_36093,N_36233);
nor U36446 (N_36446,N_36007,N_36218);
xnor U36447 (N_36447,N_36176,N_36021);
xnor U36448 (N_36448,N_36197,N_36051);
and U36449 (N_36449,N_36156,N_36146);
xnor U36450 (N_36450,N_36238,N_36151);
and U36451 (N_36451,N_36146,N_36239);
or U36452 (N_36452,N_36127,N_36023);
nor U36453 (N_36453,N_36156,N_36111);
xnor U36454 (N_36454,N_36171,N_36216);
or U36455 (N_36455,N_36138,N_36055);
xnor U36456 (N_36456,N_36059,N_36091);
and U36457 (N_36457,N_36068,N_36174);
or U36458 (N_36458,N_36172,N_36028);
nand U36459 (N_36459,N_36218,N_36112);
xor U36460 (N_36460,N_36249,N_36192);
nand U36461 (N_36461,N_36139,N_36153);
or U36462 (N_36462,N_36209,N_36127);
nor U36463 (N_36463,N_36159,N_36023);
or U36464 (N_36464,N_36206,N_36249);
and U36465 (N_36465,N_36078,N_36005);
and U36466 (N_36466,N_36054,N_36134);
or U36467 (N_36467,N_36006,N_36022);
and U36468 (N_36468,N_36119,N_36056);
or U36469 (N_36469,N_36129,N_36239);
and U36470 (N_36470,N_36036,N_36052);
nor U36471 (N_36471,N_36073,N_36236);
xnor U36472 (N_36472,N_36173,N_36035);
nand U36473 (N_36473,N_36207,N_36090);
nor U36474 (N_36474,N_36207,N_36035);
nand U36475 (N_36475,N_36080,N_36138);
and U36476 (N_36476,N_36076,N_36235);
xor U36477 (N_36477,N_36197,N_36227);
nand U36478 (N_36478,N_36166,N_36039);
nand U36479 (N_36479,N_36143,N_36239);
and U36480 (N_36480,N_36134,N_36164);
nor U36481 (N_36481,N_36069,N_36018);
nor U36482 (N_36482,N_36178,N_36079);
xnor U36483 (N_36483,N_36141,N_36195);
nor U36484 (N_36484,N_36067,N_36172);
xor U36485 (N_36485,N_36000,N_36184);
or U36486 (N_36486,N_36109,N_36092);
nor U36487 (N_36487,N_36188,N_36141);
or U36488 (N_36488,N_36169,N_36158);
and U36489 (N_36489,N_36007,N_36026);
or U36490 (N_36490,N_36235,N_36138);
xor U36491 (N_36491,N_36193,N_36196);
nand U36492 (N_36492,N_36141,N_36235);
or U36493 (N_36493,N_36212,N_36057);
nand U36494 (N_36494,N_36101,N_36167);
nand U36495 (N_36495,N_36108,N_36221);
and U36496 (N_36496,N_36085,N_36122);
xor U36497 (N_36497,N_36128,N_36207);
or U36498 (N_36498,N_36133,N_36073);
and U36499 (N_36499,N_36094,N_36176);
or U36500 (N_36500,N_36379,N_36401);
nor U36501 (N_36501,N_36256,N_36477);
xor U36502 (N_36502,N_36283,N_36381);
or U36503 (N_36503,N_36461,N_36429);
xor U36504 (N_36504,N_36475,N_36455);
or U36505 (N_36505,N_36359,N_36324);
or U36506 (N_36506,N_36273,N_36462);
and U36507 (N_36507,N_36496,N_36438);
xor U36508 (N_36508,N_36377,N_36444);
nor U36509 (N_36509,N_36297,N_36451);
nor U36510 (N_36510,N_36287,N_36322);
and U36511 (N_36511,N_36412,N_36345);
nor U36512 (N_36512,N_36485,N_36408);
or U36513 (N_36513,N_36267,N_36436);
nor U36514 (N_36514,N_36358,N_36487);
nor U36515 (N_36515,N_36342,N_36355);
nor U36516 (N_36516,N_36285,N_36383);
or U36517 (N_36517,N_36361,N_36327);
or U36518 (N_36518,N_36263,N_36473);
or U36519 (N_36519,N_36474,N_36304);
xnor U36520 (N_36520,N_36398,N_36385);
xor U36521 (N_36521,N_36426,N_36282);
nor U36522 (N_36522,N_36292,N_36458);
and U36523 (N_36523,N_36492,N_36499);
or U36524 (N_36524,N_36378,N_36270);
nor U36525 (N_36525,N_36319,N_36454);
nand U36526 (N_36526,N_36321,N_36400);
and U36527 (N_36527,N_36331,N_36332);
nand U36528 (N_36528,N_36465,N_36483);
nand U36529 (N_36529,N_36390,N_36480);
nand U36530 (N_36530,N_36305,N_36494);
and U36531 (N_36531,N_36330,N_36456);
nor U36532 (N_36532,N_36391,N_36310);
or U36533 (N_36533,N_36435,N_36303);
xnor U36534 (N_36534,N_36493,N_36349);
nor U36535 (N_36535,N_36411,N_36313);
nand U36536 (N_36536,N_36449,N_36404);
or U36537 (N_36537,N_36286,N_36427);
or U36538 (N_36538,N_36314,N_36479);
nor U36539 (N_36539,N_36459,N_36328);
nand U36540 (N_36540,N_36284,N_36353);
nor U36541 (N_36541,N_36279,N_36323);
nor U36542 (N_36542,N_36251,N_36344);
or U36543 (N_36543,N_36301,N_36470);
or U36544 (N_36544,N_36464,N_36271);
nor U36545 (N_36545,N_36443,N_36296);
and U36546 (N_36546,N_36374,N_36335);
nand U36547 (N_36547,N_36422,N_36482);
and U36548 (N_36548,N_36424,N_36341);
nand U36549 (N_36549,N_36394,N_36269);
xnor U36550 (N_36550,N_36329,N_36347);
nand U36551 (N_36551,N_36425,N_36430);
nor U36552 (N_36552,N_36418,N_36302);
nor U36553 (N_36553,N_36318,N_36491);
xor U36554 (N_36554,N_36300,N_36354);
xor U36555 (N_36555,N_36261,N_36498);
nor U36556 (N_36556,N_36441,N_36295);
nand U36557 (N_36557,N_36417,N_36281);
nand U36558 (N_36558,N_36316,N_36363);
xnor U36559 (N_36559,N_36309,N_36439);
nor U36560 (N_36560,N_36376,N_36440);
xnor U36561 (N_36561,N_36315,N_36397);
nand U36562 (N_36562,N_36333,N_36357);
or U36563 (N_36563,N_36372,N_36336);
or U36564 (N_36564,N_36460,N_36340);
xor U36565 (N_36565,N_36258,N_36471);
nor U36566 (N_36566,N_36288,N_36467);
xnor U36567 (N_36567,N_36469,N_36350);
nand U36568 (N_36568,N_36446,N_36403);
and U36569 (N_36569,N_36291,N_36277);
xor U36570 (N_36570,N_36339,N_36362);
xor U36571 (N_36571,N_36396,N_36389);
or U36572 (N_36572,N_36490,N_36432);
or U36573 (N_36573,N_36268,N_36265);
xor U36574 (N_36574,N_36266,N_36275);
or U36575 (N_36575,N_36253,N_36497);
nor U36576 (N_36576,N_36366,N_36452);
nor U36577 (N_36577,N_36343,N_36307);
and U36578 (N_36578,N_36364,N_36447);
xor U36579 (N_36579,N_36457,N_36402);
or U36580 (N_36580,N_36337,N_36448);
and U36581 (N_36581,N_36254,N_36421);
and U36582 (N_36582,N_36367,N_36259);
or U36583 (N_36583,N_36407,N_36453);
and U36584 (N_36584,N_36413,N_36356);
xor U36585 (N_36585,N_36476,N_36278);
nand U36586 (N_36586,N_36320,N_36368);
and U36587 (N_36587,N_36442,N_36393);
or U36588 (N_36588,N_36410,N_36405);
nor U36589 (N_36589,N_36365,N_36437);
nor U36590 (N_36590,N_36280,N_36386);
or U36591 (N_36591,N_36370,N_36274);
nor U36592 (N_36592,N_36463,N_36478);
and U36593 (N_36593,N_36317,N_36415);
and U36594 (N_36594,N_36346,N_36488);
and U36595 (N_36595,N_36388,N_36360);
xor U36596 (N_36596,N_36466,N_36352);
xnor U36597 (N_36597,N_36250,N_36484);
and U36598 (N_36598,N_36406,N_36375);
nor U36599 (N_36599,N_36252,N_36416);
nor U36600 (N_36600,N_36308,N_36290);
or U36601 (N_36601,N_36293,N_36481);
nand U36602 (N_36602,N_36276,N_36348);
nor U36603 (N_36603,N_36338,N_36373);
or U36604 (N_36604,N_36294,N_36369);
xor U36605 (N_36605,N_36380,N_36395);
and U36606 (N_36606,N_36486,N_36472);
xnor U36607 (N_36607,N_36409,N_36257);
and U36608 (N_36608,N_36423,N_36312);
or U36609 (N_36609,N_36384,N_36351);
xnor U36610 (N_36610,N_36419,N_36289);
or U36611 (N_36611,N_36382,N_36371);
nand U36612 (N_36612,N_36420,N_36431);
xor U36613 (N_36613,N_36306,N_36445);
and U36614 (N_36614,N_36262,N_36325);
or U36615 (N_36615,N_36264,N_36414);
and U36616 (N_36616,N_36495,N_36299);
or U36617 (N_36617,N_36428,N_36433);
and U36618 (N_36618,N_36489,N_36399);
xor U36619 (N_36619,N_36387,N_36260);
nand U36620 (N_36620,N_36298,N_36334);
and U36621 (N_36621,N_36311,N_36468);
or U36622 (N_36622,N_36272,N_36392);
or U36623 (N_36623,N_36450,N_36255);
or U36624 (N_36624,N_36434,N_36326);
nor U36625 (N_36625,N_36369,N_36362);
and U36626 (N_36626,N_36437,N_36369);
or U36627 (N_36627,N_36366,N_36470);
xor U36628 (N_36628,N_36252,N_36271);
xor U36629 (N_36629,N_36271,N_36385);
and U36630 (N_36630,N_36451,N_36321);
nor U36631 (N_36631,N_36471,N_36288);
and U36632 (N_36632,N_36275,N_36495);
nor U36633 (N_36633,N_36316,N_36453);
nand U36634 (N_36634,N_36458,N_36301);
xnor U36635 (N_36635,N_36267,N_36406);
xnor U36636 (N_36636,N_36340,N_36430);
and U36637 (N_36637,N_36287,N_36363);
nand U36638 (N_36638,N_36251,N_36407);
nor U36639 (N_36639,N_36445,N_36414);
xor U36640 (N_36640,N_36253,N_36428);
xor U36641 (N_36641,N_36394,N_36418);
and U36642 (N_36642,N_36425,N_36273);
nor U36643 (N_36643,N_36410,N_36376);
xor U36644 (N_36644,N_36492,N_36264);
nand U36645 (N_36645,N_36281,N_36478);
xor U36646 (N_36646,N_36420,N_36277);
nor U36647 (N_36647,N_36453,N_36470);
nor U36648 (N_36648,N_36369,N_36275);
or U36649 (N_36649,N_36290,N_36427);
nand U36650 (N_36650,N_36290,N_36403);
xor U36651 (N_36651,N_36323,N_36381);
nor U36652 (N_36652,N_36346,N_36481);
and U36653 (N_36653,N_36405,N_36280);
or U36654 (N_36654,N_36275,N_36389);
xnor U36655 (N_36655,N_36435,N_36341);
and U36656 (N_36656,N_36431,N_36407);
nor U36657 (N_36657,N_36392,N_36381);
or U36658 (N_36658,N_36432,N_36365);
nor U36659 (N_36659,N_36283,N_36318);
nor U36660 (N_36660,N_36263,N_36349);
or U36661 (N_36661,N_36431,N_36378);
nor U36662 (N_36662,N_36316,N_36260);
nor U36663 (N_36663,N_36360,N_36333);
or U36664 (N_36664,N_36342,N_36418);
xor U36665 (N_36665,N_36450,N_36272);
and U36666 (N_36666,N_36334,N_36486);
nand U36667 (N_36667,N_36258,N_36330);
nand U36668 (N_36668,N_36286,N_36480);
xnor U36669 (N_36669,N_36470,N_36310);
and U36670 (N_36670,N_36488,N_36362);
nand U36671 (N_36671,N_36343,N_36313);
and U36672 (N_36672,N_36317,N_36319);
xnor U36673 (N_36673,N_36480,N_36434);
nor U36674 (N_36674,N_36483,N_36382);
or U36675 (N_36675,N_36313,N_36414);
or U36676 (N_36676,N_36280,N_36417);
nand U36677 (N_36677,N_36458,N_36378);
nand U36678 (N_36678,N_36299,N_36487);
nor U36679 (N_36679,N_36492,N_36409);
xor U36680 (N_36680,N_36434,N_36346);
xnor U36681 (N_36681,N_36350,N_36313);
xor U36682 (N_36682,N_36439,N_36392);
or U36683 (N_36683,N_36428,N_36361);
nor U36684 (N_36684,N_36448,N_36298);
or U36685 (N_36685,N_36442,N_36301);
and U36686 (N_36686,N_36296,N_36321);
or U36687 (N_36687,N_36485,N_36276);
and U36688 (N_36688,N_36276,N_36414);
nor U36689 (N_36689,N_36439,N_36259);
or U36690 (N_36690,N_36482,N_36294);
and U36691 (N_36691,N_36252,N_36439);
or U36692 (N_36692,N_36419,N_36404);
nor U36693 (N_36693,N_36391,N_36448);
xnor U36694 (N_36694,N_36301,N_36324);
or U36695 (N_36695,N_36359,N_36310);
or U36696 (N_36696,N_36471,N_36363);
xnor U36697 (N_36697,N_36472,N_36295);
xnor U36698 (N_36698,N_36387,N_36434);
nand U36699 (N_36699,N_36485,N_36422);
nor U36700 (N_36700,N_36471,N_36278);
nand U36701 (N_36701,N_36263,N_36261);
nor U36702 (N_36702,N_36453,N_36388);
nand U36703 (N_36703,N_36376,N_36447);
nand U36704 (N_36704,N_36347,N_36266);
nor U36705 (N_36705,N_36437,N_36349);
nand U36706 (N_36706,N_36493,N_36292);
or U36707 (N_36707,N_36296,N_36376);
nand U36708 (N_36708,N_36259,N_36322);
nand U36709 (N_36709,N_36291,N_36468);
xnor U36710 (N_36710,N_36347,N_36408);
and U36711 (N_36711,N_36464,N_36261);
or U36712 (N_36712,N_36437,N_36276);
nand U36713 (N_36713,N_36400,N_36357);
nor U36714 (N_36714,N_36367,N_36382);
and U36715 (N_36715,N_36386,N_36332);
or U36716 (N_36716,N_36254,N_36284);
nand U36717 (N_36717,N_36339,N_36389);
nor U36718 (N_36718,N_36391,N_36414);
xor U36719 (N_36719,N_36487,N_36348);
xnor U36720 (N_36720,N_36293,N_36378);
and U36721 (N_36721,N_36299,N_36462);
and U36722 (N_36722,N_36366,N_36485);
xor U36723 (N_36723,N_36338,N_36395);
xnor U36724 (N_36724,N_36374,N_36389);
nand U36725 (N_36725,N_36438,N_36408);
nand U36726 (N_36726,N_36398,N_36258);
and U36727 (N_36727,N_36263,N_36387);
and U36728 (N_36728,N_36355,N_36325);
nand U36729 (N_36729,N_36344,N_36333);
nand U36730 (N_36730,N_36425,N_36346);
and U36731 (N_36731,N_36352,N_36360);
or U36732 (N_36732,N_36327,N_36394);
nand U36733 (N_36733,N_36428,N_36453);
and U36734 (N_36734,N_36469,N_36289);
xor U36735 (N_36735,N_36454,N_36390);
nor U36736 (N_36736,N_36345,N_36288);
nor U36737 (N_36737,N_36345,N_36370);
or U36738 (N_36738,N_36286,N_36328);
nor U36739 (N_36739,N_36487,N_36369);
nand U36740 (N_36740,N_36343,N_36359);
or U36741 (N_36741,N_36337,N_36450);
and U36742 (N_36742,N_36309,N_36254);
xnor U36743 (N_36743,N_36487,N_36467);
xor U36744 (N_36744,N_36426,N_36314);
nand U36745 (N_36745,N_36279,N_36280);
nor U36746 (N_36746,N_36369,N_36305);
nand U36747 (N_36747,N_36271,N_36466);
and U36748 (N_36748,N_36264,N_36397);
and U36749 (N_36749,N_36440,N_36268);
nor U36750 (N_36750,N_36601,N_36550);
xnor U36751 (N_36751,N_36571,N_36714);
and U36752 (N_36752,N_36628,N_36684);
and U36753 (N_36753,N_36677,N_36686);
xor U36754 (N_36754,N_36653,N_36594);
xor U36755 (N_36755,N_36683,N_36622);
nor U36756 (N_36756,N_36608,N_36685);
or U36757 (N_36757,N_36738,N_36737);
and U36758 (N_36758,N_36717,N_36671);
and U36759 (N_36759,N_36611,N_36740);
xnor U36760 (N_36760,N_36513,N_36690);
or U36761 (N_36761,N_36675,N_36617);
xnor U36762 (N_36762,N_36674,N_36710);
nand U36763 (N_36763,N_36635,N_36544);
nor U36764 (N_36764,N_36521,N_36606);
nor U36765 (N_36765,N_36732,N_36734);
xnor U36766 (N_36766,N_36668,N_36552);
and U36767 (N_36767,N_36657,N_36697);
or U36768 (N_36768,N_36573,N_36565);
and U36769 (N_36769,N_36621,N_36695);
nand U36770 (N_36770,N_36508,N_36620);
nor U36771 (N_36771,N_36649,N_36700);
xor U36772 (N_36772,N_36560,N_36665);
and U36773 (N_36773,N_36587,N_36520);
nand U36774 (N_36774,N_36575,N_36637);
nand U36775 (N_36775,N_36626,N_36512);
nand U36776 (N_36776,N_36563,N_36669);
nand U36777 (N_36777,N_36543,N_36569);
xor U36778 (N_36778,N_36527,N_36539);
xor U36779 (N_36779,N_36519,N_36701);
xnor U36780 (N_36780,N_36647,N_36748);
or U36781 (N_36781,N_36591,N_36522);
xor U36782 (N_36782,N_36676,N_36625);
and U36783 (N_36783,N_36578,N_36613);
xnor U36784 (N_36784,N_36659,N_36707);
nand U36785 (N_36785,N_36615,N_36724);
nor U36786 (N_36786,N_36561,N_36517);
nand U36787 (N_36787,N_36504,N_36553);
xnor U36788 (N_36788,N_36627,N_36693);
and U36789 (N_36789,N_36632,N_36688);
nor U36790 (N_36790,N_36722,N_36631);
nor U36791 (N_36791,N_36534,N_36548);
or U36792 (N_36792,N_36689,N_36730);
or U36793 (N_36793,N_36554,N_36597);
or U36794 (N_36794,N_36535,N_36630);
and U36795 (N_36795,N_36579,N_36696);
and U36796 (N_36796,N_36698,N_36602);
and U36797 (N_36797,N_36633,N_36680);
nand U36798 (N_36798,N_36589,N_36540);
xor U36799 (N_36799,N_36682,N_36514);
nand U36800 (N_36800,N_36741,N_36726);
xor U36801 (N_36801,N_36727,N_36725);
or U36802 (N_36802,N_36557,N_36749);
or U36803 (N_36803,N_36663,N_36547);
nand U36804 (N_36804,N_36618,N_36619);
nand U36805 (N_36805,N_36712,N_36533);
nand U36806 (N_36806,N_36501,N_36716);
nor U36807 (N_36807,N_36546,N_36654);
xor U36808 (N_36808,N_36744,N_36624);
nand U36809 (N_36809,N_36721,N_36559);
and U36810 (N_36810,N_36541,N_36582);
and U36811 (N_36811,N_36596,N_36564);
nor U36812 (N_36812,N_36545,N_36593);
or U36813 (N_36813,N_36703,N_36584);
nand U36814 (N_36814,N_36645,N_36708);
and U36815 (N_36815,N_36572,N_36644);
xor U36816 (N_36816,N_36523,N_36656);
xnor U36817 (N_36817,N_36590,N_36581);
xnor U36818 (N_36818,N_36713,N_36576);
nand U36819 (N_36819,N_36664,N_36706);
or U36820 (N_36820,N_36640,N_36530);
xnor U36821 (N_36821,N_36542,N_36711);
or U36822 (N_36822,N_36537,N_36643);
and U36823 (N_36823,N_36729,N_36610);
nand U36824 (N_36824,N_36648,N_36516);
nor U36825 (N_36825,N_36743,N_36646);
or U36826 (N_36826,N_36662,N_36655);
or U36827 (N_36827,N_36658,N_36719);
and U36828 (N_36828,N_36679,N_36673);
and U36829 (N_36829,N_36667,N_36642);
nor U36830 (N_36830,N_36702,N_36623);
and U36831 (N_36831,N_36506,N_36709);
nor U36832 (N_36832,N_36636,N_36574);
and U36833 (N_36833,N_36718,N_36670);
or U36834 (N_36834,N_36507,N_36598);
nor U36835 (N_36835,N_36531,N_36583);
or U36836 (N_36836,N_36692,N_36605);
and U36837 (N_36837,N_36604,N_36733);
xor U36838 (N_36838,N_36705,N_36715);
or U36839 (N_36839,N_36629,N_36528);
nand U36840 (N_36840,N_36588,N_36525);
and U36841 (N_36841,N_36551,N_36731);
or U36842 (N_36842,N_36687,N_36699);
xor U36843 (N_36843,N_36652,N_36566);
and U36844 (N_36844,N_36612,N_36568);
xor U36845 (N_36845,N_36746,N_36651);
nor U36846 (N_36846,N_36529,N_36728);
xnor U36847 (N_36847,N_36500,N_36577);
nand U36848 (N_36848,N_36595,N_36704);
or U36849 (N_36849,N_36720,N_36502);
or U36850 (N_36850,N_36641,N_36607);
nor U36851 (N_36851,N_36660,N_36723);
or U36852 (N_36852,N_36599,N_36678);
xnor U36853 (N_36853,N_36614,N_36558);
and U36854 (N_36854,N_36538,N_36515);
xnor U36855 (N_36855,N_36616,N_36585);
and U36856 (N_36856,N_36634,N_36609);
xor U36857 (N_36857,N_36639,N_36567);
nor U36858 (N_36858,N_36526,N_36736);
or U36859 (N_36859,N_36739,N_36518);
xor U36860 (N_36860,N_36532,N_36661);
xnor U36861 (N_36861,N_36556,N_36681);
xor U36862 (N_36862,N_36509,N_36650);
or U36863 (N_36863,N_36549,N_36510);
nor U36864 (N_36864,N_36742,N_36600);
or U36865 (N_36865,N_36603,N_36592);
or U36866 (N_36866,N_36691,N_36666);
nand U36867 (N_36867,N_36672,N_36586);
or U36868 (N_36868,N_36638,N_36580);
nor U36869 (N_36869,N_36570,N_36735);
nand U36870 (N_36870,N_36524,N_36511);
nand U36871 (N_36871,N_36555,N_36503);
or U36872 (N_36872,N_36562,N_36694);
xor U36873 (N_36873,N_36745,N_36747);
nor U36874 (N_36874,N_36536,N_36505);
and U36875 (N_36875,N_36661,N_36592);
nor U36876 (N_36876,N_36703,N_36517);
and U36877 (N_36877,N_36595,N_36622);
nor U36878 (N_36878,N_36672,N_36502);
nor U36879 (N_36879,N_36553,N_36543);
nor U36880 (N_36880,N_36660,N_36590);
xor U36881 (N_36881,N_36598,N_36645);
nor U36882 (N_36882,N_36613,N_36671);
and U36883 (N_36883,N_36610,N_36503);
or U36884 (N_36884,N_36695,N_36657);
nand U36885 (N_36885,N_36617,N_36724);
or U36886 (N_36886,N_36723,N_36672);
nor U36887 (N_36887,N_36718,N_36508);
or U36888 (N_36888,N_36658,N_36520);
and U36889 (N_36889,N_36531,N_36664);
nand U36890 (N_36890,N_36616,N_36569);
or U36891 (N_36891,N_36548,N_36526);
xnor U36892 (N_36892,N_36707,N_36729);
or U36893 (N_36893,N_36549,N_36677);
or U36894 (N_36894,N_36705,N_36532);
and U36895 (N_36895,N_36501,N_36731);
or U36896 (N_36896,N_36711,N_36645);
nand U36897 (N_36897,N_36514,N_36540);
nor U36898 (N_36898,N_36555,N_36721);
xor U36899 (N_36899,N_36539,N_36568);
nand U36900 (N_36900,N_36664,N_36537);
or U36901 (N_36901,N_36650,N_36589);
or U36902 (N_36902,N_36642,N_36553);
nand U36903 (N_36903,N_36512,N_36580);
nor U36904 (N_36904,N_36609,N_36645);
and U36905 (N_36905,N_36551,N_36651);
xor U36906 (N_36906,N_36510,N_36714);
nor U36907 (N_36907,N_36585,N_36684);
nand U36908 (N_36908,N_36693,N_36518);
nand U36909 (N_36909,N_36672,N_36734);
xor U36910 (N_36910,N_36664,N_36629);
xor U36911 (N_36911,N_36522,N_36589);
xor U36912 (N_36912,N_36530,N_36513);
nor U36913 (N_36913,N_36580,N_36691);
or U36914 (N_36914,N_36599,N_36675);
or U36915 (N_36915,N_36730,N_36663);
or U36916 (N_36916,N_36513,N_36728);
nand U36917 (N_36917,N_36616,N_36653);
nor U36918 (N_36918,N_36596,N_36708);
nor U36919 (N_36919,N_36513,N_36599);
nor U36920 (N_36920,N_36634,N_36633);
nand U36921 (N_36921,N_36724,N_36727);
and U36922 (N_36922,N_36729,N_36670);
or U36923 (N_36923,N_36590,N_36553);
xnor U36924 (N_36924,N_36514,N_36645);
nor U36925 (N_36925,N_36743,N_36647);
and U36926 (N_36926,N_36662,N_36549);
or U36927 (N_36927,N_36566,N_36574);
nand U36928 (N_36928,N_36657,N_36723);
xor U36929 (N_36929,N_36563,N_36512);
xnor U36930 (N_36930,N_36541,N_36548);
nor U36931 (N_36931,N_36525,N_36598);
xnor U36932 (N_36932,N_36559,N_36601);
or U36933 (N_36933,N_36640,N_36701);
nand U36934 (N_36934,N_36654,N_36742);
or U36935 (N_36935,N_36623,N_36600);
nor U36936 (N_36936,N_36719,N_36574);
xnor U36937 (N_36937,N_36689,N_36578);
or U36938 (N_36938,N_36686,N_36519);
or U36939 (N_36939,N_36587,N_36624);
or U36940 (N_36940,N_36744,N_36687);
and U36941 (N_36941,N_36746,N_36604);
xor U36942 (N_36942,N_36736,N_36738);
nor U36943 (N_36943,N_36543,N_36551);
nor U36944 (N_36944,N_36718,N_36597);
nand U36945 (N_36945,N_36715,N_36589);
nand U36946 (N_36946,N_36572,N_36693);
and U36947 (N_36947,N_36663,N_36591);
xor U36948 (N_36948,N_36670,N_36663);
and U36949 (N_36949,N_36587,N_36714);
nor U36950 (N_36950,N_36548,N_36725);
nor U36951 (N_36951,N_36518,N_36543);
or U36952 (N_36952,N_36607,N_36565);
or U36953 (N_36953,N_36528,N_36721);
or U36954 (N_36954,N_36682,N_36573);
nor U36955 (N_36955,N_36598,N_36576);
nand U36956 (N_36956,N_36719,N_36542);
or U36957 (N_36957,N_36638,N_36679);
or U36958 (N_36958,N_36653,N_36606);
and U36959 (N_36959,N_36500,N_36682);
nor U36960 (N_36960,N_36559,N_36666);
or U36961 (N_36961,N_36528,N_36675);
xor U36962 (N_36962,N_36607,N_36573);
xnor U36963 (N_36963,N_36576,N_36573);
nand U36964 (N_36964,N_36686,N_36533);
nand U36965 (N_36965,N_36680,N_36561);
xor U36966 (N_36966,N_36717,N_36666);
xnor U36967 (N_36967,N_36620,N_36613);
nand U36968 (N_36968,N_36586,N_36657);
or U36969 (N_36969,N_36548,N_36515);
or U36970 (N_36970,N_36564,N_36550);
nor U36971 (N_36971,N_36680,N_36656);
xnor U36972 (N_36972,N_36667,N_36508);
or U36973 (N_36973,N_36561,N_36508);
or U36974 (N_36974,N_36692,N_36676);
nand U36975 (N_36975,N_36641,N_36626);
and U36976 (N_36976,N_36640,N_36536);
nand U36977 (N_36977,N_36625,N_36503);
or U36978 (N_36978,N_36671,N_36523);
or U36979 (N_36979,N_36521,N_36740);
and U36980 (N_36980,N_36545,N_36621);
xnor U36981 (N_36981,N_36717,N_36509);
nand U36982 (N_36982,N_36679,N_36695);
xor U36983 (N_36983,N_36662,N_36632);
nand U36984 (N_36984,N_36586,N_36741);
nor U36985 (N_36985,N_36589,N_36727);
and U36986 (N_36986,N_36723,N_36636);
nand U36987 (N_36987,N_36742,N_36539);
and U36988 (N_36988,N_36562,N_36551);
nand U36989 (N_36989,N_36721,N_36711);
nand U36990 (N_36990,N_36502,N_36664);
xor U36991 (N_36991,N_36712,N_36529);
nand U36992 (N_36992,N_36707,N_36607);
nand U36993 (N_36993,N_36533,N_36734);
and U36994 (N_36994,N_36593,N_36702);
nand U36995 (N_36995,N_36549,N_36508);
xnor U36996 (N_36996,N_36686,N_36601);
and U36997 (N_36997,N_36713,N_36654);
or U36998 (N_36998,N_36658,N_36512);
nor U36999 (N_36999,N_36593,N_36563);
and U37000 (N_37000,N_36788,N_36836);
or U37001 (N_37001,N_36781,N_36909);
and U37002 (N_37002,N_36897,N_36921);
or U37003 (N_37003,N_36879,N_36859);
nor U37004 (N_37004,N_36850,N_36922);
xnor U37005 (N_37005,N_36794,N_36901);
nor U37006 (N_37006,N_36840,N_36929);
nor U37007 (N_37007,N_36967,N_36905);
nand U37008 (N_37008,N_36977,N_36946);
xor U37009 (N_37009,N_36894,N_36777);
nand U37010 (N_37010,N_36959,N_36970);
xor U37011 (N_37011,N_36899,N_36933);
nand U37012 (N_37012,N_36838,N_36751);
nor U37013 (N_37013,N_36934,N_36754);
and U37014 (N_37014,N_36883,N_36942);
nand U37015 (N_37015,N_36990,N_36862);
nand U37016 (N_37016,N_36795,N_36957);
or U37017 (N_37017,N_36891,N_36952);
nand U37018 (N_37018,N_36984,N_36848);
xor U37019 (N_37019,N_36855,N_36779);
nor U37020 (N_37020,N_36837,N_36821);
xor U37021 (N_37021,N_36902,N_36780);
and U37022 (N_37022,N_36976,N_36756);
nor U37023 (N_37023,N_36808,N_36907);
or U37024 (N_37024,N_36962,N_36864);
and U37025 (N_37025,N_36960,N_36982);
nand U37026 (N_37026,N_36896,N_36940);
or U37027 (N_37027,N_36928,N_36988);
or U37028 (N_37028,N_36853,N_36812);
nor U37029 (N_37029,N_36983,N_36965);
or U37030 (N_37030,N_36820,N_36816);
nand U37031 (N_37031,N_36852,N_36886);
and U37032 (N_37032,N_36866,N_36893);
or U37033 (N_37033,N_36935,N_36923);
nor U37034 (N_37034,N_36870,N_36802);
nor U37035 (N_37035,N_36760,N_36937);
nor U37036 (N_37036,N_36955,N_36904);
xor U37037 (N_37037,N_36775,N_36813);
xor U37038 (N_37038,N_36771,N_36767);
or U37039 (N_37039,N_36986,N_36787);
xnor U37040 (N_37040,N_36772,N_36755);
nand U37041 (N_37041,N_36969,N_36898);
or U37042 (N_37042,N_36919,N_36763);
and U37043 (N_37043,N_36811,N_36791);
xnor U37044 (N_37044,N_36931,N_36951);
nor U37045 (N_37045,N_36911,N_36809);
nand U37046 (N_37046,N_36880,N_36915);
nor U37047 (N_37047,N_36930,N_36861);
and U37048 (N_37048,N_36810,N_36953);
and U37049 (N_37049,N_36949,N_36968);
nand U37050 (N_37050,N_36826,N_36914);
nor U37051 (N_37051,N_36993,N_36818);
nor U37052 (N_37052,N_36770,N_36888);
xor U37053 (N_37053,N_36871,N_36844);
and U37054 (N_37054,N_36819,N_36956);
nor U37055 (N_37055,N_36798,N_36964);
nand U37056 (N_37056,N_36989,N_36801);
and U37057 (N_37057,N_36858,N_36831);
nand U37058 (N_37058,N_36958,N_36878);
xnor U37059 (N_37059,N_36881,N_36830);
nand U37060 (N_37060,N_36913,N_36804);
or U37061 (N_37061,N_36807,N_36924);
and U37062 (N_37062,N_36884,N_36991);
nand U37063 (N_37063,N_36889,N_36793);
xnor U37064 (N_37064,N_36823,N_36761);
and U37065 (N_37065,N_36774,N_36912);
or U37066 (N_37066,N_36841,N_36789);
nand U37067 (N_37067,N_36786,N_36766);
and U37068 (N_37068,N_36975,N_36857);
xor U37069 (N_37069,N_36764,N_36917);
or U37070 (N_37070,N_36963,N_36803);
or U37071 (N_37071,N_36784,N_36945);
and U37072 (N_37072,N_36918,N_36835);
xnor U37073 (N_37073,N_36900,N_36932);
xnor U37074 (N_37074,N_36948,N_36867);
or U37075 (N_37075,N_36815,N_36938);
nand U37076 (N_37076,N_36790,N_36758);
or U37077 (N_37077,N_36822,N_36797);
xnor U37078 (N_37078,N_36910,N_36842);
and U37079 (N_37079,N_36979,N_36971);
and U37080 (N_37080,N_36849,N_36868);
nand U37081 (N_37081,N_36769,N_36757);
and U37082 (N_37082,N_36863,N_36874);
or U37083 (N_37083,N_36851,N_36806);
or U37084 (N_37084,N_36825,N_36997);
or U37085 (N_37085,N_36752,N_36999);
and U37086 (N_37086,N_36936,N_36994);
nor U37087 (N_37087,N_36865,N_36943);
nand U37088 (N_37088,N_36805,N_36854);
nand U37089 (N_37089,N_36985,N_36765);
nor U37090 (N_37090,N_36890,N_36856);
and U37091 (N_37091,N_36872,N_36973);
xor U37092 (N_37092,N_36814,N_36869);
xnor U37093 (N_37093,N_36980,N_36978);
or U37094 (N_37094,N_36873,N_36882);
nand U37095 (N_37095,N_36753,N_36776);
or U37096 (N_37096,N_36799,N_36783);
nand U37097 (N_37097,N_36992,N_36885);
nor U37098 (N_37098,N_36939,N_36908);
xnor U37099 (N_37099,N_36916,N_36778);
or U37100 (N_37100,N_36839,N_36974);
and U37101 (N_37101,N_36944,N_36876);
and U37102 (N_37102,N_36827,N_36860);
and U37103 (N_37103,N_36954,N_36906);
nor U37104 (N_37104,N_36950,N_36996);
nand U37105 (N_37105,N_36995,N_36824);
xnor U37106 (N_37106,N_36877,N_36966);
and U37107 (N_37107,N_36972,N_36750);
nand U37108 (N_37108,N_36759,N_36895);
nand U37109 (N_37109,N_36828,N_36817);
xor U37110 (N_37110,N_36834,N_36785);
or U37111 (N_37111,N_36773,N_36927);
xnor U37112 (N_37112,N_36875,N_36903);
or U37113 (N_37113,N_36926,N_36768);
nand U37114 (N_37114,N_36845,N_36832);
nand U37115 (N_37115,N_36847,N_36920);
nor U37116 (N_37116,N_36843,N_36846);
xor U37117 (N_37117,N_36800,N_36961);
nor U37118 (N_37118,N_36925,N_36981);
xor U37119 (N_37119,N_36887,N_36941);
nor U37120 (N_37120,N_36998,N_36987);
nor U37121 (N_37121,N_36782,N_36947);
and U37122 (N_37122,N_36892,N_36792);
nand U37123 (N_37123,N_36796,N_36762);
nor U37124 (N_37124,N_36829,N_36833);
xor U37125 (N_37125,N_36851,N_36977);
xor U37126 (N_37126,N_36864,N_36937);
xnor U37127 (N_37127,N_36965,N_36942);
and U37128 (N_37128,N_36954,N_36923);
xor U37129 (N_37129,N_36923,N_36961);
or U37130 (N_37130,N_36922,N_36758);
or U37131 (N_37131,N_36839,N_36754);
xor U37132 (N_37132,N_36997,N_36967);
or U37133 (N_37133,N_36752,N_36940);
xor U37134 (N_37134,N_36858,N_36886);
nor U37135 (N_37135,N_36775,N_36790);
xor U37136 (N_37136,N_36901,N_36810);
or U37137 (N_37137,N_36808,N_36879);
xor U37138 (N_37138,N_36982,N_36808);
or U37139 (N_37139,N_36919,N_36868);
nand U37140 (N_37140,N_36898,N_36869);
and U37141 (N_37141,N_36969,N_36899);
nand U37142 (N_37142,N_36808,N_36766);
xnor U37143 (N_37143,N_36977,N_36961);
and U37144 (N_37144,N_36932,N_36936);
xor U37145 (N_37145,N_36836,N_36782);
nand U37146 (N_37146,N_36918,N_36956);
nand U37147 (N_37147,N_36958,N_36948);
and U37148 (N_37148,N_36987,N_36755);
or U37149 (N_37149,N_36895,N_36988);
or U37150 (N_37150,N_36819,N_36790);
xor U37151 (N_37151,N_36892,N_36771);
xnor U37152 (N_37152,N_36820,N_36759);
nor U37153 (N_37153,N_36902,N_36798);
or U37154 (N_37154,N_36786,N_36900);
nor U37155 (N_37155,N_36830,N_36859);
nand U37156 (N_37156,N_36849,N_36782);
or U37157 (N_37157,N_36824,N_36988);
nand U37158 (N_37158,N_36770,N_36776);
xor U37159 (N_37159,N_36752,N_36789);
nor U37160 (N_37160,N_36847,N_36902);
or U37161 (N_37161,N_36760,N_36923);
xor U37162 (N_37162,N_36994,N_36964);
and U37163 (N_37163,N_36984,N_36918);
nand U37164 (N_37164,N_36913,N_36982);
and U37165 (N_37165,N_36874,N_36892);
nand U37166 (N_37166,N_36904,N_36817);
and U37167 (N_37167,N_36796,N_36963);
xnor U37168 (N_37168,N_36888,N_36930);
nor U37169 (N_37169,N_36880,N_36758);
nand U37170 (N_37170,N_36785,N_36867);
nand U37171 (N_37171,N_36775,N_36859);
xnor U37172 (N_37172,N_36817,N_36987);
nand U37173 (N_37173,N_36774,N_36857);
or U37174 (N_37174,N_36819,N_36914);
nor U37175 (N_37175,N_36812,N_36880);
xnor U37176 (N_37176,N_36834,N_36998);
xnor U37177 (N_37177,N_36875,N_36822);
or U37178 (N_37178,N_36792,N_36763);
and U37179 (N_37179,N_36934,N_36790);
nand U37180 (N_37180,N_36785,N_36789);
nor U37181 (N_37181,N_36996,N_36905);
or U37182 (N_37182,N_36913,N_36936);
or U37183 (N_37183,N_36958,N_36830);
or U37184 (N_37184,N_36947,N_36766);
or U37185 (N_37185,N_36989,N_36886);
xor U37186 (N_37186,N_36752,N_36872);
and U37187 (N_37187,N_36894,N_36814);
xor U37188 (N_37188,N_36917,N_36955);
nand U37189 (N_37189,N_36954,N_36878);
nand U37190 (N_37190,N_36805,N_36888);
xnor U37191 (N_37191,N_36967,N_36806);
or U37192 (N_37192,N_36980,N_36795);
nand U37193 (N_37193,N_36810,N_36948);
nand U37194 (N_37194,N_36887,N_36803);
nor U37195 (N_37195,N_36780,N_36899);
nand U37196 (N_37196,N_36965,N_36800);
or U37197 (N_37197,N_36826,N_36964);
or U37198 (N_37198,N_36856,N_36829);
and U37199 (N_37199,N_36930,N_36935);
nor U37200 (N_37200,N_36974,N_36854);
nor U37201 (N_37201,N_36861,N_36891);
xnor U37202 (N_37202,N_36890,N_36897);
xor U37203 (N_37203,N_36784,N_36835);
or U37204 (N_37204,N_36793,N_36896);
or U37205 (N_37205,N_36919,N_36997);
nand U37206 (N_37206,N_36946,N_36792);
nor U37207 (N_37207,N_36857,N_36855);
or U37208 (N_37208,N_36975,N_36822);
nor U37209 (N_37209,N_36892,N_36809);
and U37210 (N_37210,N_36842,N_36838);
nand U37211 (N_37211,N_36787,N_36804);
and U37212 (N_37212,N_36873,N_36993);
nand U37213 (N_37213,N_36949,N_36861);
and U37214 (N_37214,N_36976,N_36988);
xnor U37215 (N_37215,N_36890,N_36923);
nand U37216 (N_37216,N_36868,N_36909);
xnor U37217 (N_37217,N_36787,N_36968);
xor U37218 (N_37218,N_36925,N_36847);
or U37219 (N_37219,N_36986,N_36947);
nand U37220 (N_37220,N_36754,N_36824);
nand U37221 (N_37221,N_36804,N_36992);
or U37222 (N_37222,N_36971,N_36854);
xor U37223 (N_37223,N_36919,N_36865);
xor U37224 (N_37224,N_36835,N_36772);
nor U37225 (N_37225,N_36801,N_36911);
xor U37226 (N_37226,N_36902,N_36979);
nor U37227 (N_37227,N_36945,N_36825);
xor U37228 (N_37228,N_36981,N_36961);
xor U37229 (N_37229,N_36857,N_36870);
xor U37230 (N_37230,N_36967,N_36887);
nand U37231 (N_37231,N_36799,N_36985);
nand U37232 (N_37232,N_36780,N_36754);
and U37233 (N_37233,N_36948,N_36980);
and U37234 (N_37234,N_36761,N_36866);
nor U37235 (N_37235,N_36887,N_36764);
or U37236 (N_37236,N_36839,N_36872);
xor U37237 (N_37237,N_36754,N_36975);
nor U37238 (N_37238,N_36792,N_36764);
nor U37239 (N_37239,N_36806,N_36873);
and U37240 (N_37240,N_36815,N_36822);
or U37241 (N_37241,N_36865,N_36880);
nor U37242 (N_37242,N_36796,N_36983);
xnor U37243 (N_37243,N_36825,N_36762);
nor U37244 (N_37244,N_36887,N_36786);
and U37245 (N_37245,N_36866,N_36988);
nor U37246 (N_37246,N_36834,N_36806);
nand U37247 (N_37247,N_36878,N_36911);
nand U37248 (N_37248,N_36797,N_36770);
or U37249 (N_37249,N_36757,N_36765);
nand U37250 (N_37250,N_37166,N_37170);
nand U37251 (N_37251,N_37175,N_37001);
and U37252 (N_37252,N_37173,N_37050);
nor U37253 (N_37253,N_37153,N_37079);
xor U37254 (N_37254,N_37114,N_37220);
xor U37255 (N_37255,N_37201,N_37051);
nand U37256 (N_37256,N_37168,N_37128);
and U37257 (N_37257,N_37010,N_37126);
xor U37258 (N_37258,N_37217,N_37098);
nand U37259 (N_37259,N_37102,N_37228);
nand U37260 (N_37260,N_37149,N_37065);
xor U37261 (N_37261,N_37024,N_37034);
nor U37262 (N_37262,N_37179,N_37009);
or U37263 (N_37263,N_37136,N_37143);
nor U37264 (N_37264,N_37177,N_37124);
or U37265 (N_37265,N_37160,N_37091);
or U37266 (N_37266,N_37020,N_37222);
or U37267 (N_37267,N_37074,N_37142);
or U37268 (N_37268,N_37130,N_37018);
and U37269 (N_37269,N_37071,N_37125);
and U37270 (N_37270,N_37104,N_37185);
xnor U37271 (N_37271,N_37108,N_37209);
xnor U37272 (N_37272,N_37047,N_37033);
nor U37273 (N_37273,N_37238,N_37080);
or U37274 (N_37274,N_37097,N_37200);
and U37275 (N_37275,N_37016,N_37061);
xnor U37276 (N_37276,N_37014,N_37094);
nand U37277 (N_37277,N_37215,N_37123);
and U37278 (N_37278,N_37239,N_37083);
or U37279 (N_37279,N_37183,N_37150);
nand U37280 (N_37280,N_37187,N_37105);
and U37281 (N_37281,N_37169,N_37205);
and U37282 (N_37282,N_37146,N_37129);
nor U37283 (N_37283,N_37022,N_37006);
nor U37284 (N_37284,N_37062,N_37219);
nor U37285 (N_37285,N_37172,N_37158);
and U37286 (N_37286,N_37147,N_37140);
and U37287 (N_37287,N_37037,N_37015);
nand U37288 (N_37288,N_37161,N_37157);
and U37289 (N_37289,N_37087,N_37188);
xor U37290 (N_37290,N_37145,N_37095);
xor U37291 (N_37291,N_37133,N_37052);
xor U37292 (N_37292,N_37107,N_37197);
xor U37293 (N_37293,N_37196,N_37237);
and U37294 (N_37294,N_37029,N_37093);
xor U37295 (N_37295,N_37035,N_37084);
and U37296 (N_37296,N_37089,N_37182);
xor U37297 (N_37297,N_37132,N_37085);
or U37298 (N_37298,N_37243,N_37163);
or U37299 (N_37299,N_37151,N_37101);
and U37300 (N_37300,N_37195,N_37206);
nor U37301 (N_37301,N_37106,N_37059);
xnor U37302 (N_37302,N_37000,N_37152);
and U37303 (N_37303,N_37025,N_37218);
nand U37304 (N_37304,N_37072,N_37230);
nand U37305 (N_37305,N_37224,N_37223);
or U37306 (N_37306,N_37139,N_37077);
nand U37307 (N_37307,N_37180,N_37056);
and U37308 (N_37308,N_37210,N_37075);
xnor U37309 (N_37309,N_37086,N_37067);
nand U37310 (N_37310,N_37171,N_37088);
xor U37311 (N_37311,N_37144,N_37235);
or U37312 (N_37312,N_37127,N_37057);
nor U37313 (N_37313,N_37135,N_37023);
and U37314 (N_37314,N_37043,N_37227);
and U37315 (N_37315,N_37026,N_37194);
or U37316 (N_37316,N_37100,N_37045);
or U37317 (N_37317,N_37007,N_37005);
or U37318 (N_37318,N_37245,N_37027);
and U37319 (N_37319,N_37081,N_37120);
nand U37320 (N_37320,N_37221,N_37028);
or U37321 (N_37321,N_37110,N_37049);
or U37322 (N_37322,N_37092,N_37058);
or U37323 (N_37323,N_37113,N_37040);
xnor U37324 (N_37324,N_37240,N_37032);
nand U37325 (N_37325,N_37116,N_37162);
nor U37326 (N_37326,N_37031,N_37207);
nand U37327 (N_37327,N_37190,N_37021);
xnor U37328 (N_37328,N_37193,N_37041);
and U37329 (N_37329,N_37118,N_37036);
or U37330 (N_37330,N_37122,N_37233);
and U37331 (N_37331,N_37076,N_37068);
or U37332 (N_37332,N_37241,N_37138);
and U37333 (N_37333,N_37246,N_37191);
or U37334 (N_37334,N_37042,N_37174);
nand U37335 (N_37335,N_37017,N_37167);
nand U37336 (N_37336,N_37204,N_37211);
nand U37337 (N_37337,N_37244,N_37069);
nand U37338 (N_37338,N_37054,N_37082);
nand U37339 (N_37339,N_37159,N_37198);
or U37340 (N_37340,N_37156,N_37231);
nor U37341 (N_37341,N_37039,N_37066);
or U37342 (N_37342,N_37060,N_37214);
xnor U37343 (N_37343,N_37013,N_37019);
and U37344 (N_37344,N_37008,N_37121);
nor U37345 (N_37345,N_37148,N_37112);
or U37346 (N_37346,N_37248,N_37225);
and U37347 (N_37347,N_37096,N_37055);
nand U37348 (N_37348,N_37099,N_37109);
nand U37349 (N_37349,N_37053,N_37137);
or U37350 (N_37350,N_37063,N_37213);
xnor U37351 (N_37351,N_37119,N_37134);
and U37352 (N_37352,N_37002,N_37003);
xor U37353 (N_37353,N_37154,N_37046);
nand U37354 (N_37354,N_37189,N_37178);
or U37355 (N_37355,N_37090,N_37155);
nor U37356 (N_37356,N_37186,N_37199);
and U37357 (N_37357,N_37111,N_37216);
or U37358 (N_37358,N_37249,N_37011);
nor U37359 (N_37359,N_37073,N_37004);
nand U37360 (N_37360,N_37038,N_37203);
xnor U37361 (N_37361,N_37131,N_37184);
and U37362 (N_37362,N_37064,N_37048);
or U37363 (N_37363,N_37012,N_37070);
and U37364 (N_37364,N_37234,N_37078);
xor U37365 (N_37365,N_37202,N_37044);
xnor U37366 (N_37366,N_37164,N_37103);
nand U37367 (N_37367,N_37232,N_37141);
nor U37368 (N_37368,N_37165,N_37176);
and U37369 (N_37369,N_37030,N_37192);
xor U37370 (N_37370,N_37229,N_37212);
or U37371 (N_37371,N_37117,N_37247);
nor U37372 (N_37372,N_37208,N_37236);
xor U37373 (N_37373,N_37115,N_37226);
xnor U37374 (N_37374,N_37242,N_37181);
nand U37375 (N_37375,N_37242,N_37172);
xor U37376 (N_37376,N_37107,N_37217);
xnor U37377 (N_37377,N_37224,N_37084);
nor U37378 (N_37378,N_37063,N_37111);
nand U37379 (N_37379,N_37244,N_37097);
xor U37380 (N_37380,N_37032,N_37209);
or U37381 (N_37381,N_37164,N_37019);
nand U37382 (N_37382,N_37165,N_37212);
or U37383 (N_37383,N_37137,N_37081);
or U37384 (N_37384,N_37224,N_37003);
and U37385 (N_37385,N_37119,N_37099);
or U37386 (N_37386,N_37225,N_37023);
nand U37387 (N_37387,N_37035,N_37243);
nor U37388 (N_37388,N_37050,N_37141);
nand U37389 (N_37389,N_37133,N_37069);
or U37390 (N_37390,N_37082,N_37140);
xor U37391 (N_37391,N_37166,N_37204);
nor U37392 (N_37392,N_37135,N_37018);
nor U37393 (N_37393,N_37055,N_37003);
nor U37394 (N_37394,N_37049,N_37034);
xor U37395 (N_37395,N_37039,N_37236);
nor U37396 (N_37396,N_37223,N_37085);
and U37397 (N_37397,N_37091,N_37054);
nor U37398 (N_37398,N_37002,N_37083);
xor U37399 (N_37399,N_37195,N_37029);
or U37400 (N_37400,N_37039,N_37099);
xnor U37401 (N_37401,N_37047,N_37090);
or U37402 (N_37402,N_37066,N_37160);
xor U37403 (N_37403,N_37154,N_37089);
nor U37404 (N_37404,N_37181,N_37038);
and U37405 (N_37405,N_37227,N_37139);
xor U37406 (N_37406,N_37071,N_37130);
nand U37407 (N_37407,N_37083,N_37156);
and U37408 (N_37408,N_37111,N_37039);
nand U37409 (N_37409,N_37018,N_37065);
nor U37410 (N_37410,N_37070,N_37180);
or U37411 (N_37411,N_37169,N_37019);
and U37412 (N_37412,N_37205,N_37070);
nor U37413 (N_37413,N_37073,N_37123);
nor U37414 (N_37414,N_37009,N_37122);
nand U37415 (N_37415,N_37092,N_37093);
xor U37416 (N_37416,N_37159,N_37089);
nor U37417 (N_37417,N_37204,N_37203);
xor U37418 (N_37418,N_37092,N_37066);
nand U37419 (N_37419,N_37124,N_37222);
xor U37420 (N_37420,N_37197,N_37113);
xor U37421 (N_37421,N_37018,N_37053);
or U37422 (N_37422,N_37213,N_37120);
and U37423 (N_37423,N_37113,N_37139);
or U37424 (N_37424,N_37133,N_37139);
and U37425 (N_37425,N_37195,N_37218);
nor U37426 (N_37426,N_37195,N_37197);
or U37427 (N_37427,N_37161,N_37129);
xor U37428 (N_37428,N_37188,N_37169);
nor U37429 (N_37429,N_37037,N_37234);
nor U37430 (N_37430,N_37111,N_37080);
or U37431 (N_37431,N_37225,N_37175);
nand U37432 (N_37432,N_37115,N_37036);
xnor U37433 (N_37433,N_37152,N_37010);
nand U37434 (N_37434,N_37032,N_37239);
and U37435 (N_37435,N_37089,N_37004);
nand U37436 (N_37436,N_37195,N_37140);
xor U37437 (N_37437,N_37067,N_37029);
xor U37438 (N_37438,N_37133,N_37115);
xor U37439 (N_37439,N_37229,N_37219);
nor U37440 (N_37440,N_37240,N_37236);
nand U37441 (N_37441,N_37188,N_37118);
nor U37442 (N_37442,N_37178,N_37075);
nand U37443 (N_37443,N_37139,N_37210);
nor U37444 (N_37444,N_37238,N_37216);
nand U37445 (N_37445,N_37041,N_37154);
and U37446 (N_37446,N_37087,N_37169);
nor U37447 (N_37447,N_37216,N_37054);
nor U37448 (N_37448,N_37160,N_37051);
nor U37449 (N_37449,N_37228,N_37005);
xor U37450 (N_37450,N_37210,N_37017);
or U37451 (N_37451,N_37206,N_37156);
nand U37452 (N_37452,N_37076,N_37072);
and U37453 (N_37453,N_37096,N_37134);
nor U37454 (N_37454,N_37109,N_37058);
or U37455 (N_37455,N_37221,N_37180);
and U37456 (N_37456,N_37112,N_37150);
and U37457 (N_37457,N_37107,N_37127);
and U37458 (N_37458,N_37083,N_37070);
and U37459 (N_37459,N_37174,N_37241);
nor U37460 (N_37460,N_37193,N_37222);
xor U37461 (N_37461,N_37093,N_37205);
nor U37462 (N_37462,N_37217,N_37197);
nor U37463 (N_37463,N_37069,N_37057);
and U37464 (N_37464,N_37113,N_37073);
nor U37465 (N_37465,N_37188,N_37174);
nor U37466 (N_37466,N_37049,N_37162);
nor U37467 (N_37467,N_37164,N_37026);
and U37468 (N_37468,N_37215,N_37120);
nand U37469 (N_37469,N_37016,N_37219);
and U37470 (N_37470,N_37074,N_37054);
xnor U37471 (N_37471,N_37124,N_37076);
nor U37472 (N_37472,N_37185,N_37220);
nor U37473 (N_37473,N_37037,N_37031);
or U37474 (N_37474,N_37044,N_37102);
nor U37475 (N_37475,N_37181,N_37043);
nand U37476 (N_37476,N_37048,N_37248);
or U37477 (N_37477,N_37016,N_37213);
nand U37478 (N_37478,N_37089,N_37206);
and U37479 (N_37479,N_37208,N_37018);
nor U37480 (N_37480,N_37182,N_37042);
and U37481 (N_37481,N_37196,N_37105);
nor U37482 (N_37482,N_37242,N_37117);
nor U37483 (N_37483,N_37091,N_37050);
and U37484 (N_37484,N_37155,N_37006);
nor U37485 (N_37485,N_37139,N_37224);
xnor U37486 (N_37486,N_37222,N_37170);
nand U37487 (N_37487,N_37220,N_37247);
nor U37488 (N_37488,N_37000,N_37183);
nand U37489 (N_37489,N_37164,N_37191);
nand U37490 (N_37490,N_37038,N_37097);
nand U37491 (N_37491,N_37039,N_37175);
or U37492 (N_37492,N_37169,N_37015);
nand U37493 (N_37493,N_37045,N_37243);
xor U37494 (N_37494,N_37024,N_37022);
and U37495 (N_37495,N_37048,N_37154);
nor U37496 (N_37496,N_37048,N_37216);
xnor U37497 (N_37497,N_37247,N_37208);
and U37498 (N_37498,N_37056,N_37120);
nor U37499 (N_37499,N_37070,N_37148);
nand U37500 (N_37500,N_37287,N_37401);
xor U37501 (N_37501,N_37342,N_37369);
xor U37502 (N_37502,N_37368,N_37371);
xor U37503 (N_37503,N_37468,N_37402);
nor U37504 (N_37504,N_37323,N_37400);
and U37505 (N_37505,N_37357,N_37376);
nor U37506 (N_37506,N_37485,N_37335);
nand U37507 (N_37507,N_37333,N_37378);
or U37508 (N_37508,N_37326,N_37263);
xor U37509 (N_37509,N_37275,N_37288);
nand U37510 (N_37510,N_37447,N_37470);
and U37511 (N_37511,N_37346,N_37487);
nor U37512 (N_37512,N_37471,N_37435);
nor U37513 (N_37513,N_37334,N_37386);
nor U37514 (N_37514,N_37458,N_37367);
nand U37515 (N_37515,N_37395,N_37441);
xor U37516 (N_37516,N_37261,N_37362);
nand U37517 (N_37517,N_37469,N_37492);
nand U37518 (N_37518,N_37297,N_37459);
or U37519 (N_37519,N_37310,N_37457);
nand U37520 (N_37520,N_37390,N_37494);
xnor U37521 (N_37521,N_37432,N_37350);
nor U37522 (N_37522,N_37489,N_37405);
xor U37523 (N_37523,N_37354,N_37394);
or U37524 (N_37524,N_37324,N_37317);
nand U37525 (N_37525,N_37497,N_37416);
nand U37526 (N_37526,N_37407,N_37271);
or U37527 (N_37527,N_37391,N_37437);
or U37528 (N_37528,N_37251,N_37296);
nor U37529 (N_37529,N_37365,N_37482);
or U37530 (N_37530,N_37414,N_37294);
xnor U37531 (N_37531,N_37498,N_37388);
or U37532 (N_37532,N_37383,N_37270);
xnor U37533 (N_37533,N_37257,N_37421);
nand U37534 (N_37534,N_37403,N_37284);
xor U37535 (N_37535,N_37360,N_37477);
nand U37536 (N_37536,N_37439,N_37499);
nor U37537 (N_37537,N_37266,N_37277);
nand U37538 (N_37538,N_37313,N_37254);
nand U37539 (N_37539,N_37472,N_37344);
xnor U37540 (N_37540,N_37483,N_37281);
xnor U37541 (N_37541,N_37486,N_37348);
nand U37542 (N_37542,N_37260,N_37349);
xnor U37543 (N_37543,N_37495,N_37479);
nand U37544 (N_37544,N_37409,N_37375);
xor U37545 (N_37545,N_37268,N_37279);
nand U37546 (N_37546,N_37474,N_37436);
or U37547 (N_37547,N_37422,N_37370);
and U37548 (N_37548,N_37444,N_37273);
and U37549 (N_37549,N_37373,N_37314);
or U37550 (N_37550,N_37475,N_37345);
or U37551 (N_37551,N_37265,N_37452);
xor U37552 (N_37552,N_37253,N_37358);
and U37553 (N_37553,N_37473,N_37456);
nor U37554 (N_37554,N_37425,N_37319);
nand U37555 (N_37555,N_37276,N_37262);
xnor U37556 (N_37556,N_37478,N_37359);
nor U37557 (N_37557,N_37430,N_37413);
nand U37558 (N_37558,N_37476,N_37488);
nor U37559 (N_37559,N_37330,N_37351);
and U37560 (N_37560,N_37293,N_37454);
nor U37561 (N_37561,N_37321,N_37315);
or U37562 (N_37562,N_37418,N_37340);
or U37563 (N_37563,N_37372,N_37466);
and U37564 (N_37564,N_37496,N_37366);
and U37565 (N_37565,N_37312,N_37434);
xor U37566 (N_37566,N_37460,N_37338);
xnor U37567 (N_37567,N_37289,N_37406);
and U37568 (N_37568,N_37404,N_37309);
or U37569 (N_37569,N_37264,N_37387);
nand U37570 (N_37570,N_37399,N_37461);
nand U37571 (N_37571,N_37355,N_37448);
nor U37572 (N_37572,N_37412,N_37290);
or U37573 (N_37573,N_37361,N_37303);
or U37574 (N_37574,N_37337,N_37385);
nor U37575 (N_37575,N_37252,N_37347);
or U37576 (N_37576,N_37327,N_37480);
and U37577 (N_37577,N_37446,N_37256);
and U37578 (N_37578,N_37305,N_37462);
nand U37579 (N_37579,N_37481,N_37322);
or U37580 (N_37580,N_37339,N_37298);
nand U37581 (N_37581,N_37427,N_37286);
xor U37582 (N_37582,N_37445,N_37274);
xor U37583 (N_37583,N_37397,N_37301);
and U37584 (N_37584,N_37374,N_37396);
or U37585 (N_37585,N_37299,N_37398);
nand U37586 (N_37586,N_37484,N_37311);
xor U37587 (N_37587,N_37295,N_37415);
nand U37588 (N_37588,N_37258,N_37491);
or U37589 (N_37589,N_37438,N_37442);
and U37590 (N_37590,N_37431,N_37331);
or U37591 (N_37591,N_37352,N_37308);
nor U37592 (N_37592,N_37463,N_37449);
nor U37593 (N_37593,N_37267,N_37420);
nand U37594 (N_37594,N_37408,N_37364);
xnor U37595 (N_37595,N_37259,N_37329);
xnor U37596 (N_37596,N_37363,N_37332);
and U37597 (N_37597,N_37316,N_37419);
and U37598 (N_37598,N_37451,N_37379);
and U37599 (N_37599,N_37307,N_37389);
nor U37600 (N_37600,N_37380,N_37353);
or U37601 (N_37601,N_37467,N_37343);
nand U37602 (N_37602,N_37382,N_37411);
and U37603 (N_37603,N_37443,N_37280);
nor U37604 (N_37604,N_37285,N_37490);
nand U37605 (N_37605,N_37250,N_37306);
nand U37606 (N_37606,N_37393,N_37304);
and U37607 (N_37607,N_37450,N_37328);
xnor U37608 (N_37608,N_37377,N_37428);
nand U37609 (N_37609,N_37336,N_37384);
nor U37610 (N_37610,N_37278,N_37392);
nor U37611 (N_37611,N_37455,N_37341);
xnor U37612 (N_37612,N_37493,N_37283);
xnor U37613 (N_37613,N_37291,N_37417);
nor U37614 (N_37614,N_37464,N_37423);
or U37615 (N_37615,N_37429,N_37272);
nor U37616 (N_37616,N_37325,N_37465);
or U37617 (N_37617,N_37255,N_37410);
or U37618 (N_37618,N_37424,N_37433);
nor U37619 (N_37619,N_37440,N_37453);
and U37620 (N_37620,N_37320,N_37300);
nand U37621 (N_37621,N_37318,N_37426);
and U37622 (N_37622,N_37302,N_37269);
xnor U37623 (N_37623,N_37282,N_37381);
and U37624 (N_37624,N_37356,N_37292);
and U37625 (N_37625,N_37388,N_37378);
and U37626 (N_37626,N_37366,N_37274);
xor U37627 (N_37627,N_37281,N_37442);
and U37628 (N_37628,N_37291,N_37270);
xnor U37629 (N_37629,N_37350,N_37409);
xor U37630 (N_37630,N_37348,N_37318);
nor U37631 (N_37631,N_37427,N_37283);
and U37632 (N_37632,N_37336,N_37438);
and U37633 (N_37633,N_37493,N_37364);
xor U37634 (N_37634,N_37279,N_37295);
xor U37635 (N_37635,N_37397,N_37476);
and U37636 (N_37636,N_37304,N_37454);
or U37637 (N_37637,N_37373,N_37316);
nand U37638 (N_37638,N_37269,N_37275);
and U37639 (N_37639,N_37314,N_37336);
and U37640 (N_37640,N_37458,N_37354);
nand U37641 (N_37641,N_37263,N_37427);
nand U37642 (N_37642,N_37461,N_37498);
nand U37643 (N_37643,N_37398,N_37397);
nand U37644 (N_37644,N_37349,N_37331);
xnor U37645 (N_37645,N_37373,N_37351);
or U37646 (N_37646,N_37380,N_37456);
and U37647 (N_37647,N_37383,N_37257);
and U37648 (N_37648,N_37492,N_37456);
or U37649 (N_37649,N_37451,N_37442);
nand U37650 (N_37650,N_37487,N_37252);
or U37651 (N_37651,N_37363,N_37334);
xnor U37652 (N_37652,N_37474,N_37259);
or U37653 (N_37653,N_37451,N_37358);
nor U37654 (N_37654,N_37364,N_37259);
or U37655 (N_37655,N_37264,N_37440);
and U37656 (N_37656,N_37251,N_37289);
or U37657 (N_37657,N_37370,N_37264);
or U37658 (N_37658,N_37262,N_37441);
nand U37659 (N_37659,N_37298,N_37252);
or U37660 (N_37660,N_37482,N_37382);
xor U37661 (N_37661,N_37302,N_37308);
nand U37662 (N_37662,N_37277,N_37474);
xnor U37663 (N_37663,N_37404,N_37364);
nand U37664 (N_37664,N_37264,N_37355);
nand U37665 (N_37665,N_37365,N_37360);
or U37666 (N_37666,N_37310,N_37322);
nand U37667 (N_37667,N_37471,N_37459);
xor U37668 (N_37668,N_37419,N_37409);
and U37669 (N_37669,N_37292,N_37310);
nand U37670 (N_37670,N_37375,N_37301);
and U37671 (N_37671,N_37494,N_37333);
nor U37672 (N_37672,N_37472,N_37314);
nor U37673 (N_37673,N_37297,N_37492);
nand U37674 (N_37674,N_37429,N_37329);
xnor U37675 (N_37675,N_37334,N_37370);
nor U37676 (N_37676,N_37418,N_37440);
nor U37677 (N_37677,N_37442,N_37476);
nor U37678 (N_37678,N_37333,N_37266);
or U37679 (N_37679,N_37463,N_37370);
xor U37680 (N_37680,N_37255,N_37424);
and U37681 (N_37681,N_37394,N_37333);
nor U37682 (N_37682,N_37418,N_37478);
nor U37683 (N_37683,N_37484,N_37265);
xnor U37684 (N_37684,N_37421,N_37274);
nor U37685 (N_37685,N_37426,N_37298);
and U37686 (N_37686,N_37252,N_37309);
nor U37687 (N_37687,N_37464,N_37340);
and U37688 (N_37688,N_37301,N_37454);
xor U37689 (N_37689,N_37428,N_37342);
and U37690 (N_37690,N_37464,N_37368);
xnor U37691 (N_37691,N_37387,N_37388);
or U37692 (N_37692,N_37376,N_37274);
xnor U37693 (N_37693,N_37416,N_37259);
or U37694 (N_37694,N_37452,N_37380);
and U37695 (N_37695,N_37250,N_37479);
nand U37696 (N_37696,N_37316,N_37478);
nor U37697 (N_37697,N_37483,N_37481);
and U37698 (N_37698,N_37499,N_37471);
nor U37699 (N_37699,N_37286,N_37431);
and U37700 (N_37700,N_37476,N_37432);
or U37701 (N_37701,N_37332,N_37373);
nand U37702 (N_37702,N_37493,N_37308);
nor U37703 (N_37703,N_37410,N_37428);
and U37704 (N_37704,N_37405,N_37301);
nand U37705 (N_37705,N_37460,N_37264);
or U37706 (N_37706,N_37270,N_37314);
or U37707 (N_37707,N_37439,N_37421);
or U37708 (N_37708,N_37392,N_37356);
nor U37709 (N_37709,N_37348,N_37293);
nand U37710 (N_37710,N_37261,N_37395);
xor U37711 (N_37711,N_37288,N_37322);
and U37712 (N_37712,N_37375,N_37383);
nand U37713 (N_37713,N_37324,N_37458);
nor U37714 (N_37714,N_37331,N_37314);
xnor U37715 (N_37715,N_37395,N_37351);
nand U37716 (N_37716,N_37323,N_37294);
xor U37717 (N_37717,N_37470,N_37378);
nand U37718 (N_37718,N_37271,N_37458);
nand U37719 (N_37719,N_37332,N_37266);
and U37720 (N_37720,N_37298,N_37361);
or U37721 (N_37721,N_37379,N_37284);
xnor U37722 (N_37722,N_37253,N_37296);
and U37723 (N_37723,N_37417,N_37423);
nand U37724 (N_37724,N_37448,N_37437);
or U37725 (N_37725,N_37285,N_37399);
and U37726 (N_37726,N_37312,N_37399);
nand U37727 (N_37727,N_37392,N_37439);
xor U37728 (N_37728,N_37290,N_37315);
and U37729 (N_37729,N_37439,N_37374);
nand U37730 (N_37730,N_37489,N_37454);
or U37731 (N_37731,N_37463,N_37438);
xor U37732 (N_37732,N_37480,N_37424);
nand U37733 (N_37733,N_37300,N_37414);
and U37734 (N_37734,N_37259,N_37254);
nor U37735 (N_37735,N_37258,N_37421);
and U37736 (N_37736,N_37255,N_37379);
and U37737 (N_37737,N_37419,N_37339);
nand U37738 (N_37738,N_37379,N_37258);
xor U37739 (N_37739,N_37339,N_37295);
or U37740 (N_37740,N_37460,N_37431);
or U37741 (N_37741,N_37250,N_37254);
or U37742 (N_37742,N_37272,N_37261);
and U37743 (N_37743,N_37380,N_37436);
nor U37744 (N_37744,N_37422,N_37272);
or U37745 (N_37745,N_37414,N_37485);
xor U37746 (N_37746,N_37272,N_37289);
or U37747 (N_37747,N_37403,N_37442);
xor U37748 (N_37748,N_37469,N_37319);
nand U37749 (N_37749,N_37341,N_37442);
and U37750 (N_37750,N_37590,N_37718);
nor U37751 (N_37751,N_37686,N_37715);
or U37752 (N_37752,N_37615,N_37614);
nor U37753 (N_37753,N_37570,N_37719);
or U37754 (N_37754,N_37707,N_37623);
nor U37755 (N_37755,N_37678,N_37542);
xor U37756 (N_37756,N_37717,N_37531);
or U37757 (N_37757,N_37700,N_37647);
and U37758 (N_37758,N_37720,N_37515);
nand U37759 (N_37759,N_37651,N_37706);
nand U37760 (N_37760,N_37714,N_37666);
nor U37761 (N_37761,N_37598,N_37710);
nor U37762 (N_37762,N_37640,N_37600);
or U37763 (N_37763,N_37699,N_37543);
nand U37764 (N_37764,N_37726,N_37596);
or U37765 (N_37765,N_37525,N_37535);
and U37766 (N_37766,N_37549,N_37704);
xnor U37767 (N_37767,N_37695,N_37721);
xnor U37768 (N_37768,N_37561,N_37573);
xnor U37769 (N_37769,N_37737,N_37551);
xnor U37770 (N_37770,N_37635,N_37612);
or U37771 (N_37771,N_37603,N_37519);
and U37772 (N_37772,N_37656,N_37583);
xnor U37773 (N_37773,N_37736,N_37581);
nor U37774 (N_37774,N_37712,N_37601);
nor U37775 (N_37775,N_37526,N_37681);
xnor U37776 (N_37776,N_37709,N_37654);
nor U37777 (N_37777,N_37610,N_37571);
nand U37778 (N_37778,N_37637,N_37741);
and U37779 (N_37779,N_37554,N_37655);
or U37780 (N_37780,N_37547,N_37522);
xnor U37781 (N_37781,N_37611,N_37553);
nand U37782 (N_37782,N_37546,N_37703);
and U37783 (N_37783,N_37684,N_37634);
and U37784 (N_37784,N_37698,N_37577);
or U37785 (N_37785,N_37602,N_37643);
and U37786 (N_37786,N_37722,N_37729);
or U37787 (N_37787,N_37509,N_37680);
xnor U37788 (N_37788,N_37540,N_37731);
nor U37789 (N_37789,N_37727,N_37733);
and U37790 (N_37790,N_37552,N_37557);
nor U37791 (N_37791,N_37550,N_37641);
and U37792 (N_37792,N_37565,N_37742);
nor U37793 (N_37793,N_37625,N_37572);
and U37794 (N_37794,N_37642,N_37576);
nand U37795 (N_37795,N_37595,N_37740);
or U37796 (N_37796,N_37575,N_37677);
nor U37797 (N_37797,N_37597,N_37708);
nor U37798 (N_37798,N_37588,N_37532);
xnor U37799 (N_37799,N_37563,N_37599);
or U37800 (N_37800,N_37728,N_37702);
xor U37801 (N_37801,N_37653,N_37591);
nor U37802 (N_37802,N_37559,N_37616);
nor U37803 (N_37803,N_37613,N_37523);
nor U37804 (N_37804,N_37660,N_37619);
nand U37805 (N_37805,N_37667,N_37620);
and U37806 (N_37806,N_37582,N_37690);
or U37807 (N_37807,N_37569,N_37617);
nor U37808 (N_37808,N_37661,N_37633);
nor U37809 (N_37809,N_37604,N_37606);
and U37810 (N_37810,N_37508,N_37505);
nor U37811 (N_37811,N_37638,N_37669);
nand U37812 (N_37812,N_37734,N_37558);
xor U37813 (N_37813,N_37705,N_37659);
nor U37814 (N_37814,N_37668,N_37608);
and U37815 (N_37815,N_37632,N_37739);
or U37816 (N_37816,N_37511,N_37555);
nor U37817 (N_37817,N_37743,N_37594);
and U37818 (N_37818,N_37744,N_37513);
and U37819 (N_37819,N_37676,N_37748);
or U37820 (N_37820,N_37738,N_37618);
xor U37821 (N_37821,N_37517,N_37512);
nand U37822 (N_37822,N_37504,N_37630);
or U37823 (N_37823,N_37693,N_37538);
or U37824 (N_37824,N_37745,N_37566);
xor U37825 (N_37825,N_37537,N_37567);
nand U37826 (N_37826,N_37645,N_37732);
or U37827 (N_37827,N_37688,N_37541);
xor U37828 (N_37828,N_37545,N_37533);
nand U37829 (N_37829,N_37670,N_37510);
nand U37830 (N_37830,N_37749,N_37539);
or U37831 (N_37831,N_37665,N_37564);
nor U37832 (N_37832,N_37578,N_37725);
nor U37833 (N_37833,N_37521,N_37713);
or U37834 (N_37834,N_37652,N_37674);
or U37835 (N_37835,N_37534,N_37607);
nand U37836 (N_37836,N_37514,N_37664);
nand U37837 (N_37837,N_37548,N_37735);
nor U37838 (N_37838,N_37696,N_37675);
or U37839 (N_37839,N_37692,N_37579);
xor U37840 (N_37840,N_37589,N_37662);
and U37841 (N_37841,N_37568,N_37621);
nand U37842 (N_37842,N_37500,N_37516);
nand U37843 (N_37843,N_37746,N_37502);
nand U37844 (N_37844,N_37530,N_37730);
and U37845 (N_37845,N_37631,N_37747);
xor U37846 (N_37846,N_37679,N_37649);
nand U37847 (N_37847,N_37622,N_37518);
nor U37848 (N_37848,N_37624,N_37574);
nor U37849 (N_37849,N_37501,N_37691);
and U37850 (N_37850,N_37711,N_37689);
and U37851 (N_37851,N_37627,N_37646);
or U37852 (N_37852,N_37560,N_37592);
xor U37853 (N_37853,N_37657,N_37650);
xor U37854 (N_37854,N_37687,N_37609);
or U37855 (N_37855,N_37639,N_37685);
or U37856 (N_37856,N_37644,N_37671);
xnor U37857 (N_37857,N_37701,N_37580);
nor U37858 (N_37858,N_37520,N_37723);
xor U37859 (N_37859,N_37636,N_37586);
xnor U37860 (N_37860,N_37694,N_37562);
or U37861 (N_37861,N_37697,N_37528);
or U37862 (N_37862,N_37663,N_37658);
nor U37863 (N_37863,N_37536,N_37629);
and U37864 (N_37864,N_37556,N_37503);
nor U37865 (N_37865,N_37527,N_37529);
nand U37866 (N_37866,N_37626,N_37673);
and U37867 (N_37867,N_37585,N_37587);
nand U37868 (N_37868,N_37593,N_37716);
and U37869 (N_37869,N_37584,N_37683);
nor U37870 (N_37870,N_37724,N_37648);
and U37871 (N_37871,N_37628,N_37544);
nand U37872 (N_37872,N_37524,N_37682);
nand U37873 (N_37873,N_37507,N_37605);
nor U37874 (N_37874,N_37506,N_37672);
nand U37875 (N_37875,N_37604,N_37561);
nand U37876 (N_37876,N_37519,N_37666);
and U37877 (N_37877,N_37528,N_37609);
nor U37878 (N_37878,N_37634,N_37665);
xnor U37879 (N_37879,N_37737,N_37599);
nor U37880 (N_37880,N_37612,N_37575);
nand U37881 (N_37881,N_37522,N_37617);
nor U37882 (N_37882,N_37660,N_37547);
or U37883 (N_37883,N_37576,N_37731);
nand U37884 (N_37884,N_37599,N_37736);
and U37885 (N_37885,N_37630,N_37662);
or U37886 (N_37886,N_37687,N_37654);
or U37887 (N_37887,N_37590,N_37545);
nand U37888 (N_37888,N_37500,N_37736);
xor U37889 (N_37889,N_37746,N_37683);
or U37890 (N_37890,N_37576,N_37579);
or U37891 (N_37891,N_37719,N_37631);
or U37892 (N_37892,N_37715,N_37660);
nand U37893 (N_37893,N_37649,N_37548);
and U37894 (N_37894,N_37562,N_37728);
nor U37895 (N_37895,N_37553,N_37665);
nand U37896 (N_37896,N_37715,N_37545);
or U37897 (N_37897,N_37573,N_37732);
nor U37898 (N_37898,N_37738,N_37556);
or U37899 (N_37899,N_37639,N_37621);
nand U37900 (N_37900,N_37501,N_37588);
nand U37901 (N_37901,N_37537,N_37643);
nand U37902 (N_37902,N_37700,N_37544);
xnor U37903 (N_37903,N_37666,N_37605);
nand U37904 (N_37904,N_37638,N_37582);
and U37905 (N_37905,N_37531,N_37721);
or U37906 (N_37906,N_37616,N_37506);
or U37907 (N_37907,N_37721,N_37544);
nand U37908 (N_37908,N_37571,N_37572);
or U37909 (N_37909,N_37655,N_37500);
nand U37910 (N_37910,N_37549,N_37523);
nand U37911 (N_37911,N_37506,N_37628);
nor U37912 (N_37912,N_37564,N_37572);
or U37913 (N_37913,N_37633,N_37728);
nand U37914 (N_37914,N_37569,N_37613);
or U37915 (N_37915,N_37568,N_37687);
nand U37916 (N_37916,N_37607,N_37522);
xnor U37917 (N_37917,N_37708,N_37671);
and U37918 (N_37918,N_37527,N_37576);
xor U37919 (N_37919,N_37743,N_37624);
xnor U37920 (N_37920,N_37509,N_37608);
or U37921 (N_37921,N_37697,N_37699);
nand U37922 (N_37922,N_37748,N_37594);
or U37923 (N_37923,N_37685,N_37679);
or U37924 (N_37924,N_37524,N_37749);
xor U37925 (N_37925,N_37520,N_37664);
nand U37926 (N_37926,N_37722,N_37614);
nor U37927 (N_37927,N_37696,N_37642);
nor U37928 (N_37928,N_37556,N_37528);
and U37929 (N_37929,N_37640,N_37727);
nor U37930 (N_37930,N_37717,N_37725);
and U37931 (N_37931,N_37539,N_37686);
nand U37932 (N_37932,N_37529,N_37724);
or U37933 (N_37933,N_37635,N_37583);
xor U37934 (N_37934,N_37697,N_37509);
xnor U37935 (N_37935,N_37532,N_37748);
nand U37936 (N_37936,N_37698,N_37617);
xnor U37937 (N_37937,N_37604,N_37689);
nand U37938 (N_37938,N_37643,N_37738);
or U37939 (N_37939,N_37667,N_37644);
nand U37940 (N_37940,N_37660,N_37657);
xor U37941 (N_37941,N_37523,N_37615);
and U37942 (N_37942,N_37714,N_37575);
and U37943 (N_37943,N_37688,N_37518);
and U37944 (N_37944,N_37584,N_37651);
xnor U37945 (N_37945,N_37655,N_37539);
nor U37946 (N_37946,N_37637,N_37711);
and U37947 (N_37947,N_37664,N_37656);
nor U37948 (N_37948,N_37627,N_37535);
nor U37949 (N_37949,N_37549,N_37593);
xnor U37950 (N_37950,N_37566,N_37521);
xor U37951 (N_37951,N_37519,N_37698);
nand U37952 (N_37952,N_37604,N_37566);
and U37953 (N_37953,N_37724,N_37566);
and U37954 (N_37954,N_37638,N_37537);
or U37955 (N_37955,N_37553,N_37644);
or U37956 (N_37956,N_37644,N_37560);
nand U37957 (N_37957,N_37713,N_37501);
or U37958 (N_37958,N_37532,N_37702);
nor U37959 (N_37959,N_37596,N_37677);
nand U37960 (N_37960,N_37541,N_37500);
nor U37961 (N_37961,N_37542,N_37612);
nor U37962 (N_37962,N_37729,N_37732);
and U37963 (N_37963,N_37636,N_37716);
nand U37964 (N_37964,N_37617,N_37610);
xor U37965 (N_37965,N_37632,N_37737);
nor U37966 (N_37966,N_37541,N_37723);
or U37967 (N_37967,N_37523,N_37501);
or U37968 (N_37968,N_37617,N_37518);
and U37969 (N_37969,N_37658,N_37509);
xor U37970 (N_37970,N_37632,N_37671);
and U37971 (N_37971,N_37518,N_37706);
and U37972 (N_37972,N_37526,N_37742);
xnor U37973 (N_37973,N_37734,N_37657);
or U37974 (N_37974,N_37672,N_37619);
nor U37975 (N_37975,N_37597,N_37577);
or U37976 (N_37976,N_37590,N_37530);
xor U37977 (N_37977,N_37590,N_37611);
or U37978 (N_37978,N_37659,N_37628);
nor U37979 (N_37979,N_37569,N_37527);
or U37980 (N_37980,N_37614,N_37685);
or U37981 (N_37981,N_37747,N_37726);
nor U37982 (N_37982,N_37504,N_37644);
and U37983 (N_37983,N_37724,N_37504);
and U37984 (N_37984,N_37550,N_37743);
and U37985 (N_37985,N_37633,N_37687);
and U37986 (N_37986,N_37569,N_37608);
or U37987 (N_37987,N_37739,N_37647);
xnor U37988 (N_37988,N_37553,N_37552);
or U37989 (N_37989,N_37568,N_37714);
xnor U37990 (N_37990,N_37631,N_37525);
nand U37991 (N_37991,N_37560,N_37655);
nand U37992 (N_37992,N_37505,N_37651);
and U37993 (N_37993,N_37588,N_37503);
nor U37994 (N_37994,N_37741,N_37736);
xnor U37995 (N_37995,N_37561,N_37539);
nand U37996 (N_37996,N_37648,N_37665);
nand U37997 (N_37997,N_37581,N_37662);
xor U37998 (N_37998,N_37604,N_37590);
nor U37999 (N_37999,N_37593,N_37624);
and U38000 (N_38000,N_37961,N_37778);
xor U38001 (N_38001,N_37821,N_37762);
nor U38002 (N_38002,N_37872,N_37839);
and U38003 (N_38003,N_37811,N_37789);
and U38004 (N_38004,N_37858,N_37819);
nand U38005 (N_38005,N_37825,N_37935);
and U38006 (N_38006,N_37909,N_37879);
xnor U38007 (N_38007,N_37865,N_37930);
or U38008 (N_38008,N_37950,N_37781);
or U38009 (N_38009,N_37992,N_37797);
nand U38010 (N_38010,N_37916,N_37970);
or U38011 (N_38011,N_37750,N_37860);
nor U38012 (N_38012,N_37818,N_37991);
and U38013 (N_38013,N_37886,N_37849);
or U38014 (N_38014,N_37840,N_37875);
or U38015 (N_38015,N_37948,N_37921);
or U38016 (N_38016,N_37812,N_37851);
and U38017 (N_38017,N_37842,N_37994);
or U38018 (N_38018,N_37843,N_37826);
and U38019 (N_38019,N_37969,N_37967);
and U38020 (N_38020,N_37862,N_37890);
and U38021 (N_38021,N_37814,N_37755);
xor U38022 (N_38022,N_37847,N_37771);
or U38023 (N_38023,N_37867,N_37897);
nand U38024 (N_38024,N_37864,N_37975);
xor U38025 (N_38025,N_37901,N_37866);
nor U38026 (N_38026,N_37989,N_37915);
xnor U38027 (N_38027,N_37968,N_37759);
nand U38028 (N_38028,N_37913,N_37808);
xor U38029 (N_38029,N_37936,N_37923);
or U38030 (N_38030,N_37955,N_37926);
or U38031 (N_38031,N_37845,N_37774);
nand U38032 (N_38032,N_37775,N_37827);
or U38033 (N_38033,N_37908,N_37919);
nand U38034 (N_38034,N_37883,N_37785);
nor U38035 (N_38035,N_37894,N_37939);
and U38036 (N_38036,N_37871,N_37979);
nor U38037 (N_38037,N_37941,N_37996);
and U38038 (N_38038,N_37780,N_37922);
nand U38039 (N_38039,N_37786,N_37873);
or U38040 (N_38040,N_37784,N_37777);
nand U38041 (N_38041,N_37960,N_37804);
xor U38042 (N_38042,N_37971,N_37795);
and U38043 (N_38043,N_37947,N_37856);
or U38044 (N_38044,N_37987,N_37768);
and U38045 (N_38045,N_37892,N_37918);
nand U38046 (N_38046,N_37816,N_37881);
or U38047 (N_38047,N_37751,N_37815);
and U38048 (N_38048,N_37752,N_37964);
nand U38049 (N_38049,N_37927,N_37942);
or U38050 (N_38050,N_37929,N_37857);
and U38051 (N_38051,N_37912,N_37834);
and U38052 (N_38052,N_37905,N_37809);
or U38053 (N_38053,N_37853,N_37829);
or U38054 (N_38054,N_37803,N_37760);
nand U38055 (N_38055,N_37754,N_37823);
nand U38056 (N_38056,N_37972,N_37928);
nor U38057 (N_38057,N_37914,N_37766);
and U38058 (N_38058,N_37830,N_37874);
xor U38059 (N_38059,N_37907,N_37962);
xor U38060 (N_38060,N_37999,N_37764);
nor U38061 (N_38061,N_37863,N_37954);
and U38062 (N_38062,N_37973,N_37765);
or U38063 (N_38063,N_37799,N_37917);
xnor U38064 (N_38064,N_37822,N_37798);
nor U38065 (N_38065,N_37938,N_37887);
nor U38066 (N_38066,N_37995,N_37833);
and U38067 (N_38067,N_37876,N_37753);
xnor U38068 (N_38068,N_37769,N_37956);
xnor U38069 (N_38069,N_37931,N_37761);
and U38070 (N_38070,N_37877,N_37899);
xnor U38071 (N_38071,N_37945,N_37924);
xnor U38072 (N_38072,N_37800,N_37966);
nand U38073 (N_38073,N_37852,N_37824);
nand U38074 (N_38074,N_37813,N_37934);
and U38075 (N_38075,N_37779,N_37984);
xor U38076 (N_38076,N_37997,N_37895);
and U38077 (N_38077,N_37859,N_37891);
nand U38078 (N_38078,N_37980,N_37990);
and U38079 (N_38079,N_37846,N_37952);
nand U38080 (N_38080,N_37787,N_37788);
xnor U38081 (N_38081,N_37898,N_37802);
and U38082 (N_38082,N_37817,N_37885);
xor U38083 (N_38083,N_37906,N_37981);
and U38084 (N_38084,N_37835,N_37937);
nor U38085 (N_38085,N_37807,N_37820);
nand U38086 (N_38086,N_37783,N_37793);
xor U38087 (N_38087,N_37953,N_37933);
or U38088 (N_38088,N_37903,N_37998);
nand U38089 (N_38089,N_37756,N_37869);
xor U38090 (N_38090,N_37828,N_37882);
xor U38091 (N_38091,N_37838,N_37889);
xor U38092 (N_38092,N_37986,N_37958);
nor U38093 (N_38093,N_37925,N_37884);
nor U38094 (N_38094,N_37893,N_37957);
and U38095 (N_38095,N_37932,N_37757);
and U38096 (N_38096,N_37910,N_37782);
or U38097 (N_38097,N_37848,N_37844);
xnor U38098 (N_38098,N_37792,N_37965);
or U38099 (N_38099,N_37772,N_37988);
nand U38100 (N_38100,N_37763,N_37837);
and U38101 (N_38101,N_37943,N_37861);
nand U38102 (N_38102,N_37770,N_37878);
nor U38103 (N_38103,N_37758,N_37790);
or U38104 (N_38104,N_37794,N_37911);
and U38105 (N_38105,N_37810,N_37902);
or U38106 (N_38106,N_37801,N_37946);
or U38107 (N_38107,N_37868,N_37767);
or U38108 (N_38108,N_37806,N_37896);
or U38109 (N_38109,N_37854,N_37949);
or U38110 (N_38110,N_37951,N_37855);
nor U38111 (N_38111,N_37776,N_37880);
or U38112 (N_38112,N_37982,N_37831);
and U38113 (N_38113,N_37805,N_37963);
nand U38114 (N_38114,N_37888,N_37850);
nor U38115 (N_38115,N_37836,N_37940);
or U38116 (N_38116,N_37904,N_37920);
or U38117 (N_38117,N_37900,N_37985);
nor U38118 (N_38118,N_37796,N_37976);
nand U38119 (N_38119,N_37978,N_37993);
xnor U38120 (N_38120,N_37959,N_37832);
nor U38121 (N_38121,N_37944,N_37791);
nand U38122 (N_38122,N_37983,N_37841);
xor U38123 (N_38123,N_37773,N_37977);
xnor U38124 (N_38124,N_37974,N_37870);
nand U38125 (N_38125,N_37847,N_37804);
and U38126 (N_38126,N_37984,N_37827);
nor U38127 (N_38127,N_37906,N_37773);
and U38128 (N_38128,N_37873,N_37764);
or U38129 (N_38129,N_37779,N_37999);
xnor U38130 (N_38130,N_37877,N_37819);
or U38131 (N_38131,N_37835,N_37790);
and U38132 (N_38132,N_37772,N_37909);
or U38133 (N_38133,N_37854,N_37994);
nand U38134 (N_38134,N_37844,N_37893);
nor U38135 (N_38135,N_37958,N_37834);
or U38136 (N_38136,N_37911,N_37822);
or U38137 (N_38137,N_37990,N_37823);
and U38138 (N_38138,N_37917,N_37957);
nand U38139 (N_38139,N_37985,N_37924);
nand U38140 (N_38140,N_37867,N_37817);
xor U38141 (N_38141,N_37928,N_37803);
xor U38142 (N_38142,N_37809,N_37997);
nor U38143 (N_38143,N_37895,N_37876);
nor U38144 (N_38144,N_37840,N_37862);
nand U38145 (N_38145,N_37797,N_37775);
nor U38146 (N_38146,N_37864,N_37964);
and U38147 (N_38147,N_37937,N_37871);
nor U38148 (N_38148,N_37810,N_37755);
xor U38149 (N_38149,N_37774,N_37853);
nor U38150 (N_38150,N_37853,N_37761);
xor U38151 (N_38151,N_37814,N_37757);
nor U38152 (N_38152,N_37834,N_37793);
or U38153 (N_38153,N_37854,N_37802);
or U38154 (N_38154,N_37767,N_37882);
xnor U38155 (N_38155,N_37919,N_37759);
and U38156 (N_38156,N_37945,N_37880);
nand U38157 (N_38157,N_37782,N_37849);
and U38158 (N_38158,N_37869,N_37778);
nor U38159 (N_38159,N_37915,N_37887);
and U38160 (N_38160,N_37817,N_37914);
or U38161 (N_38161,N_37994,N_37830);
and U38162 (N_38162,N_37856,N_37828);
and U38163 (N_38163,N_37805,N_37750);
xor U38164 (N_38164,N_37821,N_37939);
nor U38165 (N_38165,N_37965,N_37836);
and U38166 (N_38166,N_37953,N_37770);
nand U38167 (N_38167,N_37798,N_37815);
xor U38168 (N_38168,N_37833,N_37881);
or U38169 (N_38169,N_37939,N_37984);
xor U38170 (N_38170,N_37752,N_37877);
or U38171 (N_38171,N_37847,N_37782);
nor U38172 (N_38172,N_37791,N_37903);
nor U38173 (N_38173,N_37875,N_37856);
nand U38174 (N_38174,N_37952,N_37925);
nand U38175 (N_38175,N_37908,N_37891);
nor U38176 (N_38176,N_37776,N_37797);
nand U38177 (N_38177,N_37989,N_37836);
or U38178 (N_38178,N_37819,N_37907);
or U38179 (N_38179,N_37971,N_37949);
and U38180 (N_38180,N_37870,N_37758);
or U38181 (N_38181,N_37766,N_37882);
nand U38182 (N_38182,N_37750,N_37977);
or U38183 (N_38183,N_37902,N_37985);
nand U38184 (N_38184,N_37821,N_37851);
nand U38185 (N_38185,N_37883,N_37835);
xor U38186 (N_38186,N_37896,N_37776);
and U38187 (N_38187,N_37980,N_37925);
and U38188 (N_38188,N_37837,N_37808);
and U38189 (N_38189,N_37794,N_37775);
or U38190 (N_38190,N_37892,N_37755);
and U38191 (N_38191,N_37787,N_37823);
and U38192 (N_38192,N_37815,N_37789);
and U38193 (N_38193,N_37913,N_37767);
nand U38194 (N_38194,N_37824,N_37776);
and U38195 (N_38195,N_37883,N_37959);
or U38196 (N_38196,N_37811,N_37783);
nand U38197 (N_38197,N_37873,N_37947);
or U38198 (N_38198,N_37941,N_37793);
nor U38199 (N_38199,N_37943,N_37989);
nand U38200 (N_38200,N_37988,N_37974);
nor U38201 (N_38201,N_37907,N_37772);
nand U38202 (N_38202,N_37803,N_37756);
nand U38203 (N_38203,N_37907,N_37911);
xnor U38204 (N_38204,N_37832,N_37943);
and U38205 (N_38205,N_37892,N_37994);
and U38206 (N_38206,N_37898,N_37814);
nand U38207 (N_38207,N_37856,N_37866);
nand U38208 (N_38208,N_37947,N_37998);
and U38209 (N_38209,N_37835,N_37762);
xnor U38210 (N_38210,N_37944,N_37999);
nand U38211 (N_38211,N_37938,N_37768);
or U38212 (N_38212,N_37759,N_37980);
and U38213 (N_38213,N_37784,N_37977);
xor U38214 (N_38214,N_37978,N_37965);
nand U38215 (N_38215,N_37966,N_37802);
or U38216 (N_38216,N_37954,N_37756);
nand U38217 (N_38217,N_37765,N_37840);
nand U38218 (N_38218,N_37977,N_37971);
xor U38219 (N_38219,N_37837,N_37824);
or U38220 (N_38220,N_37841,N_37928);
nor U38221 (N_38221,N_37931,N_37866);
nor U38222 (N_38222,N_37783,N_37777);
xor U38223 (N_38223,N_37773,N_37873);
nand U38224 (N_38224,N_37780,N_37991);
nor U38225 (N_38225,N_37919,N_37822);
or U38226 (N_38226,N_37940,N_37855);
nand U38227 (N_38227,N_37925,N_37883);
nor U38228 (N_38228,N_37904,N_37905);
xor U38229 (N_38229,N_37792,N_37976);
or U38230 (N_38230,N_37751,N_37762);
xnor U38231 (N_38231,N_37899,N_37780);
nor U38232 (N_38232,N_37904,N_37832);
or U38233 (N_38233,N_37815,N_37944);
nor U38234 (N_38234,N_37900,N_37987);
xor U38235 (N_38235,N_37924,N_37765);
and U38236 (N_38236,N_37797,N_37853);
xor U38237 (N_38237,N_37753,N_37825);
and U38238 (N_38238,N_37979,N_37762);
xor U38239 (N_38239,N_37924,N_37782);
nor U38240 (N_38240,N_37825,N_37843);
or U38241 (N_38241,N_37773,N_37978);
nand U38242 (N_38242,N_37791,N_37860);
nand U38243 (N_38243,N_37944,N_37758);
and U38244 (N_38244,N_37976,N_37999);
nor U38245 (N_38245,N_37876,N_37862);
nand U38246 (N_38246,N_37834,N_37797);
and U38247 (N_38247,N_37807,N_37984);
nor U38248 (N_38248,N_37958,N_37869);
xnor U38249 (N_38249,N_37883,N_37794);
nand U38250 (N_38250,N_38180,N_38201);
xnor U38251 (N_38251,N_38135,N_38025);
and U38252 (N_38252,N_38038,N_38030);
nand U38253 (N_38253,N_38168,N_38238);
or U38254 (N_38254,N_38119,N_38214);
nand U38255 (N_38255,N_38106,N_38227);
nand U38256 (N_38256,N_38126,N_38163);
nor U38257 (N_38257,N_38023,N_38008);
nand U38258 (N_38258,N_38215,N_38095);
nor U38259 (N_38259,N_38047,N_38129);
nand U38260 (N_38260,N_38173,N_38149);
nand U38261 (N_38261,N_38084,N_38154);
or U38262 (N_38262,N_38088,N_38140);
xor U38263 (N_38263,N_38145,N_38178);
nor U38264 (N_38264,N_38010,N_38114);
and U38265 (N_38265,N_38086,N_38108);
and U38266 (N_38266,N_38220,N_38041);
nor U38267 (N_38267,N_38111,N_38228);
nor U38268 (N_38268,N_38059,N_38068);
or U38269 (N_38269,N_38222,N_38132);
and U38270 (N_38270,N_38170,N_38175);
nor U38271 (N_38271,N_38062,N_38174);
nand U38272 (N_38272,N_38065,N_38031);
nand U38273 (N_38273,N_38165,N_38057);
nor U38274 (N_38274,N_38157,N_38167);
nand U38275 (N_38275,N_38051,N_38247);
nor U38276 (N_38276,N_38039,N_38120);
xnor U38277 (N_38277,N_38211,N_38133);
xor U38278 (N_38278,N_38054,N_38033);
xnor U38279 (N_38279,N_38061,N_38105);
nand U38280 (N_38280,N_38182,N_38002);
and U38281 (N_38281,N_38009,N_38052);
xor U38282 (N_38282,N_38164,N_38118);
and U38283 (N_38283,N_38124,N_38171);
or U38284 (N_38284,N_38102,N_38172);
and U38285 (N_38285,N_38055,N_38050);
and U38286 (N_38286,N_38148,N_38067);
xnor U38287 (N_38287,N_38212,N_38240);
nand U38288 (N_38288,N_38185,N_38001);
xor U38289 (N_38289,N_38027,N_38045);
and U38290 (N_38290,N_38071,N_38166);
xnor U38291 (N_38291,N_38152,N_38037);
xnor U38292 (N_38292,N_38053,N_38121);
or U38293 (N_38293,N_38090,N_38199);
xnor U38294 (N_38294,N_38198,N_38181);
nand U38295 (N_38295,N_38122,N_38007);
nand U38296 (N_38296,N_38083,N_38018);
or U38297 (N_38297,N_38242,N_38116);
xor U38298 (N_38298,N_38161,N_38158);
nor U38299 (N_38299,N_38094,N_38239);
or U38300 (N_38300,N_38013,N_38097);
or U38301 (N_38301,N_38249,N_38003);
nand U38302 (N_38302,N_38006,N_38017);
or U38303 (N_38303,N_38169,N_38110);
nand U38304 (N_38304,N_38075,N_38064);
nor U38305 (N_38305,N_38237,N_38021);
xor U38306 (N_38306,N_38024,N_38049);
nand U38307 (N_38307,N_38096,N_38142);
nand U38308 (N_38308,N_38179,N_38139);
xor U38309 (N_38309,N_38034,N_38011);
nor U38310 (N_38310,N_38012,N_38123);
and U38311 (N_38311,N_38066,N_38107);
nand U38312 (N_38312,N_38223,N_38153);
and U38313 (N_38313,N_38141,N_38207);
nor U38314 (N_38314,N_38208,N_38104);
nor U38315 (N_38315,N_38092,N_38243);
or U38316 (N_38316,N_38127,N_38109);
xnor U38317 (N_38317,N_38248,N_38087);
xnor U38318 (N_38318,N_38245,N_38091);
nor U38319 (N_38319,N_38156,N_38078);
nand U38320 (N_38320,N_38103,N_38230);
nand U38321 (N_38321,N_38194,N_38098);
nor U38322 (N_38322,N_38079,N_38246);
xnor U38323 (N_38323,N_38115,N_38204);
xor U38324 (N_38324,N_38085,N_38082);
xnor U38325 (N_38325,N_38004,N_38183);
nand U38326 (N_38326,N_38042,N_38036);
or U38327 (N_38327,N_38138,N_38216);
nand U38328 (N_38328,N_38048,N_38128);
xor U38329 (N_38329,N_38044,N_38219);
and U38330 (N_38330,N_38229,N_38077);
and U38331 (N_38331,N_38160,N_38159);
nor U38332 (N_38332,N_38100,N_38040);
or U38333 (N_38333,N_38224,N_38162);
nor U38334 (N_38334,N_38187,N_38234);
xnor U38335 (N_38335,N_38236,N_38069);
or U38336 (N_38336,N_38020,N_38137);
nand U38337 (N_38337,N_38093,N_38203);
nor U38338 (N_38338,N_38029,N_38113);
nor U38339 (N_38339,N_38131,N_38101);
or U38340 (N_38340,N_38231,N_38213);
or U38341 (N_38341,N_38080,N_38150);
and U38342 (N_38342,N_38112,N_38184);
and U38343 (N_38343,N_38176,N_38015);
or U38344 (N_38344,N_38043,N_38233);
xor U38345 (N_38345,N_38019,N_38209);
or U38346 (N_38346,N_38076,N_38028);
and U38347 (N_38347,N_38151,N_38221);
xnor U38348 (N_38348,N_38130,N_38196);
xnor U38349 (N_38349,N_38155,N_38144);
nand U38350 (N_38350,N_38060,N_38205);
or U38351 (N_38351,N_38026,N_38063);
nand U38352 (N_38352,N_38195,N_38058);
or U38353 (N_38353,N_38192,N_38190);
or U38354 (N_38354,N_38188,N_38210);
nand U38355 (N_38355,N_38022,N_38032);
or U38356 (N_38356,N_38218,N_38125);
xnor U38357 (N_38357,N_38191,N_38226);
nor U38358 (N_38358,N_38016,N_38073);
nand U38359 (N_38359,N_38056,N_38147);
and U38360 (N_38360,N_38134,N_38005);
nor U38361 (N_38361,N_38225,N_38177);
nand U38362 (N_38362,N_38081,N_38197);
nand U38363 (N_38363,N_38193,N_38202);
and U38364 (N_38364,N_38244,N_38143);
nand U38365 (N_38365,N_38186,N_38072);
and U38366 (N_38366,N_38206,N_38136);
nand U38367 (N_38367,N_38099,N_38200);
xor U38368 (N_38368,N_38014,N_38089);
nand U38369 (N_38369,N_38046,N_38117);
and U38370 (N_38370,N_38189,N_38035);
xnor U38371 (N_38371,N_38232,N_38235);
nor U38372 (N_38372,N_38217,N_38070);
or U38373 (N_38373,N_38241,N_38146);
nand U38374 (N_38374,N_38074,N_38000);
or U38375 (N_38375,N_38209,N_38208);
nand U38376 (N_38376,N_38034,N_38138);
nor U38377 (N_38377,N_38060,N_38227);
nand U38378 (N_38378,N_38144,N_38170);
xnor U38379 (N_38379,N_38052,N_38182);
and U38380 (N_38380,N_38222,N_38147);
nor U38381 (N_38381,N_38209,N_38197);
or U38382 (N_38382,N_38231,N_38024);
nor U38383 (N_38383,N_38008,N_38016);
nand U38384 (N_38384,N_38082,N_38132);
and U38385 (N_38385,N_38139,N_38147);
xnor U38386 (N_38386,N_38173,N_38012);
xnor U38387 (N_38387,N_38090,N_38099);
and U38388 (N_38388,N_38171,N_38209);
xnor U38389 (N_38389,N_38039,N_38227);
or U38390 (N_38390,N_38159,N_38134);
nand U38391 (N_38391,N_38038,N_38231);
or U38392 (N_38392,N_38114,N_38116);
nand U38393 (N_38393,N_38220,N_38238);
nand U38394 (N_38394,N_38120,N_38112);
nand U38395 (N_38395,N_38061,N_38121);
and U38396 (N_38396,N_38109,N_38101);
nor U38397 (N_38397,N_38185,N_38111);
or U38398 (N_38398,N_38162,N_38148);
xor U38399 (N_38399,N_38114,N_38183);
or U38400 (N_38400,N_38170,N_38222);
nor U38401 (N_38401,N_38008,N_38159);
and U38402 (N_38402,N_38058,N_38002);
nand U38403 (N_38403,N_38043,N_38175);
or U38404 (N_38404,N_38037,N_38119);
nor U38405 (N_38405,N_38112,N_38077);
or U38406 (N_38406,N_38041,N_38053);
and U38407 (N_38407,N_38059,N_38000);
and U38408 (N_38408,N_38189,N_38129);
nor U38409 (N_38409,N_38050,N_38166);
nand U38410 (N_38410,N_38082,N_38078);
nor U38411 (N_38411,N_38198,N_38230);
nand U38412 (N_38412,N_38155,N_38013);
nand U38413 (N_38413,N_38122,N_38224);
xor U38414 (N_38414,N_38249,N_38063);
or U38415 (N_38415,N_38036,N_38025);
nor U38416 (N_38416,N_38066,N_38247);
and U38417 (N_38417,N_38063,N_38111);
nand U38418 (N_38418,N_38114,N_38038);
nor U38419 (N_38419,N_38121,N_38023);
nor U38420 (N_38420,N_38128,N_38075);
nor U38421 (N_38421,N_38200,N_38188);
nor U38422 (N_38422,N_38146,N_38155);
nor U38423 (N_38423,N_38138,N_38002);
and U38424 (N_38424,N_38238,N_38040);
or U38425 (N_38425,N_38130,N_38199);
nand U38426 (N_38426,N_38024,N_38017);
and U38427 (N_38427,N_38027,N_38059);
nor U38428 (N_38428,N_38039,N_38007);
xnor U38429 (N_38429,N_38021,N_38150);
and U38430 (N_38430,N_38182,N_38054);
or U38431 (N_38431,N_38197,N_38242);
or U38432 (N_38432,N_38219,N_38218);
nor U38433 (N_38433,N_38074,N_38220);
nor U38434 (N_38434,N_38148,N_38005);
and U38435 (N_38435,N_38008,N_38029);
nor U38436 (N_38436,N_38011,N_38232);
and U38437 (N_38437,N_38052,N_38096);
or U38438 (N_38438,N_38068,N_38125);
xor U38439 (N_38439,N_38029,N_38035);
nand U38440 (N_38440,N_38248,N_38072);
or U38441 (N_38441,N_38139,N_38115);
xnor U38442 (N_38442,N_38116,N_38245);
xor U38443 (N_38443,N_38071,N_38171);
xor U38444 (N_38444,N_38175,N_38229);
or U38445 (N_38445,N_38013,N_38211);
xnor U38446 (N_38446,N_38146,N_38035);
nor U38447 (N_38447,N_38145,N_38046);
and U38448 (N_38448,N_38239,N_38009);
or U38449 (N_38449,N_38068,N_38212);
or U38450 (N_38450,N_38124,N_38170);
xor U38451 (N_38451,N_38225,N_38135);
or U38452 (N_38452,N_38221,N_38038);
nand U38453 (N_38453,N_38112,N_38001);
nor U38454 (N_38454,N_38039,N_38080);
and U38455 (N_38455,N_38087,N_38158);
nor U38456 (N_38456,N_38075,N_38193);
nor U38457 (N_38457,N_38207,N_38197);
nand U38458 (N_38458,N_38028,N_38080);
xor U38459 (N_38459,N_38126,N_38145);
and U38460 (N_38460,N_38229,N_38118);
nor U38461 (N_38461,N_38046,N_38072);
or U38462 (N_38462,N_38034,N_38064);
xor U38463 (N_38463,N_38135,N_38204);
nand U38464 (N_38464,N_38236,N_38171);
nand U38465 (N_38465,N_38187,N_38201);
and U38466 (N_38466,N_38074,N_38008);
nand U38467 (N_38467,N_38058,N_38190);
nand U38468 (N_38468,N_38006,N_38196);
and U38469 (N_38469,N_38098,N_38248);
nor U38470 (N_38470,N_38247,N_38016);
nor U38471 (N_38471,N_38011,N_38248);
nand U38472 (N_38472,N_38081,N_38223);
or U38473 (N_38473,N_38203,N_38248);
and U38474 (N_38474,N_38022,N_38102);
nand U38475 (N_38475,N_38133,N_38224);
xor U38476 (N_38476,N_38089,N_38204);
nor U38477 (N_38477,N_38090,N_38151);
and U38478 (N_38478,N_38108,N_38137);
nand U38479 (N_38479,N_38175,N_38124);
xnor U38480 (N_38480,N_38111,N_38219);
nand U38481 (N_38481,N_38104,N_38021);
or U38482 (N_38482,N_38062,N_38116);
nor U38483 (N_38483,N_38150,N_38087);
or U38484 (N_38484,N_38155,N_38185);
or U38485 (N_38485,N_38008,N_38001);
or U38486 (N_38486,N_38037,N_38012);
xor U38487 (N_38487,N_38099,N_38183);
nand U38488 (N_38488,N_38181,N_38050);
nor U38489 (N_38489,N_38073,N_38082);
nand U38490 (N_38490,N_38053,N_38057);
and U38491 (N_38491,N_38040,N_38133);
nor U38492 (N_38492,N_38232,N_38031);
xor U38493 (N_38493,N_38063,N_38017);
xor U38494 (N_38494,N_38157,N_38120);
nor U38495 (N_38495,N_38166,N_38082);
xor U38496 (N_38496,N_38110,N_38123);
or U38497 (N_38497,N_38204,N_38113);
nand U38498 (N_38498,N_38075,N_38160);
xnor U38499 (N_38499,N_38026,N_38155);
nor U38500 (N_38500,N_38426,N_38444);
xor U38501 (N_38501,N_38445,N_38411);
nand U38502 (N_38502,N_38391,N_38295);
nand U38503 (N_38503,N_38493,N_38376);
nor U38504 (N_38504,N_38433,N_38382);
nand U38505 (N_38505,N_38451,N_38386);
xnor U38506 (N_38506,N_38319,N_38264);
or U38507 (N_38507,N_38372,N_38306);
nor U38508 (N_38508,N_38487,N_38374);
nand U38509 (N_38509,N_38480,N_38318);
and U38510 (N_38510,N_38257,N_38277);
or U38511 (N_38511,N_38349,N_38390);
or U38512 (N_38512,N_38404,N_38330);
xor U38513 (N_38513,N_38356,N_38428);
or U38514 (N_38514,N_38381,N_38465);
xnor U38515 (N_38515,N_38308,N_38347);
and U38516 (N_38516,N_38410,N_38271);
and U38517 (N_38517,N_38394,N_38345);
nor U38518 (N_38518,N_38405,N_38299);
nand U38519 (N_38519,N_38393,N_38291);
or U38520 (N_38520,N_38418,N_38352);
or U38521 (N_38521,N_38425,N_38348);
or U38522 (N_38522,N_38430,N_38340);
and U38523 (N_38523,N_38378,N_38303);
nand U38524 (N_38524,N_38252,N_38407);
xor U38525 (N_38525,N_38469,N_38471);
or U38526 (N_38526,N_38259,N_38324);
nand U38527 (N_38527,N_38311,N_38290);
and U38528 (N_38528,N_38305,N_38287);
xor U38529 (N_38529,N_38454,N_38423);
and U38530 (N_38530,N_38379,N_38281);
or U38531 (N_38531,N_38440,N_38265);
nand U38532 (N_38532,N_38457,N_38355);
and U38533 (N_38533,N_38398,N_38453);
nor U38534 (N_38534,N_38496,N_38293);
nand U38535 (N_38535,N_38263,N_38338);
nor U38536 (N_38536,N_38343,N_38432);
nor U38537 (N_38537,N_38392,N_38399);
and U38538 (N_38538,N_38498,N_38365);
nand U38539 (N_38539,N_38371,N_38409);
nand U38540 (N_38540,N_38422,N_38307);
or U38541 (N_38541,N_38304,N_38342);
and U38542 (N_38542,N_38479,N_38364);
xor U38543 (N_38543,N_38312,N_38437);
nand U38544 (N_38544,N_38276,N_38475);
xnor U38545 (N_38545,N_38359,N_38270);
and U38546 (N_38546,N_38412,N_38462);
nand U38547 (N_38547,N_38461,N_38325);
or U38548 (N_38548,N_38280,N_38383);
nor U38549 (N_38549,N_38458,N_38310);
nor U38550 (N_38550,N_38344,N_38492);
or U38551 (N_38551,N_38297,N_38488);
or U38552 (N_38552,N_38401,N_38414);
xnor U38553 (N_38553,N_38357,N_38363);
or U38554 (N_38554,N_38258,N_38354);
nand U38555 (N_38555,N_38387,N_38251);
xor U38556 (N_38556,N_38341,N_38370);
and U38557 (N_38557,N_38402,N_38420);
or U38558 (N_38558,N_38294,N_38368);
nor U38559 (N_38559,N_38255,N_38460);
nor U38560 (N_38560,N_38415,N_38283);
nand U38561 (N_38561,N_38384,N_38400);
or U38562 (N_38562,N_38267,N_38464);
or U38563 (N_38563,N_38482,N_38334);
and U38564 (N_38564,N_38327,N_38473);
and U38565 (N_38565,N_38266,N_38360);
nor U38566 (N_38566,N_38362,N_38250);
or U38567 (N_38567,N_38323,N_38431);
nor U38568 (N_38568,N_38481,N_38439);
and U38569 (N_38569,N_38260,N_38302);
xnor U38570 (N_38570,N_38388,N_38494);
and U38571 (N_38571,N_38315,N_38463);
and U38572 (N_38572,N_38467,N_38489);
nand U38573 (N_38573,N_38328,N_38477);
nand U38574 (N_38574,N_38397,N_38375);
and U38575 (N_38575,N_38320,N_38421);
and U38576 (N_38576,N_38274,N_38403);
nor U38577 (N_38577,N_38455,N_38335);
nor U38578 (N_38578,N_38326,N_38373);
and U38579 (N_38579,N_38329,N_38485);
xor U38580 (N_38580,N_38497,N_38256);
nand U38581 (N_38581,N_38450,N_38486);
nor U38582 (N_38582,N_38316,N_38272);
nand U38583 (N_38583,N_38275,N_38322);
and U38584 (N_38584,N_38446,N_38495);
nor U38585 (N_38585,N_38476,N_38361);
xor U38586 (N_38586,N_38254,N_38483);
and U38587 (N_38587,N_38491,N_38478);
nand U38588 (N_38588,N_38351,N_38292);
nor U38589 (N_38589,N_38434,N_38273);
nand U38590 (N_38590,N_38380,N_38435);
xnor U38591 (N_38591,N_38484,N_38331);
xor U38592 (N_38592,N_38296,N_38253);
xnor U38593 (N_38593,N_38332,N_38313);
or U38594 (N_38594,N_38456,N_38416);
nor U38595 (N_38595,N_38366,N_38474);
nand U38596 (N_38596,N_38395,N_38468);
or U38597 (N_38597,N_38408,N_38289);
nor U38598 (N_38598,N_38470,N_38429);
or U38599 (N_38599,N_38309,N_38314);
and U38600 (N_38600,N_38499,N_38406);
nor U38601 (N_38601,N_38419,N_38377);
and U38602 (N_38602,N_38353,N_38427);
or U38603 (N_38603,N_38438,N_38336);
xnor U38604 (N_38604,N_38449,N_38300);
xnor U38605 (N_38605,N_38369,N_38396);
or U38606 (N_38606,N_38358,N_38284);
and U38607 (N_38607,N_38333,N_38459);
nor U38608 (N_38608,N_38301,N_38443);
or U38609 (N_38609,N_38472,N_38413);
nand U38610 (N_38610,N_38288,N_38262);
nor U38611 (N_38611,N_38448,N_38279);
or U38612 (N_38612,N_38317,N_38346);
xor U38613 (N_38613,N_38268,N_38466);
nand U38614 (N_38614,N_38282,N_38367);
nand U38615 (N_38615,N_38339,N_38337);
nor U38616 (N_38616,N_38442,N_38285);
nand U38617 (N_38617,N_38441,N_38261);
or U38618 (N_38618,N_38385,N_38278);
xnor U38619 (N_38619,N_38452,N_38436);
xor U38620 (N_38620,N_38286,N_38269);
nand U38621 (N_38621,N_38350,N_38321);
or U38622 (N_38622,N_38298,N_38490);
nand U38623 (N_38623,N_38447,N_38417);
or U38624 (N_38624,N_38389,N_38424);
nand U38625 (N_38625,N_38330,N_38351);
xnor U38626 (N_38626,N_38495,N_38276);
nor U38627 (N_38627,N_38332,N_38489);
and U38628 (N_38628,N_38306,N_38388);
or U38629 (N_38629,N_38357,N_38369);
or U38630 (N_38630,N_38499,N_38305);
xor U38631 (N_38631,N_38401,N_38317);
nor U38632 (N_38632,N_38250,N_38402);
nand U38633 (N_38633,N_38274,N_38278);
and U38634 (N_38634,N_38414,N_38381);
nor U38635 (N_38635,N_38492,N_38376);
xnor U38636 (N_38636,N_38461,N_38280);
or U38637 (N_38637,N_38423,N_38384);
or U38638 (N_38638,N_38462,N_38273);
nor U38639 (N_38639,N_38258,N_38415);
xor U38640 (N_38640,N_38261,N_38326);
nor U38641 (N_38641,N_38256,N_38456);
nand U38642 (N_38642,N_38288,N_38411);
and U38643 (N_38643,N_38420,N_38446);
xor U38644 (N_38644,N_38496,N_38485);
nor U38645 (N_38645,N_38279,N_38420);
or U38646 (N_38646,N_38305,N_38298);
nand U38647 (N_38647,N_38435,N_38283);
or U38648 (N_38648,N_38455,N_38331);
nor U38649 (N_38649,N_38323,N_38460);
nand U38650 (N_38650,N_38420,N_38479);
xnor U38651 (N_38651,N_38429,N_38250);
or U38652 (N_38652,N_38260,N_38379);
xnor U38653 (N_38653,N_38499,N_38324);
xnor U38654 (N_38654,N_38283,N_38270);
and U38655 (N_38655,N_38442,N_38454);
nor U38656 (N_38656,N_38413,N_38336);
nor U38657 (N_38657,N_38303,N_38263);
nor U38658 (N_38658,N_38306,N_38450);
or U38659 (N_38659,N_38438,N_38375);
nand U38660 (N_38660,N_38456,N_38294);
and U38661 (N_38661,N_38340,N_38289);
or U38662 (N_38662,N_38351,N_38461);
or U38663 (N_38663,N_38421,N_38404);
or U38664 (N_38664,N_38282,N_38285);
nand U38665 (N_38665,N_38279,N_38289);
xor U38666 (N_38666,N_38485,N_38479);
and U38667 (N_38667,N_38274,N_38430);
xor U38668 (N_38668,N_38434,N_38265);
nand U38669 (N_38669,N_38315,N_38485);
xnor U38670 (N_38670,N_38322,N_38498);
nor U38671 (N_38671,N_38436,N_38272);
or U38672 (N_38672,N_38252,N_38342);
and U38673 (N_38673,N_38344,N_38324);
and U38674 (N_38674,N_38413,N_38384);
or U38675 (N_38675,N_38417,N_38271);
nor U38676 (N_38676,N_38357,N_38383);
or U38677 (N_38677,N_38269,N_38367);
nand U38678 (N_38678,N_38447,N_38267);
nor U38679 (N_38679,N_38393,N_38461);
xnor U38680 (N_38680,N_38446,N_38342);
nand U38681 (N_38681,N_38258,N_38478);
xor U38682 (N_38682,N_38415,N_38334);
nand U38683 (N_38683,N_38322,N_38437);
nand U38684 (N_38684,N_38378,N_38270);
and U38685 (N_38685,N_38486,N_38341);
and U38686 (N_38686,N_38252,N_38280);
xnor U38687 (N_38687,N_38448,N_38443);
nand U38688 (N_38688,N_38310,N_38398);
nand U38689 (N_38689,N_38392,N_38293);
nor U38690 (N_38690,N_38440,N_38395);
xor U38691 (N_38691,N_38370,N_38429);
and U38692 (N_38692,N_38346,N_38459);
or U38693 (N_38693,N_38399,N_38259);
nand U38694 (N_38694,N_38402,N_38317);
nand U38695 (N_38695,N_38319,N_38350);
or U38696 (N_38696,N_38324,N_38270);
xor U38697 (N_38697,N_38436,N_38492);
xnor U38698 (N_38698,N_38385,N_38376);
or U38699 (N_38699,N_38358,N_38327);
xor U38700 (N_38700,N_38497,N_38412);
and U38701 (N_38701,N_38360,N_38415);
xnor U38702 (N_38702,N_38443,N_38262);
or U38703 (N_38703,N_38349,N_38363);
xor U38704 (N_38704,N_38414,N_38293);
nor U38705 (N_38705,N_38356,N_38301);
nand U38706 (N_38706,N_38258,N_38261);
and U38707 (N_38707,N_38330,N_38467);
or U38708 (N_38708,N_38399,N_38378);
nor U38709 (N_38709,N_38337,N_38472);
nor U38710 (N_38710,N_38481,N_38277);
xnor U38711 (N_38711,N_38305,N_38423);
nand U38712 (N_38712,N_38278,N_38416);
and U38713 (N_38713,N_38343,N_38459);
nor U38714 (N_38714,N_38383,N_38296);
or U38715 (N_38715,N_38488,N_38374);
and U38716 (N_38716,N_38310,N_38288);
or U38717 (N_38717,N_38282,N_38422);
nand U38718 (N_38718,N_38328,N_38465);
or U38719 (N_38719,N_38311,N_38482);
nand U38720 (N_38720,N_38445,N_38308);
xnor U38721 (N_38721,N_38274,N_38379);
nor U38722 (N_38722,N_38313,N_38436);
or U38723 (N_38723,N_38397,N_38417);
or U38724 (N_38724,N_38398,N_38417);
xor U38725 (N_38725,N_38470,N_38283);
nor U38726 (N_38726,N_38406,N_38285);
nor U38727 (N_38727,N_38447,N_38420);
or U38728 (N_38728,N_38327,N_38436);
xnor U38729 (N_38729,N_38455,N_38423);
nand U38730 (N_38730,N_38337,N_38353);
and U38731 (N_38731,N_38417,N_38285);
or U38732 (N_38732,N_38305,N_38292);
nor U38733 (N_38733,N_38274,N_38344);
nor U38734 (N_38734,N_38483,N_38407);
or U38735 (N_38735,N_38287,N_38259);
or U38736 (N_38736,N_38466,N_38497);
or U38737 (N_38737,N_38430,N_38306);
nor U38738 (N_38738,N_38463,N_38313);
xnor U38739 (N_38739,N_38386,N_38499);
nand U38740 (N_38740,N_38291,N_38259);
nand U38741 (N_38741,N_38447,N_38373);
xnor U38742 (N_38742,N_38349,N_38428);
xor U38743 (N_38743,N_38430,N_38390);
nand U38744 (N_38744,N_38343,N_38455);
or U38745 (N_38745,N_38423,N_38312);
and U38746 (N_38746,N_38404,N_38331);
nor U38747 (N_38747,N_38384,N_38498);
nor U38748 (N_38748,N_38476,N_38371);
xnor U38749 (N_38749,N_38371,N_38282);
or U38750 (N_38750,N_38657,N_38654);
or U38751 (N_38751,N_38627,N_38676);
xor U38752 (N_38752,N_38622,N_38641);
nand U38753 (N_38753,N_38561,N_38644);
nor U38754 (N_38754,N_38541,N_38574);
nand U38755 (N_38755,N_38702,N_38546);
or U38756 (N_38756,N_38637,N_38557);
nor U38757 (N_38757,N_38513,N_38519);
nand U38758 (N_38758,N_38636,N_38577);
nand U38759 (N_38759,N_38529,N_38616);
and U38760 (N_38760,N_38647,N_38549);
and U38761 (N_38761,N_38500,N_38727);
nand U38762 (N_38762,N_38722,N_38655);
xor U38763 (N_38763,N_38720,N_38586);
or U38764 (N_38764,N_38712,N_38645);
nor U38765 (N_38765,N_38539,N_38594);
xnor U38766 (N_38766,N_38692,N_38560);
xnor U38767 (N_38767,N_38666,N_38584);
nor U38768 (N_38768,N_38661,N_38569);
or U38769 (N_38769,N_38599,N_38682);
xor U38770 (N_38770,N_38679,N_38533);
or U38771 (N_38771,N_38619,N_38538);
and U38772 (N_38772,N_38648,N_38521);
nor U38773 (N_38773,N_38638,N_38597);
and U38774 (N_38774,N_38534,N_38578);
nand U38775 (N_38775,N_38608,N_38553);
or U38776 (N_38776,N_38680,N_38516);
nor U38777 (N_38777,N_38536,N_38741);
nor U38778 (N_38778,N_38512,N_38522);
and U38779 (N_38779,N_38517,N_38677);
xor U38780 (N_38780,N_38663,N_38691);
nand U38781 (N_38781,N_38545,N_38664);
nand U38782 (N_38782,N_38709,N_38523);
xnor U38783 (N_38783,N_38734,N_38703);
and U38784 (N_38784,N_38711,N_38504);
nor U38785 (N_38785,N_38724,N_38650);
or U38786 (N_38786,N_38547,N_38592);
nor U38787 (N_38787,N_38696,N_38564);
and U38788 (N_38788,N_38740,N_38742);
nand U38789 (N_38789,N_38640,N_38572);
or U38790 (N_38790,N_38503,N_38735);
nor U38791 (N_38791,N_38704,N_38725);
nand U38792 (N_38792,N_38581,N_38714);
nand U38793 (N_38793,N_38531,N_38507);
and U38794 (N_38794,N_38672,N_38675);
xnor U38795 (N_38795,N_38548,N_38625);
nor U38796 (N_38796,N_38745,N_38566);
and U38797 (N_38797,N_38543,N_38552);
xnor U38798 (N_38798,N_38623,N_38733);
nand U38799 (N_38799,N_38726,N_38731);
nand U38800 (N_38800,N_38620,N_38532);
or U38801 (N_38801,N_38631,N_38652);
nor U38802 (N_38802,N_38690,N_38550);
nor U38803 (N_38803,N_38715,N_38705);
nand U38804 (N_38804,N_38514,N_38662);
nor U38805 (N_38805,N_38748,N_38670);
and U38806 (N_38806,N_38593,N_38567);
nand U38807 (N_38807,N_38525,N_38573);
or U38808 (N_38808,N_38602,N_38686);
or U38809 (N_38809,N_38687,N_38565);
and U38810 (N_38810,N_38669,N_38646);
xor U38811 (N_38811,N_38626,N_38629);
or U38812 (N_38812,N_38511,N_38613);
nand U38813 (N_38813,N_38717,N_38684);
nor U38814 (N_38814,N_38737,N_38501);
xor U38815 (N_38815,N_38580,N_38698);
nor U38816 (N_38816,N_38506,N_38674);
nand U38817 (N_38817,N_38718,N_38747);
xnor U38818 (N_38818,N_38535,N_38634);
nor U38819 (N_38819,N_38743,N_38660);
xor U38820 (N_38820,N_38744,N_38510);
nand U38821 (N_38821,N_38695,N_38587);
nand U38822 (N_38822,N_38739,N_38524);
nor U38823 (N_38823,N_38571,N_38697);
and U38824 (N_38824,N_38632,N_38746);
and U38825 (N_38825,N_38505,N_38683);
nor U38826 (N_38826,N_38502,N_38716);
nand U38827 (N_38827,N_38551,N_38609);
and U38828 (N_38828,N_38685,N_38527);
nor U38829 (N_38829,N_38656,N_38729);
and U38830 (N_38830,N_38618,N_38673);
xnor U38831 (N_38831,N_38563,N_38537);
nand U38832 (N_38832,N_38630,N_38598);
nor U38833 (N_38833,N_38699,N_38558);
and U38834 (N_38834,N_38518,N_38736);
nor U38835 (N_38835,N_38689,N_38542);
nor U38836 (N_38836,N_38605,N_38540);
nand U38837 (N_38837,N_38611,N_38708);
and U38838 (N_38838,N_38665,N_38570);
nor U38839 (N_38839,N_38642,N_38728);
or U38840 (N_38840,N_38607,N_38612);
xor U38841 (N_38841,N_38738,N_38701);
nand U38842 (N_38842,N_38589,N_38603);
or U38843 (N_38843,N_38600,N_38582);
nor U38844 (N_38844,N_38635,N_38653);
xor U38845 (N_38845,N_38617,N_38633);
and U38846 (N_38846,N_38554,N_38568);
nor U38847 (N_38847,N_38508,N_38601);
nor U38848 (N_38848,N_38713,N_38678);
and U38849 (N_38849,N_38596,N_38710);
and U38850 (N_38850,N_38693,N_38667);
nor U38851 (N_38851,N_38528,N_38749);
nand U38852 (N_38852,N_38604,N_38610);
or U38853 (N_38853,N_38556,N_38681);
xnor U38854 (N_38854,N_38575,N_38526);
xnor U38855 (N_38855,N_38591,N_38595);
and U38856 (N_38856,N_38583,N_38730);
nor U38857 (N_38857,N_38621,N_38732);
or U38858 (N_38858,N_38588,N_38515);
xnor U38859 (N_38859,N_38723,N_38559);
and U38860 (N_38860,N_38606,N_38530);
or U38861 (N_38861,N_38658,N_38659);
nand U38862 (N_38862,N_38688,N_38614);
xnor U38863 (N_38863,N_38628,N_38562);
or U38864 (N_38864,N_38579,N_38624);
nor U38865 (N_38865,N_38585,N_38706);
xnor U38866 (N_38866,N_38700,N_38668);
nand U38867 (N_38867,N_38590,N_38671);
and U38868 (N_38868,N_38576,N_38639);
nor U38869 (N_38869,N_38694,N_38707);
xor U38870 (N_38870,N_38555,N_38719);
or U38871 (N_38871,N_38544,N_38615);
and U38872 (N_38872,N_38520,N_38643);
nand U38873 (N_38873,N_38721,N_38651);
nand U38874 (N_38874,N_38649,N_38509);
or U38875 (N_38875,N_38677,N_38706);
or U38876 (N_38876,N_38518,N_38657);
or U38877 (N_38877,N_38524,N_38726);
xor U38878 (N_38878,N_38628,N_38679);
nand U38879 (N_38879,N_38675,N_38577);
nor U38880 (N_38880,N_38608,N_38631);
nor U38881 (N_38881,N_38517,N_38671);
xnor U38882 (N_38882,N_38713,N_38564);
nand U38883 (N_38883,N_38572,N_38513);
nand U38884 (N_38884,N_38688,N_38537);
nand U38885 (N_38885,N_38683,N_38658);
nand U38886 (N_38886,N_38610,N_38568);
xnor U38887 (N_38887,N_38668,N_38691);
and U38888 (N_38888,N_38670,N_38577);
xor U38889 (N_38889,N_38572,N_38510);
nand U38890 (N_38890,N_38649,N_38641);
xor U38891 (N_38891,N_38507,N_38749);
xnor U38892 (N_38892,N_38525,N_38524);
nor U38893 (N_38893,N_38697,N_38600);
nand U38894 (N_38894,N_38559,N_38685);
and U38895 (N_38895,N_38720,N_38638);
or U38896 (N_38896,N_38664,N_38513);
nor U38897 (N_38897,N_38594,N_38587);
nor U38898 (N_38898,N_38564,N_38623);
xor U38899 (N_38899,N_38724,N_38623);
and U38900 (N_38900,N_38691,N_38660);
nand U38901 (N_38901,N_38566,N_38550);
and U38902 (N_38902,N_38662,N_38635);
or U38903 (N_38903,N_38605,N_38541);
xor U38904 (N_38904,N_38511,N_38726);
xnor U38905 (N_38905,N_38565,N_38740);
nand U38906 (N_38906,N_38591,N_38574);
or U38907 (N_38907,N_38639,N_38749);
nand U38908 (N_38908,N_38742,N_38547);
xor U38909 (N_38909,N_38570,N_38722);
nor U38910 (N_38910,N_38654,N_38604);
nand U38911 (N_38911,N_38744,N_38601);
and U38912 (N_38912,N_38668,N_38704);
and U38913 (N_38913,N_38660,N_38713);
and U38914 (N_38914,N_38538,N_38696);
xnor U38915 (N_38915,N_38590,N_38523);
and U38916 (N_38916,N_38513,N_38620);
and U38917 (N_38917,N_38579,N_38649);
or U38918 (N_38918,N_38663,N_38687);
nand U38919 (N_38919,N_38606,N_38583);
xor U38920 (N_38920,N_38641,N_38521);
or U38921 (N_38921,N_38572,N_38691);
or U38922 (N_38922,N_38562,N_38541);
xnor U38923 (N_38923,N_38671,N_38544);
nand U38924 (N_38924,N_38528,N_38735);
xor U38925 (N_38925,N_38692,N_38639);
xnor U38926 (N_38926,N_38623,N_38583);
nor U38927 (N_38927,N_38686,N_38670);
nand U38928 (N_38928,N_38656,N_38631);
xor U38929 (N_38929,N_38620,N_38689);
or U38930 (N_38930,N_38529,N_38701);
xor U38931 (N_38931,N_38663,N_38505);
or U38932 (N_38932,N_38614,N_38549);
and U38933 (N_38933,N_38554,N_38749);
or U38934 (N_38934,N_38613,N_38538);
nand U38935 (N_38935,N_38674,N_38676);
nand U38936 (N_38936,N_38736,N_38650);
nand U38937 (N_38937,N_38625,N_38559);
nand U38938 (N_38938,N_38598,N_38613);
nor U38939 (N_38939,N_38510,N_38606);
nand U38940 (N_38940,N_38646,N_38528);
nor U38941 (N_38941,N_38618,N_38691);
and U38942 (N_38942,N_38593,N_38710);
and U38943 (N_38943,N_38628,N_38534);
xnor U38944 (N_38944,N_38732,N_38631);
nand U38945 (N_38945,N_38580,N_38517);
and U38946 (N_38946,N_38584,N_38655);
and U38947 (N_38947,N_38509,N_38547);
nor U38948 (N_38948,N_38649,N_38553);
or U38949 (N_38949,N_38697,N_38502);
xor U38950 (N_38950,N_38595,N_38749);
nand U38951 (N_38951,N_38728,N_38714);
xor U38952 (N_38952,N_38613,N_38586);
or U38953 (N_38953,N_38683,N_38626);
nor U38954 (N_38954,N_38696,N_38628);
nand U38955 (N_38955,N_38659,N_38730);
nand U38956 (N_38956,N_38547,N_38677);
nand U38957 (N_38957,N_38716,N_38613);
xnor U38958 (N_38958,N_38649,N_38685);
or U38959 (N_38959,N_38665,N_38692);
and U38960 (N_38960,N_38734,N_38744);
and U38961 (N_38961,N_38585,N_38502);
nor U38962 (N_38962,N_38568,N_38555);
or U38963 (N_38963,N_38504,N_38530);
nand U38964 (N_38964,N_38540,N_38601);
and U38965 (N_38965,N_38666,N_38564);
and U38966 (N_38966,N_38594,N_38573);
nor U38967 (N_38967,N_38619,N_38693);
nor U38968 (N_38968,N_38513,N_38694);
nand U38969 (N_38969,N_38501,N_38562);
xnor U38970 (N_38970,N_38692,N_38699);
xnor U38971 (N_38971,N_38661,N_38646);
nor U38972 (N_38972,N_38593,N_38617);
or U38973 (N_38973,N_38715,N_38732);
nand U38974 (N_38974,N_38560,N_38631);
and U38975 (N_38975,N_38626,N_38663);
nand U38976 (N_38976,N_38737,N_38619);
xor U38977 (N_38977,N_38648,N_38667);
nand U38978 (N_38978,N_38546,N_38574);
nand U38979 (N_38979,N_38650,N_38526);
or U38980 (N_38980,N_38541,N_38737);
or U38981 (N_38981,N_38506,N_38690);
nor U38982 (N_38982,N_38651,N_38598);
nand U38983 (N_38983,N_38685,N_38548);
nand U38984 (N_38984,N_38713,N_38728);
nand U38985 (N_38985,N_38571,N_38629);
nand U38986 (N_38986,N_38613,N_38542);
and U38987 (N_38987,N_38517,N_38565);
and U38988 (N_38988,N_38502,N_38685);
xor U38989 (N_38989,N_38608,N_38647);
or U38990 (N_38990,N_38748,N_38687);
xor U38991 (N_38991,N_38579,N_38739);
xnor U38992 (N_38992,N_38721,N_38643);
or U38993 (N_38993,N_38643,N_38687);
and U38994 (N_38994,N_38534,N_38538);
nor U38995 (N_38995,N_38641,N_38555);
and U38996 (N_38996,N_38704,N_38739);
and U38997 (N_38997,N_38735,N_38741);
or U38998 (N_38998,N_38593,N_38520);
or U38999 (N_38999,N_38645,N_38706);
xor U39000 (N_39000,N_38763,N_38784);
nor U39001 (N_39001,N_38987,N_38884);
and U39002 (N_39002,N_38762,N_38998);
and U39003 (N_39003,N_38855,N_38807);
xnor U39004 (N_39004,N_38859,N_38983);
or U39005 (N_39005,N_38902,N_38873);
nor U39006 (N_39006,N_38792,N_38759);
xnor U39007 (N_39007,N_38797,N_38803);
or U39008 (N_39008,N_38761,N_38949);
nor U39009 (N_39009,N_38903,N_38913);
and U39010 (N_39010,N_38918,N_38965);
or U39011 (N_39011,N_38769,N_38868);
xor U39012 (N_39012,N_38930,N_38989);
xnor U39013 (N_39013,N_38799,N_38962);
nor U39014 (N_39014,N_38751,N_38959);
and U39015 (N_39015,N_38975,N_38856);
nand U39016 (N_39016,N_38924,N_38900);
or U39017 (N_39017,N_38804,N_38914);
and U39018 (N_39018,N_38828,N_38781);
xnor U39019 (N_39019,N_38775,N_38858);
nand U39020 (N_39020,N_38844,N_38752);
and U39021 (N_39021,N_38888,N_38841);
or U39022 (N_39022,N_38936,N_38907);
nand U39023 (N_39023,N_38942,N_38860);
and U39024 (N_39024,N_38765,N_38866);
or U39025 (N_39025,N_38820,N_38978);
or U39026 (N_39026,N_38847,N_38849);
and U39027 (N_39027,N_38899,N_38883);
xor U39028 (N_39028,N_38819,N_38980);
or U39029 (N_39029,N_38995,N_38864);
nand U39030 (N_39030,N_38810,N_38985);
and U39031 (N_39031,N_38920,N_38910);
xnor U39032 (N_39032,N_38808,N_38970);
xnor U39033 (N_39033,N_38997,N_38906);
nand U39034 (N_39034,N_38824,N_38778);
or U39035 (N_39035,N_38948,N_38986);
nor U39036 (N_39036,N_38893,N_38785);
xnor U39037 (N_39037,N_38954,N_38815);
nand U39038 (N_39038,N_38938,N_38935);
xor U39039 (N_39039,N_38836,N_38791);
and U39040 (N_39040,N_38939,N_38817);
or U39041 (N_39041,N_38961,N_38904);
nand U39042 (N_39042,N_38922,N_38905);
or U39043 (N_39043,N_38839,N_38779);
nor U39044 (N_39044,N_38890,N_38827);
or U39045 (N_39045,N_38974,N_38758);
nor U39046 (N_39046,N_38812,N_38943);
and U39047 (N_39047,N_38934,N_38821);
or U39048 (N_39048,N_38921,N_38843);
xor U39049 (N_39049,N_38805,N_38816);
and U39050 (N_39050,N_38916,N_38862);
and U39051 (N_39051,N_38981,N_38990);
and U39052 (N_39052,N_38760,N_38867);
or U39053 (N_39053,N_38915,N_38952);
nor U39054 (N_39054,N_38848,N_38796);
nor U39055 (N_39055,N_38857,N_38953);
nor U39056 (N_39056,N_38994,N_38876);
nor U39057 (N_39057,N_38988,N_38802);
xnor U39058 (N_39058,N_38957,N_38929);
xnor U39059 (N_39059,N_38754,N_38901);
xor U39060 (N_39060,N_38895,N_38753);
or U39061 (N_39061,N_38854,N_38911);
nand U39062 (N_39062,N_38880,N_38830);
nor U39063 (N_39063,N_38833,N_38832);
nor U39064 (N_39064,N_38840,N_38772);
and U39065 (N_39065,N_38960,N_38941);
and U39066 (N_39066,N_38874,N_38813);
or U39067 (N_39067,N_38823,N_38842);
and U39068 (N_39068,N_38966,N_38885);
or U39069 (N_39069,N_38976,N_38798);
or U39070 (N_39070,N_38909,N_38897);
xnor U39071 (N_39071,N_38818,N_38825);
and U39072 (N_39072,N_38889,N_38877);
nor U39073 (N_39073,N_38756,N_38996);
nor U39074 (N_39074,N_38834,N_38919);
nor U39075 (N_39075,N_38984,N_38958);
nand U39076 (N_39076,N_38956,N_38879);
and U39077 (N_39077,N_38882,N_38853);
nand U39078 (N_39078,N_38999,N_38972);
nand U39079 (N_39079,N_38871,N_38932);
and U39080 (N_39080,N_38845,N_38992);
and U39081 (N_39081,N_38814,N_38928);
or U39082 (N_39082,N_38969,N_38806);
nand U39083 (N_39083,N_38837,N_38771);
nand U39084 (N_39084,N_38982,N_38773);
or U39085 (N_39085,N_38933,N_38795);
and U39086 (N_39086,N_38822,N_38755);
xor U39087 (N_39087,N_38863,N_38835);
nor U39088 (N_39088,N_38967,N_38898);
and U39089 (N_39089,N_38782,N_38878);
or U39090 (N_39090,N_38777,N_38931);
and U39091 (N_39091,N_38783,N_38977);
nand U39092 (N_39092,N_38945,N_38892);
nor U39093 (N_39093,N_38894,N_38951);
nor U39094 (N_39094,N_38846,N_38927);
xor U39095 (N_39095,N_38800,N_38908);
nor U39096 (N_39096,N_38912,N_38869);
nand U39097 (N_39097,N_38809,N_38979);
nor U39098 (N_39098,N_38770,N_38964);
or U39099 (N_39099,N_38787,N_38946);
or U39100 (N_39100,N_38790,N_38944);
xor U39101 (N_39101,N_38950,N_38923);
nand U39102 (N_39102,N_38764,N_38793);
xnor U39103 (N_39103,N_38786,N_38870);
and U39104 (N_39104,N_38774,N_38750);
and U39105 (N_39105,N_38872,N_38851);
or U39106 (N_39106,N_38766,N_38757);
and U39107 (N_39107,N_38937,N_38973);
or U39108 (N_39108,N_38917,N_38780);
or U39109 (N_39109,N_38852,N_38865);
and U39110 (N_39110,N_38991,N_38850);
xor U39111 (N_39111,N_38789,N_38794);
or U39112 (N_39112,N_38891,N_38896);
nand U39113 (N_39113,N_38955,N_38925);
and U39114 (N_39114,N_38801,N_38971);
nand U39115 (N_39115,N_38768,N_38926);
or U39116 (N_39116,N_38767,N_38940);
nand U39117 (N_39117,N_38963,N_38826);
and U39118 (N_39118,N_38838,N_38886);
or U39119 (N_39119,N_38776,N_38861);
or U39120 (N_39120,N_38881,N_38829);
nor U39121 (N_39121,N_38831,N_38887);
xor U39122 (N_39122,N_38947,N_38811);
nand U39123 (N_39123,N_38968,N_38875);
nand U39124 (N_39124,N_38788,N_38993);
nand U39125 (N_39125,N_38867,N_38778);
nand U39126 (N_39126,N_38993,N_38875);
or U39127 (N_39127,N_38798,N_38778);
or U39128 (N_39128,N_38934,N_38899);
and U39129 (N_39129,N_38880,N_38966);
nor U39130 (N_39130,N_38953,N_38779);
nand U39131 (N_39131,N_38958,N_38783);
and U39132 (N_39132,N_38831,N_38789);
xor U39133 (N_39133,N_38763,N_38920);
or U39134 (N_39134,N_38996,N_38811);
nand U39135 (N_39135,N_38835,N_38918);
or U39136 (N_39136,N_38936,N_38978);
nand U39137 (N_39137,N_38962,N_38828);
or U39138 (N_39138,N_38773,N_38948);
or U39139 (N_39139,N_38880,N_38791);
and U39140 (N_39140,N_38804,N_38907);
nand U39141 (N_39141,N_38865,N_38888);
nor U39142 (N_39142,N_38803,N_38821);
nand U39143 (N_39143,N_38756,N_38900);
or U39144 (N_39144,N_38827,N_38868);
and U39145 (N_39145,N_38922,N_38868);
xnor U39146 (N_39146,N_38809,N_38900);
and U39147 (N_39147,N_38884,N_38842);
and U39148 (N_39148,N_38852,N_38985);
nor U39149 (N_39149,N_38869,N_38969);
xnor U39150 (N_39150,N_38806,N_38830);
and U39151 (N_39151,N_38757,N_38760);
xor U39152 (N_39152,N_38845,N_38885);
nand U39153 (N_39153,N_38909,N_38808);
xor U39154 (N_39154,N_38791,N_38766);
xor U39155 (N_39155,N_38754,N_38991);
nor U39156 (N_39156,N_38787,N_38923);
or U39157 (N_39157,N_38980,N_38759);
nor U39158 (N_39158,N_38781,N_38888);
or U39159 (N_39159,N_38779,N_38798);
nor U39160 (N_39160,N_38772,N_38984);
xnor U39161 (N_39161,N_38777,N_38972);
nor U39162 (N_39162,N_38770,N_38942);
xnor U39163 (N_39163,N_38972,N_38966);
nand U39164 (N_39164,N_38959,N_38984);
nor U39165 (N_39165,N_38935,N_38761);
or U39166 (N_39166,N_38943,N_38763);
nor U39167 (N_39167,N_38841,N_38756);
xnor U39168 (N_39168,N_38868,N_38791);
nand U39169 (N_39169,N_38846,N_38980);
or U39170 (N_39170,N_38957,N_38857);
and U39171 (N_39171,N_38878,N_38791);
nand U39172 (N_39172,N_38962,N_38993);
nand U39173 (N_39173,N_38792,N_38835);
and U39174 (N_39174,N_38955,N_38785);
xnor U39175 (N_39175,N_38940,N_38950);
nor U39176 (N_39176,N_38871,N_38850);
or U39177 (N_39177,N_38862,N_38995);
and U39178 (N_39178,N_38788,N_38850);
or U39179 (N_39179,N_38878,N_38794);
xor U39180 (N_39180,N_38973,N_38914);
or U39181 (N_39181,N_38847,N_38832);
xor U39182 (N_39182,N_38950,N_38879);
nand U39183 (N_39183,N_38928,N_38760);
and U39184 (N_39184,N_38939,N_38941);
nand U39185 (N_39185,N_38806,N_38910);
nand U39186 (N_39186,N_38944,N_38991);
xnor U39187 (N_39187,N_38791,N_38901);
xor U39188 (N_39188,N_38809,N_38844);
nand U39189 (N_39189,N_38937,N_38928);
or U39190 (N_39190,N_38867,N_38790);
nor U39191 (N_39191,N_38983,N_38791);
or U39192 (N_39192,N_38779,N_38879);
xor U39193 (N_39193,N_38888,N_38956);
or U39194 (N_39194,N_38802,N_38920);
and U39195 (N_39195,N_38918,N_38913);
nor U39196 (N_39196,N_38884,N_38928);
xnor U39197 (N_39197,N_38979,N_38832);
or U39198 (N_39198,N_38800,N_38874);
nor U39199 (N_39199,N_38854,N_38982);
nand U39200 (N_39200,N_38877,N_38866);
nor U39201 (N_39201,N_38866,N_38792);
xnor U39202 (N_39202,N_38793,N_38837);
xor U39203 (N_39203,N_38780,N_38953);
and U39204 (N_39204,N_38942,N_38990);
nand U39205 (N_39205,N_38772,N_38943);
xor U39206 (N_39206,N_38821,N_38893);
nand U39207 (N_39207,N_38751,N_38912);
nand U39208 (N_39208,N_38855,N_38779);
or U39209 (N_39209,N_38846,N_38789);
or U39210 (N_39210,N_38922,N_38862);
nand U39211 (N_39211,N_38935,N_38754);
nor U39212 (N_39212,N_38970,N_38871);
xor U39213 (N_39213,N_38845,N_38801);
and U39214 (N_39214,N_38898,N_38943);
and U39215 (N_39215,N_38818,N_38887);
xnor U39216 (N_39216,N_38952,N_38770);
and U39217 (N_39217,N_38839,N_38939);
and U39218 (N_39218,N_38952,N_38971);
nor U39219 (N_39219,N_38795,N_38848);
nor U39220 (N_39220,N_38996,N_38896);
nand U39221 (N_39221,N_38801,N_38985);
nor U39222 (N_39222,N_38838,N_38837);
or U39223 (N_39223,N_38914,N_38760);
nor U39224 (N_39224,N_38902,N_38777);
or U39225 (N_39225,N_38922,N_38860);
xnor U39226 (N_39226,N_38767,N_38768);
xnor U39227 (N_39227,N_38990,N_38886);
nor U39228 (N_39228,N_38807,N_38844);
or U39229 (N_39229,N_38934,N_38907);
nor U39230 (N_39230,N_38761,N_38836);
xor U39231 (N_39231,N_38750,N_38804);
xor U39232 (N_39232,N_38848,N_38886);
nor U39233 (N_39233,N_38954,N_38941);
xnor U39234 (N_39234,N_38986,N_38880);
and U39235 (N_39235,N_38766,N_38952);
or U39236 (N_39236,N_38786,N_38992);
nand U39237 (N_39237,N_38934,N_38768);
or U39238 (N_39238,N_38908,N_38858);
xor U39239 (N_39239,N_38984,N_38970);
nor U39240 (N_39240,N_38844,N_38947);
and U39241 (N_39241,N_38860,N_38838);
nor U39242 (N_39242,N_38769,N_38815);
xor U39243 (N_39243,N_38996,N_38779);
nand U39244 (N_39244,N_38827,N_38903);
nor U39245 (N_39245,N_38969,N_38771);
nor U39246 (N_39246,N_38794,N_38854);
xnor U39247 (N_39247,N_38985,N_38802);
nor U39248 (N_39248,N_38751,N_38990);
xor U39249 (N_39249,N_38840,N_38803);
xor U39250 (N_39250,N_39227,N_39242);
and U39251 (N_39251,N_39166,N_39116);
and U39252 (N_39252,N_39169,N_39104);
nand U39253 (N_39253,N_39066,N_39143);
or U39254 (N_39254,N_39076,N_39014);
or U39255 (N_39255,N_39145,N_39004);
nor U39256 (N_39256,N_39086,N_39148);
or U39257 (N_39257,N_39056,N_39247);
nand U39258 (N_39258,N_39174,N_39065);
xor U39259 (N_39259,N_39141,N_39200);
and U39260 (N_39260,N_39221,N_39126);
and U39261 (N_39261,N_39155,N_39090);
nand U39262 (N_39262,N_39098,N_39198);
nor U39263 (N_39263,N_39167,N_39186);
nor U39264 (N_39264,N_39027,N_39151);
or U39265 (N_39265,N_39049,N_39134);
nor U39266 (N_39266,N_39067,N_39108);
nor U39267 (N_39267,N_39006,N_39159);
xnor U39268 (N_39268,N_39222,N_39057);
xor U39269 (N_39269,N_39038,N_39007);
or U39270 (N_39270,N_39241,N_39017);
xnor U39271 (N_39271,N_39030,N_39059);
xnor U39272 (N_39272,N_39081,N_39226);
xnor U39273 (N_39273,N_39153,N_39248);
nand U39274 (N_39274,N_39101,N_39249);
and U39275 (N_39275,N_39084,N_39190);
xnor U39276 (N_39276,N_39161,N_39185);
nand U39277 (N_39277,N_39183,N_39233);
nand U39278 (N_39278,N_39131,N_39188);
xnor U39279 (N_39279,N_39130,N_39121);
nor U39280 (N_39280,N_39100,N_39064);
or U39281 (N_39281,N_39205,N_39078);
and U39282 (N_39282,N_39018,N_39207);
nor U39283 (N_39283,N_39041,N_39176);
or U39284 (N_39284,N_39193,N_39127);
and U39285 (N_39285,N_39039,N_39094);
nor U39286 (N_39286,N_39036,N_39058);
and U39287 (N_39287,N_39063,N_39000);
nor U39288 (N_39288,N_39154,N_39011);
xnor U39289 (N_39289,N_39146,N_39005);
nor U39290 (N_39290,N_39157,N_39234);
or U39291 (N_39291,N_39105,N_39070);
xor U39292 (N_39292,N_39228,N_39085);
nand U39293 (N_39293,N_39016,N_39182);
and U39294 (N_39294,N_39158,N_39211);
and U39295 (N_39295,N_39135,N_39229);
nor U39296 (N_39296,N_39220,N_39195);
or U39297 (N_39297,N_39140,N_39118);
xnor U39298 (N_39298,N_39162,N_39173);
xnor U39299 (N_39299,N_39034,N_39003);
nand U39300 (N_39300,N_39156,N_39061);
nor U39301 (N_39301,N_39212,N_39133);
nand U39302 (N_39302,N_39037,N_39075);
xor U39303 (N_39303,N_39050,N_39232);
or U39304 (N_39304,N_39123,N_39028);
or U39305 (N_39305,N_39107,N_39015);
nor U39306 (N_39306,N_39072,N_39128);
nor U39307 (N_39307,N_39223,N_39053);
nor U39308 (N_39308,N_39138,N_39119);
nand U39309 (N_39309,N_39165,N_39106);
nand U39310 (N_39310,N_39178,N_39199);
or U39311 (N_39311,N_39111,N_39042);
or U39312 (N_39312,N_39020,N_39073);
or U39313 (N_39313,N_39093,N_39026);
nor U39314 (N_39314,N_39044,N_39088);
nand U39315 (N_39315,N_39087,N_39150);
and U39316 (N_39316,N_39060,N_39139);
or U39317 (N_39317,N_39021,N_39208);
nand U39318 (N_39318,N_39092,N_39068);
or U39319 (N_39319,N_39206,N_39160);
xor U39320 (N_39320,N_39201,N_39080);
nand U39321 (N_39321,N_39112,N_39124);
or U39322 (N_39322,N_39191,N_39051);
nor U39323 (N_39323,N_39091,N_39180);
nand U39324 (N_39324,N_39244,N_39192);
xnor U39325 (N_39325,N_39102,N_39025);
and U39326 (N_39326,N_39024,N_39032);
xor U39327 (N_39327,N_39202,N_39132);
or U39328 (N_39328,N_39008,N_39079);
or U39329 (N_39329,N_39196,N_39137);
and U39330 (N_39330,N_39109,N_39043);
nor U39331 (N_39331,N_39069,N_39194);
nor U39332 (N_39332,N_39187,N_39113);
xnor U39333 (N_39333,N_39235,N_39055);
and U39334 (N_39334,N_39103,N_39013);
nor U39335 (N_39335,N_39129,N_39033);
and U39336 (N_39336,N_39114,N_39164);
xnor U39337 (N_39337,N_39149,N_39074);
nand U39338 (N_39338,N_39239,N_39009);
and U39339 (N_39339,N_39095,N_39179);
nor U39340 (N_39340,N_39082,N_39031);
xor U39341 (N_39341,N_39181,N_39010);
nor U39342 (N_39342,N_39177,N_39225);
nand U39343 (N_39343,N_39122,N_39046);
and U39344 (N_39344,N_39152,N_39172);
or U39345 (N_39345,N_39052,N_39029);
nand U39346 (N_39346,N_39184,N_39035);
nand U39347 (N_39347,N_39217,N_39083);
nor U39348 (N_39348,N_39231,N_39045);
and U39349 (N_39349,N_39230,N_39048);
nor U39350 (N_39350,N_39213,N_39023);
and U39351 (N_39351,N_39209,N_39175);
xnor U39352 (N_39352,N_39246,N_39089);
xnor U39353 (N_39353,N_39022,N_39215);
nand U39354 (N_39354,N_39054,N_39071);
nor U39355 (N_39355,N_39163,N_39243);
nor U39356 (N_39356,N_39117,N_39245);
nand U39357 (N_39357,N_39189,N_39218);
nand U39358 (N_39358,N_39099,N_39197);
nand U39359 (N_39359,N_39040,N_39019);
nor U39360 (N_39360,N_39110,N_39002);
and U39361 (N_39361,N_39115,N_39204);
nand U39362 (N_39362,N_39224,N_39170);
and U39363 (N_39363,N_39238,N_39125);
xor U39364 (N_39364,N_39001,N_39062);
xor U39365 (N_39365,N_39012,N_39214);
nand U39366 (N_39366,N_39142,N_39077);
nand U39367 (N_39367,N_39219,N_39240);
nand U39368 (N_39368,N_39120,N_39236);
and U39369 (N_39369,N_39210,N_39237);
xnor U39370 (N_39370,N_39144,N_39203);
and U39371 (N_39371,N_39047,N_39168);
nand U39372 (N_39372,N_39216,N_39136);
or U39373 (N_39373,N_39096,N_39147);
xnor U39374 (N_39374,N_39097,N_39171);
nand U39375 (N_39375,N_39030,N_39072);
xor U39376 (N_39376,N_39084,N_39086);
and U39377 (N_39377,N_39121,N_39066);
nand U39378 (N_39378,N_39011,N_39083);
nor U39379 (N_39379,N_39204,N_39032);
xor U39380 (N_39380,N_39087,N_39035);
nand U39381 (N_39381,N_39190,N_39164);
nor U39382 (N_39382,N_39184,N_39036);
nand U39383 (N_39383,N_39172,N_39133);
or U39384 (N_39384,N_39044,N_39080);
and U39385 (N_39385,N_39035,N_39211);
or U39386 (N_39386,N_39131,N_39035);
nor U39387 (N_39387,N_39178,N_39098);
or U39388 (N_39388,N_39180,N_39114);
nand U39389 (N_39389,N_39161,N_39100);
nor U39390 (N_39390,N_39036,N_39055);
and U39391 (N_39391,N_39211,N_39145);
nand U39392 (N_39392,N_39023,N_39050);
and U39393 (N_39393,N_39098,N_39044);
or U39394 (N_39394,N_39112,N_39171);
or U39395 (N_39395,N_39139,N_39021);
nand U39396 (N_39396,N_39124,N_39109);
nand U39397 (N_39397,N_39197,N_39175);
and U39398 (N_39398,N_39026,N_39033);
or U39399 (N_39399,N_39044,N_39126);
and U39400 (N_39400,N_39165,N_39167);
and U39401 (N_39401,N_39042,N_39133);
xnor U39402 (N_39402,N_39006,N_39095);
or U39403 (N_39403,N_39090,N_39179);
nand U39404 (N_39404,N_39226,N_39234);
and U39405 (N_39405,N_39147,N_39011);
or U39406 (N_39406,N_39201,N_39109);
nand U39407 (N_39407,N_39170,N_39200);
nand U39408 (N_39408,N_39031,N_39229);
nand U39409 (N_39409,N_39068,N_39019);
xnor U39410 (N_39410,N_39051,N_39230);
and U39411 (N_39411,N_39104,N_39005);
and U39412 (N_39412,N_39125,N_39137);
xor U39413 (N_39413,N_39024,N_39100);
nand U39414 (N_39414,N_39181,N_39105);
nor U39415 (N_39415,N_39035,N_39011);
nand U39416 (N_39416,N_39088,N_39049);
nor U39417 (N_39417,N_39088,N_39164);
and U39418 (N_39418,N_39001,N_39153);
and U39419 (N_39419,N_39012,N_39075);
nor U39420 (N_39420,N_39054,N_39228);
nor U39421 (N_39421,N_39107,N_39020);
xnor U39422 (N_39422,N_39228,N_39009);
nand U39423 (N_39423,N_39101,N_39109);
xnor U39424 (N_39424,N_39215,N_39234);
or U39425 (N_39425,N_39248,N_39017);
xnor U39426 (N_39426,N_39030,N_39104);
nor U39427 (N_39427,N_39028,N_39052);
xor U39428 (N_39428,N_39176,N_39229);
nand U39429 (N_39429,N_39015,N_39127);
xor U39430 (N_39430,N_39072,N_39163);
and U39431 (N_39431,N_39061,N_39095);
and U39432 (N_39432,N_39107,N_39234);
or U39433 (N_39433,N_39033,N_39109);
and U39434 (N_39434,N_39036,N_39142);
xnor U39435 (N_39435,N_39246,N_39151);
or U39436 (N_39436,N_39063,N_39028);
or U39437 (N_39437,N_39247,N_39097);
nand U39438 (N_39438,N_39106,N_39017);
xnor U39439 (N_39439,N_39124,N_39079);
nand U39440 (N_39440,N_39153,N_39099);
nor U39441 (N_39441,N_39066,N_39217);
and U39442 (N_39442,N_39031,N_39208);
nor U39443 (N_39443,N_39055,N_39107);
or U39444 (N_39444,N_39190,N_39105);
or U39445 (N_39445,N_39035,N_39138);
nand U39446 (N_39446,N_39102,N_39232);
nand U39447 (N_39447,N_39051,N_39236);
xor U39448 (N_39448,N_39116,N_39030);
nor U39449 (N_39449,N_39102,N_39045);
xnor U39450 (N_39450,N_39018,N_39178);
nor U39451 (N_39451,N_39102,N_39060);
nor U39452 (N_39452,N_39111,N_39062);
nor U39453 (N_39453,N_39142,N_39188);
xnor U39454 (N_39454,N_39210,N_39038);
nand U39455 (N_39455,N_39232,N_39190);
or U39456 (N_39456,N_39111,N_39165);
and U39457 (N_39457,N_39110,N_39142);
or U39458 (N_39458,N_39223,N_39071);
nor U39459 (N_39459,N_39218,N_39118);
xnor U39460 (N_39460,N_39184,N_39030);
nand U39461 (N_39461,N_39040,N_39111);
nor U39462 (N_39462,N_39102,N_39247);
and U39463 (N_39463,N_39143,N_39021);
nor U39464 (N_39464,N_39047,N_39113);
and U39465 (N_39465,N_39120,N_39233);
xnor U39466 (N_39466,N_39014,N_39010);
nor U39467 (N_39467,N_39211,N_39207);
and U39468 (N_39468,N_39244,N_39145);
and U39469 (N_39469,N_39074,N_39196);
nand U39470 (N_39470,N_39077,N_39048);
or U39471 (N_39471,N_39020,N_39005);
xnor U39472 (N_39472,N_39185,N_39012);
nor U39473 (N_39473,N_39039,N_39149);
and U39474 (N_39474,N_39098,N_39126);
nand U39475 (N_39475,N_39020,N_39180);
xor U39476 (N_39476,N_39203,N_39066);
or U39477 (N_39477,N_39089,N_39006);
and U39478 (N_39478,N_39199,N_39099);
and U39479 (N_39479,N_39124,N_39078);
and U39480 (N_39480,N_39196,N_39235);
or U39481 (N_39481,N_39069,N_39021);
and U39482 (N_39482,N_39244,N_39089);
nand U39483 (N_39483,N_39229,N_39215);
nor U39484 (N_39484,N_39169,N_39167);
or U39485 (N_39485,N_39177,N_39001);
nand U39486 (N_39486,N_39136,N_39022);
nand U39487 (N_39487,N_39007,N_39207);
xor U39488 (N_39488,N_39065,N_39116);
and U39489 (N_39489,N_39208,N_39164);
or U39490 (N_39490,N_39215,N_39028);
or U39491 (N_39491,N_39110,N_39241);
nor U39492 (N_39492,N_39188,N_39079);
or U39493 (N_39493,N_39004,N_39084);
xor U39494 (N_39494,N_39080,N_39046);
xnor U39495 (N_39495,N_39202,N_39146);
nand U39496 (N_39496,N_39228,N_39052);
or U39497 (N_39497,N_39063,N_39219);
nor U39498 (N_39498,N_39199,N_39105);
nand U39499 (N_39499,N_39140,N_39012);
nand U39500 (N_39500,N_39494,N_39492);
and U39501 (N_39501,N_39469,N_39320);
or U39502 (N_39502,N_39266,N_39422);
nor U39503 (N_39503,N_39263,N_39351);
and U39504 (N_39504,N_39375,N_39466);
nor U39505 (N_39505,N_39497,N_39420);
or U39506 (N_39506,N_39419,N_39468);
nand U39507 (N_39507,N_39450,N_39486);
nand U39508 (N_39508,N_39369,N_39341);
xor U39509 (N_39509,N_39355,N_39253);
or U39510 (N_39510,N_39289,N_39410);
nor U39511 (N_39511,N_39498,N_39275);
nor U39512 (N_39512,N_39380,N_39405);
or U39513 (N_39513,N_39311,N_39386);
or U39514 (N_39514,N_39315,N_39269);
nor U39515 (N_39515,N_39377,N_39361);
nand U39516 (N_39516,N_39448,N_39424);
nor U39517 (N_39517,N_39276,N_39324);
nor U39518 (N_39518,N_39251,N_39307);
and U39519 (N_39519,N_39303,N_39490);
or U39520 (N_39520,N_39401,N_39270);
or U39521 (N_39521,N_39316,N_39476);
and U39522 (N_39522,N_39328,N_39478);
nand U39523 (N_39523,N_39383,N_39406);
nor U39524 (N_39524,N_39400,N_39274);
nand U39525 (N_39525,N_39317,N_39321);
nand U39526 (N_39526,N_39449,N_39398);
xor U39527 (N_39527,N_39396,N_39447);
xnor U39528 (N_39528,N_39337,N_39338);
xor U39529 (N_39529,N_39363,N_39425);
and U39530 (N_39530,N_39254,N_39479);
nand U39531 (N_39531,N_39451,N_39305);
xnor U39532 (N_39532,N_39314,N_39257);
and U39533 (N_39533,N_39368,N_39376);
and U39534 (N_39534,N_39300,N_39331);
or U39535 (N_39535,N_39473,N_39343);
or U39536 (N_39536,N_39282,N_39259);
nor U39537 (N_39537,N_39477,N_39260);
nor U39538 (N_39538,N_39288,N_39379);
nand U39539 (N_39539,N_39378,N_39336);
and U39540 (N_39540,N_39442,N_39278);
xor U39541 (N_39541,N_39471,N_39347);
or U39542 (N_39542,N_39280,N_39397);
nand U39543 (N_39543,N_39455,N_39434);
or U39544 (N_39544,N_39443,N_39322);
nand U39545 (N_39545,N_39250,N_39463);
nor U39546 (N_39546,N_39346,N_39467);
xor U39547 (N_39547,N_39393,N_39252);
or U39548 (N_39548,N_39413,N_39362);
and U39549 (N_39549,N_39441,N_39489);
and U39550 (N_39550,N_39273,N_39319);
xnor U39551 (N_39551,N_39428,N_39432);
and U39552 (N_39552,N_39329,N_39293);
xor U39553 (N_39553,N_39256,N_39404);
nor U39554 (N_39554,N_39394,N_39487);
xnor U39555 (N_39555,N_39277,N_39310);
xor U39556 (N_39556,N_39299,N_39265);
nand U39557 (N_39557,N_39399,N_39342);
nand U39558 (N_39558,N_39358,N_39408);
or U39559 (N_39559,N_39418,N_39426);
nand U39560 (N_39560,N_39440,N_39423);
or U39561 (N_39561,N_39284,N_39353);
nand U39562 (N_39562,N_39359,N_39495);
and U39563 (N_39563,N_39453,N_39365);
xnor U39564 (N_39564,N_39381,N_39412);
nand U39565 (N_39565,N_39482,N_39334);
xnor U39566 (N_39566,N_39344,N_39429);
nor U39567 (N_39567,N_39444,N_39366);
and U39568 (N_39568,N_39389,N_39433);
or U39569 (N_39569,N_39382,N_39255);
nand U39570 (N_39570,N_39335,N_39301);
xnor U39571 (N_39571,N_39414,N_39330);
or U39572 (N_39572,N_39313,N_39281);
or U39573 (N_39573,N_39390,N_39437);
and U39574 (N_39574,N_39261,N_39360);
and U39575 (N_39575,N_39430,N_39287);
xnor U39576 (N_39576,N_39385,N_39395);
and U39577 (N_39577,N_39445,N_39304);
nor U39578 (N_39578,N_39371,N_39294);
xor U39579 (N_39579,N_39354,N_39459);
and U39580 (N_39580,N_39364,N_39391);
nand U39581 (N_39581,N_39460,N_39472);
nor U39582 (N_39582,N_39348,N_39387);
nor U39583 (N_39583,N_39295,N_39465);
nor U39584 (N_39584,N_39388,N_39392);
or U39585 (N_39585,N_39367,N_39318);
or U39586 (N_39586,N_39285,N_39286);
nand U39587 (N_39587,N_39403,N_39271);
nor U39588 (N_39588,N_39483,N_39446);
nor U39589 (N_39589,N_39349,N_39323);
xor U39590 (N_39590,N_39456,N_39279);
xor U39591 (N_39591,N_39496,N_39427);
xnor U39592 (N_39592,N_39435,N_39438);
or U39593 (N_39593,N_39480,N_39488);
xor U39594 (N_39594,N_39290,N_39373);
and U39595 (N_39595,N_39291,N_39484);
xnor U39596 (N_39596,N_39372,N_39475);
nor U39597 (N_39597,N_39407,N_39327);
or U39598 (N_39598,N_39417,N_39332);
nand U39599 (N_39599,N_39499,N_39302);
nand U39600 (N_39600,N_39308,N_39339);
or U39601 (N_39601,N_39333,N_39340);
or U39602 (N_39602,N_39491,N_39452);
xor U39603 (N_39603,N_39309,N_39350);
and U39604 (N_39604,N_39431,N_39415);
nand U39605 (N_39605,N_39352,N_39298);
and U39606 (N_39606,N_39374,N_39457);
and U39607 (N_39607,N_39345,N_39264);
or U39608 (N_39608,N_39283,N_39470);
and U39609 (N_39609,N_39312,N_39421);
xor U39610 (N_39610,N_39384,N_39297);
xnor U39611 (N_39611,N_39292,N_39326);
nand U39612 (N_39612,N_39409,N_39411);
nand U39613 (N_39613,N_39296,N_39416);
nor U39614 (N_39614,N_39439,N_39325);
xnor U39615 (N_39615,N_39258,N_39370);
nand U39616 (N_39616,N_39462,N_39356);
nand U39617 (N_39617,N_39485,N_39436);
and U39618 (N_39618,N_39262,N_39461);
nand U39619 (N_39619,N_39268,N_39357);
and U39620 (N_39620,N_39474,N_39493);
nand U39621 (N_39621,N_39272,N_39458);
nor U39622 (N_39622,N_39402,N_39267);
xor U39623 (N_39623,N_39306,N_39481);
or U39624 (N_39624,N_39454,N_39464);
xnor U39625 (N_39625,N_39270,N_39321);
and U39626 (N_39626,N_39287,N_39378);
nor U39627 (N_39627,N_39255,N_39372);
nor U39628 (N_39628,N_39311,N_39381);
nand U39629 (N_39629,N_39329,N_39444);
or U39630 (N_39630,N_39483,N_39416);
and U39631 (N_39631,N_39284,N_39446);
and U39632 (N_39632,N_39384,N_39430);
or U39633 (N_39633,N_39369,N_39407);
nor U39634 (N_39634,N_39388,N_39344);
xor U39635 (N_39635,N_39294,N_39448);
nor U39636 (N_39636,N_39360,N_39398);
or U39637 (N_39637,N_39250,N_39366);
and U39638 (N_39638,N_39410,N_39486);
xor U39639 (N_39639,N_39415,N_39375);
xor U39640 (N_39640,N_39447,N_39362);
nand U39641 (N_39641,N_39307,N_39283);
or U39642 (N_39642,N_39259,N_39351);
nor U39643 (N_39643,N_39290,N_39417);
nand U39644 (N_39644,N_39483,N_39362);
or U39645 (N_39645,N_39480,N_39492);
and U39646 (N_39646,N_39261,N_39263);
or U39647 (N_39647,N_39392,N_39370);
nand U39648 (N_39648,N_39286,N_39479);
and U39649 (N_39649,N_39437,N_39404);
or U39650 (N_39650,N_39393,N_39477);
xor U39651 (N_39651,N_39444,N_39499);
xnor U39652 (N_39652,N_39259,N_39421);
nand U39653 (N_39653,N_39431,N_39499);
xnor U39654 (N_39654,N_39334,N_39441);
xor U39655 (N_39655,N_39348,N_39279);
and U39656 (N_39656,N_39296,N_39482);
nor U39657 (N_39657,N_39304,N_39365);
and U39658 (N_39658,N_39269,N_39287);
nor U39659 (N_39659,N_39451,N_39431);
and U39660 (N_39660,N_39364,N_39410);
nor U39661 (N_39661,N_39253,N_39338);
xnor U39662 (N_39662,N_39359,N_39287);
nand U39663 (N_39663,N_39430,N_39398);
nor U39664 (N_39664,N_39346,N_39320);
and U39665 (N_39665,N_39428,N_39426);
nand U39666 (N_39666,N_39356,N_39336);
nand U39667 (N_39667,N_39364,N_39303);
xor U39668 (N_39668,N_39371,N_39491);
and U39669 (N_39669,N_39375,N_39385);
and U39670 (N_39670,N_39387,N_39362);
nand U39671 (N_39671,N_39359,N_39346);
and U39672 (N_39672,N_39431,N_39444);
and U39673 (N_39673,N_39283,N_39392);
xnor U39674 (N_39674,N_39357,N_39406);
or U39675 (N_39675,N_39255,N_39465);
nor U39676 (N_39676,N_39471,N_39318);
nor U39677 (N_39677,N_39335,N_39313);
or U39678 (N_39678,N_39398,N_39289);
and U39679 (N_39679,N_39340,N_39443);
and U39680 (N_39680,N_39415,N_39433);
nand U39681 (N_39681,N_39374,N_39479);
and U39682 (N_39682,N_39471,N_39285);
xor U39683 (N_39683,N_39357,N_39400);
and U39684 (N_39684,N_39267,N_39440);
and U39685 (N_39685,N_39499,N_39350);
xor U39686 (N_39686,N_39315,N_39494);
xor U39687 (N_39687,N_39367,N_39437);
xnor U39688 (N_39688,N_39336,N_39412);
xnor U39689 (N_39689,N_39354,N_39294);
and U39690 (N_39690,N_39365,N_39483);
or U39691 (N_39691,N_39409,N_39436);
nor U39692 (N_39692,N_39314,N_39344);
nand U39693 (N_39693,N_39339,N_39338);
and U39694 (N_39694,N_39423,N_39419);
xnor U39695 (N_39695,N_39440,N_39332);
and U39696 (N_39696,N_39390,N_39395);
and U39697 (N_39697,N_39342,N_39370);
and U39698 (N_39698,N_39457,N_39387);
and U39699 (N_39699,N_39474,N_39321);
nand U39700 (N_39700,N_39397,N_39325);
and U39701 (N_39701,N_39401,N_39383);
xor U39702 (N_39702,N_39272,N_39363);
nor U39703 (N_39703,N_39381,N_39498);
nor U39704 (N_39704,N_39359,N_39264);
and U39705 (N_39705,N_39333,N_39312);
nor U39706 (N_39706,N_39273,N_39460);
nor U39707 (N_39707,N_39300,N_39272);
nor U39708 (N_39708,N_39445,N_39428);
or U39709 (N_39709,N_39396,N_39305);
xnor U39710 (N_39710,N_39377,N_39484);
and U39711 (N_39711,N_39371,N_39287);
nor U39712 (N_39712,N_39312,N_39271);
nor U39713 (N_39713,N_39394,N_39473);
nand U39714 (N_39714,N_39350,N_39312);
nand U39715 (N_39715,N_39373,N_39417);
nor U39716 (N_39716,N_39456,N_39296);
nor U39717 (N_39717,N_39285,N_39347);
nor U39718 (N_39718,N_39295,N_39452);
or U39719 (N_39719,N_39449,N_39418);
and U39720 (N_39720,N_39364,N_39354);
xnor U39721 (N_39721,N_39414,N_39267);
and U39722 (N_39722,N_39312,N_39456);
xnor U39723 (N_39723,N_39443,N_39329);
nor U39724 (N_39724,N_39347,N_39410);
nand U39725 (N_39725,N_39442,N_39326);
nor U39726 (N_39726,N_39311,N_39297);
nand U39727 (N_39727,N_39291,N_39481);
and U39728 (N_39728,N_39404,N_39278);
or U39729 (N_39729,N_39304,N_39356);
nand U39730 (N_39730,N_39261,N_39269);
nor U39731 (N_39731,N_39431,N_39335);
or U39732 (N_39732,N_39438,N_39479);
and U39733 (N_39733,N_39496,N_39482);
and U39734 (N_39734,N_39455,N_39269);
nand U39735 (N_39735,N_39491,N_39442);
nand U39736 (N_39736,N_39354,N_39440);
xor U39737 (N_39737,N_39432,N_39474);
nand U39738 (N_39738,N_39265,N_39397);
nand U39739 (N_39739,N_39367,N_39294);
nand U39740 (N_39740,N_39466,N_39404);
xor U39741 (N_39741,N_39408,N_39319);
xor U39742 (N_39742,N_39287,N_39328);
xnor U39743 (N_39743,N_39448,N_39342);
nand U39744 (N_39744,N_39308,N_39463);
or U39745 (N_39745,N_39254,N_39454);
xnor U39746 (N_39746,N_39433,N_39258);
nor U39747 (N_39747,N_39486,N_39404);
nand U39748 (N_39748,N_39253,N_39313);
nand U39749 (N_39749,N_39459,N_39495);
and U39750 (N_39750,N_39578,N_39719);
and U39751 (N_39751,N_39540,N_39530);
nand U39752 (N_39752,N_39640,N_39724);
or U39753 (N_39753,N_39589,N_39737);
nor U39754 (N_39754,N_39745,N_39703);
xor U39755 (N_39755,N_39594,N_39707);
and U39756 (N_39756,N_39646,N_39639);
nor U39757 (N_39757,N_39579,N_39522);
or U39758 (N_39758,N_39658,N_39688);
nand U39759 (N_39759,N_39531,N_39544);
xnor U39760 (N_39760,N_39571,N_39588);
or U39761 (N_39761,N_39702,N_39536);
nor U39762 (N_39762,N_39603,N_39717);
nor U39763 (N_39763,N_39558,N_39657);
xnor U39764 (N_39764,N_39636,N_39504);
or U39765 (N_39765,N_39666,N_39701);
and U39766 (N_39766,N_39642,N_39650);
and U39767 (N_39767,N_39574,N_39532);
xnor U39768 (N_39768,N_39534,N_39700);
and U39769 (N_39769,N_39705,N_39549);
or U39770 (N_39770,N_39747,N_39721);
and U39771 (N_39771,N_39723,N_39545);
and U39772 (N_39772,N_39572,N_39541);
and U39773 (N_39773,N_39628,N_39718);
nor U39774 (N_39774,N_39546,N_39749);
or U39775 (N_39775,N_39599,N_39525);
nand U39776 (N_39776,N_39601,N_39733);
xnor U39777 (N_39777,N_39606,N_39735);
and U39778 (N_39778,N_39738,N_39561);
and U39779 (N_39779,N_39643,N_39526);
nand U39780 (N_39780,N_39533,N_39664);
or U39781 (N_39781,N_39654,N_39568);
and U39782 (N_39782,N_39740,N_39648);
nor U39783 (N_39783,N_39722,N_39619);
and U39784 (N_39784,N_39593,N_39629);
and U39785 (N_39785,N_39617,N_39612);
or U39786 (N_39786,N_39502,N_39644);
and U39787 (N_39787,N_39684,N_39668);
nand U39788 (N_39788,N_39653,N_39509);
nor U39789 (N_39789,N_39590,N_39624);
xnor U39790 (N_39790,N_39575,N_39596);
or U39791 (N_39791,N_39667,N_39686);
xor U39792 (N_39792,N_39520,N_39560);
xnor U39793 (N_39793,N_39517,N_39535);
nor U39794 (N_39794,N_39656,N_39672);
xor U39795 (N_39795,N_39548,N_39630);
and U39796 (N_39796,N_39676,N_39725);
or U39797 (N_39797,N_39713,N_39675);
or U39798 (N_39798,N_39584,N_39691);
xnor U39799 (N_39799,N_39655,N_39739);
or U39800 (N_39800,N_39746,N_39623);
and U39801 (N_39801,N_39716,N_39573);
and U39802 (N_39802,N_39663,N_39690);
or U39803 (N_39803,N_39613,N_39547);
or U39804 (N_39804,N_39741,N_39711);
nor U39805 (N_39805,N_39508,N_39687);
nand U39806 (N_39806,N_39678,N_39500);
xnor U39807 (N_39807,N_39567,N_39514);
nand U39808 (N_39808,N_39627,N_39528);
xor U39809 (N_39809,N_39591,N_39555);
and U39810 (N_39810,N_39742,N_39734);
nand U39811 (N_39811,N_39556,N_39564);
xnor U39812 (N_39812,N_39682,N_39679);
xor U39813 (N_39813,N_39622,N_39685);
and U39814 (N_39814,N_39602,N_39507);
and U39815 (N_39815,N_39552,N_39595);
nor U39816 (N_39816,N_39582,N_39566);
or U39817 (N_39817,N_39683,N_39538);
nand U39818 (N_39818,N_39677,N_39600);
and U39819 (N_39819,N_39694,N_39581);
or U39820 (N_39820,N_39576,N_39647);
nor U39821 (N_39821,N_39543,N_39516);
or U39822 (N_39822,N_39693,N_39637);
nand U39823 (N_39823,N_39689,N_39704);
nand U39824 (N_39824,N_39583,N_39597);
nor U39825 (N_39825,N_39661,N_39699);
nand U39826 (N_39826,N_39651,N_39681);
nand U39827 (N_39827,N_39598,N_39563);
or U39828 (N_39828,N_39550,N_39732);
nor U39829 (N_39829,N_39569,N_39551);
nor U39830 (N_39830,N_39673,N_39510);
or U39831 (N_39831,N_39662,N_39539);
or U39832 (N_39832,N_39634,N_39720);
and U39833 (N_39833,N_39632,N_39665);
xnor U39834 (N_39834,N_39585,N_39503);
and U39835 (N_39835,N_39743,N_39680);
or U39836 (N_39836,N_39641,N_39635);
and U39837 (N_39837,N_39529,N_39674);
nor U39838 (N_39838,N_39744,N_39626);
xor U39839 (N_39839,N_39715,N_39638);
nor U39840 (N_39840,N_39748,N_39727);
nor U39841 (N_39841,N_39607,N_39570);
nor U39842 (N_39842,N_39586,N_39580);
nand U39843 (N_39843,N_39706,N_39587);
or U39844 (N_39844,N_39542,N_39515);
or U39845 (N_39845,N_39671,N_39537);
nor U39846 (N_39846,N_39604,N_39554);
or U39847 (N_39847,N_39649,N_39519);
xor U39848 (N_39848,N_39731,N_39660);
and U39849 (N_39849,N_39736,N_39559);
nor U39850 (N_39850,N_39695,N_39692);
nand U39851 (N_39851,N_39506,N_39730);
nand U39852 (N_39852,N_39527,N_39728);
nand U39853 (N_39853,N_39512,N_39611);
or U39854 (N_39854,N_39610,N_39631);
nand U39855 (N_39855,N_39505,N_39621);
or U39856 (N_39856,N_39501,N_39645);
and U39857 (N_39857,N_39696,N_39616);
xnor U39858 (N_39858,N_39523,N_39709);
nor U39859 (N_39859,N_39670,N_39513);
and U39860 (N_39860,N_39710,N_39614);
nor U39861 (N_39861,N_39708,N_39669);
or U39862 (N_39862,N_39553,N_39608);
nor U39863 (N_39863,N_39615,N_39562);
and U39864 (N_39864,N_39518,N_39577);
nor U39865 (N_39865,N_39511,N_39659);
or U39866 (N_39866,N_39618,N_39609);
xnor U39867 (N_39867,N_39605,N_39524);
nor U39868 (N_39868,N_39565,N_39712);
nand U39869 (N_39869,N_39697,N_39652);
and U39870 (N_39870,N_39625,N_39714);
xor U39871 (N_39871,N_39729,N_39592);
or U39872 (N_39872,N_39726,N_39521);
nand U39873 (N_39873,N_39620,N_39557);
or U39874 (N_39874,N_39633,N_39698);
nor U39875 (N_39875,N_39716,N_39597);
nor U39876 (N_39876,N_39662,N_39745);
and U39877 (N_39877,N_39739,N_39646);
or U39878 (N_39878,N_39538,N_39586);
nand U39879 (N_39879,N_39603,N_39508);
nor U39880 (N_39880,N_39500,N_39508);
nand U39881 (N_39881,N_39597,N_39677);
xnor U39882 (N_39882,N_39625,N_39727);
and U39883 (N_39883,N_39583,N_39603);
nand U39884 (N_39884,N_39678,N_39699);
or U39885 (N_39885,N_39575,N_39595);
xnor U39886 (N_39886,N_39553,N_39671);
nor U39887 (N_39887,N_39578,N_39548);
or U39888 (N_39888,N_39687,N_39748);
and U39889 (N_39889,N_39637,N_39568);
xor U39890 (N_39890,N_39718,N_39674);
and U39891 (N_39891,N_39681,N_39641);
and U39892 (N_39892,N_39607,N_39552);
or U39893 (N_39893,N_39563,N_39601);
and U39894 (N_39894,N_39695,N_39702);
xor U39895 (N_39895,N_39640,N_39725);
xnor U39896 (N_39896,N_39628,N_39594);
xor U39897 (N_39897,N_39580,N_39504);
and U39898 (N_39898,N_39684,N_39600);
nor U39899 (N_39899,N_39582,N_39698);
nand U39900 (N_39900,N_39525,N_39699);
and U39901 (N_39901,N_39599,N_39745);
xor U39902 (N_39902,N_39631,N_39704);
or U39903 (N_39903,N_39535,N_39650);
nand U39904 (N_39904,N_39714,N_39613);
nand U39905 (N_39905,N_39512,N_39714);
nand U39906 (N_39906,N_39652,N_39639);
xnor U39907 (N_39907,N_39747,N_39596);
or U39908 (N_39908,N_39745,N_39543);
xnor U39909 (N_39909,N_39547,N_39687);
nor U39910 (N_39910,N_39682,N_39548);
nand U39911 (N_39911,N_39536,N_39562);
nor U39912 (N_39912,N_39708,N_39686);
nand U39913 (N_39913,N_39615,N_39581);
nor U39914 (N_39914,N_39555,N_39554);
nor U39915 (N_39915,N_39743,N_39655);
nand U39916 (N_39916,N_39555,N_39722);
and U39917 (N_39917,N_39509,N_39500);
nor U39918 (N_39918,N_39746,N_39530);
nor U39919 (N_39919,N_39739,N_39711);
nor U39920 (N_39920,N_39516,N_39705);
and U39921 (N_39921,N_39721,N_39671);
xnor U39922 (N_39922,N_39660,N_39738);
xnor U39923 (N_39923,N_39509,N_39602);
and U39924 (N_39924,N_39718,N_39699);
xor U39925 (N_39925,N_39555,N_39699);
nor U39926 (N_39926,N_39736,N_39535);
nor U39927 (N_39927,N_39530,N_39733);
or U39928 (N_39928,N_39501,N_39544);
or U39929 (N_39929,N_39606,N_39529);
nand U39930 (N_39930,N_39545,N_39636);
and U39931 (N_39931,N_39682,N_39553);
nand U39932 (N_39932,N_39536,N_39664);
and U39933 (N_39933,N_39626,N_39530);
nand U39934 (N_39934,N_39546,N_39706);
and U39935 (N_39935,N_39547,N_39742);
and U39936 (N_39936,N_39689,N_39608);
nand U39937 (N_39937,N_39565,N_39704);
nor U39938 (N_39938,N_39669,N_39664);
and U39939 (N_39939,N_39661,N_39729);
nor U39940 (N_39940,N_39735,N_39688);
nand U39941 (N_39941,N_39588,N_39523);
nor U39942 (N_39942,N_39720,N_39737);
or U39943 (N_39943,N_39508,N_39618);
nor U39944 (N_39944,N_39533,N_39697);
nor U39945 (N_39945,N_39587,N_39583);
nand U39946 (N_39946,N_39715,N_39543);
nor U39947 (N_39947,N_39717,N_39605);
nand U39948 (N_39948,N_39686,N_39596);
nor U39949 (N_39949,N_39537,N_39563);
or U39950 (N_39950,N_39517,N_39740);
and U39951 (N_39951,N_39713,N_39638);
and U39952 (N_39952,N_39643,N_39527);
or U39953 (N_39953,N_39583,N_39614);
nand U39954 (N_39954,N_39612,N_39736);
nand U39955 (N_39955,N_39515,N_39713);
or U39956 (N_39956,N_39608,N_39636);
xor U39957 (N_39957,N_39514,N_39668);
or U39958 (N_39958,N_39725,N_39570);
or U39959 (N_39959,N_39555,N_39706);
nor U39960 (N_39960,N_39633,N_39637);
xor U39961 (N_39961,N_39645,N_39566);
nor U39962 (N_39962,N_39516,N_39696);
or U39963 (N_39963,N_39508,N_39528);
nor U39964 (N_39964,N_39638,N_39504);
nor U39965 (N_39965,N_39669,N_39633);
nand U39966 (N_39966,N_39741,N_39583);
or U39967 (N_39967,N_39608,N_39598);
nor U39968 (N_39968,N_39693,N_39692);
or U39969 (N_39969,N_39658,N_39656);
or U39970 (N_39970,N_39528,N_39622);
nor U39971 (N_39971,N_39698,N_39554);
xnor U39972 (N_39972,N_39563,N_39646);
or U39973 (N_39973,N_39743,N_39660);
nor U39974 (N_39974,N_39540,N_39605);
nor U39975 (N_39975,N_39548,N_39681);
nor U39976 (N_39976,N_39512,N_39563);
or U39977 (N_39977,N_39538,N_39743);
nand U39978 (N_39978,N_39742,N_39602);
nor U39979 (N_39979,N_39537,N_39595);
and U39980 (N_39980,N_39713,N_39731);
xnor U39981 (N_39981,N_39692,N_39746);
xnor U39982 (N_39982,N_39513,N_39702);
nor U39983 (N_39983,N_39572,N_39612);
and U39984 (N_39984,N_39649,N_39678);
and U39985 (N_39985,N_39610,N_39552);
or U39986 (N_39986,N_39546,N_39525);
or U39987 (N_39987,N_39535,N_39709);
nand U39988 (N_39988,N_39529,N_39636);
nand U39989 (N_39989,N_39627,N_39634);
and U39990 (N_39990,N_39665,N_39630);
and U39991 (N_39991,N_39620,N_39731);
or U39992 (N_39992,N_39572,N_39705);
nand U39993 (N_39993,N_39688,N_39631);
or U39994 (N_39994,N_39724,N_39654);
and U39995 (N_39995,N_39634,N_39571);
nor U39996 (N_39996,N_39505,N_39696);
nor U39997 (N_39997,N_39616,N_39559);
nand U39998 (N_39998,N_39744,N_39734);
nand U39999 (N_39999,N_39694,N_39510);
nand U40000 (N_40000,N_39782,N_39815);
or U40001 (N_40001,N_39963,N_39813);
nor U40002 (N_40002,N_39766,N_39923);
nand U40003 (N_40003,N_39860,N_39854);
and U40004 (N_40004,N_39855,N_39762);
nand U40005 (N_40005,N_39957,N_39886);
xor U40006 (N_40006,N_39806,N_39992);
nor U40007 (N_40007,N_39770,N_39793);
xor U40008 (N_40008,N_39752,N_39897);
and U40009 (N_40009,N_39881,N_39982);
and U40010 (N_40010,N_39929,N_39787);
or U40011 (N_40011,N_39814,N_39755);
nor U40012 (N_40012,N_39911,N_39900);
or U40013 (N_40013,N_39800,N_39893);
xor U40014 (N_40014,N_39899,N_39954);
and U40015 (N_40015,N_39940,N_39934);
nor U40016 (N_40016,N_39767,N_39820);
nor U40017 (N_40017,N_39908,N_39827);
xor U40018 (N_40018,N_39865,N_39780);
or U40019 (N_40019,N_39887,N_39965);
nand U40020 (N_40020,N_39987,N_39856);
nor U40021 (N_40021,N_39816,N_39792);
nor U40022 (N_40022,N_39933,N_39975);
and U40023 (N_40023,N_39844,N_39794);
nor U40024 (N_40024,N_39817,N_39990);
nand U40025 (N_40025,N_39882,N_39790);
and U40026 (N_40026,N_39909,N_39830);
xnor U40027 (N_40027,N_39907,N_39935);
xnor U40028 (N_40028,N_39845,N_39759);
nor U40029 (N_40029,N_39979,N_39952);
nor U40030 (N_40030,N_39843,N_39864);
nand U40031 (N_40031,N_39809,N_39930);
and U40032 (N_40032,N_39981,N_39924);
xor U40033 (N_40033,N_39773,N_39905);
or U40034 (N_40034,N_39758,N_39871);
xnor U40035 (N_40035,N_39776,N_39959);
xor U40036 (N_40036,N_39869,N_39873);
and U40037 (N_40037,N_39898,N_39995);
and U40038 (N_40038,N_39999,N_39892);
and U40039 (N_40039,N_39837,N_39942);
and U40040 (N_40040,N_39821,N_39764);
and U40041 (N_40041,N_39789,N_39956);
and U40042 (N_40042,N_39788,N_39926);
xor U40043 (N_40043,N_39966,N_39944);
or U40044 (N_40044,N_39941,N_39996);
nand U40045 (N_40045,N_39802,N_39832);
nand U40046 (N_40046,N_39947,N_39994);
or U40047 (N_40047,N_39874,N_39868);
xor U40048 (N_40048,N_39939,N_39936);
xnor U40049 (N_40049,N_39819,N_39977);
nand U40050 (N_40050,N_39901,N_39812);
nand U40051 (N_40051,N_39914,N_39804);
or U40052 (N_40052,N_39807,N_39991);
nand U40053 (N_40053,N_39839,N_39961);
nor U40054 (N_40054,N_39904,N_39811);
and U40055 (N_40055,N_39875,N_39796);
or U40056 (N_40056,N_39958,N_39912);
nor U40057 (N_40057,N_39877,N_39921);
nor U40058 (N_40058,N_39920,N_39797);
nor U40059 (N_40059,N_39879,N_39862);
xnor U40060 (N_40060,N_39784,N_39867);
and U40061 (N_40061,N_39988,N_39880);
and U40062 (N_40062,N_39943,N_39998);
nor U40063 (N_40063,N_39910,N_39824);
and U40064 (N_40064,N_39876,N_39989);
nand U40065 (N_40065,N_39883,N_39857);
or U40066 (N_40066,N_39971,N_39949);
nor U40067 (N_40067,N_39919,N_39891);
or U40068 (N_40068,N_39783,N_39772);
or U40069 (N_40069,N_39872,N_39795);
nor U40070 (N_40070,N_39848,N_39834);
or U40071 (N_40071,N_39851,N_39931);
and U40072 (N_40072,N_39937,N_39853);
nand U40073 (N_40073,N_39791,N_39778);
or U40074 (N_40074,N_39774,N_39779);
or U40075 (N_40075,N_39889,N_39754);
nand U40076 (N_40076,N_39927,N_39970);
or U40077 (N_40077,N_39974,N_39849);
or U40078 (N_40078,N_39928,N_39753);
or U40079 (N_40079,N_39948,N_39946);
and U40080 (N_40080,N_39808,N_39895);
or U40081 (N_40081,N_39953,N_39925);
and U40082 (N_40082,N_39976,N_39969);
nor U40083 (N_40083,N_39801,N_39859);
nand U40084 (N_40084,N_39922,N_39818);
or U40085 (N_40085,N_39822,N_39968);
and U40086 (N_40086,N_39960,N_39913);
nor U40087 (N_40087,N_39918,N_39978);
nor U40088 (N_40088,N_39842,N_39785);
and U40089 (N_40089,N_39993,N_39878);
or U40090 (N_40090,N_39866,N_39805);
xnor U40091 (N_40091,N_39841,N_39983);
nand U40092 (N_40092,N_39964,N_39972);
nor U40093 (N_40093,N_39831,N_39984);
or U40094 (N_40094,N_39771,N_39894);
nor U40095 (N_40095,N_39786,N_39756);
or U40096 (N_40096,N_39829,N_39769);
and U40097 (N_40097,N_39915,N_39836);
nor U40098 (N_40098,N_39938,N_39823);
nand U40099 (N_40099,N_39850,N_39828);
nor U40100 (N_40100,N_39750,N_39945);
nor U40101 (N_40101,N_39825,N_39775);
nand U40102 (N_40102,N_39798,N_39847);
and U40103 (N_40103,N_39835,N_39858);
and U40104 (N_40104,N_39751,N_39799);
and U40105 (N_40105,N_39863,N_39917);
and U40106 (N_40106,N_39962,N_39951);
xnor U40107 (N_40107,N_39763,N_39840);
and U40108 (N_40108,N_39838,N_39760);
nor U40109 (N_40109,N_39803,N_39826);
and U40110 (N_40110,N_39903,N_39870);
or U40111 (N_40111,N_39852,N_39896);
xnor U40112 (N_40112,N_39985,N_39757);
nand U40113 (N_40113,N_39781,N_39980);
nand U40114 (N_40114,N_39932,N_39997);
xnor U40115 (N_40115,N_39846,N_39861);
and U40116 (N_40116,N_39768,N_39967);
and U40117 (N_40117,N_39890,N_39884);
or U40118 (N_40118,N_39761,N_39906);
nand U40119 (N_40119,N_39765,N_39833);
xor U40120 (N_40120,N_39986,N_39777);
and U40121 (N_40121,N_39916,N_39888);
xnor U40122 (N_40122,N_39950,N_39902);
xnor U40123 (N_40123,N_39810,N_39955);
and U40124 (N_40124,N_39973,N_39885);
nand U40125 (N_40125,N_39870,N_39893);
xnor U40126 (N_40126,N_39790,N_39848);
and U40127 (N_40127,N_39863,N_39889);
nor U40128 (N_40128,N_39750,N_39826);
and U40129 (N_40129,N_39905,N_39782);
xnor U40130 (N_40130,N_39890,N_39765);
or U40131 (N_40131,N_39889,N_39990);
nor U40132 (N_40132,N_39872,N_39959);
xnor U40133 (N_40133,N_39888,N_39977);
and U40134 (N_40134,N_39896,N_39816);
nor U40135 (N_40135,N_39967,N_39887);
nor U40136 (N_40136,N_39868,N_39788);
or U40137 (N_40137,N_39783,N_39834);
or U40138 (N_40138,N_39889,N_39877);
and U40139 (N_40139,N_39933,N_39854);
nor U40140 (N_40140,N_39796,N_39930);
and U40141 (N_40141,N_39858,N_39968);
nand U40142 (N_40142,N_39989,N_39918);
xnor U40143 (N_40143,N_39913,N_39959);
xnor U40144 (N_40144,N_39850,N_39936);
xor U40145 (N_40145,N_39866,N_39953);
or U40146 (N_40146,N_39820,N_39995);
xor U40147 (N_40147,N_39769,N_39764);
xnor U40148 (N_40148,N_39844,N_39928);
or U40149 (N_40149,N_39916,N_39811);
or U40150 (N_40150,N_39773,N_39856);
and U40151 (N_40151,N_39894,N_39799);
nand U40152 (N_40152,N_39858,N_39788);
and U40153 (N_40153,N_39925,N_39986);
or U40154 (N_40154,N_39902,N_39829);
xnor U40155 (N_40155,N_39988,N_39979);
nand U40156 (N_40156,N_39906,N_39943);
or U40157 (N_40157,N_39905,N_39864);
nor U40158 (N_40158,N_39900,N_39923);
nand U40159 (N_40159,N_39941,N_39903);
nor U40160 (N_40160,N_39929,N_39896);
or U40161 (N_40161,N_39784,N_39992);
nand U40162 (N_40162,N_39962,N_39847);
nor U40163 (N_40163,N_39853,N_39945);
nor U40164 (N_40164,N_39959,N_39869);
nor U40165 (N_40165,N_39984,N_39756);
nand U40166 (N_40166,N_39836,N_39971);
or U40167 (N_40167,N_39817,N_39776);
nand U40168 (N_40168,N_39951,N_39918);
nand U40169 (N_40169,N_39910,N_39864);
or U40170 (N_40170,N_39872,N_39756);
or U40171 (N_40171,N_39845,N_39957);
or U40172 (N_40172,N_39907,N_39894);
and U40173 (N_40173,N_39821,N_39880);
nand U40174 (N_40174,N_39784,N_39801);
nand U40175 (N_40175,N_39756,N_39912);
xnor U40176 (N_40176,N_39953,N_39948);
nor U40177 (N_40177,N_39882,N_39772);
or U40178 (N_40178,N_39848,N_39767);
xor U40179 (N_40179,N_39929,N_39967);
nor U40180 (N_40180,N_39922,N_39867);
nand U40181 (N_40181,N_39832,N_39938);
nand U40182 (N_40182,N_39780,N_39938);
nor U40183 (N_40183,N_39889,N_39766);
xor U40184 (N_40184,N_39870,N_39788);
and U40185 (N_40185,N_39790,N_39885);
nand U40186 (N_40186,N_39900,N_39957);
xor U40187 (N_40187,N_39842,N_39792);
nand U40188 (N_40188,N_39793,N_39823);
xnor U40189 (N_40189,N_39757,N_39892);
or U40190 (N_40190,N_39890,N_39920);
nor U40191 (N_40191,N_39952,N_39799);
or U40192 (N_40192,N_39851,N_39771);
and U40193 (N_40193,N_39891,N_39980);
xor U40194 (N_40194,N_39770,N_39939);
or U40195 (N_40195,N_39928,N_39932);
nor U40196 (N_40196,N_39830,N_39764);
or U40197 (N_40197,N_39948,N_39757);
and U40198 (N_40198,N_39941,N_39951);
nand U40199 (N_40199,N_39992,N_39947);
or U40200 (N_40200,N_39874,N_39928);
nand U40201 (N_40201,N_39897,N_39852);
and U40202 (N_40202,N_39890,N_39752);
nor U40203 (N_40203,N_39840,N_39769);
or U40204 (N_40204,N_39849,N_39794);
xnor U40205 (N_40205,N_39921,N_39913);
and U40206 (N_40206,N_39750,N_39806);
nand U40207 (N_40207,N_39847,N_39876);
and U40208 (N_40208,N_39817,N_39986);
xor U40209 (N_40209,N_39853,N_39926);
nor U40210 (N_40210,N_39954,N_39965);
nand U40211 (N_40211,N_39817,N_39947);
nor U40212 (N_40212,N_39973,N_39992);
nor U40213 (N_40213,N_39887,N_39962);
nor U40214 (N_40214,N_39875,N_39926);
nor U40215 (N_40215,N_39814,N_39841);
nand U40216 (N_40216,N_39996,N_39821);
or U40217 (N_40217,N_39970,N_39796);
or U40218 (N_40218,N_39959,N_39987);
nand U40219 (N_40219,N_39759,N_39828);
and U40220 (N_40220,N_39764,N_39868);
nand U40221 (N_40221,N_39776,N_39862);
xnor U40222 (N_40222,N_39766,N_39950);
nor U40223 (N_40223,N_39752,N_39922);
nand U40224 (N_40224,N_39879,N_39926);
nor U40225 (N_40225,N_39769,N_39947);
xnor U40226 (N_40226,N_39760,N_39862);
or U40227 (N_40227,N_39841,N_39807);
nor U40228 (N_40228,N_39983,N_39845);
and U40229 (N_40229,N_39755,N_39897);
and U40230 (N_40230,N_39868,N_39754);
nor U40231 (N_40231,N_39988,N_39845);
nand U40232 (N_40232,N_39796,N_39954);
nor U40233 (N_40233,N_39808,N_39962);
or U40234 (N_40234,N_39840,N_39750);
nand U40235 (N_40235,N_39902,N_39839);
or U40236 (N_40236,N_39904,N_39992);
nand U40237 (N_40237,N_39969,N_39782);
xor U40238 (N_40238,N_39787,N_39978);
and U40239 (N_40239,N_39808,N_39876);
or U40240 (N_40240,N_39956,N_39836);
xor U40241 (N_40241,N_39824,N_39924);
or U40242 (N_40242,N_39838,N_39909);
and U40243 (N_40243,N_39903,N_39897);
nand U40244 (N_40244,N_39812,N_39979);
nor U40245 (N_40245,N_39959,N_39860);
and U40246 (N_40246,N_39863,N_39817);
nor U40247 (N_40247,N_39804,N_39846);
and U40248 (N_40248,N_39910,N_39888);
or U40249 (N_40249,N_39826,N_39875);
xor U40250 (N_40250,N_40151,N_40211);
nand U40251 (N_40251,N_40246,N_40011);
nand U40252 (N_40252,N_40181,N_40120);
nor U40253 (N_40253,N_40056,N_40185);
xor U40254 (N_40254,N_40145,N_40160);
and U40255 (N_40255,N_40022,N_40131);
nor U40256 (N_40256,N_40086,N_40112);
or U40257 (N_40257,N_40183,N_40029);
nand U40258 (N_40258,N_40105,N_40113);
nand U40259 (N_40259,N_40073,N_40219);
or U40260 (N_40260,N_40161,N_40241);
and U40261 (N_40261,N_40116,N_40005);
nor U40262 (N_40262,N_40212,N_40249);
nor U40263 (N_40263,N_40013,N_40202);
nand U40264 (N_40264,N_40166,N_40052);
or U40265 (N_40265,N_40077,N_40053);
xor U40266 (N_40266,N_40067,N_40223);
and U40267 (N_40267,N_40118,N_40242);
or U40268 (N_40268,N_40025,N_40061);
xnor U40269 (N_40269,N_40066,N_40104);
nand U40270 (N_40270,N_40082,N_40179);
nor U40271 (N_40271,N_40169,N_40142);
nor U40272 (N_40272,N_40075,N_40174);
nor U40273 (N_40273,N_40002,N_40156);
or U40274 (N_40274,N_40058,N_40038);
nand U40275 (N_40275,N_40081,N_40159);
or U40276 (N_40276,N_40230,N_40232);
nand U40277 (N_40277,N_40115,N_40057);
or U40278 (N_40278,N_40214,N_40041);
or U40279 (N_40279,N_40088,N_40102);
and U40280 (N_40280,N_40182,N_40243);
and U40281 (N_40281,N_40172,N_40020);
or U40282 (N_40282,N_40195,N_40090);
nor U40283 (N_40283,N_40042,N_40247);
and U40284 (N_40284,N_40039,N_40175);
nand U40285 (N_40285,N_40089,N_40125);
and U40286 (N_40286,N_40111,N_40193);
nor U40287 (N_40287,N_40083,N_40010);
and U40288 (N_40288,N_40107,N_40079);
and U40289 (N_40289,N_40101,N_40017);
nand U40290 (N_40290,N_40206,N_40154);
or U40291 (N_40291,N_40031,N_40098);
and U40292 (N_40292,N_40237,N_40198);
xor U40293 (N_40293,N_40205,N_40244);
nand U40294 (N_40294,N_40229,N_40108);
xor U40295 (N_40295,N_40036,N_40018);
xor U40296 (N_40296,N_40167,N_40070);
or U40297 (N_40297,N_40177,N_40171);
nand U40298 (N_40298,N_40173,N_40149);
nor U40299 (N_40299,N_40140,N_40046);
nor U40300 (N_40300,N_40139,N_40059);
xnor U40301 (N_40301,N_40144,N_40069);
and U40302 (N_40302,N_40204,N_40027);
nand U40303 (N_40303,N_40092,N_40133);
xor U40304 (N_40304,N_40040,N_40095);
nor U40305 (N_40305,N_40076,N_40187);
nor U40306 (N_40306,N_40191,N_40132);
xor U40307 (N_40307,N_40163,N_40049);
and U40308 (N_40308,N_40155,N_40016);
nand U40309 (N_40309,N_40080,N_40138);
xor U40310 (N_40310,N_40033,N_40085);
nand U40311 (N_40311,N_40134,N_40148);
and U40312 (N_40312,N_40128,N_40162);
nand U40313 (N_40313,N_40137,N_40119);
and U40314 (N_40314,N_40186,N_40099);
nand U40315 (N_40315,N_40201,N_40216);
or U40316 (N_40316,N_40045,N_40051);
nor U40317 (N_40317,N_40019,N_40188);
nor U40318 (N_40318,N_40235,N_40153);
nand U40319 (N_40319,N_40117,N_40096);
xor U40320 (N_40320,N_40034,N_40192);
nand U40321 (N_40321,N_40130,N_40184);
and U40322 (N_40322,N_40164,N_40078);
nand U40323 (N_40323,N_40215,N_40122);
or U40324 (N_40324,N_40109,N_40150);
nor U40325 (N_40325,N_40209,N_40103);
nand U40326 (N_40326,N_40063,N_40176);
and U40327 (N_40327,N_40068,N_40165);
xor U40328 (N_40328,N_40030,N_40009);
nand U40329 (N_40329,N_40127,N_40054);
nor U40330 (N_40330,N_40231,N_40129);
and U40331 (N_40331,N_40240,N_40157);
nor U40332 (N_40332,N_40087,N_40071);
and U40333 (N_40333,N_40210,N_40032);
nand U40334 (N_40334,N_40004,N_40222);
or U40335 (N_40335,N_40012,N_40190);
xor U40336 (N_40336,N_40000,N_40218);
or U40337 (N_40337,N_40028,N_40100);
nor U40338 (N_40338,N_40136,N_40084);
xor U40339 (N_40339,N_40094,N_40143);
nor U40340 (N_40340,N_40228,N_40170);
and U40341 (N_40341,N_40245,N_40147);
or U40342 (N_40342,N_40014,N_40008);
nor U40343 (N_40343,N_40225,N_40065);
nand U40344 (N_40344,N_40220,N_40234);
xnor U40345 (N_40345,N_40224,N_40236);
xnor U40346 (N_40346,N_40123,N_40091);
xnor U40347 (N_40347,N_40152,N_40048);
xnor U40348 (N_40348,N_40064,N_40007);
or U40349 (N_40349,N_40178,N_40097);
and U40350 (N_40350,N_40168,N_40248);
nand U40351 (N_40351,N_40203,N_40003);
nand U40352 (N_40352,N_40044,N_40114);
nor U40353 (N_40353,N_40110,N_40026);
xor U40354 (N_40354,N_40238,N_40126);
nor U40355 (N_40355,N_40021,N_40050);
xnor U40356 (N_40356,N_40001,N_40106);
and U40357 (N_40357,N_40074,N_40227);
xnor U40358 (N_40358,N_40146,N_40207);
nand U40359 (N_40359,N_40072,N_40208);
and U40360 (N_40360,N_40217,N_40141);
and U40361 (N_40361,N_40189,N_40043);
or U40362 (N_40362,N_40194,N_40180);
or U40363 (N_40363,N_40055,N_40015);
and U40364 (N_40364,N_40226,N_40062);
or U40365 (N_40365,N_40124,N_40199);
nand U40366 (N_40366,N_40135,N_40197);
nor U40367 (N_40367,N_40037,N_40060);
or U40368 (N_40368,N_40093,N_40047);
nor U40369 (N_40369,N_40024,N_40200);
nand U40370 (N_40370,N_40121,N_40006);
nand U40371 (N_40371,N_40196,N_40023);
nand U40372 (N_40372,N_40233,N_40221);
nand U40373 (N_40373,N_40035,N_40213);
and U40374 (N_40374,N_40158,N_40239);
nor U40375 (N_40375,N_40050,N_40204);
nand U40376 (N_40376,N_40139,N_40157);
or U40377 (N_40377,N_40036,N_40212);
nand U40378 (N_40378,N_40057,N_40042);
or U40379 (N_40379,N_40203,N_40150);
nand U40380 (N_40380,N_40170,N_40154);
or U40381 (N_40381,N_40014,N_40158);
nor U40382 (N_40382,N_40058,N_40163);
nor U40383 (N_40383,N_40139,N_40167);
xor U40384 (N_40384,N_40220,N_40002);
xnor U40385 (N_40385,N_40105,N_40131);
or U40386 (N_40386,N_40047,N_40087);
nor U40387 (N_40387,N_40037,N_40090);
nor U40388 (N_40388,N_40115,N_40068);
nor U40389 (N_40389,N_40082,N_40187);
and U40390 (N_40390,N_40121,N_40133);
xor U40391 (N_40391,N_40207,N_40244);
or U40392 (N_40392,N_40106,N_40090);
nand U40393 (N_40393,N_40232,N_40018);
and U40394 (N_40394,N_40234,N_40209);
and U40395 (N_40395,N_40112,N_40148);
nand U40396 (N_40396,N_40007,N_40146);
and U40397 (N_40397,N_40148,N_40078);
nand U40398 (N_40398,N_40176,N_40234);
nand U40399 (N_40399,N_40168,N_40145);
xor U40400 (N_40400,N_40061,N_40041);
nor U40401 (N_40401,N_40131,N_40000);
or U40402 (N_40402,N_40137,N_40123);
or U40403 (N_40403,N_40063,N_40156);
nor U40404 (N_40404,N_40006,N_40205);
xor U40405 (N_40405,N_40249,N_40007);
xor U40406 (N_40406,N_40021,N_40018);
xnor U40407 (N_40407,N_40178,N_40143);
or U40408 (N_40408,N_40197,N_40103);
nand U40409 (N_40409,N_40175,N_40047);
nand U40410 (N_40410,N_40232,N_40209);
or U40411 (N_40411,N_40233,N_40101);
xor U40412 (N_40412,N_40075,N_40221);
or U40413 (N_40413,N_40127,N_40036);
nor U40414 (N_40414,N_40203,N_40205);
nand U40415 (N_40415,N_40089,N_40131);
and U40416 (N_40416,N_40004,N_40040);
nor U40417 (N_40417,N_40012,N_40206);
nand U40418 (N_40418,N_40136,N_40213);
nand U40419 (N_40419,N_40136,N_40024);
nor U40420 (N_40420,N_40056,N_40142);
nand U40421 (N_40421,N_40127,N_40073);
xnor U40422 (N_40422,N_40146,N_40201);
xnor U40423 (N_40423,N_40187,N_40101);
or U40424 (N_40424,N_40006,N_40164);
nor U40425 (N_40425,N_40098,N_40041);
and U40426 (N_40426,N_40152,N_40070);
nand U40427 (N_40427,N_40183,N_40100);
nand U40428 (N_40428,N_40205,N_40218);
nand U40429 (N_40429,N_40110,N_40167);
and U40430 (N_40430,N_40086,N_40196);
nor U40431 (N_40431,N_40056,N_40014);
xnor U40432 (N_40432,N_40188,N_40169);
xor U40433 (N_40433,N_40139,N_40134);
and U40434 (N_40434,N_40245,N_40082);
xor U40435 (N_40435,N_40129,N_40197);
or U40436 (N_40436,N_40043,N_40244);
nor U40437 (N_40437,N_40180,N_40159);
nor U40438 (N_40438,N_40214,N_40030);
xnor U40439 (N_40439,N_40211,N_40102);
nor U40440 (N_40440,N_40245,N_40039);
xnor U40441 (N_40441,N_40178,N_40009);
nand U40442 (N_40442,N_40098,N_40205);
and U40443 (N_40443,N_40216,N_40071);
xor U40444 (N_40444,N_40015,N_40217);
xnor U40445 (N_40445,N_40114,N_40205);
nor U40446 (N_40446,N_40062,N_40197);
nand U40447 (N_40447,N_40088,N_40074);
nor U40448 (N_40448,N_40119,N_40002);
nor U40449 (N_40449,N_40114,N_40240);
nand U40450 (N_40450,N_40048,N_40228);
or U40451 (N_40451,N_40126,N_40237);
xnor U40452 (N_40452,N_40067,N_40114);
and U40453 (N_40453,N_40167,N_40143);
nor U40454 (N_40454,N_40164,N_40024);
nand U40455 (N_40455,N_40144,N_40143);
nor U40456 (N_40456,N_40224,N_40134);
xnor U40457 (N_40457,N_40077,N_40132);
or U40458 (N_40458,N_40155,N_40061);
nor U40459 (N_40459,N_40013,N_40097);
xor U40460 (N_40460,N_40137,N_40207);
nor U40461 (N_40461,N_40106,N_40065);
xnor U40462 (N_40462,N_40038,N_40233);
or U40463 (N_40463,N_40115,N_40061);
xnor U40464 (N_40464,N_40044,N_40010);
and U40465 (N_40465,N_40219,N_40121);
xnor U40466 (N_40466,N_40245,N_40065);
or U40467 (N_40467,N_40199,N_40052);
xor U40468 (N_40468,N_40128,N_40126);
nor U40469 (N_40469,N_40218,N_40197);
xnor U40470 (N_40470,N_40087,N_40076);
nand U40471 (N_40471,N_40011,N_40249);
nor U40472 (N_40472,N_40168,N_40057);
xnor U40473 (N_40473,N_40063,N_40104);
xor U40474 (N_40474,N_40029,N_40210);
nand U40475 (N_40475,N_40064,N_40045);
nor U40476 (N_40476,N_40119,N_40052);
xnor U40477 (N_40477,N_40187,N_40147);
xnor U40478 (N_40478,N_40127,N_40106);
nand U40479 (N_40479,N_40233,N_40183);
or U40480 (N_40480,N_40189,N_40065);
xor U40481 (N_40481,N_40201,N_40184);
and U40482 (N_40482,N_40052,N_40004);
or U40483 (N_40483,N_40241,N_40126);
nand U40484 (N_40484,N_40232,N_40079);
or U40485 (N_40485,N_40120,N_40183);
or U40486 (N_40486,N_40048,N_40248);
xor U40487 (N_40487,N_40035,N_40144);
or U40488 (N_40488,N_40003,N_40245);
or U40489 (N_40489,N_40224,N_40122);
nor U40490 (N_40490,N_40043,N_40186);
and U40491 (N_40491,N_40199,N_40197);
nand U40492 (N_40492,N_40107,N_40152);
nand U40493 (N_40493,N_40051,N_40244);
or U40494 (N_40494,N_40216,N_40192);
xor U40495 (N_40495,N_40086,N_40065);
or U40496 (N_40496,N_40085,N_40177);
nor U40497 (N_40497,N_40013,N_40016);
nand U40498 (N_40498,N_40078,N_40127);
nand U40499 (N_40499,N_40025,N_40147);
nor U40500 (N_40500,N_40432,N_40421);
and U40501 (N_40501,N_40343,N_40291);
and U40502 (N_40502,N_40358,N_40366);
or U40503 (N_40503,N_40331,N_40373);
or U40504 (N_40504,N_40292,N_40313);
nor U40505 (N_40505,N_40499,N_40319);
and U40506 (N_40506,N_40463,N_40411);
nor U40507 (N_40507,N_40274,N_40272);
and U40508 (N_40508,N_40384,N_40419);
and U40509 (N_40509,N_40307,N_40295);
and U40510 (N_40510,N_40452,N_40412);
nand U40511 (N_40511,N_40333,N_40380);
xnor U40512 (N_40512,N_40265,N_40455);
xnor U40513 (N_40513,N_40271,N_40376);
nand U40514 (N_40514,N_40461,N_40396);
nor U40515 (N_40515,N_40318,N_40270);
xor U40516 (N_40516,N_40392,N_40442);
and U40517 (N_40517,N_40334,N_40298);
xnor U40518 (N_40518,N_40449,N_40390);
and U40519 (N_40519,N_40278,N_40382);
nor U40520 (N_40520,N_40320,N_40394);
xor U40521 (N_40521,N_40266,N_40363);
nand U40522 (N_40522,N_40341,N_40375);
and U40523 (N_40523,N_40325,N_40410);
or U40524 (N_40524,N_40460,N_40342);
nand U40525 (N_40525,N_40494,N_40405);
nand U40526 (N_40526,N_40422,N_40316);
nor U40527 (N_40527,N_40258,N_40389);
or U40528 (N_40528,N_40283,N_40254);
xnor U40529 (N_40529,N_40415,N_40381);
nor U40530 (N_40530,N_40427,N_40487);
or U40531 (N_40531,N_40330,N_40281);
nor U40532 (N_40532,N_40475,N_40468);
nor U40533 (N_40533,N_40482,N_40485);
or U40534 (N_40534,N_40413,N_40273);
and U40535 (N_40535,N_40473,N_40369);
nand U40536 (N_40536,N_40260,N_40399);
nand U40537 (N_40537,N_40267,N_40378);
xor U40538 (N_40538,N_40483,N_40256);
or U40539 (N_40539,N_40275,N_40374);
or U40540 (N_40540,N_40466,N_40430);
xnor U40541 (N_40541,N_40417,N_40329);
nor U40542 (N_40542,N_40255,N_40490);
and U40543 (N_40543,N_40416,N_40403);
nand U40544 (N_40544,N_40350,N_40439);
and U40545 (N_40545,N_40303,N_40336);
nand U40546 (N_40546,N_40454,N_40406);
and U40547 (N_40547,N_40304,N_40289);
nand U40548 (N_40548,N_40491,N_40429);
or U40549 (N_40549,N_40264,N_40301);
and U40550 (N_40550,N_40328,N_40477);
nor U40551 (N_40551,N_40326,N_40359);
xor U40552 (N_40552,N_40495,N_40445);
and U40553 (N_40553,N_40252,N_40493);
or U40554 (N_40554,N_40250,N_40424);
nand U40555 (N_40555,N_40288,N_40352);
nand U40556 (N_40556,N_40367,N_40294);
and U40557 (N_40557,N_40443,N_40268);
or U40558 (N_40558,N_40299,N_40306);
nor U40559 (N_40559,N_40441,N_40437);
xnor U40560 (N_40560,N_40465,N_40492);
and U40561 (N_40561,N_40447,N_40314);
or U40562 (N_40562,N_40279,N_40277);
and U40563 (N_40563,N_40310,N_40261);
or U40564 (N_40564,N_40347,N_40300);
or U40565 (N_40565,N_40311,N_40446);
and U40566 (N_40566,N_40354,N_40425);
and U40567 (N_40567,N_40282,N_40349);
xnor U40568 (N_40568,N_40462,N_40297);
xnor U40569 (N_40569,N_40324,N_40387);
nor U40570 (N_40570,N_40469,N_40420);
nand U40571 (N_40571,N_40386,N_40379);
nor U40572 (N_40572,N_40440,N_40346);
nor U40573 (N_40573,N_40385,N_40315);
nor U40574 (N_40574,N_40404,N_40259);
nor U40575 (N_40575,N_40401,N_40371);
xnor U40576 (N_40576,N_40251,N_40428);
nand U40577 (N_40577,N_40484,N_40340);
nor U40578 (N_40578,N_40489,N_40434);
or U40579 (N_40579,N_40409,N_40360);
and U40580 (N_40580,N_40348,N_40456);
or U40581 (N_40581,N_40305,N_40418);
nor U40582 (N_40582,N_40481,N_40457);
nor U40583 (N_40583,N_40388,N_40312);
nand U40584 (N_40584,N_40276,N_40269);
nand U40585 (N_40585,N_40280,N_40486);
or U40586 (N_40586,N_40414,N_40368);
and U40587 (N_40587,N_40393,N_40471);
or U40588 (N_40588,N_40309,N_40370);
or U40589 (N_40589,N_40391,N_40339);
nor U40590 (N_40590,N_40450,N_40408);
nand U40591 (N_40591,N_40356,N_40436);
or U40592 (N_40592,N_40286,N_40488);
xor U40593 (N_40593,N_40407,N_40361);
and U40594 (N_40594,N_40365,N_40480);
and U40595 (N_40595,N_40497,N_40496);
xnor U40596 (N_40596,N_40476,N_40364);
nor U40597 (N_40597,N_40345,N_40284);
and U40598 (N_40598,N_40435,N_40332);
and U40599 (N_40599,N_40317,N_40453);
nand U40600 (N_40600,N_40262,N_40383);
nor U40601 (N_40601,N_40400,N_40423);
and U40602 (N_40602,N_40478,N_40451);
xnor U40603 (N_40603,N_40335,N_40458);
nand U40604 (N_40604,N_40438,N_40397);
nor U40605 (N_40605,N_40377,N_40431);
xnor U40606 (N_40606,N_40470,N_40327);
nand U40607 (N_40607,N_40293,N_40308);
xor U40608 (N_40608,N_40321,N_40474);
nand U40609 (N_40609,N_40302,N_40287);
nand U40610 (N_40610,N_40444,N_40402);
or U40611 (N_40611,N_40296,N_40337);
nor U40612 (N_40612,N_40498,N_40323);
or U40613 (N_40613,N_40257,N_40433);
nand U40614 (N_40614,N_40322,N_40448);
and U40615 (N_40615,N_40338,N_40467);
nor U40616 (N_40616,N_40355,N_40362);
or U40617 (N_40617,N_40395,N_40357);
nand U40618 (N_40618,N_40263,N_40351);
and U40619 (N_40619,N_40353,N_40459);
and U40620 (N_40620,N_40464,N_40472);
nor U40621 (N_40621,N_40344,N_40398);
xnor U40622 (N_40622,N_40285,N_40290);
nand U40623 (N_40623,N_40372,N_40479);
nor U40624 (N_40624,N_40253,N_40426);
or U40625 (N_40625,N_40255,N_40284);
or U40626 (N_40626,N_40368,N_40281);
nand U40627 (N_40627,N_40367,N_40495);
nor U40628 (N_40628,N_40376,N_40311);
xor U40629 (N_40629,N_40423,N_40344);
and U40630 (N_40630,N_40255,N_40411);
nor U40631 (N_40631,N_40277,N_40497);
and U40632 (N_40632,N_40349,N_40352);
nand U40633 (N_40633,N_40406,N_40296);
and U40634 (N_40634,N_40288,N_40331);
nor U40635 (N_40635,N_40475,N_40314);
and U40636 (N_40636,N_40373,N_40252);
nor U40637 (N_40637,N_40349,N_40367);
xnor U40638 (N_40638,N_40495,N_40259);
and U40639 (N_40639,N_40470,N_40268);
nand U40640 (N_40640,N_40260,N_40443);
xor U40641 (N_40641,N_40468,N_40474);
nor U40642 (N_40642,N_40429,N_40378);
nor U40643 (N_40643,N_40328,N_40456);
nor U40644 (N_40644,N_40406,N_40409);
nand U40645 (N_40645,N_40492,N_40419);
nor U40646 (N_40646,N_40321,N_40363);
and U40647 (N_40647,N_40252,N_40432);
or U40648 (N_40648,N_40467,N_40369);
xor U40649 (N_40649,N_40419,N_40334);
nand U40650 (N_40650,N_40454,N_40423);
nor U40651 (N_40651,N_40416,N_40371);
and U40652 (N_40652,N_40367,N_40423);
or U40653 (N_40653,N_40479,N_40333);
nand U40654 (N_40654,N_40275,N_40442);
nor U40655 (N_40655,N_40496,N_40430);
nor U40656 (N_40656,N_40315,N_40380);
nor U40657 (N_40657,N_40251,N_40352);
and U40658 (N_40658,N_40370,N_40477);
and U40659 (N_40659,N_40277,N_40420);
xnor U40660 (N_40660,N_40418,N_40346);
or U40661 (N_40661,N_40377,N_40468);
and U40662 (N_40662,N_40258,N_40445);
and U40663 (N_40663,N_40409,N_40385);
xor U40664 (N_40664,N_40477,N_40405);
nor U40665 (N_40665,N_40482,N_40471);
nand U40666 (N_40666,N_40390,N_40417);
or U40667 (N_40667,N_40355,N_40470);
nand U40668 (N_40668,N_40268,N_40385);
and U40669 (N_40669,N_40422,N_40303);
or U40670 (N_40670,N_40405,N_40423);
or U40671 (N_40671,N_40458,N_40464);
nand U40672 (N_40672,N_40295,N_40279);
xor U40673 (N_40673,N_40318,N_40269);
or U40674 (N_40674,N_40254,N_40361);
nor U40675 (N_40675,N_40405,N_40253);
nor U40676 (N_40676,N_40403,N_40393);
or U40677 (N_40677,N_40423,N_40461);
or U40678 (N_40678,N_40279,N_40371);
and U40679 (N_40679,N_40466,N_40272);
nor U40680 (N_40680,N_40469,N_40472);
and U40681 (N_40681,N_40309,N_40416);
and U40682 (N_40682,N_40292,N_40382);
nand U40683 (N_40683,N_40491,N_40394);
and U40684 (N_40684,N_40259,N_40386);
or U40685 (N_40685,N_40288,N_40376);
or U40686 (N_40686,N_40286,N_40460);
or U40687 (N_40687,N_40330,N_40275);
xnor U40688 (N_40688,N_40371,N_40251);
and U40689 (N_40689,N_40463,N_40382);
or U40690 (N_40690,N_40256,N_40300);
nand U40691 (N_40691,N_40446,N_40371);
xnor U40692 (N_40692,N_40479,N_40474);
or U40693 (N_40693,N_40469,N_40299);
or U40694 (N_40694,N_40475,N_40424);
nor U40695 (N_40695,N_40257,N_40286);
xnor U40696 (N_40696,N_40486,N_40410);
nor U40697 (N_40697,N_40474,N_40415);
nor U40698 (N_40698,N_40377,N_40456);
xnor U40699 (N_40699,N_40482,N_40404);
xor U40700 (N_40700,N_40336,N_40488);
or U40701 (N_40701,N_40440,N_40389);
and U40702 (N_40702,N_40287,N_40439);
nand U40703 (N_40703,N_40387,N_40472);
nand U40704 (N_40704,N_40427,N_40441);
or U40705 (N_40705,N_40347,N_40361);
xnor U40706 (N_40706,N_40492,N_40287);
nand U40707 (N_40707,N_40488,N_40283);
nor U40708 (N_40708,N_40417,N_40300);
and U40709 (N_40709,N_40428,N_40427);
and U40710 (N_40710,N_40463,N_40406);
and U40711 (N_40711,N_40349,N_40358);
or U40712 (N_40712,N_40257,N_40381);
nor U40713 (N_40713,N_40485,N_40484);
nor U40714 (N_40714,N_40477,N_40273);
or U40715 (N_40715,N_40436,N_40412);
and U40716 (N_40716,N_40444,N_40446);
xnor U40717 (N_40717,N_40426,N_40274);
nand U40718 (N_40718,N_40372,N_40324);
nand U40719 (N_40719,N_40256,N_40335);
nand U40720 (N_40720,N_40444,N_40358);
xor U40721 (N_40721,N_40485,N_40440);
and U40722 (N_40722,N_40396,N_40490);
and U40723 (N_40723,N_40279,N_40485);
nor U40724 (N_40724,N_40386,N_40488);
and U40725 (N_40725,N_40434,N_40362);
nor U40726 (N_40726,N_40467,N_40456);
nor U40727 (N_40727,N_40265,N_40304);
or U40728 (N_40728,N_40498,N_40427);
xor U40729 (N_40729,N_40498,N_40384);
and U40730 (N_40730,N_40403,N_40473);
and U40731 (N_40731,N_40260,N_40297);
nand U40732 (N_40732,N_40447,N_40275);
xnor U40733 (N_40733,N_40432,N_40403);
or U40734 (N_40734,N_40346,N_40442);
and U40735 (N_40735,N_40444,N_40485);
nand U40736 (N_40736,N_40253,N_40276);
xnor U40737 (N_40737,N_40329,N_40274);
and U40738 (N_40738,N_40354,N_40265);
and U40739 (N_40739,N_40389,N_40418);
or U40740 (N_40740,N_40426,N_40291);
and U40741 (N_40741,N_40333,N_40447);
nand U40742 (N_40742,N_40324,N_40336);
nor U40743 (N_40743,N_40252,N_40372);
or U40744 (N_40744,N_40352,N_40401);
xnor U40745 (N_40745,N_40488,N_40253);
nor U40746 (N_40746,N_40262,N_40270);
or U40747 (N_40747,N_40407,N_40288);
nor U40748 (N_40748,N_40389,N_40335);
nand U40749 (N_40749,N_40426,N_40282);
and U40750 (N_40750,N_40591,N_40604);
and U40751 (N_40751,N_40624,N_40527);
or U40752 (N_40752,N_40528,N_40581);
and U40753 (N_40753,N_40608,N_40565);
and U40754 (N_40754,N_40689,N_40532);
or U40755 (N_40755,N_40630,N_40582);
nor U40756 (N_40756,N_40718,N_40526);
nand U40757 (N_40757,N_40702,N_40674);
xnor U40758 (N_40758,N_40700,N_40658);
nor U40759 (N_40759,N_40536,N_40668);
xor U40760 (N_40760,N_40729,N_40676);
or U40761 (N_40761,N_40697,N_40715);
or U40762 (N_40762,N_40606,N_40551);
xnor U40763 (N_40763,N_40745,N_40519);
xor U40764 (N_40764,N_40726,N_40665);
xnor U40765 (N_40765,N_40614,N_40675);
nand U40766 (N_40766,N_40727,N_40612);
or U40767 (N_40767,N_40620,N_40688);
nand U40768 (N_40768,N_40503,N_40705);
and U40769 (N_40769,N_40661,N_40592);
nand U40770 (N_40770,N_40641,N_40576);
xor U40771 (N_40771,N_40615,N_40564);
and U40772 (N_40772,N_40647,N_40741);
and U40773 (N_40773,N_40701,N_40622);
and U40774 (N_40774,N_40690,N_40586);
xnor U40775 (N_40775,N_40550,N_40708);
and U40776 (N_40776,N_40596,N_40502);
nor U40777 (N_40777,N_40618,N_40706);
nand U40778 (N_40778,N_40556,N_40724);
nor U40779 (N_40779,N_40572,N_40723);
xnor U40780 (N_40780,N_40683,N_40573);
and U40781 (N_40781,N_40522,N_40544);
or U40782 (N_40782,N_40590,N_40664);
nor U40783 (N_40783,N_40553,N_40722);
xnor U40784 (N_40784,N_40598,N_40512);
xnor U40785 (N_40785,N_40506,N_40578);
nor U40786 (N_40786,N_40625,N_40559);
or U40787 (N_40787,N_40687,N_40525);
nor U40788 (N_40788,N_40692,N_40736);
xor U40789 (N_40789,N_40574,N_40577);
nor U40790 (N_40790,N_40611,N_40558);
and U40791 (N_40791,N_40533,N_40694);
and U40792 (N_40792,N_40734,N_40509);
nand U40793 (N_40793,N_40642,N_40575);
and U40794 (N_40794,N_40584,N_40735);
nand U40795 (N_40795,N_40613,N_40709);
and U40796 (N_40796,N_40748,N_40649);
and U40797 (N_40797,N_40634,N_40560);
and U40798 (N_40798,N_40524,N_40638);
and U40799 (N_40799,N_40535,N_40684);
nand U40800 (N_40800,N_40742,N_40656);
nand U40801 (N_40801,N_40554,N_40653);
and U40802 (N_40802,N_40510,N_40585);
and U40803 (N_40803,N_40643,N_40568);
nor U40804 (N_40804,N_40731,N_40739);
and U40805 (N_40805,N_40547,N_40626);
or U40806 (N_40806,N_40507,N_40746);
or U40807 (N_40807,N_40707,N_40639);
xor U40808 (N_40808,N_40539,N_40619);
nor U40809 (N_40809,N_40511,N_40691);
nand U40810 (N_40810,N_40666,N_40599);
nand U40811 (N_40811,N_40579,N_40737);
nand U40812 (N_40812,N_40717,N_40500);
nor U40813 (N_40813,N_40686,N_40749);
nor U40814 (N_40814,N_40607,N_40588);
xnor U40815 (N_40815,N_40652,N_40567);
xnor U40816 (N_40816,N_40616,N_40569);
nor U40817 (N_40817,N_40530,N_40645);
or U40818 (N_40818,N_40555,N_40663);
nor U40819 (N_40819,N_40738,N_40546);
nor U40820 (N_40820,N_40662,N_40504);
and U40821 (N_40821,N_40679,N_40635);
nand U40822 (N_40822,N_40601,N_40719);
nand U40823 (N_40823,N_40670,N_40610);
nor U40824 (N_40824,N_40659,N_40743);
xnor U40825 (N_40825,N_40672,N_40721);
or U40826 (N_40826,N_40529,N_40628);
and U40827 (N_40827,N_40651,N_40521);
and U40828 (N_40828,N_40673,N_40637);
nor U40829 (N_40829,N_40516,N_40654);
xor U40830 (N_40830,N_40667,N_40699);
xor U40831 (N_40831,N_40671,N_40677);
nand U40832 (N_40832,N_40580,N_40540);
or U40833 (N_40833,N_40696,N_40703);
xor U40834 (N_40834,N_40557,N_40548);
nor U40835 (N_40835,N_40597,N_40720);
nand U40836 (N_40836,N_40605,N_40640);
and U40837 (N_40837,N_40583,N_40698);
xnor U40838 (N_40838,N_40531,N_40514);
nor U40839 (N_40839,N_40728,N_40534);
nor U40840 (N_40840,N_40595,N_40543);
xor U40841 (N_40841,N_40632,N_40566);
and U40842 (N_40842,N_40695,N_40571);
or U40843 (N_40843,N_40562,N_40740);
nand U40844 (N_40844,N_40680,N_40593);
nor U40845 (N_40845,N_40505,N_40549);
xor U40846 (N_40846,N_40542,N_40747);
nor U40847 (N_40847,N_40730,N_40693);
xor U40848 (N_40848,N_40657,N_40520);
nand U40849 (N_40849,N_40681,N_40552);
and U40850 (N_40850,N_40609,N_40600);
nor U40851 (N_40851,N_40712,N_40603);
xor U40852 (N_40852,N_40733,N_40711);
nor U40853 (N_40853,N_40660,N_40508);
and U40854 (N_40854,N_40650,N_40669);
nor U40855 (N_40855,N_40501,N_40629);
or U40856 (N_40856,N_40725,N_40631);
xor U40857 (N_40857,N_40732,N_40627);
and U40858 (N_40858,N_40716,N_40682);
nand U40859 (N_40859,N_40621,N_40713);
nor U40860 (N_40860,N_40644,N_40646);
nor U40861 (N_40861,N_40538,N_40655);
xor U40862 (N_40862,N_40537,N_40594);
and U40863 (N_40863,N_40602,N_40633);
nor U40864 (N_40864,N_40587,N_40589);
or U40865 (N_40865,N_40517,N_40561);
nor U40866 (N_40866,N_40710,N_40541);
nor U40867 (N_40867,N_40545,N_40515);
and U40868 (N_40868,N_40704,N_40563);
nand U40869 (N_40869,N_40744,N_40570);
xor U40870 (N_40870,N_40523,N_40714);
nor U40871 (N_40871,N_40648,N_40513);
nor U40872 (N_40872,N_40518,N_40685);
xor U40873 (N_40873,N_40617,N_40623);
nor U40874 (N_40874,N_40636,N_40678);
nand U40875 (N_40875,N_40737,N_40562);
or U40876 (N_40876,N_40698,N_40584);
nand U40877 (N_40877,N_40535,N_40567);
and U40878 (N_40878,N_40534,N_40746);
nand U40879 (N_40879,N_40572,N_40619);
nand U40880 (N_40880,N_40645,N_40749);
nand U40881 (N_40881,N_40571,N_40600);
nor U40882 (N_40882,N_40566,N_40523);
or U40883 (N_40883,N_40734,N_40604);
or U40884 (N_40884,N_40589,N_40684);
or U40885 (N_40885,N_40638,N_40670);
nand U40886 (N_40886,N_40735,N_40511);
nand U40887 (N_40887,N_40603,N_40651);
or U40888 (N_40888,N_40518,N_40661);
or U40889 (N_40889,N_40580,N_40742);
nand U40890 (N_40890,N_40530,N_40727);
and U40891 (N_40891,N_40545,N_40536);
xnor U40892 (N_40892,N_40742,N_40684);
xnor U40893 (N_40893,N_40558,N_40543);
nor U40894 (N_40894,N_40520,N_40629);
xnor U40895 (N_40895,N_40532,N_40707);
xnor U40896 (N_40896,N_40684,N_40717);
xor U40897 (N_40897,N_40608,N_40542);
nand U40898 (N_40898,N_40730,N_40691);
or U40899 (N_40899,N_40536,N_40588);
nor U40900 (N_40900,N_40668,N_40528);
nand U40901 (N_40901,N_40749,N_40625);
and U40902 (N_40902,N_40621,N_40636);
xor U40903 (N_40903,N_40672,N_40688);
xnor U40904 (N_40904,N_40723,N_40684);
xor U40905 (N_40905,N_40571,N_40731);
xnor U40906 (N_40906,N_40606,N_40689);
or U40907 (N_40907,N_40685,N_40721);
nand U40908 (N_40908,N_40654,N_40682);
nor U40909 (N_40909,N_40609,N_40548);
xnor U40910 (N_40910,N_40746,N_40703);
xor U40911 (N_40911,N_40735,N_40533);
or U40912 (N_40912,N_40577,N_40737);
nor U40913 (N_40913,N_40648,N_40711);
or U40914 (N_40914,N_40623,N_40697);
or U40915 (N_40915,N_40658,N_40608);
and U40916 (N_40916,N_40665,N_40591);
nand U40917 (N_40917,N_40551,N_40675);
or U40918 (N_40918,N_40596,N_40720);
xnor U40919 (N_40919,N_40703,N_40594);
and U40920 (N_40920,N_40689,N_40742);
or U40921 (N_40921,N_40681,N_40558);
nand U40922 (N_40922,N_40523,N_40560);
and U40923 (N_40923,N_40540,N_40705);
and U40924 (N_40924,N_40510,N_40749);
nor U40925 (N_40925,N_40694,N_40574);
nand U40926 (N_40926,N_40547,N_40536);
or U40927 (N_40927,N_40722,N_40558);
nor U40928 (N_40928,N_40614,N_40520);
nand U40929 (N_40929,N_40642,N_40523);
or U40930 (N_40930,N_40713,N_40648);
or U40931 (N_40931,N_40523,N_40661);
nand U40932 (N_40932,N_40625,N_40660);
xor U40933 (N_40933,N_40645,N_40649);
and U40934 (N_40934,N_40576,N_40670);
nor U40935 (N_40935,N_40545,N_40592);
nand U40936 (N_40936,N_40587,N_40623);
and U40937 (N_40937,N_40569,N_40582);
xor U40938 (N_40938,N_40552,N_40663);
and U40939 (N_40939,N_40589,N_40601);
or U40940 (N_40940,N_40536,N_40505);
or U40941 (N_40941,N_40657,N_40687);
nor U40942 (N_40942,N_40644,N_40504);
nor U40943 (N_40943,N_40554,N_40720);
nor U40944 (N_40944,N_40588,N_40676);
or U40945 (N_40945,N_40639,N_40738);
nand U40946 (N_40946,N_40535,N_40550);
xnor U40947 (N_40947,N_40617,N_40538);
nand U40948 (N_40948,N_40663,N_40591);
and U40949 (N_40949,N_40656,N_40651);
or U40950 (N_40950,N_40553,N_40693);
or U40951 (N_40951,N_40542,N_40601);
nor U40952 (N_40952,N_40727,N_40590);
nor U40953 (N_40953,N_40700,N_40634);
nand U40954 (N_40954,N_40657,N_40689);
xor U40955 (N_40955,N_40704,N_40669);
xnor U40956 (N_40956,N_40745,N_40657);
and U40957 (N_40957,N_40527,N_40594);
and U40958 (N_40958,N_40572,N_40536);
nand U40959 (N_40959,N_40724,N_40735);
nand U40960 (N_40960,N_40696,N_40561);
nor U40961 (N_40961,N_40740,N_40511);
nand U40962 (N_40962,N_40740,N_40617);
xnor U40963 (N_40963,N_40718,N_40565);
nor U40964 (N_40964,N_40577,N_40554);
nand U40965 (N_40965,N_40510,N_40528);
or U40966 (N_40966,N_40667,N_40694);
xnor U40967 (N_40967,N_40615,N_40554);
and U40968 (N_40968,N_40502,N_40660);
and U40969 (N_40969,N_40545,N_40652);
nand U40970 (N_40970,N_40664,N_40582);
or U40971 (N_40971,N_40503,N_40690);
xor U40972 (N_40972,N_40647,N_40700);
and U40973 (N_40973,N_40682,N_40589);
nand U40974 (N_40974,N_40505,N_40736);
or U40975 (N_40975,N_40739,N_40568);
or U40976 (N_40976,N_40627,N_40728);
nand U40977 (N_40977,N_40591,N_40660);
or U40978 (N_40978,N_40545,N_40569);
nand U40979 (N_40979,N_40525,N_40715);
or U40980 (N_40980,N_40691,N_40629);
or U40981 (N_40981,N_40508,N_40607);
or U40982 (N_40982,N_40554,N_40541);
and U40983 (N_40983,N_40658,N_40539);
or U40984 (N_40984,N_40579,N_40620);
or U40985 (N_40985,N_40666,N_40543);
or U40986 (N_40986,N_40682,N_40693);
or U40987 (N_40987,N_40533,N_40595);
nand U40988 (N_40988,N_40710,N_40517);
xor U40989 (N_40989,N_40583,N_40659);
nand U40990 (N_40990,N_40629,N_40632);
nor U40991 (N_40991,N_40611,N_40633);
xor U40992 (N_40992,N_40638,N_40533);
xnor U40993 (N_40993,N_40653,N_40557);
xnor U40994 (N_40994,N_40647,N_40547);
or U40995 (N_40995,N_40555,N_40556);
xor U40996 (N_40996,N_40535,N_40591);
nand U40997 (N_40997,N_40533,N_40555);
nor U40998 (N_40998,N_40597,N_40608);
nand U40999 (N_40999,N_40746,N_40743);
nand U41000 (N_41000,N_40849,N_40884);
nand U41001 (N_41001,N_40998,N_40876);
xor U41002 (N_41002,N_40861,N_40960);
nor U41003 (N_41003,N_40898,N_40970);
xor U41004 (N_41004,N_40770,N_40992);
and U41005 (N_41005,N_40886,N_40972);
or U41006 (N_41006,N_40855,N_40757);
nand U41007 (N_41007,N_40950,N_40881);
nor U41008 (N_41008,N_40979,N_40807);
and U41009 (N_41009,N_40987,N_40949);
and U41010 (N_41010,N_40818,N_40847);
or U41011 (N_41011,N_40827,N_40872);
and U41012 (N_41012,N_40813,N_40988);
nand U41013 (N_41013,N_40942,N_40844);
nand U41014 (N_41014,N_40840,N_40865);
nand U41015 (N_41015,N_40773,N_40793);
xnor U41016 (N_41016,N_40777,N_40943);
nor U41017 (N_41017,N_40941,N_40864);
nor U41018 (N_41018,N_40801,N_40805);
xor U41019 (N_41019,N_40869,N_40779);
or U41020 (N_41020,N_40764,N_40944);
nand U41021 (N_41021,N_40791,N_40752);
and U41022 (N_41022,N_40857,N_40919);
nand U41023 (N_41023,N_40897,N_40913);
and U41024 (N_41024,N_40802,N_40846);
and U41025 (N_41025,N_40783,N_40894);
xnor U41026 (N_41026,N_40831,N_40775);
and U41027 (N_41027,N_40940,N_40974);
or U41028 (N_41028,N_40795,N_40803);
nand U41029 (N_41029,N_40951,N_40910);
nor U41030 (N_41030,N_40934,N_40880);
or U41031 (N_41031,N_40997,N_40809);
nor U41032 (N_41032,N_40952,N_40948);
xor U41033 (N_41033,N_40959,N_40933);
nand U41034 (N_41034,N_40854,N_40769);
nand U41035 (N_41035,N_40782,N_40984);
nand U41036 (N_41036,N_40771,N_40772);
xnor U41037 (N_41037,N_40879,N_40895);
or U41038 (N_41038,N_40848,N_40945);
xnor U41039 (N_41039,N_40780,N_40800);
nand U41040 (N_41040,N_40862,N_40936);
or U41041 (N_41041,N_40923,N_40906);
nand U41042 (N_41042,N_40975,N_40843);
nor U41043 (N_41043,N_40928,N_40902);
nand U41044 (N_41044,N_40999,N_40893);
or U41045 (N_41045,N_40868,N_40834);
xnor U41046 (N_41046,N_40908,N_40796);
nor U41047 (N_41047,N_40966,N_40912);
or U41048 (N_41048,N_40790,N_40882);
nand U41049 (N_41049,N_40787,N_40765);
nand U41050 (N_41050,N_40767,N_40859);
nor U41051 (N_41051,N_40874,N_40851);
nand U41052 (N_41052,N_40798,N_40863);
nand U41053 (N_41053,N_40870,N_40852);
xor U41054 (N_41054,N_40938,N_40826);
nor U41055 (N_41055,N_40873,N_40930);
or U41056 (N_41056,N_40958,N_40836);
nor U41057 (N_41057,N_40918,N_40927);
and U41058 (N_41058,N_40778,N_40962);
or U41059 (N_41059,N_40968,N_40954);
xor U41060 (N_41060,N_40786,N_40808);
and U41061 (N_41061,N_40794,N_40837);
or U41062 (N_41062,N_40887,N_40961);
nor U41063 (N_41063,N_40850,N_40986);
xor U41064 (N_41064,N_40867,N_40911);
nor U41065 (N_41065,N_40955,N_40822);
and U41066 (N_41066,N_40768,N_40956);
or U41067 (N_41067,N_40866,N_40892);
nor U41068 (N_41068,N_40947,N_40996);
and U41069 (N_41069,N_40830,N_40832);
xor U41070 (N_41070,N_40839,N_40788);
nand U41071 (N_41071,N_40891,N_40842);
xor U41072 (N_41072,N_40921,N_40817);
nor U41073 (N_41073,N_40835,N_40946);
nand U41074 (N_41074,N_40823,N_40753);
or U41075 (N_41075,N_40792,N_40990);
or U41076 (N_41076,N_40751,N_40776);
or U41077 (N_41077,N_40819,N_40816);
nand U41078 (N_41078,N_40814,N_40820);
or U41079 (N_41079,N_40926,N_40759);
nor U41080 (N_41080,N_40985,N_40899);
or U41081 (N_41081,N_40905,N_40829);
xnor U41082 (N_41082,N_40924,N_40883);
nand U41083 (N_41083,N_40756,N_40754);
nand U41084 (N_41084,N_40917,N_40871);
xnor U41085 (N_41085,N_40815,N_40903);
nor U41086 (N_41086,N_40904,N_40939);
or U41087 (N_41087,N_40799,N_40824);
nor U41088 (N_41088,N_40901,N_40781);
nor U41089 (N_41089,N_40877,N_40875);
and U41090 (N_41090,N_40789,N_40810);
and U41091 (N_41091,N_40841,N_40925);
or U41092 (N_41092,N_40853,N_40878);
nand U41093 (N_41093,N_40978,N_40991);
or U41094 (N_41094,N_40900,N_40828);
or U41095 (N_41095,N_40983,N_40995);
nand U41096 (N_41096,N_40758,N_40971);
and U41097 (N_41097,N_40755,N_40856);
and U41098 (N_41098,N_40922,N_40896);
or U41099 (N_41099,N_40965,N_40797);
nor U41100 (N_41100,N_40774,N_40931);
xnor U41101 (N_41101,N_40860,N_40953);
xor U41102 (N_41102,N_40907,N_40993);
or U41103 (N_41103,N_40750,N_40785);
or U41104 (N_41104,N_40957,N_40964);
xor U41105 (N_41105,N_40760,N_40762);
and U41106 (N_41106,N_40982,N_40806);
xnor U41107 (N_41107,N_40838,N_40937);
and U41108 (N_41108,N_40890,N_40821);
nor U41109 (N_41109,N_40833,N_40812);
nand U41110 (N_41110,N_40967,N_40914);
nand U41111 (N_41111,N_40858,N_40973);
xnor U41112 (N_41112,N_40981,N_40916);
nor U41113 (N_41113,N_40784,N_40763);
xnor U41114 (N_41114,N_40845,N_40920);
xor U41115 (N_41115,N_40980,N_40889);
or U41116 (N_41116,N_40932,N_40888);
or U41117 (N_41117,N_40963,N_40929);
nor U41118 (N_41118,N_40885,N_40977);
nor U41119 (N_41119,N_40811,N_40825);
nor U41120 (N_41120,N_40766,N_40935);
nand U41121 (N_41121,N_40989,N_40976);
nor U41122 (N_41122,N_40994,N_40969);
xor U41123 (N_41123,N_40804,N_40761);
or U41124 (N_41124,N_40909,N_40915);
or U41125 (N_41125,N_40869,N_40850);
and U41126 (N_41126,N_40817,N_40887);
nand U41127 (N_41127,N_40773,N_40809);
or U41128 (N_41128,N_40954,N_40901);
and U41129 (N_41129,N_40843,N_40915);
xnor U41130 (N_41130,N_40815,N_40943);
nand U41131 (N_41131,N_40990,N_40870);
and U41132 (N_41132,N_40853,N_40843);
nor U41133 (N_41133,N_40788,N_40751);
nand U41134 (N_41134,N_40951,N_40978);
and U41135 (N_41135,N_40836,N_40979);
xnor U41136 (N_41136,N_40996,N_40755);
nor U41137 (N_41137,N_40831,N_40855);
or U41138 (N_41138,N_40830,N_40870);
nand U41139 (N_41139,N_40874,N_40918);
xor U41140 (N_41140,N_40810,N_40806);
nor U41141 (N_41141,N_40805,N_40928);
nor U41142 (N_41142,N_40777,N_40800);
nand U41143 (N_41143,N_40864,N_40903);
xor U41144 (N_41144,N_40765,N_40807);
and U41145 (N_41145,N_40789,N_40761);
nor U41146 (N_41146,N_40849,N_40787);
nor U41147 (N_41147,N_40954,N_40866);
nor U41148 (N_41148,N_40933,N_40856);
nor U41149 (N_41149,N_40860,N_40999);
and U41150 (N_41150,N_40774,N_40908);
and U41151 (N_41151,N_40923,N_40986);
xnor U41152 (N_41152,N_40985,N_40915);
or U41153 (N_41153,N_40969,N_40984);
and U41154 (N_41154,N_40933,N_40777);
and U41155 (N_41155,N_40997,N_40965);
nor U41156 (N_41156,N_40819,N_40854);
or U41157 (N_41157,N_40766,N_40872);
nor U41158 (N_41158,N_40915,N_40819);
xnor U41159 (N_41159,N_40989,N_40845);
and U41160 (N_41160,N_40845,N_40858);
or U41161 (N_41161,N_40904,N_40982);
or U41162 (N_41162,N_40891,N_40986);
and U41163 (N_41163,N_40855,N_40888);
or U41164 (N_41164,N_40831,N_40832);
nor U41165 (N_41165,N_40996,N_40778);
nor U41166 (N_41166,N_40984,N_40935);
xnor U41167 (N_41167,N_40763,N_40937);
xor U41168 (N_41168,N_40971,N_40905);
xnor U41169 (N_41169,N_40798,N_40924);
nand U41170 (N_41170,N_40986,N_40963);
or U41171 (N_41171,N_40766,N_40821);
nor U41172 (N_41172,N_40989,N_40804);
xnor U41173 (N_41173,N_40965,N_40770);
nor U41174 (N_41174,N_40792,N_40915);
nor U41175 (N_41175,N_40880,N_40864);
or U41176 (N_41176,N_40926,N_40951);
nand U41177 (N_41177,N_40787,N_40807);
or U41178 (N_41178,N_40764,N_40840);
nor U41179 (N_41179,N_40971,N_40937);
or U41180 (N_41180,N_40950,N_40882);
xor U41181 (N_41181,N_40774,N_40922);
xnor U41182 (N_41182,N_40986,N_40977);
and U41183 (N_41183,N_40851,N_40950);
nor U41184 (N_41184,N_40941,N_40758);
or U41185 (N_41185,N_40869,N_40971);
nand U41186 (N_41186,N_40808,N_40993);
or U41187 (N_41187,N_40921,N_40874);
or U41188 (N_41188,N_40840,N_40841);
nor U41189 (N_41189,N_40863,N_40770);
or U41190 (N_41190,N_40980,N_40841);
nand U41191 (N_41191,N_40898,N_40821);
nor U41192 (N_41192,N_40880,N_40767);
nor U41193 (N_41193,N_40904,N_40926);
nand U41194 (N_41194,N_40766,N_40801);
and U41195 (N_41195,N_40830,N_40958);
xnor U41196 (N_41196,N_40896,N_40872);
or U41197 (N_41197,N_40938,N_40903);
xor U41198 (N_41198,N_40760,N_40759);
nor U41199 (N_41199,N_40776,N_40917);
xor U41200 (N_41200,N_40816,N_40869);
and U41201 (N_41201,N_40953,N_40935);
nand U41202 (N_41202,N_40777,N_40849);
or U41203 (N_41203,N_40849,N_40985);
and U41204 (N_41204,N_40930,N_40931);
nor U41205 (N_41205,N_40835,N_40967);
xnor U41206 (N_41206,N_40840,N_40774);
nand U41207 (N_41207,N_40846,N_40923);
nand U41208 (N_41208,N_40861,N_40903);
nand U41209 (N_41209,N_40918,N_40957);
xnor U41210 (N_41210,N_40788,N_40835);
xor U41211 (N_41211,N_40996,N_40792);
nand U41212 (N_41212,N_40884,N_40821);
or U41213 (N_41213,N_40769,N_40917);
and U41214 (N_41214,N_40756,N_40765);
nor U41215 (N_41215,N_40812,N_40948);
nand U41216 (N_41216,N_40758,N_40896);
nand U41217 (N_41217,N_40815,N_40782);
xnor U41218 (N_41218,N_40971,N_40962);
xor U41219 (N_41219,N_40896,N_40771);
or U41220 (N_41220,N_40947,N_40862);
and U41221 (N_41221,N_40969,N_40790);
xor U41222 (N_41222,N_40812,N_40964);
xor U41223 (N_41223,N_40965,N_40897);
and U41224 (N_41224,N_40931,N_40902);
nand U41225 (N_41225,N_40973,N_40970);
nand U41226 (N_41226,N_40938,N_40900);
and U41227 (N_41227,N_40973,N_40977);
nor U41228 (N_41228,N_40878,N_40758);
xnor U41229 (N_41229,N_40952,N_40774);
nand U41230 (N_41230,N_40933,N_40807);
xor U41231 (N_41231,N_40826,N_40798);
nor U41232 (N_41232,N_40803,N_40859);
nor U41233 (N_41233,N_40782,N_40830);
nor U41234 (N_41234,N_40915,N_40988);
and U41235 (N_41235,N_40942,N_40753);
xor U41236 (N_41236,N_40882,N_40870);
or U41237 (N_41237,N_40824,N_40911);
nor U41238 (N_41238,N_40905,N_40757);
or U41239 (N_41239,N_40777,N_40981);
or U41240 (N_41240,N_40941,N_40966);
and U41241 (N_41241,N_40781,N_40907);
nand U41242 (N_41242,N_40901,N_40839);
and U41243 (N_41243,N_40986,N_40826);
nand U41244 (N_41244,N_40933,N_40957);
xor U41245 (N_41245,N_40755,N_40997);
nor U41246 (N_41246,N_40871,N_40987);
or U41247 (N_41247,N_40792,N_40987);
nand U41248 (N_41248,N_40922,N_40785);
or U41249 (N_41249,N_40956,N_40754);
nor U41250 (N_41250,N_41151,N_41036);
xor U41251 (N_41251,N_41218,N_41249);
nor U41252 (N_41252,N_41243,N_41008);
nand U41253 (N_41253,N_41100,N_41232);
xor U41254 (N_41254,N_41124,N_41179);
nand U41255 (N_41255,N_41067,N_41031);
nand U41256 (N_41256,N_41180,N_41012);
nor U41257 (N_41257,N_41207,N_41188);
nor U41258 (N_41258,N_41087,N_41234);
or U41259 (N_41259,N_41119,N_41158);
xnor U41260 (N_41260,N_41189,N_41101);
xor U41261 (N_41261,N_41061,N_41133);
xnor U41262 (N_41262,N_41168,N_41051);
and U41263 (N_41263,N_41090,N_41111);
nand U41264 (N_41264,N_41171,N_41149);
nor U41265 (N_41265,N_41023,N_41214);
nand U41266 (N_41266,N_41088,N_41058);
nand U41267 (N_41267,N_41081,N_41070);
nand U41268 (N_41268,N_41182,N_41103);
or U41269 (N_41269,N_41178,N_41127);
or U41270 (N_41270,N_41046,N_41230);
and U41271 (N_41271,N_41219,N_41229);
xnor U41272 (N_41272,N_41037,N_41237);
xnor U41273 (N_41273,N_41113,N_41045);
nand U41274 (N_41274,N_41160,N_41241);
nor U41275 (N_41275,N_41123,N_41130);
nand U41276 (N_41276,N_41034,N_41060);
nor U41277 (N_41277,N_41244,N_41152);
nor U41278 (N_41278,N_41122,N_41226);
nor U41279 (N_41279,N_41108,N_41195);
and U41280 (N_41280,N_41215,N_41005);
nor U41281 (N_41281,N_41246,N_41161);
nand U41282 (N_41282,N_41013,N_41191);
nand U41283 (N_41283,N_41135,N_41239);
nand U41284 (N_41284,N_41131,N_41083);
and U41285 (N_41285,N_41173,N_41212);
or U41286 (N_41286,N_41099,N_41233);
nand U41287 (N_41287,N_41148,N_41019);
xor U41288 (N_41288,N_41063,N_41002);
or U41289 (N_41289,N_41021,N_41150);
xnor U41290 (N_41290,N_41086,N_41194);
nand U41291 (N_41291,N_41221,N_41129);
xor U41292 (N_41292,N_41105,N_41136);
or U41293 (N_41293,N_41145,N_41084);
nand U41294 (N_41294,N_41153,N_41039);
xnor U41295 (N_41295,N_41052,N_41071);
nand U41296 (N_41296,N_41033,N_41196);
or U41297 (N_41297,N_41177,N_41096);
nor U41298 (N_41298,N_41125,N_41154);
nand U41299 (N_41299,N_41020,N_41128);
nor U41300 (N_41300,N_41235,N_41211);
nand U41301 (N_41301,N_41059,N_41042);
or U41302 (N_41302,N_41216,N_41174);
xor U41303 (N_41303,N_41007,N_41104);
xor U41304 (N_41304,N_41015,N_41139);
nor U41305 (N_41305,N_41077,N_41082);
or U41306 (N_41306,N_41075,N_41032);
or U41307 (N_41307,N_41176,N_41202);
and U41308 (N_41308,N_41028,N_41132);
and U41309 (N_41309,N_41134,N_41085);
or U41310 (N_41310,N_41035,N_41025);
or U41311 (N_41311,N_41116,N_41026);
and U41312 (N_41312,N_41224,N_41048);
and U41313 (N_41313,N_41047,N_41172);
xor U41314 (N_41314,N_41198,N_41022);
nor U41315 (N_41315,N_41240,N_41092);
nand U41316 (N_41316,N_41068,N_41017);
xnor U41317 (N_41317,N_41199,N_41155);
nor U41318 (N_41318,N_41109,N_41112);
nor U41319 (N_41319,N_41044,N_41187);
or U41320 (N_41320,N_41225,N_41089);
or U41321 (N_41321,N_41078,N_41009);
nand U41322 (N_41322,N_41102,N_41016);
or U41323 (N_41323,N_41091,N_41076);
nor U41324 (N_41324,N_41064,N_41098);
nand U41325 (N_41325,N_41049,N_41030);
xor U41326 (N_41326,N_41093,N_41223);
and U41327 (N_41327,N_41117,N_41118);
nand U41328 (N_41328,N_41186,N_41231);
nand U41329 (N_41329,N_41114,N_41120);
and U41330 (N_41330,N_41062,N_41065);
nand U41331 (N_41331,N_41000,N_41011);
or U41332 (N_41332,N_41147,N_41001);
xor U41333 (N_41333,N_41192,N_41073);
or U41334 (N_41334,N_41209,N_41074);
nand U41335 (N_41335,N_41213,N_41069);
nand U41336 (N_41336,N_41228,N_41167);
xnor U41337 (N_41337,N_41054,N_41126);
xor U41338 (N_41338,N_41175,N_41050);
nor U41339 (N_41339,N_41157,N_41055);
nor U41340 (N_41340,N_41095,N_41041);
nand U41341 (N_41341,N_41185,N_41138);
and U41342 (N_41342,N_41197,N_41206);
nor U41343 (N_41343,N_41003,N_41027);
or U41344 (N_41344,N_41205,N_41204);
xor U41345 (N_41345,N_41066,N_41115);
xnor U41346 (N_41346,N_41220,N_41106);
or U41347 (N_41347,N_41018,N_41043);
and U41348 (N_41348,N_41137,N_41165);
nor U41349 (N_41349,N_41024,N_41222);
nor U41350 (N_41350,N_41181,N_41142);
and U41351 (N_41351,N_41203,N_41164);
xor U41352 (N_41352,N_41163,N_41201);
or U41353 (N_41353,N_41227,N_41004);
xnor U41354 (N_41354,N_41038,N_41040);
nor U41355 (N_41355,N_41121,N_41238);
and U41356 (N_41356,N_41006,N_41242);
and U41357 (N_41357,N_41146,N_41190);
or U41358 (N_41358,N_41208,N_41079);
or U41359 (N_41359,N_41236,N_41141);
nand U41360 (N_41360,N_41169,N_41144);
xnor U41361 (N_41361,N_41248,N_41210);
nand U41362 (N_41362,N_41056,N_41053);
xnor U41363 (N_41363,N_41094,N_41072);
nand U41364 (N_41364,N_41110,N_41247);
or U41365 (N_41365,N_41097,N_41200);
and U41366 (N_41366,N_41080,N_41159);
nor U41367 (N_41367,N_41010,N_41183);
nand U41368 (N_41368,N_41166,N_41140);
nand U41369 (N_41369,N_41156,N_41029);
nand U41370 (N_41370,N_41107,N_41193);
or U41371 (N_41371,N_41245,N_41162);
xnor U41372 (N_41372,N_41170,N_41143);
nand U41373 (N_41373,N_41217,N_41184);
and U41374 (N_41374,N_41057,N_41014);
nand U41375 (N_41375,N_41063,N_41186);
nand U41376 (N_41376,N_41145,N_41066);
nor U41377 (N_41377,N_41130,N_41093);
and U41378 (N_41378,N_41068,N_41089);
nand U41379 (N_41379,N_41203,N_41108);
or U41380 (N_41380,N_41103,N_41029);
and U41381 (N_41381,N_41236,N_41248);
and U41382 (N_41382,N_41190,N_41140);
nor U41383 (N_41383,N_41153,N_41192);
xnor U41384 (N_41384,N_41152,N_41221);
and U41385 (N_41385,N_41134,N_41028);
nor U41386 (N_41386,N_41139,N_41221);
xnor U41387 (N_41387,N_41089,N_41116);
nor U41388 (N_41388,N_41235,N_41204);
or U41389 (N_41389,N_41103,N_41159);
nand U41390 (N_41390,N_41078,N_41187);
xor U41391 (N_41391,N_41052,N_41244);
xnor U41392 (N_41392,N_41069,N_41178);
or U41393 (N_41393,N_41049,N_41037);
xor U41394 (N_41394,N_41157,N_41034);
nand U41395 (N_41395,N_41036,N_41125);
or U41396 (N_41396,N_41083,N_41212);
or U41397 (N_41397,N_41223,N_41167);
xor U41398 (N_41398,N_41062,N_41071);
and U41399 (N_41399,N_41206,N_41054);
xnor U41400 (N_41400,N_41108,N_41199);
and U41401 (N_41401,N_41239,N_41220);
or U41402 (N_41402,N_41094,N_41073);
and U41403 (N_41403,N_41057,N_41044);
nor U41404 (N_41404,N_41018,N_41111);
or U41405 (N_41405,N_41132,N_41234);
nand U41406 (N_41406,N_41053,N_41033);
nand U41407 (N_41407,N_41070,N_41113);
and U41408 (N_41408,N_41167,N_41247);
or U41409 (N_41409,N_41232,N_41111);
or U41410 (N_41410,N_41026,N_41193);
and U41411 (N_41411,N_41072,N_41103);
nor U41412 (N_41412,N_41185,N_41058);
xnor U41413 (N_41413,N_41139,N_41151);
and U41414 (N_41414,N_41111,N_41210);
or U41415 (N_41415,N_41142,N_41198);
xnor U41416 (N_41416,N_41231,N_41044);
or U41417 (N_41417,N_41202,N_41174);
nand U41418 (N_41418,N_41227,N_41070);
nor U41419 (N_41419,N_41031,N_41190);
and U41420 (N_41420,N_41003,N_41036);
nor U41421 (N_41421,N_41201,N_41249);
xor U41422 (N_41422,N_41079,N_41163);
or U41423 (N_41423,N_41199,N_41022);
nor U41424 (N_41424,N_41190,N_41112);
or U41425 (N_41425,N_41232,N_41124);
and U41426 (N_41426,N_41007,N_41008);
or U41427 (N_41427,N_41230,N_41146);
or U41428 (N_41428,N_41021,N_41104);
nor U41429 (N_41429,N_41040,N_41136);
xor U41430 (N_41430,N_41192,N_41246);
nor U41431 (N_41431,N_41191,N_41105);
or U41432 (N_41432,N_41194,N_41060);
and U41433 (N_41433,N_41090,N_41083);
and U41434 (N_41434,N_41003,N_41183);
xor U41435 (N_41435,N_41066,N_41161);
xor U41436 (N_41436,N_41086,N_41180);
xor U41437 (N_41437,N_41015,N_41009);
nor U41438 (N_41438,N_41036,N_41178);
nor U41439 (N_41439,N_41210,N_41162);
nand U41440 (N_41440,N_41041,N_41182);
nand U41441 (N_41441,N_41010,N_41169);
nand U41442 (N_41442,N_41134,N_41111);
or U41443 (N_41443,N_41017,N_41045);
nor U41444 (N_41444,N_41158,N_41140);
or U41445 (N_41445,N_41178,N_41061);
nand U41446 (N_41446,N_41235,N_41210);
and U41447 (N_41447,N_41246,N_41049);
nor U41448 (N_41448,N_41243,N_41070);
or U41449 (N_41449,N_41158,N_41202);
nand U41450 (N_41450,N_41200,N_41236);
nand U41451 (N_41451,N_41138,N_41021);
nor U41452 (N_41452,N_41248,N_41146);
and U41453 (N_41453,N_41086,N_41178);
and U41454 (N_41454,N_41213,N_41242);
nand U41455 (N_41455,N_41127,N_41041);
nor U41456 (N_41456,N_41091,N_41097);
xor U41457 (N_41457,N_41177,N_41061);
nor U41458 (N_41458,N_41002,N_41125);
nand U41459 (N_41459,N_41137,N_41122);
or U41460 (N_41460,N_41004,N_41233);
nand U41461 (N_41461,N_41059,N_41197);
and U41462 (N_41462,N_41241,N_41083);
or U41463 (N_41463,N_41011,N_41043);
or U41464 (N_41464,N_41034,N_41089);
and U41465 (N_41465,N_41081,N_41146);
nand U41466 (N_41466,N_41002,N_41034);
nand U41467 (N_41467,N_41004,N_41175);
nand U41468 (N_41468,N_41034,N_41131);
and U41469 (N_41469,N_41046,N_41223);
and U41470 (N_41470,N_41181,N_41225);
or U41471 (N_41471,N_41121,N_41158);
and U41472 (N_41472,N_41232,N_41198);
xnor U41473 (N_41473,N_41207,N_41235);
and U41474 (N_41474,N_41140,N_41012);
nand U41475 (N_41475,N_41133,N_41060);
nor U41476 (N_41476,N_41054,N_41207);
xor U41477 (N_41477,N_41113,N_41046);
nand U41478 (N_41478,N_41249,N_41185);
nor U41479 (N_41479,N_41097,N_41215);
nand U41480 (N_41480,N_41039,N_41048);
nor U41481 (N_41481,N_41154,N_41214);
nand U41482 (N_41482,N_41044,N_41176);
xnor U41483 (N_41483,N_41067,N_41178);
xor U41484 (N_41484,N_41205,N_41198);
or U41485 (N_41485,N_41194,N_41203);
and U41486 (N_41486,N_41009,N_41017);
or U41487 (N_41487,N_41245,N_41126);
nand U41488 (N_41488,N_41035,N_41075);
nor U41489 (N_41489,N_41057,N_41142);
nand U41490 (N_41490,N_41053,N_41184);
nand U41491 (N_41491,N_41156,N_41201);
xnor U41492 (N_41492,N_41116,N_41140);
nor U41493 (N_41493,N_41178,N_41084);
xnor U41494 (N_41494,N_41119,N_41052);
or U41495 (N_41495,N_41165,N_41055);
or U41496 (N_41496,N_41110,N_41240);
nand U41497 (N_41497,N_41246,N_41191);
xnor U41498 (N_41498,N_41229,N_41168);
xor U41499 (N_41499,N_41136,N_41109);
and U41500 (N_41500,N_41395,N_41329);
xnor U41501 (N_41501,N_41385,N_41382);
and U41502 (N_41502,N_41433,N_41496);
xnor U41503 (N_41503,N_41250,N_41441);
or U41504 (N_41504,N_41414,N_41381);
or U41505 (N_41505,N_41430,N_41324);
or U41506 (N_41506,N_41447,N_41343);
nand U41507 (N_41507,N_41471,N_41393);
or U41508 (N_41508,N_41478,N_41431);
xor U41509 (N_41509,N_41336,N_41341);
xnor U41510 (N_41510,N_41256,N_41263);
or U41511 (N_41511,N_41379,N_41428);
nor U41512 (N_41512,N_41436,N_41299);
nand U41513 (N_41513,N_41347,N_41339);
and U41514 (N_41514,N_41309,N_41439);
and U41515 (N_41515,N_41365,N_41456);
or U41516 (N_41516,N_41357,N_41330);
nor U41517 (N_41517,N_41313,N_41396);
or U41518 (N_41518,N_41260,N_41335);
xnor U41519 (N_41519,N_41409,N_41432);
or U41520 (N_41520,N_41371,N_41278);
nor U41521 (N_41521,N_41453,N_41367);
nor U41522 (N_41522,N_41298,N_41307);
xnor U41523 (N_41523,N_41295,N_41283);
or U41524 (N_41524,N_41304,N_41454);
or U41525 (N_41525,N_41477,N_41459);
nand U41526 (N_41526,N_41391,N_41362);
nand U41527 (N_41527,N_41464,N_41406);
nand U41528 (N_41528,N_41261,N_41269);
or U41529 (N_41529,N_41489,N_41467);
and U41530 (N_41530,N_41272,N_41302);
nor U41531 (N_41531,N_41444,N_41384);
and U41532 (N_41532,N_41495,N_41306);
or U41533 (N_41533,N_41415,N_41413);
nor U41534 (N_41534,N_41325,N_41494);
nand U41535 (N_41535,N_41290,N_41344);
nor U41536 (N_41536,N_41401,N_41312);
xor U41537 (N_41537,N_41280,N_41363);
nand U41538 (N_41538,N_41294,N_41271);
or U41539 (N_41539,N_41282,N_41277);
and U41540 (N_41540,N_41317,N_41468);
and U41541 (N_41541,N_41403,N_41398);
nand U41542 (N_41542,N_41326,N_41355);
xnor U41543 (N_41543,N_41440,N_41493);
or U41544 (N_41544,N_41268,N_41319);
xnor U41545 (N_41545,N_41276,N_41389);
xnor U41546 (N_41546,N_41476,N_41497);
or U41547 (N_41547,N_41498,N_41419);
and U41548 (N_41548,N_41404,N_41418);
nor U41549 (N_41549,N_41351,N_41486);
or U41550 (N_41550,N_41472,N_41321);
and U41551 (N_41551,N_41352,N_41469);
and U41552 (N_41552,N_41342,N_41303);
nand U41553 (N_41553,N_41264,N_41460);
nor U41554 (N_41554,N_41289,N_41411);
xnor U41555 (N_41555,N_41465,N_41358);
or U41556 (N_41556,N_41443,N_41457);
xor U41557 (N_41557,N_41254,N_41296);
or U41558 (N_41558,N_41338,N_41425);
or U41559 (N_41559,N_41253,N_41373);
xor U41560 (N_41560,N_41463,N_41259);
nor U41561 (N_41561,N_41257,N_41458);
xor U41562 (N_41562,N_41314,N_41420);
and U41563 (N_41563,N_41349,N_41387);
and U41564 (N_41564,N_41388,N_41446);
or U41565 (N_41565,N_41286,N_41340);
nand U41566 (N_41566,N_41499,N_41482);
nor U41567 (N_41567,N_41328,N_41399);
nand U41568 (N_41568,N_41251,N_41354);
xor U41569 (N_41569,N_41284,N_41374);
or U41570 (N_41570,N_41356,N_41265);
nand U41571 (N_41571,N_41270,N_41485);
nor U41572 (N_41572,N_41466,N_41273);
nand U41573 (N_41573,N_41287,N_41490);
and U41574 (N_41574,N_41410,N_41455);
and U41575 (N_41575,N_41305,N_41377);
xnor U41576 (N_41576,N_41421,N_41332);
and U41577 (N_41577,N_41293,N_41318);
and U41578 (N_41578,N_41434,N_41281);
nor U41579 (N_41579,N_41474,N_41424);
nand U41580 (N_41580,N_41255,N_41450);
nor U41581 (N_41581,N_41481,N_41488);
and U41582 (N_41582,N_41400,N_41479);
nand U41583 (N_41583,N_41375,N_41442);
and U41584 (N_41584,N_41475,N_41452);
xor U41585 (N_41585,N_41266,N_41274);
or U41586 (N_41586,N_41372,N_41405);
xor U41587 (N_41587,N_41445,N_41364);
xnor U41588 (N_41588,N_41423,N_41448);
and U41589 (N_41589,N_41470,N_41297);
xor U41590 (N_41590,N_41315,N_41383);
xor U41591 (N_41591,N_41291,N_41386);
and U41592 (N_41592,N_41300,N_41333);
nand U41593 (N_41593,N_41369,N_41301);
and U41594 (N_41594,N_41310,N_41361);
nor U41595 (N_41595,N_41451,N_41360);
xnor U41596 (N_41596,N_41334,N_41473);
or U41597 (N_41597,N_41359,N_41327);
nand U41598 (N_41598,N_41368,N_41353);
and U41599 (N_41599,N_41480,N_41461);
nand U41600 (N_41600,N_41412,N_41346);
xor U41601 (N_41601,N_41279,N_41438);
nor U41602 (N_41602,N_41366,N_41275);
nand U41603 (N_41603,N_41390,N_41392);
xnor U41604 (N_41604,N_41427,N_41402);
nand U41605 (N_41605,N_41417,N_41378);
nor U41606 (N_41606,N_41311,N_41337);
nand U41607 (N_41607,N_41380,N_41331);
and U41608 (N_41608,N_41348,N_41487);
nand U41609 (N_41609,N_41350,N_41394);
and U41610 (N_41610,N_41437,N_41407);
xnor U41611 (N_41611,N_41462,N_41397);
and U41612 (N_41612,N_41252,N_41370);
and U41613 (N_41613,N_41345,N_41376);
nand U41614 (N_41614,N_41416,N_41323);
and U41615 (N_41615,N_41449,N_41316);
nand U41616 (N_41616,N_41320,N_41491);
and U41617 (N_41617,N_41408,N_41262);
or U41618 (N_41618,N_41484,N_41288);
and U41619 (N_41619,N_41483,N_41426);
nand U41620 (N_41620,N_41322,N_41422);
nand U41621 (N_41621,N_41435,N_41267);
nand U41622 (N_41622,N_41308,N_41292);
nor U41623 (N_41623,N_41258,N_41285);
nand U41624 (N_41624,N_41492,N_41429);
nor U41625 (N_41625,N_41431,N_41385);
nor U41626 (N_41626,N_41294,N_41490);
nor U41627 (N_41627,N_41383,N_41349);
xor U41628 (N_41628,N_41383,N_41302);
nor U41629 (N_41629,N_41256,N_41435);
and U41630 (N_41630,N_41307,N_41390);
xnor U41631 (N_41631,N_41277,N_41488);
xnor U41632 (N_41632,N_41498,N_41416);
xor U41633 (N_41633,N_41306,N_41419);
nand U41634 (N_41634,N_41333,N_41471);
xor U41635 (N_41635,N_41338,N_41367);
nand U41636 (N_41636,N_41381,N_41257);
nor U41637 (N_41637,N_41293,N_41334);
and U41638 (N_41638,N_41347,N_41318);
xnor U41639 (N_41639,N_41307,N_41364);
xor U41640 (N_41640,N_41494,N_41363);
and U41641 (N_41641,N_41349,N_41400);
and U41642 (N_41642,N_41269,N_41277);
and U41643 (N_41643,N_41356,N_41361);
or U41644 (N_41644,N_41443,N_41290);
and U41645 (N_41645,N_41290,N_41404);
xor U41646 (N_41646,N_41479,N_41401);
or U41647 (N_41647,N_41308,N_41487);
nand U41648 (N_41648,N_41272,N_41491);
xnor U41649 (N_41649,N_41284,N_41473);
nor U41650 (N_41650,N_41345,N_41493);
nand U41651 (N_41651,N_41415,N_41469);
or U41652 (N_41652,N_41434,N_41277);
nor U41653 (N_41653,N_41449,N_41298);
and U41654 (N_41654,N_41348,N_41443);
and U41655 (N_41655,N_41391,N_41289);
or U41656 (N_41656,N_41484,N_41342);
xnor U41657 (N_41657,N_41470,N_41347);
nand U41658 (N_41658,N_41318,N_41458);
nor U41659 (N_41659,N_41397,N_41316);
xnor U41660 (N_41660,N_41266,N_41370);
or U41661 (N_41661,N_41269,N_41310);
or U41662 (N_41662,N_41498,N_41478);
nor U41663 (N_41663,N_41291,N_41437);
nand U41664 (N_41664,N_41440,N_41460);
or U41665 (N_41665,N_41492,N_41482);
xor U41666 (N_41666,N_41462,N_41296);
nand U41667 (N_41667,N_41252,N_41303);
and U41668 (N_41668,N_41284,N_41458);
nand U41669 (N_41669,N_41420,N_41389);
xor U41670 (N_41670,N_41289,N_41382);
or U41671 (N_41671,N_41444,N_41291);
or U41672 (N_41672,N_41349,N_41462);
nor U41673 (N_41673,N_41286,N_41392);
xnor U41674 (N_41674,N_41417,N_41343);
nand U41675 (N_41675,N_41297,N_41433);
and U41676 (N_41676,N_41413,N_41342);
and U41677 (N_41677,N_41345,N_41492);
or U41678 (N_41678,N_41477,N_41367);
nor U41679 (N_41679,N_41460,N_41491);
xnor U41680 (N_41680,N_41364,N_41428);
and U41681 (N_41681,N_41303,N_41391);
nand U41682 (N_41682,N_41333,N_41402);
and U41683 (N_41683,N_41462,N_41300);
or U41684 (N_41684,N_41477,N_41438);
nor U41685 (N_41685,N_41346,N_41336);
nor U41686 (N_41686,N_41428,N_41393);
and U41687 (N_41687,N_41403,N_41466);
or U41688 (N_41688,N_41417,N_41407);
and U41689 (N_41689,N_41325,N_41464);
nand U41690 (N_41690,N_41484,N_41388);
xor U41691 (N_41691,N_41326,N_41397);
nor U41692 (N_41692,N_41346,N_41252);
and U41693 (N_41693,N_41299,N_41252);
nor U41694 (N_41694,N_41270,N_41312);
nor U41695 (N_41695,N_41492,N_41480);
and U41696 (N_41696,N_41301,N_41306);
nand U41697 (N_41697,N_41427,N_41417);
nor U41698 (N_41698,N_41261,N_41330);
nand U41699 (N_41699,N_41449,N_41269);
and U41700 (N_41700,N_41328,N_41257);
or U41701 (N_41701,N_41253,N_41391);
and U41702 (N_41702,N_41486,N_41496);
nor U41703 (N_41703,N_41456,N_41400);
nor U41704 (N_41704,N_41384,N_41406);
xor U41705 (N_41705,N_41277,N_41337);
or U41706 (N_41706,N_41494,N_41468);
nand U41707 (N_41707,N_41342,N_41458);
nor U41708 (N_41708,N_41323,N_41451);
nand U41709 (N_41709,N_41265,N_41456);
nor U41710 (N_41710,N_41444,N_41455);
nand U41711 (N_41711,N_41387,N_41481);
xnor U41712 (N_41712,N_41358,N_41254);
and U41713 (N_41713,N_41355,N_41354);
nor U41714 (N_41714,N_41356,N_41381);
xor U41715 (N_41715,N_41406,N_41454);
nor U41716 (N_41716,N_41461,N_41302);
xnor U41717 (N_41717,N_41305,N_41252);
or U41718 (N_41718,N_41278,N_41368);
or U41719 (N_41719,N_41281,N_41478);
xor U41720 (N_41720,N_41388,N_41335);
nand U41721 (N_41721,N_41308,N_41415);
nand U41722 (N_41722,N_41250,N_41310);
nand U41723 (N_41723,N_41484,N_41363);
and U41724 (N_41724,N_41416,N_41277);
or U41725 (N_41725,N_41382,N_41431);
nand U41726 (N_41726,N_41489,N_41373);
xnor U41727 (N_41727,N_41331,N_41349);
xor U41728 (N_41728,N_41341,N_41311);
nor U41729 (N_41729,N_41303,N_41329);
nand U41730 (N_41730,N_41333,N_41449);
nor U41731 (N_41731,N_41421,N_41309);
xnor U41732 (N_41732,N_41484,N_41298);
and U41733 (N_41733,N_41264,N_41263);
nand U41734 (N_41734,N_41279,N_41422);
or U41735 (N_41735,N_41390,N_41304);
nor U41736 (N_41736,N_41283,N_41431);
and U41737 (N_41737,N_41400,N_41407);
and U41738 (N_41738,N_41265,N_41294);
or U41739 (N_41739,N_41358,N_41415);
nor U41740 (N_41740,N_41324,N_41322);
nand U41741 (N_41741,N_41275,N_41386);
nand U41742 (N_41742,N_41372,N_41495);
xor U41743 (N_41743,N_41312,N_41366);
nand U41744 (N_41744,N_41471,N_41272);
nor U41745 (N_41745,N_41294,N_41291);
and U41746 (N_41746,N_41393,N_41275);
nand U41747 (N_41747,N_41277,N_41464);
or U41748 (N_41748,N_41325,N_41339);
xor U41749 (N_41749,N_41279,N_41355);
or U41750 (N_41750,N_41538,N_41653);
or U41751 (N_41751,N_41605,N_41522);
or U41752 (N_41752,N_41564,N_41740);
xnor U41753 (N_41753,N_41700,N_41717);
nor U41754 (N_41754,N_41612,N_41649);
nor U41755 (N_41755,N_41594,N_41609);
nor U41756 (N_41756,N_41579,N_41725);
and U41757 (N_41757,N_41550,N_41684);
nor U41758 (N_41758,N_41505,N_41610);
nor U41759 (N_41759,N_41566,N_41542);
nor U41760 (N_41760,N_41628,N_41697);
xor U41761 (N_41761,N_41748,N_41694);
or U41762 (N_41762,N_41691,N_41651);
or U41763 (N_41763,N_41529,N_41576);
or U41764 (N_41764,N_41709,N_41570);
or U41765 (N_41765,N_41561,N_41670);
or U41766 (N_41766,N_41549,N_41531);
nor U41767 (N_41767,N_41701,N_41723);
or U41768 (N_41768,N_41568,N_41682);
or U41769 (N_41769,N_41585,N_41686);
xor U41770 (N_41770,N_41577,N_41619);
nand U41771 (N_41771,N_41597,N_41571);
and U41772 (N_41772,N_41702,N_41528);
nor U41773 (N_41773,N_41526,N_41679);
and U41774 (N_41774,N_41535,N_41506);
xor U41775 (N_41775,N_41690,N_41616);
or U41776 (N_41776,N_41518,N_41569);
or U41777 (N_41777,N_41642,N_41687);
xnor U41778 (N_41778,N_41662,N_41710);
xor U41779 (N_41779,N_41713,N_41510);
and U41780 (N_41780,N_41689,N_41606);
and U41781 (N_41781,N_41509,N_41530);
xnor U41782 (N_41782,N_41501,N_41553);
and U41783 (N_41783,N_41622,N_41504);
or U41784 (N_41784,N_41695,N_41588);
and U41785 (N_41785,N_41673,N_41692);
and U41786 (N_41786,N_41560,N_41574);
and U41787 (N_41787,N_41627,N_41672);
and U41788 (N_41788,N_41696,N_41615);
or U41789 (N_41789,N_41527,N_41693);
nor U41790 (N_41790,N_41500,N_41507);
xnor U41791 (N_41791,N_41715,N_41688);
and U41792 (N_41792,N_41720,N_41664);
and U41793 (N_41793,N_41646,N_41533);
nor U41794 (N_41794,N_41729,N_41556);
and U41795 (N_41795,N_41681,N_41573);
or U41796 (N_41796,N_41513,N_41659);
nor U41797 (N_41797,N_41599,N_41661);
or U41798 (N_41798,N_41674,N_41601);
nand U41799 (N_41799,N_41708,N_41562);
xnor U41800 (N_41800,N_41704,N_41727);
nor U41801 (N_41801,N_41584,N_41743);
nand U41802 (N_41802,N_41544,N_41712);
and U41803 (N_41803,N_41706,N_41563);
nand U41804 (N_41804,N_41637,N_41516);
or U41805 (N_41805,N_41617,N_41521);
or U41806 (N_41806,N_41738,N_41671);
nand U41807 (N_41807,N_41640,N_41532);
xor U41808 (N_41808,N_41590,N_41534);
or U41809 (N_41809,N_41719,N_41714);
nand U41810 (N_41810,N_41592,N_41643);
nor U41811 (N_41811,N_41678,N_41536);
and U41812 (N_41812,N_41677,N_41554);
nor U41813 (N_41813,N_41520,N_41578);
or U41814 (N_41814,N_41555,N_41647);
nand U41815 (N_41815,N_41508,N_41722);
nor U41816 (N_41816,N_41613,N_41596);
or U41817 (N_41817,N_41517,N_41567);
or U41818 (N_41818,N_41648,N_41663);
nor U41819 (N_41819,N_41511,N_41650);
nor U41820 (N_41820,N_41730,N_41739);
nor U41821 (N_41821,N_41742,N_41565);
nor U41822 (N_41822,N_41666,N_41707);
xor U41823 (N_41823,N_41736,N_41598);
nor U41824 (N_41824,N_41749,N_41698);
nand U41825 (N_41825,N_41502,N_41669);
and U41826 (N_41826,N_41623,N_41515);
or U41827 (N_41827,N_41558,N_41525);
nor U41828 (N_41828,N_41635,N_41658);
or U41829 (N_41829,N_41572,N_41524);
xnor U41830 (N_41830,N_41726,N_41718);
xor U41831 (N_41831,N_41523,N_41741);
or U41832 (N_41832,N_41639,N_41655);
or U41833 (N_41833,N_41582,N_41746);
nor U41834 (N_41834,N_41614,N_41620);
and U41835 (N_41835,N_41607,N_41641);
and U41836 (N_41836,N_41699,N_41625);
nor U41837 (N_41837,N_41675,N_41703);
nor U41838 (N_41838,N_41512,N_41589);
or U41839 (N_41839,N_41546,N_41668);
and U41840 (N_41840,N_41548,N_41733);
nand U41841 (N_41841,N_41737,N_41503);
and U41842 (N_41842,N_41618,N_41514);
and U41843 (N_41843,N_41735,N_41552);
nor U41844 (N_41844,N_41747,N_41541);
or U41845 (N_41845,N_41645,N_41630);
and U41846 (N_41846,N_41543,N_41745);
xnor U41847 (N_41847,N_41629,N_41634);
and U41848 (N_41848,N_41636,N_41665);
xor U41849 (N_41849,N_41683,N_41680);
xor U41850 (N_41850,N_41657,N_41652);
and U41851 (N_41851,N_41644,N_41731);
and U41852 (N_41852,N_41600,N_41575);
xor U41853 (N_41853,N_41581,N_41580);
nor U41854 (N_41854,N_41602,N_41728);
and U41855 (N_41855,N_41586,N_41631);
xnor U41856 (N_41856,N_41626,N_41608);
nand U41857 (N_41857,N_41557,N_41545);
or U41858 (N_41858,N_41732,N_41721);
nand U41859 (N_41859,N_41667,N_41595);
nand U41860 (N_41860,N_41711,N_41724);
and U41861 (N_41861,N_41583,N_41624);
xor U41862 (N_41862,N_41734,N_41559);
nor U41863 (N_41863,N_41537,N_41654);
and U41864 (N_41864,N_41638,N_41676);
or U41865 (N_41865,N_41632,N_41685);
nor U41866 (N_41866,N_41539,N_41587);
nand U41867 (N_41867,N_41705,N_41611);
nand U41868 (N_41868,N_41547,N_41656);
and U41869 (N_41869,N_41633,N_41744);
nor U41870 (N_41870,N_41519,N_41591);
or U41871 (N_41871,N_41603,N_41540);
nand U41872 (N_41872,N_41604,N_41551);
nand U41873 (N_41873,N_41716,N_41621);
and U41874 (N_41874,N_41593,N_41660);
nor U41875 (N_41875,N_41664,N_41739);
nor U41876 (N_41876,N_41732,N_41701);
nand U41877 (N_41877,N_41548,N_41737);
nor U41878 (N_41878,N_41701,N_41665);
nand U41879 (N_41879,N_41610,N_41604);
and U41880 (N_41880,N_41705,N_41712);
xor U41881 (N_41881,N_41525,N_41706);
nand U41882 (N_41882,N_41718,N_41607);
or U41883 (N_41883,N_41735,N_41509);
and U41884 (N_41884,N_41703,N_41623);
or U41885 (N_41885,N_41672,N_41543);
and U41886 (N_41886,N_41601,N_41669);
nor U41887 (N_41887,N_41707,N_41638);
nand U41888 (N_41888,N_41630,N_41525);
nand U41889 (N_41889,N_41730,N_41625);
and U41890 (N_41890,N_41722,N_41562);
nand U41891 (N_41891,N_41691,N_41502);
and U41892 (N_41892,N_41623,N_41564);
nor U41893 (N_41893,N_41735,N_41622);
or U41894 (N_41894,N_41645,N_41716);
xnor U41895 (N_41895,N_41558,N_41596);
nor U41896 (N_41896,N_41686,N_41587);
or U41897 (N_41897,N_41586,N_41703);
and U41898 (N_41898,N_41673,N_41704);
nand U41899 (N_41899,N_41722,N_41526);
and U41900 (N_41900,N_41724,N_41732);
nand U41901 (N_41901,N_41612,N_41595);
and U41902 (N_41902,N_41633,N_41575);
and U41903 (N_41903,N_41708,N_41557);
nor U41904 (N_41904,N_41678,N_41675);
nand U41905 (N_41905,N_41522,N_41616);
xnor U41906 (N_41906,N_41650,N_41515);
and U41907 (N_41907,N_41667,N_41728);
nor U41908 (N_41908,N_41590,N_41660);
nand U41909 (N_41909,N_41647,N_41579);
or U41910 (N_41910,N_41693,N_41576);
nand U41911 (N_41911,N_41618,N_41644);
nor U41912 (N_41912,N_41747,N_41684);
xnor U41913 (N_41913,N_41709,N_41749);
and U41914 (N_41914,N_41586,N_41592);
xnor U41915 (N_41915,N_41547,N_41732);
nand U41916 (N_41916,N_41541,N_41708);
xnor U41917 (N_41917,N_41629,N_41748);
or U41918 (N_41918,N_41542,N_41748);
or U41919 (N_41919,N_41602,N_41509);
and U41920 (N_41920,N_41605,N_41550);
and U41921 (N_41921,N_41664,N_41506);
xnor U41922 (N_41922,N_41539,N_41739);
nor U41923 (N_41923,N_41646,N_41539);
xnor U41924 (N_41924,N_41569,N_41690);
or U41925 (N_41925,N_41531,N_41537);
nand U41926 (N_41926,N_41525,N_41567);
nor U41927 (N_41927,N_41533,N_41620);
nor U41928 (N_41928,N_41599,N_41550);
or U41929 (N_41929,N_41640,N_41641);
xor U41930 (N_41930,N_41737,N_41657);
nand U41931 (N_41931,N_41503,N_41683);
or U41932 (N_41932,N_41574,N_41730);
nor U41933 (N_41933,N_41726,N_41544);
xnor U41934 (N_41934,N_41700,N_41568);
xnor U41935 (N_41935,N_41588,N_41671);
xor U41936 (N_41936,N_41602,N_41549);
xnor U41937 (N_41937,N_41598,N_41611);
and U41938 (N_41938,N_41657,N_41605);
or U41939 (N_41939,N_41721,N_41612);
xor U41940 (N_41940,N_41691,N_41684);
nor U41941 (N_41941,N_41500,N_41516);
nor U41942 (N_41942,N_41746,N_41633);
nand U41943 (N_41943,N_41611,N_41559);
xor U41944 (N_41944,N_41637,N_41718);
or U41945 (N_41945,N_41546,N_41633);
and U41946 (N_41946,N_41550,N_41570);
and U41947 (N_41947,N_41547,N_41596);
nor U41948 (N_41948,N_41747,N_41555);
xnor U41949 (N_41949,N_41723,N_41532);
nor U41950 (N_41950,N_41530,N_41692);
nor U41951 (N_41951,N_41711,N_41607);
xnor U41952 (N_41952,N_41608,N_41662);
nor U41953 (N_41953,N_41601,N_41528);
nor U41954 (N_41954,N_41626,N_41578);
nor U41955 (N_41955,N_41630,N_41625);
and U41956 (N_41956,N_41678,N_41671);
nand U41957 (N_41957,N_41518,N_41675);
nor U41958 (N_41958,N_41623,N_41505);
nand U41959 (N_41959,N_41552,N_41582);
or U41960 (N_41960,N_41532,N_41625);
nand U41961 (N_41961,N_41641,N_41603);
nor U41962 (N_41962,N_41602,N_41543);
nand U41963 (N_41963,N_41732,N_41696);
nand U41964 (N_41964,N_41670,N_41739);
nand U41965 (N_41965,N_41654,N_41711);
and U41966 (N_41966,N_41642,N_41683);
or U41967 (N_41967,N_41550,N_41572);
or U41968 (N_41968,N_41509,N_41589);
or U41969 (N_41969,N_41559,N_41612);
nand U41970 (N_41970,N_41548,N_41542);
nor U41971 (N_41971,N_41545,N_41663);
nand U41972 (N_41972,N_41565,N_41537);
nor U41973 (N_41973,N_41630,N_41739);
nor U41974 (N_41974,N_41510,N_41670);
and U41975 (N_41975,N_41689,N_41588);
xor U41976 (N_41976,N_41659,N_41698);
and U41977 (N_41977,N_41713,N_41738);
nor U41978 (N_41978,N_41633,N_41624);
xor U41979 (N_41979,N_41579,N_41563);
nand U41980 (N_41980,N_41600,N_41578);
nand U41981 (N_41981,N_41679,N_41518);
or U41982 (N_41982,N_41657,N_41677);
or U41983 (N_41983,N_41540,N_41654);
or U41984 (N_41984,N_41655,N_41604);
xnor U41985 (N_41985,N_41570,N_41631);
nand U41986 (N_41986,N_41510,N_41743);
nand U41987 (N_41987,N_41738,N_41661);
nand U41988 (N_41988,N_41512,N_41736);
and U41989 (N_41989,N_41547,N_41634);
or U41990 (N_41990,N_41667,N_41555);
or U41991 (N_41991,N_41679,N_41741);
or U41992 (N_41992,N_41621,N_41503);
nand U41993 (N_41993,N_41514,N_41629);
xor U41994 (N_41994,N_41677,N_41710);
nand U41995 (N_41995,N_41525,N_41522);
nand U41996 (N_41996,N_41668,N_41523);
or U41997 (N_41997,N_41613,N_41721);
nand U41998 (N_41998,N_41585,N_41604);
nor U41999 (N_41999,N_41615,N_41565);
and U42000 (N_42000,N_41833,N_41761);
xor U42001 (N_42001,N_41880,N_41824);
and U42002 (N_42002,N_41940,N_41918);
or U42003 (N_42003,N_41827,N_41831);
and U42004 (N_42004,N_41976,N_41887);
or U42005 (N_42005,N_41960,N_41832);
nand U42006 (N_42006,N_41840,N_41790);
or U42007 (N_42007,N_41920,N_41900);
or U42008 (N_42008,N_41990,N_41971);
and U42009 (N_42009,N_41907,N_41891);
or U42010 (N_42010,N_41843,N_41966);
and U42011 (N_42011,N_41893,N_41859);
xnor U42012 (N_42012,N_41755,N_41888);
nor U42013 (N_42013,N_41818,N_41985);
nor U42014 (N_42014,N_41801,N_41965);
or U42015 (N_42015,N_41870,N_41879);
nor U42016 (N_42016,N_41961,N_41875);
nand U42017 (N_42017,N_41867,N_41871);
and U42018 (N_42018,N_41989,N_41792);
xor U42019 (N_42019,N_41922,N_41873);
and U42020 (N_42020,N_41781,N_41786);
xnor U42021 (N_42021,N_41980,N_41766);
nand U42022 (N_42022,N_41968,N_41860);
nor U42023 (N_42023,N_41890,N_41830);
or U42024 (N_42024,N_41881,N_41776);
nand U42025 (N_42025,N_41908,N_41858);
or U42026 (N_42026,N_41946,N_41914);
nand U42027 (N_42027,N_41779,N_41789);
nand U42028 (N_42028,N_41905,N_41934);
xnor U42029 (N_42029,N_41967,N_41864);
or U42030 (N_42030,N_41872,N_41901);
and U42031 (N_42031,N_41816,N_41984);
nand U42032 (N_42032,N_41760,N_41802);
nand U42033 (N_42033,N_41862,N_41983);
and U42034 (N_42034,N_41770,N_41812);
nand U42035 (N_42035,N_41787,N_41834);
and U42036 (N_42036,N_41993,N_41811);
xnor U42037 (N_42037,N_41931,N_41794);
and U42038 (N_42038,N_41958,N_41795);
xnor U42039 (N_42039,N_41951,N_41850);
xnor U42040 (N_42040,N_41895,N_41838);
and U42041 (N_42041,N_41884,N_41957);
or U42042 (N_42042,N_41911,N_41942);
xnor U42043 (N_42043,N_41977,N_41925);
nand U42044 (N_42044,N_41782,N_41857);
or U42045 (N_42045,N_41919,N_41823);
and U42046 (N_42046,N_41974,N_41944);
and U42047 (N_42047,N_41807,N_41963);
and U42048 (N_42048,N_41924,N_41927);
nand U42049 (N_42049,N_41756,N_41987);
nor U42050 (N_42050,N_41959,N_41866);
nand U42051 (N_42051,N_41762,N_41785);
nor U42052 (N_42052,N_41981,N_41798);
xnor U42053 (N_42053,N_41948,N_41771);
xnor U42054 (N_42054,N_41943,N_41751);
xor U42055 (N_42055,N_41998,N_41758);
nand U42056 (N_42056,N_41841,N_41869);
or U42057 (N_42057,N_41820,N_41986);
xnor U42058 (N_42058,N_41903,N_41842);
and U42059 (N_42059,N_41775,N_41906);
xor U42060 (N_42060,N_41883,N_41932);
nor U42061 (N_42061,N_41999,N_41910);
nand U42062 (N_42062,N_41791,N_41973);
nand U42063 (N_42063,N_41979,N_41757);
nor U42064 (N_42064,N_41803,N_41753);
nor U42065 (N_42065,N_41933,N_41952);
xnor U42066 (N_42066,N_41797,N_41897);
xnor U42067 (N_42067,N_41839,N_41904);
nand U42068 (N_42068,N_41926,N_41796);
and U42069 (N_42069,N_41975,N_41923);
and U42070 (N_42070,N_41784,N_41874);
and U42071 (N_42071,N_41750,N_41829);
nand U42072 (N_42072,N_41972,N_41815);
xor U42073 (N_42073,N_41821,N_41962);
or U42074 (N_42074,N_41765,N_41805);
nand U42075 (N_42075,N_41844,N_41778);
nor U42076 (N_42076,N_41854,N_41828);
or U42077 (N_42077,N_41767,N_41945);
nor U42078 (N_42078,N_41915,N_41892);
xnor U42079 (N_42079,N_41814,N_41941);
nand U42080 (N_42080,N_41947,N_41835);
nand U42081 (N_42081,N_41982,N_41970);
or U42082 (N_42082,N_41774,N_41938);
or U42083 (N_42083,N_41764,N_41817);
nand U42084 (N_42084,N_41936,N_41819);
and U42085 (N_42085,N_41885,N_41991);
xnor U42086 (N_42086,N_41769,N_41894);
nand U42087 (N_42087,N_41950,N_41878);
and U42088 (N_42088,N_41899,N_41988);
xnor U42089 (N_42089,N_41754,N_41955);
and U42090 (N_42090,N_41825,N_41909);
nor U42091 (N_42091,N_41772,N_41921);
nand U42092 (N_42092,N_41783,N_41916);
and U42093 (N_42093,N_41865,N_41763);
and U42094 (N_42094,N_41773,N_41759);
and U42095 (N_42095,N_41995,N_41954);
xor U42096 (N_42096,N_41929,N_41939);
or U42097 (N_42097,N_41836,N_41928);
nor U42098 (N_42098,N_41804,N_41996);
and U42099 (N_42099,N_41964,N_41902);
or U42100 (N_42100,N_41949,N_41809);
xor U42101 (N_42101,N_41777,N_41953);
nand U42102 (N_42102,N_41846,N_41806);
and U42103 (N_42103,N_41913,N_41793);
xnor U42104 (N_42104,N_41855,N_41800);
xor U42105 (N_42105,N_41861,N_41780);
or U42106 (N_42106,N_41912,N_41847);
xnor U42107 (N_42107,N_41810,N_41930);
nor U42108 (N_42108,N_41768,N_41845);
and U42109 (N_42109,N_41956,N_41853);
nand U42110 (N_42110,N_41978,N_41826);
or U42111 (N_42111,N_41886,N_41808);
and U42112 (N_42112,N_41849,N_41896);
or U42113 (N_42113,N_41889,N_41937);
nand U42114 (N_42114,N_41868,N_41994);
or U42115 (N_42115,N_41877,N_41837);
and U42116 (N_42116,N_41882,N_41852);
nand U42117 (N_42117,N_41876,N_41935);
or U42118 (N_42118,N_41898,N_41788);
and U42119 (N_42119,N_41856,N_41851);
nor U42120 (N_42120,N_41822,N_41917);
nand U42121 (N_42121,N_41969,N_41813);
nand U42122 (N_42122,N_41992,N_41848);
nor U42123 (N_42123,N_41997,N_41752);
and U42124 (N_42124,N_41799,N_41863);
nand U42125 (N_42125,N_41917,N_41773);
nor U42126 (N_42126,N_41751,N_41932);
nor U42127 (N_42127,N_41894,N_41942);
xnor U42128 (N_42128,N_41906,N_41997);
or U42129 (N_42129,N_41972,N_41896);
nor U42130 (N_42130,N_41962,N_41970);
nand U42131 (N_42131,N_41824,N_41757);
or U42132 (N_42132,N_41962,N_41802);
nor U42133 (N_42133,N_41757,N_41846);
and U42134 (N_42134,N_41916,N_41803);
and U42135 (N_42135,N_41931,N_41757);
nand U42136 (N_42136,N_41907,N_41906);
or U42137 (N_42137,N_41857,N_41833);
or U42138 (N_42138,N_41773,N_41777);
and U42139 (N_42139,N_41918,N_41901);
xor U42140 (N_42140,N_41802,N_41775);
xor U42141 (N_42141,N_41853,N_41827);
nand U42142 (N_42142,N_41792,N_41805);
or U42143 (N_42143,N_41860,N_41820);
and U42144 (N_42144,N_41935,N_41857);
or U42145 (N_42145,N_41986,N_41982);
nand U42146 (N_42146,N_41956,N_41862);
nand U42147 (N_42147,N_41868,N_41959);
or U42148 (N_42148,N_41878,N_41790);
and U42149 (N_42149,N_41812,N_41829);
and U42150 (N_42150,N_41938,N_41950);
or U42151 (N_42151,N_41895,N_41787);
nor U42152 (N_42152,N_41927,N_41815);
nand U42153 (N_42153,N_41777,N_41845);
or U42154 (N_42154,N_41791,N_41907);
nand U42155 (N_42155,N_41834,N_41753);
nand U42156 (N_42156,N_41920,N_41790);
nand U42157 (N_42157,N_41987,N_41979);
or U42158 (N_42158,N_41907,N_41806);
nor U42159 (N_42159,N_41932,N_41861);
nand U42160 (N_42160,N_41963,N_41974);
and U42161 (N_42161,N_41851,N_41877);
xnor U42162 (N_42162,N_41903,N_41870);
nand U42163 (N_42163,N_41824,N_41812);
and U42164 (N_42164,N_41941,N_41855);
nor U42165 (N_42165,N_41788,N_41832);
or U42166 (N_42166,N_41773,N_41874);
or U42167 (N_42167,N_41855,N_41774);
nor U42168 (N_42168,N_41877,N_41872);
xor U42169 (N_42169,N_41883,N_41969);
xor U42170 (N_42170,N_41865,N_41984);
xor U42171 (N_42171,N_41770,N_41855);
or U42172 (N_42172,N_41874,N_41980);
or U42173 (N_42173,N_41971,N_41977);
and U42174 (N_42174,N_41868,N_41865);
or U42175 (N_42175,N_41913,N_41843);
nand U42176 (N_42176,N_41948,N_41997);
and U42177 (N_42177,N_41929,N_41897);
or U42178 (N_42178,N_41869,N_41891);
nand U42179 (N_42179,N_41865,N_41968);
and U42180 (N_42180,N_41929,N_41806);
xor U42181 (N_42181,N_41884,N_41974);
nor U42182 (N_42182,N_41912,N_41763);
nand U42183 (N_42183,N_41856,N_41996);
nor U42184 (N_42184,N_41889,N_41785);
xnor U42185 (N_42185,N_41987,N_41764);
nor U42186 (N_42186,N_41834,N_41885);
or U42187 (N_42187,N_41877,N_41875);
nand U42188 (N_42188,N_41833,N_41829);
or U42189 (N_42189,N_41991,N_41960);
nand U42190 (N_42190,N_41753,N_41862);
nor U42191 (N_42191,N_41766,N_41934);
nor U42192 (N_42192,N_41893,N_41855);
nor U42193 (N_42193,N_41944,N_41864);
nor U42194 (N_42194,N_41832,N_41883);
and U42195 (N_42195,N_41990,N_41819);
or U42196 (N_42196,N_41972,N_41764);
xor U42197 (N_42197,N_41777,N_41800);
xnor U42198 (N_42198,N_41908,N_41826);
xor U42199 (N_42199,N_41778,N_41983);
and U42200 (N_42200,N_41896,N_41799);
xor U42201 (N_42201,N_41840,N_41920);
nor U42202 (N_42202,N_41951,N_41995);
xnor U42203 (N_42203,N_41867,N_41956);
and U42204 (N_42204,N_41881,N_41790);
and U42205 (N_42205,N_41797,N_41940);
and U42206 (N_42206,N_41839,N_41951);
nand U42207 (N_42207,N_41779,N_41923);
or U42208 (N_42208,N_41928,N_41967);
nor U42209 (N_42209,N_41805,N_41836);
nand U42210 (N_42210,N_41924,N_41871);
or U42211 (N_42211,N_41804,N_41912);
xor U42212 (N_42212,N_41765,N_41839);
nor U42213 (N_42213,N_41994,N_41761);
or U42214 (N_42214,N_41922,N_41768);
or U42215 (N_42215,N_41820,N_41922);
or U42216 (N_42216,N_41894,N_41908);
or U42217 (N_42217,N_41972,N_41763);
xnor U42218 (N_42218,N_41819,N_41754);
nand U42219 (N_42219,N_41946,N_41887);
and U42220 (N_42220,N_41894,N_41798);
nand U42221 (N_42221,N_41773,N_41965);
xor U42222 (N_42222,N_41759,N_41986);
nor U42223 (N_42223,N_41817,N_41827);
nor U42224 (N_42224,N_41927,N_41770);
nand U42225 (N_42225,N_41959,N_41898);
xor U42226 (N_42226,N_41781,N_41856);
and U42227 (N_42227,N_41806,N_41974);
xnor U42228 (N_42228,N_41889,N_41871);
or U42229 (N_42229,N_41847,N_41952);
and U42230 (N_42230,N_41903,N_41824);
or U42231 (N_42231,N_41913,N_41801);
nor U42232 (N_42232,N_41774,N_41977);
or U42233 (N_42233,N_41938,N_41784);
xor U42234 (N_42234,N_41796,N_41906);
xor U42235 (N_42235,N_41937,N_41950);
nor U42236 (N_42236,N_41926,N_41835);
and U42237 (N_42237,N_41857,N_41813);
and U42238 (N_42238,N_41845,N_41872);
xor U42239 (N_42239,N_41892,N_41919);
or U42240 (N_42240,N_41844,N_41810);
xnor U42241 (N_42241,N_41901,N_41882);
xnor U42242 (N_42242,N_41856,N_41774);
nand U42243 (N_42243,N_41816,N_41993);
xor U42244 (N_42244,N_41932,N_41914);
and U42245 (N_42245,N_41936,N_41924);
xnor U42246 (N_42246,N_41944,N_41792);
or U42247 (N_42247,N_41966,N_41880);
nor U42248 (N_42248,N_41799,N_41814);
xor U42249 (N_42249,N_41856,N_41820);
nand U42250 (N_42250,N_42198,N_42084);
or U42251 (N_42251,N_42200,N_42211);
nor U42252 (N_42252,N_42229,N_42079);
and U42253 (N_42253,N_42156,N_42096);
or U42254 (N_42254,N_42159,N_42125);
nor U42255 (N_42255,N_42134,N_42145);
xor U42256 (N_42256,N_42165,N_42107);
xnor U42257 (N_42257,N_42246,N_42009);
nand U42258 (N_42258,N_42204,N_42228);
nand U42259 (N_42259,N_42213,N_42036);
and U42260 (N_42260,N_42160,N_42183);
or U42261 (N_42261,N_42238,N_42008);
and U42262 (N_42262,N_42090,N_42112);
nor U42263 (N_42263,N_42053,N_42061);
or U42264 (N_42264,N_42066,N_42173);
xor U42265 (N_42265,N_42216,N_42058);
nor U42266 (N_42266,N_42197,N_42064);
xor U42267 (N_42267,N_42138,N_42062);
and U42268 (N_42268,N_42052,N_42056);
nand U42269 (N_42269,N_42194,N_42143);
or U42270 (N_42270,N_42024,N_42039);
and U42271 (N_42271,N_42076,N_42214);
xor U42272 (N_42272,N_42130,N_42093);
and U42273 (N_42273,N_42069,N_42167);
nand U42274 (N_42274,N_42025,N_42007);
nand U42275 (N_42275,N_42043,N_42029);
and U42276 (N_42276,N_42203,N_42181);
nand U42277 (N_42277,N_42120,N_42179);
and U42278 (N_42278,N_42004,N_42201);
or U42279 (N_42279,N_42136,N_42026);
xnor U42280 (N_42280,N_42182,N_42234);
nor U42281 (N_42281,N_42158,N_42142);
and U42282 (N_42282,N_42241,N_42117);
nor U42283 (N_42283,N_42144,N_42176);
or U42284 (N_42284,N_42018,N_42155);
or U42285 (N_42285,N_42190,N_42154);
or U42286 (N_42286,N_42087,N_42209);
nand U42287 (N_42287,N_42038,N_42129);
and U42288 (N_42288,N_42016,N_42085);
xnor U42289 (N_42289,N_42041,N_42010);
nor U42290 (N_42290,N_42207,N_42098);
or U42291 (N_42291,N_42175,N_42146);
xnor U42292 (N_42292,N_42195,N_42172);
nand U42293 (N_42293,N_42170,N_42192);
xnor U42294 (N_42294,N_42242,N_42070);
and U42295 (N_42295,N_42180,N_42001);
nand U42296 (N_42296,N_42219,N_42071);
or U42297 (N_42297,N_42208,N_42051);
nand U42298 (N_42298,N_42037,N_42121);
or U42299 (N_42299,N_42082,N_42030);
xor U42300 (N_42300,N_42050,N_42011);
xor U42301 (N_42301,N_42106,N_42065);
xnor U42302 (N_42302,N_42149,N_42123);
xnor U42303 (N_42303,N_42196,N_42225);
and U42304 (N_42304,N_42021,N_42217);
nand U42305 (N_42305,N_42000,N_42083);
and U42306 (N_42306,N_42248,N_42060);
and U42307 (N_42307,N_42028,N_42072);
xnor U42308 (N_42308,N_42063,N_42247);
xor U42309 (N_42309,N_42014,N_42151);
nor U42310 (N_42310,N_42086,N_42091);
nor U42311 (N_42311,N_42218,N_42013);
and U42312 (N_42312,N_42105,N_42095);
nor U42313 (N_42313,N_42224,N_42193);
and U42314 (N_42314,N_42178,N_42075);
xor U42315 (N_42315,N_42152,N_42057);
nor U42316 (N_42316,N_42045,N_42137);
xnor U42317 (N_42317,N_42124,N_42177);
xnor U42318 (N_42318,N_42141,N_42080);
xnor U42319 (N_42319,N_42059,N_42113);
nand U42320 (N_42320,N_42102,N_42027);
nand U42321 (N_42321,N_42118,N_42081);
or U42322 (N_42322,N_42103,N_42020);
nand U42323 (N_42323,N_42088,N_42089);
and U42324 (N_42324,N_42068,N_42115);
xnor U42325 (N_42325,N_42168,N_42153);
nand U42326 (N_42326,N_42185,N_42135);
or U42327 (N_42327,N_42017,N_42223);
xnor U42328 (N_42328,N_42131,N_42157);
nand U42329 (N_42329,N_42139,N_42077);
xnor U42330 (N_42330,N_42171,N_42033);
nor U42331 (N_42331,N_42235,N_42169);
xor U42332 (N_42332,N_42127,N_42005);
nand U42333 (N_42333,N_42122,N_42140);
xnor U42334 (N_42334,N_42236,N_42015);
xnor U42335 (N_42335,N_42116,N_42163);
xor U42336 (N_42336,N_42003,N_42249);
nand U42337 (N_42337,N_42230,N_42002);
or U42338 (N_42338,N_42092,N_42101);
and U42339 (N_42339,N_42222,N_42100);
or U42340 (N_42340,N_42109,N_42162);
and U42341 (N_42341,N_42023,N_42094);
nor U42342 (N_42342,N_42110,N_42232);
nor U42343 (N_42343,N_42074,N_42184);
or U42344 (N_42344,N_42047,N_42220);
xor U42345 (N_42345,N_42243,N_42244);
and U42346 (N_42346,N_42233,N_42191);
and U42347 (N_42347,N_42187,N_42245);
and U42348 (N_42348,N_42126,N_42111);
and U42349 (N_42349,N_42231,N_42221);
and U42350 (N_42350,N_42148,N_42227);
nand U42351 (N_42351,N_42044,N_42032);
nand U42352 (N_42352,N_42166,N_42202);
and U42353 (N_42353,N_42054,N_42239);
nor U42354 (N_42354,N_42040,N_42205);
or U42355 (N_42355,N_42199,N_42073);
nor U42356 (N_42356,N_42161,N_42189);
and U42357 (N_42357,N_42150,N_42035);
nor U42358 (N_42358,N_42237,N_42164);
nor U42359 (N_42359,N_42210,N_42078);
or U42360 (N_42360,N_42186,N_42006);
and U42361 (N_42361,N_42108,N_42215);
and U42362 (N_42362,N_42133,N_42188);
and U42363 (N_42363,N_42049,N_42132);
nor U42364 (N_42364,N_42067,N_42104);
nand U42365 (N_42365,N_42055,N_42099);
nand U42366 (N_42366,N_42226,N_42012);
xor U42367 (N_42367,N_42114,N_42128);
xnor U42368 (N_42368,N_42147,N_42019);
nand U42369 (N_42369,N_42046,N_42119);
nor U42370 (N_42370,N_42048,N_42206);
nor U42371 (N_42371,N_42212,N_42034);
or U42372 (N_42372,N_42042,N_42022);
xnor U42373 (N_42373,N_42174,N_42097);
nor U42374 (N_42374,N_42031,N_42240);
nand U42375 (N_42375,N_42118,N_42153);
nand U42376 (N_42376,N_42155,N_42029);
nor U42377 (N_42377,N_42001,N_42150);
nor U42378 (N_42378,N_42186,N_42228);
nand U42379 (N_42379,N_42083,N_42202);
and U42380 (N_42380,N_42001,N_42229);
nor U42381 (N_42381,N_42123,N_42033);
nand U42382 (N_42382,N_42047,N_42175);
nand U42383 (N_42383,N_42069,N_42117);
nand U42384 (N_42384,N_42124,N_42239);
or U42385 (N_42385,N_42072,N_42185);
nor U42386 (N_42386,N_42195,N_42078);
nor U42387 (N_42387,N_42126,N_42099);
and U42388 (N_42388,N_42066,N_42229);
and U42389 (N_42389,N_42023,N_42015);
xor U42390 (N_42390,N_42217,N_42166);
nand U42391 (N_42391,N_42090,N_42092);
nand U42392 (N_42392,N_42070,N_42058);
nor U42393 (N_42393,N_42030,N_42002);
nor U42394 (N_42394,N_42085,N_42132);
or U42395 (N_42395,N_42205,N_42057);
nor U42396 (N_42396,N_42130,N_42135);
nand U42397 (N_42397,N_42121,N_42056);
xnor U42398 (N_42398,N_42239,N_42213);
xor U42399 (N_42399,N_42170,N_42040);
xnor U42400 (N_42400,N_42021,N_42191);
nand U42401 (N_42401,N_42233,N_42213);
nand U42402 (N_42402,N_42202,N_42017);
nand U42403 (N_42403,N_42207,N_42236);
nand U42404 (N_42404,N_42240,N_42044);
nor U42405 (N_42405,N_42042,N_42086);
and U42406 (N_42406,N_42231,N_42193);
nand U42407 (N_42407,N_42079,N_42190);
nor U42408 (N_42408,N_42136,N_42116);
nor U42409 (N_42409,N_42191,N_42105);
nor U42410 (N_42410,N_42006,N_42099);
xor U42411 (N_42411,N_42018,N_42180);
nor U42412 (N_42412,N_42052,N_42181);
nand U42413 (N_42413,N_42141,N_42162);
nand U42414 (N_42414,N_42012,N_42229);
nand U42415 (N_42415,N_42031,N_42036);
xnor U42416 (N_42416,N_42186,N_42234);
or U42417 (N_42417,N_42229,N_42097);
xnor U42418 (N_42418,N_42235,N_42118);
xnor U42419 (N_42419,N_42154,N_42034);
nor U42420 (N_42420,N_42234,N_42228);
xnor U42421 (N_42421,N_42013,N_42100);
or U42422 (N_42422,N_42196,N_42137);
and U42423 (N_42423,N_42112,N_42145);
and U42424 (N_42424,N_42041,N_42166);
nand U42425 (N_42425,N_42155,N_42160);
xnor U42426 (N_42426,N_42222,N_42035);
nor U42427 (N_42427,N_42067,N_42234);
nor U42428 (N_42428,N_42038,N_42050);
nand U42429 (N_42429,N_42186,N_42080);
nand U42430 (N_42430,N_42053,N_42140);
xnor U42431 (N_42431,N_42092,N_42034);
xor U42432 (N_42432,N_42154,N_42159);
nand U42433 (N_42433,N_42087,N_42167);
or U42434 (N_42434,N_42137,N_42239);
or U42435 (N_42435,N_42055,N_42227);
xnor U42436 (N_42436,N_42032,N_42025);
nor U42437 (N_42437,N_42032,N_42020);
xnor U42438 (N_42438,N_42122,N_42094);
or U42439 (N_42439,N_42185,N_42142);
xor U42440 (N_42440,N_42230,N_42075);
and U42441 (N_42441,N_42074,N_42153);
nor U42442 (N_42442,N_42123,N_42023);
and U42443 (N_42443,N_42231,N_42173);
and U42444 (N_42444,N_42079,N_42129);
nor U42445 (N_42445,N_42139,N_42212);
nand U42446 (N_42446,N_42092,N_42028);
or U42447 (N_42447,N_42096,N_42135);
and U42448 (N_42448,N_42061,N_42033);
or U42449 (N_42449,N_42071,N_42014);
or U42450 (N_42450,N_42003,N_42080);
or U42451 (N_42451,N_42046,N_42141);
or U42452 (N_42452,N_42057,N_42162);
or U42453 (N_42453,N_42197,N_42030);
or U42454 (N_42454,N_42174,N_42247);
nor U42455 (N_42455,N_42003,N_42014);
xor U42456 (N_42456,N_42148,N_42063);
xor U42457 (N_42457,N_42002,N_42105);
or U42458 (N_42458,N_42013,N_42112);
nor U42459 (N_42459,N_42165,N_42244);
or U42460 (N_42460,N_42121,N_42067);
and U42461 (N_42461,N_42133,N_42031);
and U42462 (N_42462,N_42044,N_42051);
nand U42463 (N_42463,N_42170,N_42183);
nand U42464 (N_42464,N_42240,N_42146);
nor U42465 (N_42465,N_42162,N_42220);
xnor U42466 (N_42466,N_42121,N_42155);
nor U42467 (N_42467,N_42072,N_42012);
nand U42468 (N_42468,N_42028,N_42246);
or U42469 (N_42469,N_42031,N_42055);
xor U42470 (N_42470,N_42167,N_42045);
or U42471 (N_42471,N_42171,N_42139);
and U42472 (N_42472,N_42006,N_42108);
xor U42473 (N_42473,N_42102,N_42160);
and U42474 (N_42474,N_42144,N_42119);
nor U42475 (N_42475,N_42088,N_42086);
nor U42476 (N_42476,N_42230,N_42159);
nand U42477 (N_42477,N_42103,N_42229);
nand U42478 (N_42478,N_42220,N_42118);
and U42479 (N_42479,N_42180,N_42063);
or U42480 (N_42480,N_42101,N_42236);
nor U42481 (N_42481,N_42082,N_42216);
xor U42482 (N_42482,N_42141,N_42000);
nor U42483 (N_42483,N_42100,N_42043);
or U42484 (N_42484,N_42076,N_42050);
xnor U42485 (N_42485,N_42051,N_42242);
nand U42486 (N_42486,N_42056,N_42243);
or U42487 (N_42487,N_42230,N_42173);
and U42488 (N_42488,N_42086,N_42241);
or U42489 (N_42489,N_42121,N_42185);
nand U42490 (N_42490,N_42213,N_42175);
nor U42491 (N_42491,N_42043,N_42057);
nor U42492 (N_42492,N_42002,N_42022);
xnor U42493 (N_42493,N_42063,N_42109);
xnor U42494 (N_42494,N_42091,N_42065);
nor U42495 (N_42495,N_42051,N_42073);
or U42496 (N_42496,N_42101,N_42114);
or U42497 (N_42497,N_42249,N_42223);
and U42498 (N_42498,N_42016,N_42089);
nor U42499 (N_42499,N_42002,N_42073);
nand U42500 (N_42500,N_42279,N_42269);
xor U42501 (N_42501,N_42340,N_42286);
nor U42502 (N_42502,N_42478,N_42425);
and U42503 (N_42503,N_42285,N_42332);
xor U42504 (N_42504,N_42380,N_42392);
or U42505 (N_42505,N_42367,N_42295);
nor U42506 (N_42506,N_42453,N_42433);
nand U42507 (N_42507,N_42360,N_42293);
xnor U42508 (N_42508,N_42282,N_42485);
nand U42509 (N_42509,N_42298,N_42251);
nand U42510 (N_42510,N_42297,N_42307);
xor U42511 (N_42511,N_42371,N_42264);
and U42512 (N_42512,N_42377,N_42400);
and U42513 (N_42513,N_42494,N_42475);
and U42514 (N_42514,N_42443,N_42361);
nor U42515 (N_42515,N_42404,N_42407);
nor U42516 (N_42516,N_42335,N_42312);
or U42517 (N_42517,N_42257,N_42368);
or U42518 (N_42518,N_42468,N_42353);
nor U42519 (N_42519,N_42271,N_42393);
or U42520 (N_42520,N_42397,N_42351);
and U42521 (N_42521,N_42499,N_42266);
xor U42522 (N_42522,N_42341,N_42262);
xor U42523 (N_42523,N_42369,N_42418);
or U42524 (N_42524,N_42398,N_42473);
and U42525 (N_42525,N_42394,N_42436);
xnor U42526 (N_42526,N_42465,N_42291);
or U42527 (N_42527,N_42490,N_42336);
and U42528 (N_42528,N_42489,N_42480);
xnor U42529 (N_42529,N_42402,N_42464);
or U42530 (N_42530,N_42498,N_42421);
and U42531 (N_42531,N_42313,N_42409);
xor U42532 (N_42532,N_42370,N_42469);
and U42533 (N_42533,N_42319,N_42310);
nor U42534 (N_42534,N_42429,N_42456);
or U42535 (N_42535,N_42482,N_42449);
nor U42536 (N_42536,N_42350,N_42386);
or U42537 (N_42537,N_42303,N_42455);
xnor U42538 (N_42538,N_42428,N_42322);
nand U42539 (N_42539,N_42497,N_42403);
or U42540 (N_42540,N_42388,N_42261);
and U42541 (N_42541,N_42381,N_42311);
nand U42542 (N_42542,N_42284,N_42444);
or U42543 (N_42543,N_42256,N_42346);
and U42544 (N_42544,N_42253,N_42294);
nor U42545 (N_42545,N_42434,N_42445);
xnor U42546 (N_42546,N_42383,N_42334);
nand U42547 (N_42547,N_42389,N_42347);
and U42548 (N_42548,N_42304,N_42470);
nor U42549 (N_42549,N_42488,N_42454);
xnor U42550 (N_42550,N_42385,N_42439);
or U42551 (N_42551,N_42375,N_42265);
or U42552 (N_42552,N_42450,N_42337);
nor U42553 (N_42553,N_42276,N_42323);
xnor U42554 (N_42554,N_42345,N_42376);
nand U42555 (N_42555,N_42273,N_42280);
xnor U42556 (N_42556,N_42440,N_42315);
xor U42557 (N_42557,N_42474,N_42476);
and U42558 (N_42558,N_42274,N_42382);
or U42559 (N_42559,N_42372,N_42270);
or U42560 (N_42560,N_42272,N_42320);
xor U42561 (N_42561,N_42493,N_42447);
or U42562 (N_42562,N_42331,N_42462);
xor U42563 (N_42563,N_42481,N_42422);
nand U42564 (N_42564,N_42329,N_42487);
nand U42565 (N_42565,N_42365,N_42305);
or U42566 (N_42566,N_42352,N_42472);
xnor U42567 (N_42567,N_42354,N_42259);
xor U42568 (N_42568,N_42484,N_42399);
nor U42569 (N_42569,N_42491,N_42287);
and U42570 (N_42570,N_42301,N_42258);
or U42571 (N_42571,N_42441,N_42255);
and U42572 (N_42572,N_42486,N_42314);
nor U42573 (N_42573,N_42451,N_42395);
or U42574 (N_42574,N_42326,N_42359);
nand U42575 (N_42575,N_42357,N_42289);
xnor U42576 (N_42576,N_42325,N_42281);
and U42577 (N_42577,N_42415,N_42495);
and U42578 (N_42578,N_42417,N_42288);
and U42579 (N_42579,N_42316,N_42327);
and U42580 (N_42580,N_42349,N_42308);
nand U42581 (N_42581,N_42254,N_42467);
and U42582 (N_42582,N_42411,N_42379);
nor U42583 (N_42583,N_42330,N_42408);
nand U42584 (N_42584,N_42448,N_42356);
xor U42585 (N_42585,N_42460,N_42466);
nor U42586 (N_42586,N_42390,N_42426);
and U42587 (N_42587,N_42463,N_42496);
nand U42588 (N_42588,N_42406,N_42452);
nand U42589 (N_42589,N_42416,N_42405);
or U42590 (N_42590,N_42435,N_42283);
or U42591 (N_42591,N_42355,N_42260);
nor U42592 (N_42592,N_42492,N_42431);
and U42593 (N_42593,N_42424,N_42401);
nand U42594 (N_42594,N_42414,N_42339);
and U42595 (N_42595,N_42343,N_42396);
or U42596 (N_42596,N_42364,N_42438);
and U42597 (N_42597,N_42328,N_42479);
nand U42598 (N_42598,N_42344,N_42446);
and U42599 (N_42599,N_42423,N_42292);
nand U42600 (N_42600,N_42362,N_42317);
xor U42601 (N_42601,N_42442,N_42309);
nand U42602 (N_42602,N_42324,N_42358);
or U42603 (N_42603,N_42373,N_42296);
nor U42604 (N_42604,N_42277,N_42457);
xnor U42605 (N_42605,N_42366,N_42413);
nor U42606 (N_42606,N_42302,N_42267);
or U42607 (N_42607,N_42477,N_42459);
xnor U42608 (N_42608,N_42348,N_42275);
nor U42609 (N_42609,N_42471,N_42321);
xnor U42610 (N_42610,N_42458,N_42461);
nand U42611 (N_42611,N_42342,N_42263);
nor U42612 (N_42612,N_42430,N_42427);
nand U42613 (N_42613,N_42278,N_42378);
nand U42614 (N_42614,N_42290,N_42384);
nand U42615 (N_42615,N_42410,N_42437);
and U42616 (N_42616,N_42387,N_42432);
and U42617 (N_42617,N_42374,N_42300);
xor U42618 (N_42618,N_42420,N_42268);
nand U42619 (N_42619,N_42363,N_42419);
or U42620 (N_42620,N_42391,N_42338);
nand U42621 (N_42621,N_42483,N_42299);
nor U42622 (N_42622,N_42412,N_42333);
xor U42623 (N_42623,N_42306,N_42318);
nor U42624 (N_42624,N_42252,N_42250);
nor U42625 (N_42625,N_42429,N_42398);
nand U42626 (N_42626,N_42380,N_42269);
nor U42627 (N_42627,N_42257,N_42468);
and U42628 (N_42628,N_42428,N_42309);
and U42629 (N_42629,N_42469,N_42495);
xor U42630 (N_42630,N_42426,N_42317);
xnor U42631 (N_42631,N_42265,N_42352);
xnor U42632 (N_42632,N_42428,N_42275);
or U42633 (N_42633,N_42454,N_42343);
nor U42634 (N_42634,N_42304,N_42320);
and U42635 (N_42635,N_42398,N_42378);
nor U42636 (N_42636,N_42251,N_42399);
nand U42637 (N_42637,N_42466,N_42344);
and U42638 (N_42638,N_42455,N_42285);
and U42639 (N_42639,N_42418,N_42268);
nand U42640 (N_42640,N_42486,N_42266);
xor U42641 (N_42641,N_42328,N_42347);
and U42642 (N_42642,N_42444,N_42469);
or U42643 (N_42643,N_42331,N_42383);
xor U42644 (N_42644,N_42264,N_42254);
nand U42645 (N_42645,N_42421,N_42295);
xor U42646 (N_42646,N_42468,N_42384);
or U42647 (N_42647,N_42373,N_42457);
or U42648 (N_42648,N_42324,N_42306);
and U42649 (N_42649,N_42277,N_42285);
nand U42650 (N_42650,N_42358,N_42417);
nor U42651 (N_42651,N_42336,N_42381);
nor U42652 (N_42652,N_42394,N_42402);
nand U42653 (N_42653,N_42462,N_42425);
and U42654 (N_42654,N_42330,N_42419);
xor U42655 (N_42655,N_42345,N_42407);
nand U42656 (N_42656,N_42389,N_42349);
or U42657 (N_42657,N_42289,N_42406);
or U42658 (N_42658,N_42339,N_42286);
nand U42659 (N_42659,N_42356,N_42390);
or U42660 (N_42660,N_42348,N_42283);
or U42661 (N_42661,N_42336,N_42279);
or U42662 (N_42662,N_42324,N_42316);
and U42663 (N_42663,N_42485,N_42479);
or U42664 (N_42664,N_42404,N_42454);
and U42665 (N_42665,N_42293,N_42409);
or U42666 (N_42666,N_42473,N_42256);
xnor U42667 (N_42667,N_42483,N_42381);
nand U42668 (N_42668,N_42344,N_42418);
and U42669 (N_42669,N_42471,N_42333);
or U42670 (N_42670,N_42331,N_42389);
nor U42671 (N_42671,N_42305,N_42326);
or U42672 (N_42672,N_42425,N_42330);
or U42673 (N_42673,N_42396,N_42436);
nand U42674 (N_42674,N_42476,N_42493);
nand U42675 (N_42675,N_42255,N_42451);
nor U42676 (N_42676,N_42265,N_42336);
nand U42677 (N_42677,N_42287,N_42424);
nor U42678 (N_42678,N_42371,N_42426);
and U42679 (N_42679,N_42448,N_42371);
or U42680 (N_42680,N_42361,N_42295);
xnor U42681 (N_42681,N_42255,N_42426);
xor U42682 (N_42682,N_42456,N_42361);
or U42683 (N_42683,N_42319,N_42439);
nor U42684 (N_42684,N_42384,N_42252);
nor U42685 (N_42685,N_42309,N_42324);
or U42686 (N_42686,N_42467,N_42437);
and U42687 (N_42687,N_42319,N_42296);
nor U42688 (N_42688,N_42442,N_42413);
nor U42689 (N_42689,N_42432,N_42494);
or U42690 (N_42690,N_42251,N_42448);
or U42691 (N_42691,N_42345,N_42296);
and U42692 (N_42692,N_42399,N_42394);
nor U42693 (N_42693,N_42375,N_42423);
or U42694 (N_42694,N_42412,N_42336);
xor U42695 (N_42695,N_42478,N_42296);
or U42696 (N_42696,N_42305,N_42399);
or U42697 (N_42697,N_42391,N_42354);
nand U42698 (N_42698,N_42262,N_42427);
xor U42699 (N_42699,N_42323,N_42352);
nor U42700 (N_42700,N_42350,N_42352);
or U42701 (N_42701,N_42330,N_42477);
xor U42702 (N_42702,N_42429,N_42454);
and U42703 (N_42703,N_42253,N_42465);
or U42704 (N_42704,N_42368,N_42450);
and U42705 (N_42705,N_42357,N_42312);
or U42706 (N_42706,N_42474,N_42407);
nor U42707 (N_42707,N_42261,N_42329);
nor U42708 (N_42708,N_42268,N_42453);
nor U42709 (N_42709,N_42416,N_42309);
or U42710 (N_42710,N_42336,N_42296);
and U42711 (N_42711,N_42328,N_42471);
and U42712 (N_42712,N_42362,N_42462);
xnor U42713 (N_42713,N_42335,N_42437);
nor U42714 (N_42714,N_42382,N_42339);
nor U42715 (N_42715,N_42437,N_42395);
nor U42716 (N_42716,N_42365,N_42492);
xor U42717 (N_42717,N_42312,N_42402);
xor U42718 (N_42718,N_42408,N_42363);
or U42719 (N_42719,N_42440,N_42441);
or U42720 (N_42720,N_42259,N_42394);
and U42721 (N_42721,N_42457,N_42427);
nor U42722 (N_42722,N_42312,N_42406);
xnor U42723 (N_42723,N_42297,N_42337);
nor U42724 (N_42724,N_42325,N_42373);
or U42725 (N_42725,N_42442,N_42429);
nor U42726 (N_42726,N_42434,N_42376);
nand U42727 (N_42727,N_42458,N_42311);
nor U42728 (N_42728,N_42376,N_42328);
or U42729 (N_42729,N_42499,N_42272);
xor U42730 (N_42730,N_42466,N_42453);
nor U42731 (N_42731,N_42437,N_42289);
nor U42732 (N_42732,N_42416,N_42323);
or U42733 (N_42733,N_42308,N_42310);
nor U42734 (N_42734,N_42429,N_42394);
nand U42735 (N_42735,N_42317,N_42343);
or U42736 (N_42736,N_42393,N_42325);
or U42737 (N_42737,N_42456,N_42330);
nor U42738 (N_42738,N_42425,N_42312);
xor U42739 (N_42739,N_42425,N_42372);
xor U42740 (N_42740,N_42401,N_42493);
xnor U42741 (N_42741,N_42260,N_42393);
nand U42742 (N_42742,N_42281,N_42349);
and U42743 (N_42743,N_42341,N_42346);
xnor U42744 (N_42744,N_42316,N_42404);
nand U42745 (N_42745,N_42434,N_42279);
nor U42746 (N_42746,N_42351,N_42364);
and U42747 (N_42747,N_42260,N_42343);
or U42748 (N_42748,N_42378,N_42291);
or U42749 (N_42749,N_42477,N_42419);
or U42750 (N_42750,N_42667,N_42744);
nand U42751 (N_42751,N_42612,N_42504);
nand U42752 (N_42752,N_42657,N_42737);
nor U42753 (N_42753,N_42548,N_42546);
nor U42754 (N_42754,N_42526,N_42694);
and U42755 (N_42755,N_42528,N_42601);
or U42756 (N_42756,N_42530,N_42693);
nor U42757 (N_42757,N_42571,N_42676);
and U42758 (N_42758,N_42592,N_42642);
nand U42759 (N_42759,N_42649,N_42515);
or U42760 (N_42760,N_42525,N_42552);
nor U42761 (N_42761,N_42691,N_42585);
nand U42762 (N_42762,N_42729,N_42644);
nand U42763 (N_42763,N_42618,N_42578);
nand U42764 (N_42764,N_42554,N_42653);
nor U42765 (N_42765,N_42576,N_42698);
and U42766 (N_42766,N_42595,N_42710);
or U42767 (N_42767,N_42619,N_42568);
or U42768 (N_42768,N_42725,N_42678);
xnor U42769 (N_42769,N_42715,N_42641);
nand U42770 (N_42770,N_42722,N_42703);
xor U42771 (N_42771,N_42610,N_42524);
and U42772 (N_42772,N_42536,N_42719);
nand U42773 (N_42773,N_42532,N_42549);
and U42774 (N_42774,N_42531,N_42599);
nand U42775 (N_42775,N_42579,N_42664);
nor U42776 (N_42776,N_42740,N_42523);
nor U42777 (N_42777,N_42519,N_42735);
xor U42778 (N_42778,N_42604,N_42606);
nand U42779 (N_42779,N_42645,N_42603);
or U42780 (N_42780,N_42590,N_42724);
or U42781 (N_42781,N_42584,N_42608);
nand U42782 (N_42782,N_42656,N_42638);
xor U42783 (N_42783,N_42630,N_42516);
and U42784 (N_42784,N_42743,N_42747);
nand U42785 (N_42785,N_42648,N_42632);
xnor U42786 (N_42786,N_42502,N_42701);
nand U42787 (N_42787,N_42637,N_42570);
nand U42788 (N_42788,N_42511,N_42721);
xor U42789 (N_42789,N_42687,N_42503);
and U42790 (N_42790,N_42541,N_42643);
xor U42791 (N_42791,N_42628,N_42688);
or U42792 (N_42792,N_42707,N_42651);
nand U42793 (N_42793,N_42586,N_42500);
or U42794 (N_42794,N_42537,N_42544);
nor U42795 (N_42795,N_42646,N_42673);
nor U42796 (N_42796,N_42535,N_42711);
or U42797 (N_42797,N_42666,N_42605);
and U42798 (N_42798,N_42509,N_42663);
and U42799 (N_42799,N_42633,N_42654);
xnor U42800 (N_42800,N_42668,N_42501);
nand U42801 (N_42801,N_42695,N_42561);
nor U42802 (N_42802,N_42510,N_42506);
nand U42803 (N_42803,N_42679,N_42686);
nand U42804 (N_42804,N_42683,N_42508);
xnor U42805 (N_42805,N_42738,N_42527);
or U42806 (N_42806,N_42690,N_42672);
or U42807 (N_42807,N_42702,N_42569);
and U42808 (N_42808,N_42700,N_42681);
or U42809 (N_42809,N_42658,N_42514);
nor U42810 (N_42810,N_42682,N_42680);
nor U42811 (N_42811,N_42538,N_42505);
nor U42812 (N_42812,N_42594,N_42611);
and U42813 (N_42813,N_42709,N_42621);
or U42814 (N_42814,N_42613,N_42674);
or U42815 (N_42815,N_42718,N_42669);
xnor U42816 (N_42816,N_42749,N_42671);
and U42817 (N_42817,N_42574,N_42615);
nor U42818 (N_42818,N_42627,N_42728);
xor U42819 (N_42819,N_42575,N_42635);
nand U42820 (N_42820,N_42513,N_42677);
and U42821 (N_42821,N_42727,N_42731);
and U42822 (N_42822,N_42588,N_42675);
and U42823 (N_42823,N_42597,N_42733);
xor U42824 (N_42824,N_42726,N_42614);
nor U42825 (N_42825,N_42716,N_42563);
xnor U42826 (N_42826,N_42547,N_42662);
nand U42827 (N_42827,N_42684,N_42553);
nor U42828 (N_42828,N_42562,N_42580);
and U42829 (N_42829,N_42564,N_42634);
nor U42830 (N_42830,N_42607,N_42636);
or U42831 (N_42831,N_42732,N_42520);
xor U42832 (N_42832,N_42631,N_42739);
xnor U42833 (N_42833,N_42652,N_42730);
xor U42834 (N_42834,N_42577,N_42540);
nand U42835 (N_42835,N_42745,N_42624);
or U42836 (N_42836,N_42589,N_42512);
or U42837 (N_42837,N_42567,N_42661);
nor U42838 (N_42838,N_42581,N_42660);
nand U42839 (N_42839,N_42622,N_42556);
nand U42840 (N_42840,N_42517,N_42625);
nand U42841 (N_42841,N_42543,N_42717);
xor U42842 (N_42842,N_42640,N_42723);
or U42843 (N_42843,N_42697,N_42551);
or U42844 (N_42844,N_42655,N_42529);
nor U42845 (N_42845,N_42713,N_42692);
nor U42846 (N_42846,N_42629,N_42602);
nand U42847 (N_42847,N_42720,N_42598);
or U42848 (N_42848,N_42689,N_42734);
or U42849 (N_42849,N_42708,N_42696);
and U42850 (N_42850,N_42600,N_42558);
nor U42851 (N_42851,N_42573,N_42566);
xnor U42852 (N_42852,N_42704,N_42557);
xnor U42853 (N_42853,N_42587,N_42714);
and U42854 (N_42854,N_42522,N_42670);
and U42855 (N_42855,N_42736,N_42593);
nor U42856 (N_42856,N_42623,N_42539);
and U42857 (N_42857,N_42659,N_42705);
nand U42858 (N_42858,N_42560,N_42706);
and U42859 (N_42859,N_42533,N_42565);
or U42860 (N_42860,N_42582,N_42685);
xnor U42861 (N_42861,N_42555,N_42699);
nor U42862 (N_42862,N_42521,N_42559);
xor U42863 (N_42863,N_42518,N_42741);
nor U42864 (N_42864,N_42617,N_42550);
nand U42865 (N_42865,N_42620,N_42591);
and U42866 (N_42866,N_42748,N_42572);
xnor U42867 (N_42867,N_42583,N_42639);
or U42868 (N_42868,N_42545,N_42647);
and U42869 (N_42869,N_42626,N_42665);
xor U42870 (N_42870,N_42507,N_42542);
nor U42871 (N_42871,N_42534,N_42712);
or U42872 (N_42872,N_42616,N_42742);
and U42873 (N_42873,N_42746,N_42650);
xnor U42874 (N_42874,N_42596,N_42609);
xor U42875 (N_42875,N_42501,N_42677);
or U42876 (N_42876,N_42608,N_42662);
xor U42877 (N_42877,N_42638,N_42633);
or U42878 (N_42878,N_42613,N_42668);
nor U42879 (N_42879,N_42677,N_42631);
xor U42880 (N_42880,N_42718,N_42662);
nor U42881 (N_42881,N_42614,N_42611);
nand U42882 (N_42882,N_42694,N_42683);
nor U42883 (N_42883,N_42633,N_42552);
xor U42884 (N_42884,N_42640,N_42576);
nor U42885 (N_42885,N_42647,N_42571);
or U42886 (N_42886,N_42707,N_42540);
and U42887 (N_42887,N_42534,N_42521);
and U42888 (N_42888,N_42544,N_42547);
or U42889 (N_42889,N_42709,N_42643);
xor U42890 (N_42890,N_42535,N_42717);
xor U42891 (N_42891,N_42613,N_42607);
and U42892 (N_42892,N_42581,N_42602);
nand U42893 (N_42893,N_42529,N_42724);
nor U42894 (N_42894,N_42548,N_42583);
xor U42895 (N_42895,N_42562,N_42618);
or U42896 (N_42896,N_42625,N_42609);
or U42897 (N_42897,N_42515,N_42733);
nor U42898 (N_42898,N_42683,N_42538);
or U42899 (N_42899,N_42633,N_42524);
or U42900 (N_42900,N_42606,N_42605);
nand U42901 (N_42901,N_42598,N_42589);
xnor U42902 (N_42902,N_42507,N_42730);
and U42903 (N_42903,N_42619,N_42516);
and U42904 (N_42904,N_42722,N_42626);
or U42905 (N_42905,N_42745,N_42554);
nand U42906 (N_42906,N_42749,N_42555);
xor U42907 (N_42907,N_42514,N_42551);
xnor U42908 (N_42908,N_42539,N_42686);
and U42909 (N_42909,N_42532,N_42613);
nand U42910 (N_42910,N_42554,N_42585);
nand U42911 (N_42911,N_42529,N_42508);
nand U42912 (N_42912,N_42539,N_42636);
xor U42913 (N_42913,N_42737,N_42517);
and U42914 (N_42914,N_42614,N_42691);
xnor U42915 (N_42915,N_42646,N_42655);
nand U42916 (N_42916,N_42592,N_42739);
nor U42917 (N_42917,N_42715,N_42619);
nor U42918 (N_42918,N_42550,N_42595);
or U42919 (N_42919,N_42610,N_42718);
and U42920 (N_42920,N_42739,N_42566);
or U42921 (N_42921,N_42675,N_42556);
nor U42922 (N_42922,N_42670,N_42545);
nor U42923 (N_42923,N_42694,N_42549);
and U42924 (N_42924,N_42508,N_42565);
nor U42925 (N_42925,N_42680,N_42675);
nor U42926 (N_42926,N_42640,N_42698);
nor U42927 (N_42927,N_42737,N_42632);
or U42928 (N_42928,N_42514,N_42724);
xnor U42929 (N_42929,N_42656,N_42522);
nor U42930 (N_42930,N_42533,N_42684);
nand U42931 (N_42931,N_42689,N_42579);
xnor U42932 (N_42932,N_42615,N_42555);
nor U42933 (N_42933,N_42640,N_42516);
xnor U42934 (N_42934,N_42674,N_42638);
or U42935 (N_42935,N_42728,N_42586);
and U42936 (N_42936,N_42682,N_42552);
nand U42937 (N_42937,N_42681,N_42748);
xor U42938 (N_42938,N_42509,N_42717);
nand U42939 (N_42939,N_42506,N_42587);
or U42940 (N_42940,N_42531,N_42712);
nor U42941 (N_42941,N_42609,N_42531);
and U42942 (N_42942,N_42503,N_42505);
nand U42943 (N_42943,N_42651,N_42548);
xor U42944 (N_42944,N_42626,N_42633);
and U42945 (N_42945,N_42550,N_42628);
and U42946 (N_42946,N_42505,N_42696);
nor U42947 (N_42947,N_42593,N_42599);
or U42948 (N_42948,N_42727,N_42601);
nand U42949 (N_42949,N_42734,N_42585);
and U42950 (N_42950,N_42522,N_42643);
or U42951 (N_42951,N_42652,N_42573);
nor U42952 (N_42952,N_42730,N_42552);
or U42953 (N_42953,N_42606,N_42742);
and U42954 (N_42954,N_42518,N_42695);
and U42955 (N_42955,N_42657,N_42569);
nand U42956 (N_42956,N_42574,N_42510);
nand U42957 (N_42957,N_42617,N_42636);
xnor U42958 (N_42958,N_42596,N_42656);
and U42959 (N_42959,N_42706,N_42745);
and U42960 (N_42960,N_42589,N_42623);
or U42961 (N_42961,N_42625,N_42716);
xor U42962 (N_42962,N_42515,N_42619);
xnor U42963 (N_42963,N_42592,N_42547);
nand U42964 (N_42964,N_42510,N_42655);
or U42965 (N_42965,N_42680,N_42502);
and U42966 (N_42966,N_42691,N_42625);
nand U42967 (N_42967,N_42613,N_42602);
or U42968 (N_42968,N_42595,N_42715);
nor U42969 (N_42969,N_42644,N_42632);
nor U42970 (N_42970,N_42531,N_42513);
nand U42971 (N_42971,N_42697,N_42607);
nand U42972 (N_42972,N_42676,N_42583);
xnor U42973 (N_42973,N_42605,N_42740);
xnor U42974 (N_42974,N_42675,N_42536);
nor U42975 (N_42975,N_42734,N_42559);
or U42976 (N_42976,N_42707,N_42567);
xnor U42977 (N_42977,N_42747,N_42636);
xor U42978 (N_42978,N_42507,N_42656);
nand U42979 (N_42979,N_42699,N_42735);
nand U42980 (N_42980,N_42535,N_42579);
nor U42981 (N_42981,N_42501,N_42557);
nand U42982 (N_42982,N_42573,N_42721);
xnor U42983 (N_42983,N_42685,N_42608);
xor U42984 (N_42984,N_42742,N_42667);
nand U42985 (N_42985,N_42594,N_42596);
xor U42986 (N_42986,N_42613,N_42727);
nand U42987 (N_42987,N_42530,N_42523);
nor U42988 (N_42988,N_42608,N_42635);
nor U42989 (N_42989,N_42616,N_42528);
xor U42990 (N_42990,N_42532,N_42514);
or U42991 (N_42991,N_42742,N_42531);
and U42992 (N_42992,N_42546,N_42676);
xnor U42993 (N_42993,N_42707,N_42664);
and U42994 (N_42994,N_42562,N_42592);
or U42995 (N_42995,N_42518,N_42633);
xnor U42996 (N_42996,N_42686,N_42620);
nor U42997 (N_42997,N_42668,N_42649);
nand U42998 (N_42998,N_42513,N_42649);
or U42999 (N_42999,N_42526,N_42537);
or U43000 (N_43000,N_42960,N_42841);
nor U43001 (N_43001,N_42787,N_42817);
and U43002 (N_43002,N_42823,N_42938);
xor U43003 (N_43003,N_42861,N_42965);
nor U43004 (N_43004,N_42935,N_42788);
nor U43005 (N_43005,N_42846,N_42837);
nand U43006 (N_43006,N_42816,N_42862);
xnor U43007 (N_43007,N_42864,N_42835);
or U43008 (N_43008,N_42998,N_42912);
nor U43009 (N_43009,N_42848,N_42959);
and U43010 (N_43010,N_42875,N_42954);
nor U43011 (N_43011,N_42932,N_42867);
xor U43012 (N_43012,N_42770,N_42913);
nor U43013 (N_43013,N_42865,N_42961);
xnor U43014 (N_43014,N_42888,N_42974);
nand U43015 (N_43015,N_42937,N_42901);
nor U43016 (N_43016,N_42766,N_42811);
nor U43017 (N_43017,N_42898,N_42880);
and U43018 (N_43018,N_42863,N_42918);
and U43019 (N_43019,N_42869,N_42903);
nand U43020 (N_43020,N_42765,N_42896);
and U43021 (N_43021,N_42893,N_42845);
xnor U43022 (N_43022,N_42904,N_42849);
xor U43023 (N_43023,N_42943,N_42806);
and U43024 (N_43024,N_42897,N_42923);
or U43025 (N_43025,N_42884,N_42828);
xor U43026 (N_43026,N_42762,N_42815);
or U43027 (N_43027,N_42881,N_42900);
or U43028 (N_43028,N_42831,N_42751);
and U43029 (N_43029,N_42919,N_42885);
nand U43030 (N_43030,N_42907,N_42836);
nor U43031 (N_43031,N_42874,N_42780);
or U43032 (N_43032,N_42839,N_42908);
and U43033 (N_43033,N_42833,N_42922);
xnor U43034 (N_43034,N_42814,N_42752);
nand U43035 (N_43035,N_42853,N_42826);
xor U43036 (N_43036,N_42995,N_42952);
xor U43037 (N_43037,N_42772,N_42796);
nand U43038 (N_43038,N_42980,N_42967);
nand U43039 (N_43039,N_42777,N_42911);
or U43040 (N_43040,N_42971,N_42802);
nor U43041 (N_43041,N_42946,N_42989);
nand U43042 (N_43042,N_42887,N_42803);
nand U43043 (N_43043,N_42969,N_42930);
xnor U43044 (N_43044,N_42857,N_42992);
xor U43045 (N_43045,N_42829,N_42789);
nor U43046 (N_43046,N_42855,N_42760);
nor U43047 (N_43047,N_42868,N_42878);
nor U43048 (N_43048,N_42753,N_42889);
nor U43049 (N_43049,N_42798,N_42939);
xnor U43050 (N_43050,N_42776,N_42944);
and U43051 (N_43051,N_42936,N_42822);
xor U43052 (N_43052,N_42977,N_42894);
and U43053 (N_43053,N_42758,N_42956);
or U43054 (N_43054,N_42851,N_42941);
xor U43055 (N_43055,N_42914,N_42764);
xor U43056 (N_43056,N_42994,N_42993);
xor U43057 (N_43057,N_42949,N_42856);
nor U43058 (N_43058,N_42926,N_42870);
xnor U43059 (N_43059,N_42999,N_42834);
xnor U43060 (N_43060,N_42779,N_42882);
and U43061 (N_43061,N_42808,N_42792);
nor U43062 (N_43062,N_42842,N_42825);
xor U43063 (N_43063,N_42850,N_42830);
or U43064 (N_43064,N_42920,N_42940);
and U43065 (N_43065,N_42948,N_42866);
nor U43066 (N_43066,N_42951,N_42966);
and U43067 (N_43067,N_42810,N_42942);
xor U43068 (N_43068,N_42793,N_42947);
and U43069 (N_43069,N_42860,N_42891);
or U43070 (N_43070,N_42791,N_42819);
xor U43071 (N_43071,N_42763,N_42872);
nand U43072 (N_43072,N_42988,N_42986);
nor U43073 (N_43073,N_42858,N_42818);
xnor U43074 (N_43074,N_42976,N_42963);
xor U43075 (N_43075,N_42964,N_42783);
nor U43076 (N_43076,N_42812,N_42854);
nand U43077 (N_43077,N_42924,N_42945);
nor U43078 (N_43078,N_42785,N_42928);
or U43079 (N_43079,N_42794,N_42757);
xor U43080 (N_43080,N_42800,N_42782);
nor U43081 (N_43081,N_42982,N_42955);
nor U43082 (N_43082,N_42805,N_42756);
xnor U43083 (N_43083,N_42997,N_42990);
or U43084 (N_43084,N_42905,N_42821);
and U43085 (N_43085,N_42934,N_42877);
nand U43086 (N_43086,N_42917,N_42767);
xnor U43087 (N_43087,N_42979,N_42873);
nor U43088 (N_43088,N_42902,N_42886);
nand U43089 (N_43089,N_42844,N_42883);
nor U43090 (N_43090,N_42786,N_42983);
nand U43091 (N_43091,N_42771,N_42859);
and U43092 (N_43092,N_42892,N_42968);
nand U43093 (N_43093,N_42820,N_42784);
or U43094 (N_43094,N_42950,N_42921);
nor U43095 (N_43095,N_42809,N_42754);
or U43096 (N_43096,N_42832,N_42987);
and U43097 (N_43097,N_42958,N_42906);
nand U43098 (N_43098,N_42797,N_42929);
xnor U43099 (N_43099,N_42962,N_42985);
xnor U43100 (N_43100,N_42807,N_42996);
nor U43101 (N_43101,N_42775,N_42773);
or U43102 (N_43102,N_42978,N_42991);
or U43103 (N_43103,N_42953,N_42824);
nand U43104 (N_43104,N_42895,N_42790);
nor U43105 (N_43105,N_42876,N_42970);
or U43106 (N_43106,N_42761,N_42843);
nor U43107 (N_43107,N_42910,N_42774);
and U43108 (N_43108,N_42890,N_42781);
and U43109 (N_43109,N_42871,N_42750);
or U43110 (N_43110,N_42768,N_42759);
or U43111 (N_43111,N_42957,N_42847);
and U43112 (N_43112,N_42972,N_42931);
xnor U43113 (N_43113,N_42840,N_42838);
and U43114 (N_43114,N_42925,N_42981);
xor U43115 (N_43115,N_42769,N_42813);
and U43116 (N_43116,N_42909,N_42795);
nor U43117 (N_43117,N_42801,N_42804);
nor U43118 (N_43118,N_42827,N_42933);
nor U43119 (N_43119,N_42755,N_42975);
nor U43120 (N_43120,N_42799,N_42879);
or U43121 (N_43121,N_42852,N_42915);
or U43122 (N_43122,N_42973,N_42927);
or U43123 (N_43123,N_42778,N_42899);
and U43124 (N_43124,N_42916,N_42984);
xnor U43125 (N_43125,N_42830,N_42910);
xnor U43126 (N_43126,N_42763,N_42797);
nand U43127 (N_43127,N_42946,N_42819);
xnor U43128 (N_43128,N_42957,N_42858);
xnor U43129 (N_43129,N_42889,N_42756);
nand U43130 (N_43130,N_42754,N_42757);
xor U43131 (N_43131,N_42876,N_42998);
xor U43132 (N_43132,N_42816,N_42779);
or U43133 (N_43133,N_42946,N_42950);
nand U43134 (N_43134,N_42803,N_42920);
xor U43135 (N_43135,N_42955,N_42952);
nor U43136 (N_43136,N_42787,N_42889);
nand U43137 (N_43137,N_42948,N_42913);
nor U43138 (N_43138,N_42908,N_42817);
or U43139 (N_43139,N_42879,N_42826);
and U43140 (N_43140,N_42788,N_42940);
nand U43141 (N_43141,N_42959,N_42922);
nand U43142 (N_43142,N_42932,N_42830);
nor U43143 (N_43143,N_42990,N_42920);
and U43144 (N_43144,N_42895,N_42819);
xor U43145 (N_43145,N_42945,N_42995);
nand U43146 (N_43146,N_42930,N_42964);
xnor U43147 (N_43147,N_42955,N_42860);
and U43148 (N_43148,N_42945,N_42830);
and U43149 (N_43149,N_42804,N_42883);
xor U43150 (N_43150,N_42988,N_42980);
or U43151 (N_43151,N_42753,N_42820);
nor U43152 (N_43152,N_42815,N_42868);
nand U43153 (N_43153,N_42949,N_42901);
nand U43154 (N_43154,N_42906,N_42865);
xor U43155 (N_43155,N_42843,N_42776);
nand U43156 (N_43156,N_42819,N_42816);
or U43157 (N_43157,N_42776,N_42823);
and U43158 (N_43158,N_42966,N_42758);
nor U43159 (N_43159,N_42902,N_42965);
nor U43160 (N_43160,N_42845,N_42932);
nand U43161 (N_43161,N_42910,N_42806);
xor U43162 (N_43162,N_42973,N_42865);
xor U43163 (N_43163,N_42797,N_42989);
nor U43164 (N_43164,N_42927,N_42901);
xnor U43165 (N_43165,N_42902,N_42850);
or U43166 (N_43166,N_42917,N_42786);
nand U43167 (N_43167,N_42850,N_42946);
xor U43168 (N_43168,N_42842,N_42984);
and U43169 (N_43169,N_42760,N_42751);
and U43170 (N_43170,N_42823,N_42957);
or U43171 (N_43171,N_42874,N_42950);
or U43172 (N_43172,N_42908,N_42968);
and U43173 (N_43173,N_42801,N_42891);
nand U43174 (N_43174,N_42774,N_42864);
xor U43175 (N_43175,N_42951,N_42760);
and U43176 (N_43176,N_42801,N_42824);
xor U43177 (N_43177,N_42994,N_42846);
and U43178 (N_43178,N_42839,N_42826);
xnor U43179 (N_43179,N_42786,N_42752);
xor U43180 (N_43180,N_42927,N_42964);
xor U43181 (N_43181,N_42989,N_42985);
xor U43182 (N_43182,N_42953,N_42978);
nand U43183 (N_43183,N_42989,N_42840);
xor U43184 (N_43184,N_42845,N_42902);
and U43185 (N_43185,N_42990,N_42928);
xor U43186 (N_43186,N_42838,N_42836);
and U43187 (N_43187,N_42895,N_42942);
and U43188 (N_43188,N_42911,N_42967);
nand U43189 (N_43189,N_42946,N_42774);
xor U43190 (N_43190,N_42910,N_42983);
and U43191 (N_43191,N_42834,N_42788);
nor U43192 (N_43192,N_42964,N_42943);
xnor U43193 (N_43193,N_42761,N_42803);
or U43194 (N_43194,N_42873,N_42905);
xor U43195 (N_43195,N_42818,N_42813);
or U43196 (N_43196,N_42977,N_42998);
nor U43197 (N_43197,N_42937,N_42796);
and U43198 (N_43198,N_42823,N_42834);
xor U43199 (N_43199,N_42760,N_42977);
xor U43200 (N_43200,N_42824,N_42787);
or U43201 (N_43201,N_42958,N_42881);
or U43202 (N_43202,N_42861,N_42856);
or U43203 (N_43203,N_42792,N_42996);
nand U43204 (N_43204,N_42941,N_42885);
xor U43205 (N_43205,N_42854,N_42821);
nor U43206 (N_43206,N_42756,N_42812);
xnor U43207 (N_43207,N_42807,N_42828);
and U43208 (N_43208,N_42781,N_42846);
nand U43209 (N_43209,N_42938,N_42812);
or U43210 (N_43210,N_42785,N_42837);
or U43211 (N_43211,N_42759,N_42941);
or U43212 (N_43212,N_42818,N_42884);
or U43213 (N_43213,N_42870,N_42878);
and U43214 (N_43214,N_42942,N_42933);
xor U43215 (N_43215,N_42861,N_42763);
nand U43216 (N_43216,N_42782,N_42949);
or U43217 (N_43217,N_42926,N_42820);
or U43218 (N_43218,N_42753,N_42956);
and U43219 (N_43219,N_42827,N_42856);
nor U43220 (N_43220,N_42839,N_42767);
and U43221 (N_43221,N_42951,N_42946);
or U43222 (N_43222,N_42893,N_42903);
nand U43223 (N_43223,N_42759,N_42751);
nor U43224 (N_43224,N_42885,N_42782);
or U43225 (N_43225,N_42978,N_42764);
and U43226 (N_43226,N_42940,N_42903);
or U43227 (N_43227,N_42875,N_42832);
and U43228 (N_43228,N_42891,N_42842);
and U43229 (N_43229,N_42844,N_42905);
nand U43230 (N_43230,N_42796,N_42863);
nand U43231 (N_43231,N_42957,N_42922);
nand U43232 (N_43232,N_42794,N_42993);
or U43233 (N_43233,N_42936,N_42783);
and U43234 (N_43234,N_42796,N_42821);
or U43235 (N_43235,N_42965,N_42914);
or U43236 (N_43236,N_42762,N_42870);
and U43237 (N_43237,N_42987,N_42761);
nor U43238 (N_43238,N_42902,N_42814);
nor U43239 (N_43239,N_42812,N_42814);
xnor U43240 (N_43240,N_42775,N_42854);
or U43241 (N_43241,N_42835,N_42935);
or U43242 (N_43242,N_42796,N_42835);
nor U43243 (N_43243,N_42849,N_42919);
or U43244 (N_43244,N_42924,N_42800);
nor U43245 (N_43245,N_42956,N_42905);
and U43246 (N_43246,N_42761,N_42807);
nand U43247 (N_43247,N_42968,N_42933);
xor U43248 (N_43248,N_42861,N_42857);
xor U43249 (N_43249,N_42894,N_42831);
nor U43250 (N_43250,N_43128,N_43054);
nand U43251 (N_43251,N_43105,N_43033);
nor U43252 (N_43252,N_43204,N_43151);
and U43253 (N_43253,N_43032,N_43131);
nand U43254 (N_43254,N_43188,N_43114);
xnor U43255 (N_43255,N_43202,N_43162);
nor U43256 (N_43256,N_43058,N_43019);
nor U43257 (N_43257,N_43022,N_43107);
and U43258 (N_43258,N_43067,N_43237);
and U43259 (N_43259,N_43226,N_43144);
xnor U43260 (N_43260,N_43175,N_43078);
nand U43261 (N_43261,N_43129,N_43183);
or U43262 (N_43262,N_43243,N_43005);
nand U43263 (N_43263,N_43222,N_43241);
xor U43264 (N_43264,N_43136,N_43220);
xnor U43265 (N_43265,N_43205,N_43004);
or U43266 (N_43266,N_43198,N_43135);
nand U43267 (N_43267,N_43166,N_43024);
and U43268 (N_43268,N_43191,N_43096);
nand U43269 (N_43269,N_43210,N_43133);
xnor U43270 (N_43270,N_43130,N_43164);
xnor U43271 (N_43271,N_43057,N_43224);
or U43272 (N_43272,N_43139,N_43143);
xor U43273 (N_43273,N_43091,N_43169);
nand U43274 (N_43274,N_43152,N_43190);
nor U43275 (N_43275,N_43213,N_43120);
and U43276 (N_43276,N_43235,N_43141);
or U43277 (N_43277,N_43048,N_43148);
xnor U43278 (N_43278,N_43047,N_43240);
xor U43279 (N_43279,N_43097,N_43159);
and U43280 (N_43280,N_43248,N_43092);
nand U43281 (N_43281,N_43084,N_43149);
nand U43282 (N_43282,N_43008,N_43249);
nor U43283 (N_43283,N_43095,N_43112);
and U43284 (N_43284,N_43173,N_43037);
nor U43285 (N_43285,N_43014,N_43116);
xnor U43286 (N_43286,N_43167,N_43045);
and U43287 (N_43287,N_43117,N_43232);
xor U43288 (N_43288,N_43077,N_43076);
nand U43289 (N_43289,N_43200,N_43036);
nor U43290 (N_43290,N_43034,N_43225);
and U43291 (N_43291,N_43184,N_43062);
or U43292 (N_43292,N_43000,N_43214);
nor U43293 (N_43293,N_43061,N_43111);
nand U43294 (N_43294,N_43073,N_43104);
or U43295 (N_43295,N_43127,N_43216);
or U43296 (N_43296,N_43098,N_43158);
or U43297 (N_43297,N_43094,N_43020);
or U43298 (N_43298,N_43182,N_43121);
and U43299 (N_43299,N_43247,N_43060);
and U43300 (N_43300,N_43163,N_43132);
nand U43301 (N_43301,N_43203,N_43142);
xnor U43302 (N_43302,N_43042,N_43122);
nor U43303 (N_43303,N_43012,N_43137);
nor U43304 (N_43304,N_43089,N_43177);
nand U43305 (N_43305,N_43160,N_43046);
or U43306 (N_43306,N_43108,N_43103);
nor U43307 (N_43307,N_43236,N_43170);
and U43308 (N_43308,N_43211,N_43195);
or U43309 (N_43309,N_43192,N_43146);
nand U43310 (N_43310,N_43126,N_43038);
or U43311 (N_43311,N_43185,N_43118);
or U43312 (N_43312,N_43081,N_43233);
nand U43313 (N_43313,N_43099,N_43178);
nand U43314 (N_43314,N_43083,N_43113);
xnor U43315 (N_43315,N_43219,N_43080);
nor U43316 (N_43316,N_43196,N_43199);
nor U43317 (N_43317,N_43172,N_43227);
nor U43318 (N_43318,N_43231,N_43056);
xnor U43319 (N_43319,N_43215,N_43015);
and U43320 (N_43320,N_43055,N_43059);
nand U43321 (N_43321,N_43110,N_43119);
nand U43322 (N_43322,N_43171,N_43180);
and U43323 (N_43323,N_43193,N_43039);
nand U43324 (N_43324,N_43138,N_43230);
or U43325 (N_43325,N_43018,N_43074);
nand U43326 (N_43326,N_43168,N_43026);
or U43327 (N_43327,N_43041,N_43245);
xnor U43328 (N_43328,N_43246,N_43154);
xor U43329 (N_43329,N_43021,N_43006);
nor U43330 (N_43330,N_43102,N_43157);
xnor U43331 (N_43331,N_43066,N_43176);
xor U43332 (N_43332,N_43106,N_43187);
xor U43333 (N_43333,N_43050,N_43063);
nand U43334 (N_43334,N_43031,N_43186);
and U43335 (N_43335,N_43189,N_43082);
or U43336 (N_43336,N_43001,N_43075);
and U43337 (N_43337,N_43044,N_43239);
nor U43338 (N_43338,N_43155,N_43016);
nand U43339 (N_43339,N_43011,N_43147);
and U43340 (N_43340,N_43087,N_43124);
nor U43341 (N_43341,N_43068,N_43065);
or U43342 (N_43342,N_43028,N_43093);
nand U43343 (N_43343,N_43051,N_43145);
and U43344 (N_43344,N_43052,N_43197);
or U43345 (N_43345,N_43156,N_43221);
nand U43346 (N_43346,N_43072,N_43207);
nor U43347 (N_43347,N_43115,N_43174);
or U43348 (N_43348,N_43194,N_43070);
or U43349 (N_43349,N_43201,N_43181);
nor U43350 (N_43350,N_43134,N_43242);
and U43351 (N_43351,N_43085,N_43064);
xnor U43352 (N_43352,N_43040,N_43209);
and U43353 (N_43353,N_43208,N_43053);
nor U43354 (N_43354,N_43140,N_43086);
and U43355 (N_43355,N_43234,N_43030);
nand U43356 (N_43356,N_43244,N_43007);
and U43357 (N_43357,N_43238,N_43017);
or U43358 (N_43358,N_43218,N_43043);
nand U43359 (N_43359,N_43079,N_43229);
nand U43360 (N_43360,N_43013,N_43153);
or U43361 (N_43361,N_43002,N_43150);
and U43362 (N_43362,N_43101,N_43090);
and U43363 (N_43363,N_43009,N_43010);
or U43364 (N_43364,N_43165,N_43025);
nand U43365 (N_43365,N_43125,N_43027);
nor U43366 (N_43366,N_43109,N_43217);
or U43367 (N_43367,N_43049,N_43023);
nand U43368 (N_43368,N_43071,N_43223);
or U43369 (N_43369,N_43228,N_43123);
and U43370 (N_43370,N_43179,N_43035);
and U43371 (N_43371,N_43029,N_43003);
nor U43372 (N_43372,N_43161,N_43100);
xor U43373 (N_43373,N_43206,N_43088);
nand U43374 (N_43374,N_43069,N_43212);
or U43375 (N_43375,N_43111,N_43150);
nor U43376 (N_43376,N_43120,N_43228);
nand U43377 (N_43377,N_43180,N_43185);
nor U43378 (N_43378,N_43087,N_43044);
nand U43379 (N_43379,N_43043,N_43102);
xnor U43380 (N_43380,N_43036,N_43223);
nor U43381 (N_43381,N_43223,N_43106);
and U43382 (N_43382,N_43215,N_43192);
and U43383 (N_43383,N_43184,N_43012);
or U43384 (N_43384,N_43071,N_43092);
or U43385 (N_43385,N_43173,N_43202);
xor U43386 (N_43386,N_43087,N_43225);
nand U43387 (N_43387,N_43214,N_43084);
and U43388 (N_43388,N_43242,N_43078);
nor U43389 (N_43389,N_43043,N_43172);
nor U43390 (N_43390,N_43066,N_43168);
or U43391 (N_43391,N_43115,N_43037);
nand U43392 (N_43392,N_43224,N_43053);
xnor U43393 (N_43393,N_43230,N_43058);
nand U43394 (N_43394,N_43061,N_43033);
nand U43395 (N_43395,N_43195,N_43210);
nor U43396 (N_43396,N_43223,N_43244);
and U43397 (N_43397,N_43046,N_43175);
or U43398 (N_43398,N_43164,N_43048);
and U43399 (N_43399,N_43034,N_43033);
nor U43400 (N_43400,N_43171,N_43231);
nor U43401 (N_43401,N_43062,N_43112);
nand U43402 (N_43402,N_43154,N_43228);
nor U43403 (N_43403,N_43160,N_43201);
or U43404 (N_43404,N_43106,N_43152);
and U43405 (N_43405,N_43097,N_43118);
and U43406 (N_43406,N_43035,N_43149);
xnor U43407 (N_43407,N_43232,N_43176);
or U43408 (N_43408,N_43186,N_43045);
or U43409 (N_43409,N_43142,N_43168);
and U43410 (N_43410,N_43083,N_43102);
or U43411 (N_43411,N_43071,N_43062);
and U43412 (N_43412,N_43122,N_43033);
or U43413 (N_43413,N_43132,N_43062);
xor U43414 (N_43414,N_43036,N_43164);
and U43415 (N_43415,N_43177,N_43094);
nand U43416 (N_43416,N_43031,N_43246);
xnor U43417 (N_43417,N_43052,N_43147);
or U43418 (N_43418,N_43113,N_43245);
nand U43419 (N_43419,N_43171,N_43217);
and U43420 (N_43420,N_43037,N_43154);
nor U43421 (N_43421,N_43172,N_43088);
nand U43422 (N_43422,N_43177,N_43133);
nor U43423 (N_43423,N_43122,N_43209);
or U43424 (N_43424,N_43157,N_43123);
and U43425 (N_43425,N_43141,N_43125);
and U43426 (N_43426,N_43154,N_43044);
or U43427 (N_43427,N_43103,N_43172);
or U43428 (N_43428,N_43078,N_43003);
or U43429 (N_43429,N_43062,N_43214);
xnor U43430 (N_43430,N_43002,N_43053);
and U43431 (N_43431,N_43225,N_43006);
or U43432 (N_43432,N_43073,N_43035);
nand U43433 (N_43433,N_43208,N_43150);
xor U43434 (N_43434,N_43161,N_43099);
nor U43435 (N_43435,N_43197,N_43113);
and U43436 (N_43436,N_43165,N_43245);
nor U43437 (N_43437,N_43085,N_43241);
or U43438 (N_43438,N_43147,N_43056);
nand U43439 (N_43439,N_43246,N_43008);
nor U43440 (N_43440,N_43035,N_43167);
and U43441 (N_43441,N_43186,N_43134);
or U43442 (N_43442,N_43112,N_43056);
and U43443 (N_43443,N_43138,N_43080);
nor U43444 (N_43444,N_43179,N_43207);
nor U43445 (N_43445,N_43034,N_43036);
nand U43446 (N_43446,N_43049,N_43048);
nand U43447 (N_43447,N_43121,N_43148);
nor U43448 (N_43448,N_43205,N_43046);
and U43449 (N_43449,N_43007,N_43150);
nor U43450 (N_43450,N_43126,N_43138);
or U43451 (N_43451,N_43133,N_43044);
and U43452 (N_43452,N_43161,N_43154);
or U43453 (N_43453,N_43179,N_43191);
or U43454 (N_43454,N_43171,N_43029);
xnor U43455 (N_43455,N_43006,N_43229);
or U43456 (N_43456,N_43196,N_43108);
and U43457 (N_43457,N_43151,N_43168);
xor U43458 (N_43458,N_43183,N_43209);
nor U43459 (N_43459,N_43068,N_43033);
xor U43460 (N_43460,N_43092,N_43236);
xnor U43461 (N_43461,N_43046,N_43247);
xor U43462 (N_43462,N_43138,N_43140);
and U43463 (N_43463,N_43218,N_43243);
nand U43464 (N_43464,N_43081,N_43247);
xnor U43465 (N_43465,N_43052,N_43072);
nor U43466 (N_43466,N_43065,N_43027);
nor U43467 (N_43467,N_43068,N_43185);
xnor U43468 (N_43468,N_43073,N_43111);
nand U43469 (N_43469,N_43115,N_43105);
and U43470 (N_43470,N_43215,N_43070);
nor U43471 (N_43471,N_43207,N_43206);
and U43472 (N_43472,N_43106,N_43236);
nor U43473 (N_43473,N_43050,N_43173);
xor U43474 (N_43474,N_43008,N_43213);
and U43475 (N_43475,N_43126,N_43178);
xor U43476 (N_43476,N_43210,N_43216);
nand U43477 (N_43477,N_43095,N_43087);
nand U43478 (N_43478,N_43017,N_43145);
xor U43479 (N_43479,N_43019,N_43201);
and U43480 (N_43480,N_43132,N_43087);
xnor U43481 (N_43481,N_43213,N_43238);
or U43482 (N_43482,N_43237,N_43226);
or U43483 (N_43483,N_43128,N_43214);
nand U43484 (N_43484,N_43234,N_43105);
nor U43485 (N_43485,N_43244,N_43162);
nand U43486 (N_43486,N_43150,N_43198);
and U43487 (N_43487,N_43052,N_43207);
or U43488 (N_43488,N_43054,N_43018);
nor U43489 (N_43489,N_43234,N_43091);
and U43490 (N_43490,N_43036,N_43183);
nand U43491 (N_43491,N_43027,N_43159);
or U43492 (N_43492,N_43069,N_43183);
or U43493 (N_43493,N_43222,N_43186);
and U43494 (N_43494,N_43244,N_43035);
nor U43495 (N_43495,N_43242,N_43030);
xor U43496 (N_43496,N_43078,N_43080);
nand U43497 (N_43497,N_43169,N_43194);
and U43498 (N_43498,N_43218,N_43176);
and U43499 (N_43499,N_43249,N_43055);
nor U43500 (N_43500,N_43471,N_43404);
nor U43501 (N_43501,N_43464,N_43498);
nor U43502 (N_43502,N_43463,N_43439);
or U43503 (N_43503,N_43452,N_43408);
or U43504 (N_43504,N_43405,N_43455);
xnor U43505 (N_43505,N_43328,N_43494);
and U43506 (N_43506,N_43353,N_43359);
nand U43507 (N_43507,N_43436,N_43312);
nor U43508 (N_43508,N_43289,N_43402);
nor U43509 (N_43509,N_43496,N_43443);
nor U43510 (N_43510,N_43298,N_43357);
and U43511 (N_43511,N_43480,N_43479);
nor U43512 (N_43512,N_43485,N_43320);
xnor U43513 (N_43513,N_43414,N_43447);
nand U43514 (N_43514,N_43432,N_43440);
or U43515 (N_43515,N_43341,N_43456);
and U43516 (N_43516,N_43273,N_43412);
or U43517 (N_43517,N_43415,N_43269);
nor U43518 (N_43518,N_43453,N_43295);
or U43519 (N_43519,N_43347,N_43260);
and U43520 (N_43520,N_43316,N_43278);
and U43521 (N_43521,N_43346,N_43286);
or U43522 (N_43522,N_43251,N_43259);
or U43523 (N_43523,N_43399,N_43338);
nand U43524 (N_43524,N_43313,N_43390);
xor U43525 (N_43525,N_43413,N_43499);
nor U43526 (N_43526,N_43334,N_43311);
nor U43527 (N_43527,N_43491,N_43336);
xor U43528 (N_43528,N_43488,N_43290);
nand U43529 (N_43529,N_43300,N_43431);
nor U43530 (N_43530,N_43417,N_43492);
nand U43531 (N_43531,N_43296,N_43352);
xnor U43532 (N_43532,N_43287,N_43477);
and U43533 (N_43533,N_43327,N_43301);
or U43534 (N_43534,N_43457,N_43377);
nand U43535 (N_43535,N_43279,N_43356);
nand U43536 (N_43536,N_43406,N_43403);
and U43537 (N_43537,N_43398,N_43258);
nor U43538 (N_43538,N_43324,N_43389);
and U43539 (N_43539,N_43252,N_43283);
xor U43540 (N_43540,N_43428,N_43281);
or U43541 (N_43541,N_43266,N_43315);
and U43542 (N_43542,N_43388,N_43309);
nand U43543 (N_43543,N_43468,N_43305);
nand U43544 (N_43544,N_43411,N_43449);
nand U43545 (N_43545,N_43433,N_43358);
nor U43546 (N_43546,N_43255,N_43416);
or U43547 (N_43547,N_43424,N_43372);
nand U43548 (N_43548,N_43318,N_43459);
and U43549 (N_43549,N_43350,N_43345);
xnor U43550 (N_43550,N_43288,N_43284);
or U43551 (N_43551,N_43470,N_43486);
or U43552 (N_43552,N_43314,N_43280);
or U43553 (N_43553,N_43454,N_43422);
or U43554 (N_43554,N_43319,N_43257);
nand U43555 (N_43555,N_43325,N_43374);
or U43556 (N_43556,N_43302,N_43339);
and U43557 (N_43557,N_43475,N_43282);
or U43558 (N_43558,N_43265,N_43364);
or U43559 (N_43559,N_43385,N_43426);
nand U43560 (N_43560,N_43275,N_43423);
nor U43561 (N_43561,N_43310,N_43365);
or U43562 (N_43562,N_43418,N_43373);
nor U43563 (N_43563,N_43493,N_43382);
nor U43564 (N_43564,N_43410,N_43349);
and U43565 (N_43565,N_43381,N_43355);
nor U43566 (N_43566,N_43285,N_43458);
nor U43567 (N_43567,N_43393,N_43421);
nor U43568 (N_43568,N_43461,N_43437);
nor U43569 (N_43569,N_43380,N_43321);
xor U43570 (N_43570,N_43386,N_43267);
nor U43571 (N_43571,N_43445,N_43329);
xor U43572 (N_43572,N_43473,N_43253);
nor U43573 (N_43573,N_43323,N_43474);
and U43574 (N_43574,N_43333,N_43348);
or U43575 (N_43575,N_43276,N_43481);
or U43576 (N_43576,N_43497,N_43427);
nor U43577 (N_43577,N_43397,N_43489);
xnor U43578 (N_43578,N_43272,N_43340);
xor U43579 (N_43579,N_43277,N_43256);
or U43580 (N_43580,N_43262,N_43375);
nor U43581 (N_43581,N_43335,N_43483);
nand U43582 (N_43582,N_43351,N_43342);
xnor U43583 (N_43583,N_43343,N_43448);
and U43584 (N_43584,N_43303,N_43434);
xnor U43585 (N_43585,N_43425,N_43344);
and U43586 (N_43586,N_43482,N_43444);
xor U43587 (N_43587,N_43330,N_43370);
nor U43588 (N_43588,N_43383,N_43307);
nor U43589 (N_43589,N_43490,N_43420);
nor U43590 (N_43590,N_43304,N_43270);
or U43591 (N_43591,N_43419,N_43438);
nor U43592 (N_43592,N_43291,N_43297);
or U43593 (N_43593,N_43429,N_43361);
xor U43594 (N_43594,N_43469,N_43326);
and U43595 (N_43595,N_43441,N_43409);
xor U43596 (N_43596,N_43495,N_43317);
nor U43597 (N_43597,N_43261,N_43379);
or U43598 (N_43598,N_43466,N_43371);
nor U43599 (N_43599,N_43360,N_43299);
nor U43600 (N_43600,N_43430,N_43363);
xnor U43601 (N_43601,N_43391,N_43460);
and U43602 (N_43602,N_43332,N_43368);
xor U43603 (N_43603,N_43442,N_43293);
nand U43604 (N_43604,N_43366,N_43331);
xnor U43605 (N_43605,N_43376,N_43450);
nand U43606 (N_43606,N_43392,N_43484);
or U43607 (N_43607,N_43387,N_43472);
xor U43608 (N_43608,N_43292,N_43263);
nand U43609 (N_43609,N_43487,N_43308);
nor U43610 (N_43610,N_43435,N_43250);
nand U43611 (N_43611,N_43476,N_43294);
or U43612 (N_43612,N_43362,N_43446);
nand U43613 (N_43613,N_43400,N_43254);
and U43614 (N_43614,N_43367,N_43271);
nand U43615 (N_43615,N_43395,N_43274);
nor U43616 (N_43616,N_43369,N_43401);
or U43617 (N_43617,N_43467,N_43384);
or U43618 (N_43618,N_43394,N_43306);
nor U43619 (N_43619,N_43451,N_43378);
nand U43620 (N_43620,N_43264,N_43268);
nand U43621 (N_43621,N_43407,N_43354);
and U43622 (N_43622,N_43322,N_43462);
nor U43623 (N_43623,N_43478,N_43396);
nand U43624 (N_43624,N_43337,N_43465);
or U43625 (N_43625,N_43456,N_43353);
or U43626 (N_43626,N_43261,N_43331);
and U43627 (N_43627,N_43466,N_43308);
nand U43628 (N_43628,N_43268,N_43352);
and U43629 (N_43629,N_43329,N_43268);
nor U43630 (N_43630,N_43289,N_43486);
or U43631 (N_43631,N_43428,N_43384);
or U43632 (N_43632,N_43443,N_43487);
and U43633 (N_43633,N_43427,N_43318);
nor U43634 (N_43634,N_43390,N_43416);
or U43635 (N_43635,N_43446,N_43381);
and U43636 (N_43636,N_43490,N_43293);
xor U43637 (N_43637,N_43271,N_43382);
nor U43638 (N_43638,N_43375,N_43393);
or U43639 (N_43639,N_43455,N_43361);
nand U43640 (N_43640,N_43401,N_43455);
or U43641 (N_43641,N_43266,N_43463);
nor U43642 (N_43642,N_43282,N_43290);
nor U43643 (N_43643,N_43299,N_43399);
or U43644 (N_43644,N_43441,N_43387);
or U43645 (N_43645,N_43421,N_43416);
nand U43646 (N_43646,N_43363,N_43467);
and U43647 (N_43647,N_43429,N_43344);
nor U43648 (N_43648,N_43362,N_43325);
nand U43649 (N_43649,N_43293,N_43444);
nor U43650 (N_43650,N_43391,N_43287);
nand U43651 (N_43651,N_43421,N_43413);
nor U43652 (N_43652,N_43360,N_43478);
xnor U43653 (N_43653,N_43397,N_43463);
xnor U43654 (N_43654,N_43276,N_43297);
nand U43655 (N_43655,N_43431,N_43317);
nor U43656 (N_43656,N_43423,N_43433);
xnor U43657 (N_43657,N_43277,N_43341);
and U43658 (N_43658,N_43306,N_43319);
and U43659 (N_43659,N_43268,N_43387);
or U43660 (N_43660,N_43420,N_43425);
nand U43661 (N_43661,N_43401,N_43310);
nor U43662 (N_43662,N_43335,N_43274);
nand U43663 (N_43663,N_43375,N_43377);
nor U43664 (N_43664,N_43382,N_43302);
or U43665 (N_43665,N_43296,N_43295);
or U43666 (N_43666,N_43320,N_43421);
xor U43667 (N_43667,N_43318,N_43428);
nand U43668 (N_43668,N_43491,N_43412);
xnor U43669 (N_43669,N_43426,N_43391);
or U43670 (N_43670,N_43419,N_43424);
nand U43671 (N_43671,N_43422,N_43473);
and U43672 (N_43672,N_43323,N_43335);
nand U43673 (N_43673,N_43301,N_43474);
and U43674 (N_43674,N_43271,N_43392);
and U43675 (N_43675,N_43434,N_43346);
and U43676 (N_43676,N_43319,N_43251);
and U43677 (N_43677,N_43478,N_43394);
nand U43678 (N_43678,N_43314,N_43273);
nand U43679 (N_43679,N_43351,N_43326);
nand U43680 (N_43680,N_43464,N_43443);
xor U43681 (N_43681,N_43402,N_43328);
nor U43682 (N_43682,N_43453,N_43387);
and U43683 (N_43683,N_43476,N_43379);
nand U43684 (N_43684,N_43404,N_43325);
nor U43685 (N_43685,N_43294,N_43312);
nor U43686 (N_43686,N_43440,N_43363);
or U43687 (N_43687,N_43271,N_43357);
and U43688 (N_43688,N_43456,N_43480);
nand U43689 (N_43689,N_43333,N_43316);
nand U43690 (N_43690,N_43495,N_43295);
or U43691 (N_43691,N_43298,N_43341);
nand U43692 (N_43692,N_43323,N_43283);
xnor U43693 (N_43693,N_43314,N_43328);
xor U43694 (N_43694,N_43469,N_43266);
and U43695 (N_43695,N_43427,N_43320);
xnor U43696 (N_43696,N_43275,N_43362);
and U43697 (N_43697,N_43390,N_43496);
nor U43698 (N_43698,N_43472,N_43378);
or U43699 (N_43699,N_43418,N_43354);
or U43700 (N_43700,N_43421,N_43353);
and U43701 (N_43701,N_43383,N_43267);
nand U43702 (N_43702,N_43313,N_43405);
nor U43703 (N_43703,N_43351,N_43439);
nand U43704 (N_43704,N_43442,N_43462);
nor U43705 (N_43705,N_43443,N_43482);
xor U43706 (N_43706,N_43375,N_43479);
xnor U43707 (N_43707,N_43460,N_43382);
xor U43708 (N_43708,N_43387,N_43426);
xor U43709 (N_43709,N_43362,N_43425);
and U43710 (N_43710,N_43320,N_43334);
nor U43711 (N_43711,N_43413,N_43305);
xnor U43712 (N_43712,N_43293,N_43314);
or U43713 (N_43713,N_43408,N_43467);
nor U43714 (N_43714,N_43273,N_43428);
and U43715 (N_43715,N_43321,N_43452);
and U43716 (N_43716,N_43286,N_43287);
and U43717 (N_43717,N_43299,N_43336);
and U43718 (N_43718,N_43400,N_43475);
nand U43719 (N_43719,N_43397,N_43414);
or U43720 (N_43720,N_43496,N_43366);
or U43721 (N_43721,N_43273,N_43281);
nor U43722 (N_43722,N_43470,N_43403);
xor U43723 (N_43723,N_43401,N_43333);
or U43724 (N_43724,N_43259,N_43393);
and U43725 (N_43725,N_43430,N_43461);
nand U43726 (N_43726,N_43359,N_43290);
nand U43727 (N_43727,N_43374,N_43353);
or U43728 (N_43728,N_43457,N_43321);
nor U43729 (N_43729,N_43494,N_43429);
nand U43730 (N_43730,N_43345,N_43424);
nor U43731 (N_43731,N_43395,N_43400);
nor U43732 (N_43732,N_43475,N_43429);
nor U43733 (N_43733,N_43252,N_43269);
nand U43734 (N_43734,N_43493,N_43316);
nor U43735 (N_43735,N_43353,N_43269);
xor U43736 (N_43736,N_43499,N_43389);
xnor U43737 (N_43737,N_43459,N_43340);
and U43738 (N_43738,N_43393,N_43308);
or U43739 (N_43739,N_43434,N_43289);
nor U43740 (N_43740,N_43380,N_43332);
nand U43741 (N_43741,N_43272,N_43360);
xor U43742 (N_43742,N_43481,N_43414);
and U43743 (N_43743,N_43325,N_43496);
and U43744 (N_43744,N_43470,N_43353);
xor U43745 (N_43745,N_43296,N_43326);
nand U43746 (N_43746,N_43386,N_43379);
nor U43747 (N_43747,N_43320,N_43395);
xnor U43748 (N_43748,N_43397,N_43351);
nand U43749 (N_43749,N_43265,N_43399);
and U43750 (N_43750,N_43617,N_43577);
nor U43751 (N_43751,N_43509,N_43678);
xor U43752 (N_43752,N_43558,N_43560);
or U43753 (N_43753,N_43581,N_43597);
nor U43754 (N_43754,N_43694,N_43653);
nor U43755 (N_43755,N_43710,N_43663);
nand U43756 (N_43756,N_43570,N_43749);
xor U43757 (N_43757,N_43507,N_43588);
and U43758 (N_43758,N_43609,N_43546);
nor U43759 (N_43759,N_43566,N_43649);
and U43760 (N_43760,N_43642,N_43720);
and U43761 (N_43761,N_43547,N_43590);
and U43762 (N_43762,N_43729,N_43575);
nor U43763 (N_43763,N_43563,N_43564);
and U43764 (N_43764,N_43671,N_43626);
and U43765 (N_43765,N_43629,N_43701);
and U43766 (N_43766,N_43711,N_43550);
or U43767 (N_43767,N_43668,N_43623);
nand U43768 (N_43768,N_43722,N_43639);
or U43769 (N_43769,N_43565,N_43712);
xnor U43770 (N_43770,N_43508,N_43601);
or U43771 (N_43771,N_43600,N_43510);
or U43772 (N_43772,N_43709,N_43530);
nand U43773 (N_43773,N_43704,N_43674);
xnor U43774 (N_43774,N_43614,N_43714);
xnor U43775 (N_43775,N_43519,N_43692);
and U43776 (N_43776,N_43611,N_43612);
and U43777 (N_43777,N_43595,N_43707);
nand U43778 (N_43778,N_43531,N_43659);
or U43779 (N_43779,N_43514,N_43666);
nor U43780 (N_43780,N_43598,N_43706);
xor U43781 (N_43781,N_43624,N_43680);
xnor U43782 (N_43782,N_43567,N_43632);
and U43783 (N_43783,N_43693,N_43677);
nand U43784 (N_43784,N_43580,N_43502);
nor U43785 (N_43785,N_43596,N_43736);
nand U43786 (N_43786,N_43535,N_43602);
or U43787 (N_43787,N_43543,N_43631);
and U43788 (N_43788,N_43643,N_43544);
nor U43789 (N_43789,N_43527,N_43583);
and U43790 (N_43790,N_43638,N_43613);
and U43791 (N_43791,N_43656,N_43696);
xor U43792 (N_43792,N_43599,N_43702);
and U43793 (N_43793,N_43705,N_43584);
nor U43794 (N_43794,N_43553,N_43670);
xor U43795 (N_43795,N_43529,N_43726);
and U43796 (N_43796,N_43526,N_43516);
nand U43797 (N_43797,N_43603,N_43651);
nand U43798 (N_43798,N_43619,N_43699);
nor U43799 (N_43799,N_43719,N_43524);
or U43800 (N_43800,N_43733,N_43608);
xor U43801 (N_43801,N_43748,N_43591);
xnor U43802 (N_43802,N_43732,N_43627);
or U43803 (N_43803,N_43579,N_43679);
and U43804 (N_43804,N_43605,N_43673);
nor U43805 (N_43805,N_43697,N_43664);
xor U43806 (N_43806,N_43637,N_43582);
xnor U43807 (N_43807,N_43645,N_43534);
nand U43808 (N_43808,N_43585,N_43685);
or U43809 (N_43809,N_43522,N_43630);
nand U43810 (N_43810,N_43505,N_43655);
and U43811 (N_43811,N_43647,N_43703);
xnor U43812 (N_43812,N_43744,N_43718);
nand U43813 (N_43813,N_43513,N_43503);
or U43814 (N_43814,N_43650,N_43561);
nor U43815 (N_43815,N_43686,N_43657);
nor U43816 (N_43816,N_43745,N_43644);
or U43817 (N_43817,N_43658,N_43594);
or U43818 (N_43818,N_43700,N_43532);
or U43819 (N_43819,N_43646,N_43607);
nor U43820 (N_43820,N_43727,N_43568);
and U43821 (N_43821,N_43549,N_43545);
nor U43822 (N_43822,N_43675,N_43698);
nand U43823 (N_43823,N_43708,N_43569);
and U43824 (N_43824,N_43654,N_43592);
or U43825 (N_43825,N_43572,N_43593);
nand U43826 (N_43826,N_43716,N_43690);
or U43827 (N_43827,N_43735,N_43511);
nor U43828 (N_43828,N_43523,N_43557);
and U43829 (N_43829,N_43578,N_43576);
xnor U43830 (N_43830,N_43731,N_43689);
xor U43831 (N_43831,N_43552,N_43676);
or U43832 (N_43832,N_43562,N_43660);
nor U43833 (N_43833,N_43525,N_43715);
and U43834 (N_43834,N_43661,N_43682);
or U43835 (N_43835,N_43621,N_43728);
and U43836 (N_43836,N_43539,N_43628);
xor U43837 (N_43837,N_43536,N_43622);
nand U43838 (N_43838,N_43742,N_43652);
nand U43839 (N_43839,N_43610,N_43695);
nor U43840 (N_43840,N_43641,N_43625);
xnor U43841 (N_43841,N_43504,N_43648);
nor U43842 (N_43842,N_43683,N_43542);
nor U43843 (N_43843,N_43589,N_43687);
nand U43844 (N_43844,N_43517,N_43633);
xor U43845 (N_43845,N_43747,N_43616);
and U43846 (N_43846,N_43672,N_43515);
nand U43847 (N_43847,N_43541,N_43734);
nand U43848 (N_43848,N_43606,N_43512);
and U43849 (N_43849,N_43571,N_43554);
xnor U43850 (N_43850,N_43620,N_43713);
nand U43851 (N_43851,N_43533,N_43500);
nand U43852 (N_43852,N_43640,N_43501);
xor U43853 (N_43853,N_43555,N_43586);
nand U43854 (N_43854,N_43634,N_43520);
and U43855 (N_43855,N_43725,N_43743);
or U43856 (N_43856,N_43665,N_43506);
nor U43857 (N_43857,N_43730,N_43741);
or U43858 (N_43858,N_43662,N_43739);
or U43859 (N_43859,N_43688,N_43556);
nor U43860 (N_43860,N_43667,N_43740);
nand U43861 (N_43861,N_43684,N_43587);
nor U43862 (N_43862,N_43538,N_43717);
and U43863 (N_43863,N_43669,N_43537);
and U43864 (N_43864,N_43615,N_43635);
nor U43865 (N_43865,N_43721,N_43540);
nor U43866 (N_43866,N_43573,N_43604);
nor U43867 (N_43867,N_43551,N_43746);
or U43868 (N_43868,N_43724,N_43691);
and U43869 (N_43869,N_43738,N_43521);
xor U43870 (N_43870,N_43618,N_43737);
nor U43871 (N_43871,N_43528,N_43723);
nand U43872 (N_43872,N_43559,N_43518);
or U43873 (N_43873,N_43574,N_43548);
and U43874 (N_43874,N_43681,N_43636);
and U43875 (N_43875,N_43521,N_43667);
or U43876 (N_43876,N_43621,N_43648);
xor U43877 (N_43877,N_43580,N_43640);
and U43878 (N_43878,N_43687,N_43666);
or U43879 (N_43879,N_43622,N_43636);
or U43880 (N_43880,N_43618,N_43650);
xor U43881 (N_43881,N_43627,N_43649);
nand U43882 (N_43882,N_43622,N_43529);
and U43883 (N_43883,N_43577,N_43579);
nand U43884 (N_43884,N_43513,N_43500);
or U43885 (N_43885,N_43697,N_43527);
and U43886 (N_43886,N_43611,N_43565);
or U43887 (N_43887,N_43509,N_43520);
and U43888 (N_43888,N_43691,N_43504);
or U43889 (N_43889,N_43638,N_43713);
nor U43890 (N_43890,N_43740,N_43515);
and U43891 (N_43891,N_43720,N_43669);
nand U43892 (N_43892,N_43699,N_43583);
and U43893 (N_43893,N_43593,N_43612);
and U43894 (N_43894,N_43642,N_43511);
xnor U43895 (N_43895,N_43617,N_43532);
nor U43896 (N_43896,N_43717,N_43614);
xnor U43897 (N_43897,N_43599,N_43653);
xnor U43898 (N_43898,N_43500,N_43733);
nor U43899 (N_43899,N_43500,N_43623);
nor U43900 (N_43900,N_43513,N_43624);
or U43901 (N_43901,N_43589,N_43672);
xor U43902 (N_43902,N_43591,N_43513);
xor U43903 (N_43903,N_43580,N_43639);
xnor U43904 (N_43904,N_43668,N_43716);
nor U43905 (N_43905,N_43547,N_43531);
nor U43906 (N_43906,N_43620,N_43521);
xor U43907 (N_43907,N_43551,N_43583);
and U43908 (N_43908,N_43725,N_43548);
and U43909 (N_43909,N_43553,N_43555);
or U43910 (N_43910,N_43556,N_43639);
nor U43911 (N_43911,N_43613,N_43705);
nand U43912 (N_43912,N_43562,N_43620);
nand U43913 (N_43913,N_43680,N_43746);
nor U43914 (N_43914,N_43708,N_43513);
xor U43915 (N_43915,N_43527,N_43540);
and U43916 (N_43916,N_43546,N_43603);
nand U43917 (N_43917,N_43748,N_43725);
or U43918 (N_43918,N_43613,N_43530);
and U43919 (N_43919,N_43597,N_43520);
xnor U43920 (N_43920,N_43723,N_43568);
nand U43921 (N_43921,N_43610,N_43551);
or U43922 (N_43922,N_43631,N_43623);
nand U43923 (N_43923,N_43630,N_43727);
nand U43924 (N_43924,N_43715,N_43615);
nand U43925 (N_43925,N_43729,N_43640);
or U43926 (N_43926,N_43680,N_43600);
or U43927 (N_43927,N_43537,N_43506);
nor U43928 (N_43928,N_43578,N_43508);
xnor U43929 (N_43929,N_43651,N_43639);
xnor U43930 (N_43930,N_43723,N_43629);
xnor U43931 (N_43931,N_43638,N_43691);
or U43932 (N_43932,N_43676,N_43664);
or U43933 (N_43933,N_43728,N_43742);
nor U43934 (N_43934,N_43580,N_43693);
nand U43935 (N_43935,N_43565,N_43517);
nor U43936 (N_43936,N_43691,N_43690);
or U43937 (N_43937,N_43546,N_43625);
nor U43938 (N_43938,N_43592,N_43660);
nand U43939 (N_43939,N_43670,N_43588);
nand U43940 (N_43940,N_43720,N_43673);
and U43941 (N_43941,N_43745,N_43648);
nor U43942 (N_43942,N_43695,N_43697);
nor U43943 (N_43943,N_43554,N_43585);
and U43944 (N_43944,N_43536,N_43720);
or U43945 (N_43945,N_43745,N_43578);
nor U43946 (N_43946,N_43742,N_43686);
or U43947 (N_43947,N_43694,N_43591);
or U43948 (N_43948,N_43589,N_43574);
and U43949 (N_43949,N_43618,N_43503);
or U43950 (N_43950,N_43567,N_43564);
or U43951 (N_43951,N_43602,N_43732);
nor U43952 (N_43952,N_43526,N_43710);
nor U43953 (N_43953,N_43618,N_43620);
or U43954 (N_43954,N_43684,N_43656);
and U43955 (N_43955,N_43729,N_43520);
or U43956 (N_43956,N_43589,N_43743);
nor U43957 (N_43957,N_43642,N_43594);
and U43958 (N_43958,N_43621,N_43590);
nand U43959 (N_43959,N_43510,N_43567);
xor U43960 (N_43960,N_43645,N_43654);
nor U43961 (N_43961,N_43693,N_43622);
nor U43962 (N_43962,N_43605,N_43524);
nand U43963 (N_43963,N_43505,N_43610);
xnor U43964 (N_43964,N_43593,N_43574);
or U43965 (N_43965,N_43569,N_43745);
nand U43966 (N_43966,N_43737,N_43679);
nand U43967 (N_43967,N_43708,N_43687);
nand U43968 (N_43968,N_43598,N_43731);
xor U43969 (N_43969,N_43539,N_43703);
nand U43970 (N_43970,N_43702,N_43643);
nand U43971 (N_43971,N_43511,N_43545);
and U43972 (N_43972,N_43719,N_43551);
or U43973 (N_43973,N_43513,N_43564);
nor U43974 (N_43974,N_43558,N_43509);
xnor U43975 (N_43975,N_43702,N_43534);
nor U43976 (N_43976,N_43586,N_43529);
xor U43977 (N_43977,N_43699,N_43748);
or U43978 (N_43978,N_43746,N_43687);
or U43979 (N_43979,N_43504,N_43518);
and U43980 (N_43980,N_43684,N_43631);
and U43981 (N_43981,N_43684,N_43676);
or U43982 (N_43982,N_43613,N_43741);
or U43983 (N_43983,N_43535,N_43581);
or U43984 (N_43984,N_43563,N_43513);
nor U43985 (N_43985,N_43691,N_43562);
and U43986 (N_43986,N_43676,N_43570);
nand U43987 (N_43987,N_43507,N_43555);
or U43988 (N_43988,N_43684,N_43673);
xnor U43989 (N_43989,N_43685,N_43622);
xor U43990 (N_43990,N_43504,N_43748);
and U43991 (N_43991,N_43582,N_43740);
and U43992 (N_43992,N_43528,N_43748);
xor U43993 (N_43993,N_43549,N_43734);
or U43994 (N_43994,N_43622,N_43507);
nor U43995 (N_43995,N_43546,N_43649);
nor U43996 (N_43996,N_43530,N_43612);
and U43997 (N_43997,N_43693,N_43701);
and U43998 (N_43998,N_43658,N_43747);
nand U43999 (N_43999,N_43572,N_43611);
and U44000 (N_44000,N_43959,N_43877);
nand U44001 (N_44001,N_43817,N_43908);
and U44002 (N_44002,N_43952,N_43890);
nand U44003 (N_44003,N_43963,N_43823);
and U44004 (N_44004,N_43879,N_43836);
nand U44005 (N_44005,N_43931,N_43752);
nand U44006 (N_44006,N_43770,N_43772);
nor U44007 (N_44007,N_43985,N_43843);
xnor U44008 (N_44008,N_43925,N_43809);
and U44009 (N_44009,N_43827,N_43808);
or U44010 (N_44010,N_43788,N_43926);
or U44011 (N_44011,N_43793,N_43922);
or U44012 (N_44012,N_43794,N_43833);
xnor U44013 (N_44013,N_43928,N_43927);
nor U44014 (N_44014,N_43935,N_43854);
nand U44015 (N_44015,N_43986,N_43953);
or U44016 (N_44016,N_43807,N_43870);
xnor U44017 (N_44017,N_43763,N_43914);
and U44018 (N_44018,N_43769,N_43901);
and U44019 (N_44019,N_43897,N_43797);
xor U44020 (N_44020,N_43767,N_43940);
or U44021 (N_44021,N_43891,N_43924);
nor U44022 (N_44022,N_43904,N_43838);
xnor U44023 (N_44023,N_43830,N_43791);
or U44024 (N_44024,N_43875,N_43903);
xor U44025 (N_44025,N_43937,N_43782);
nand U44026 (N_44026,N_43934,N_43810);
and U44027 (N_44027,N_43896,N_43811);
or U44028 (N_44028,N_43834,N_43846);
nor U44029 (N_44029,N_43972,N_43863);
nor U44030 (N_44030,N_43813,N_43932);
xnor U44031 (N_44031,N_43929,N_43967);
xor U44032 (N_44032,N_43961,N_43852);
or U44033 (N_44033,N_43756,N_43945);
or U44034 (N_44034,N_43910,N_43882);
nor U44035 (N_44035,N_43858,N_43885);
or U44036 (N_44036,N_43824,N_43894);
and U44037 (N_44037,N_43980,N_43857);
nor U44038 (N_44038,N_43778,N_43965);
nor U44039 (N_44039,N_43995,N_43899);
nor U44040 (N_44040,N_43977,N_43783);
nor U44041 (N_44041,N_43913,N_43835);
xnor U44042 (N_44042,N_43760,N_43888);
and U44043 (N_44043,N_43851,N_43792);
nor U44044 (N_44044,N_43774,N_43768);
or U44045 (N_44045,N_43943,N_43976);
or U44046 (N_44046,N_43765,N_43887);
nor U44047 (N_44047,N_43900,N_43873);
nor U44048 (N_44048,N_43942,N_43859);
or U44049 (N_44049,N_43975,N_43822);
xnor U44050 (N_44050,N_43821,N_43862);
or U44051 (N_44051,N_43758,N_43939);
nand U44052 (N_44052,N_43915,N_43773);
nand U44053 (N_44053,N_43969,N_43892);
nand U44054 (N_44054,N_43964,N_43856);
or U44055 (N_44055,N_43802,N_43983);
and U44056 (N_44056,N_43757,N_43991);
nor U44057 (N_44057,N_43920,N_43771);
nand U44058 (N_44058,N_43907,N_43909);
xnor U44059 (N_44059,N_43867,N_43981);
and U44060 (N_44060,N_43803,N_43849);
xor U44061 (N_44061,N_43979,N_43962);
nor U44062 (N_44062,N_43974,N_43918);
nand U44063 (N_44063,N_43855,N_43871);
nand U44064 (N_44064,N_43841,N_43801);
xnor U44065 (N_44065,N_43881,N_43831);
nor U44066 (N_44066,N_43828,N_43916);
nor U44067 (N_44067,N_43987,N_43800);
nand U44068 (N_44068,N_43820,N_43753);
nand U44069 (N_44069,N_43776,N_43826);
nand U44070 (N_44070,N_43997,N_43837);
and U44071 (N_44071,N_43805,N_43895);
or U44072 (N_44072,N_43872,N_43984);
or U44073 (N_44073,N_43750,N_43842);
or U44074 (N_44074,N_43876,N_43957);
or U44075 (N_44075,N_43777,N_43861);
nand U44076 (N_44076,N_43960,N_43886);
nor U44077 (N_44077,N_43804,N_43906);
or U44078 (N_44078,N_43951,N_43898);
or U44079 (N_44079,N_43998,N_43884);
nor U44080 (N_44080,N_43844,N_43850);
and U44081 (N_44081,N_43923,N_43847);
nand U44082 (N_44082,N_43874,N_43762);
nand U44083 (N_44083,N_43883,N_43790);
or U44084 (N_44084,N_43996,N_43795);
xor U44085 (N_44085,N_43958,N_43815);
nor U44086 (N_44086,N_43988,N_43759);
and U44087 (N_44087,N_43785,N_43912);
xnor U44088 (N_44088,N_43966,N_43866);
xor U44089 (N_44089,N_43968,N_43799);
nand U44090 (N_44090,N_43825,N_43814);
nor U44091 (N_44091,N_43950,N_43798);
nand U44092 (N_44092,N_43938,N_43919);
nor U44093 (N_44093,N_43954,N_43819);
nor U44094 (N_44094,N_43990,N_43993);
nor U44095 (N_44095,N_43973,N_43970);
nand U44096 (N_44096,N_43982,N_43880);
or U44097 (N_44097,N_43971,N_43829);
and U44098 (N_44098,N_43911,N_43947);
nor U44099 (N_44099,N_43917,N_43775);
or U44100 (N_44100,N_43839,N_43787);
xor U44101 (N_44101,N_43781,N_43806);
nor U44102 (N_44102,N_43860,N_43944);
or U44103 (N_44103,N_43978,N_43832);
or U44104 (N_44104,N_43864,N_43766);
and U44105 (N_44105,N_43789,N_43868);
xnor U44106 (N_44106,N_43812,N_43936);
and U44107 (N_44107,N_43889,N_43994);
and U44108 (N_44108,N_43946,N_43955);
nor U44109 (N_44109,N_43869,N_43754);
and U44110 (N_44110,N_43786,N_43755);
nor U44111 (N_44111,N_43779,N_43865);
and U44112 (N_44112,N_43848,N_43780);
xor U44113 (N_44113,N_43751,N_43902);
nor U44114 (N_44114,N_43796,N_43948);
or U44115 (N_44115,N_43999,N_43818);
xor U44116 (N_44116,N_43989,N_43893);
nor U44117 (N_44117,N_43933,N_43949);
and U44118 (N_44118,N_43992,N_43853);
or U44119 (N_44119,N_43840,N_43764);
nand U44120 (N_44120,N_43761,N_43921);
nand U44121 (N_44121,N_43878,N_43941);
or U44122 (N_44122,N_43930,N_43905);
or U44123 (N_44123,N_43845,N_43956);
xor U44124 (N_44124,N_43784,N_43816);
xnor U44125 (N_44125,N_43854,N_43985);
nand U44126 (N_44126,N_43936,N_43865);
or U44127 (N_44127,N_43984,N_43871);
xnor U44128 (N_44128,N_43848,N_43813);
nor U44129 (N_44129,N_43875,N_43885);
nor U44130 (N_44130,N_43936,N_43973);
nand U44131 (N_44131,N_43774,N_43890);
nor U44132 (N_44132,N_43969,N_43752);
or U44133 (N_44133,N_43822,N_43989);
or U44134 (N_44134,N_43852,N_43994);
or U44135 (N_44135,N_43925,N_43959);
and U44136 (N_44136,N_43836,N_43953);
xnor U44137 (N_44137,N_43936,N_43875);
and U44138 (N_44138,N_43957,N_43958);
xor U44139 (N_44139,N_43951,N_43857);
or U44140 (N_44140,N_43828,N_43933);
and U44141 (N_44141,N_43821,N_43930);
nor U44142 (N_44142,N_43757,N_43962);
nand U44143 (N_44143,N_43773,N_43865);
xor U44144 (N_44144,N_43890,N_43768);
nor U44145 (N_44145,N_43779,N_43927);
nor U44146 (N_44146,N_43998,N_43801);
and U44147 (N_44147,N_43840,N_43899);
and U44148 (N_44148,N_43825,N_43773);
nor U44149 (N_44149,N_43788,N_43830);
or U44150 (N_44150,N_43797,N_43966);
nor U44151 (N_44151,N_43774,N_43913);
or U44152 (N_44152,N_43852,N_43990);
or U44153 (N_44153,N_43871,N_43955);
nor U44154 (N_44154,N_43795,N_43853);
xor U44155 (N_44155,N_43942,N_43799);
nand U44156 (N_44156,N_43769,N_43812);
xnor U44157 (N_44157,N_43841,N_43959);
nor U44158 (N_44158,N_43914,N_43950);
and U44159 (N_44159,N_43802,N_43818);
nand U44160 (N_44160,N_43756,N_43908);
and U44161 (N_44161,N_43913,N_43807);
nand U44162 (N_44162,N_43943,N_43887);
and U44163 (N_44163,N_43839,N_43775);
xor U44164 (N_44164,N_43792,N_43754);
or U44165 (N_44165,N_43988,N_43786);
nor U44166 (N_44166,N_43762,N_43872);
nor U44167 (N_44167,N_43897,N_43750);
xnor U44168 (N_44168,N_43980,N_43969);
nor U44169 (N_44169,N_43764,N_43779);
nor U44170 (N_44170,N_43772,N_43915);
and U44171 (N_44171,N_43782,N_43761);
or U44172 (N_44172,N_43930,N_43901);
nand U44173 (N_44173,N_43943,N_43850);
or U44174 (N_44174,N_43823,N_43943);
xor U44175 (N_44175,N_43964,N_43980);
nor U44176 (N_44176,N_43773,N_43969);
nand U44177 (N_44177,N_43880,N_43864);
nor U44178 (N_44178,N_43861,N_43908);
nor U44179 (N_44179,N_43888,N_43829);
or U44180 (N_44180,N_43856,N_43808);
xor U44181 (N_44181,N_43962,N_43897);
and U44182 (N_44182,N_43937,N_43786);
nor U44183 (N_44183,N_43799,N_43965);
or U44184 (N_44184,N_43885,N_43976);
and U44185 (N_44185,N_43998,N_43832);
and U44186 (N_44186,N_43807,N_43899);
nor U44187 (N_44187,N_43815,N_43810);
or U44188 (N_44188,N_43987,N_43780);
nor U44189 (N_44189,N_43862,N_43799);
or U44190 (N_44190,N_43787,N_43784);
and U44191 (N_44191,N_43979,N_43867);
nor U44192 (N_44192,N_43856,N_43866);
and U44193 (N_44193,N_43897,N_43886);
nand U44194 (N_44194,N_43821,N_43819);
nand U44195 (N_44195,N_43883,N_43967);
nand U44196 (N_44196,N_43937,N_43900);
nor U44197 (N_44197,N_43934,N_43902);
and U44198 (N_44198,N_43768,N_43897);
or U44199 (N_44199,N_43807,N_43818);
and U44200 (N_44200,N_43939,N_43909);
or U44201 (N_44201,N_43874,N_43772);
nand U44202 (N_44202,N_43870,N_43955);
nand U44203 (N_44203,N_43760,N_43957);
nand U44204 (N_44204,N_43801,N_43880);
and U44205 (N_44205,N_43855,N_43988);
or U44206 (N_44206,N_43824,N_43832);
or U44207 (N_44207,N_43783,N_43999);
and U44208 (N_44208,N_43828,N_43982);
nor U44209 (N_44209,N_43912,N_43987);
nand U44210 (N_44210,N_43909,N_43931);
nand U44211 (N_44211,N_43842,N_43821);
and U44212 (N_44212,N_43756,N_43854);
nor U44213 (N_44213,N_43790,N_43933);
or U44214 (N_44214,N_43823,N_43984);
xor U44215 (N_44215,N_43860,N_43863);
and U44216 (N_44216,N_43811,N_43945);
nor U44217 (N_44217,N_43938,N_43953);
xor U44218 (N_44218,N_43818,N_43979);
or U44219 (N_44219,N_43860,N_43896);
or U44220 (N_44220,N_43841,N_43937);
nor U44221 (N_44221,N_43887,N_43968);
nand U44222 (N_44222,N_43825,N_43837);
nor U44223 (N_44223,N_43944,N_43951);
nor U44224 (N_44224,N_43967,N_43818);
and U44225 (N_44225,N_43954,N_43978);
or U44226 (N_44226,N_43873,N_43920);
and U44227 (N_44227,N_43784,N_43908);
and U44228 (N_44228,N_43893,N_43886);
nor U44229 (N_44229,N_43859,N_43806);
or U44230 (N_44230,N_43942,N_43975);
or U44231 (N_44231,N_43902,N_43890);
xnor U44232 (N_44232,N_43837,N_43770);
or U44233 (N_44233,N_43792,N_43755);
nor U44234 (N_44234,N_43800,N_43888);
xor U44235 (N_44235,N_43886,N_43828);
and U44236 (N_44236,N_43956,N_43943);
nand U44237 (N_44237,N_43868,N_43856);
or U44238 (N_44238,N_43953,N_43970);
nor U44239 (N_44239,N_43960,N_43970);
xor U44240 (N_44240,N_43877,N_43986);
nand U44241 (N_44241,N_43930,N_43825);
nand U44242 (N_44242,N_43898,N_43880);
xor U44243 (N_44243,N_43947,N_43913);
nand U44244 (N_44244,N_43932,N_43894);
or U44245 (N_44245,N_43788,N_43901);
nand U44246 (N_44246,N_43776,N_43972);
nand U44247 (N_44247,N_43911,N_43905);
nand U44248 (N_44248,N_43888,N_43823);
nand U44249 (N_44249,N_43801,N_43849);
and U44250 (N_44250,N_44189,N_44248);
or U44251 (N_44251,N_44092,N_44134);
or U44252 (N_44252,N_44119,N_44048);
or U44253 (N_44253,N_44003,N_44246);
and U44254 (N_44254,N_44074,N_44070);
and U44255 (N_44255,N_44115,N_44036);
and U44256 (N_44256,N_44133,N_44167);
nor U44257 (N_44257,N_44200,N_44208);
and U44258 (N_44258,N_44179,N_44129);
xnor U44259 (N_44259,N_44131,N_44242);
nor U44260 (N_44260,N_44053,N_44109);
and U44261 (N_44261,N_44061,N_44030);
nand U44262 (N_44262,N_44226,N_44192);
xor U44263 (N_44263,N_44060,N_44197);
or U44264 (N_44264,N_44183,N_44210);
or U44265 (N_44265,N_44148,N_44214);
xor U44266 (N_44266,N_44233,N_44076);
or U44267 (N_44267,N_44223,N_44040);
and U44268 (N_44268,N_44080,N_44161);
nor U44269 (N_44269,N_44238,N_44121);
and U44270 (N_44270,N_44169,N_44056);
xnor U44271 (N_44271,N_44237,N_44105);
nand U44272 (N_44272,N_44088,N_44178);
nand U44273 (N_44273,N_44099,N_44023);
xnor U44274 (N_44274,N_44045,N_44004);
and U44275 (N_44275,N_44173,N_44033);
nand U44276 (N_44276,N_44010,N_44151);
nand U44277 (N_44277,N_44247,N_44239);
nor U44278 (N_44278,N_44194,N_44217);
and U44279 (N_44279,N_44149,N_44145);
nand U44280 (N_44280,N_44128,N_44084);
and U44281 (N_44281,N_44155,N_44107);
or U44282 (N_44282,N_44232,N_44202);
nand U44283 (N_44283,N_44199,N_44021);
nor U44284 (N_44284,N_44042,N_44240);
nor U44285 (N_44285,N_44014,N_44142);
nand U44286 (N_44286,N_44153,N_44209);
and U44287 (N_44287,N_44012,N_44071);
or U44288 (N_44288,N_44102,N_44069);
nor U44289 (N_44289,N_44049,N_44147);
and U44290 (N_44290,N_44090,N_44245);
nand U44291 (N_44291,N_44244,N_44164);
xor U44292 (N_44292,N_44104,N_44022);
nor U44293 (N_44293,N_44018,N_44195);
xor U44294 (N_44294,N_44198,N_44124);
nor U44295 (N_44295,N_44072,N_44097);
or U44296 (N_44296,N_44028,N_44002);
nor U44297 (N_44297,N_44222,N_44039);
and U44298 (N_44298,N_44007,N_44186);
and U44299 (N_44299,N_44229,N_44083);
and U44300 (N_44300,N_44127,N_44116);
and U44301 (N_44301,N_44181,N_44228);
nor U44302 (N_44302,N_44000,N_44230);
xor U44303 (N_44303,N_44034,N_44073);
nand U44304 (N_44304,N_44137,N_44243);
and U44305 (N_44305,N_44057,N_44201);
and U44306 (N_44306,N_44035,N_44207);
xnor U44307 (N_44307,N_44086,N_44219);
nor U44308 (N_44308,N_44082,N_44130);
and U44309 (N_44309,N_44171,N_44235);
nand U44310 (N_44310,N_44011,N_44100);
nand U44311 (N_44311,N_44110,N_44132);
nand U44312 (N_44312,N_44038,N_44106);
nor U44313 (N_44313,N_44085,N_44117);
nor U44314 (N_44314,N_44170,N_44047);
or U44315 (N_44315,N_44139,N_44172);
and U44316 (N_44316,N_44087,N_44013);
and U44317 (N_44317,N_44093,N_44046);
or U44318 (N_44318,N_44188,N_44215);
nand U44319 (N_44319,N_44075,N_44234);
and U44320 (N_44320,N_44190,N_44025);
xor U44321 (N_44321,N_44096,N_44218);
xnor U44322 (N_44322,N_44043,N_44206);
and U44323 (N_44323,N_44138,N_44196);
nor U44324 (N_44324,N_44205,N_44182);
nand U44325 (N_44325,N_44236,N_44051);
or U44326 (N_44326,N_44152,N_44063);
nand U44327 (N_44327,N_44032,N_44123);
or U44328 (N_44328,N_44118,N_44135);
or U44329 (N_44329,N_44054,N_44143);
and U44330 (N_44330,N_44225,N_44091);
nor U44331 (N_44331,N_44220,N_44058);
or U44332 (N_44332,N_44185,N_44005);
and U44333 (N_44333,N_44166,N_44094);
or U44334 (N_44334,N_44211,N_44160);
or U44335 (N_44335,N_44213,N_44079);
xnor U44336 (N_44336,N_44077,N_44146);
or U44337 (N_44337,N_44156,N_44176);
nor U44338 (N_44338,N_44216,N_44017);
xor U44339 (N_44339,N_44125,N_44221);
xnor U44340 (N_44340,N_44175,N_44020);
xnor U44341 (N_44341,N_44016,N_44065);
nor U44342 (N_44342,N_44204,N_44095);
xnor U44343 (N_44343,N_44191,N_44184);
nand U44344 (N_44344,N_44067,N_44052);
nor U44345 (N_44345,N_44203,N_44024);
nor U44346 (N_44346,N_44026,N_44136);
or U44347 (N_44347,N_44019,N_44108);
and U44348 (N_44348,N_44029,N_44168);
or U44349 (N_44349,N_44006,N_44141);
and U44350 (N_44350,N_44174,N_44098);
nor U44351 (N_44351,N_44177,N_44111);
nand U44352 (N_44352,N_44224,N_44154);
nor U44353 (N_44353,N_44180,N_44120);
nand U44354 (N_44354,N_44081,N_44044);
xnor U44355 (N_44355,N_44187,N_44140);
and U44356 (N_44356,N_44068,N_44031);
or U44357 (N_44357,N_44157,N_44050);
nor U44358 (N_44358,N_44103,N_44126);
nand U44359 (N_44359,N_44163,N_44008);
and U44360 (N_44360,N_44037,N_44101);
xor U44361 (N_44361,N_44078,N_44015);
xor U44362 (N_44362,N_44041,N_44162);
or U44363 (N_44363,N_44001,N_44122);
xor U44364 (N_44364,N_44064,N_44165);
nand U44365 (N_44365,N_44227,N_44158);
xnor U44366 (N_44366,N_44150,N_44009);
nor U44367 (N_44367,N_44193,N_44159);
or U44368 (N_44368,N_44055,N_44089);
and U44369 (N_44369,N_44112,N_44066);
nand U44370 (N_44370,N_44062,N_44212);
nor U44371 (N_44371,N_44249,N_44113);
xor U44372 (N_44372,N_44144,N_44027);
or U44373 (N_44373,N_44114,N_44241);
nor U44374 (N_44374,N_44059,N_44231);
or U44375 (N_44375,N_44196,N_44164);
xor U44376 (N_44376,N_44043,N_44240);
nor U44377 (N_44377,N_44097,N_44173);
or U44378 (N_44378,N_44191,N_44128);
or U44379 (N_44379,N_44140,N_44152);
and U44380 (N_44380,N_44128,N_44122);
and U44381 (N_44381,N_44120,N_44024);
xor U44382 (N_44382,N_44005,N_44021);
nand U44383 (N_44383,N_44117,N_44038);
nor U44384 (N_44384,N_44180,N_44234);
nand U44385 (N_44385,N_44197,N_44147);
nand U44386 (N_44386,N_44025,N_44093);
or U44387 (N_44387,N_44046,N_44135);
nand U44388 (N_44388,N_44170,N_44085);
nand U44389 (N_44389,N_44168,N_44153);
nand U44390 (N_44390,N_44106,N_44167);
nor U44391 (N_44391,N_44106,N_44123);
and U44392 (N_44392,N_44218,N_44137);
nor U44393 (N_44393,N_44051,N_44008);
and U44394 (N_44394,N_44224,N_44090);
nand U44395 (N_44395,N_44010,N_44241);
xor U44396 (N_44396,N_44188,N_44098);
nor U44397 (N_44397,N_44157,N_44015);
or U44398 (N_44398,N_44094,N_44013);
or U44399 (N_44399,N_44127,N_44005);
nand U44400 (N_44400,N_44225,N_44178);
or U44401 (N_44401,N_44246,N_44179);
xnor U44402 (N_44402,N_44240,N_44104);
nor U44403 (N_44403,N_44208,N_44158);
nand U44404 (N_44404,N_44030,N_44144);
nor U44405 (N_44405,N_44098,N_44033);
or U44406 (N_44406,N_44186,N_44178);
nand U44407 (N_44407,N_44202,N_44168);
or U44408 (N_44408,N_44007,N_44139);
nand U44409 (N_44409,N_44243,N_44110);
and U44410 (N_44410,N_44228,N_44089);
xor U44411 (N_44411,N_44109,N_44093);
and U44412 (N_44412,N_44220,N_44188);
nand U44413 (N_44413,N_44135,N_44074);
xor U44414 (N_44414,N_44218,N_44138);
and U44415 (N_44415,N_44248,N_44171);
nor U44416 (N_44416,N_44229,N_44234);
xnor U44417 (N_44417,N_44023,N_44018);
xnor U44418 (N_44418,N_44016,N_44149);
or U44419 (N_44419,N_44166,N_44207);
nand U44420 (N_44420,N_44249,N_44162);
xnor U44421 (N_44421,N_44068,N_44056);
xor U44422 (N_44422,N_44194,N_44037);
xnor U44423 (N_44423,N_44159,N_44227);
and U44424 (N_44424,N_44095,N_44044);
nand U44425 (N_44425,N_44223,N_44181);
xor U44426 (N_44426,N_44109,N_44240);
nor U44427 (N_44427,N_44138,N_44121);
nand U44428 (N_44428,N_44033,N_44175);
nand U44429 (N_44429,N_44242,N_44125);
and U44430 (N_44430,N_44091,N_44055);
nand U44431 (N_44431,N_44006,N_44173);
xor U44432 (N_44432,N_44202,N_44240);
and U44433 (N_44433,N_44023,N_44169);
nor U44434 (N_44434,N_44178,N_44026);
nand U44435 (N_44435,N_44080,N_44084);
or U44436 (N_44436,N_44020,N_44195);
and U44437 (N_44437,N_44178,N_44002);
xor U44438 (N_44438,N_44149,N_44108);
and U44439 (N_44439,N_44144,N_44172);
and U44440 (N_44440,N_44138,N_44099);
nand U44441 (N_44441,N_44009,N_44075);
nor U44442 (N_44442,N_44183,N_44179);
nand U44443 (N_44443,N_44121,N_44110);
and U44444 (N_44444,N_44229,N_44060);
or U44445 (N_44445,N_44224,N_44142);
xor U44446 (N_44446,N_44154,N_44235);
and U44447 (N_44447,N_44237,N_44213);
or U44448 (N_44448,N_44083,N_44133);
nand U44449 (N_44449,N_44129,N_44082);
or U44450 (N_44450,N_44012,N_44073);
nor U44451 (N_44451,N_44197,N_44052);
nand U44452 (N_44452,N_44224,N_44180);
nand U44453 (N_44453,N_44067,N_44234);
or U44454 (N_44454,N_44070,N_44115);
and U44455 (N_44455,N_44077,N_44244);
or U44456 (N_44456,N_44067,N_44197);
nor U44457 (N_44457,N_44028,N_44052);
nand U44458 (N_44458,N_44185,N_44023);
or U44459 (N_44459,N_44241,N_44139);
xnor U44460 (N_44460,N_44130,N_44212);
or U44461 (N_44461,N_44155,N_44017);
and U44462 (N_44462,N_44007,N_44015);
and U44463 (N_44463,N_44197,N_44189);
xnor U44464 (N_44464,N_44006,N_44244);
nor U44465 (N_44465,N_44190,N_44070);
nor U44466 (N_44466,N_44218,N_44205);
xor U44467 (N_44467,N_44086,N_44000);
or U44468 (N_44468,N_44160,N_44049);
or U44469 (N_44469,N_44161,N_44246);
nand U44470 (N_44470,N_44219,N_44047);
nand U44471 (N_44471,N_44148,N_44132);
nand U44472 (N_44472,N_44221,N_44138);
nor U44473 (N_44473,N_44234,N_44157);
nand U44474 (N_44474,N_44060,N_44125);
and U44475 (N_44475,N_44077,N_44058);
nand U44476 (N_44476,N_44229,N_44093);
or U44477 (N_44477,N_44101,N_44094);
or U44478 (N_44478,N_44197,N_44210);
xor U44479 (N_44479,N_44187,N_44083);
and U44480 (N_44480,N_44108,N_44229);
nand U44481 (N_44481,N_44219,N_44185);
nand U44482 (N_44482,N_44099,N_44144);
nand U44483 (N_44483,N_44028,N_44193);
nand U44484 (N_44484,N_44241,N_44106);
nand U44485 (N_44485,N_44215,N_44132);
and U44486 (N_44486,N_44138,N_44162);
and U44487 (N_44487,N_44227,N_44003);
nor U44488 (N_44488,N_44087,N_44035);
nor U44489 (N_44489,N_44121,N_44061);
xnor U44490 (N_44490,N_44052,N_44016);
xnor U44491 (N_44491,N_44099,N_44227);
and U44492 (N_44492,N_44023,N_44027);
nand U44493 (N_44493,N_44039,N_44114);
and U44494 (N_44494,N_44055,N_44240);
and U44495 (N_44495,N_44158,N_44190);
nand U44496 (N_44496,N_44020,N_44035);
nand U44497 (N_44497,N_44245,N_44080);
or U44498 (N_44498,N_44085,N_44073);
nand U44499 (N_44499,N_44035,N_44078);
nor U44500 (N_44500,N_44283,N_44343);
and U44501 (N_44501,N_44256,N_44304);
and U44502 (N_44502,N_44417,N_44345);
nand U44503 (N_44503,N_44379,N_44481);
xnor U44504 (N_44504,N_44468,N_44255);
and U44505 (N_44505,N_44313,N_44350);
nor U44506 (N_44506,N_44431,N_44428);
nand U44507 (N_44507,N_44399,N_44330);
or U44508 (N_44508,N_44465,N_44405);
or U44509 (N_44509,N_44294,N_44496);
nand U44510 (N_44510,N_44418,N_44480);
nor U44511 (N_44511,N_44498,N_44309);
nand U44512 (N_44512,N_44329,N_44288);
nor U44513 (N_44513,N_44378,N_44412);
nor U44514 (N_44514,N_44395,N_44293);
nand U44515 (N_44515,N_44447,N_44254);
and U44516 (N_44516,N_44339,N_44440);
or U44517 (N_44517,N_44367,N_44272);
nor U44518 (N_44518,N_44344,N_44289);
or U44519 (N_44519,N_44355,N_44260);
nor U44520 (N_44520,N_44491,N_44466);
nand U44521 (N_44521,N_44411,N_44450);
and U44522 (N_44522,N_44432,N_44443);
or U44523 (N_44523,N_44348,N_44451);
nand U44524 (N_44524,N_44323,N_44453);
and U44525 (N_44525,N_44285,N_44427);
or U44526 (N_44526,N_44274,N_44259);
nor U44527 (N_44527,N_44488,N_44499);
nand U44528 (N_44528,N_44403,N_44277);
nor U44529 (N_44529,N_44384,N_44271);
and U44530 (N_44530,N_44300,N_44360);
xor U44531 (N_44531,N_44477,N_44317);
xnor U44532 (N_44532,N_44448,N_44335);
nor U44533 (N_44533,N_44484,N_44486);
and U44534 (N_44534,N_44327,N_44490);
nand U44535 (N_44535,N_44303,N_44333);
and U44536 (N_44536,N_44485,N_44322);
nand U44537 (N_44537,N_44365,N_44337);
or U44538 (N_44538,N_44470,N_44471);
nor U44539 (N_44539,N_44456,N_44282);
nor U44540 (N_44540,N_44262,N_44364);
nand U44541 (N_44541,N_44420,N_44297);
xnor U44542 (N_44542,N_44354,N_44483);
and U44543 (N_44543,N_44280,N_44353);
or U44544 (N_44544,N_44454,N_44316);
and U44545 (N_44545,N_44479,N_44253);
or U44546 (N_44546,N_44352,N_44371);
or U44547 (N_44547,N_44299,N_44381);
xnor U44548 (N_44548,N_44325,N_44269);
nor U44549 (N_44549,N_44407,N_44312);
or U44550 (N_44550,N_44292,N_44263);
and U44551 (N_44551,N_44425,N_44482);
and U44552 (N_44552,N_44424,N_44287);
nand U44553 (N_44553,N_44409,N_44359);
nor U44554 (N_44554,N_44445,N_44332);
nor U44555 (N_44555,N_44318,N_44497);
nand U44556 (N_44556,N_44326,N_44494);
and U44557 (N_44557,N_44415,N_44388);
or U44558 (N_44558,N_44434,N_44389);
nor U44559 (N_44559,N_44422,N_44438);
and U44560 (N_44560,N_44314,N_44449);
and U44561 (N_44561,N_44446,N_44433);
nand U44562 (N_44562,N_44268,N_44386);
nand U44563 (N_44563,N_44338,N_44377);
nand U44564 (N_44564,N_44492,N_44306);
xnor U44565 (N_44565,N_44398,N_44375);
nand U44566 (N_44566,N_44401,N_44489);
xnor U44567 (N_44567,N_44475,N_44429);
xor U44568 (N_44568,N_44495,N_44387);
xnor U44569 (N_44569,N_44402,N_44279);
xnor U44570 (N_44570,N_44426,N_44290);
xor U44571 (N_44571,N_44362,N_44472);
and U44572 (N_44572,N_44408,N_44382);
nor U44573 (N_44573,N_44473,N_44436);
or U44574 (N_44574,N_44423,N_44455);
or U44575 (N_44575,N_44257,N_44459);
nand U44576 (N_44576,N_44410,N_44394);
and U44577 (N_44577,N_44462,N_44286);
xor U44578 (N_44578,N_44307,N_44273);
xnor U44579 (N_44579,N_44474,N_44342);
xnor U44580 (N_44580,N_44310,N_44349);
nor U44581 (N_44581,N_44464,N_44369);
or U44582 (N_44582,N_44311,N_44376);
nand U44583 (N_44583,N_44328,N_44366);
and U44584 (N_44584,N_44457,N_44264);
nand U44585 (N_44585,N_44298,N_44356);
or U44586 (N_44586,N_44251,N_44467);
xnor U44587 (N_44587,N_44258,N_44295);
nand U44588 (N_44588,N_44458,N_44331);
and U44589 (N_44589,N_44324,N_44421);
nand U44590 (N_44590,N_44266,N_44373);
xor U44591 (N_44591,N_44390,N_44361);
and U44592 (N_44592,N_44270,N_44250);
xnor U44593 (N_44593,N_44275,N_44393);
and U44594 (N_44594,N_44351,N_44452);
or U44595 (N_44595,N_44441,N_44414);
xnor U44596 (N_44596,N_44374,N_44302);
nand U44597 (N_44597,N_44276,N_44261);
xor U44598 (N_44598,N_44476,N_44340);
or U44599 (N_44599,N_44397,N_44413);
and U44600 (N_44600,N_44308,N_44278);
xnor U44601 (N_44601,N_44370,N_44334);
nor U44602 (N_44602,N_44320,N_44493);
nand U44603 (N_44603,N_44315,N_44444);
xor U44604 (N_44604,N_44430,N_44460);
xor U44605 (N_44605,N_44358,N_44442);
nor U44606 (N_44606,N_44291,N_44487);
and U44607 (N_44607,N_44346,N_44461);
or U44608 (N_44608,N_44336,N_44305);
and U44609 (N_44609,N_44296,N_44435);
and U44610 (N_44610,N_44372,N_44284);
or U44611 (N_44611,N_44368,N_44419);
nor U44612 (N_44612,N_44463,N_44383);
and U44613 (N_44613,N_44347,N_44406);
xor U44614 (N_44614,N_44439,N_44469);
or U44615 (N_44615,N_44357,N_44380);
or U44616 (N_44616,N_44437,N_44301);
nor U44617 (N_44617,N_44391,N_44281);
nor U44618 (N_44618,N_44319,N_44478);
xnor U44619 (N_44619,N_44416,N_44265);
nand U44620 (N_44620,N_44392,N_44321);
nor U44621 (N_44621,N_44396,N_44400);
xor U44622 (N_44622,N_44385,N_44267);
and U44623 (N_44623,N_44404,N_44363);
and U44624 (N_44624,N_44341,N_44252);
or U44625 (N_44625,N_44337,N_44318);
or U44626 (N_44626,N_44422,N_44498);
xnor U44627 (N_44627,N_44259,N_44382);
xnor U44628 (N_44628,N_44362,N_44465);
xor U44629 (N_44629,N_44288,N_44353);
or U44630 (N_44630,N_44377,N_44459);
or U44631 (N_44631,N_44304,N_44356);
and U44632 (N_44632,N_44327,N_44395);
nor U44633 (N_44633,N_44429,N_44336);
and U44634 (N_44634,N_44468,N_44482);
nor U44635 (N_44635,N_44324,N_44358);
or U44636 (N_44636,N_44344,N_44466);
and U44637 (N_44637,N_44476,N_44331);
nand U44638 (N_44638,N_44283,N_44408);
xnor U44639 (N_44639,N_44271,N_44421);
and U44640 (N_44640,N_44307,N_44287);
nor U44641 (N_44641,N_44473,N_44443);
or U44642 (N_44642,N_44373,N_44478);
or U44643 (N_44643,N_44494,N_44414);
xnor U44644 (N_44644,N_44387,N_44423);
nor U44645 (N_44645,N_44364,N_44444);
nor U44646 (N_44646,N_44439,N_44332);
xnor U44647 (N_44647,N_44459,N_44260);
or U44648 (N_44648,N_44372,N_44417);
or U44649 (N_44649,N_44430,N_44481);
or U44650 (N_44650,N_44355,N_44266);
xnor U44651 (N_44651,N_44309,N_44466);
or U44652 (N_44652,N_44454,N_44318);
or U44653 (N_44653,N_44437,N_44486);
xor U44654 (N_44654,N_44279,N_44342);
and U44655 (N_44655,N_44476,N_44485);
or U44656 (N_44656,N_44326,N_44464);
nor U44657 (N_44657,N_44416,N_44316);
nand U44658 (N_44658,N_44496,N_44279);
and U44659 (N_44659,N_44270,N_44416);
and U44660 (N_44660,N_44351,N_44250);
xnor U44661 (N_44661,N_44252,N_44308);
and U44662 (N_44662,N_44337,N_44394);
xor U44663 (N_44663,N_44273,N_44281);
or U44664 (N_44664,N_44402,N_44331);
xor U44665 (N_44665,N_44489,N_44403);
and U44666 (N_44666,N_44409,N_44387);
xnor U44667 (N_44667,N_44378,N_44470);
xor U44668 (N_44668,N_44258,N_44349);
or U44669 (N_44669,N_44467,N_44465);
xor U44670 (N_44670,N_44368,N_44468);
and U44671 (N_44671,N_44417,N_44446);
nor U44672 (N_44672,N_44262,N_44477);
or U44673 (N_44673,N_44287,N_44314);
nor U44674 (N_44674,N_44272,N_44389);
nor U44675 (N_44675,N_44280,N_44383);
nor U44676 (N_44676,N_44306,N_44272);
or U44677 (N_44677,N_44412,N_44417);
or U44678 (N_44678,N_44254,N_44265);
xnor U44679 (N_44679,N_44357,N_44360);
xnor U44680 (N_44680,N_44402,N_44287);
xnor U44681 (N_44681,N_44260,N_44336);
or U44682 (N_44682,N_44436,N_44456);
and U44683 (N_44683,N_44499,N_44321);
and U44684 (N_44684,N_44407,N_44256);
nand U44685 (N_44685,N_44477,N_44305);
and U44686 (N_44686,N_44444,N_44284);
xnor U44687 (N_44687,N_44295,N_44476);
or U44688 (N_44688,N_44361,N_44462);
nand U44689 (N_44689,N_44422,N_44409);
xnor U44690 (N_44690,N_44457,N_44300);
nand U44691 (N_44691,N_44448,N_44468);
nor U44692 (N_44692,N_44285,N_44435);
nand U44693 (N_44693,N_44388,N_44469);
nor U44694 (N_44694,N_44301,N_44312);
nor U44695 (N_44695,N_44370,N_44306);
nand U44696 (N_44696,N_44308,N_44445);
or U44697 (N_44697,N_44302,N_44481);
nor U44698 (N_44698,N_44352,N_44350);
xnor U44699 (N_44699,N_44379,N_44495);
or U44700 (N_44700,N_44406,N_44475);
xnor U44701 (N_44701,N_44466,N_44498);
nand U44702 (N_44702,N_44342,N_44365);
and U44703 (N_44703,N_44430,N_44413);
nor U44704 (N_44704,N_44289,N_44357);
nand U44705 (N_44705,N_44324,N_44381);
xnor U44706 (N_44706,N_44262,N_44379);
nor U44707 (N_44707,N_44260,N_44380);
nand U44708 (N_44708,N_44283,N_44357);
or U44709 (N_44709,N_44472,N_44413);
nand U44710 (N_44710,N_44378,N_44380);
nor U44711 (N_44711,N_44297,N_44494);
nand U44712 (N_44712,N_44406,N_44400);
nor U44713 (N_44713,N_44446,N_44448);
xnor U44714 (N_44714,N_44419,N_44470);
or U44715 (N_44715,N_44285,N_44347);
and U44716 (N_44716,N_44339,N_44338);
nor U44717 (N_44717,N_44401,N_44492);
and U44718 (N_44718,N_44351,N_44257);
nand U44719 (N_44719,N_44432,N_44401);
and U44720 (N_44720,N_44460,N_44303);
and U44721 (N_44721,N_44324,N_44477);
nor U44722 (N_44722,N_44441,N_44310);
nand U44723 (N_44723,N_44369,N_44281);
nor U44724 (N_44724,N_44266,N_44296);
or U44725 (N_44725,N_44455,N_44400);
xor U44726 (N_44726,N_44441,N_44367);
or U44727 (N_44727,N_44349,N_44305);
and U44728 (N_44728,N_44383,N_44430);
xnor U44729 (N_44729,N_44322,N_44378);
and U44730 (N_44730,N_44452,N_44366);
xor U44731 (N_44731,N_44284,N_44475);
xnor U44732 (N_44732,N_44456,N_44281);
nand U44733 (N_44733,N_44284,N_44410);
and U44734 (N_44734,N_44367,N_44394);
or U44735 (N_44735,N_44336,N_44495);
nor U44736 (N_44736,N_44369,N_44328);
nand U44737 (N_44737,N_44492,N_44293);
or U44738 (N_44738,N_44425,N_44312);
and U44739 (N_44739,N_44464,N_44333);
nor U44740 (N_44740,N_44485,N_44403);
or U44741 (N_44741,N_44473,N_44376);
xor U44742 (N_44742,N_44491,N_44262);
nand U44743 (N_44743,N_44384,N_44391);
and U44744 (N_44744,N_44305,N_44485);
nand U44745 (N_44745,N_44274,N_44290);
nor U44746 (N_44746,N_44439,N_44430);
nand U44747 (N_44747,N_44397,N_44482);
xor U44748 (N_44748,N_44394,N_44439);
nand U44749 (N_44749,N_44298,N_44410);
nand U44750 (N_44750,N_44536,N_44593);
and U44751 (N_44751,N_44529,N_44736);
nand U44752 (N_44752,N_44683,N_44570);
nand U44753 (N_44753,N_44578,N_44638);
or U44754 (N_44754,N_44547,N_44707);
xnor U44755 (N_44755,N_44675,N_44558);
and U44756 (N_44756,N_44733,N_44676);
nor U44757 (N_44757,N_44711,N_44620);
and U44758 (N_44758,N_44745,N_44521);
or U44759 (N_44759,N_44662,N_44660);
xor U44760 (N_44760,N_44746,N_44514);
xor U44761 (N_44761,N_44621,N_44569);
or U44762 (N_44762,N_44664,N_44566);
nor U44763 (N_44763,N_44627,N_44618);
nor U44764 (N_44764,N_44568,N_44582);
nor U44765 (N_44765,N_44518,N_44643);
or U44766 (N_44766,N_44614,N_44712);
nand U44767 (N_44767,N_44599,N_44647);
nand U44768 (N_44768,N_44500,N_44623);
nor U44769 (N_44769,N_44598,N_44653);
nand U44770 (N_44770,N_44549,N_44531);
and U44771 (N_44771,N_44523,N_44553);
or U44772 (N_44772,N_44505,N_44648);
nor U44773 (N_44773,N_44586,N_44655);
and U44774 (N_44774,N_44693,N_44677);
xnor U44775 (N_44775,N_44635,N_44741);
xnor U44776 (N_44776,N_44510,N_44530);
nor U44777 (N_44777,N_44613,N_44674);
or U44778 (N_44778,N_44658,N_44645);
or U44779 (N_44779,N_44519,N_44555);
nor U44780 (N_44780,N_44633,N_44603);
or U44781 (N_44781,N_44744,N_44665);
nor U44782 (N_44782,N_44546,N_44526);
nand U44783 (N_44783,N_44737,N_44626);
nand U44784 (N_44784,N_44577,N_44564);
nand U44785 (N_44785,N_44628,N_44605);
or U44786 (N_44786,N_44720,N_44501);
nand U44787 (N_44787,N_44701,N_44503);
nor U44788 (N_44788,N_44601,N_44739);
nor U44789 (N_44789,N_44725,N_44571);
xor U44790 (N_44790,N_44583,N_44592);
and U44791 (N_44791,N_44612,N_44574);
nand U44792 (N_44792,N_44535,N_44669);
and U44793 (N_44793,N_44650,N_44509);
or U44794 (N_44794,N_44636,N_44522);
xnor U44795 (N_44795,N_44600,N_44727);
nor U44796 (N_44796,N_44715,N_44532);
nor U44797 (N_44797,N_44515,N_44731);
or U44798 (N_44798,N_44534,N_44579);
and U44799 (N_44799,N_44575,N_44724);
xor U44800 (N_44800,N_44584,N_44559);
xor U44801 (N_44801,N_44723,N_44544);
and U44802 (N_44802,N_44630,N_44670);
or U44803 (N_44803,N_44685,N_44661);
nor U44804 (N_44804,N_44691,N_44730);
xnor U44805 (N_44805,N_44719,N_44668);
or U44806 (N_44806,N_44710,N_44550);
xor U44807 (N_44807,N_44507,N_44610);
or U44808 (N_44808,N_44651,N_44709);
and U44809 (N_44809,N_44562,N_44684);
and U44810 (N_44810,N_44732,N_44697);
or U44811 (N_44811,N_44690,N_44702);
or U44812 (N_44812,N_44513,N_44718);
and U44813 (N_44813,N_44556,N_44649);
nand U44814 (N_44814,N_44572,N_44615);
nor U44815 (N_44815,N_44657,N_44573);
or U44816 (N_44816,N_44588,N_44540);
nor U44817 (N_44817,N_44704,N_44678);
nor U44818 (N_44818,N_44703,N_44680);
or U44819 (N_44819,N_44742,N_44671);
or U44820 (N_44820,N_44672,N_44548);
or U44821 (N_44821,N_44506,N_44517);
and U44822 (N_44822,N_44524,N_44642);
and U44823 (N_44823,N_44692,N_44595);
and U44824 (N_44824,N_44644,N_44525);
and U44825 (N_44825,N_44698,N_44729);
nor U44826 (N_44826,N_44726,N_44551);
nor U44827 (N_44827,N_44576,N_44625);
nand U44828 (N_44828,N_44748,N_44622);
nand U44829 (N_44829,N_44689,N_44616);
and U44830 (N_44830,N_44713,N_44656);
and U44831 (N_44831,N_44594,N_44735);
or U44832 (N_44832,N_44502,N_44527);
xor U44833 (N_44833,N_44688,N_44663);
nand U44834 (N_44834,N_44596,N_44541);
nor U44835 (N_44835,N_44717,N_44696);
xnor U44836 (N_44836,N_44722,N_44667);
nand U44837 (N_44837,N_44587,N_44740);
or U44838 (N_44838,N_44659,N_44539);
or U44839 (N_44839,N_44557,N_44542);
and U44840 (N_44840,N_44654,N_44552);
xnor U44841 (N_44841,N_44631,N_44609);
nand U44842 (N_44842,N_44567,N_44511);
and U44843 (N_44843,N_44516,N_44581);
nand U44844 (N_44844,N_44607,N_44561);
nor U44845 (N_44845,N_44589,N_44560);
or U44846 (N_44846,N_44646,N_44512);
and U44847 (N_44847,N_44528,N_44632);
nand U44848 (N_44848,N_44624,N_44545);
nand U44849 (N_44849,N_44641,N_44714);
or U44850 (N_44850,N_44679,N_44619);
nand U44851 (N_44851,N_44695,N_44694);
xor U44852 (N_44852,N_44743,N_44682);
xnor U44853 (N_44853,N_44591,N_44716);
nor U44854 (N_44854,N_44687,N_44590);
xnor U44855 (N_44855,N_44681,N_44520);
xnor U44856 (N_44856,N_44673,N_44734);
xor U44857 (N_44857,N_44639,N_44606);
or U44858 (N_44858,N_44700,N_44634);
or U44859 (N_44859,N_44554,N_44597);
xor U44860 (N_44860,N_44604,N_44533);
or U44861 (N_44861,N_44611,N_44580);
nand U44862 (N_44862,N_44666,N_44602);
or U44863 (N_44863,N_44637,N_44537);
nor U44864 (N_44864,N_44705,N_44504);
or U44865 (N_44865,N_44728,N_44585);
nor U44866 (N_44866,N_44563,N_44617);
or U44867 (N_44867,N_44686,N_44640);
and U44868 (N_44868,N_44543,N_44738);
and U44869 (N_44869,N_44708,N_44706);
xnor U44870 (N_44870,N_44652,N_44508);
and U44871 (N_44871,N_44565,N_44629);
nor U44872 (N_44872,N_44538,N_44608);
and U44873 (N_44873,N_44721,N_44699);
nor U44874 (N_44874,N_44749,N_44747);
and U44875 (N_44875,N_44684,N_44561);
xor U44876 (N_44876,N_44724,N_44640);
or U44877 (N_44877,N_44696,N_44529);
nand U44878 (N_44878,N_44563,N_44676);
xnor U44879 (N_44879,N_44571,N_44684);
xnor U44880 (N_44880,N_44564,N_44600);
and U44881 (N_44881,N_44683,N_44529);
and U44882 (N_44882,N_44536,N_44541);
nor U44883 (N_44883,N_44507,N_44657);
nor U44884 (N_44884,N_44645,N_44522);
and U44885 (N_44885,N_44509,N_44687);
xnor U44886 (N_44886,N_44743,N_44607);
nand U44887 (N_44887,N_44743,N_44565);
or U44888 (N_44888,N_44571,N_44740);
nand U44889 (N_44889,N_44601,N_44501);
nor U44890 (N_44890,N_44540,N_44600);
and U44891 (N_44891,N_44541,N_44668);
and U44892 (N_44892,N_44705,N_44569);
nor U44893 (N_44893,N_44713,N_44514);
xor U44894 (N_44894,N_44746,N_44691);
nand U44895 (N_44895,N_44675,N_44655);
and U44896 (N_44896,N_44516,N_44680);
xor U44897 (N_44897,N_44554,N_44564);
xor U44898 (N_44898,N_44579,N_44549);
nand U44899 (N_44899,N_44735,N_44704);
or U44900 (N_44900,N_44548,N_44663);
xor U44901 (N_44901,N_44509,N_44748);
and U44902 (N_44902,N_44571,N_44565);
nor U44903 (N_44903,N_44676,N_44514);
nand U44904 (N_44904,N_44733,N_44703);
and U44905 (N_44905,N_44635,N_44522);
or U44906 (N_44906,N_44584,N_44689);
or U44907 (N_44907,N_44501,N_44607);
nand U44908 (N_44908,N_44727,N_44527);
nor U44909 (N_44909,N_44707,N_44507);
and U44910 (N_44910,N_44603,N_44652);
xnor U44911 (N_44911,N_44609,N_44563);
nand U44912 (N_44912,N_44661,N_44648);
xnor U44913 (N_44913,N_44749,N_44659);
nand U44914 (N_44914,N_44544,N_44508);
xnor U44915 (N_44915,N_44669,N_44561);
nor U44916 (N_44916,N_44715,N_44530);
xor U44917 (N_44917,N_44688,N_44687);
nand U44918 (N_44918,N_44569,N_44582);
nor U44919 (N_44919,N_44698,N_44651);
nor U44920 (N_44920,N_44734,N_44652);
or U44921 (N_44921,N_44742,N_44591);
and U44922 (N_44922,N_44722,N_44725);
nand U44923 (N_44923,N_44657,N_44702);
xor U44924 (N_44924,N_44667,N_44663);
and U44925 (N_44925,N_44512,N_44609);
nand U44926 (N_44926,N_44554,N_44704);
xor U44927 (N_44927,N_44742,N_44520);
xnor U44928 (N_44928,N_44591,N_44644);
nand U44929 (N_44929,N_44571,N_44587);
and U44930 (N_44930,N_44613,N_44618);
and U44931 (N_44931,N_44665,N_44575);
nor U44932 (N_44932,N_44539,N_44567);
or U44933 (N_44933,N_44550,N_44556);
or U44934 (N_44934,N_44704,N_44626);
and U44935 (N_44935,N_44514,N_44525);
nor U44936 (N_44936,N_44516,N_44531);
and U44937 (N_44937,N_44559,N_44649);
xnor U44938 (N_44938,N_44592,N_44555);
xor U44939 (N_44939,N_44703,N_44611);
or U44940 (N_44940,N_44724,N_44728);
nor U44941 (N_44941,N_44726,N_44643);
xnor U44942 (N_44942,N_44598,N_44524);
or U44943 (N_44943,N_44545,N_44587);
nor U44944 (N_44944,N_44575,N_44504);
nand U44945 (N_44945,N_44706,N_44699);
and U44946 (N_44946,N_44543,N_44718);
or U44947 (N_44947,N_44590,N_44588);
nor U44948 (N_44948,N_44593,N_44564);
xor U44949 (N_44949,N_44610,N_44552);
nor U44950 (N_44950,N_44605,N_44507);
and U44951 (N_44951,N_44584,N_44734);
xor U44952 (N_44952,N_44731,N_44595);
nand U44953 (N_44953,N_44600,N_44615);
nand U44954 (N_44954,N_44509,N_44575);
and U44955 (N_44955,N_44602,N_44627);
and U44956 (N_44956,N_44608,N_44559);
or U44957 (N_44957,N_44618,N_44533);
nand U44958 (N_44958,N_44747,N_44706);
xnor U44959 (N_44959,N_44701,N_44709);
or U44960 (N_44960,N_44640,N_44558);
nand U44961 (N_44961,N_44544,N_44736);
nor U44962 (N_44962,N_44652,N_44630);
nand U44963 (N_44963,N_44568,N_44649);
nand U44964 (N_44964,N_44741,N_44734);
and U44965 (N_44965,N_44638,N_44705);
nor U44966 (N_44966,N_44677,N_44617);
xor U44967 (N_44967,N_44702,N_44635);
or U44968 (N_44968,N_44544,N_44534);
nand U44969 (N_44969,N_44731,N_44635);
xnor U44970 (N_44970,N_44690,N_44584);
nor U44971 (N_44971,N_44732,N_44715);
nand U44972 (N_44972,N_44550,N_44547);
nand U44973 (N_44973,N_44652,N_44657);
or U44974 (N_44974,N_44555,N_44619);
or U44975 (N_44975,N_44730,N_44630);
nor U44976 (N_44976,N_44500,N_44731);
nand U44977 (N_44977,N_44677,N_44579);
nor U44978 (N_44978,N_44558,N_44631);
nand U44979 (N_44979,N_44703,N_44540);
xor U44980 (N_44980,N_44647,N_44637);
xor U44981 (N_44981,N_44652,N_44505);
and U44982 (N_44982,N_44660,N_44681);
or U44983 (N_44983,N_44635,N_44546);
and U44984 (N_44984,N_44703,N_44515);
nor U44985 (N_44985,N_44548,N_44525);
and U44986 (N_44986,N_44501,N_44669);
or U44987 (N_44987,N_44686,N_44519);
or U44988 (N_44988,N_44569,N_44596);
and U44989 (N_44989,N_44619,N_44598);
or U44990 (N_44990,N_44579,N_44504);
xor U44991 (N_44991,N_44691,N_44559);
and U44992 (N_44992,N_44589,N_44699);
and U44993 (N_44993,N_44688,N_44694);
xor U44994 (N_44994,N_44637,N_44560);
and U44995 (N_44995,N_44621,N_44653);
xor U44996 (N_44996,N_44685,N_44663);
and U44997 (N_44997,N_44607,N_44700);
or U44998 (N_44998,N_44676,N_44544);
or U44999 (N_44999,N_44678,N_44514);
or U45000 (N_45000,N_44808,N_44852);
nor U45001 (N_45001,N_44860,N_44883);
and U45002 (N_45002,N_44982,N_44838);
nor U45003 (N_45003,N_44907,N_44919);
nand U45004 (N_45004,N_44878,N_44990);
xor U45005 (N_45005,N_44758,N_44822);
nor U45006 (N_45006,N_44840,N_44966);
xor U45007 (N_45007,N_44825,N_44991);
xnor U45008 (N_45008,N_44987,N_44955);
nor U45009 (N_45009,N_44951,N_44917);
or U45010 (N_45010,N_44930,N_44816);
nor U45011 (N_45011,N_44913,N_44809);
nand U45012 (N_45012,N_44944,N_44847);
or U45013 (N_45013,N_44821,N_44996);
nor U45014 (N_45014,N_44999,N_44804);
or U45015 (N_45015,N_44993,N_44826);
xnor U45016 (N_45016,N_44882,N_44935);
and U45017 (N_45017,N_44752,N_44945);
and U45018 (N_45018,N_44842,N_44908);
or U45019 (N_45019,N_44768,N_44801);
nor U45020 (N_45020,N_44756,N_44875);
or U45021 (N_45021,N_44950,N_44839);
nand U45022 (N_45022,N_44880,N_44851);
or U45023 (N_45023,N_44976,N_44932);
or U45024 (N_45024,N_44832,N_44906);
xnor U45025 (N_45025,N_44977,N_44869);
nand U45026 (N_45026,N_44947,N_44909);
xnor U45027 (N_45027,N_44873,N_44904);
xnor U45028 (N_45028,N_44943,N_44787);
or U45029 (N_45029,N_44953,N_44823);
xor U45030 (N_45030,N_44819,N_44785);
nand U45031 (N_45031,N_44759,N_44974);
xor U45032 (N_45032,N_44762,N_44896);
nor U45033 (N_45033,N_44862,N_44789);
xnor U45034 (N_45034,N_44845,N_44771);
xor U45035 (N_45035,N_44778,N_44940);
or U45036 (N_45036,N_44864,N_44939);
nor U45037 (N_45037,N_44782,N_44961);
and U45038 (N_45038,N_44824,N_44918);
and U45039 (N_45039,N_44971,N_44854);
and U45040 (N_45040,N_44774,N_44897);
nand U45041 (N_45041,N_44853,N_44829);
and U45042 (N_45042,N_44973,N_44921);
or U45043 (N_45043,N_44901,N_44928);
xnor U45044 (N_45044,N_44751,N_44857);
nand U45045 (N_45045,N_44894,N_44879);
nor U45046 (N_45046,N_44992,N_44949);
and U45047 (N_45047,N_44886,N_44929);
and U45048 (N_45048,N_44763,N_44969);
and U45049 (N_45049,N_44946,N_44855);
nand U45050 (N_45050,N_44810,N_44916);
xor U45051 (N_45051,N_44858,N_44892);
nor U45052 (N_45052,N_44900,N_44877);
xnor U45053 (N_45053,N_44807,N_44849);
or U45054 (N_45054,N_44794,N_44898);
nor U45055 (N_45055,N_44958,N_44948);
nor U45056 (N_45056,N_44871,N_44750);
and U45057 (N_45057,N_44942,N_44910);
nand U45058 (N_45058,N_44815,N_44830);
and U45059 (N_45059,N_44802,N_44952);
and U45060 (N_45060,N_44786,N_44970);
xnor U45061 (N_45061,N_44818,N_44861);
and U45062 (N_45062,N_44905,N_44914);
or U45063 (N_45063,N_44784,N_44983);
xnor U45064 (N_45064,N_44941,N_44937);
nand U45065 (N_45065,N_44988,N_44841);
xnor U45066 (N_45066,N_44820,N_44781);
xor U45067 (N_45067,N_44817,N_44846);
xnor U45068 (N_45068,N_44985,N_44803);
and U45069 (N_45069,N_44856,N_44757);
and U45070 (N_45070,N_44795,N_44979);
nand U45071 (N_45071,N_44779,N_44933);
xnor U45072 (N_45072,N_44872,N_44911);
or U45073 (N_45073,N_44780,N_44798);
nor U45074 (N_45074,N_44960,N_44866);
and U45075 (N_45075,N_44967,N_44868);
nand U45076 (N_45076,N_44926,N_44931);
nor U45077 (N_45077,N_44790,N_44893);
xnor U45078 (N_45078,N_44850,N_44765);
or U45079 (N_45079,N_44938,N_44814);
and U45080 (N_45080,N_44890,N_44833);
nand U45081 (N_45081,N_44895,N_44859);
xnor U45082 (N_45082,N_44773,N_44902);
and U45083 (N_45083,N_44954,N_44792);
xnor U45084 (N_45084,N_44806,N_44793);
nand U45085 (N_45085,N_44865,N_44783);
or U45086 (N_45086,N_44831,N_44903);
xor U45087 (N_45087,N_44891,N_44796);
xor U45088 (N_45088,N_44776,N_44925);
nand U45089 (N_45089,N_44981,N_44964);
nand U45090 (N_45090,N_44837,N_44835);
or U45091 (N_45091,N_44767,N_44995);
and U45092 (N_45092,N_44811,N_44912);
nand U45093 (N_45093,N_44956,N_44848);
and U45094 (N_45094,N_44770,N_44936);
nand U45095 (N_45095,N_44797,N_44876);
nor U45096 (N_45096,N_44994,N_44959);
xor U45097 (N_45097,N_44965,N_44927);
nand U45098 (N_45098,N_44834,N_44915);
and U45099 (N_45099,N_44799,N_44836);
xor U45100 (N_45100,N_44764,N_44889);
xor U45101 (N_45101,N_44885,N_44828);
nor U45102 (N_45102,N_44957,N_44769);
nand U45103 (N_45103,N_44844,N_44874);
xor U45104 (N_45104,N_44899,N_44761);
xnor U45105 (N_45105,N_44755,N_44968);
nand U45106 (N_45106,N_44772,N_44997);
nor U45107 (N_45107,N_44887,N_44863);
nor U45108 (N_45108,N_44867,N_44975);
and U45109 (N_45109,N_44881,N_44980);
and U45110 (N_45110,N_44813,N_44800);
nor U45111 (N_45111,N_44998,N_44753);
and U45112 (N_45112,N_44888,N_44978);
and U45113 (N_45113,N_44924,N_44754);
nor U45114 (N_45114,N_44920,N_44963);
nand U45115 (N_45115,N_44870,N_44989);
nand U45116 (N_45116,N_44805,N_44775);
nand U45117 (N_45117,N_44934,N_44984);
and U45118 (N_45118,N_44986,N_44812);
xor U45119 (N_45119,N_44972,N_44923);
nand U45120 (N_45120,N_44788,N_44884);
and U45121 (N_45121,N_44760,N_44791);
or U45122 (N_45122,N_44843,N_44962);
xnor U45123 (N_45123,N_44766,N_44827);
xor U45124 (N_45124,N_44777,N_44922);
nor U45125 (N_45125,N_44881,N_44771);
or U45126 (N_45126,N_44791,N_44962);
nor U45127 (N_45127,N_44874,N_44752);
xor U45128 (N_45128,N_44809,N_44963);
and U45129 (N_45129,N_44857,N_44865);
nor U45130 (N_45130,N_44997,N_44863);
and U45131 (N_45131,N_44852,N_44768);
xnor U45132 (N_45132,N_44978,N_44906);
or U45133 (N_45133,N_44894,N_44900);
and U45134 (N_45134,N_44852,N_44837);
xor U45135 (N_45135,N_44825,N_44899);
nand U45136 (N_45136,N_44870,N_44968);
nor U45137 (N_45137,N_44858,N_44957);
and U45138 (N_45138,N_44857,N_44769);
xnor U45139 (N_45139,N_44933,N_44920);
or U45140 (N_45140,N_44768,N_44909);
xnor U45141 (N_45141,N_44785,N_44845);
nor U45142 (N_45142,N_44841,N_44874);
xor U45143 (N_45143,N_44964,N_44842);
xor U45144 (N_45144,N_44870,N_44820);
xor U45145 (N_45145,N_44883,N_44780);
and U45146 (N_45146,N_44806,N_44779);
nand U45147 (N_45147,N_44937,N_44826);
nor U45148 (N_45148,N_44952,N_44853);
and U45149 (N_45149,N_44921,N_44754);
nor U45150 (N_45150,N_44986,N_44963);
or U45151 (N_45151,N_44763,N_44965);
nor U45152 (N_45152,N_44894,N_44995);
xor U45153 (N_45153,N_44926,N_44859);
or U45154 (N_45154,N_44954,N_44904);
nor U45155 (N_45155,N_44910,N_44763);
or U45156 (N_45156,N_44913,N_44893);
and U45157 (N_45157,N_44768,N_44896);
xnor U45158 (N_45158,N_44755,N_44919);
nor U45159 (N_45159,N_44901,N_44798);
or U45160 (N_45160,N_44989,N_44764);
or U45161 (N_45161,N_44805,N_44940);
or U45162 (N_45162,N_44887,N_44814);
and U45163 (N_45163,N_44864,N_44905);
nand U45164 (N_45164,N_44802,N_44907);
xnor U45165 (N_45165,N_44844,N_44955);
xor U45166 (N_45166,N_44760,N_44775);
or U45167 (N_45167,N_44807,N_44817);
and U45168 (N_45168,N_44786,N_44962);
xor U45169 (N_45169,N_44820,N_44894);
nor U45170 (N_45170,N_44927,N_44999);
nand U45171 (N_45171,N_44782,N_44849);
and U45172 (N_45172,N_44956,N_44937);
nand U45173 (N_45173,N_44944,N_44783);
nand U45174 (N_45174,N_44841,N_44927);
xnor U45175 (N_45175,N_44814,N_44753);
xnor U45176 (N_45176,N_44826,N_44759);
nand U45177 (N_45177,N_44795,N_44912);
nor U45178 (N_45178,N_44971,N_44921);
nand U45179 (N_45179,N_44971,N_44966);
nand U45180 (N_45180,N_44962,N_44890);
nor U45181 (N_45181,N_44770,N_44803);
nor U45182 (N_45182,N_44787,N_44867);
nor U45183 (N_45183,N_44880,N_44763);
and U45184 (N_45184,N_44809,N_44985);
nor U45185 (N_45185,N_44950,N_44987);
nand U45186 (N_45186,N_44854,N_44887);
nor U45187 (N_45187,N_44795,N_44847);
xnor U45188 (N_45188,N_44788,N_44984);
nand U45189 (N_45189,N_44898,N_44757);
and U45190 (N_45190,N_44964,N_44786);
and U45191 (N_45191,N_44972,N_44947);
xor U45192 (N_45192,N_44911,N_44821);
and U45193 (N_45193,N_44948,N_44994);
and U45194 (N_45194,N_44840,N_44921);
nand U45195 (N_45195,N_44927,N_44922);
or U45196 (N_45196,N_44871,N_44889);
or U45197 (N_45197,N_44798,N_44763);
nand U45198 (N_45198,N_44879,N_44795);
nor U45199 (N_45199,N_44986,N_44989);
nand U45200 (N_45200,N_44838,N_44888);
xor U45201 (N_45201,N_44851,N_44762);
or U45202 (N_45202,N_44998,N_44800);
xor U45203 (N_45203,N_44846,N_44795);
and U45204 (N_45204,N_44867,N_44965);
nor U45205 (N_45205,N_44939,N_44918);
xnor U45206 (N_45206,N_44877,N_44979);
nand U45207 (N_45207,N_44803,N_44978);
or U45208 (N_45208,N_44843,N_44774);
xnor U45209 (N_45209,N_44993,N_44918);
xnor U45210 (N_45210,N_44956,N_44923);
and U45211 (N_45211,N_44987,N_44910);
nor U45212 (N_45212,N_44892,N_44819);
or U45213 (N_45213,N_44985,N_44901);
nand U45214 (N_45214,N_44818,N_44886);
and U45215 (N_45215,N_44883,N_44759);
and U45216 (N_45216,N_44944,N_44827);
nand U45217 (N_45217,N_44867,N_44805);
nor U45218 (N_45218,N_44881,N_44993);
nand U45219 (N_45219,N_44802,N_44951);
xnor U45220 (N_45220,N_44862,N_44823);
nand U45221 (N_45221,N_44941,N_44954);
xor U45222 (N_45222,N_44872,N_44776);
and U45223 (N_45223,N_44824,N_44921);
or U45224 (N_45224,N_44939,N_44961);
xor U45225 (N_45225,N_44900,N_44918);
xnor U45226 (N_45226,N_44832,N_44850);
or U45227 (N_45227,N_44804,N_44867);
nor U45228 (N_45228,N_44792,N_44797);
and U45229 (N_45229,N_44865,N_44918);
and U45230 (N_45230,N_44878,N_44814);
nand U45231 (N_45231,N_44922,N_44867);
xnor U45232 (N_45232,N_44802,N_44857);
xor U45233 (N_45233,N_44950,N_44799);
nand U45234 (N_45234,N_44852,N_44755);
or U45235 (N_45235,N_44940,N_44820);
nor U45236 (N_45236,N_44878,N_44779);
or U45237 (N_45237,N_44765,N_44763);
xnor U45238 (N_45238,N_44897,N_44931);
or U45239 (N_45239,N_44772,N_44979);
nand U45240 (N_45240,N_44883,N_44889);
nand U45241 (N_45241,N_44763,N_44791);
nand U45242 (N_45242,N_44882,N_44857);
or U45243 (N_45243,N_44843,N_44790);
and U45244 (N_45244,N_44936,N_44957);
or U45245 (N_45245,N_44885,N_44901);
nand U45246 (N_45246,N_44883,N_44827);
and U45247 (N_45247,N_44765,N_44937);
or U45248 (N_45248,N_44751,N_44891);
nand U45249 (N_45249,N_44866,N_44783);
nand U45250 (N_45250,N_45098,N_45111);
or U45251 (N_45251,N_45039,N_45007);
nand U45252 (N_45252,N_45165,N_45191);
nand U45253 (N_45253,N_45203,N_45090);
and U45254 (N_45254,N_45018,N_45229);
nor U45255 (N_45255,N_45127,N_45179);
or U45256 (N_45256,N_45215,N_45072);
and U45257 (N_45257,N_45190,N_45074);
nor U45258 (N_45258,N_45233,N_45133);
xor U45259 (N_45259,N_45146,N_45226);
nor U45260 (N_45260,N_45125,N_45021);
nand U45261 (N_45261,N_45145,N_45049);
or U45262 (N_45262,N_45202,N_45153);
or U45263 (N_45263,N_45106,N_45249);
and U45264 (N_45264,N_45036,N_45065);
nor U45265 (N_45265,N_45161,N_45167);
nand U45266 (N_45266,N_45015,N_45112);
xor U45267 (N_45267,N_45200,N_45010);
nor U45268 (N_45268,N_45030,N_45119);
or U45269 (N_45269,N_45023,N_45037);
nand U45270 (N_45270,N_45062,N_45210);
xor U45271 (N_45271,N_45033,N_45124);
nor U45272 (N_45272,N_45101,N_45014);
nand U45273 (N_45273,N_45143,N_45162);
nor U45274 (N_45274,N_45194,N_45219);
nor U45275 (N_45275,N_45198,N_45011);
nor U45276 (N_45276,N_45199,N_45218);
nor U45277 (N_45277,N_45099,N_45151);
or U45278 (N_45278,N_45044,N_45178);
nor U45279 (N_45279,N_45135,N_45168);
nor U45280 (N_45280,N_45078,N_45000);
and U45281 (N_45281,N_45116,N_45117);
nor U45282 (N_45282,N_45164,N_45017);
nand U45283 (N_45283,N_45042,N_45245);
and U45284 (N_45284,N_45114,N_45103);
nand U45285 (N_45285,N_45080,N_45139);
nand U45286 (N_45286,N_45189,N_45123);
xnor U45287 (N_45287,N_45100,N_45142);
nand U45288 (N_45288,N_45003,N_45175);
and U45289 (N_45289,N_45009,N_45087);
or U45290 (N_45290,N_45109,N_45154);
nor U45291 (N_45291,N_45110,N_45188);
nand U45292 (N_45292,N_45056,N_45217);
nor U45293 (N_45293,N_45152,N_45070);
and U45294 (N_45294,N_45132,N_45025);
nor U45295 (N_45295,N_45184,N_45107);
and U45296 (N_45296,N_45158,N_45144);
nand U45297 (N_45297,N_45169,N_45211);
or U45298 (N_45298,N_45005,N_45108);
and U45299 (N_45299,N_45081,N_45063);
and U45300 (N_45300,N_45008,N_45197);
xnor U45301 (N_45301,N_45013,N_45136);
nor U45302 (N_45302,N_45032,N_45075);
or U45303 (N_45303,N_45035,N_45246);
nand U45304 (N_45304,N_45243,N_45248);
nor U45305 (N_45305,N_45223,N_45242);
or U45306 (N_45306,N_45174,N_45232);
or U45307 (N_45307,N_45069,N_45201);
nand U45308 (N_45308,N_45216,N_45076);
xnor U45309 (N_45309,N_45064,N_45137);
xnor U45310 (N_45310,N_45182,N_45066);
nand U45311 (N_45311,N_45237,N_45170);
nand U45312 (N_45312,N_45068,N_45057);
and U45313 (N_45313,N_45016,N_45053);
nand U45314 (N_45314,N_45160,N_45140);
and U45315 (N_45315,N_45047,N_45061);
nor U45316 (N_45316,N_45083,N_45067);
and U45317 (N_45317,N_45102,N_45084);
and U45318 (N_45318,N_45048,N_45038);
and U45319 (N_45319,N_45028,N_45089);
nand U45320 (N_45320,N_45180,N_45227);
nor U45321 (N_45321,N_45094,N_45024);
nand U45322 (N_45322,N_45236,N_45026);
nand U45323 (N_45323,N_45001,N_45212);
and U45324 (N_45324,N_45234,N_45045);
or U45325 (N_45325,N_45171,N_45131);
nor U45326 (N_45326,N_45091,N_45181);
and U45327 (N_45327,N_45221,N_45029);
and U45328 (N_45328,N_45156,N_45041);
nor U45329 (N_45329,N_45134,N_45240);
xor U45330 (N_45330,N_45079,N_45238);
and U45331 (N_45331,N_45173,N_45247);
nor U45332 (N_45332,N_45088,N_45196);
and U45333 (N_45333,N_45052,N_45126);
nor U45334 (N_45334,N_45043,N_45166);
nor U45335 (N_45335,N_45115,N_45129);
nor U45336 (N_45336,N_45128,N_45224);
nor U45337 (N_45337,N_45239,N_45022);
and U45338 (N_45338,N_45244,N_45130);
nand U45339 (N_45339,N_45207,N_45209);
xor U45340 (N_45340,N_45138,N_45230);
xnor U45341 (N_45341,N_45159,N_45002);
nand U45342 (N_45342,N_45222,N_45085);
xnor U45343 (N_45343,N_45104,N_45141);
xnor U45344 (N_45344,N_45241,N_45147);
xor U45345 (N_45345,N_45185,N_45172);
and U45346 (N_45346,N_45118,N_45235);
or U45347 (N_45347,N_45095,N_45177);
xnor U45348 (N_45348,N_45205,N_45097);
and U45349 (N_45349,N_45213,N_45073);
nand U45350 (N_45350,N_45077,N_45071);
nand U45351 (N_45351,N_45148,N_45020);
nand U45352 (N_45352,N_45086,N_45155);
and U45353 (N_45353,N_45113,N_45157);
xnor U45354 (N_45354,N_45006,N_45208);
xnor U45355 (N_45355,N_45206,N_45040);
xor U45356 (N_45356,N_45004,N_45060);
nand U45357 (N_45357,N_45187,N_45150);
xor U45358 (N_45358,N_45120,N_45050);
xor U45359 (N_45359,N_45193,N_45058);
and U45360 (N_45360,N_45122,N_45046);
xor U45361 (N_45361,N_45228,N_45163);
nor U45362 (N_45362,N_45220,N_45092);
and U45363 (N_45363,N_45192,N_45082);
nor U45364 (N_45364,N_45176,N_45186);
nand U45365 (N_45365,N_45195,N_45096);
xor U45366 (N_45366,N_45204,N_45019);
and U45367 (N_45367,N_45121,N_45183);
and U45368 (N_45368,N_45059,N_45105);
and U45369 (N_45369,N_45225,N_45055);
nor U45370 (N_45370,N_45034,N_45093);
and U45371 (N_45371,N_45149,N_45214);
nand U45372 (N_45372,N_45231,N_45031);
nand U45373 (N_45373,N_45051,N_45027);
and U45374 (N_45374,N_45054,N_45012);
or U45375 (N_45375,N_45209,N_45186);
or U45376 (N_45376,N_45115,N_45074);
nor U45377 (N_45377,N_45156,N_45220);
nand U45378 (N_45378,N_45048,N_45020);
or U45379 (N_45379,N_45133,N_45043);
and U45380 (N_45380,N_45002,N_45160);
nor U45381 (N_45381,N_45195,N_45158);
or U45382 (N_45382,N_45065,N_45239);
or U45383 (N_45383,N_45144,N_45093);
and U45384 (N_45384,N_45178,N_45113);
nor U45385 (N_45385,N_45074,N_45123);
nor U45386 (N_45386,N_45078,N_45059);
nor U45387 (N_45387,N_45071,N_45037);
or U45388 (N_45388,N_45058,N_45209);
and U45389 (N_45389,N_45115,N_45140);
nand U45390 (N_45390,N_45110,N_45239);
xnor U45391 (N_45391,N_45086,N_45123);
or U45392 (N_45392,N_45045,N_45078);
nor U45393 (N_45393,N_45022,N_45071);
xor U45394 (N_45394,N_45236,N_45040);
or U45395 (N_45395,N_45189,N_45068);
xnor U45396 (N_45396,N_45145,N_45150);
nand U45397 (N_45397,N_45039,N_45030);
or U45398 (N_45398,N_45188,N_45186);
and U45399 (N_45399,N_45039,N_45052);
or U45400 (N_45400,N_45041,N_45031);
nor U45401 (N_45401,N_45033,N_45056);
nor U45402 (N_45402,N_45133,N_45234);
and U45403 (N_45403,N_45109,N_45086);
nand U45404 (N_45404,N_45145,N_45126);
or U45405 (N_45405,N_45048,N_45004);
or U45406 (N_45406,N_45168,N_45021);
nand U45407 (N_45407,N_45239,N_45249);
or U45408 (N_45408,N_45111,N_45197);
nor U45409 (N_45409,N_45225,N_45137);
or U45410 (N_45410,N_45094,N_45150);
and U45411 (N_45411,N_45014,N_45086);
nor U45412 (N_45412,N_45189,N_45210);
xor U45413 (N_45413,N_45001,N_45151);
nand U45414 (N_45414,N_45049,N_45141);
xor U45415 (N_45415,N_45128,N_45238);
nand U45416 (N_45416,N_45035,N_45127);
nand U45417 (N_45417,N_45199,N_45156);
and U45418 (N_45418,N_45060,N_45188);
xor U45419 (N_45419,N_45000,N_45054);
or U45420 (N_45420,N_45029,N_45018);
nor U45421 (N_45421,N_45044,N_45015);
nor U45422 (N_45422,N_45077,N_45120);
nand U45423 (N_45423,N_45229,N_45035);
and U45424 (N_45424,N_45133,N_45247);
or U45425 (N_45425,N_45075,N_45232);
or U45426 (N_45426,N_45218,N_45147);
nor U45427 (N_45427,N_45047,N_45003);
nor U45428 (N_45428,N_45084,N_45071);
nor U45429 (N_45429,N_45161,N_45235);
nand U45430 (N_45430,N_45010,N_45092);
and U45431 (N_45431,N_45204,N_45178);
nand U45432 (N_45432,N_45156,N_45113);
or U45433 (N_45433,N_45243,N_45089);
nor U45434 (N_45434,N_45037,N_45113);
nor U45435 (N_45435,N_45193,N_45075);
nand U45436 (N_45436,N_45018,N_45158);
and U45437 (N_45437,N_45017,N_45183);
or U45438 (N_45438,N_45202,N_45026);
and U45439 (N_45439,N_45101,N_45209);
nor U45440 (N_45440,N_45064,N_45216);
nor U45441 (N_45441,N_45181,N_45174);
xor U45442 (N_45442,N_45028,N_45040);
and U45443 (N_45443,N_45190,N_45122);
nor U45444 (N_45444,N_45130,N_45008);
or U45445 (N_45445,N_45236,N_45041);
and U45446 (N_45446,N_45080,N_45092);
or U45447 (N_45447,N_45047,N_45046);
and U45448 (N_45448,N_45005,N_45020);
nor U45449 (N_45449,N_45039,N_45100);
nand U45450 (N_45450,N_45024,N_45206);
xnor U45451 (N_45451,N_45181,N_45210);
nor U45452 (N_45452,N_45046,N_45147);
or U45453 (N_45453,N_45038,N_45000);
xor U45454 (N_45454,N_45077,N_45033);
and U45455 (N_45455,N_45078,N_45052);
nand U45456 (N_45456,N_45195,N_45088);
xnor U45457 (N_45457,N_45137,N_45228);
xnor U45458 (N_45458,N_45095,N_45243);
xnor U45459 (N_45459,N_45101,N_45241);
and U45460 (N_45460,N_45185,N_45039);
or U45461 (N_45461,N_45106,N_45064);
xor U45462 (N_45462,N_45030,N_45111);
and U45463 (N_45463,N_45010,N_45085);
or U45464 (N_45464,N_45157,N_45159);
or U45465 (N_45465,N_45173,N_45207);
nor U45466 (N_45466,N_45000,N_45216);
nor U45467 (N_45467,N_45048,N_45212);
xnor U45468 (N_45468,N_45149,N_45078);
or U45469 (N_45469,N_45235,N_45099);
nor U45470 (N_45470,N_45074,N_45185);
xnor U45471 (N_45471,N_45021,N_45100);
xnor U45472 (N_45472,N_45078,N_45230);
or U45473 (N_45473,N_45174,N_45017);
nand U45474 (N_45474,N_45110,N_45218);
and U45475 (N_45475,N_45192,N_45128);
and U45476 (N_45476,N_45123,N_45242);
xnor U45477 (N_45477,N_45245,N_45237);
or U45478 (N_45478,N_45013,N_45228);
xnor U45479 (N_45479,N_45237,N_45249);
nand U45480 (N_45480,N_45111,N_45168);
xnor U45481 (N_45481,N_45122,N_45221);
xnor U45482 (N_45482,N_45234,N_45155);
nor U45483 (N_45483,N_45070,N_45048);
xor U45484 (N_45484,N_45141,N_45144);
xnor U45485 (N_45485,N_45008,N_45096);
xnor U45486 (N_45486,N_45125,N_45030);
nor U45487 (N_45487,N_45051,N_45129);
nand U45488 (N_45488,N_45198,N_45190);
or U45489 (N_45489,N_45140,N_45187);
and U45490 (N_45490,N_45115,N_45235);
and U45491 (N_45491,N_45021,N_45051);
nand U45492 (N_45492,N_45103,N_45047);
or U45493 (N_45493,N_45236,N_45192);
and U45494 (N_45494,N_45220,N_45155);
xnor U45495 (N_45495,N_45059,N_45227);
nand U45496 (N_45496,N_45177,N_45022);
nand U45497 (N_45497,N_45120,N_45142);
or U45498 (N_45498,N_45052,N_45017);
nor U45499 (N_45499,N_45108,N_45043);
nand U45500 (N_45500,N_45449,N_45346);
xnor U45501 (N_45501,N_45323,N_45385);
nand U45502 (N_45502,N_45444,N_45276);
nand U45503 (N_45503,N_45339,N_45314);
xnor U45504 (N_45504,N_45312,N_45362);
nand U45505 (N_45505,N_45496,N_45391);
or U45506 (N_45506,N_45471,N_45465);
and U45507 (N_45507,N_45288,N_45354);
xor U45508 (N_45508,N_45369,N_45324);
xnor U45509 (N_45509,N_45364,N_45454);
nand U45510 (N_45510,N_45292,N_45371);
nor U45511 (N_45511,N_45280,N_45299);
xor U45512 (N_45512,N_45421,N_45394);
nor U45513 (N_45513,N_45309,N_45481);
nor U45514 (N_45514,N_45416,N_45350);
and U45515 (N_45515,N_45376,N_45396);
and U45516 (N_45516,N_45414,N_45410);
xor U45517 (N_45517,N_45261,N_45306);
nor U45518 (N_45518,N_45353,N_45476);
xor U45519 (N_45519,N_45315,N_45466);
nand U45520 (N_45520,N_45310,N_45426);
xor U45521 (N_45521,N_45372,N_45401);
nor U45522 (N_45522,N_45268,N_45266);
xnor U45523 (N_45523,N_45408,N_45267);
and U45524 (N_45524,N_45365,N_45457);
or U45525 (N_45525,N_45291,N_45419);
or U45526 (N_45526,N_45434,N_45258);
xor U45527 (N_45527,N_45286,N_45327);
nand U45528 (N_45528,N_45432,N_45497);
and U45529 (N_45529,N_45265,N_45326);
xnor U45530 (N_45530,N_45355,N_45322);
xnor U45531 (N_45531,N_45460,N_45431);
and U45532 (N_45532,N_45274,N_45285);
and U45533 (N_45533,N_45341,N_45435);
nor U45534 (N_45534,N_45433,N_45424);
nor U45535 (N_45535,N_45332,N_45422);
xor U45536 (N_45536,N_45379,N_45380);
or U45537 (N_45537,N_45320,N_45482);
and U45538 (N_45538,N_45490,N_45305);
xnor U45539 (N_45539,N_45361,N_45281);
nand U45540 (N_45540,N_45381,N_45415);
xor U45541 (N_45541,N_45319,N_45253);
nand U45542 (N_45542,N_45384,N_45483);
xnor U45543 (N_45543,N_45260,N_45284);
nand U45544 (N_45544,N_45297,N_45360);
or U45545 (N_45545,N_45373,N_45272);
xnor U45546 (N_45546,N_45256,N_45455);
xor U45547 (N_45547,N_45448,N_45287);
or U45548 (N_45548,N_45321,N_45464);
xnor U45549 (N_45549,N_45366,N_45349);
nor U45550 (N_45550,N_45450,N_45472);
or U45551 (N_45551,N_45270,N_45377);
and U45552 (N_45552,N_45337,N_45283);
nor U45553 (N_45553,N_45345,N_45289);
nor U45554 (N_45554,N_45404,N_45313);
nor U45555 (N_45555,N_45370,N_45342);
xnor U45556 (N_45556,N_45441,N_45395);
nor U45557 (N_45557,N_45255,N_45367);
xnor U45558 (N_45558,N_45328,N_45397);
xnor U45559 (N_45559,N_45439,N_45375);
nand U45560 (N_45560,N_45279,N_45290);
xor U45561 (N_45561,N_45257,N_45277);
xor U45562 (N_45562,N_45462,N_45458);
xor U45563 (N_45563,N_45393,N_45269);
xor U45564 (N_45564,N_45440,N_45495);
and U45565 (N_45565,N_45417,N_45390);
xor U45566 (N_45566,N_45488,N_45344);
or U45567 (N_45567,N_45438,N_45402);
and U45568 (N_45568,N_45333,N_45445);
or U45569 (N_45569,N_45386,N_45493);
nor U45570 (N_45570,N_45485,N_45318);
or U45571 (N_45571,N_45251,N_45461);
or U45572 (N_45572,N_45356,N_45301);
nor U45573 (N_45573,N_45335,N_45378);
xor U45574 (N_45574,N_45275,N_45363);
nor U45575 (N_45575,N_45352,N_45316);
and U45576 (N_45576,N_45409,N_45311);
nand U45577 (N_45577,N_45451,N_45442);
xnor U45578 (N_45578,N_45329,N_45368);
nor U45579 (N_45579,N_45358,N_45492);
xor U45580 (N_45580,N_45308,N_45413);
nand U45581 (N_45581,N_45259,N_45498);
nor U45582 (N_45582,N_45262,N_45427);
xnor U45583 (N_45583,N_45452,N_45307);
nor U45584 (N_45584,N_45294,N_45343);
xnor U45585 (N_45585,N_45263,N_45347);
nor U45586 (N_45586,N_45499,N_45486);
nand U45587 (N_45587,N_45374,N_45487);
or U45588 (N_45588,N_45475,N_45389);
or U45589 (N_45589,N_45340,N_45304);
nand U45590 (N_45590,N_45298,N_45250);
xor U45591 (N_45591,N_45477,N_45484);
nor U45592 (N_45592,N_45479,N_45491);
or U45593 (N_45593,N_45405,N_45403);
and U45594 (N_45594,N_45383,N_45467);
xnor U45595 (N_45595,N_45423,N_45334);
and U45596 (N_45596,N_45398,N_45446);
or U45597 (N_45597,N_45428,N_45348);
and U45598 (N_45598,N_45480,N_45425);
or U45599 (N_45599,N_45437,N_45325);
nand U45600 (N_45600,N_45468,N_45387);
and U45601 (N_45601,N_45336,N_45436);
xor U45602 (N_45602,N_45469,N_45478);
nand U45603 (N_45603,N_45411,N_45494);
nor U45604 (N_45604,N_45302,N_45392);
and U45605 (N_45605,N_45382,N_45473);
nand U45606 (N_45606,N_45303,N_45443);
xnor U45607 (N_45607,N_45282,N_45273);
or U45608 (N_45608,N_45463,N_45459);
or U45609 (N_45609,N_45447,N_45338);
nand U45610 (N_45610,N_45399,N_45296);
nand U45611 (N_45611,N_45293,N_45317);
nand U45612 (N_45612,N_45295,N_45418);
or U45613 (N_45613,N_45351,N_45254);
nor U45614 (N_45614,N_45412,N_45489);
nand U45615 (N_45615,N_45300,N_45357);
nand U45616 (N_45616,N_45264,N_45456);
and U45617 (N_45617,N_45407,N_45330);
and U45618 (N_45618,N_45406,N_45400);
nand U45619 (N_45619,N_45474,N_45252);
nand U45620 (N_45620,N_45453,N_45359);
and U45621 (N_45621,N_45388,N_45429);
nor U45622 (N_45622,N_45278,N_45430);
xor U45623 (N_45623,N_45331,N_45271);
xor U45624 (N_45624,N_45470,N_45420);
and U45625 (N_45625,N_45458,N_45252);
and U45626 (N_45626,N_45414,N_45297);
and U45627 (N_45627,N_45361,N_45260);
or U45628 (N_45628,N_45467,N_45415);
nand U45629 (N_45629,N_45357,N_45407);
nand U45630 (N_45630,N_45409,N_45459);
or U45631 (N_45631,N_45273,N_45355);
nor U45632 (N_45632,N_45326,N_45282);
and U45633 (N_45633,N_45384,N_45490);
nor U45634 (N_45634,N_45270,N_45362);
xnor U45635 (N_45635,N_45320,N_45311);
xor U45636 (N_45636,N_45289,N_45262);
nand U45637 (N_45637,N_45488,N_45454);
nor U45638 (N_45638,N_45390,N_45495);
xor U45639 (N_45639,N_45352,N_45262);
nand U45640 (N_45640,N_45346,N_45493);
nand U45641 (N_45641,N_45461,N_45479);
xor U45642 (N_45642,N_45329,N_45312);
and U45643 (N_45643,N_45406,N_45277);
nand U45644 (N_45644,N_45499,N_45335);
nor U45645 (N_45645,N_45427,N_45305);
xnor U45646 (N_45646,N_45387,N_45330);
or U45647 (N_45647,N_45473,N_45387);
and U45648 (N_45648,N_45469,N_45256);
or U45649 (N_45649,N_45458,N_45392);
and U45650 (N_45650,N_45283,N_45488);
and U45651 (N_45651,N_45377,N_45341);
and U45652 (N_45652,N_45477,N_45464);
nor U45653 (N_45653,N_45469,N_45255);
nor U45654 (N_45654,N_45290,N_45427);
or U45655 (N_45655,N_45499,N_45295);
xnor U45656 (N_45656,N_45256,N_45275);
or U45657 (N_45657,N_45353,N_45439);
or U45658 (N_45658,N_45476,N_45429);
and U45659 (N_45659,N_45464,N_45263);
and U45660 (N_45660,N_45358,N_45283);
nand U45661 (N_45661,N_45259,N_45253);
nor U45662 (N_45662,N_45302,N_45391);
nand U45663 (N_45663,N_45363,N_45309);
and U45664 (N_45664,N_45473,N_45266);
nor U45665 (N_45665,N_45341,N_45418);
nand U45666 (N_45666,N_45427,N_45283);
nand U45667 (N_45667,N_45408,N_45353);
and U45668 (N_45668,N_45364,N_45433);
or U45669 (N_45669,N_45456,N_45472);
xnor U45670 (N_45670,N_45286,N_45328);
xor U45671 (N_45671,N_45318,N_45323);
nor U45672 (N_45672,N_45335,N_45444);
xnor U45673 (N_45673,N_45459,N_45320);
nand U45674 (N_45674,N_45407,N_45476);
or U45675 (N_45675,N_45415,N_45423);
and U45676 (N_45676,N_45466,N_45406);
xnor U45677 (N_45677,N_45412,N_45335);
and U45678 (N_45678,N_45367,N_45312);
xor U45679 (N_45679,N_45414,N_45266);
and U45680 (N_45680,N_45315,N_45488);
xor U45681 (N_45681,N_45493,N_45410);
or U45682 (N_45682,N_45286,N_45364);
and U45683 (N_45683,N_45492,N_45356);
or U45684 (N_45684,N_45359,N_45299);
and U45685 (N_45685,N_45267,N_45411);
nor U45686 (N_45686,N_45338,N_45463);
nand U45687 (N_45687,N_45263,N_45362);
xor U45688 (N_45688,N_45388,N_45495);
xnor U45689 (N_45689,N_45292,N_45490);
nand U45690 (N_45690,N_45389,N_45303);
or U45691 (N_45691,N_45471,N_45479);
nand U45692 (N_45692,N_45498,N_45287);
nor U45693 (N_45693,N_45319,N_45402);
and U45694 (N_45694,N_45464,N_45453);
nand U45695 (N_45695,N_45461,N_45434);
nor U45696 (N_45696,N_45315,N_45260);
nor U45697 (N_45697,N_45279,N_45392);
nor U45698 (N_45698,N_45380,N_45374);
nand U45699 (N_45699,N_45497,N_45408);
and U45700 (N_45700,N_45417,N_45372);
xor U45701 (N_45701,N_45324,N_45306);
nor U45702 (N_45702,N_45341,N_45452);
nor U45703 (N_45703,N_45422,N_45499);
or U45704 (N_45704,N_45422,N_45338);
nor U45705 (N_45705,N_45429,N_45410);
nor U45706 (N_45706,N_45388,N_45254);
nand U45707 (N_45707,N_45264,N_45357);
and U45708 (N_45708,N_45481,N_45303);
xnor U45709 (N_45709,N_45299,N_45448);
or U45710 (N_45710,N_45401,N_45260);
nand U45711 (N_45711,N_45339,N_45288);
nand U45712 (N_45712,N_45431,N_45492);
or U45713 (N_45713,N_45461,N_45266);
xnor U45714 (N_45714,N_45250,N_45438);
nor U45715 (N_45715,N_45477,N_45362);
and U45716 (N_45716,N_45467,N_45345);
nor U45717 (N_45717,N_45387,N_45435);
xor U45718 (N_45718,N_45421,N_45291);
xnor U45719 (N_45719,N_45266,N_45310);
nor U45720 (N_45720,N_45388,N_45305);
nor U45721 (N_45721,N_45392,N_45451);
xor U45722 (N_45722,N_45270,N_45363);
nand U45723 (N_45723,N_45450,N_45413);
xor U45724 (N_45724,N_45330,N_45480);
and U45725 (N_45725,N_45345,N_45259);
xor U45726 (N_45726,N_45277,N_45297);
nand U45727 (N_45727,N_45370,N_45315);
nor U45728 (N_45728,N_45441,N_45416);
nor U45729 (N_45729,N_45466,N_45357);
and U45730 (N_45730,N_45348,N_45331);
or U45731 (N_45731,N_45486,N_45415);
xor U45732 (N_45732,N_45272,N_45440);
xnor U45733 (N_45733,N_45492,N_45284);
nand U45734 (N_45734,N_45443,N_45461);
or U45735 (N_45735,N_45336,N_45255);
and U45736 (N_45736,N_45450,N_45359);
xnor U45737 (N_45737,N_45497,N_45315);
and U45738 (N_45738,N_45464,N_45430);
or U45739 (N_45739,N_45350,N_45382);
or U45740 (N_45740,N_45252,N_45389);
nor U45741 (N_45741,N_45286,N_45387);
or U45742 (N_45742,N_45493,N_45277);
nand U45743 (N_45743,N_45479,N_45336);
and U45744 (N_45744,N_45332,N_45451);
nor U45745 (N_45745,N_45448,N_45293);
or U45746 (N_45746,N_45400,N_45430);
and U45747 (N_45747,N_45399,N_45370);
or U45748 (N_45748,N_45377,N_45397);
nand U45749 (N_45749,N_45475,N_45368);
nor U45750 (N_45750,N_45712,N_45627);
nand U45751 (N_45751,N_45704,N_45662);
nand U45752 (N_45752,N_45713,N_45723);
nor U45753 (N_45753,N_45587,N_45707);
or U45754 (N_45754,N_45520,N_45694);
nor U45755 (N_45755,N_45552,N_45680);
and U45756 (N_45756,N_45700,N_45626);
and U45757 (N_45757,N_45669,N_45628);
nor U45758 (N_45758,N_45687,N_45548);
nand U45759 (N_45759,N_45543,N_45584);
or U45760 (N_45760,N_45651,N_45732);
and U45761 (N_45761,N_45741,N_45632);
xnor U45762 (N_45762,N_45560,N_45597);
and U45763 (N_45763,N_45648,N_45519);
nor U45764 (N_45764,N_45736,N_45657);
nand U45765 (N_45765,N_45720,N_45544);
and U45766 (N_45766,N_45722,N_45529);
nor U45767 (N_45767,N_45624,N_45563);
nor U45768 (N_45768,N_45703,N_45592);
or U45769 (N_45769,N_45638,N_45616);
nor U45770 (N_45770,N_45571,N_45532);
and U45771 (N_45771,N_45649,N_45598);
or U45772 (N_45772,N_45709,N_45664);
and U45773 (N_45773,N_45689,N_45677);
and U45774 (N_45774,N_45555,N_45611);
nand U45775 (N_45775,N_45710,N_45581);
nor U45776 (N_45776,N_45576,N_45533);
nand U45777 (N_45777,N_45727,N_45537);
and U45778 (N_45778,N_45526,N_45614);
or U45779 (N_45779,N_45575,N_45623);
nand U45780 (N_45780,N_45594,N_45735);
xnor U45781 (N_45781,N_45605,N_45553);
and U45782 (N_45782,N_45595,N_45679);
or U45783 (N_45783,N_45517,N_45582);
xor U45784 (N_45784,N_45522,N_45535);
and U45785 (N_45785,N_45633,N_45599);
xnor U45786 (N_45786,N_45591,N_45647);
nor U45787 (N_45787,N_45618,N_45536);
and U45788 (N_45788,N_45566,N_45600);
and U45789 (N_45789,N_45534,N_45644);
or U45790 (N_45790,N_45564,N_45739);
or U45791 (N_45791,N_45593,N_45745);
or U45792 (N_45792,N_45615,N_45637);
xor U45793 (N_45793,N_45681,N_45556);
and U45794 (N_45794,N_45507,N_45684);
nor U45795 (N_45795,N_45572,N_45646);
and U45796 (N_45796,N_45653,N_45683);
and U45797 (N_45797,N_45728,N_45740);
or U45798 (N_45798,N_45510,N_45641);
nor U45799 (N_45799,N_45719,N_45516);
nor U45800 (N_45800,N_45559,N_45521);
xnor U45801 (N_45801,N_45539,N_45691);
xnor U45802 (N_45802,N_45718,N_45506);
nor U45803 (N_45803,N_45749,N_45569);
nand U45804 (N_45804,N_45642,N_45668);
nor U45805 (N_45805,N_45607,N_45578);
nand U45806 (N_45806,N_45549,N_45730);
and U45807 (N_45807,N_45655,N_45562);
or U45808 (N_45808,N_45588,N_45692);
nor U45809 (N_45809,N_45630,N_45667);
nand U45810 (N_45810,N_45746,N_45635);
nand U45811 (N_45811,N_45579,N_45685);
xnor U45812 (N_45812,N_45501,N_45620);
nand U45813 (N_45813,N_45554,N_45702);
or U45814 (N_45814,N_45613,N_45701);
or U45815 (N_45815,N_45511,N_45663);
or U45816 (N_45816,N_45608,N_45733);
xor U45817 (N_45817,N_45688,N_45546);
or U45818 (N_45818,N_45551,N_45666);
xnor U45819 (N_45819,N_45557,N_45545);
nand U45820 (N_45820,N_45738,N_45531);
or U45821 (N_45821,N_45512,N_45699);
nor U45822 (N_45822,N_45527,N_45636);
and U45823 (N_45823,N_45603,N_45696);
nor U45824 (N_45824,N_45604,N_45590);
or U45825 (N_45825,N_45612,N_45742);
nor U45826 (N_45826,N_45565,N_45602);
xnor U45827 (N_45827,N_45672,N_45671);
or U45828 (N_45828,N_45660,N_45729);
or U45829 (N_45829,N_45747,N_45693);
nor U45830 (N_45830,N_45528,N_45670);
and U45831 (N_45831,N_45540,N_45695);
xnor U45832 (N_45832,N_45731,N_45715);
xor U45833 (N_45833,N_45558,N_45639);
or U45834 (N_45834,N_45568,N_45634);
xnor U45835 (N_45835,N_45580,N_45659);
nor U45836 (N_45836,N_45711,N_45690);
nor U45837 (N_45837,N_45518,N_45622);
and U45838 (N_45838,N_45547,N_45734);
or U45839 (N_45839,N_45744,N_45708);
or U45840 (N_45840,N_45714,N_45585);
nand U45841 (N_45841,N_45619,N_45724);
nand U45842 (N_45842,N_45538,N_45686);
nor U45843 (N_45843,N_45721,N_45661);
nor U45844 (N_45844,N_45525,N_45503);
nand U45845 (N_45845,N_45643,N_45596);
xor U45846 (N_45846,N_45541,N_45513);
nand U45847 (N_45847,N_45698,N_45743);
nand U45848 (N_45848,N_45629,N_45645);
nand U45849 (N_45849,N_45561,N_45678);
nand U45850 (N_45850,N_45676,N_45654);
and U45851 (N_45851,N_45682,N_45586);
xor U45852 (N_45852,N_45567,N_45748);
or U45853 (N_45853,N_45675,N_45514);
nand U45854 (N_45854,N_45658,N_45500);
xor U45855 (N_45855,N_45573,N_45502);
nand U45856 (N_45856,N_45674,N_45515);
nand U45857 (N_45857,N_45665,N_45673);
and U45858 (N_45858,N_45574,N_45589);
xor U45859 (N_45859,N_45705,N_45650);
nand U45860 (N_45860,N_45524,N_45716);
xnor U45861 (N_45861,N_45652,N_45523);
nor U45862 (N_45862,N_45509,N_45656);
nor U45863 (N_45863,N_45601,N_45583);
nor U45864 (N_45864,N_45570,N_45530);
and U45865 (N_45865,N_45617,N_45606);
xnor U45866 (N_45866,N_45717,N_45625);
xnor U45867 (N_45867,N_45725,N_45610);
nand U45868 (N_45868,N_45505,N_45706);
xnor U45869 (N_45869,N_45640,N_45577);
and U45870 (N_45870,N_45726,N_45550);
nand U45871 (N_45871,N_45504,N_45621);
or U45872 (N_45872,N_45737,N_45609);
nand U45873 (N_45873,N_45508,N_45542);
nor U45874 (N_45874,N_45697,N_45631);
nand U45875 (N_45875,N_45710,N_45744);
or U45876 (N_45876,N_45713,N_45566);
or U45877 (N_45877,N_45577,N_45516);
nand U45878 (N_45878,N_45656,N_45712);
or U45879 (N_45879,N_45503,N_45563);
xor U45880 (N_45880,N_45500,N_45647);
nand U45881 (N_45881,N_45611,N_45613);
or U45882 (N_45882,N_45519,N_45514);
nor U45883 (N_45883,N_45508,N_45607);
and U45884 (N_45884,N_45583,N_45519);
and U45885 (N_45885,N_45517,N_45588);
xor U45886 (N_45886,N_45622,N_45567);
nand U45887 (N_45887,N_45682,N_45541);
nor U45888 (N_45888,N_45616,N_45651);
or U45889 (N_45889,N_45590,N_45672);
xor U45890 (N_45890,N_45507,N_45673);
and U45891 (N_45891,N_45747,N_45675);
nand U45892 (N_45892,N_45514,N_45600);
nor U45893 (N_45893,N_45525,N_45615);
xor U45894 (N_45894,N_45682,N_45724);
or U45895 (N_45895,N_45729,N_45516);
xor U45896 (N_45896,N_45591,N_45700);
nand U45897 (N_45897,N_45550,N_45631);
nand U45898 (N_45898,N_45563,N_45682);
xor U45899 (N_45899,N_45564,N_45717);
nor U45900 (N_45900,N_45686,N_45625);
xor U45901 (N_45901,N_45736,N_45520);
nand U45902 (N_45902,N_45554,N_45669);
xor U45903 (N_45903,N_45538,N_45598);
or U45904 (N_45904,N_45618,N_45694);
and U45905 (N_45905,N_45519,N_45728);
nor U45906 (N_45906,N_45547,N_45722);
and U45907 (N_45907,N_45673,N_45580);
nand U45908 (N_45908,N_45740,N_45685);
nor U45909 (N_45909,N_45516,N_45661);
xor U45910 (N_45910,N_45558,N_45506);
xor U45911 (N_45911,N_45722,N_45708);
xor U45912 (N_45912,N_45643,N_45661);
xor U45913 (N_45913,N_45512,N_45645);
nand U45914 (N_45914,N_45724,N_45725);
nor U45915 (N_45915,N_45687,N_45657);
nand U45916 (N_45916,N_45535,N_45577);
nand U45917 (N_45917,N_45652,N_45611);
and U45918 (N_45918,N_45552,N_45723);
or U45919 (N_45919,N_45534,N_45611);
xnor U45920 (N_45920,N_45736,N_45522);
xor U45921 (N_45921,N_45565,N_45519);
xnor U45922 (N_45922,N_45641,N_45746);
nor U45923 (N_45923,N_45618,N_45520);
xor U45924 (N_45924,N_45613,N_45521);
and U45925 (N_45925,N_45702,N_45551);
nor U45926 (N_45926,N_45697,N_45705);
xor U45927 (N_45927,N_45630,N_45504);
and U45928 (N_45928,N_45633,N_45578);
and U45929 (N_45929,N_45635,N_45738);
nor U45930 (N_45930,N_45510,N_45694);
xor U45931 (N_45931,N_45661,N_45707);
or U45932 (N_45932,N_45514,N_45683);
and U45933 (N_45933,N_45599,N_45573);
xnor U45934 (N_45934,N_45711,N_45637);
nor U45935 (N_45935,N_45508,N_45748);
and U45936 (N_45936,N_45653,N_45702);
nand U45937 (N_45937,N_45722,N_45682);
and U45938 (N_45938,N_45637,N_45680);
nor U45939 (N_45939,N_45743,N_45726);
nor U45940 (N_45940,N_45598,N_45620);
nor U45941 (N_45941,N_45616,N_45505);
nor U45942 (N_45942,N_45629,N_45698);
or U45943 (N_45943,N_45647,N_45576);
and U45944 (N_45944,N_45701,N_45687);
and U45945 (N_45945,N_45659,N_45735);
xnor U45946 (N_45946,N_45731,N_45702);
xor U45947 (N_45947,N_45584,N_45700);
nand U45948 (N_45948,N_45696,N_45583);
nor U45949 (N_45949,N_45709,N_45626);
nor U45950 (N_45950,N_45576,N_45555);
nand U45951 (N_45951,N_45561,N_45598);
xnor U45952 (N_45952,N_45624,N_45734);
nor U45953 (N_45953,N_45526,N_45594);
or U45954 (N_45954,N_45666,N_45626);
nand U45955 (N_45955,N_45644,N_45612);
or U45956 (N_45956,N_45541,N_45687);
or U45957 (N_45957,N_45717,N_45612);
xor U45958 (N_45958,N_45600,N_45728);
and U45959 (N_45959,N_45607,N_45697);
nor U45960 (N_45960,N_45649,N_45654);
or U45961 (N_45961,N_45663,N_45729);
nand U45962 (N_45962,N_45544,N_45614);
nand U45963 (N_45963,N_45732,N_45659);
xor U45964 (N_45964,N_45582,N_45600);
or U45965 (N_45965,N_45693,N_45721);
nand U45966 (N_45966,N_45614,N_45514);
nand U45967 (N_45967,N_45545,N_45555);
or U45968 (N_45968,N_45608,N_45698);
nand U45969 (N_45969,N_45529,N_45604);
and U45970 (N_45970,N_45532,N_45593);
xor U45971 (N_45971,N_45500,N_45687);
or U45972 (N_45972,N_45539,N_45740);
nand U45973 (N_45973,N_45664,N_45513);
nor U45974 (N_45974,N_45584,N_45741);
and U45975 (N_45975,N_45680,N_45725);
xnor U45976 (N_45976,N_45525,N_45617);
nand U45977 (N_45977,N_45514,N_45736);
and U45978 (N_45978,N_45647,N_45601);
xor U45979 (N_45979,N_45645,N_45591);
nor U45980 (N_45980,N_45528,N_45536);
xnor U45981 (N_45981,N_45727,N_45589);
or U45982 (N_45982,N_45573,N_45729);
or U45983 (N_45983,N_45696,N_45632);
xor U45984 (N_45984,N_45592,N_45649);
xor U45985 (N_45985,N_45505,N_45523);
and U45986 (N_45986,N_45504,N_45561);
and U45987 (N_45987,N_45561,N_45702);
nor U45988 (N_45988,N_45621,N_45629);
nand U45989 (N_45989,N_45621,N_45640);
nor U45990 (N_45990,N_45542,N_45630);
nand U45991 (N_45991,N_45572,N_45520);
xor U45992 (N_45992,N_45511,N_45569);
and U45993 (N_45993,N_45581,N_45611);
nor U45994 (N_45994,N_45519,N_45531);
nor U45995 (N_45995,N_45615,N_45719);
nor U45996 (N_45996,N_45674,N_45557);
nand U45997 (N_45997,N_45556,N_45672);
nand U45998 (N_45998,N_45564,N_45734);
or U45999 (N_45999,N_45572,N_45674);
xnor U46000 (N_46000,N_45881,N_45979);
nand U46001 (N_46001,N_45770,N_45994);
xor U46002 (N_46002,N_45966,N_45781);
nor U46003 (N_46003,N_45952,N_45927);
nor U46004 (N_46004,N_45824,N_45884);
xor U46005 (N_46005,N_45838,N_45969);
xor U46006 (N_46006,N_45799,N_45803);
nor U46007 (N_46007,N_45834,N_45914);
nand U46008 (N_46008,N_45996,N_45883);
xor U46009 (N_46009,N_45783,N_45916);
nand U46010 (N_46010,N_45864,N_45887);
and U46011 (N_46011,N_45907,N_45797);
and U46012 (N_46012,N_45840,N_45868);
or U46013 (N_46013,N_45905,N_45791);
nor U46014 (N_46014,N_45826,N_45938);
and U46015 (N_46015,N_45839,N_45876);
nor U46016 (N_46016,N_45847,N_45829);
or U46017 (N_46017,N_45874,N_45936);
or U46018 (N_46018,N_45766,N_45873);
nand U46019 (N_46019,N_45946,N_45830);
or U46020 (N_46020,N_45971,N_45819);
nor U46021 (N_46021,N_45993,N_45769);
nor U46022 (N_46022,N_45764,N_45937);
xnor U46023 (N_46023,N_45816,N_45929);
nor U46024 (N_46024,N_45999,N_45855);
and U46025 (N_46025,N_45939,N_45871);
and U46026 (N_46026,N_45815,N_45942);
and U46027 (N_46027,N_45768,N_45856);
xor U46028 (N_46028,N_45957,N_45800);
and U46029 (N_46029,N_45825,N_45922);
nand U46030 (N_46030,N_45804,N_45915);
nand U46031 (N_46031,N_45885,N_45888);
nor U46032 (N_46032,N_45857,N_45982);
nand U46033 (N_46033,N_45980,N_45964);
or U46034 (N_46034,N_45755,N_45774);
and U46035 (N_46035,N_45894,N_45836);
nor U46036 (N_46036,N_45860,N_45763);
nor U46037 (N_46037,N_45990,N_45893);
and U46038 (N_46038,N_45794,N_45779);
nor U46039 (N_46039,N_45812,N_45924);
xnor U46040 (N_46040,N_45869,N_45778);
and U46041 (N_46041,N_45932,N_45806);
xor U46042 (N_46042,N_45817,N_45809);
xnor U46043 (N_46043,N_45968,N_45786);
nand U46044 (N_46044,N_45902,N_45911);
nor U46045 (N_46045,N_45882,N_45897);
nand U46046 (N_46046,N_45921,N_45933);
xor U46047 (N_46047,N_45899,N_45919);
xor U46048 (N_46048,N_45997,N_45841);
or U46049 (N_46049,N_45866,N_45992);
and U46050 (N_46050,N_45820,N_45962);
or U46051 (N_46051,N_45789,N_45947);
and U46052 (N_46052,N_45810,N_45998);
and U46053 (N_46053,N_45858,N_45782);
or U46054 (N_46054,N_45843,N_45772);
or U46055 (N_46055,N_45904,N_45891);
nand U46056 (N_46056,N_45879,N_45908);
and U46057 (N_46057,N_45977,N_45944);
xnor U46058 (N_46058,N_45945,N_45991);
and U46059 (N_46059,N_45978,N_45795);
nor U46060 (N_46060,N_45948,N_45928);
nor U46061 (N_46061,N_45961,N_45970);
or U46062 (N_46062,N_45975,N_45972);
nand U46063 (N_46063,N_45986,N_45833);
or U46064 (N_46064,N_45958,N_45818);
nand U46065 (N_46065,N_45828,N_45984);
nor U46066 (N_46066,N_45845,N_45777);
or U46067 (N_46067,N_45956,N_45935);
nand U46068 (N_46068,N_45923,N_45877);
nor U46069 (N_46069,N_45988,N_45918);
or U46070 (N_46070,N_45805,N_45790);
and U46071 (N_46071,N_45900,N_45762);
xor U46072 (N_46072,N_45949,N_45793);
and U46073 (N_46073,N_45852,N_45775);
nor U46074 (N_46074,N_45848,N_45925);
or U46075 (N_46075,N_45784,N_45951);
and U46076 (N_46076,N_45853,N_45807);
nand U46077 (N_46077,N_45837,N_45889);
xor U46078 (N_46078,N_45875,N_45759);
xnor U46079 (N_46079,N_45954,N_45813);
and U46080 (N_46080,N_45758,N_45796);
xor U46081 (N_46081,N_45880,N_45896);
nor U46082 (N_46082,N_45967,N_45846);
and U46083 (N_46083,N_45878,N_45859);
and U46084 (N_46084,N_45950,N_45854);
xor U46085 (N_46085,N_45771,N_45917);
and U46086 (N_46086,N_45912,N_45792);
nor U46087 (N_46087,N_45862,N_45913);
and U46088 (N_46088,N_45808,N_45898);
and U46089 (N_46089,N_45973,N_45785);
and U46090 (N_46090,N_45960,N_45821);
or U46091 (N_46091,N_45987,N_45850);
nand U46092 (N_46092,N_45831,N_45943);
nor U46093 (N_46093,N_45765,N_45801);
nand U46094 (N_46094,N_45940,N_45757);
xnor U46095 (N_46095,N_45963,N_45823);
xor U46096 (N_46096,N_45811,N_45776);
nor U46097 (N_46097,N_45865,N_45863);
or U46098 (N_46098,N_45798,N_45872);
or U46099 (N_46099,N_45959,N_45934);
and U46100 (N_46100,N_45985,N_45753);
or U46101 (N_46101,N_45751,N_45760);
xor U46102 (N_46102,N_45780,N_45903);
xor U46103 (N_46103,N_45920,N_45910);
nor U46104 (N_46104,N_45974,N_45953);
xnor U46105 (N_46105,N_45886,N_45761);
nor U46106 (N_46106,N_45835,N_45851);
and U46107 (N_46107,N_45981,N_45955);
and U46108 (N_46108,N_45754,N_45849);
nor U46109 (N_46109,N_45788,N_45983);
nand U46110 (N_46110,N_45767,N_45931);
or U46111 (N_46111,N_45895,N_45832);
or U46112 (N_46112,N_45909,N_45870);
and U46113 (N_46113,N_45890,N_45802);
or U46114 (N_46114,N_45756,N_45941);
nand U46115 (N_46115,N_45842,N_45787);
nand U46116 (N_46116,N_45827,N_45930);
nor U46117 (N_46117,N_45901,N_45822);
or U46118 (N_46118,N_45989,N_45861);
nand U46119 (N_46119,N_45892,N_45976);
and U46120 (N_46120,N_45965,N_45906);
nor U46121 (N_46121,N_45752,N_45844);
nor U46122 (N_46122,N_45814,N_45750);
xor U46123 (N_46123,N_45926,N_45867);
nand U46124 (N_46124,N_45773,N_45995);
xor U46125 (N_46125,N_45761,N_45920);
nand U46126 (N_46126,N_45937,N_45765);
nor U46127 (N_46127,N_45957,N_45987);
xor U46128 (N_46128,N_45912,N_45828);
nand U46129 (N_46129,N_45849,N_45819);
and U46130 (N_46130,N_45848,N_45775);
and U46131 (N_46131,N_45946,N_45808);
or U46132 (N_46132,N_45945,N_45759);
nand U46133 (N_46133,N_45912,N_45995);
nand U46134 (N_46134,N_45843,N_45756);
nand U46135 (N_46135,N_45891,N_45760);
nand U46136 (N_46136,N_45891,N_45814);
nor U46137 (N_46137,N_45824,N_45883);
nand U46138 (N_46138,N_45751,N_45842);
or U46139 (N_46139,N_45940,N_45810);
xor U46140 (N_46140,N_45808,N_45966);
or U46141 (N_46141,N_45827,N_45830);
xnor U46142 (N_46142,N_45756,N_45764);
nor U46143 (N_46143,N_45837,N_45792);
or U46144 (N_46144,N_45838,N_45976);
xor U46145 (N_46145,N_45896,N_45939);
xnor U46146 (N_46146,N_45798,N_45911);
xnor U46147 (N_46147,N_45985,N_45820);
or U46148 (N_46148,N_45784,N_45933);
nor U46149 (N_46149,N_45772,N_45783);
nor U46150 (N_46150,N_45784,N_45759);
or U46151 (N_46151,N_45998,N_45991);
and U46152 (N_46152,N_45962,N_45822);
and U46153 (N_46153,N_45914,N_45806);
and U46154 (N_46154,N_45871,N_45994);
or U46155 (N_46155,N_45807,N_45901);
or U46156 (N_46156,N_45788,N_45992);
or U46157 (N_46157,N_45910,N_45851);
or U46158 (N_46158,N_45963,N_45872);
nor U46159 (N_46159,N_45957,N_45771);
nor U46160 (N_46160,N_45878,N_45752);
xor U46161 (N_46161,N_45900,N_45996);
nor U46162 (N_46162,N_45947,N_45906);
nor U46163 (N_46163,N_45946,N_45956);
or U46164 (N_46164,N_45965,N_45818);
or U46165 (N_46165,N_45870,N_45897);
and U46166 (N_46166,N_45976,N_45822);
and U46167 (N_46167,N_45830,N_45860);
and U46168 (N_46168,N_45828,N_45842);
nand U46169 (N_46169,N_45854,N_45808);
xor U46170 (N_46170,N_45994,N_45896);
nor U46171 (N_46171,N_45930,N_45955);
or U46172 (N_46172,N_45929,N_45761);
xor U46173 (N_46173,N_45912,N_45965);
xnor U46174 (N_46174,N_45808,N_45846);
nand U46175 (N_46175,N_45963,N_45878);
nor U46176 (N_46176,N_45830,N_45954);
nor U46177 (N_46177,N_45773,N_45985);
xor U46178 (N_46178,N_45944,N_45813);
and U46179 (N_46179,N_45925,N_45856);
and U46180 (N_46180,N_45949,N_45890);
nor U46181 (N_46181,N_45936,N_45998);
nor U46182 (N_46182,N_45897,N_45943);
or U46183 (N_46183,N_45893,N_45922);
and U46184 (N_46184,N_45779,N_45808);
xnor U46185 (N_46185,N_45813,N_45872);
nor U46186 (N_46186,N_45983,N_45949);
or U46187 (N_46187,N_45925,N_45992);
or U46188 (N_46188,N_45803,N_45772);
or U46189 (N_46189,N_45789,N_45980);
nor U46190 (N_46190,N_45932,N_45824);
nand U46191 (N_46191,N_45761,N_45825);
and U46192 (N_46192,N_45876,N_45924);
nand U46193 (N_46193,N_45889,N_45929);
or U46194 (N_46194,N_45883,N_45832);
or U46195 (N_46195,N_45987,N_45782);
or U46196 (N_46196,N_45851,N_45994);
or U46197 (N_46197,N_45763,N_45764);
nand U46198 (N_46198,N_45757,N_45882);
and U46199 (N_46199,N_45758,N_45800);
xnor U46200 (N_46200,N_45891,N_45862);
xor U46201 (N_46201,N_45819,N_45775);
xor U46202 (N_46202,N_45823,N_45995);
xor U46203 (N_46203,N_45886,N_45955);
nor U46204 (N_46204,N_45902,N_45915);
xor U46205 (N_46205,N_45819,N_45796);
nand U46206 (N_46206,N_45806,N_45794);
or U46207 (N_46207,N_45819,N_45915);
or U46208 (N_46208,N_45840,N_45879);
xor U46209 (N_46209,N_45819,N_45936);
or U46210 (N_46210,N_45825,N_45752);
or U46211 (N_46211,N_45793,N_45859);
nor U46212 (N_46212,N_45841,N_45874);
or U46213 (N_46213,N_45936,N_45905);
and U46214 (N_46214,N_45891,N_45906);
nand U46215 (N_46215,N_45808,N_45954);
nand U46216 (N_46216,N_45978,N_45800);
or U46217 (N_46217,N_45791,N_45906);
nand U46218 (N_46218,N_45751,N_45840);
or U46219 (N_46219,N_45877,N_45934);
or U46220 (N_46220,N_45896,N_45782);
nor U46221 (N_46221,N_45945,N_45890);
or U46222 (N_46222,N_45982,N_45847);
nand U46223 (N_46223,N_45796,N_45929);
and U46224 (N_46224,N_45927,N_45892);
nand U46225 (N_46225,N_45756,N_45897);
nand U46226 (N_46226,N_45819,N_45784);
nor U46227 (N_46227,N_45889,N_45999);
nor U46228 (N_46228,N_45933,N_45853);
or U46229 (N_46229,N_45919,N_45864);
or U46230 (N_46230,N_45955,N_45986);
xnor U46231 (N_46231,N_45977,N_45961);
and U46232 (N_46232,N_45867,N_45954);
xor U46233 (N_46233,N_45789,N_45780);
nor U46234 (N_46234,N_45912,N_45832);
and U46235 (N_46235,N_45884,N_45878);
xnor U46236 (N_46236,N_45900,N_45903);
or U46237 (N_46237,N_45816,N_45796);
nor U46238 (N_46238,N_45911,N_45837);
or U46239 (N_46239,N_45996,N_45766);
and U46240 (N_46240,N_45912,N_45839);
xor U46241 (N_46241,N_45818,N_45891);
or U46242 (N_46242,N_45818,N_45780);
or U46243 (N_46243,N_45783,N_45924);
nand U46244 (N_46244,N_45818,N_45882);
xor U46245 (N_46245,N_45793,N_45751);
nor U46246 (N_46246,N_45791,N_45944);
or U46247 (N_46247,N_45786,N_45801);
nor U46248 (N_46248,N_45761,N_45758);
xnor U46249 (N_46249,N_45776,N_45751);
nand U46250 (N_46250,N_46083,N_46119);
or U46251 (N_46251,N_46167,N_46131);
and U46252 (N_46252,N_46244,N_46220);
or U46253 (N_46253,N_46198,N_46004);
and U46254 (N_46254,N_46005,N_46028);
nor U46255 (N_46255,N_46066,N_46030);
and U46256 (N_46256,N_46090,N_46176);
nand U46257 (N_46257,N_46128,N_46126);
nor U46258 (N_46258,N_46000,N_46201);
or U46259 (N_46259,N_46029,N_46241);
or U46260 (N_46260,N_46008,N_46155);
nand U46261 (N_46261,N_46067,N_46037);
xor U46262 (N_46262,N_46209,N_46001);
or U46263 (N_46263,N_46012,N_46200);
and U46264 (N_46264,N_46020,N_46211);
nor U46265 (N_46265,N_46084,N_46183);
or U46266 (N_46266,N_46044,N_46113);
or U46267 (N_46267,N_46153,N_46073);
xor U46268 (N_46268,N_46069,N_46058);
nor U46269 (N_46269,N_46196,N_46237);
nand U46270 (N_46270,N_46009,N_46079);
or U46271 (N_46271,N_46230,N_46129);
nand U46272 (N_46272,N_46227,N_46181);
nor U46273 (N_46273,N_46208,N_46043);
nor U46274 (N_46274,N_46135,N_46142);
nand U46275 (N_46275,N_46236,N_46015);
nor U46276 (N_46276,N_46110,N_46192);
nor U46277 (N_46277,N_46248,N_46242);
or U46278 (N_46278,N_46074,N_46007);
nor U46279 (N_46279,N_46046,N_46111);
nand U46280 (N_46280,N_46053,N_46089);
xor U46281 (N_46281,N_46085,N_46228);
and U46282 (N_46282,N_46166,N_46042);
or U46283 (N_46283,N_46162,N_46086);
nand U46284 (N_46284,N_46231,N_46062);
nand U46285 (N_46285,N_46134,N_46077);
and U46286 (N_46286,N_46050,N_46082);
nor U46287 (N_46287,N_46097,N_46114);
nor U46288 (N_46288,N_46213,N_46061);
nand U46289 (N_46289,N_46212,N_46091);
nor U46290 (N_46290,N_46202,N_46027);
or U46291 (N_46291,N_46179,N_46094);
or U46292 (N_46292,N_46141,N_46187);
nor U46293 (N_46293,N_46222,N_46099);
nor U46294 (N_46294,N_46139,N_46022);
nand U46295 (N_46295,N_46133,N_46239);
nor U46296 (N_46296,N_46055,N_46190);
nor U46297 (N_46297,N_46019,N_46123);
and U46298 (N_46298,N_46217,N_46189);
xnor U46299 (N_46299,N_46148,N_46108);
nor U46300 (N_46300,N_46151,N_46138);
or U46301 (N_46301,N_46117,N_46068);
or U46302 (N_46302,N_46021,N_46040);
xnor U46303 (N_46303,N_46188,N_46232);
xnor U46304 (N_46304,N_46011,N_46218);
xor U46305 (N_46305,N_46240,N_46064);
or U46306 (N_46306,N_46223,N_46057);
nand U46307 (N_46307,N_46178,N_46070);
nor U46308 (N_46308,N_46080,N_46137);
or U46309 (N_46309,N_46168,N_46229);
nor U46310 (N_46310,N_46049,N_46101);
or U46311 (N_46311,N_46034,N_46159);
or U46312 (N_46312,N_46075,N_46249);
xnor U46313 (N_46313,N_46130,N_46065);
and U46314 (N_46314,N_46197,N_46087);
nand U46315 (N_46315,N_46127,N_46039);
and U46316 (N_46316,N_46225,N_46163);
and U46317 (N_46317,N_46165,N_46018);
or U46318 (N_46318,N_46184,N_46052);
nand U46319 (N_46319,N_46059,N_46194);
nor U46320 (N_46320,N_46045,N_46247);
nand U46321 (N_46321,N_46032,N_46072);
xnor U46322 (N_46322,N_46233,N_46016);
nor U46323 (N_46323,N_46054,N_46103);
or U46324 (N_46324,N_46243,N_46010);
nor U46325 (N_46325,N_46149,N_46164);
nor U46326 (N_46326,N_46150,N_46100);
and U46327 (N_46327,N_46158,N_46105);
and U46328 (N_46328,N_46206,N_46109);
nand U46329 (N_46329,N_46203,N_46026);
xor U46330 (N_46330,N_46112,N_46060);
nor U46331 (N_46331,N_46122,N_46098);
xnor U46332 (N_46332,N_46219,N_46147);
and U46333 (N_46333,N_46156,N_46003);
nand U46334 (N_46334,N_46047,N_46199);
xor U46335 (N_46335,N_46093,N_46014);
nor U46336 (N_46336,N_46170,N_46136);
nand U46337 (N_46337,N_46171,N_46144);
and U46338 (N_46338,N_46246,N_46193);
and U46339 (N_46339,N_46025,N_46107);
xnor U46340 (N_46340,N_46140,N_46116);
xor U46341 (N_46341,N_46121,N_46161);
nor U46342 (N_46342,N_46185,N_46175);
or U46343 (N_46343,N_46132,N_46186);
nand U46344 (N_46344,N_46235,N_46088);
nand U46345 (N_46345,N_46157,N_46017);
xnor U46346 (N_46346,N_46048,N_46078);
nor U46347 (N_46347,N_46238,N_46195);
and U46348 (N_46348,N_46013,N_46115);
or U46349 (N_46349,N_46102,N_46031);
nor U46350 (N_46350,N_46104,N_46076);
nor U46351 (N_46351,N_46146,N_46180);
or U46352 (N_46352,N_46063,N_46124);
or U46353 (N_46353,N_46224,N_46154);
and U46354 (N_46354,N_46174,N_46120);
and U46355 (N_46355,N_46071,N_46033);
nor U46356 (N_46356,N_46152,N_46036);
nor U46357 (N_46357,N_46056,N_46081);
nand U46358 (N_46358,N_46177,N_46118);
xnor U46359 (N_46359,N_46172,N_46234);
and U46360 (N_46360,N_46207,N_46051);
and U46361 (N_46361,N_46173,N_46226);
nand U46362 (N_46362,N_46041,N_46214);
xnor U46363 (N_46363,N_46216,N_46160);
nor U46364 (N_46364,N_46095,N_46002);
nand U46365 (N_46365,N_46023,N_46169);
and U46366 (N_46366,N_46096,N_46205);
nor U46367 (N_46367,N_46245,N_46215);
xor U46368 (N_46368,N_46092,N_46035);
xnor U46369 (N_46369,N_46024,N_46143);
nand U46370 (N_46370,N_46210,N_46182);
xnor U46371 (N_46371,N_46204,N_46038);
nor U46372 (N_46372,N_46191,N_46106);
and U46373 (N_46373,N_46125,N_46006);
or U46374 (N_46374,N_46145,N_46221);
and U46375 (N_46375,N_46247,N_46022);
nor U46376 (N_46376,N_46204,N_46048);
nor U46377 (N_46377,N_46034,N_46009);
or U46378 (N_46378,N_46234,N_46089);
xnor U46379 (N_46379,N_46242,N_46030);
nand U46380 (N_46380,N_46054,N_46186);
nand U46381 (N_46381,N_46173,N_46042);
or U46382 (N_46382,N_46127,N_46194);
and U46383 (N_46383,N_46072,N_46156);
nand U46384 (N_46384,N_46188,N_46215);
and U46385 (N_46385,N_46065,N_46207);
nand U46386 (N_46386,N_46237,N_46212);
nor U46387 (N_46387,N_46067,N_46083);
or U46388 (N_46388,N_46050,N_46159);
or U46389 (N_46389,N_46193,N_46112);
nand U46390 (N_46390,N_46123,N_46119);
or U46391 (N_46391,N_46060,N_46036);
or U46392 (N_46392,N_46199,N_46114);
nor U46393 (N_46393,N_46239,N_46169);
nand U46394 (N_46394,N_46167,N_46038);
nand U46395 (N_46395,N_46216,N_46243);
or U46396 (N_46396,N_46244,N_46144);
nor U46397 (N_46397,N_46034,N_46237);
nand U46398 (N_46398,N_46034,N_46153);
xnor U46399 (N_46399,N_46080,N_46204);
nand U46400 (N_46400,N_46067,N_46124);
or U46401 (N_46401,N_46025,N_46177);
or U46402 (N_46402,N_46239,N_46030);
nor U46403 (N_46403,N_46175,N_46096);
and U46404 (N_46404,N_46087,N_46084);
xor U46405 (N_46405,N_46082,N_46249);
nand U46406 (N_46406,N_46249,N_46045);
nand U46407 (N_46407,N_46234,N_46222);
nor U46408 (N_46408,N_46029,N_46224);
nor U46409 (N_46409,N_46125,N_46164);
and U46410 (N_46410,N_46033,N_46045);
xnor U46411 (N_46411,N_46156,N_46181);
xor U46412 (N_46412,N_46225,N_46051);
and U46413 (N_46413,N_46241,N_46151);
xnor U46414 (N_46414,N_46135,N_46198);
nor U46415 (N_46415,N_46020,N_46100);
nand U46416 (N_46416,N_46012,N_46209);
xor U46417 (N_46417,N_46151,N_46226);
nor U46418 (N_46418,N_46100,N_46104);
or U46419 (N_46419,N_46127,N_46213);
nand U46420 (N_46420,N_46233,N_46057);
xor U46421 (N_46421,N_46224,N_46203);
nand U46422 (N_46422,N_46019,N_46085);
and U46423 (N_46423,N_46199,N_46090);
and U46424 (N_46424,N_46044,N_46110);
xor U46425 (N_46425,N_46199,N_46239);
nand U46426 (N_46426,N_46136,N_46040);
or U46427 (N_46427,N_46054,N_46094);
and U46428 (N_46428,N_46207,N_46102);
and U46429 (N_46429,N_46238,N_46206);
nor U46430 (N_46430,N_46180,N_46122);
xor U46431 (N_46431,N_46183,N_46094);
xnor U46432 (N_46432,N_46039,N_46146);
or U46433 (N_46433,N_46069,N_46245);
or U46434 (N_46434,N_46133,N_46020);
nand U46435 (N_46435,N_46018,N_46228);
xnor U46436 (N_46436,N_46100,N_46230);
and U46437 (N_46437,N_46021,N_46126);
or U46438 (N_46438,N_46200,N_46036);
xnor U46439 (N_46439,N_46027,N_46056);
xnor U46440 (N_46440,N_46040,N_46236);
or U46441 (N_46441,N_46206,N_46210);
nor U46442 (N_46442,N_46238,N_46091);
and U46443 (N_46443,N_46015,N_46110);
and U46444 (N_46444,N_46245,N_46140);
nand U46445 (N_46445,N_46052,N_46042);
nor U46446 (N_46446,N_46095,N_46121);
and U46447 (N_46447,N_46149,N_46228);
or U46448 (N_46448,N_46150,N_46096);
and U46449 (N_46449,N_46001,N_46124);
nand U46450 (N_46450,N_46001,N_46195);
nand U46451 (N_46451,N_46085,N_46174);
and U46452 (N_46452,N_46155,N_46150);
or U46453 (N_46453,N_46115,N_46113);
and U46454 (N_46454,N_46142,N_46005);
xor U46455 (N_46455,N_46051,N_46196);
and U46456 (N_46456,N_46030,N_46043);
or U46457 (N_46457,N_46086,N_46082);
xor U46458 (N_46458,N_46110,N_46161);
or U46459 (N_46459,N_46006,N_46248);
xor U46460 (N_46460,N_46151,N_46014);
nor U46461 (N_46461,N_46044,N_46187);
nor U46462 (N_46462,N_46000,N_46048);
nor U46463 (N_46463,N_46060,N_46081);
or U46464 (N_46464,N_46216,N_46061);
and U46465 (N_46465,N_46126,N_46012);
or U46466 (N_46466,N_46231,N_46027);
nor U46467 (N_46467,N_46146,N_46036);
xor U46468 (N_46468,N_46070,N_46200);
xor U46469 (N_46469,N_46004,N_46235);
nor U46470 (N_46470,N_46227,N_46062);
or U46471 (N_46471,N_46004,N_46212);
nor U46472 (N_46472,N_46220,N_46229);
or U46473 (N_46473,N_46211,N_46213);
xor U46474 (N_46474,N_46187,N_46247);
xor U46475 (N_46475,N_46242,N_46218);
nor U46476 (N_46476,N_46030,N_46188);
xor U46477 (N_46477,N_46108,N_46092);
xnor U46478 (N_46478,N_46216,N_46186);
and U46479 (N_46479,N_46235,N_46114);
or U46480 (N_46480,N_46031,N_46188);
nor U46481 (N_46481,N_46228,N_46208);
nand U46482 (N_46482,N_46054,N_46073);
xor U46483 (N_46483,N_46233,N_46241);
nand U46484 (N_46484,N_46072,N_46041);
and U46485 (N_46485,N_46155,N_46196);
nand U46486 (N_46486,N_46056,N_46181);
and U46487 (N_46487,N_46031,N_46158);
xnor U46488 (N_46488,N_46205,N_46005);
or U46489 (N_46489,N_46006,N_46141);
nor U46490 (N_46490,N_46096,N_46117);
nor U46491 (N_46491,N_46089,N_46130);
nand U46492 (N_46492,N_46025,N_46225);
or U46493 (N_46493,N_46069,N_46201);
xnor U46494 (N_46494,N_46162,N_46051);
nand U46495 (N_46495,N_46058,N_46192);
xor U46496 (N_46496,N_46108,N_46219);
or U46497 (N_46497,N_46249,N_46027);
xnor U46498 (N_46498,N_46182,N_46126);
nand U46499 (N_46499,N_46247,N_46100);
nor U46500 (N_46500,N_46448,N_46263);
xor U46501 (N_46501,N_46378,N_46363);
or U46502 (N_46502,N_46458,N_46439);
nand U46503 (N_46503,N_46321,N_46408);
nand U46504 (N_46504,N_46401,N_46487);
or U46505 (N_46505,N_46306,N_46445);
nand U46506 (N_46506,N_46496,N_46340);
or U46507 (N_46507,N_46261,N_46283);
nand U46508 (N_46508,N_46426,N_46260);
or U46509 (N_46509,N_46419,N_46277);
or U46510 (N_46510,N_46392,N_46383);
nor U46511 (N_46511,N_46410,N_46351);
xnor U46512 (N_46512,N_46387,N_46299);
or U46513 (N_46513,N_46380,N_46343);
or U46514 (N_46514,N_46362,N_46279);
nor U46515 (N_46515,N_46434,N_46313);
nand U46516 (N_46516,N_46368,N_46305);
xor U46517 (N_46517,N_46457,N_46379);
and U46518 (N_46518,N_46270,N_46485);
nor U46519 (N_46519,N_46269,N_46477);
xor U46520 (N_46520,N_46395,N_46294);
nor U46521 (N_46521,N_46451,N_46338);
nand U46522 (N_46522,N_46390,N_46267);
and U46523 (N_46523,N_46266,N_46255);
nor U46524 (N_46524,N_46280,N_46354);
or U46525 (N_46525,N_46455,N_46394);
or U46526 (N_46526,N_46365,N_46356);
nor U46527 (N_46527,N_46274,N_46484);
nand U46528 (N_46528,N_46251,N_46353);
or U46529 (N_46529,N_46418,N_46323);
and U46530 (N_46530,N_46435,N_46403);
nor U46531 (N_46531,N_46406,N_46427);
and U46532 (N_46532,N_46495,N_46300);
xnor U46533 (N_46533,N_46320,N_46254);
nand U46534 (N_46534,N_46428,N_46498);
nor U46535 (N_46535,N_46326,N_46311);
or U46536 (N_46536,N_46259,N_46480);
nor U46537 (N_46537,N_46492,N_46405);
and U46538 (N_46538,N_46440,N_46465);
nor U46539 (N_46539,N_46339,N_46268);
xor U46540 (N_46540,N_46384,N_46472);
xnor U46541 (N_46541,N_46296,N_46377);
or U46542 (N_46542,N_46331,N_46358);
and U46543 (N_46543,N_46497,N_46286);
and U46544 (N_46544,N_46417,N_46437);
and U46545 (N_46545,N_46290,N_46342);
nand U46546 (N_46546,N_46402,N_46415);
nor U46547 (N_46547,N_46275,N_46471);
nand U46548 (N_46548,N_46337,N_46468);
or U46549 (N_46549,N_46292,N_46304);
and U46550 (N_46550,N_46287,N_46295);
nand U46551 (N_46551,N_46470,N_46348);
nand U46552 (N_46552,N_46398,N_46493);
xor U46553 (N_46553,N_46265,N_46316);
and U46554 (N_46554,N_46454,N_46341);
and U46555 (N_46555,N_46271,N_46360);
nor U46556 (N_46556,N_46324,N_46361);
xnor U46557 (N_46557,N_46346,N_46258);
and U46558 (N_46558,N_46312,N_46262);
or U46559 (N_46559,N_46281,N_46335);
nor U46560 (N_46560,N_46463,N_46499);
or U46561 (N_46561,N_46278,N_46328);
nand U46562 (N_46562,N_46310,N_46303);
or U46563 (N_46563,N_46476,N_46386);
or U46564 (N_46564,N_46462,N_46433);
and U46565 (N_46565,N_46489,N_46413);
xnor U46566 (N_46566,N_46332,N_46317);
nor U46567 (N_46567,N_46293,N_46357);
and U46568 (N_46568,N_46285,N_46309);
and U46569 (N_46569,N_46449,N_46284);
or U46570 (N_46570,N_46443,N_46336);
nand U46571 (N_46571,N_46441,N_46432);
nand U46572 (N_46572,N_46371,N_46327);
or U46573 (N_46573,N_46399,N_46344);
nor U46574 (N_46574,N_46431,N_46416);
nor U46575 (N_46575,N_46414,N_46474);
xnor U46576 (N_46576,N_46404,N_46456);
and U46577 (N_46577,N_46264,N_46375);
nand U46578 (N_46578,N_46481,N_46400);
or U46579 (N_46579,N_46486,N_46257);
xor U46580 (N_46580,N_46430,N_46425);
or U46581 (N_46581,N_46393,N_46288);
nand U46582 (N_46582,N_46330,N_46314);
xnor U46583 (N_46583,N_46355,N_46478);
nand U46584 (N_46584,N_46315,N_46301);
xor U46585 (N_46585,N_46420,N_46329);
nor U46586 (N_46586,N_46396,N_46411);
xnor U46587 (N_46587,N_46479,N_46372);
or U46588 (N_46588,N_46482,N_46429);
nand U46589 (N_46589,N_46438,N_46494);
nor U46590 (N_46590,N_46289,N_46488);
nand U46591 (N_46591,N_46446,N_46407);
nand U46592 (N_46592,N_46308,N_46307);
and U46593 (N_46593,N_46453,N_46318);
xor U46594 (N_46594,N_46276,N_46412);
or U46595 (N_46595,N_46272,N_46391);
nand U46596 (N_46596,N_46349,N_46491);
or U46597 (N_46597,N_46347,N_46452);
nand U46598 (N_46598,N_46469,N_46250);
nand U46599 (N_46599,N_46352,N_46291);
or U46600 (N_46600,N_46388,N_46381);
and U46601 (N_46601,N_46422,N_46459);
xnor U46602 (N_46602,N_46373,N_46298);
nor U46603 (N_46603,N_46334,N_46302);
or U46604 (N_46604,N_46376,N_46467);
nand U46605 (N_46605,N_46366,N_46442);
nand U46606 (N_46606,N_46475,N_46370);
nand U46607 (N_46607,N_46333,N_46367);
xnor U46608 (N_46608,N_46460,N_46483);
nand U46609 (N_46609,N_46444,N_46350);
nand U46610 (N_46610,N_46450,N_46421);
xor U46611 (N_46611,N_46447,N_46273);
and U46612 (N_46612,N_46461,N_46374);
and U46613 (N_46613,N_46466,N_46490);
nor U46614 (N_46614,N_46424,N_46389);
nor U46615 (N_46615,N_46385,N_46282);
nand U46616 (N_46616,N_46297,N_46359);
or U46617 (N_46617,N_46256,N_46436);
xor U46618 (N_46618,N_46397,N_46319);
xor U46619 (N_46619,N_46252,N_46325);
or U46620 (N_46620,N_46322,N_46382);
nand U46621 (N_46621,N_46369,N_46409);
and U46622 (N_46622,N_46464,N_46345);
and U46623 (N_46623,N_46364,N_46253);
nor U46624 (N_46624,N_46423,N_46473);
nand U46625 (N_46625,N_46489,N_46336);
nor U46626 (N_46626,N_46457,N_46389);
and U46627 (N_46627,N_46491,N_46485);
nor U46628 (N_46628,N_46498,N_46283);
and U46629 (N_46629,N_46463,N_46293);
xnor U46630 (N_46630,N_46419,N_46267);
and U46631 (N_46631,N_46454,N_46312);
nor U46632 (N_46632,N_46380,N_46315);
or U46633 (N_46633,N_46479,N_46348);
xnor U46634 (N_46634,N_46280,N_46305);
and U46635 (N_46635,N_46436,N_46468);
and U46636 (N_46636,N_46406,N_46432);
and U46637 (N_46637,N_46359,N_46344);
nand U46638 (N_46638,N_46281,N_46493);
and U46639 (N_46639,N_46262,N_46320);
nand U46640 (N_46640,N_46274,N_46494);
xnor U46641 (N_46641,N_46282,N_46439);
nor U46642 (N_46642,N_46372,N_46250);
and U46643 (N_46643,N_46409,N_46482);
nand U46644 (N_46644,N_46479,N_46487);
or U46645 (N_46645,N_46282,N_46493);
or U46646 (N_46646,N_46261,N_46300);
and U46647 (N_46647,N_46484,N_46363);
and U46648 (N_46648,N_46306,N_46444);
xnor U46649 (N_46649,N_46400,N_46272);
nor U46650 (N_46650,N_46438,N_46282);
or U46651 (N_46651,N_46466,N_46471);
nor U46652 (N_46652,N_46272,N_46350);
nand U46653 (N_46653,N_46466,N_46497);
and U46654 (N_46654,N_46443,N_46354);
or U46655 (N_46655,N_46351,N_46298);
xor U46656 (N_46656,N_46338,N_46259);
nor U46657 (N_46657,N_46262,N_46406);
and U46658 (N_46658,N_46313,N_46262);
or U46659 (N_46659,N_46393,N_46476);
or U46660 (N_46660,N_46456,N_46366);
xor U46661 (N_46661,N_46352,N_46283);
or U46662 (N_46662,N_46323,N_46425);
xor U46663 (N_46663,N_46305,N_46285);
xnor U46664 (N_46664,N_46405,N_46254);
xnor U46665 (N_46665,N_46410,N_46438);
xor U46666 (N_46666,N_46289,N_46446);
and U46667 (N_46667,N_46395,N_46470);
nor U46668 (N_46668,N_46303,N_46367);
and U46669 (N_46669,N_46430,N_46474);
nand U46670 (N_46670,N_46315,N_46480);
nand U46671 (N_46671,N_46484,N_46277);
and U46672 (N_46672,N_46268,N_46406);
or U46673 (N_46673,N_46325,N_46469);
nand U46674 (N_46674,N_46329,N_46476);
or U46675 (N_46675,N_46352,N_46447);
and U46676 (N_46676,N_46289,N_46485);
or U46677 (N_46677,N_46276,N_46336);
and U46678 (N_46678,N_46308,N_46354);
xor U46679 (N_46679,N_46484,N_46469);
xor U46680 (N_46680,N_46449,N_46393);
nand U46681 (N_46681,N_46255,N_46360);
nand U46682 (N_46682,N_46481,N_46407);
and U46683 (N_46683,N_46492,N_46255);
xnor U46684 (N_46684,N_46361,N_46275);
or U46685 (N_46685,N_46385,N_46287);
and U46686 (N_46686,N_46416,N_46483);
or U46687 (N_46687,N_46489,N_46396);
nor U46688 (N_46688,N_46435,N_46313);
and U46689 (N_46689,N_46450,N_46268);
and U46690 (N_46690,N_46388,N_46429);
xor U46691 (N_46691,N_46460,N_46492);
and U46692 (N_46692,N_46279,N_46433);
and U46693 (N_46693,N_46346,N_46388);
xnor U46694 (N_46694,N_46479,N_46374);
and U46695 (N_46695,N_46369,N_46330);
nor U46696 (N_46696,N_46456,N_46350);
nor U46697 (N_46697,N_46430,N_46435);
xor U46698 (N_46698,N_46251,N_46422);
or U46699 (N_46699,N_46264,N_46294);
nand U46700 (N_46700,N_46302,N_46482);
xnor U46701 (N_46701,N_46321,N_46457);
or U46702 (N_46702,N_46272,N_46279);
nor U46703 (N_46703,N_46309,N_46292);
xor U46704 (N_46704,N_46295,N_46290);
and U46705 (N_46705,N_46375,N_46418);
xor U46706 (N_46706,N_46301,N_46337);
nand U46707 (N_46707,N_46258,N_46298);
xor U46708 (N_46708,N_46457,N_46316);
nand U46709 (N_46709,N_46307,N_46362);
nand U46710 (N_46710,N_46463,N_46259);
nor U46711 (N_46711,N_46351,N_46282);
or U46712 (N_46712,N_46250,N_46394);
and U46713 (N_46713,N_46397,N_46436);
or U46714 (N_46714,N_46392,N_46256);
or U46715 (N_46715,N_46399,N_46435);
nand U46716 (N_46716,N_46270,N_46301);
and U46717 (N_46717,N_46404,N_46410);
xnor U46718 (N_46718,N_46435,N_46340);
nor U46719 (N_46719,N_46435,N_46492);
and U46720 (N_46720,N_46315,N_46430);
nor U46721 (N_46721,N_46381,N_46484);
and U46722 (N_46722,N_46286,N_46343);
xor U46723 (N_46723,N_46407,N_46444);
nand U46724 (N_46724,N_46401,N_46362);
xnor U46725 (N_46725,N_46468,N_46489);
xnor U46726 (N_46726,N_46444,N_46420);
and U46727 (N_46727,N_46401,N_46336);
or U46728 (N_46728,N_46461,N_46457);
xnor U46729 (N_46729,N_46260,N_46466);
nor U46730 (N_46730,N_46372,N_46354);
or U46731 (N_46731,N_46480,N_46442);
and U46732 (N_46732,N_46349,N_46266);
or U46733 (N_46733,N_46357,N_46485);
nand U46734 (N_46734,N_46415,N_46394);
nand U46735 (N_46735,N_46271,N_46411);
xnor U46736 (N_46736,N_46286,N_46455);
nand U46737 (N_46737,N_46380,N_46273);
and U46738 (N_46738,N_46287,N_46338);
and U46739 (N_46739,N_46353,N_46284);
nand U46740 (N_46740,N_46456,N_46483);
or U46741 (N_46741,N_46401,N_46333);
nor U46742 (N_46742,N_46455,N_46328);
nand U46743 (N_46743,N_46496,N_46390);
nand U46744 (N_46744,N_46437,N_46485);
and U46745 (N_46745,N_46346,N_46430);
and U46746 (N_46746,N_46400,N_46366);
nand U46747 (N_46747,N_46325,N_46392);
xnor U46748 (N_46748,N_46443,N_46462);
nor U46749 (N_46749,N_46488,N_46359);
nor U46750 (N_46750,N_46748,N_46681);
nor U46751 (N_46751,N_46527,N_46691);
or U46752 (N_46752,N_46725,N_46513);
or U46753 (N_46753,N_46721,N_46720);
and U46754 (N_46754,N_46517,N_46736);
or U46755 (N_46755,N_46652,N_46533);
nor U46756 (N_46756,N_46603,N_46653);
nor U46757 (N_46757,N_46698,N_46616);
nand U46758 (N_46758,N_46705,N_46742);
xor U46759 (N_46759,N_46545,N_46581);
nand U46760 (N_46760,N_46638,N_46628);
or U46761 (N_46761,N_46646,N_46554);
xor U46762 (N_46762,N_46682,N_46683);
nand U46763 (N_46763,N_46696,N_46669);
and U46764 (N_46764,N_46728,N_46663);
and U46765 (N_46765,N_46589,N_46650);
nand U46766 (N_46766,N_46621,N_46578);
nor U46767 (N_46767,N_46654,N_46657);
nand U46768 (N_46768,N_46609,N_46747);
xnor U46769 (N_46769,N_46717,N_46511);
and U46770 (N_46770,N_46604,N_46636);
xor U46771 (N_46771,N_46695,N_46660);
xnor U46772 (N_46772,N_46735,N_46532);
xnor U46773 (N_46773,N_46711,N_46679);
xnor U46774 (N_46774,N_46600,N_46644);
and U46775 (N_46775,N_46559,N_46744);
or U46776 (N_46776,N_46643,N_46536);
and U46777 (N_46777,N_46686,N_46521);
or U46778 (N_46778,N_46631,N_46667);
nand U46779 (N_46779,N_46731,N_46700);
xor U46780 (N_46780,N_46633,N_46706);
nand U46781 (N_46781,N_46671,N_46707);
and U46782 (N_46782,N_46719,N_46535);
nand U46783 (N_46783,N_46557,N_46541);
xnor U46784 (N_46784,N_46555,N_46592);
or U46785 (N_46785,N_46526,N_46516);
nand U46786 (N_46786,N_46637,N_46551);
nand U46787 (N_46787,N_46503,N_46568);
nor U46788 (N_46788,N_46739,N_46576);
nor U46789 (N_46789,N_46531,N_46656);
and U46790 (N_46790,N_46665,N_46699);
xor U46791 (N_46791,N_46632,N_46709);
nor U46792 (N_46792,N_46522,N_46701);
nand U46793 (N_46793,N_46585,N_46680);
nand U46794 (N_46794,N_46710,N_46666);
nand U46795 (N_46795,N_46583,N_46587);
nand U46796 (N_46796,N_46602,N_46546);
or U46797 (N_46797,N_46722,N_46505);
nor U46798 (N_46798,N_46726,N_46595);
xnor U46799 (N_46799,N_46718,N_46504);
nand U46800 (N_46800,N_46509,N_46528);
nand U46801 (N_46801,N_46740,N_46689);
nand U46802 (N_46802,N_46525,N_46569);
nor U46803 (N_46803,N_46712,N_46534);
nand U46804 (N_46804,N_46713,N_46601);
and U46805 (N_46805,N_46745,N_46529);
nand U46806 (N_46806,N_46561,N_46574);
nand U46807 (N_46807,N_46606,N_46550);
or U46808 (N_46808,N_46512,N_46625);
xor U46809 (N_46809,N_46743,N_46539);
and U46810 (N_46810,N_46641,N_46697);
xor U46811 (N_46811,N_46708,N_46501);
nand U46812 (N_46812,N_46730,N_46684);
and U46813 (N_46813,N_46618,N_46677);
xor U46814 (N_46814,N_46664,N_46548);
nand U46815 (N_46815,N_46508,N_46577);
nand U46816 (N_46816,N_46614,N_46579);
or U46817 (N_46817,N_46615,N_46540);
nand U46818 (N_46818,N_46630,N_46693);
nand U46819 (N_46819,N_46692,N_46611);
nor U46820 (N_46820,N_46596,N_46694);
or U46821 (N_46821,N_46746,N_46563);
or U46822 (N_46822,N_46582,N_46562);
and U46823 (N_46823,N_46715,N_46586);
nor U46824 (N_46824,N_46688,N_46560);
and U46825 (N_46825,N_46594,N_46617);
xor U46826 (N_46826,N_46515,N_46507);
or U46827 (N_46827,N_46510,N_46659);
or U46828 (N_46828,N_46687,N_46553);
nor U46829 (N_46829,N_46599,N_46538);
xor U46830 (N_46830,N_46724,N_46518);
xor U46831 (N_46831,N_46607,N_46702);
xor U46832 (N_46832,N_46678,N_46704);
nand U46833 (N_46833,N_46591,N_46658);
or U46834 (N_46834,N_46627,N_46542);
xnor U46835 (N_46835,N_46703,N_46670);
or U46836 (N_46836,N_46514,N_46613);
xnor U46837 (N_46837,N_46619,N_46610);
and U46838 (N_46838,N_46634,N_46584);
nor U46839 (N_46839,N_46737,N_46523);
and U46840 (N_46840,N_46570,N_46575);
xor U46841 (N_46841,N_46605,N_46598);
and U46842 (N_46842,N_46620,N_46661);
nand U46843 (N_46843,N_46676,N_46572);
xnor U46844 (N_46844,N_46567,N_46558);
or U46845 (N_46845,N_46723,N_46672);
or U46846 (N_46846,N_46651,N_46624);
nand U46847 (N_46847,N_46506,N_46571);
nor U46848 (N_46848,N_46524,N_46588);
nand U46849 (N_46849,N_46716,N_46675);
xnor U46850 (N_46850,N_46727,N_46655);
nor U46851 (N_46851,N_46608,N_46639);
nor U46852 (N_46852,N_46690,N_46668);
and U46853 (N_46853,N_46738,N_46729);
and U46854 (N_46854,N_46580,N_46549);
nor U46855 (N_46855,N_46566,N_46649);
nand U46856 (N_46856,N_46593,N_46635);
nor U46857 (N_46857,N_46547,N_46597);
or U46858 (N_46858,N_46674,N_46612);
or U46859 (N_46859,N_46648,N_46732);
and U46860 (N_46860,N_46673,N_46520);
nor U46861 (N_46861,N_46543,N_46556);
and U46862 (N_46862,N_46502,N_46565);
or U46863 (N_46863,N_46645,N_46685);
xnor U46864 (N_46864,N_46662,N_46622);
nor U46865 (N_46865,N_46626,N_46629);
or U46866 (N_46866,N_46564,N_46623);
nor U46867 (N_46867,N_46530,N_46733);
and U46868 (N_46868,N_46734,N_46714);
xor U46869 (N_46869,N_46573,N_46647);
nor U46870 (N_46870,N_46640,N_46544);
nor U46871 (N_46871,N_46537,N_46519);
or U46872 (N_46872,N_46749,N_46552);
or U46873 (N_46873,N_46590,N_46500);
nor U46874 (N_46874,N_46642,N_46741);
xnor U46875 (N_46875,N_46577,N_46737);
or U46876 (N_46876,N_46681,N_46667);
nand U46877 (N_46877,N_46583,N_46677);
xor U46878 (N_46878,N_46543,N_46724);
and U46879 (N_46879,N_46648,N_46714);
and U46880 (N_46880,N_46626,N_46712);
nand U46881 (N_46881,N_46728,N_46647);
xor U46882 (N_46882,N_46536,N_46686);
and U46883 (N_46883,N_46544,N_46547);
or U46884 (N_46884,N_46526,N_46725);
nand U46885 (N_46885,N_46622,N_46713);
nand U46886 (N_46886,N_46653,N_46729);
nand U46887 (N_46887,N_46590,N_46688);
xor U46888 (N_46888,N_46677,N_46675);
nand U46889 (N_46889,N_46706,N_46558);
nand U46890 (N_46890,N_46530,N_46500);
nor U46891 (N_46891,N_46584,N_46717);
nand U46892 (N_46892,N_46544,N_46691);
and U46893 (N_46893,N_46640,N_46510);
nand U46894 (N_46894,N_46676,N_46612);
nor U46895 (N_46895,N_46679,N_46653);
and U46896 (N_46896,N_46735,N_46727);
nand U46897 (N_46897,N_46517,N_46741);
or U46898 (N_46898,N_46675,N_46546);
nor U46899 (N_46899,N_46747,N_46501);
and U46900 (N_46900,N_46527,N_46681);
nor U46901 (N_46901,N_46574,N_46580);
nor U46902 (N_46902,N_46652,N_46574);
xor U46903 (N_46903,N_46723,N_46561);
and U46904 (N_46904,N_46701,N_46579);
nor U46905 (N_46905,N_46506,N_46592);
and U46906 (N_46906,N_46579,N_46708);
nand U46907 (N_46907,N_46593,N_46581);
nor U46908 (N_46908,N_46502,N_46698);
xnor U46909 (N_46909,N_46618,N_46667);
and U46910 (N_46910,N_46640,N_46735);
xnor U46911 (N_46911,N_46644,N_46522);
nand U46912 (N_46912,N_46593,N_46564);
nor U46913 (N_46913,N_46665,N_46709);
and U46914 (N_46914,N_46571,N_46655);
nor U46915 (N_46915,N_46690,N_46697);
nand U46916 (N_46916,N_46711,N_46720);
xnor U46917 (N_46917,N_46736,N_46717);
nand U46918 (N_46918,N_46625,N_46614);
nor U46919 (N_46919,N_46705,N_46625);
nor U46920 (N_46920,N_46626,N_46676);
or U46921 (N_46921,N_46559,N_46536);
and U46922 (N_46922,N_46661,N_46573);
or U46923 (N_46923,N_46723,N_46595);
nor U46924 (N_46924,N_46512,N_46517);
xnor U46925 (N_46925,N_46655,N_46685);
nand U46926 (N_46926,N_46743,N_46610);
nor U46927 (N_46927,N_46716,N_46709);
nor U46928 (N_46928,N_46679,N_46575);
nand U46929 (N_46929,N_46595,N_46517);
and U46930 (N_46930,N_46589,N_46538);
nor U46931 (N_46931,N_46502,N_46677);
and U46932 (N_46932,N_46665,N_46716);
and U46933 (N_46933,N_46627,N_46607);
nor U46934 (N_46934,N_46724,N_46671);
nor U46935 (N_46935,N_46715,N_46742);
nor U46936 (N_46936,N_46577,N_46667);
or U46937 (N_46937,N_46684,N_46694);
xor U46938 (N_46938,N_46579,N_46553);
nand U46939 (N_46939,N_46718,N_46634);
nor U46940 (N_46940,N_46511,N_46743);
or U46941 (N_46941,N_46679,N_46584);
xnor U46942 (N_46942,N_46699,N_46524);
xnor U46943 (N_46943,N_46598,N_46667);
and U46944 (N_46944,N_46513,N_46683);
nor U46945 (N_46945,N_46718,N_46520);
and U46946 (N_46946,N_46716,N_46728);
nand U46947 (N_46947,N_46565,N_46552);
and U46948 (N_46948,N_46559,N_46513);
or U46949 (N_46949,N_46546,N_46617);
xor U46950 (N_46950,N_46559,N_46556);
nor U46951 (N_46951,N_46597,N_46719);
nor U46952 (N_46952,N_46734,N_46562);
or U46953 (N_46953,N_46627,N_46685);
nand U46954 (N_46954,N_46631,N_46708);
and U46955 (N_46955,N_46641,N_46736);
nor U46956 (N_46956,N_46556,N_46542);
nand U46957 (N_46957,N_46550,N_46511);
nor U46958 (N_46958,N_46601,N_46551);
xor U46959 (N_46959,N_46639,N_46701);
nor U46960 (N_46960,N_46614,N_46657);
nor U46961 (N_46961,N_46696,N_46507);
or U46962 (N_46962,N_46673,N_46572);
nand U46963 (N_46963,N_46727,N_46567);
nor U46964 (N_46964,N_46600,N_46621);
xnor U46965 (N_46965,N_46558,N_46529);
and U46966 (N_46966,N_46686,N_46699);
nand U46967 (N_46967,N_46631,N_46736);
nand U46968 (N_46968,N_46535,N_46623);
nand U46969 (N_46969,N_46624,N_46563);
and U46970 (N_46970,N_46577,N_46708);
or U46971 (N_46971,N_46646,N_46533);
xor U46972 (N_46972,N_46677,N_46708);
and U46973 (N_46973,N_46645,N_46656);
or U46974 (N_46974,N_46668,N_46604);
nand U46975 (N_46975,N_46735,N_46633);
or U46976 (N_46976,N_46596,N_46578);
and U46977 (N_46977,N_46535,N_46574);
xnor U46978 (N_46978,N_46673,N_46591);
nor U46979 (N_46979,N_46629,N_46523);
xnor U46980 (N_46980,N_46590,N_46634);
xor U46981 (N_46981,N_46723,N_46615);
nor U46982 (N_46982,N_46713,N_46612);
nor U46983 (N_46983,N_46579,N_46523);
nand U46984 (N_46984,N_46696,N_46589);
or U46985 (N_46985,N_46622,N_46684);
and U46986 (N_46986,N_46547,N_46677);
nor U46987 (N_46987,N_46728,N_46542);
nand U46988 (N_46988,N_46504,N_46579);
nor U46989 (N_46989,N_46721,N_46691);
xor U46990 (N_46990,N_46658,N_46586);
or U46991 (N_46991,N_46719,N_46676);
nor U46992 (N_46992,N_46690,N_46656);
and U46993 (N_46993,N_46715,N_46516);
or U46994 (N_46994,N_46555,N_46560);
and U46995 (N_46995,N_46566,N_46666);
or U46996 (N_46996,N_46599,N_46734);
and U46997 (N_46997,N_46682,N_46501);
and U46998 (N_46998,N_46644,N_46636);
xnor U46999 (N_46999,N_46666,N_46551);
xnor U47000 (N_47000,N_46931,N_46991);
nand U47001 (N_47001,N_46944,N_46998);
and U47002 (N_47002,N_46832,N_46992);
nand U47003 (N_47003,N_46799,N_46906);
nand U47004 (N_47004,N_46864,N_46898);
nor U47005 (N_47005,N_46926,N_46943);
or U47006 (N_47006,N_46753,N_46997);
or U47007 (N_47007,N_46960,N_46867);
nand U47008 (N_47008,N_46825,N_46887);
nand U47009 (N_47009,N_46860,N_46941);
xnor U47010 (N_47010,N_46759,N_46801);
or U47011 (N_47011,N_46827,N_46904);
and U47012 (N_47012,N_46818,N_46861);
xnor U47013 (N_47013,N_46889,N_46976);
nor U47014 (N_47014,N_46972,N_46762);
nor U47015 (N_47015,N_46988,N_46975);
xnor U47016 (N_47016,N_46798,N_46752);
nor U47017 (N_47017,N_46881,N_46769);
xor U47018 (N_47018,N_46828,N_46844);
nand U47019 (N_47019,N_46968,N_46761);
or U47020 (N_47020,N_46862,N_46876);
xnor U47021 (N_47021,N_46901,N_46873);
and U47022 (N_47022,N_46900,N_46894);
or U47023 (N_47023,N_46826,N_46952);
or U47024 (N_47024,N_46806,N_46804);
or U47025 (N_47025,N_46927,N_46786);
and U47026 (N_47026,N_46956,N_46961);
xnor U47027 (N_47027,N_46866,N_46750);
nor U47028 (N_47028,N_46802,N_46882);
nor U47029 (N_47029,N_46883,N_46817);
nand U47030 (N_47030,N_46781,N_46850);
or U47031 (N_47031,N_46948,N_46830);
or U47032 (N_47032,N_46925,N_46777);
and U47033 (N_47033,N_46824,N_46831);
nor U47034 (N_47034,N_46884,N_46986);
and U47035 (N_47035,N_46839,N_46836);
or U47036 (N_47036,N_46792,N_46970);
nand U47037 (N_47037,N_46980,N_46978);
nor U47038 (N_47038,N_46751,N_46954);
or U47039 (N_47039,N_46913,N_46985);
xor U47040 (N_47040,N_46963,N_46989);
xnor U47041 (N_47041,N_46812,N_46914);
xnor U47042 (N_47042,N_46923,N_46964);
nand U47043 (N_47043,N_46758,N_46819);
nor U47044 (N_47044,N_46892,N_46754);
and U47045 (N_47045,N_46994,N_46919);
or U47046 (N_47046,N_46787,N_46955);
and U47047 (N_47047,N_46885,N_46971);
nand U47048 (N_47048,N_46767,N_46909);
and U47049 (N_47049,N_46987,N_46796);
or U47050 (N_47050,N_46805,N_46915);
xnor U47051 (N_47051,N_46911,N_46999);
or U47052 (N_47052,N_46807,N_46973);
nand U47053 (N_47053,N_46765,N_46966);
xor U47054 (N_47054,N_46924,N_46778);
and U47055 (N_47055,N_46848,N_46780);
nand U47056 (N_47056,N_46953,N_46859);
nand U47057 (N_47057,N_46764,N_46854);
or U47058 (N_47058,N_46916,N_46810);
nand U47059 (N_47059,N_46995,N_46803);
or U47060 (N_47060,N_46766,N_46789);
nand U47061 (N_47061,N_46790,N_46933);
nand U47062 (N_47062,N_46783,N_46929);
and U47063 (N_47063,N_46815,N_46895);
and U47064 (N_47064,N_46782,N_46903);
nand U47065 (N_47065,N_46846,N_46771);
nor U47066 (N_47066,N_46756,N_46930);
nand U47067 (N_47067,N_46856,N_46870);
and U47068 (N_47068,N_46833,N_46775);
or U47069 (N_47069,N_46865,N_46977);
nand U47070 (N_47070,N_46935,N_46829);
xor U47071 (N_47071,N_46993,N_46945);
nand U47072 (N_47072,N_46772,N_46852);
nor U47073 (N_47073,N_46875,N_46962);
or U47074 (N_47074,N_46811,N_46910);
nand U47075 (N_47075,N_46842,N_46957);
or U47076 (N_47076,N_46982,N_46816);
xor U47077 (N_47077,N_46845,N_46981);
and U47078 (N_47078,N_46908,N_46851);
xor U47079 (N_47079,N_46905,N_46809);
xor U47080 (N_47080,N_46763,N_46984);
xnor U47081 (N_47081,N_46857,N_46785);
nand U47082 (N_47082,N_46928,N_46879);
nand U47083 (N_47083,N_46969,N_46899);
nor U47084 (N_47084,N_46918,N_46947);
nor U47085 (N_47085,N_46990,N_46808);
and U47086 (N_47086,N_46820,N_46814);
or U47087 (N_47087,N_46821,N_46912);
nor U47088 (N_47088,N_46907,N_46784);
nand U47089 (N_47089,N_46940,N_46958);
or U47090 (N_47090,N_46967,N_46880);
xor U47091 (N_47091,N_46779,N_46788);
nor U47092 (N_47092,N_46773,N_46822);
nand U47093 (N_47093,N_46949,N_46942);
nand U47094 (N_47094,N_46946,N_46950);
xnor U47095 (N_47095,N_46872,N_46877);
or U47096 (N_47096,N_46874,N_46890);
xor U47097 (N_47097,N_46797,N_46840);
nor U47098 (N_47098,N_46791,N_46886);
nand U47099 (N_47099,N_46868,N_46849);
or U47100 (N_47100,N_46858,N_46841);
or U47101 (N_47101,N_46893,N_46863);
nor U47102 (N_47102,N_46939,N_46776);
and U47103 (N_47103,N_46834,N_46847);
nor U47104 (N_47104,N_46768,N_46871);
nand U47105 (N_47105,N_46891,N_46853);
nor U47106 (N_47106,N_46800,N_46774);
xnor U47107 (N_47107,N_46755,N_46888);
or U47108 (N_47108,N_46878,N_46770);
nand U47109 (N_47109,N_46897,N_46902);
xnor U47110 (N_47110,N_46793,N_46951);
xor U47111 (N_47111,N_46921,N_46920);
or U47112 (N_47112,N_46843,N_46959);
and U47113 (N_47113,N_46794,N_46835);
and U47114 (N_47114,N_46760,N_46938);
nor U47115 (N_47115,N_46823,N_46965);
or U47116 (N_47116,N_46974,N_46869);
and U47117 (N_47117,N_46983,N_46838);
xor U47118 (N_47118,N_46932,N_46917);
or U47119 (N_47119,N_46813,N_46934);
and U47120 (N_47120,N_46936,N_46757);
or U47121 (N_47121,N_46922,N_46795);
or U47122 (N_47122,N_46979,N_46996);
nor U47123 (N_47123,N_46896,N_46855);
nor U47124 (N_47124,N_46937,N_46837);
and U47125 (N_47125,N_46785,N_46937);
nor U47126 (N_47126,N_46831,N_46973);
or U47127 (N_47127,N_46909,N_46973);
and U47128 (N_47128,N_46910,N_46892);
and U47129 (N_47129,N_46759,N_46804);
xor U47130 (N_47130,N_46752,N_46783);
xnor U47131 (N_47131,N_46928,N_46792);
nor U47132 (N_47132,N_46977,N_46869);
nor U47133 (N_47133,N_46814,N_46757);
and U47134 (N_47134,N_46787,N_46877);
nor U47135 (N_47135,N_46951,N_46991);
nor U47136 (N_47136,N_46764,N_46949);
or U47137 (N_47137,N_46778,N_46765);
or U47138 (N_47138,N_46918,N_46807);
nor U47139 (N_47139,N_46812,N_46858);
nand U47140 (N_47140,N_46912,N_46799);
or U47141 (N_47141,N_46938,N_46866);
nand U47142 (N_47142,N_46827,N_46781);
or U47143 (N_47143,N_46758,N_46939);
and U47144 (N_47144,N_46919,N_46895);
xor U47145 (N_47145,N_46799,N_46910);
and U47146 (N_47146,N_46754,N_46959);
and U47147 (N_47147,N_46981,N_46882);
and U47148 (N_47148,N_46951,N_46880);
nand U47149 (N_47149,N_46920,N_46807);
xnor U47150 (N_47150,N_46808,N_46981);
nor U47151 (N_47151,N_46869,N_46983);
nand U47152 (N_47152,N_46894,N_46954);
nor U47153 (N_47153,N_46868,N_46800);
or U47154 (N_47154,N_46849,N_46957);
nand U47155 (N_47155,N_46891,N_46978);
and U47156 (N_47156,N_46807,N_46960);
or U47157 (N_47157,N_46831,N_46816);
nor U47158 (N_47158,N_46782,N_46917);
and U47159 (N_47159,N_46834,N_46910);
nand U47160 (N_47160,N_46847,N_46804);
nand U47161 (N_47161,N_46928,N_46833);
xnor U47162 (N_47162,N_46983,N_46789);
xor U47163 (N_47163,N_46934,N_46755);
and U47164 (N_47164,N_46789,N_46857);
nand U47165 (N_47165,N_46972,N_46756);
nor U47166 (N_47166,N_46971,N_46844);
xnor U47167 (N_47167,N_46862,N_46885);
nand U47168 (N_47168,N_46928,N_46924);
and U47169 (N_47169,N_46769,N_46961);
or U47170 (N_47170,N_46857,N_46855);
nand U47171 (N_47171,N_46818,N_46812);
or U47172 (N_47172,N_46871,N_46945);
and U47173 (N_47173,N_46827,N_46892);
nor U47174 (N_47174,N_46997,N_46881);
xnor U47175 (N_47175,N_46853,N_46826);
and U47176 (N_47176,N_46832,N_46962);
nand U47177 (N_47177,N_46998,N_46915);
nand U47178 (N_47178,N_46939,N_46971);
nand U47179 (N_47179,N_46768,N_46999);
nand U47180 (N_47180,N_46885,N_46771);
nor U47181 (N_47181,N_46840,N_46770);
nor U47182 (N_47182,N_46991,N_46822);
xnor U47183 (N_47183,N_46991,N_46753);
or U47184 (N_47184,N_46792,N_46926);
nor U47185 (N_47185,N_46864,N_46911);
xnor U47186 (N_47186,N_46870,N_46965);
or U47187 (N_47187,N_46860,N_46787);
or U47188 (N_47188,N_46963,N_46984);
xnor U47189 (N_47189,N_46901,N_46865);
nor U47190 (N_47190,N_46836,N_46900);
nand U47191 (N_47191,N_46824,N_46929);
nor U47192 (N_47192,N_46955,N_46879);
and U47193 (N_47193,N_46876,N_46810);
xor U47194 (N_47194,N_46896,N_46757);
and U47195 (N_47195,N_46807,N_46842);
or U47196 (N_47196,N_46769,N_46843);
nor U47197 (N_47197,N_46902,N_46936);
nand U47198 (N_47198,N_46998,N_46939);
xnor U47199 (N_47199,N_46834,N_46768);
xnor U47200 (N_47200,N_46855,N_46943);
or U47201 (N_47201,N_46776,N_46854);
and U47202 (N_47202,N_46793,N_46921);
xor U47203 (N_47203,N_46908,N_46999);
nor U47204 (N_47204,N_46856,N_46952);
or U47205 (N_47205,N_46957,N_46904);
nor U47206 (N_47206,N_46869,N_46857);
and U47207 (N_47207,N_46766,N_46892);
nand U47208 (N_47208,N_46915,N_46985);
or U47209 (N_47209,N_46900,N_46796);
and U47210 (N_47210,N_46838,N_46830);
or U47211 (N_47211,N_46754,N_46827);
and U47212 (N_47212,N_46870,N_46907);
nand U47213 (N_47213,N_46890,N_46838);
xnor U47214 (N_47214,N_46823,N_46899);
or U47215 (N_47215,N_46946,N_46919);
nand U47216 (N_47216,N_46960,N_46902);
or U47217 (N_47217,N_46949,N_46882);
nand U47218 (N_47218,N_46784,N_46951);
and U47219 (N_47219,N_46987,N_46908);
nor U47220 (N_47220,N_46834,N_46912);
nor U47221 (N_47221,N_46857,N_46772);
nor U47222 (N_47222,N_46871,N_46940);
xnor U47223 (N_47223,N_46834,N_46933);
or U47224 (N_47224,N_46778,N_46784);
and U47225 (N_47225,N_46971,N_46761);
nor U47226 (N_47226,N_46927,N_46928);
and U47227 (N_47227,N_46870,N_46890);
or U47228 (N_47228,N_46755,N_46778);
xnor U47229 (N_47229,N_46761,N_46861);
and U47230 (N_47230,N_46790,N_46775);
nand U47231 (N_47231,N_46942,N_46779);
and U47232 (N_47232,N_46813,N_46876);
nand U47233 (N_47233,N_46762,N_46926);
xnor U47234 (N_47234,N_46853,N_46772);
or U47235 (N_47235,N_46875,N_46953);
and U47236 (N_47236,N_46958,N_46815);
nand U47237 (N_47237,N_46820,N_46893);
and U47238 (N_47238,N_46946,N_46833);
nand U47239 (N_47239,N_46873,N_46911);
nor U47240 (N_47240,N_46836,N_46846);
xor U47241 (N_47241,N_46944,N_46975);
or U47242 (N_47242,N_46822,N_46782);
and U47243 (N_47243,N_46839,N_46797);
and U47244 (N_47244,N_46918,N_46780);
and U47245 (N_47245,N_46890,N_46982);
xnor U47246 (N_47246,N_46989,N_46898);
nand U47247 (N_47247,N_46990,N_46884);
and U47248 (N_47248,N_46953,N_46800);
nand U47249 (N_47249,N_46985,N_46858);
xnor U47250 (N_47250,N_47065,N_47058);
and U47251 (N_47251,N_47129,N_47092);
xor U47252 (N_47252,N_47206,N_47228);
nand U47253 (N_47253,N_47241,N_47214);
nand U47254 (N_47254,N_47013,N_47114);
or U47255 (N_47255,N_47128,N_47244);
or U47256 (N_47256,N_47017,N_47024);
xnor U47257 (N_47257,N_47026,N_47083);
and U47258 (N_47258,N_47201,N_47127);
or U47259 (N_47259,N_47196,N_47099);
and U47260 (N_47260,N_47219,N_47086);
and U47261 (N_47261,N_47081,N_47121);
nor U47262 (N_47262,N_47073,N_47022);
nand U47263 (N_47263,N_47234,N_47134);
xor U47264 (N_47264,N_47146,N_47240);
and U47265 (N_47265,N_47185,N_47225);
and U47266 (N_47266,N_47018,N_47015);
nor U47267 (N_47267,N_47130,N_47235);
and U47268 (N_47268,N_47115,N_47061);
nand U47269 (N_47269,N_47060,N_47047);
nand U47270 (N_47270,N_47052,N_47156);
and U47271 (N_47271,N_47221,N_47195);
or U47272 (N_47272,N_47070,N_47067);
nand U47273 (N_47273,N_47102,N_47216);
xor U47274 (N_47274,N_47220,N_47066);
xor U47275 (N_47275,N_47105,N_47120);
and U47276 (N_47276,N_47093,N_47123);
or U47277 (N_47277,N_47182,N_47176);
xor U47278 (N_47278,N_47135,N_47029);
nor U47279 (N_47279,N_47245,N_47054);
or U47280 (N_47280,N_47207,N_47124);
nor U47281 (N_47281,N_47012,N_47160);
xnor U47282 (N_47282,N_47137,N_47154);
and U47283 (N_47283,N_47224,N_47091);
nor U47284 (N_47284,N_47183,N_47243);
nand U47285 (N_47285,N_47162,N_47033);
or U47286 (N_47286,N_47143,N_47095);
nor U47287 (N_47287,N_47180,N_47164);
and U47288 (N_47288,N_47088,N_47181);
or U47289 (N_47289,N_47056,N_47075);
nand U47290 (N_47290,N_47157,N_47050);
xnor U47291 (N_47291,N_47098,N_47167);
xor U47292 (N_47292,N_47163,N_47155);
and U47293 (N_47293,N_47215,N_47064);
nor U47294 (N_47294,N_47229,N_47147);
and U47295 (N_47295,N_47204,N_47142);
and U47296 (N_47296,N_47021,N_47097);
nand U47297 (N_47297,N_47011,N_47037);
nand U47298 (N_47298,N_47209,N_47108);
xor U47299 (N_47299,N_47222,N_47144);
nand U47300 (N_47300,N_47110,N_47169);
or U47301 (N_47301,N_47051,N_47149);
nand U47302 (N_47302,N_47090,N_47186);
xnor U47303 (N_47303,N_47072,N_47117);
xor U47304 (N_47304,N_47170,N_47200);
nor U47305 (N_47305,N_47153,N_47223);
and U47306 (N_47306,N_47212,N_47084);
and U47307 (N_47307,N_47131,N_47014);
nor U47308 (N_47308,N_47236,N_47198);
and U47309 (N_47309,N_47008,N_47116);
xor U47310 (N_47310,N_47044,N_47028);
nor U47311 (N_47311,N_47139,N_47217);
nand U47312 (N_47312,N_47071,N_47035);
nor U47313 (N_47313,N_47055,N_47172);
or U47314 (N_47314,N_47249,N_47082);
nand U47315 (N_47315,N_47004,N_47173);
nand U47316 (N_47316,N_47096,N_47046);
nand U47317 (N_47317,N_47074,N_47062);
nor U47318 (N_47318,N_47208,N_47001);
or U47319 (N_47319,N_47175,N_47193);
and U47320 (N_47320,N_47166,N_47042);
nor U47321 (N_47321,N_47232,N_47152);
and U47322 (N_47322,N_47192,N_47202);
nor U47323 (N_47323,N_47184,N_47048);
nor U47324 (N_47324,N_47133,N_47161);
or U47325 (N_47325,N_47069,N_47002);
xnor U47326 (N_47326,N_47125,N_47112);
nand U47327 (N_47327,N_47199,N_47246);
nor U47328 (N_47328,N_47159,N_47104);
nor U47329 (N_47329,N_47205,N_47165);
nand U47330 (N_47330,N_47231,N_47132);
nor U47331 (N_47331,N_47039,N_47118);
or U47332 (N_47332,N_47178,N_47031);
xor U47333 (N_47333,N_47171,N_47087);
xnor U47334 (N_47334,N_47227,N_47188);
nand U47335 (N_47335,N_47187,N_47168);
nand U47336 (N_47336,N_47059,N_47247);
and U47337 (N_47337,N_47238,N_47136);
nand U47338 (N_47338,N_47106,N_47109);
and U47339 (N_47339,N_47145,N_47080);
xnor U47340 (N_47340,N_47043,N_47141);
xnor U47341 (N_47341,N_47158,N_47203);
xnor U47342 (N_47342,N_47211,N_47094);
and U47343 (N_47343,N_47041,N_47010);
xor U47344 (N_47344,N_47045,N_47113);
or U47345 (N_47345,N_47148,N_47138);
or U47346 (N_47346,N_47079,N_47076);
xnor U47347 (N_47347,N_47077,N_47101);
and U47348 (N_47348,N_47003,N_47210);
xnor U47349 (N_47349,N_47009,N_47151);
xnor U47350 (N_47350,N_47036,N_47078);
nor U47351 (N_47351,N_47213,N_47242);
or U47352 (N_47352,N_47030,N_47007);
and U47353 (N_47353,N_47177,N_47230);
and U47354 (N_47354,N_47190,N_47068);
or U47355 (N_47355,N_47107,N_47150);
and U47356 (N_47356,N_47233,N_47023);
nand U47357 (N_47357,N_47119,N_47034);
nand U47358 (N_47358,N_47085,N_47040);
xnor U47359 (N_47359,N_47197,N_47025);
or U47360 (N_47360,N_47239,N_47038);
and U47361 (N_47361,N_47140,N_47020);
and U47362 (N_47362,N_47218,N_47191);
nor U47363 (N_47363,N_47032,N_47174);
nor U47364 (N_47364,N_47053,N_47027);
xor U47365 (N_47365,N_47100,N_47111);
and U47366 (N_47366,N_47049,N_47006);
nor U47367 (N_47367,N_47019,N_47016);
and U47368 (N_47368,N_47226,N_47122);
and U47369 (N_47369,N_47237,N_47005);
or U47370 (N_47370,N_47000,N_47057);
xnor U47371 (N_47371,N_47089,N_47179);
or U47372 (N_47372,N_47063,N_47248);
nand U47373 (N_47373,N_47103,N_47189);
and U47374 (N_47374,N_47194,N_47126);
xnor U47375 (N_47375,N_47152,N_47191);
nor U47376 (N_47376,N_47042,N_47120);
or U47377 (N_47377,N_47092,N_47114);
xor U47378 (N_47378,N_47076,N_47192);
xnor U47379 (N_47379,N_47102,N_47178);
or U47380 (N_47380,N_47110,N_47221);
and U47381 (N_47381,N_47217,N_47102);
nand U47382 (N_47382,N_47175,N_47086);
and U47383 (N_47383,N_47229,N_47019);
nor U47384 (N_47384,N_47177,N_47063);
and U47385 (N_47385,N_47052,N_47016);
nand U47386 (N_47386,N_47105,N_47089);
nor U47387 (N_47387,N_47084,N_47131);
and U47388 (N_47388,N_47197,N_47153);
xnor U47389 (N_47389,N_47193,N_47037);
or U47390 (N_47390,N_47235,N_47187);
or U47391 (N_47391,N_47200,N_47009);
xnor U47392 (N_47392,N_47006,N_47005);
nand U47393 (N_47393,N_47189,N_47240);
xor U47394 (N_47394,N_47065,N_47149);
nand U47395 (N_47395,N_47055,N_47196);
nand U47396 (N_47396,N_47019,N_47221);
xor U47397 (N_47397,N_47236,N_47022);
and U47398 (N_47398,N_47208,N_47071);
nand U47399 (N_47399,N_47004,N_47206);
or U47400 (N_47400,N_47247,N_47012);
nand U47401 (N_47401,N_47013,N_47028);
and U47402 (N_47402,N_47070,N_47097);
nand U47403 (N_47403,N_47147,N_47222);
nand U47404 (N_47404,N_47157,N_47059);
nor U47405 (N_47405,N_47162,N_47186);
and U47406 (N_47406,N_47087,N_47242);
or U47407 (N_47407,N_47196,N_47131);
and U47408 (N_47408,N_47083,N_47042);
nand U47409 (N_47409,N_47180,N_47197);
nor U47410 (N_47410,N_47249,N_47044);
or U47411 (N_47411,N_47028,N_47145);
or U47412 (N_47412,N_47049,N_47112);
and U47413 (N_47413,N_47103,N_47154);
and U47414 (N_47414,N_47136,N_47184);
nor U47415 (N_47415,N_47144,N_47008);
nor U47416 (N_47416,N_47084,N_47226);
nor U47417 (N_47417,N_47177,N_47173);
nand U47418 (N_47418,N_47057,N_47215);
or U47419 (N_47419,N_47152,N_47076);
or U47420 (N_47420,N_47137,N_47194);
nor U47421 (N_47421,N_47174,N_47123);
xnor U47422 (N_47422,N_47196,N_47177);
or U47423 (N_47423,N_47221,N_47227);
nor U47424 (N_47424,N_47147,N_47173);
xor U47425 (N_47425,N_47083,N_47249);
nor U47426 (N_47426,N_47103,N_47079);
nand U47427 (N_47427,N_47061,N_47203);
xor U47428 (N_47428,N_47221,N_47040);
xor U47429 (N_47429,N_47230,N_47124);
or U47430 (N_47430,N_47012,N_47116);
or U47431 (N_47431,N_47024,N_47133);
nor U47432 (N_47432,N_47226,N_47140);
nand U47433 (N_47433,N_47177,N_47115);
nand U47434 (N_47434,N_47132,N_47030);
or U47435 (N_47435,N_47082,N_47025);
or U47436 (N_47436,N_47059,N_47184);
xnor U47437 (N_47437,N_47242,N_47088);
or U47438 (N_47438,N_47100,N_47039);
nor U47439 (N_47439,N_47204,N_47161);
xor U47440 (N_47440,N_47101,N_47089);
and U47441 (N_47441,N_47244,N_47088);
or U47442 (N_47442,N_47154,N_47121);
xnor U47443 (N_47443,N_47049,N_47217);
or U47444 (N_47444,N_47169,N_47081);
xor U47445 (N_47445,N_47096,N_47035);
and U47446 (N_47446,N_47083,N_47248);
and U47447 (N_47447,N_47028,N_47051);
xor U47448 (N_47448,N_47034,N_47237);
nor U47449 (N_47449,N_47044,N_47185);
nand U47450 (N_47450,N_47053,N_47068);
nand U47451 (N_47451,N_47147,N_47063);
xor U47452 (N_47452,N_47183,N_47188);
and U47453 (N_47453,N_47011,N_47203);
xor U47454 (N_47454,N_47053,N_47124);
xor U47455 (N_47455,N_47041,N_47118);
xor U47456 (N_47456,N_47036,N_47054);
nor U47457 (N_47457,N_47238,N_47064);
or U47458 (N_47458,N_47173,N_47183);
xnor U47459 (N_47459,N_47053,N_47206);
or U47460 (N_47460,N_47088,N_47213);
and U47461 (N_47461,N_47088,N_47164);
or U47462 (N_47462,N_47210,N_47074);
nor U47463 (N_47463,N_47001,N_47114);
nand U47464 (N_47464,N_47139,N_47111);
xnor U47465 (N_47465,N_47249,N_47014);
nor U47466 (N_47466,N_47016,N_47202);
and U47467 (N_47467,N_47241,N_47102);
xor U47468 (N_47468,N_47012,N_47131);
or U47469 (N_47469,N_47125,N_47106);
nor U47470 (N_47470,N_47031,N_47163);
or U47471 (N_47471,N_47149,N_47109);
nand U47472 (N_47472,N_47201,N_47204);
or U47473 (N_47473,N_47169,N_47014);
or U47474 (N_47474,N_47136,N_47211);
nor U47475 (N_47475,N_47104,N_47237);
nand U47476 (N_47476,N_47110,N_47008);
and U47477 (N_47477,N_47148,N_47200);
nor U47478 (N_47478,N_47152,N_47032);
or U47479 (N_47479,N_47181,N_47045);
nor U47480 (N_47480,N_47109,N_47081);
and U47481 (N_47481,N_47218,N_47058);
nor U47482 (N_47482,N_47101,N_47205);
or U47483 (N_47483,N_47132,N_47092);
and U47484 (N_47484,N_47138,N_47050);
and U47485 (N_47485,N_47082,N_47111);
and U47486 (N_47486,N_47058,N_47111);
nand U47487 (N_47487,N_47090,N_47037);
nor U47488 (N_47488,N_47094,N_47011);
nand U47489 (N_47489,N_47013,N_47154);
and U47490 (N_47490,N_47071,N_47157);
nand U47491 (N_47491,N_47089,N_47037);
xor U47492 (N_47492,N_47136,N_47230);
nor U47493 (N_47493,N_47191,N_47239);
xnor U47494 (N_47494,N_47151,N_47243);
nand U47495 (N_47495,N_47114,N_47065);
nor U47496 (N_47496,N_47011,N_47084);
nand U47497 (N_47497,N_47114,N_47218);
xnor U47498 (N_47498,N_47091,N_47041);
and U47499 (N_47499,N_47083,N_47003);
nand U47500 (N_47500,N_47365,N_47369);
xor U47501 (N_47501,N_47425,N_47328);
or U47502 (N_47502,N_47311,N_47489);
xnor U47503 (N_47503,N_47350,N_47347);
and U47504 (N_47504,N_47348,N_47441);
and U47505 (N_47505,N_47329,N_47297);
nor U47506 (N_47506,N_47454,N_47271);
nand U47507 (N_47507,N_47404,N_47382);
xor U47508 (N_47508,N_47331,N_47469);
and U47509 (N_47509,N_47364,N_47446);
xnor U47510 (N_47510,N_47448,N_47488);
or U47511 (N_47511,N_47252,N_47261);
nand U47512 (N_47512,N_47388,N_47357);
nor U47513 (N_47513,N_47372,N_47273);
xor U47514 (N_47514,N_47356,N_47353);
and U47515 (N_47515,N_47472,N_47420);
xnor U47516 (N_47516,N_47366,N_47456);
xor U47517 (N_47517,N_47301,N_47327);
and U47518 (N_47518,N_47264,N_47268);
nor U47519 (N_47519,N_47436,N_47282);
and U47520 (N_47520,N_47468,N_47312);
and U47521 (N_47521,N_47393,N_47487);
or U47522 (N_47522,N_47259,N_47387);
nor U47523 (N_47523,N_47477,N_47412);
nor U47524 (N_47524,N_47324,N_47392);
nand U47525 (N_47525,N_47292,N_47490);
nor U47526 (N_47526,N_47408,N_47385);
nor U47527 (N_47527,N_47342,N_47407);
xor U47528 (N_47528,N_47473,N_47346);
xnor U47529 (N_47529,N_47374,N_47431);
nor U47530 (N_47530,N_47482,N_47440);
nand U47531 (N_47531,N_47355,N_47479);
nand U47532 (N_47532,N_47422,N_47352);
xor U47533 (N_47533,N_47377,N_47411);
xnor U47534 (N_47534,N_47406,N_47316);
and U47535 (N_47535,N_47499,N_47483);
nor U47536 (N_47536,N_47314,N_47277);
and U47537 (N_47537,N_47401,N_47452);
or U47538 (N_47538,N_47266,N_47379);
nor U47539 (N_47539,N_47325,N_47383);
nand U47540 (N_47540,N_47305,N_47270);
xnor U47541 (N_47541,N_47275,N_47370);
and U47542 (N_47542,N_47474,N_47302);
xnor U47543 (N_47543,N_47323,N_47281);
nor U47544 (N_47544,N_47290,N_47416);
xor U47545 (N_47545,N_47481,N_47476);
and U47546 (N_47546,N_47315,N_47283);
and U47547 (N_47547,N_47304,N_47389);
nand U47548 (N_47548,N_47380,N_47345);
and U47549 (N_47549,N_47453,N_47437);
nand U47550 (N_47550,N_47445,N_47298);
xnor U47551 (N_47551,N_47410,N_47418);
xnor U47552 (N_47552,N_47378,N_47398);
and U47553 (N_47553,N_47486,N_47433);
nor U47554 (N_47554,N_47303,N_47285);
or U47555 (N_47555,N_47337,N_47368);
or U47556 (N_47556,N_47360,N_47376);
and U47557 (N_47557,N_47423,N_47361);
xnor U47558 (N_47558,N_47419,N_47460);
nor U47559 (N_47559,N_47466,N_47443);
nor U47560 (N_47560,N_47484,N_47467);
or U47561 (N_47561,N_47399,N_47397);
nor U47562 (N_47562,N_47288,N_47262);
and U47563 (N_47563,N_47319,N_47274);
or U47564 (N_47564,N_47384,N_47258);
xnor U47565 (N_47565,N_47309,N_47415);
nor U47566 (N_47566,N_47455,N_47332);
nor U47567 (N_47567,N_47338,N_47371);
nand U47568 (N_47568,N_47320,N_47354);
nand U47569 (N_47569,N_47351,N_47293);
xor U47570 (N_47570,N_47396,N_47394);
and U47571 (N_47571,N_47363,N_47451);
and U47572 (N_47572,N_47409,N_47336);
nand U47573 (N_47573,N_47253,N_47465);
nand U47574 (N_47574,N_47341,N_47291);
xor U47575 (N_47575,N_47308,N_47349);
or U47576 (N_47576,N_47478,N_47438);
nand U47577 (N_47577,N_47405,N_47429);
and U47578 (N_47578,N_47257,N_47296);
xor U47579 (N_47579,N_47334,N_47381);
or U47580 (N_47580,N_47439,N_47461);
nand U47581 (N_47581,N_47413,N_47459);
nand U47582 (N_47582,N_47287,N_47295);
xnor U47583 (N_47583,N_47432,N_47322);
xnor U47584 (N_47584,N_47496,N_47458);
and U47585 (N_47585,N_47497,N_47417);
nor U47586 (N_47586,N_47390,N_47256);
nand U47587 (N_47587,N_47391,N_47263);
nor U47588 (N_47588,N_47250,N_47491);
nand U47589 (N_47589,N_47278,N_47470);
xnor U47590 (N_47590,N_47485,N_47464);
nor U47591 (N_47591,N_47344,N_47318);
or U47592 (N_47592,N_47276,N_47462);
xnor U47593 (N_47593,N_47280,N_47480);
xor U47594 (N_47594,N_47330,N_47359);
or U47595 (N_47595,N_47463,N_47447);
nor U47596 (N_47596,N_47498,N_47317);
xnor U47597 (N_47597,N_47339,N_47414);
nor U47598 (N_47598,N_47251,N_47313);
xnor U47599 (N_47599,N_47272,N_47457);
nor U47600 (N_47600,N_47255,N_47335);
nor U47601 (N_47601,N_47400,N_47343);
xor U47602 (N_47602,N_47395,N_47435);
xor U47603 (N_47603,N_47299,N_47265);
nor U47604 (N_47604,N_47471,N_47358);
nor U47605 (N_47605,N_47279,N_47402);
xor U47606 (N_47606,N_47284,N_47427);
or U47607 (N_47607,N_47267,N_47321);
nor U47608 (N_47608,N_47289,N_47492);
xnor U47609 (N_47609,N_47430,N_47428);
xor U47610 (N_47610,N_47260,N_47449);
or U47611 (N_47611,N_47294,N_47269);
or U47612 (N_47612,N_47495,N_47444);
and U47613 (N_47613,N_47307,N_47434);
or U47614 (N_47614,N_47475,N_47310);
and U47615 (N_47615,N_47362,N_47286);
xnor U47616 (N_47616,N_47386,N_47306);
nand U47617 (N_47617,N_47421,N_47333);
xor U47618 (N_47618,N_47494,N_47375);
nor U47619 (N_47619,N_47424,N_47450);
nand U47620 (N_47620,N_47493,N_47442);
and U47621 (N_47621,N_47254,N_47373);
nand U47622 (N_47622,N_47426,N_47403);
xnor U47623 (N_47623,N_47340,N_47367);
nand U47624 (N_47624,N_47326,N_47300);
and U47625 (N_47625,N_47344,N_47353);
xnor U47626 (N_47626,N_47414,N_47279);
nor U47627 (N_47627,N_47426,N_47328);
nor U47628 (N_47628,N_47317,N_47258);
xnor U47629 (N_47629,N_47410,N_47452);
or U47630 (N_47630,N_47322,N_47381);
nor U47631 (N_47631,N_47467,N_47274);
nor U47632 (N_47632,N_47256,N_47448);
or U47633 (N_47633,N_47304,N_47427);
or U47634 (N_47634,N_47342,N_47333);
and U47635 (N_47635,N_47300,N_47264);
nor U47636 (N_47636,N_47475,N_47480);
nand U47637 (N_47637,N_47441,N_47366);
and U47638 (N_47638,N_47269,N_47439);
and U47639 (N_47639,N_47425,N_47260);
nand U47640 (N_47640,N_47270,N_47492);
or U47641 (N_47641,N_47289,N_47420);
nor U47642 (N_47642,N_47262,N_47279);
or U47643 (N_47643,N_47298,N_47433);
nand U47644 (N_47644,N_47291,N_47496);
xor U47645 (N_47645,N_47402,N_47425);
nand U47646 (N_47646,N_47251,N_47486);
nand U47647 (N_47647,N_47467,N_47453);
xnor U47648 (N_47648,N_47272,N_47348);
nand U47649 (N_47649,N_47335,N_47250);
xor U47650 (N_47650,N_47443,N_47278);
or U47651 (N_47651,N_47260,N_47418);
and U47652 (N_47652,N_47294,N_47480);
or U47653 (N_47653,N_47410,N_47282);
nor U47654 (N_47654,N_47267,N_47466);
xor U47655 (N_47655,N_47492,N_47268);
nand U47656 (N_47656,N_47331,N_47339);
nand U47657 (N_47657,N_47381,N_47299);
xor U47658 (N_47658,N_47293,N_47378);
nand U47659 (N_47659,N_47353,N_47260);
nor U47660 (N_47660,N_47466,N_47312);
or U47661 (N_47661,N_47311,N_47478);
xor U47662 (N_47662,N_47496,N_47326);
and U47663 (N_47663,N_47277,N_47278);
and U47664 (N_47664,N_47382,N_47366);
and U47665 (N_47665,N_47295,N_47402);
and U47666 (N_47666,N_47384,N_47347);
xnor U47667 (N_47667,N_47353,N_47282);
nor U47668 (N_47668,N_47397,N_47451);
or U47669 (N_47669,N_47412,N_47439);
nand U47670 (N_47670,N_47387,N_47492);
nor U47671 (N_47671,N_47352,N_47491);
xor U47672 (N_47672,N_47300,N_47488);
nor U47673 (N_47673,N_47476,N_47387);
nand U47674 (N_47674,N_47315,N_47479);
and U47675 (N_47675,N_47432,N_47339);
nand U47676 (N_47676,N_47350,N_47348);
nand U47677 (N_47677,N_47355,N_47289);
and U47678 (N_47678,N_47408,N_47456);
and U47679 (N_47679,N_47434,N_47374);
nor U47680 (N_47680,N_47329,N_47259);
xnor U47681 (N_47681,N_47471,N_47329);
nor U47682 (N_47682,N_47421,N_47471);
and U47683 (N_47683,N_47491,N_47313);
xnor U47684 (N_47684,N_47489,N_47280);
or U47685 (N_47685,N_47360,N_47474);
or U47686 (N_47686,N_47395,N_47376);
nand U47687 (N_47687,N_47414,N_47315);
nor U47688 (N_47688,N_47376,N_47407);
or U47689 (N_47689,N_47322,N_47405);
or U47690 (N_47690,N_47337,N_47449);
xnor U47691 (N_47691,N_47406,N_47388);
and U47692 (N_47692,N_47315,N_47299);
and U47693 (N_47693,N_47325,N_47398);
or U47694 (N_47694,N_47271,N_47379);
nand U47695 (N_47695,N_47290,N_47412);
or U47696 (N_47696,N_47427,N_47459);
or U47697 (N_47697,N_47349,N_47368);
or U47698 (N_47698,N_47262,N_47440);
or U47699 (N_47699,N_47474,N_47287);
or U47700 (N_47700,N_47465,N_47283);
or U47701 (N_47701,N_47412,N_47304);
xnor U47702 (N_47702,N_47449,N_47250);
and U47703 (N_47703,N_47428,N_47442);
nor U47704 (N_47704,N_47295,N_47379);
or U47705 (N_47705,N_47437,N_47359);
nor U47706 (N_47706,N_47467,N_47438);
or U47707 (N_47707,N_47484,N_47359);
and U47708 (N_47708,N_47419,N_47466);
nor U47709 (N_47709,N_47340,N_47341);
or U47710 (N_47710,N_47271,N_47309);
nor U47711 (N_47711,N_47350,N_47260);
or U47712 (N_47712,N_47381,N_47352);
xor U47713 (N_47713,N_47282,N_47408);
and U47714 (N_47714,N_47443,N_47399);
xor U47715 (N_47715,N_47322,N_47308);
or U47716 (N_47716,N_47423,N_47454);
xor U47717 (N_47717,N_47348,N_47302);
nand U47718 (N_47718,N_47405,N_47381);
and U47719 (N_47719,N_47322,N_47290);
xnor U47720 (N_47720,N_47341,N_47277);
xnor U47721 (N_47721,N_47358,N_47493);
or U47722 (N_47722,N_47332,N_47334);
xnor U47723 (N_47723,N_47411,N_47499);
nand U47724 (N_47724,N_47292,N_47274);
and U47725 (N_47725,N_47374,N_47443);
nor U47726 (N_47726,N_47350,N_47436);
and U47727 (N_47727,N_47346,N_47293);
nor U47728 (N_47728,N_47377,N_47361);
and U47729 (N_47729,N_47338,N_47434);
nand U47730 (N_47730,N_47406,N_47365);
nand U47731 (N_47731,N_47460,N_47414);
and U47732 (N_47732,N_47366,N_47264);
xor U47733 (N_47733,N_47368,N_47493);
and U47734 (N_47734,N_47441,N_47384);
or U47735 (N_47735,N_47279,N_47408);
and U47736 (N_47736,N_47427,N_47450);
and U47737 (N_47737,N_47493,N_47262);
xnor U47738 (N_47738,N_47458,N_47468);
nor U47739 (N_47739,N_47261,N_47420);
nor U47740 (N_47740,N_47256,N_47436);
xnor U47741 (N_47741,N_47340,N_47484);
and U47742 (N_47742,N_47401,N_47273);
or U47743 (N_47743,N_47372,N_47274);
xnor U47744 (N_47744,N_47280,N_47301);
nor U47745 (N_47745,N_47389,N_47377);
xnor U47746 (N_47746,N_47439,N_47415);
and U47747 (N_47747,N_47328,N_47309);
nand U47748 (N_47748,N_47286,N_47305);
nor U47749 (N_47749,N_47422,N_47390);
nand U47750 (N_47750,N_47513,N_47664);
nor U47751 (N_47751,N_47582,N_47581);
xnor U47752 (N_47752,N_47725,N_47539);
nor U47753 (N_47753,N_47536,N_47557);
and U47754 (N_47754,N_47745,N_47720);
nand U47755 (N_47755,N_47683,N_47625);
and U47756 (N_47756,N_47565,N_47737);
nand U47757 (N_47757,N_47503,N_47649);
xor U47758 (N_47758,N_47543,N_47738);
xor U47759 (N_47759,N_47545,N_47710);
and U47760 (N_47760,N_47595,N_47681);
xnor U47761 (N_47761,N_47680,N_47736);
nand U47762 (N_47762,N_47529,N_47514);
nand U47763 (N_47763,N_47668,N_47575);
nand U47764 (N_47764,N_47703,N_47641);
or U47765 (N_47765,N_47610,N_47685);
xor U47766 (N_47766,N_47615,N_47596);
nor U47767 (N_47767,N_47580,N_47597);
nand U47768 (N_47768,N_47642,N_47623);
nand U47769 (N_47769,N_47662,N_47541);
and U47770 (N_47770,N_47639,N_47712);
xor U47771 (N_47771,N_47748,N_47588);
nor U47772 (N_47772,N_47724,N_47635);
nor U47773 (N_47773,N_47520,N_47742);
and U47774 (N_47774,N_47714,N_47674);
and U47775 (N_47775,N_47741,N_47663);
xor U47776 (N_47776,N_47654,N_47537);
xnor U47777 (N_47777,N_47690,N_47743);
nor U47778 (N_47778,N_47591,N_47616);
xnor U47779 (N_47779,N_47508,N_47574);
or U47780 (N_47780,N_47657,N_47659);
nand U47781 (N_47781,N_47731,N_47687);
xor U47782 (N_47782,N_47593,N_47705);
and U47783 (N_47783,N_47728,N_47523);
and U47784 (N_47784,N_47673,N_47535);
nand U47785 (N_47785,N_47723,N_47599);
nor U47786 (N_47786,N_47698,N_47534);
nor U47787 (N_47787,N_47617,N_47620);
and U47788 (N_47788,N_47613,N_47586);
or U47789 (N_47789,N_47542,N_47671);
and U47790 (N_47790,N_47532,N_47700);
or U47791 (N_47791,N_47678,N_47717);
or U47792 (N_47792,N_47660,N_47515);
and U47793 (N_47793,N_47630,N_47695);
nand U47794 (N_47794,N_47524,N_47540);
xnor U47795 (N_47795,N_47563,N_47730);
or U47796 (N_47796,N_47682,N_47651);
and U47797 (N_47797,N_47567,N_47516);
or U47798 (N_47798,N_47606,N_47626);
and U47799 (N_47799,N_47722,N_47533);
and U47800 (N_47800,N_47587,N_47699);
nor U47801 (N_47801,N_47584,N_47622);
and U47802 (N_47802,N_47735,N_47502);
or U47803 (N_47803,N_47528,N_47732);
nor U47804 (N_47804,N_47538,N_47519);
nor U47805 (N_47805,N_47551,N_47509);
nand U47806 (N_47806,N_47733,N_47549);
and U47807 (N_47807,N_47653,N_47629);
nand U47808 (N_47808,N_47560,N_47527);
nand U47809 (N_47809,N_47518,N_47715);
or U47810 (N_47810,N_47638,N_47704);
or U47811 (N_47811,N_47600,N_47579);
xor U47812 (N_47812,N_47697,N_47573);
and U47813 (N_47813,N_47644,N_47564);
and U47814 (N_47814,N_47640,N_47611);
and U47815 (N_47815,N_47658,N_47628);
nand U47816 (N_47816,N_47507,N_47608);
or U47817 (N_47817,N_47583,N_47566);
nand U47818 (N_47818,N_47691,N_47585);
and U47819 (N_47819,N_47562,N_47603);
nand U47820 (N_47820,N_47627,N_47553);
xnor U47821 (N_47821,N_47729,N_47601);
and U47822 (N_47822,N_47633,N_47667);
nand U47823 (N_47823,N_47568,N_47605);
nor U47824 (N_47824,N_47648,N_47689);
and U47825 (N_47825,N_47709,N_47636);
nand U47826 (N_47826,N_47501,N_47531);
nand U47827 (N_47827,N_47684,N_47643);
and U47828 (N_47828,N_47677,N_47570);
or U47829 (N_47829,N_47544,N_47713);
and U47830 (N_47830,N_47604,N_47661);
xor U47831 (N_47831,N_47598,N_47572);
nand U47832 (N_47832,N_47594,N_47510);
nand U47833 (N_47833,N_47526,N_47696);
xor U47834 (N_47834,N_47569,N_47521);
nor U47835 (N_47835,N_47655,N_47708);
nand U47836 (N_47836,N_47688,N_47631);
xnor U47837 (N_47837,N_47727,N_47554);
or U47838 (N_47838,N_47686,N_47609);
nand U47839 (N_47839,N_47561,N_47550);
nand U47840 (N_47840,N_47692,N_47612);
xor U47841 (N_47841,N_47607,N_47707);
and U47842 (N_47842,N_47530,N_47749);
nand U47843 (N_47843,N_47676,N_47546);
xnor U47844 (N_47844,N_47719,N_47578);
nand U47845 (N_47845,N_47558,N_47701);
and U47846 (N_47846,N_47618,N_47512);
nor U47847 (N_47847,N_47632,N_47747);
or U47848 (N_47848,N_47669,N_47706);
nand U47849 (N_47849,N_47744,N_47506);
xor U47850 (N_47850,N_47548,N_47577);
nand U47851 (N_47851,N_47679,N_47702);
xnor U47852 (N_47852,N_47525,N_47589);
and U47853 (N_47853,N_47694,N_47672);
nand U47854 (N_47854,N_47517,N_47726);
nand U47855 (N_47855,N_47716,N_47740);
and U47856 (N_47856,N_47555,N_47652);
nor U47857 (N_47857,N_47734,N_47670);
nor U47858 (N_47858,N_47522,N_47571);
nand U47859 (N_47859,N_47637,N_47665);
xnor U47860 (N_47860,N_47621,N_47592);
nand U47861 (N_47861,N_47646,N_47746);
nand U47862 (N_47862,N_47511,N_47647);
nand U47863 (N_47863,N_47693,N_47576);
nand U47864 (N_47864,N_47602,N_47650);
or U47865 (N_47865,N_47504,N_47718);
xnor U47866 (N_47866,N_47675,N_47739);
or U47867 (N_47867,N_47634,N_47666);
or U47868 (N_47868,N_47556,N_47559);
nand U47869 (N_47869,N_47624,N_47645);
nor U47870 (N_47870,N_47721,N_47656);
or U47871 (N_47871,N_47711,N_47614);
or U47872 (N_47872,N_47505,N_47619);
nand U47873 (N_47873,N_47552,N_47590);
and U47874 (N_47874,N_47547,N_47500);
and U47875 (N_47875,N_47519,N_47530);
and U47876 (N_47876,N_47562,N_47599);
nor U47877 (N_47877,N_47506,N_47573);
or U47878 (N_47878,N_47582,N_47699);
or U47879 (N_47879,N_47657,N_47653);
nor U47880 (N_47880,N_47541,N_47681);
nor U47881 (N_47881,N_47648,N_47549);
nor U47882 (N_47882,N_47693,N_47515);
xnor U47883 (N_47883,N_47611,N_47517);
nand U47884 (N_47884,N_47516,N_47721);
nor U47885 (N_47885,N_47550,N_47607);
nand U47886 (N_47886,N_47662,N_47558);
xnor U47887 (N_47887,N_47653,N_47624);
nand U47888 (N_47888,N_47609,N_47641);
nor U47889 (N_47889,N_47680,N_47603);
xor U47890 (N_47890,N_47658,N_47513);
and U47891 (N_47891,N_47732,N_47522);
nor U47892 (N_47892,N_47723,N_47626);
nand U47893 (N_47893,N_47638,N_47662);
and U47894 (N_47894,N_47586,N_47590);
nand U47895 (N_47895,N_47507,N_47685);
xor U47896 (N_47896,N_47543,N_47677);
or U47897 (N_47897,N_47706,N_47704);
xor U47898 (N_47898,N_47741,N_47748);
nor U47899 (N_47899,N_47524,N_47567);
and U47900 (N_47900,N_47612,N_47669);
nand U47901 (N_47901,N_47504,N_47685);
and U47902 (N_47902,N_47631,N_47653);
or U47903 (N_47903,N_47711,N_47622);
or U47904 (N_47904,N_47583,N_47524);
xor U47905 (N_47905,N_47534,N_47681);
and U47906 (N_47906,N_47612,N_47561);
xnor U47907 (N_47907,N_47736,N_47667);
or U47908 (N_47908,N_47586,N_47633);
or U47909 (N_47909,N_47601,N_47634);
nand U47910 (N_47910,N_47675,N_47649);
and U47911 (N_47911,N_47682,N_47564);
xor U47912 (N_47912,N_47577,N_47588);
and U47913 (N_47913,N_47707,N_47681);
and U47914 (N_47914,N_47626,N_47684);
or U47915 (N_47915,N_47694,N_47572);
nor U47916 (N_47916,N_47550,N_47634);
nand U47917 (N_47917,N_47673,N_47687);
and U47918 (N_47918,N_47563,N_47560);
nor U47919 (N_47919,N_47509,N_47593);
nand U47920 (N_47920,N_47526,N_47707);
and U47921 (N_47921,N_47667,N_47570);
and U47922 (N_47922,N_47639,N_47715);
xor U47923 (N_47923,N_47547,N_47597);
xnor U47924 (N_47924,N_47612,N_47677);
or U47925 (N_47925,N_47677,N_47656);
xor U47926 (N_47926,N_47683,N_47524);
nand U47927 (N_47927,N_47568,N_47711);
or U47928 (N_47928,N_47663,N_47567);
nand U47929 (N_47929,N_47500,N_47682);
and U47930 (N_47930,N_47576,N_47700);
nand U47931 (N_47931,N_47744,N_47602);
xor U47932 (N_47932,N_47552,N_47743);
nor U47933 (N_47933,N_47530,N_47680);
or U47934 (N_47934,N_47713,N_47582);
and U47935 (N_47935,N_47562,N_47531);
xnor U47936 (N_47936,N_47670,N_47653);
nor U47937 (N_47937,N_47691,N_47674);
xor U47938 (N_47938,N_47526,N_47581);
xnor U47939 (N_47939,N_47698,N_47583);
nor U47940 (N_47940,N_47601,N_47614);
xor U47941 (N_47941,N_47659,N_47541);
xnor U47942 (N_47942,N_47566,N_47704);
xor U47943 (N_47943,N_47531,N_47657);
nor U47944 (N_47944,N_47578,N_47594);
nand U47945 (N_47945,N_47651,N_47702);
and U47946 (N_47946,N_47726,N_47564);
nand U47947 (N_47947,N_47655,N_47516);
and U47948 (N_47948,N_47522,N_47658);
and U47949 (N_47949,N_47510,N_47533);
nor U47950 (N_47950,N_47594,N_47714);
and U47951 (N_47951,N_47569,N_47557);
nand U47952 (N_47952,N_47544,N_47670);
or U47953 (N_47953,N_47540,N_47745);
xor U47954 (N_47954,N_47697,N_47525);
nand U47955 (N_47955,N_47590,N_47636);
nor U47956 (N_47956,N_47605,N_47727);
nand U47957 (N_47957,N_47577,N_47536);
and U47958 (N_47958,N_47725,N_47738);
nand U47959 (N_47959,N_47637,N_47642);
nor U47960 (N_47960,N_47550,N_47651);
and U47961 (N_47961,N_47550,N_47574);
nand U47962 (N_47962,N_47633,N_47552);
xor U47963 (N_47963,N_47737,N_47653);
or U47964 (N_47964,N_47702,N_47510);
nor U47965 (N_47965,N_47682,N_47570);
xnor U47966 (N_47966,N_47725,N_47694);
and U47967 (N_47967,N_47676,N_47588);
nor U47968 (N_47968,N_47660,N_47636);
xor U47969 (N_47969,N_47672,N_47659);
xor U47970 (N_47970,N_47701,N_47681);
nand U47971 (N_47971,N_47524,N_47646);
xnor U47972 (N_47972,N_47556,N_47534);
nor U47973 (N_47973,N_47533,N_47529);
nand U47974 (N_47974,N_47553,N_47628);
or U47975 (N_47975,N_47747,N_47540);
xnor U47976 (N_47976,N_47713,N_47556);
nor U47977 (N_47977,N_47641,N_47645);
and U47978 (N_47978,N_47690,N_47716);
xnor U47979 (N_47979,N_47545,N_47527);
nand U47980 (N_47980,N_47502,N_47594);
or U47981 (N_47981,N_47738,N_47539);
nor U47982 (N_47982,N_47560,N_47572);
xor U47983 (N_47983,N_47638,N_47745);
or U47984 (N_47984,N_47597,N_47653);
nand U47985 (N_47985,N_47509,N_47743);
xnor U47986 (N_47986,N_47514,N_47681);
or U47987 (N_47987,N_47725,N_47680);
xor U47988 (N_47988,N_47719,N_47596);
and U47989 (N_47989,N_47692,N_47583);
and U47990 (N_47990,N_47648,N_47511);
nor U47991 (N_47991,N_47533,N_47502);
and U47992 (N_47992,N_47650,N_47643);
and U47993 (N_47993,N_47697,N_47667);
and U47994 (N_47994,N_47609,N_47550);
xor U47995 (N_47995,N_47685,N_47522);
and U47996 (N_47996,N_47684,N_47589);
xor U47997 (N_47997,N_47653,N_47700);
or U47998 (N_47998,N_47585,N_47696);
nand U47999 (N_47999,N_47558,N_47501);
nand U48000 (N_48000,N_47850,N_47982);
nor U48001 (N_48001,N_47900,N_47827);
and U48002 (N_48002,N_47923,N_47851);
or U48003 (N_48003,N_47777,N_47810);
xor U48004 (N_48004,N_47908,N_47902);
xnor U48005 (N_48005,N_47882,N_47786);
and U48006 (N_48006,N_47779,N_47819);
nor U48007 (N_48007,N_47997,N_47890);
xnor U48008 (N_48008,N_47811,N_47757);
or U48009 (N_48009,N_47963,N_47826);
nand U48010 (N_48010,N_47948,N_47969);
and U48011 (N_48011,N_47848,N_47833);
or U48012 (N_48012,N_47776,N_47962);
or U48013 (N_48013,N_47822,N_47755);
nand U48014 (N_48014,N_47987,N_47775);
nor U48015 (N_48015,N_47961,N_47800);
nand U48016 (N_48016,N_47858,N_47891);
or U48017 (N_48017,N_47818,N_47876);
and U48018 (N_48018,N_47807,N_47985);
nand U48019 (N_48019,N_47844,N_47813);
nor U48020 (N_48020,N_47960,N_47880);
and U48021 (N_48021,N_47894,N_47917);
and U48022 (N_48022,N_47949,N_47935);
and U48023 (N_48023,N_47872,N_47915);
nor U48024 (N_48024,N_47954,N_47972);
nor U48025 (N_48025,N_47870,N_47874);
nand U48026 (N_48026,N_47825,N_47758);
or U48027 (N_48027,N_47845,N_47978);
nor U48028 (N_48028,N_47975,N_47835);
nand U48029 (N_48029,N_47864,N_47998);
or U48030 (N_48030,N_47938,N_47944);
and U48031 (N_48031,N_47836,N_47877);
nand U48032 (N_48032,N_47898,N_47946);
and U48033 (N_48033,N_47765,N_47842);
or U48034 (N_48034,N_47856,N_47892);
nor U48035 (N_48035,N_47869,N_47926);
xnor U48036 (N_48036,N_47752,N_47794);
nand U48037 (N_48037,N_47921,N_47909);
and U48038 (N_48038,N_47855,N_47919);
xor U48039 (N_48039,N_47847,N_47976);
nor U48040 (N_48040,N_47970,N_47971);
or U48041 (N_48041,N_47878,N_47996);
and U48042 (N_48042,N_47986,N_47980);
or U48043 (N_48043,N_47853,N_47871);
nor U48044 (N_48044,N_47884,N_47834);
xor U48045 (N_48045,N_47754,N_47801);
or U48046 (N_48046,N_47945,N_47958);
and U48047 (N_48047,N_47808,N_47965);
or U48048 (N_48048,N_47973,N_47771);
nor U48049 (N_48049,N_47803,N_47828);
or U48050 (N_48050,N_47812,N_47936);
or U48051 (N_48051,N_47814,N_47756);
or U48052 (N_48052,N_47941,N_47950);
or U48053 (N_48053,N_47957,N_47896);
nand U48054 (N_48054,N_47964,N_47860);
xor U48055 (N_48055,N_47838,N_47789);
nand U48056 (N_48056,N_47939,N_47913);
or U48057 (N_48057,N_47994,N_47859);
xnor U48058 (N_48058,N_47797,N_47966);
or U48059 (N_48059,N_47875,N_47899);
xor U48060 (N_48060,N_47889,N_47795);
xnor U48061 (N_48061,N_47861,N_47903);
xor U48062 (N_48062,N_47831,N_47798);
or U48063 (N_48063,N_47927,N_47925);
and U48064 (N_48064,N_47815,N_47796);
nand U48065 (N_48065,N_47984,N_47937);
nand U48066 (N_48066,N_47773,N_47840);
and U48067 (N_48067,N_47767,N_47955);
nand U48068 (N_48068,N_47829,N_47967);
nor U48069 (N_48069,N_47762,N_47791);
and U48070 (N_48070,N_47940,N_47934);
nor U48071 (N_48071,N_47866,N_47911);
nand U48072 (N_48072,N_47839,N_47920);
xnor U48073 (N_48073,N_47929,N_47989);
or U48074 (N_48074,N_47916,N_47922);
xor U48075 (N_48075,N_47816,N_47809);
and U48076 (N_48076,N_47897,N_47932);
nor U48077 (N_48077,N_47905,N_47865);
nand U48078 (N_48078,N_47784,N_47999);
or U48079 (N_48079,N_47783,N_47846);
or U48080 (N_48080,N_47781,N_47832);
or U48081 (N_48081,N_47914,N_47959);
xor U48082 (N_48082,N_47830,N_47764);
nand U48083 (N_48083,N_47766,N_47887);
nor U48084 (N_48084,N_47857,N_47931);
and U48085 (N_48085,N_47821,N_47912);
nor U48086 (N_48086,N_47981,N_47792);
xnor U48087 (N_48087,N_47823,N_47806);
nand U48088 (N_48088,N_47885,N_47886);
nor U48089 (N_48089,N_47895,N_47761);
xnor U48090 (N_48090,N_47873,N_47750);
nor U48091 (N_48091,N_47763,N_47849);
or U48092 (N_48092,N_47820,N_47802);
xor U48093 (N_48093,N_47804,N_47780);
nand U48094 (N_48094,N_47817,N_47953);
or U48095 (N_48095,N_47930,N_47843);
or U48096 (N_48096,N_47760,N_47863);
nand U48097 (N_48097,N_47770,N_47988);
and U48098 (N_48098,N_47906,N_47888);
nor U48099 (N_48099,N_47990,N_47837);
and U48100 (N_48100,N_47983,N_47942);
or U48101 (N_48101,N_47933,N_47951);
nand U48102 (N_48102,N_47862,N_47907);
nand U48103 (N_48103,N_47774,N_47918);
nand U48104 (N_48104,N_47824,N_47993);
nor U48105 (N_48105,N_47883,N_47879);
nand U48106 (N_48106,N_47977,N_47904);
nand U48107 (N_48107,N_47753,N_47893);
nand U48108 (N_48108,N_47782,N_47805);
nand U48109 (N_48109,N_47790,N_47854);
nor U48110 (N_48110,N_47841,N_47868);
nand U48111 (N_48111,N_47901,N_47772);
and U48112 (N_48112,N_47956,N_47924);
nand U48113 (N_48113,N_47979,N_47974);
nor U48114 (N_48114,N_47968,N_47881);
and U48115 (N_48115,N_47769,N_47785);
nor U48116 (N_48116,N_47852,N_47867);
and U48117 (N_48117,N_47751,N_47778);
or U48118 (N_48118,N_47991,N_47947);
or U48119 (N_48119,N_47995,N_47788);
or U48120 (N_48120,N_47768,N_47787);
nand U48121 (N_48121,N_47928,N_47952);
nor U48122 (N_48122,N_47943,N_47759);
or U48123 (N_48123,N_47910,N_47799);
xor U48124 (N_48124,N_47992,N_47793);
xnor U48125 (N_48125,N_47828,N_47843);
nor U48126 (N_48126,N_47999,N_47906);
nor U48127 (N_48127,N_47876,N_47995);
xor U48128 (N_48128,N_47959,N_47772);
nand U48129 (N_48129,N_47984,N_47852);
and U48130 (N_48130,N_47755,N_47887);
and U48131 (N_48131,N_47903,N_47841);
nand U48132 (N_48132,N_47793,N_47966);
nand U48133 (N_48133,N_47966,N_47755);
or U48134 (N_48134,N_47859,N_47971);
and U48135 (N_48135,N_47766,N_47952);
and U48136 (N_48136,N_47754,N_47874);
nand U48137 (N_48137,N_47986,N_47785);
and U48138 (N_48138,N_47985,N_47852);
nor U48139 (N_48139,N_47904,N_47925);
and U48140 (N_48140,N_47859,N_47781);
nor U48141 (N_48141,N_47806,N_47782);
and U48142 (N_48142,N_47785,N_47938);
nor U48143 (N_48143,N_47822,N_47989);
xnor U48144 (N_48144,N_47823,N_47928);
or U48145 (N_48145,N_47831,N_47895);
nor U48146 (N_48146,N_47911,N_47906);
or U48147 (N_48147,N_47991,N_47966);
and U48148 (N_48148,N_47850,N_47936);
nand U48149 (N_48149,N_47811,N_47936);
nor U48150 (N_48150,N_47956,N_47851);
or U48151 (N_48151,N_47855,N_47938);
xor U48152 (N_48152,N_47811,N_47820);
xnor U48153 (N_48153,N_47975,N_47767);
or U48154 (N_48154,N_47898,N_47768);
nor U48155 (N_48155,N_47791,N_47892);
or U48156 (N_48156,N_47881,N_47757);
and U48157 (N_48157,N_47868,N_47768);
nor U48158 (N_48158,N_47956,N_47878);
or U48159 (N_48159,N_47825,N_47876);
and U48160 (N_48160,N_47797,N_47894);
nor U48161 (N_48161,N_47954,N_47851);
nand U48162 (N_48162,N_47752,N_47991);
and U48163 (N_48163,N_47997,N_47847);
nand U48164 (N_48164,N_47878,N_47767);
xor U48165 (N_48165,N_47838,N_47909);
xnor U48166 (N_48166,N_47993,N_47857);
xnor U48167 (N_48167,N_47800,N_47984);
nor U48168 (N_48168,N_47754,N_47907);
or U48169 (N_48169,N_47982,N_47880);
xor U48170 (N_48170,N_47901,N_47790);
nor U48171 (N_48171,N_47967,N_47785);
nor U48172 (N_48172,N_47908,N_47759);
xnor U48173 (N_48173,N_47787,N_47767);
xnor U48174 (N_48174,N_47865,N_47959);
nor U48175 (N_48175,N_47919,N_47869);
and U48176 (N_48176,N_47961,N_47988);
xor U48177 (N_48177,N_47905,N_47875);
nor U48178 (N_48178,N_47842,N_47975);
nor U48179 (N_48179,N_47996,N_47902);
or U48180 (N_48180,N_47964,N_47880);
and U48181 (N_48181,N_47787,N_47806);
xnor U48182 (N_48182,N_47961,N_47813);
nor U48183 (N_48183,N_47932,N_47948);
or U48184 (N_48184,N_47832,N_47907);
xnor U48185 (N_48185,N_47877,N_47895);
nor U48186 (N_48186,N_47954,N_47907);
and U48187 (N_48187,N_47821,N_47871);
and U48188 (N_48188,N_47829,N_47950);
and U48189 (N_48189,N_47806,N_47940);
nand U48190 (N_48190,N_47814,N_47938);
or U48191 (N_48191,N_47977,N_47924);
or U48192 (N_48192,N_47814,N_47790);
and U48193 (N_48193,N_47886,N_47866);
nand U48194 (N_48194,N_47911,N_47936);
nand U48195 (N_48195,N_47996,N_47889);
or U48196 (N_48196,N_47825,N_47871);
xor U48197 (N_48197,N_47870,N_47967);
xor U48198 (N_48198,N_47936,N_47758);
nor U48199 (N_48199,N_47801,N_47871);
nand U48200 (N_48200,N_47856,N_47759);
or U48201 (N_48201,N_47889,N_47832);
or U48202 (N_48202,N_47838,N_47875);
xnor U48203 (N_48203,N_47837,N_47864);
or U48204 (N_48204,N_47878,N_47934);
and U48205 (N_48205,N_47773,N_47994);
xor U48206 (N_48206,N_47800,N_47790);
or U48207 (N_48207,N_47777,N_47806);
and U48208 (N_48208,N_47751,N_47942);
nor U48209 (N_48209,N_47807,N_47757);
or U48210 (N_48210,N_47916,N_47931);
nand U48211 (N_48211,N_47790,N_47972);
or U48212 (N_48212,N_47862,N_47802);
xnor U48213 (N_48213,N_47941,N_47979);
xnor U48214 (N_48214,N_47837,N_47931);
xnor U48215 (N_48215,N_47825,N_47896);
nand U48216 (N_48216,N_47953,N_47766);
xor U48217 (N_48217,N_47897,N_47970);
xor U48218 (N_48218,N_47764,N_47993);
nor U48219 (N_48219,N_47983,N_47827);
nand U48220 (N_48220,N_47756,N_47984);
nand U48221 (N_48221,N_47898,N_47982);
or U48222 (N_48222,N_47881,N_47984);
nand U48223 (N_48223,N_47768,N_47847);
nor U48224 (N_48224,N_47880,N_47966);
or U48225 (N_48225,N_47911,N_47903);
nor U48226 (N_48226,N_47996,N_47919);
nor U48227 (N_48227,N_47868,N_47878);
nand U48228 (N_48228,N_47915,N_47924);
xnor U48229 (N_48229,N_47963,N_47943);
and U48230 (N_48230,N_47875,N_47776);
and U48231 (N_48231,N_47999,N_47792);
xor U48232 (N_48232,N_47877,N_47825);
nand U48233 (N_48233,N_47818,N_47877);
xnor U48234 (N_48234,N_47946,N_47883);
nor U48235 (N_48235,N_47989,N_47955);
nand U48236 (N_48236,N_47857,N_47784);
and U48237 (N_48237,N_47956,N_47773);
or U48238 (N_48238,N_47764,N_47803);
and U48239 (N_48239,N_47987,N_47794);
or U48240 (N_48240,N_47890,N_47770);
xnor U48241 (N_48241,N_47918,N_47961);
and U48242 (N_48242,N_47937,N_47814);
nand U48243 (N_48243,N_47959,N_47800);
or U48244 (N_48244,N_47979,N_47901);
nor U48245 (N_48245,N_47857,N_47894);
and U48246 (N_48246,N_47980,N_47906);
nor U48247 (N_48247,N_47917,N_47786);
nand U48248 (N_48248,N_47753,N_47866);
nand U48249 (N_48249,N_47928,N_47842);
and U48250 (N_48250,N_48185,N_48124);
and U48251 (N_48251,N_48173,N_48143);
or U48252 (N_48252,N_48190,N_48202);
and U48253 (N_48253,N_48218,N_48150);
xnor U48254 (N_48254,N_48201,N_48176);
xor U48255 (N_48255,N_48157,N_48015);
or U48256 (N_48256,N_48147,N_48014);
nor U48257 (N_48257,N_48221,N_48138);
nand U48258 (N_48258,N_48042,N_48188);
nand U48259 (N_48259,N_48197,N_48023);
and U48260 (N_48260,N_48030,N_48179);
xor U48261 (N_48261,N_48227,N_48037);
nand U48262 (N_48262,N_48132,N_48080);
nand U48263 (N_48263,N_48210,N_48046);
xor U48264 (N_48264,N_48054,N_48027);
xor U48265 (N_48265,N_48038,N_48245);
xor U48266 (N_48266,N_48158,N_48119);
xnor U48267 (N_48267,N_48220,N_48019);
nor U48268 (N_48268,N_48191,N_48065);
nand U48269 (N_48269,N_48164,N_48223);
nand U48270 (N_48270,N_48022,N_48211);
nor U48271 (N_48271,N_48112,N_48161);
or U48272 (N_48272,N_48109,N_48171);
or U48273 (N_48273,N_48060,N_48039);
nor U48274 (N_48274,N_48144,N_48021);
and U48275 (N_48275,N_48076,N_48183);
and U48276 (N_48276,N_48230,N_48208);
nand U48277 (N_48277,N_48247,N_48070);
nand U48278 (N_48278,N_48181,N_48036);
and U48279 (N_48279,N_48074,N_48149);
or U48280 (N_48280,N_48097,N_48226);
xnor U48281 (N_48281,N_48140,N_48093);
and U48282 (N_48282,N_48040,N_48103);
nand U48283 (N_48283,N_48186,N_48126);
xnor U48284 (N_48284,N_48017,N_48152);
nand U48285 (N_48285,N_48053,N_48031);
nor U48286 (N_48286,N_48088,N_48068);
xnor U48287 (N_48287,N_48059,N_48163);
or U48288 (N_48288,N_48013,N_48091);
and U48289 (N_48289,N_48101,N_48090);
or U48290 (N_48290,N_48162,N_48155);
nor U48291 (N_48291,N_48196,N_48198);
or U48292 (N_48292,N_48209,N_48003);
nor U48293 (N_48293,N_48034,N_48011);
xnor U48294 (N_48294,N_48099,N_48078);
and U48295 (N_48295,N_48082,N_48075);
xor U48296 (N_48296,N_48224,N_48026);
xor U48297 (N_48297,N_48032,N_48113);
xnor U48298 (N_48298,N_48248,N_48241);
or U48299 (N_48299,N_48096,N_48166);
or U48300 (N_48300,N_48007,N_48085);
nor U48301 (N_48301,N_48045,N_48100);
xor U48302 (N_48302,N_48115,N_48073);
nor U48303 (N_48303,N_48170,N_48243);
xnor U48304 (N_48304,N_48172,N_48184);
or U48305 (N_48305,N_48246,N_48236);
nor U48306 (N_48306,N_48005,N_48052);
nand U48307 (N_48307,N_48094,N_48130);
xnor U48308 (N_48308,N_48135,N_48192);
or U48309 (N_48309,N_48215,N_48200);
or U48310 (N_48310,N_48089,N_48071);
nand U48311 (N_48311,N_48129,N_48092);
or U48312 (N_48312,N_48086,N_48239);
nor U48313 (N_48313,N_48237,N_48047);
or U48314 (N_48314,N_48033,N_48043);
xnor U48315 (N_48315,N_48238,N_48206);
xnor U48316 (N_48316,N_48063,N_48216);
or U48317 (N_48317,N_48105,N_48156);
nor U48318 (N_48318,N_48139,N_48009);
and U48319 (N_48319,N_48087,N_48159);
xor U48320 (N_48320,N_48167,N_48120);
nor U48321 (N_48321,N_48213,N_48145);
and U48322 (N_48322,N_48182,N_48029);
nand U48323 (N_48323,N_48204,N_48012);
xor U48324 (N_48324,N_48057,N_48232);
or U48325 (N_48325,N_48116,N_48064);
and U48326 (N_48326,N_48235,N_48069);
or U48327 (N_48327,N_48205,N_48175);
nor U48328 (N_48328,N_48217,N_48229);
and U48329 (N_48329,N_48010,N_48195);
or U48330 (N_48330,N_48234,N_48044);
and U48331 (N_48331,N_48104,N_48077);
xor U48332 (N_48332,N_48207,N_48233);
and U48333 (N_48333,N_48123,N_48110);
and U48334 (N_48334,N_48121,N_48169);
and U48335 (N_48335,N_48194,N_48131);
nand U48336 (N_48336,N_48187,N_48189);
nor U48337 (N_48337,N_48006,N_48051);
xnor U48338 (N_48338,N_48151,N_48081);
nand U48339 (N_48339,N_48098,N_48244);
and U48340 (N_48340,N_48160,N_48056);
nand U48341 (N_48341,N_48242,N_48127);
nand U48342 (N_48342,N_48102,N_48168);
xnor U48343 (N_48343,N_48136,N_48153);
xor U48344 (N_48344,N_48066,N_48001);
nor U48345 (N_48345,N_48178,N_48174);
nor U48346 (N_48346,N_48106,N_48035);
or U48347 (N_48347,N_48020,N_48025);
nand U48348 (N_48348,N_48016,N_48203);
or U48349 (N_48349,N_48212,N_48154);
nor U48350 (N_48350,N_48117,N_48024);
and U48351 (N_48351,N_48004,N_48118);
or U48352 (N_48352,N_48048,N_48122);
and U48353 (N_48353,N_48240,N_48146);
nor U48354 (N_48354,N_48002,N_48084);
and U48355 (N_48355,N_48079,N_48041);
and U48356 (N_48356,N_48049,N_48177);
nor U48357 (N_48357,N_48219,N_48008);
nor U48358 (N_48358,N_48133,N_48141);
nand U48359 (N_48359,N_48067,N_48125);
xor U48360 (N_48360,N_48199,N_48083);
xnor U48361 (N_48361,N_48062,N_48108);
xnor U48362 (N_48362,N_48050,N_48228);
nor U48363 (N_48363,N_48028,N_48018);
xnor U48364 (N_48364,N_48214,N_48134);
nor U48365 (N_48365,N_48142,N_48111);
xor U48366 (N_48366,N_48148,N_48165);
nand U48367 (N_48367,N_48107,N_48225);
nor U48368 (N_48368,N_48249,N_48055);
xor U48369 (N_48369,N_48000,N_48061);
xnor U48370 (N_48370,N_48222,N_48058);
and U48371 (N_48371,N_48114,N_48180);
and U48372 (N_48372,N_48072,N_48231);
and U48373 (N_48373,N_48137,N_48095);
xor U48374 (N_48374,N_48193,N_48128);
nand U48375 (N_48375,N_48185,N_48036);
nor U48376 (N_48376,N_48191,N_48109);
xor U48377 (N_48377,N_48022,N_48073);
and U48378 (N_48378,N_48236,N_48071);
and U48379 (N_48379,N_48025,N_48070);
nand U48380 (N_48380,N_48163,N_48138);
or U48381 (N_48381,N_48037,N_48247);
nor U48382 (N_48382,N_48028,N_48122);
or U48383 (N_48383,N_48145,N_48159);
nor U48384 (N_48384,N_48110,N_48068);
and U48385 (N_48385,N_48162,N_48142);
and U48386 (N_48386,N_48044,N_48161);
nand U48387 (N_48387,N_48079,N_48074);
nand U48388 (N_48388,N_48030,N_48227);
and U48389 (N_48389,N_48081,N_48238);
or U48390 (N_48390,N_48192,N_48058);
nand U48391 (N_48391,N_48208,N_48022);
or U48392 (N_48392,N_48219,N_48222);
xor U48393 (N_48393,N_48081,N_48164);
nor U48394 (N_48394,N_48071,N_48128);
nand U48395 (N_48395,N_48139,N_48006);
and U48396 (N_48396,N_48145,N_48033);
nand U48397 (N_48397,N_48103,N_48039);
and U48398 (N_48398,N_48076,N_48164);
nand U48399 (N_48399,N_48087,N_48106);
nor U48400 (N_48400,N_48029,N_48236);
xor U48401 (N_48401,N_48136,N_48043);
nand U48402 (N_48402,N_48103,N_48010);
or U48403 (N_48403,N_48115,N_48068);
nand U48404 (N_48404,N_48174,N_48245);
nor U48405 (N_48405,N_48207,N_48156);
xor U48406 (N_48406,N_48073,N_48075);
and U48407 (N_48407,N_48088,N_48097);
and U48408 (N_48408,N_48183,N_48130);
nor U48409 (N_48409,N_48011,N_48185);
nor U48410 (N_48410,N_48105,N_48029);
nand U48411 (N_48411,N_48094,N_48198);
or U48412 (N_48412,N_48169,N_48197);
or U48413 (N_48413,N_48076,N_48069);
nand U48414 (N_48414,N_48026,N_48165);
nor U48415 (N_48415,N_48053,N_48021);
and U48416 (N_48416,N_48243,N_48238);
xor U48417 (N_48417,N_48047,N_48165);
or U48418 (N_48418,N_48090,N_48149);
and U48419 (N_48419,N_48028,N_48204);
or U48420 (N_48420,N_48067,N_48173);
or U48421 (N_48421,N_48091,N_48011);
and U48422 (N_48422,N_48236,N_48040);
or U48423 (N_48423,N_48128,N_48100);
nor U48424 (N_48424,N_48081,N_48195);
xnor U48425 (N_48425,N_48218,N_48024);
nor U48426 (N_48426,N_48038,N_48237);
or U48427 (N_48427,N_48081,N_48249);
nor U48428 (N_48428,N_48118,N_48047);
and U48429 (N_48429,N_48096,N_48043);
nand U48430 (N_48430,N_48186,N_48168);
and U48431 (N_48431,N_48059,N_48085);
and U48432 (N_48432,N_48036,N_48016);
nand U48433 (N_48433,N_48188,N_48204);
xor U48434 (N_48434,N_48026,N_48225);
nand U48435 (N_48435,N_48078,N_48069);
or U48436 (N_48436,N_48204,N_48159);
nor U48437 (N_48437,N_48217,N_48204);
nand U48438 (N_48438,N_48201,N_48058);
and U48439 (N_48439,N_48034,N_48227);
xnor U48440 (N_48440,N_48156,N_48211);
nor U48441 (N_48441,N_48167,N_48111);
or U48442 (N_48442,N_48124,N_48095);
and U48443 (N_48443,N_48214,N_48231);
xor U48444 (N_48444,N_48105,N_48019);
xor U48445 (N_48445,N_48106,N_48135);
and U48446 (N_48446,N_48109,N_48137);
nor U48447 (N_48447,N_48017,N_48024);
nand U48448 (N_48448,N_48034,N_48186);
nand U48449 (N_48449,N_48031,N_48163);
and U48450 (N_48450,N_48031,N_48152);
nand U48451 (N_48451,N_48105,N_48202);
or U48452 (N_48452,N_48109,N_48110);
nand U48453 (N_48453,N_48006,N_48212);
xnor U48454 (N_48454,N_48058,N_48050);
nor U48455 (N_48455,N_48163,N_48029);
or U48456 (N_48456,N_48100,N_48106);
and U48457 (N_48457,N_48035,N_48034);
xor U48458 (N_48458,N_48024,N_48210);
or U48459 (N_48459,N_48203,N_48173);
and U48460 (N_48460,N_48053,N_48178);
nand U48461 (N_48461,N_48091,N_48063);
nor U48462 (N_48462,N_48042,N_48121);
and U48463 (N_48463,N_48236,N_48162);
nand U48464 (N_48464,N_48198,N_48029);
nor U48465 (N_48465,N_48245,N_48102);
and U48466 (N_48466,N_48201,N_48222);
nand U48467 (N_48467,N_48223,N_48066);
nor U48468 (N_48468,N_48004,N_48032);
nor U48469 (N_48469,N_48215,N_48203);
nor U48470 (N_48470,N_48022,N_48043);
xor U48471 (N_48471,N_48239,N_48170);
nand U48472 (N_48472,N_48153,N_48043);
or U48473 (N_48473,N_48076,N_48096);
nor U48474 (N_48474,N_48222,N_48033);
nor U48475 (N_48475,N_48158,N_48097);
or U48476 (N_48476,N_48026,N_48136);
and U48477 (N_48477,N_48083,N_48039);
nand U48478 (N_48478,N_48087,N_48248);
or U48479 (N_48479,N_48150,N_48106);
xor U48480 (N_48480,N_48084,N_48112);
nor U48481 (N_48481,N_48161,N_48248);
nor U48482 (N_48482,N_48006,N_48142);
and U48483 (N_48483,N_48099,N_48001);
and U48484 (N_48484,N_48218,N_48191);
xor U48485 (N_48485,N_48013,N_48028);
and U48486 (N_48486,N_48091,N_48140);
nor U48487 (N_48487,N_48039,N_48220);
and U48488 (N_48488,N_48230,N_48084);
nor U48489 (N_48489,N_48217,N_48009);
or U48490 (N_48490,N_48187,N_48006);
or U48491 (N_48491,N_48102,N_48114);
nor U48492 (N_48492,N_48033,N_48185);
and U48493 (N_48493,N_48076,N_48192);
xnor U48494 (N_48494,N_48136,N_48116);
nor U48495 (N_48495,N_48180,N_48153);
and U48496 (N_48496,N_48062,N_48084);
xor U48497 (N_48497,N_48136,N_48046);
and U48498 (N_48498,N_48164,N_48113);
xor U48499 (N_48499,N_48159,N_48240);
or U48500 (N_48500,N_48348,N_48396);
nand U48501 (N_48501,N_48483,N_48398);
nand U48502 (N_48502,N_48364,N_48319);
nand U48503 (N_48503,N_48495,N_48453);
and U48504 (N_48504,N_48429,N_48419);
nor U48505 (N_48505,N_48260,N_48383);
nor U48506 (N_48506,N_48257,N_48271);
nor U48507 (N_48507,N_48379,N_48387);
xor U48508 (N_48508,N_48321,N_48415);
and U48509 (N_48509,N_48275,N_48488);
or U48510 (N_48510,N_48404,N_48489);
and U48511 (N_48511,N_48427,N_48468);
nor U48512 (N_48512,N_48354,N_48268);
xor U48513 (N_48513,N_48329,N_48372);
or U48514 (N_48514,N_48279,N_48420);
or U48515 (N_48515,N_48343,N_48401);
and U48516 (N_48516,N_48425,N_48418);
nand U48517 (N_48517,N_48378,N_48400);
or U48518 (N_48518,N_48498,N_48262);
or U48519 (N_48519,N_48444,N_48433);
xor U48520 (N_48520,N_48497,N_48263);
or U48521 (N_48521,N_48403,N_48309);
xor U48522 (N_48522,N_48291,N_48426);
nor U48523 (N_48523,N_48471,N_48421);
and U48524 (N_48524,N_48395,N_48469);
or U48525 (N_48525,N_48315,N_48431);
or U48526 (N_48526,N_48454,N_48411);
and U48527 (N_48527,N_48377,N_48296);
nand U48528 (N_48528,N_48351,N_48349);
xnor U48529 (N_48529,N_48325,N_48347);
or U48530 (N_48530,N_48439,N_48371);
or U48531 (N_48531,N_48294,N_48276);
xnor U48532 (N_48532,N_48350,N_48290);
xor U48533 (N_48533,N_48310,N_48408);
nor U48534 (N_48534,N_48393,N_48442);
nand U48535 (N_48535,N_48437,N_48467);
or U48536 (N_48536,N_48269,N_48438);
or U48537 (N_48537,N_48301,N_48388);
nand U48538 (N_48538,N_48424,N_48412);
or U48539 (N_48539,N_48445,N_48284);
and U48540 (N_48540,N_48264,N_48463);
nand U48541 (N_48541,N_48289,N_48340);
nor U48542 (N_48542,N_48405,N_48344);
nor U48543 (N_48543,N_48288,N_48386);
nor U48544 (N_48544,N_48283,N_48322);
xor U48545 (N_48545,N_48417,N_48481);
nor U48546 (N_48546,N_48374,N_48479);
nor U48547 (N_48547,N_48434,N_48443);
nand U48548 (N_48548,N_48470,N_48375);
nor U48549 (N_48549,N_48464,N_48258);
or U48550 (N_48550,N_48490,N_48259);
nand U48551 (N_48551,N_48255,N_48370);
xor U48552 (N_48552,N_48475,N_48451);
xnor U48553 (N_48553,N_48380,N_48413);
nor U48554 (N_48554,N_48330,N_48256);
nor U48555 (N_48555,N_48450,N_48435);
or U48556 (N_48556,N_48474,N_48494);
or U48557 (N_48557,N_48298,N_48353);
nand U48558 (N_48558,N_48428,N_48307);
xor U48559 (N_48559,N_48391,N_48492);
and U48560 (N_48560,N_48305,N_48456);
xor U48561 (N_48561,N_48368,N_48423);
or U48562 (N_48562,N_48478,N_48384);
or U48563 (N_48563,N_48300,N_48441);
nand U48564 (N_48564,N_48267,N_48251);
nand U48565 (N_48565,N_48473,N_48360);
or U48566 (N_48566,N_48422,N_48369);
or U48567 (N_48567,N_48448,N_48452);
or U48568 (N_48568,N_48480,N_48274);
nor U48569 (N_48569,N_48366,N_48327);
and U48570 (N_48570,N_48270,N_48496);
xor U48571 (N_48571,N_48282,N_48252);
and U48572 (N_48572,N_48436,N_48280);
nor U48573 (N_48573,N_48373,N_48339);
nor U48574 (N_48574,N_48345,N_48332);
nor U48575 (N_48575,N_48485,N_48416);
nand U48576 (N_48576,N_48272,N_48286);
and U48577 (N_48577,N_48407,N_48499);
nor U48578 (N_48578,N_48397,N_48334);
or U48579 (N_48579,N_48361,N_48446);
nor U48580 (N_48580,N_48362,N_48303);
xnor U48581 (N_48581,N_48317,N_48261);
nand U48582 (N_48582,N_48466,N_48293);
and U48583 (N_48583,N_48462,N_48491);
nand U48584 (N_48584,N_48394,N_48487);
xnor U48585 (N_48585,N_48352,N_48278);
nor U48586 (N_48586,N_48363,N_48472);
or U48587 (N_48587,N_48316,N_48356);
nor U48588 (N_48588,N_48265,N_48461);
nand U48589 (N_48589,N_48311,N_48449);
or U48590 (N_48590,N_48342,N_48392);
nand U48591 (N_48591,N_48493,N_48365);
or U48592 (N_48592,N_48459,N_48254);
nor U48593 (N_48593,N_48381,N_48318);
or U48594 (N_48594,N_48359,N_48324);
nor U48595 (N_48595,N_48314,N_48266);
and U48596 (N_48596,N_48402,N_48409);
nor U48597 (N_48597,N_48367,N_48304);
nand U48598 (N_48598,N_48328,N_48432);
xor U48599 (N_48599,N_48484,N_48250);
nand U48600 (N_48600,N_48482,N_48390);
nor U48601 (N_48601,N_48306,N_48292);
nand U48602 (N_48602,N_48335,N_48458);
or U48603 (N_48603,N_48302,N_48430);
nor U48604 (N_48604,N_48287,N_48410);
nand U48605 (N_48605,N_48447,N_48465);
nor U48606 (N_48606,N_48337,N_48358);
nor U48607 (N_48607,N_48326,N_48320);
nand U48608 (N_48608,N_48336,N_48457);
nor U48609 (N_48609,N_48357,N_48273);
nand U48610 (N_48610,N_48346,N_48295);
nand U48611 (N_48611,N_48440,N_48376);
nand U48612 (N_48612,N_48382,N_48399);
or U48613 (N_48613,N_48313,N_48253);
or U48614 (N_48614,N_48385,N_48299);
nor U48615 (N_48615,N_48323,N_48476);
nand U48616 (N_48616,N_48460,N_48341);
nor U48617 (N_48617,N_48355,N_48277);
and U48618 (N_48618,N_48297,N_48455);
and U48619 (N_48619,N_48406,N_48285);
xor U48620 (N_48620,N_48281,N_48477);
nand U48621 (N_48621,N_48389,N_48308);
or U48622 (N_48622,N_48331,N_48312);
or U48623 (N_48623,N_48486,N_48333);
nand U48624 (N_48624,N_48414,N_48338);
and U48625 (N_48625,N_48371,N_48352);
or U48626 (N_48626,N_48439,N_48423);
xnor U48627 (N_48627,N_48329,N_48257);
nand U48628 (N_48628,N_48459,N_48433);
nor U48629 (N_48629,N_48309,N_48369);
nor U48630 (N_48630,N_48305,N_48272);
or U48631 (N_48631,N_48450,N_48281);
xor U48632 (N_48632,N_48332,N_48323);
or U48633 (N_48633,N_48347,N_48264);
or U48634 (N_48634,N_48455,N_48491);
or U48635 (N_48635,N_48373,N_48366);
and U48636 (N_48636,N_48437,N_48254);
or U48637 (N_48637,N_48269,N_48462);
and U48638 (N_48638,N_48337,N_48356);
nor U48639 (N_48639,N_48333,N_48282);
nand U48640 (N_48640,N_48368,N_48352);
xor U48641 (N_48641,N_48331,N_48336);
or U48642 (N_48642,N_48494,N_48468);
or U48643 (N_48643,N_48288,N_48480);
xor U48644 (N_48644,N_48473,N_48411);
and U48645 (N_48645,N_48295,N_48322);
nand U48646 (N_48646,N_48444,N_48387);
and U48647 (N_48647,N_48308,N_48464);
nand U48648 (N_48648,N_48354,N_48286);
xor U48649 (N_48649,N_48308,N_48411);
or U48650 (N_48650,N_48268,N_48330);
nand U48651 (N_48651,N_48469,N_48453);
xnor U48652 (N_48652,N_48470,N_48356);
nand U48653 (N_48653,N_48268,N_48443);
nand U48654 (N_48654,N_48423,N_48324);
and U48655 (N_48655,N_48458,N_48296);
and U48656 (N_48656,N_48339,N_48290);
and U48657 (N_48657,N_48422,N_48266);
nand U48658 (N_48658,N_48429,N_48386);
nor U48659 (N_48659,N_48390,N_48486);
xor U48660 (N_48660,N_48442,N_48445);
or U48661 (N_48661,N_48250,N_48399);
nand U48662 (N_48662,N_48436,N_48441);
nand U48663 (N_48663,N_48367,N_48396);
and U48664 (N_48664,N_48283,N_48314);
xor U48665 (N_48665,N_48313,N_48490);
nor U48666 (N_48666,N_48352,N_48329);
nand U48667 (N_48667,N_48421,N_48301);
or U48668 (N_48668,N_48483,N_48444);
nand U48669 (N_48669,N_48347,N_48465);
or U48670 (N_48670,N_48475,N_48423);
and U48671 (N_48671,N_48293,N_48315);
and U48672 (N_48672,N_48493,N_48266);
xor U48673 (N_48673,N_48303,N_48364);
nor U48674 (N_48674,N_48469,N_48338);
nand U48675 (N_48675,N_48292,N_48462);
xnor U48676 (N_48676,N_48430,N_48488);
nand U48677 (N_48677,N_48399,N_48376);
and U48678 (N_48678,N_48260,N_48371);
nand U48679 (N_48679,N_48399,N_48303);
nor U48680 (N_48680,N_48290,N_48258);
nand U48681 (N_48681,N_48479,N_48437);
nand U48682 (N_48682,N_48257,N_48375);
or U48683 (N_48683,N_48324,N_48344);
nand U48684 (N_48684,N_48378,N_48289);
nand U48685 (N_48685,N_48254,N_48320);
xnor U48686 (N_48686,N_48393,N_48288);
nand U48687 (N_48687,N_48311,N_48429);
nor U48688 (N_48688,N_48462,N_48293);
and U48689 (N_48689,N_48382,N_48464);
nand U48690 (N_48690,N_48476,N_48431);
xor U48691 (N_48691,N_48459,N_48440);
nand U48692 (N_48692,N_48301,N_48332);
nor U48693 (N_48693,N_48368,N_48382);
nor U48694 (N_48694,N_48345,N_48358);
and U48695 (N_48695,N_48256,N_48374);
nand U48696 (N_48696,N_48497,N_48499);
xnor U48697 (N_48697,N_48458,N_48440);
and U48698 (N_48698,N_48377,N_48259);
nor U48699 (N_48699,N_48264,N_48370);
and U48700 (N_48700,N_48332,N_48453);
and U48701 (N_48701,N_48355,N_48263);
or U48702 (N_48702,N_48287,N_48337);
and U48703 (N_48703,N_48491,N_48417);
or U48704 (N_48704,N_48309,N_48329);
nor U48705 (N_48705,N_48366,N_48498);
nand U48706 (N_48706,N_48348,N_48334);
or U48707 (N_48707,N_48495,N_48277);
nor U48708 (N_48708,N_48270,N_48464);
and U48709 (N_48709,N_48428,N_48290);
nand U48710 (N_48710,N_48271,N_48315);
nor U48711 (N_48711,N_48256,N_48404);
xnor U48712 (N_48712,N_48348,N_48428);
nor U48713 (N_48713,N_48387,N_48383);
nand U48714 (N_48714,N_48363,N_48378);
or U48715 (N_48715,N_48364,N_48408);
nor U48716 (N_48716,N_48311,N_48475);
nand U48717 (N_48717,N_48477,N_48391);
or U48718 (N_48718,N_48293,N_48492);
xnor U48719 (N_48719,N_48388,N_48277);
nand U48720 (N_48720,N_48471,N_48331);
and U48721 (N_48721,N_48410,N_48384);
nand U48722 (N_48722,N_48403,N_48372);
nand U48723 (N_48723,N_48472,N_48483);
or U48724 (N_48724,N_48361,N_48319);
or U48725 (N_48725,N_48488,N_48389);
and U48726 (N_48726,N_48387,N_48288);
and U48727 (N_48727,N_48261,N_48327);
or U48728 (N_48728,N_48289,N_48496);
or U48729 (N_48729,N_48408,N_48345);
nor U48730 (N_48730,N_48275,N_48493);
or U48731 (N_48731,N_48285,N_48388);
xor U48732 (N_48732,N_48414,N_48491);
nand U48733 (N_48733,N_48290,N_48492);
nor U48734 (N_48734,N_48496,N_48366);
nor U48735 (N_48735,N_48418,N_48461);
xor U48736 (N_48736,N_48334,N_48313);
nor U48737 (N_48737,N_48418,N_48263);
xor U48738 (N_48738,N_48411,N_48299);
xor U48739 (N_48739,N_48403,N_48265);
nand U48740 (N_48740,N_48396,N_48363);
and U48741 (N_48741,N_48288,N_48474);
and U48742 (N_48742,N_48425,N_48455);
nor U48743 (N_48743,N_48288,N_48353);
or U48744 (N_48744,N_48370,N_48482);
and U48745 (N_48745,N_48481,N_48444);
nor U48746 (N_48746,N_48497,N_48371);
nor U48747 (N_48747,N_48434,N_48428);
and U48748 (N_48748,N_48397,N_48383);
nor U48749 (N_48749,N_48495,N_48351);
nor U48750 (N_48750,N_48610,N_48556);
or U48751 (N_48751,N_48741,N_48734);
or U48752 (N_48752,N_48545,N_48683);
and U48753 (N_48753,N_48566,N_48512);
xnor U48754 (N_48754,N_48694,N_48646);
or U48755 (N_48755,N_48716,N_48519);
nor U48756 (N_48756,N_48507,N_48739);
nand U48757 (N_48757,N_48723,N_48749);
and U48758 (N_48758,N_48670,N_48663);
nand U48759 (N_48759,N_48641,N_48665);
xnor U48760 (N_48760,N_48551,N_48648);
nand U48761 (N_48761,N_48601,N_48713);
or U48762 (N_48762,N_48509,N_48639);
and U48763 (N_48763,N_48701,N_48652);
xnor U48764 (N_48764,N_48668,N_48732);
xnor U48765 (N_48765,N_48687,N_48692);
nand U48766 (N_48766,N_48657,N_48618);
xor U48767 (N_48767,N_48638,N_48633);
and U48768 (N_48768,N_48585,N_48684);
and U48769 (N_48769,N_48743,N_48690);
nand U48770 (N_48770,N_48651,N_48516);
or U48771 (N_48771,N_48640,N_48600);
nor U48772 (N_48772,N_48700,N_48591);
nand U48773 (N_48773,N_48505,N_48559);
and U48774 (N_48774,N_48676,N_48696);
or U48775 (N_48775,N_48605,N_48531);
xor U48776 (N_48776,N_48537,N_48720);
xor U48777 (N_48777,N_48533,N_48616);
nor U48778 (N_48778,N_48607,N_48667);
nor U48779 (N_48779,N_48688,N_48654);
nor U48780 (N_48780,N_48634,N_48587);
or U48781 (N_48781,N_48513,N_48525);
or U48782 (N_48782,N_48706,N_48745);
nand U48783 (N_48783,N_48503,N_48504);
nor U48784 (N_48784,N_48589,N_48717);
nor U48785 (N_48785,N_48558,N_48727);
or U48786 (N_48786,N_48685,N_48562);
nor U48787 (N_48787,N_48658,N_48693);
or U48788 (N_48788,N_48575,N_48673);
xor U48789 (N_48789,N_48588,N_48666);
and U48790 (N_48790,N_48742,N_48532);
nand U48791 (N_48791,N_48695,N_48594);
xor U48792 (N_48792,N_48733,N_48674);
or U48793 (N_48793,N_48748,N_48655);
and U48794 (N_48794,N_48514,N_48747);
nand U48795 (N_48795,N_48584,N_48567);
nor U48796 (N_48796,N_48738,N_48619);
nor U48797 (N_48797,N_48520,N_48719);
xor U48798 (N_48798,N_48574,N_48730);
nor U48799 (N_48799,N_48539,N_48576);
nor U48800 (N_48800,N_48708,N_48511);
or U48801 (N_48801,N_48722,N_48538);
nand U48802 (N_48802,N_48623,N_48534);
or U48803 (N_48803,N_48593,N_48729);
nand U48804 (N_48804,N_48595,N_48526);
nor U48805 (N_48805,N_48523,N_48680);
nor U48806 (N_48806,N_48647,N_48596);
xnor U48807 (N_48807,N_48582,N_48677);
or U48808 (N_48808,N_48535,N_48697);
or U48809 (N_48809,N_48645,N_48564);
and U48810 (N_48810,N_48675,N_48579);
or U48811 (N_48811,N_48698,N_48703);
nor U48812 (N_48812,N_48571,N_48548);
xor U48813 (N_48813,N_48624,N_48592);
and U48814 (N_48814,N_48608,N_48530);
and U48815 (N_48815,N_48536,N_48546);
nand U48816 (N_48816,N_48614,N_48662);
xor U48817 (N_48817,N_48678,N_48615);
nand U48818 (N_48818,N_48631,N_48500);
nor U48819 (N_48819,N_48553,N_48661);
and U48820 (N_48820,N_48554,N_48570);
and U48821 (N_48821,N_48609,N_48613);
nand U48822 (N_48822,N_48737,N_48621);
nor U48823 (N_48823,N_48656,N_48635);
and U48824 (N_48824,N_48502,N_48578);
and U48825 (N_48825,N_48515,N_48522);
and U48826 (N_48826,N_48599,N_48630);
or U48827 (N_48827,N_48524,N_48603);
xor U48828 (N_48828,N_48671,N_48714);
and U48829 (N_48829,N_48625,N_48644);
or U48830 (N_48830,N_48726,N_48707);
xnor U48831 (N_48831,N_48510,N_48577);
or U48832 (N_48832,N_48547,N_48682);
xnor U48833 (N_48833,N_48606,N_48542);
and U48834 (N_48834,N_48517,N_48724);
xor U48835 (N_48835,N_48552,N_48628);
xor U48836 (N_48836,N_48728,N_48506);
nand U48837 (N_48837,N_48629,N_48681);
nand U48838 (N_48838,N_48583,N_48598);
xnor U48839 (N_48839,N_48527,N_48710);
xnor U48840 (N_48840,N_48731,N_48543);
or U48841 (N_48841,N_48611,N_48622);
or U48842 (N_48842,N_48528,N_48541);
or U48843 (N_48843,N_48555,N_48550);
nor U48844 (N_48844,N_48508,N_48721);
and U48845 (N_48845,N_48705,N_48557);
nor U48846 (N_48846,N_48620,N_48521);
nand U48847 (N_48847,N_48540,N_48612);
or U48848 (N_48848,N_48735,N_48712);
xnor U48849 (N_48849,N_48626,N_48632);
xor U48850 (N_48850,N_48581,N_48672);
xor U48851 (N_48851,N_48560,N_48740);
nand U48852 (N_48852,N_48602,N_48649);
and U48853 (N_48853,N_48709,N_48636);
and U48854 (N_48854,N_48699,N_48660);
xor U48855 (N_48855,N_48573,N_48718);
nor U48856 (N_48856,N_48704,N_48691);
nand U48857 (N_48857,N_48586,N_48580);
or U48858 (N_48858,N_48746,N_48563);
nand U48859 (N_48859,N_48650,N_48653);
and U48860 (N_48860,N_48597,N_48617);
nand U48861 (N_48861,N_48568,N_48637);
nand U48862 (N_48862,N_48549,N_48604);
or U48863 (N_48863,N_48643,N_48669);
nor U48864 (N_48864,N_48518,N_48569);
or U48865 (N_48865,N_48561,N_48702);
nand U48866 (N_48866,N_48659,N_48572);
or U48867 (N_48867,N_48501,N_48642);
xor U48868 (N_48868,N_48686,N_48711);
xnor U48869 (N_48869,N_48627,N_48736);
nor U48870 (N_48870,N_48715,N_48725);
nand U48871 (N_48871,N_48744,N_48664);
xnor U48872 (N_48872,N_48565,N_48590);
and U48873 (N_48873,N_48689,N_48529);
nor U48874 (N_48874,N_48544,N_48679);
or U48875 (N_48875,N_48604,N_48696);
nor U48876 (N_48876,N_48612,N_48565);
nand U48877 (N_48877,N_48687,N_48677);
nand U48878 (N_48878,N_48579,N_48534);
xnor U48879 (N_48879,N_48525,N_48622);
and U48880 (N_48880,N_48618,N_48679);
or U48881 (N_48881,N_48558,N_48623);
nor U48882 (N_48882,N_48545,N_48744);
xor U48883 (N_48883,N_48546,N_48621);
and U48884 (N_48884,N_48539,N_48530);
xnor U48885 (N_48885,N_48561,N_48551);
nand U48886 (N_48886,N_48653,N_48528);
nand U48887 (N_48887,N_48617,N_48690);
or U48888 (N_48888,N_48531,N_48674);
and U48889 (N_48889,N_48625,N_48696);
xor U48890 (N_48890,N_48615,N_48688);
or U48891 (N_48891,N_48600,N_48703);
nor U48892 (N_48892,N_48517,N_48548);
or U48893 (N_48893,N_48609,N_48515);
xnor U48894 (N_48894,N_48584,N_48535);
nand U48895 (N_48895,N_48641,N_48518);
or U48896 (N_48896,N_48504,N_48663);
xnor U48897 (N_48897,N_48506,N_48700);
or U48898 (N_48898,N_48669,N_48745);
and U48899 (N_48899,N_48531,N_48722);
nand U48900 (N_48900,N_48742,N_48644);
nor U48901 (N_48901,N_48741,N_48588);
and U48902 (N_48902,N_48644,N_48629);
or U48903 (N_48903,N_48673,N_48569);
nand U48904 (N_48904,N_48555,N_48722);
or U48905 (N_48905,N_48725,N_48616);
or U48906 (N_48906,N_48620,N_48686);
nor U48907 (N_48907,N_48698,N_48673);
or U48908 (N_48908,N_48553,N_48662);
or U48909 (N_48909,N_48633,N_48673);
and U48910 (N_48910,N_48566,N_48526);
xnor U48911 (N_48911,N_48594,N_48511);
and U48912 (N_48912,N_48729,N_48530);
nand U48913 (N_48913,N_48630,N_48725);
xnor U48914 (N_48914,N_48556,N_48727);
and U48915 (N_48915,N_48507,N_48514);
nor U48916 (N_48916,N_48583,N_48521);
or U48917 (N_48917,N_48718,N_48708);
or U48918 (N_48918,N_48672,N_48556);
xor U48919 (N_48919,N_48728,N_48707);
xor U48920 (N_48920,N_48671,N_48680);
and U48921 (N_48921,N_48609,N_48675);
nor U48922 (N_48922,N_48524,N_48534);
nor U48923 (N_48923,N_48545,N_48566);
xor U48924 (N_48924,N_48633,N_48711);
and U48925 (N_48925,N_48742,N_48505);
nor U48926 (N_48926,N_48708,N_48612);
nor U48927 (N_48927,N_48701,N_48552);
nand U48928 (N_48928,N_48588,N_48592);
nand U48929 (N_48929,N_48728,N_48715);
and U48930 (N_48930,N_48706,N_48557);
nor U48931 (N_48931,N_48551,N_48660);
or U48932 (N_48932,N_48599,N_48512);
nand U48933 (N_48933,N_48670,N_48621);
xor U48934 (N_48934,N_48733,N_48506);
and U48935 (N_48935,N_48672,N_48502);
and U48936 (N_48936,N_48716,N_48654);
nor U48937 (N_48937,N_48543,N_48711);
xor U48938 (N_48938,N_48666,N_48656);
nor U48939 (N_48939,N_48550,N_48509);
nand U48940 (N_48940,N_48737,N_48590);
or U48941 (N_48941,N_48606,N_48621);
nand U48942 (N_48942,N_48612,N_48711);
xor U48943 (N_48943,N_48681,N_48727);
and U48944 (N_48944,N_48549,N_48652);
or U48945 (N_48945,N_48617,N_48588);
and U48946 (N_48946,N_48639,N_48576);
nand U48947 (N_48947,N_48691,N_48535);
nand U48948 (N_48948,N_48645,N_48547);
xor U48949 (N_48949,N_48737,N_48545);
nor U48950 (N_48950,N_48703,N_48665);
nor U48951 (N_48951,N_48721,N_48529);
and U48952 (N_48952,N_48717,N_48565);
or U48953 (N_48953,N_48509,N_48587);
xnor U48954 (N_48954,N_48748,N_48735);
nor U48955 (N_48955,N_48662,N_48586);
nor U48956 (N_48956,N_48576,N_48552);
or U48957 (N_48957,N_48745,N_48510);
or U48958 (N_48958,N_48505,N_48734);
xnor U48959 (N_48959,N_48540,N_48604);
or U48960 (N_48960,N_48681,N_48660);
nand U48961 (N_48961,N_48560,N_48504);
nand U48962 (N_48962,N_48591,N_48606);
or U48963 (N_48963,N_48558,N_48667);
xnor U48964 (N_48964,N_48694,N_48584);
and U48965 (N_48965,N_48615,N_48533);
nor U48966 (N_48966,N_48733,N_48511);
or U48967 (N_48967,N_48603,N_48636);
xor U48968 (N_48968,N_48590,N_48690);
and U48969 (N_48969,N_48572,N_48715);
or U48970 (N_48970,N_48628,N_48601);
xor U48971 (N_48971,N_48555,N_48707);
xnor U48972 (N_48972,N_48523,N_48530);
xor U48973 (N_48973,N_48679,N_48643);
xor U48974 (N_48974,N_48680,N_48542);
xnor U48975 (N_48975,N_48746,N_48573);
nand U48976 (N_48976,N_48628,N_48508);
nor U48977 (N_48977,N_48701,N_48603);
nor U48978 (N_48978,N_48615,N_48552);
nor U48979 (N_48979,N_48540,N_48500);
and U48980 (N_48980,N_48721,N_48627);
and U48981 (N_48981,N_48719,N_48652);
and U48982 (N_48982,N_48624,N_48701);
and U48983 (N_48983,N_48534,N_48739);
nor U48984 (N_48984,N_48569,N_48534);
nor U48985 (N_48985,N_48597,N_48686);
and U48986 (N_48986,N_48500,N_48684);
nor U48987 (N_48987,N_48583,N_48748);
or U48988 (N_48988,N_48538,N_48647);
xor U48989 (N_48989,N_48608,N_48598);
nor U48990 (N_48990,N_48548,N_48586);
nor U48991 (N_48991,N_48659,N_48555);
or U48992 (N_48992,N_48636,N_48595);
and U48993 (N_48993,N_48583,N_48512);
nand U48994 (N_48994,N_48702,N_48616);
nor U48995 (N_48995,N_48522,N_48704);
or U48996 (N_48996,N_48576,N_48600);
xor U48997 (N_48997,N_48714,N_48542);
or U48998 (N_48998,N_48651,N_48645);
nand U48999 (N_48999,N_48546,N_48656);
and U49000 (N_49000,N_48795,N_48988);
nand U49001 (N_49001,N_48943,N_48913);
xor U49002 (N_49002,N_48750,N_48780);
or U49003 (N_49003,N_48857,N_48965);
or U49004 (N_49004,N_48837,N_48937);
or U49005 (N_49005,N_48847,N_48761);
nor U49006 (N_49006,N_48918,N_48753);
nand U49007 (N_49007,N_48898,N_48982);
xor U49008 (N_49008,N_48910,N_48811);
xor U49009 (N_49009,N_48779,N_48916);
xor U49010 (N_49010,N_48802,N_48815);
xor U49011 (N_49011,N_48980,N_48940);
nand U49012 (N_49012,N_48759,N_48899);
xor U49013 (N_49013,N_48975,N_48853);
nand U49014 (N_49014,N_48990,N_48850);
and U49015 (N_49015,N_48941,N_48809);
and U49016 (N_49016,N_48773,N_48801);
and U49017 (N_49017,N_48754,N_48889);
nand U49018 (N_49018,N_48876,N_48823);
nor U49019 (N_49019,N_48909,N_48999);
xor U49020 (N_49020,N_48901,N_48820);
nand U49021 (N_49021,N_48917,N_48813);
and U49022 (N_49022,N_48832,N_48862);
and U49023 (N_49023,N_48954,N_48922);
nand U49024 (N_49024,N_48961,N_48814);
xor U49025 (N_49025,N_48981,N_48788);
and U49026 (N_49026,N_48984,N_48936);
or U49027 (N_49027,N_48894,N_48785);
xor U49028 (N_49028,N_48839,N_48855);
xor U49029 (N_49029,N_48828,N_48911);
xor U49030 (N_49030,N_48864,N_48849);
and U49031 (N_49031,N_48931,N_48793);
and U49032 (N_49032,N_48883,N_48893);
xor U49033 (N_49033,N_48992,N_48873);
or U49034 (N_49034,N_48960,N_48880);
xnor U49035 (N_49035,N_48778,N_48775);
or U49036 (N_49036,N_48919,N_48970);
xor U49037 (N_49037,N_48907,N_48956);
or U49038 (N_49038,N_48926,N_48781);
or U49039 (N_49039,N_48867,N_48854);
xnor U49040 (N_49040,N_48962,N_48987);
and U49041 (N_49041,N_48914,N_48900);
nor U49042 (N_49042,N_48859,N_48787);
or U49043 (N_49043,N_48957,N_48763);
or U49044 (N_49044,N_48924,N_48772);
and U49045 (N_49045,N_48797,N_48819);
or U49046 (N_49046,N_48833,N_48966);
nor U49047 (N_49047,N_48794,N_48861);
xnor U49048 (N_49048,N_48782,N_48963);
xor U49049 (N_49049,N_48929,N_48891);
nand U49050 (N_49050,N_48791,N_48969);
nor U49051 (N_49051,N_48959,N_48755);
nor U49052 (N_49052,N_48783,N_48856);
nand U49053 (N_49053,N_48824,N_48865);
and U49054 (N_49054,N_48805,N_48902);
xnor U49055 (N_49055,N_48868,N_48757);
and U49056 (N_49056,N_48946,N_48971);
xor U49057 (N_49057,N_48996,N_48774);
nor U49058 (N_49058,N_48938,N_48886);
and U49059 (N_49059,N_48756,N_48817);
and U49060 (N_49060,N_48858,N_48986);
and U49061 (N_49061,N_48766,N_48895);
nand U49062 (N_49062,N_48945,N_48993);
nor U49063 (N_49063,N_48892,N_48870);
and U49064 (N_49064,N_48994,N_48927);
xor U49065 (N_49065,N_48792,N_48968);
nor U49066 (N_49066,N_48933,N_48770);
and U49067 (N_49067,N_48767,N_48838);
and U49068 (N_49068,N_48997,N_48798);
or U49069 (N_49069,N_48897,N_48974);
xor U49070 (N_49070,N_48860,N_48950);
nand U49071 (N_49071,N_48840,N_48752);
xor U49072 (N_49072,N_48796,N_48842);
or U49073 (N_49073,N_48978,N_48942);
and U49074 (N_49074,N_48885,N_48915);
xor U49075 (N_49075,N_48808,N_48935);
and U49076 (N_49076,N_48998,N_48836);
and U49077 (N_49077,N_48863,N_48851);
and U49078 (N_49078,N_48983,N_48958);
nand U49079 (N_49079,N_48869,N_48777);
xnor U49080 (N_49080,N_48800,N_48948);
nand U49081 (N_49081,N_48769,N_48822);
nor U49082 (N_49082,N_48947,N_48989);
and U49083 (N_49083,N_48825,N_48789);
xor U49084 (N_49084,N_48920,N_48830);
and U49085 (N_49085,N_48827,N_48964);
xnor U49086 (N_49086,N_48806,N_48934);
xnor U49087 (N_49087,N_48848,N_48804);
or U49088 (N_49088,N_48818,N_48887);
nand U49089 (N_49089,N_48835,N_48829);
xnor U49090 (N_49090,N_48939,N_48955);
xor U49091 (N_49091,N_48784,N_48764);
nand U49092 (N_49092,N_48803,N_48826);
nor U49093 (N_49093,N_48786,N_48888);
xnor U49094 (N_49094,N_48921,N_48890);
or U49095 (N_49095,N_48991,N_48874);
and U49096 (N_49096,N_48768,N_48845);
or U49097 (N_49097,N_48771,N_48760);
or U49098 (N_49098,N_48758,N_48879);
nand U49099 (N_49099,N_48904,N_48765);
xor U49100 (N_49100,N_48790,N_48831);
nand U49101 (N_49101,N_48751,N_48925);
xor U49102 (N_49102,N_48967,N_48979);
or U49103 (N_49103,N_48973,N_48846);
xnor U49104 (N_49104,N_48810,N_48912);
and U49105 (N_49105,N_48816,N_48821);
xnor U49106 (N_49106,N_48812,N_48799);
nand U49107 (N_49107,N_48976,N_48896);
and U49108 (N_49108,N_48906,N_48871);
nand U49109 (N_49109,N_48951,N_48844);
nor U49110 (N_49110,N_48923,N_48977);
xnor U49111 (N_49111,N_48881,N_48877);
and U49112 (N_49112,N_48834,N_48882);
nor U49113 (N_49113,N_48884,N_48905);
or U49114 (N_49114,N_48908,N_48932);
and U49115 (N_49115,N_48843,N_48872);
and U49116 (N_49116,N_48985,N_48930);
nor U49117 (N_49117,N_48878,N_48944);
or U49118 (N_49118,N_48928,N_48866);
and U49119 (N_49119,N_48841,N_48776);
xnor U49120 (N_49120,N_48972,N_48807);
nand U49121 (N_49121,N_48762,N_48852);
nand U49122 (N_49122,N_48903,N_48953);
nor U49123 (N_49123,N_48952,N_48949);
xnor U49124 (N_49124,N_48875,N_48995);
or U49125 (N_49125,N_48946,N_48880);
nor U49126 (N_49126,N_48914,N_48932);
or U49127 (N_49127,N_48939,N_48914);
and U49128 (N_49128,N_48835,N_48916);
xnor U49129 (N_49129,N_48864,N_48859);
or U49130 (N_49130,N_48942,N_48884);
or U49131 (N_49131,N_48786,N_48814);
nor U49132 (N_49132,N_48800,N_48881);
nor U49133 (N_49133,N_48891,N_48837);
nand U49134 (N_49134,N_48843,N_48926);
or U49135 (N_49135,N_48897,N_48779);
and U49136 (N_49136,N_48984,N_48835);
nand U49137 (N_49137,N_48875,N_48963);
nand U49138 (N_49138,N_48973,N_48780);
or U49139 (N_49139,N_48791,N_48902);
nor U49140 (N_49140,N_48791,N_48779);
or U49141 (N_49141,N_48851,N_48794);
nor U49142 (N_49142,N_48911,N_48832);
or U49143 (N_49143,N_48916,N_48980);
xnor U49144 (N_49144,N_48955,N_48752);
nand U49145 (N_49145,N_48875,N_48796);
or U49146 (N_49146,N_48919,N_48827);
xor U49147 (N_49147,N_48880,N_48996);
nand U49148 (N_49148,N_48778,N_48809);
nand U49149 (N_49149,N_48870,N_48863);
xnor U49150 (N_49150,N_48909,N_48983);
and U49151 (N_49151,N_48917,N_48955);
nand U49152 (N_49152,N_48884,N_48769);
nor U49153 (N_49153,N_48908,N_48887);
or U49154 (N_49154,N_48782,N_48904);
nor U49155 (N_49155,N_48986,N_48803);
and U49156 (N_49156,N_48904,N_48833);
or U49157 (N_49157,N_48915,N_48767);
and U49158 (N_49158,N_48881,N_48785);
and U49159 (N_49159,N_48929,N_48942);
or U49160 (N_49160,N_48842,N_48770);
and U49161 (N_49161,N_48829,N_48860);
or U49162 (N_49162,N_48916,N_48816);
nand U49163 (N_49163,N_48793,N_48767);
nor U49164 (N_49164,N_48771,N_48861);
and U49165 (N_49165,N_48949,N_48904);
or U49166 (N_49166,N_48782,N_48980);
nand U49167 (N_49167,N_48793,N_48989);
and U49168 (N_49168,N_48888,N_48856);
or U49169 (N_49169,N_48761,N_48870);
nor U49170 (N_49170,N_48922,N_48968);
xor U49171 (N_49171,N_48787,N_48776);
xor U49172 (N_49172,N_48964,N_48935);
or U49173 (N_49173,N_48892,N_48896);
nand U49174 (N_49174,N_48918,N_48926);
and U49175 (N_49175,N_48769,N_48758);
nand U49176 (N_49176,N_48894,N_48927);
nand U49177 (N_49177,N_48835,N_48993);
nor U49178 (N_49178,N_48958,N_48975);
xor U49179 (N_49179,N_48830,N_48948);
or U49180 (N_49180,N_48878,N_48953);
nor U49181 (N_49181,N_48891,N_48777);
nand U49182 (N_49182,N_48977,N_48855);
xnor U49183 (N_49183,N_48787,N_48977);
nor U49184 (N_49184,N_48917,N_48841);
nor U49185 (N_49185,N_48995,N_48819);
xor U49186 (N_49186,N_48955,N_48857);
nand U49187 (N_49187,N_48940,N_48820);
or U49188 (N_49188,N_48944,N_48821);
nand U49189 (N_49189,N_48869,N_48865);
and U49190 (N_49190,N_48775,N_48932);
xor U49191 (N_49191,N_48968,N_48996);
and U49192 (N_49192,N_48952,N_48958);
and U49193 (N_49193,N_48999,N_48926);
nor U49194 (N_49194,N_48779,N_48788);
or U49195 (N_49195,N_48786,N_48843);
xnor U49196 (N_49196,N_48882,N_48855);
nor U49197 (N_49197,N_48957,N_48884);
nor U49198 (N_49198,N_48977,N_48782);
nand U49199 (N_49199,N_48847,N_48964);
nor U49200 (N_49200,N_48759,N_48926);
nor U49201 (N_49201,N_48871,N_48965);
and U49202 (N_49202,N_48885,N_48830);
nand U49203 (N_49203,N_48934,N_48940);
nor U49204 (N_49204,N_48896,N_48827);
nand U49205 (N_49205,N_48790,N_48994);
and U49206 (N_49206,N_48772,N_48783);
nor U49207 (N_49207,N_48817,N_48979);
nand U49208 (N_49208,N_48947,N_48963);
nand U49209 (N_49209,N_48934,N_48820);
nor U49210 (N_49210,N_48774,N_48892);
xnor U49211 (N_49211,N_48929,N_48949);
and U49212 (N_49212,N_48757,N_48883);
and U49213 (N_49213,N_48784,N_48935);
or U49214 (N_49214,N_48994,N_48796);
xor U49215 (N_49215,N_48817,N_48754);
or U49216 (N_49216,N_48809,N_48894);
or U49217 (N_49217,N_48920,N_48770);
xnor U49218 (N_49218,N_48961,N_48972);
nand U49219 (N_49219,N_48792,N_48923);
nand U49220 (N_49220,N_48865,N_48916);
and U49221 (N_49221,N_48841,N_48855);
and U49222 (N_49222,N_48957,N_48752);
xnor U49223 (N_49223,N_48876,N_48922);
nand U49224 (N_49224,N_48974,N_48871);
nor U49225 (N_49225,N_48985,N_48990);
nand U49226 (N_49226,N_48914,N_48786);
nor U49227 (N_49227,N_48761,N_48936);
and U49228 (N_49228,N_48938,N_48795);
and U49229 (N_49229,N_48806,N_48939);
nand U49230 (N_49230,N_48946,N_48923);
and U49231 (N_49231,N_48759,N_48988);
or U49232 (N_49232,N_48927,N_48882);
nor U49233 (N_49233,N_48843,N_48867);
nand U49234 (N_49234,N_48873,N_48860);
or U49235 (N_49235,N_48926,N_48795);
or U49236 (N_49236,N_48822,N_48837);
nor U49237 (N_49237,N_48862,N_48947);
and U49238 (N_49238,N_48812,N_48929);
nand U49239 (N_49239,N_48957,N_48933);
nand U49240 (N_49240,N_48822,N_48912);
nand U49241 (N_49241,N_48952,N_48921);
nor U49242 (N_49242,N_48899,N_48866);
and U49243 (N_49243,N_48978,N_48957);
and U49244 (N_49244,N_48987,N_48951);
nand U49245 (N_49245,N_48789,N_48759);
nand U49246 (N_49246,N_48827,N_48920);
or U49247 (N_49247,N_48871,N_48915);
or U49248 (N_49248,N_48991,N_48944);
xor U49249 (N_49249,N_48931,N_48889);
or U49250 (N_49250,N_49050,N_49230);
nor U49251 (N_49251,N_49075,N_49129);
and U49252 (N_49252,N_49150,N_49169);
nor U49253 (N_49253,N_49202,N_49176);
nand U49254 (N_49254,N_49056,N_49045);
or U49255 (N_49255,N_49030,N_49091);
or U49256 (N_49256,N_49248,N_49163);
or U49257 (N_49257,N_49022,N_49216);
nor U49258 (N_49258,N_49242,N_49212);
and U49259 (N_49259,N_49191,N_49170);
and U49260 (N_49260,N_49178,N_49117);
or U49261 (N_49261,N_49018,N_49090);
xor U49262 (N_49262,N_49138,N_49131);
xor U49263 (N_49263,N_49013,N_49246);
xor U49264 (N_49264,N_49136,N_49168);
xnor U49265 (N_49265,N_49137,N_49140);
xor U49266 (N_49266,N_49162,N_49145);
or U49267 (N_49267,N_49244,N_49128);
nand U49268 (N_49268,N_49038,N_49132);
or U49269 (N_49269,N_49002,N_49061);
xnor U49270 (N_49270,N_49243,N_49160);
nand U49271 (N_49271,N_49206,N_49194);
nand U49272 (N_49272,N_49098,N_49188);
nand U49273 (N_49273,N_49103,N_49161);
nand U49274 (N_49274,N_49070,N_49186);
nor U49275 (N_49275,N_49035,N_49153);
nand U49276 (N_49276,N_49174,N_49009);
xor U49277 (N_49277,N_49042,N_49021);
or U49278 (N_49278,N_49172,N_49029);
nand U49279 (N_49279,N_49052,N_49193);
nor U49280 (N_49280,N_49204,N_49014);
and U49281 (N_49281,N_49236,N_49184);
or U49282 (N_49282,N_49210,N_49154);
xnor U49283 (N_49283,N_49127,N_49112);
or U49284 (N_49284,N_49234,N_49100);
nand U49285 (N_49285,N_49088,N_49064);
nor U49286 (N_49286,N_49196,N_49225);
or U49287 (N_49287,N_49200,N_49177);
and U49288 (N_49288,N_49031,N_49116);
and U49289 (N_49289,N_49181,N_49007);
or U49290 (N_49290,N_49115,N_49211);
xnor U49291 (N_49291,N_49074,N_49036);
nand U49292 (N_49292,N_49123,N_49134);
xnor U49293 (N_49293,N_49054,N_49105);
nand U49294 (N_49294,N_49155,N_49060);
xor U49295 (N_49295,N_49109,N_49228);
nand U49296 (N_49296,N_49003,N_49034);
xnor U49297 (N_49297,N_49231,N_49093);
nor U49298 (N_49298,N_49240,N_49201);
nand U49299 (N_49299,N_49040,N_49152);
nor U49300 (N_49300,N_49179,N_49025);
and U49301 (N_49301,N_49151,N_49180);
and U49302 (N_49302,N_49183,N_49104);
xor U49303 (N_49303,N_49032,N_49141);
xor U49304 (N_49304,N_49110,N_49222);
nor U49305 (N_49305,N_49121,N_49187);
nor U49306 (N_49306,N_49233,N_49048);
or U49307 (N_49307,N_49023,N_49059);
nand U49308 (N_49308,N_49107,N_49096);
or U49309 (N_49309,N_49017,N_49041);
xnor U49310 (N_49310,N_49185,N_49080);
xor U49311 (N_49311,N_49111,N_49227);
xnor U49312 (N_49312,N_49192,N_49114);
xor U49313 (N_49313,N_49006,N_49232);
or U49314 (N_49314,N_49239,N_49106);
or U49315 (N_49315,N_49043,N_49218);
xnor U49316 (N_49316,N_49195,N_49076);
nor U49317 (N_49317,N_49024,N_49118);
nor U49318 (N_49318,N_49004,N_49143);
and U49319 (N_49319,N_49081,N_49078);
or U49320 (N_49320,N_49083,N_49235);
xor U49321 (N_49321,N_49000,N_49166);
nor U49322 (N_49322,N_49208,N_49011);
or U49323 (N_49323,N_49084,N_49085);
xor U49324 (N_49324,N_49010,N_49205);
nor U49325 (N_49325,N_49092,N_49245);
xnor U49326 (N_49326,N_49033,N_49207);
xor U49327 (N_49327,N_49217,N_49028);
nand U49328 (N_49328,N_49058,N_49069);
nor U49329 (N_49329,N_49005,N_49016);
xor U49330 (N_49330,N_49167,N_49126);
or U49331 (N_49331,N_49019,N_49102);
nor U49332 (N_49332,N_49214,N_49063);
nand U49333 (N_49333,N_49146,N_49125);
nor U49334 (N_49334,N_49008,N_49158);
and U49335 (N_49335,N_49237,N_49182);
nand U49336 (N_49336,N_49144,N_49148);
and U49337 (N_49337,N_49055,N_49164);
nor U49338 (N_49338,N_49097,N_49073);
or U49339 (N_49339,N_49124,N_49209);
xor U49340 (N_49340,N_49087,N_49101);
nand U49341 (N_49341,N_49213,N_49203);
xor U49342 (N_49342,N_49037,N_49071);
or U49343 (N_49343,N_49086,N_49229);
nand U49344 (N_49344,N_49047,N_49122);
xor U49345 (N_49345,N_49249,N_49119);
xor U49346 (N_49346,N_49130,N_49175);
or U49347 (N_49347,N_49051,N_49068);
nand U49348 (N_49348,N_49082,N_49039);
and U49349 (N_49349,N_49099,N_49062);
or U49350 (N_49350,N_49226,N_49215);
nor U49351 (N_49351,N_49015,N_49142);
and U49352 (N_49352,N_49089,N_49095);
nor U49353 (N_49353,N_49190,N_49113);
xor U49354 (N_49354,N_49149,N_49012);
nand U49355 (N_49355,N_49147,N_49139);
or U49356 (N_49356,N_49065,N_49156);
nor U49357 (N_49357,N_49077,N_49238);
nand U49358 (N_49358,N_49133,N_49072);
and U49359 (N_49359,N_49157,N_49057);
nor U49360 (N_49360,N_49221,N_49198);
nand U49361 (N_49361,N_49049,N_49165);
nand U49362 (N_49362,N_49197,N_49094);
and U49363 (N_49363,N_49247,N_49189);
nand U49364 (N_49364,N_49223,N_49120);
nand U49365 (N_49365,N_49219,N_49066);
nand U49366 (N_49366,N_49199,N_49108);
xor U49367 (N_49367,N_49224,N_49027);
and U49368 (N_49368,N_49053,N_49173);
or U49369 (N_49369,N_49046,N_49241);
and U49370 (N_49370,N_49001,N_49067);
and U49371 (N_49371,N_49171,N_49044);
xnor U49372 (N_49372,N_49135,N_49079);
or U49373 (N_49373,N_49159,N_49220);
nand U49374 (N_49374,N_49026,N_49020);
nor U49375 (N_49375,N_49213,N_49085);
or U49376 (N_49376,N_49017,N_49181);
xor U49377 (N_49377,N_49135,N_49239);
and U49378 (N_49378,N_49046,N_49072);
or U49379 (N_49379,N_49162,N_49194);
nand U49380 (N_49380,N_49066,N_49068);
nor U49381 (N_49381,N_49144,N_49127);
and U49382 (N_49382,N_49061,N_49117);
nor U49383 (N_49383,N_49213,N_49016);
nor U49384 (N_49384,N_49114,N_49229);
or U49385 (N_49385,N_49065,N_49110);
or U49386 (N_49386,N_49065,N_49205);
and U49387 (N_49387,N_49018,N_49110);
nor U49388 (N_49388,N_49214,N_49167);
nand U49389 (N_49389,N_49030,N_49061);
or U49390 (N_49390,N_49162,N_49140);
xor U49391 (N_49391,N_49092,N_49035);
and U49392 (N_49392,N_49200,N_49159);
and U49393 (N_49393,N_49113,N_49060);
and U49394 (N_49394,N_49223,N_49093);
xor U49395 (N_49395,N_49005,N_49227);
or U49396 (N_49396,N_49085,N_49215);
and U49397 (N_49397,N_49138,N_49086);
nand U49398 (N_49398,N_49224,N_49181);
and U49399 (N_49399,N_49111,N_49202);
and U49400 (N_49400,N_49179,N_49245);
and U49401 (N_49401,N_49217,N_49204);
and U49402 (N_49402,N_49073,N_49218);
and U49403 (N_49403,N_49159,N_49053);
nor U49404 (N_49404,N_49237,N_49230);
nand U49405 (N_49405,N_49177,N_49039);
and U49406 (N_49406,N_49186,N_49187);
nand U49407 (N_49407,N_49113,N_49017);
nand U49408 (N_49408,N_49222,N_49010);
and U49409 (N_49409,N_49042,N_49148);
nand U49410 (N_49410,N_49188,N_49195);
xnor U49411 (N_49411,N_49078,N_49029);
nand U49412 (N_49412,N_49221,N_49072);
nand U49413 (N_49413,N_49026,N_49103);
nand U49414 (N_49414,N_49138,N_49072);
nor U49415 (N_49415,N_49093,N_49159);
nor U49416 (N_49416,N_49115,N_49056);
nand U49417 (N_49417,N_49156,N_49106);
nand U49418 (N_49418,N_49165,N_49198);
nor U49419 (N_49419,N_49068,N_49031);
and U49420 (N_49420,N_49015,N_49247);
xnor U49421 (N_49421,N_49181,N_49043);
and U49422 (N_49422,N_49152,N_49098);
and U49423 (N_49423,N_49161,N_49050);
or U49424 (N_49424,N_49243,N_49195);
or U49425 (N_49425,N_49205,N_49126);
and U49426 (N_49426,N_49202,N_49057);
nor U49427 (N_49427,N_49023,N_49117);
nor U49428 (N_49428,N_49219,N_49214);
xnor U49429 (N_49429,N_49175,N_49222);
or U49430 (N_49430,N_49104,N_49163);
nor U49431 (N_49431,N_49124,N_49170);
nor U49432 (N_49432,N_49075,N_49084);
nand U49433 (N_49433,N_49241,N_49034);
nand U49434 (N_49434,N_49043,N_49184);
or U49435 (N_49435,N_49249,N_49169);
or U49436 (N_49436,N_49096,N_49223);
or U49437 (N_49437,N_49154,N_49058);
nor U49438 (N_49438,N_49093,N_49035);
xnor U49439 (N_49439,N_49142,N_49069);
or U49440 (N_49440,N_49191,N_49054);
or U49441 (N_49441,N_49227,N_49058);
nor U49442 (N_49442,N_49072,N_49086);
or U49443 (N_49443,N_49090,N_49187);
xnor U49444 (N_49444,N_49194,N_49200);
and U49445 (N_49445,N_49014,N_49128);
and U49446 (N_49446,N_49161,N_49234);
nor U49447 (N_49447,N_49198,N_49145);
nand U49448 (N_49448,N_49149,N_49192);
nor U49449 (N_49449,N_49046,N_49215);
or U49450 (N_49450,N_49008,N_49216);
or U49451 (N_49451,N_49225,N_49230);
nand U49452 (N_49452,N_49156,N_49203);
or U49453 (N_49453,N_49201,N_49096);
nand U49454 (N_49454,N_49073,N_49172);
nand U49455 (N_49455,N_49245,N_49058);
or U49456 (N_49456,N_49233,N_49038);
xor U49457 (N_49457,N_49009,N_49005);
nor U49458 (N_49458,N_49156,N_49009);
nor U49459 (N_49459,N_49066,N_49079);
xnor U49460 (N_49460,N_49241,N_49157);
nor U49461 (N_49461,N_49082,N_49232);
and U49462 (N_49462,N_49195,N_49055);
nor U49463 (N_49463,N_49174,N_49084);
nand U49464 (N_49464,N_49065,N_49028);
nand U49465 (N_49465,N_49192,N_49216);
or U49466 (N_49466,N_49203,N_49135);
or U49467 (N_49467,N_49015,N_49191);
or U49468 (N_49468,N_49033,N_49061);
nor U49469 (N_49469,N_49149,N_49190);
nand U49470 (N_49470,N_49236,N_49220);
or U49471 (N_49471,N_49195,N_49080);
and U49472 (N_49472,N_49150,N_49200);
and U49473 (N_49473,N_49058,N_49046);
nand U49474 (N_49474,N_49109,N_49011);
nor U49475 (N_49475,N_49232,N_49153);
nand U49476 (N_49476,N_49030,N_49016);
xor U49477 (N_49477,N_49148,N_49218);
or U49478 (N_49478,N_49011,N_49155);
xor U49479 (N_49479,N_49073,N_49087);
nor U49480 (N_49480,N_49152,N_49141);
xor U49481 (N_49481,N_49204,N_49187);
xor U49482 (N_49482,N_49127,N_49034);
or U49483 (N_49483,N_49035,N_49107);
nor U49484 (N_49484,N_49133,N_49099);
or U49485 (N_49485,N_49237,N_49157);
nor U49486 (N_49486,N_49023,N_49027);
nand U49487 (N_49487,N_49044,N_49124);
and U49488 (N_49488,N_49073,N_49125);
or U49489 (N_49489,N_49101,N_49224);
xor U49490 (N_49490,N_49191,N_49145);
nor U49491 (N_49491,N_49197,N_49040);
xor U49492 (N_49492,N_49112,N_49170);
and U49493 (N_49493,N_49074,N_49052);
nand U49494 (N_49494,N_49191,N_49045);
nor U49495 (N_49495,N_49144,N_49101);
xor U49496 (N_49496,N_49101,N_49219);
xnor U49497 (N_49497,N_49223,N_49177);
nor U49498 (N_49498,N_49049,N_49158);
xnor U49499 (N_49499,N_49181,N_49035);
or U49500 (N_49500,N_49497,N_49347);
and U49501 (N_49501,N_49361,N_49398);
and U49502 (N_49502,N_49300,N_49329);
xor U49503 (N_49503,N_49443,N_49385);
nand U49504 (N_49504,N_49280,N_49404);
and U49505 (N_49505,N_49486,N_49317);
xnor U49506 (N_49506,N_49344,N_49428);
and U49507 (N_49507,N_49367,N_49415);
and U49508 (N_49508,N_49402,N_49292);
nor U49509 (N_49509,N_49424,N_49348);
and U49510 (N_49510,N_49384,N_49283);
and U49511 (N_49511,N_49396,N_49430);
xnor U49512 (N_49512,N_49416,N_49250);
and U49513 (N_49513,N_49299,N_49418);
xor U49514 (N_49514,N_49407,N_49305);
or U49515 (N_49515,N_49286,N_49267);
xor U49516 (N_49516,N_49436,N_49343);
nand U49517 (N_49517,N_49442,N_49307);
xnor U49518 (N_49518,N_49293,N_49496);
and U49519 (N_49519,N_49399,N_49282);
nand U49520 (N_49520,N_49324,N_49439);
nor U49521 (N_49521,N_49391,N_49304);
or U49522 (N_49522,N_49482,N_49381);
or U49523 (N_49523,N_49359,N_49409);
or U49524 (N_49524,N_49272,N_49278);
and U49525 (N_49525,N_49448,N_49354);
and U49526 (N_49526,N_49403,N_49392);
nor U49527 (N_49527,N_49301,N_49370);
xnor U49528 (N_49528,N_49291,N_49360);
and U49529 (N_49529,N_49334,N_49472);
xor U49530 (N_49530,N_49390,N_49444);
or U49531 (N_49531,N_49440,N_49437);
xnor U49532 (N_49532,N_49376,N_49422);
or U49533 (N_49533,N_49426,N_49449);
nor U49534 (N_49534,N_49254,N_49251);
or U49535 (N_49535,N_49258,N_49308);
xnor U49536 (N_49536,N_49340,N_49289);
nor U49537 (N_49537,N_49431,N_49253);
and U49538 (N_49538,N_49413,N_49446);
and U49539 (N_49539,N_49479,N_49471);
or U49540 (N_49540,N_49260,N_49460);
and U49541 (N_49541,N_49310,N_49372);
nor U49542 (N_49542,N_49332,N_49255);
and U49543 (N_49543,N_49458,N_49447);
and U49544 (N_49544,N_49394,N_49427);
and U49545 (N_49545,N_49429,N_49388);
or U49546 (N_49546,N_49259,N_49269);
nor U49547 (N_49547,N_49397,N_49420);
nand U49548 (N_49548,N_49454,N_49288);
and U49549 (N_49549,N_49369,N_49281);
nand U49550 (N_49550,N_49349,N_49295);
xnor U49551 (N_49551,N_49457,N_49389);
xor U49552 (N_49552,N_49466,N_49461);
xor U49553 (N_49553,N_49363,N_49306);
and U49554 (N_49554,N_49355,N_49333);
nand U49555 (N_49555,N_49365,N_49277);
xor U49556 (N_49556,N_49316,N_49287);
and U49557 (N_49557,N_49284,N_49336);
xnor U49558 (N_49558,N_49473,N_49346);
and U49559 (N_49559,N_49405,N_49262);
nor U49560 (N_49560,N_49469,N_49495);
xnor U49561 (N_49561,N_49393,N_49474);
nor U49562 (N_49562,N_49483,N_49468);
xnor U49563 (N_49563,N_49445,N_49320);
or U49564 (N_49564,N_49450,N_49325);
nand U49565 (N_49565,N_49314,N_49465);
nand U49566 (N_49566,N_49331,N_49345);
or U49567 (N_49567,N_49493,N_49414);
nor U49568 (N_49568,N_49475,N_49356);
xor U49569 (N_49569,N_49432,N_49326);
or U49570 (N_49570,N_49358,N_49321);
nand U49571 (N_49571,N_49273,N_49408);
and U49572 (N_49572,N_49387,N_49480);
and U49573 (N_49573,N_49290,N_49268);
nand U49574 (N_49574,N_49476,N_49406);
nand U49575 (N_49575,N_49419,N_49338);
and U49576 (N_49576,N_49276,N_49411);
nand U49577 (N_49577,N_49341,N_49371);
xnor U49578 (N_49578,N_49382,N_49318);
nor U49579 (N_49579,N_49252,N_49484);
nor U49580 (N_49580,N_49434,N_49377);
and U49581 (N_49581,N_49279,N_49378);
or U49582 (N_49582,N_49265,N_49350);
or U49583 (N_49583,N_49417,N_49463);
nand U49584 (N_49584,N_49271,N_49395);
and U49585 (N_49585,N_49335,N_49261);
or U49586 (N_49586,N_49488,N_49491);
and U49587 (N_49587,N_49368,N_49400);
and U49588 (N_49588,N_49313,N_49297);
and U49589 (N_49589,N_49453,N_49485);
nor U49590 (N_49590,N_49353,N_49494);
nand U49591 (N_49591,N_49330,N_49380);
xor U49592 (N_49592,N_49489,N_49328);
nor U49593 (N_49593,N_49364,N_49425);
and U49594 (N_49594,N_49423,N_49303);
or U49595 (N_49595,N_49375,N_49478);
and U49596 (N_49596,N_49319,N_49256);
or U49597 (N_49597,N_49481,N_49309);
nand U49598 (N_49598,N_49302,N_49357);
nand U49599 (N_49599,N_49455,N_49492);
xor U49600 (N_49600,N_49421,N_49470);
and U49601 (N_49601,N_49459,N_49352);
xnor U49602 (N_49602,N_49477,N_49339);
or U49603 (N_49603,N_49499,N_49412);
xor U49604 (N_49604,N_49383,N_49315);
nand U49605 (N_49605,N_49337,N_49373);
or U49606 (N_49606,N_49498,N_49285);
and U49607 (N_49607,N_49327,N_49274);
xor U49608 (N_49608,N_49464,N_49467);
and U49609 (N_49609,N_49270,N_49462);
or U49610 (N_49610,N_49323,N_49401);
or U49611 (N_49611,N_49351,N_49257);
nor U49612 (N_49612,N_49266,N_49490);
nor U49613 (N_49613,N_49452,N_49379);
nor U49614 (N_49614,N_49366,N_49362);
and U49615 (N_49615,N_49322,N_49456);
and U49616 (N_49616,N_49298,N_49435);
xor U49617 (N_49617,N_49438,N_49487);
nor U49618 (N_49618,N_49294,N_49451);
or U49619 (N_49619,N_49433,N_49296);
xnor U49620 (N_49620,N_49263,N_49441);
nand U49621 (N_49621,N_49374,N_49342);
and U49622 (N_49622,N_49275,N_49311);
nor U49623 (N_49623,N_49386,N_49312);
or U49624 (N_49624,N_49410,N_49264);
and U49625 (N_49625,N_49399,N_49371);
nand U49626 (N_49626,N_49461,N_49476);
nor U49627 (N_49627,N_49361,N_49345);
xor U49628 (N_49628,N_49487,N_49302);
nand U49629 (N_49629,N_49440,N_49393);
and U49630 (N_49630,N_49436,N_49251);
or U49631 (N_49631,N_49424,N_49395);
nand U49632 (N_49632,N_49356,N_49366);
and U49633 (N_49633,N_49391,N_49373);
xnor U49634 (N_49634,N_49268,N_49296);
xor U49635 (N_49635,N_49384,N_49262);
and U49636 (N_49636,N_49335,N_49344);
or U49637 (N_49637,N_49467,N_49339);
and U49638 (N_49638,N_49482,N_49298);
nand U49639 (N_49639,N_49464,N_49325);
or U49640 (N_49640,N_49395,N_49321);
or U49641 (N_49641,N_49315,N_49318);
xnor U49642 (N_49642,N_49378,N_49486);
or U49643 (N_49643,N_49271,N_49482);
and U49644 (N_49644,N_49374,N_49499);
xor U49645 (N_49645,N_49428,N_49255);
or U49646 (N_49646,N_49272,N_49471);
xor U49647 (N_49647,N_49458,N_49493);
nand U49648 (N_49648,N_49267,N_49430);
or U49649 (N_49649,N_49252,N_49439);
nor U49650 (N_49650,N_49491,N_49332);
or U49651 (N_49651,N_49351,N_49271);
xor U49652 (N_49652,N_49403,N_49442);
or U49653 (N_49653,N_49424,N_49366);
nor U49654 (N_49654,N_49258,N_49402);
or U49655 (N_49655,N_49296,N_49498);
or U49656 (N_49656,N_49484,N_49282);
or U49657 (N_49657,N_49388,N_49392);
or U49658 (N_49658,N_49312,N_49419);
or U49659 (N_49659,N_49491,N_49396);
xnor U49660 (N_49660,N_49297,N_49428);
and U49661 (N_49661,N_49482,N_49350);
xnor U49662 (N_49662,N_49456,N_49429);
or U49663 (N_49663,N_49416,N_49426);
xnor U49664 (N_49664,N_49364,N_49374);
or U49665 (N_49665,N_49266,N_49379);
or U49666 (N_49666,N_49459,N_49476);
xor U49667 (N_49667,N_49390,N_49462);
or U49668 (N_49668,N_49458,N_49343);
nor U49669 (N_49669,N_49384,N_49263);
nor U49670 (N_49670,N_49273,N_49416);
nand U49671 (N_49671,N_49486,N_49281);
and U49672 (N_49672,N_49318,N_49280);
or U49673 (N_49673,N_49418,N_49420);
and U49674 (N_49674,N_49420,N_49292);
nor U49675 (N_49675,N_49473,N_49453);
nand U49676 (N_49676,N_49269,N_49394);
nor U49677 (N_49677,N_49430,N_49302);
nand U49678 (N_49678,N_49260,N_49294);
nor U49679 (N_49679,N_49419,N_49388);
and U49680 (N_49680,N_49384,N_49388);
or U49681 (N_49681,N_49456,N_49491);
xor U49682 (N_49682,N_49427,N_49462);
and U49683 (N_49683,N_49436,N_49483);
and U49684 (N_49684,N_49331,N_49310);
or U49685 (N_49685,N_49342,N_49432);
nor U49686 (N_49686,N_49354,N_49489);
xnor U49687 (N_49687,N_49486,N_49316);
nor U49688 (N_49688,N_49262,N_49288);
nor U49689 (N_49689,N_49419,N_49418);
and U49690 (N_49690,N_49444,N_49263);
and U49691 (N_49691,N_49255,N_49411);
nand U49692 (N_49692,N_49298,N_49465);
and U49693 (N_49693,N_49346,N_49469);
nor U49694 (N_49694,N_49477,N_49355);
nor U49695 (N_49695,N_49384,N_49443);
nor U49696 (N_49696,N_49342,N_49423);
and U49697 (N_49697,N_49319,N_49310);
and U49698 (N_49698,N_49323,N_49426);
or U49699 (N_49699,N_49463,N_49420);
nor U49700 (N_49700,N_49361,N_49338);
xor U49701 (N_49701,N_49384,N_49354);
nor U49702 (N_49702,N_49266,N_49462);
xor U49703 (N_49703,N_49329,N_49463);
nor U49704 (N_49704,N_49311,N_49430);
nand U49705 (N_49705,N_49468,N_49297);
and U49706 (N_49706,N_49297,N_49296);
or U49707 (N_49707,N_49355,N_49331);
nor U49708 (N_49708,N_49303,N_49407);
xor U49709 (N_49709,N_49327,N_49390);
nor U49710 (N_49710,N_49290,N_49425);
nor U49711 (N_49711,N_49424,N_49374);
nand U49712 (N_49712,N_49437,N_49443);
nor U49713 (N_49713,N_49476,N_49346);
nor U49714 (N_49714,N_49265,N_49392);
nor U49715 (N_49715,N_49439,N_49485);
or U49716 (N_49716,N_49380,N_49393);
or U49717 (N_49717,N_49261,N_49309);
nand U49718 (N_49718,N_49383,N_49465);
nor U49719 (N_49719,N_49314,N_49383);
or U49720 (N_49720,N_49493,N_49445);
nand U49721 (N_49721,N_49368,N_49250);
xnor U49722 (N_49722,N_49372,N_49393);
and U49723 (N_49723,N_49337,N_49429);
and U49724 (N_49724,N_49253,N_49304);
nor U49725 (N_49725,N_49327,N_49444);
nor U49726 (N_49726,N_49494,N_49399);
nand U49727 (N_49727,N_49296,N_49291);
nand U49728 (N_49728,N_49495,N_49453);
or U49729 (N_49729,N_49480,N_49349);
nor U49730 (N_49730,N_49313,N_49470);
xor U49731 (N_49731,N_49311,N_49457);
nand U49732 (N_49732,N_49444,N_49426);
or U49733 (N_49733,N_49442,N_49408);
nor U49734 (N_49734,N_49417,N_49307);
nand U49735 (N_49735,N_49463,N_49332);
and U49736 (N_49736,N_49313,N_49271);
and U49737 (N_49737,N_49417,N_49273);
nor U49738 (N_49738,N_49315,N_49381);
xor U49739 (N_49739,N_49475,N_49302);
nand U49740 (N_49740,N_49290,N_49266);
nor U49741 (N_49741,N_49326,N_49431);
nor U49742 (N_49742,N_49327,N_49420);
or U49743 (N_49743,N_49441,N_49362);
xnor U49744 (N_49744,N_49251,N_49454);
nor U49745 (N_49745,N_49358,N_49465);
or U49746 (N_49746,N_49466,N_49256);
and U49747 (N_49747,N_49345,N_49267);
or U49748 (N_49748,N_49425,N_49297);
and U49749 (N_49749,N_49275,N_49307);
xnor U49750 (N_49750,N_49509,N_49616);
nor U49751 (N_49751,N_49700,N_49698);
nor U49752 (N_49752,N_49599,N_49578);
nand U49753 (N_49753,N_49736,N_49602);
and U49754 (N_49754,N_49635,N_49615);
nand U49755 (N_49755,N_49746,N_49657);
and U49756 (N_49756,N_49683,N_49526);
nand U49757 (N_49757,N_49735,N_49690);
and U49758 (N_49758,N_49650,N_49513);
or U49759 (N_49759,N_49640,N_49653);
nor U49760 (N_49760,N_49638,N_49505);
nor U49761 (N_49761,N_49636,N_49600);
nand U49762 (N_49762,N_49612,N_49730);
nand U49763 (N_49763,N_49576,N_49745);
xnor U49764 (N_49764,N_49644,N_49579);
and U49765 (N_49765,N_49682,N_49610);
nor U49766 (N_49766,N_49622,N_49703);
and U49767 (N_49767,N_49500,N_49572);
or U49768 (N_49768,N_49715,N_49611);
xnor U49769 (N_49769,N_49727,N_49570);
nor U49770 (N_49770,N_49660,N_49627);
and U49771 (N_49771,N_49713,N_49726);
nor U49772 (N_49772,N_49580,N_49714);
nor U49773 (N_49773,N_49749,N_49641);
nand U49774 (N_49774,N_49514,N_49667);
xor U49775 (N_49775,N_49603,N_49665);
and U49776 (N_49776,N_49654,N_49606);
xor U49777 (N_49777,N_49691,N_49701);
nand U49778 (N_49778,N_49720,N_49681);
nor U49779 (N_49779,N_49569,N_49629);
and U49780 (N_49780,N_49733,N_49742);
xor U49781 (N_49781,N_49687,N_49740);
or U49782 (N_49782,N_49540,N_49567);
xnor U49783 (N_49783,N_49680,N_49621);
xnor U49784 (N_49784,N_49674,N_49577);
xor U49785 (N_49785,N_49739,N_49707);
nand U49786 (N_49786,N_49668,N_49624);
xor U49787 (N_49787,N_49520,N_49672);
and U49788 (N_49788,N_49547,N_49656);
nand U49789 (N_49789,N_49523,N_49689);
and U49790 (N_49790,N_49688,N_49573);
nor U49791 (N_49791,N_49722,N_49531);
and U49792 (N_49792,N_49702,N_49659);
and U49793 (N_49793,N_49619,N_49594);
nand U49794 (N_49794,N_49601,N_49634);
or U49795 (N_49795,N_49614,N_49537);
or U49796 (N_49796,N_49558,N_49585);
and U49797 (N_49797,N_49539,N_49504);
or U49798 (N_49798,N_49618,N_49534);
and U49799 (N_49799,N_49670,N_49632);
xnor U49800 (N_49800,N_49516,N_49512);
nand U49801 (N_49801,N_49710,N_49637);
nor U49802 (N_49802,N_49533,N_49506);
nor U49803 (N_49803,N_49661,N_49719);
nand U49804 (N_49804,N_49718,N_49507);
or U49805 (N_49805,N_49593,N_49652);
nand U49806 (N_49806,N_49598,N_49566);
xnor U49807 (N_49807,N_49518,N_49723);
nand U49808 (N_49808,N_49528,N_49519);
and U49809 (N_49809,N_49663,N_49548);
xor U49810 (N_49810,N_49625,N_49743);
xnor U49811 (N_49811,N_49527,N_49729);
nand U49812 (N_49812,N_49676,N_49511);
and U49813 (N_49813,N_49704,N_49510);
and U49814 (N_49814,N_49669,N_49550);
and U49815 (N_49815,N_49628,N_49554);
nand U49816 (N_49816,N_49515,N_49673);
xnor U49817 (N_49817,N_49604,N_49535);
xor U49818 (N_49818,N_49582,N_49648);
nand U49819 (N_49819,N_49544,N_49574);
or U49820 (N_49820,N_49725,N_49607);
nor U49821 (N_49821,N_49711,N_49524);
nor U49822 (N_49822,N_49630,N_49522);
xnor U49823 (N_49823,N_49595,N_49732);
nor U49824 (N_49824,N_49609,N_49541);
nor U49825 (N_49825,N_49590,N_49643);
or U49826 (N_49826,N_49646,N_49737);
xnor U49827 (N_49827,N_49734,N_49645);
or U49828 (N_49828,N_49555,N_49664);
xnor U49829 (N_49829,N_49716,N_49708);
nor U49830 (N_49830,N_49697,N_49561);
nor U49831 (N_49831,N_49557,N_49530);
and U49832 (N_49832,N_49532,N_49583);
nor U49833 (N_49833,N_49684,N_49542);
and U49834 (N_49834,N_49748,N_49658);
or U49835 (N_49835,N_49731,N_49695);
and U49836 (N_49836,N_49596,N_49693);
nand U49837 (N_49837,N_49545,N_49575);
or U49838 (N_49838,N_49508,N_49705);
and U49839 (N_49839,N_49696,N_49551);
nand U49840 (N_49840,N_49563,N_49623);
and U49841 (N_49841,N_49581,N_49543);
or U49842 (N_49842,N_49568,N_49562);
xnor U49843 (N_49843,N_49529,N_49503);
or U49844 (N_49844,N_49559,N_49564);
or U49845 (N_49845,N_49709,N_49571);
nor U49846 (N_49846,N_49589,N_49741);
or U49847 (N_49847,N_49592,N_49671);
and U49848 (N_49848,N_49738,N_49678);
and U49849 (N_49849,N_49662,N_49605);
xor U49850 (N_49850,N_49565,N_49501);
nor U49851 (N_49851,N_49728,N_49631);
or U49852 (N_49852,N_49620,N_49626);
or U49853 (N_49853,N_49706,N_49666);
nor U49854 (N_49854,N_49699,N_49694);
xnor U49855 (N_49855,N_49591,N_49686);
xor U49856 (N_49856,N_49608,N_49502);
or U49857 (N_49857,N_49717,N_49647);
xor U49858 (N_49858,N_49556,N_49549);
and U49859 (N_49859,N_49685,N_49552);
nor U49860 (N_49860,N_49649,N_49538);
xnor U49861 (N_49861,N_49517,N_49747);
or U49862 (N_49862,N_49642,N_49692);
nor U49863 (N_49863,N_49521,N_49724);
or U49864 (N_49864,N_49744,N_49536);
xor U49865 (N_49865,N_49546,N_49712);
xor U49866 (N_49866,N_49584,N_49553);
and U49867 (N_49867,N_49679,N_49633);
nand U49868 (N_49868,N_49721,N_49639);
nand U49869 (N_49869,N_49587,N_49525);
nor U49870 (N_49870,N_49675,N_49597);
nand U49871 (N_49871,N_49617,N_49655);
nor U49872 (N_49872,N_49651,N_49588);
xnor U49873 (N_49873,N_49677,N_49586);
nand U49874 (N_49874,N_49613,N_49560);
nand U49875 (N_49875,N_49515,N_49724);
nor U49876 (N_49876,N_49617,N_49711);
nand U49877 (N_49877,N_49676,N_49677);
nor U49878 (N_49878,N_49673,N_49716);
nor U49879 (N_49879,N_49588,N_49595);
and U49880 (N_49880,N_49719,N_49632);
nand U49881 (N_49881,N_49558,N_49523);
nand U49882 (N_49882,N_49725,N_49698);
or U49883 (N_49883,N_49545,N_49577);
nor U49884 (N_49884,N_49615,N_49645);
nor U49885 (N_49885,N_49739,N_49583);
nand U49886 (N_49886,N_49703,N_49604);
nor U49887 (N_49887,N_49517,N_49578);
and U49888 (N_49888,N_49662,N_49515);
or U49889 (N_49889,N_49708,N_49725);
nand U49890 (N_49890,N_49534,N_49555);
nand U49891 (N_49891,N_49700,N_49694);
nand U49892 (N_49892,N_49718,N_49533);
or U49893 (N_49893,N_49503,N_49581);
or U49894 (N_49894,N_49660,N_49720);
or U49895 (N_49895,N_49693,N_49658);
and U49896 (N_49896,N_49617,N_49544);
or U49897 (N_49897,N_49712,N_49566);
and U49898 (N_49898,N_49525,N_49572);
or U49899 (N_49899,N_49657,N_49651);
nor U49900 (N_49900,N_49584,N_49677);
xor U49901 (N_49901,N_49608,N_49520);
nand U49902 (N_49902,N_49734,N_49666);
and U49903 (N_49903,N_49596,N_49707);
and U49904 (N_49904,N_49743,N_49630);
nor U49905 (N_49905,N_49572,N_49564);
xnor U49906 (N_49906,N_49673,N_49698);
xor U49907 (N_49907,N_49607,N_49694);
nand U49908 (N_49908,N_49710,N_49611);
nor U49909 (N_49909,N_49586,N_49653);
and U49910 (N_49910,N_49563,N_49670);
or U49911 (N_49911,N_49609,N_49596);
xor U49912 (N_49912,N_49667,N_49548);
xnor U49913 (N_49913,N_49561,N_49518);
nand U49914 (N_49914,N_49740,N_49533);
and U49915 (N_49915,N_49586,N_49692);
nor U49916 (N_49916,N_49698,N_49622);
and U49917 (N_49917,N_49519,N_49590);
or U49918 (N_49918,N_49510,N_49526);
and U49919 (N_49919,N_49615,N_49643);
nand U49920 (N_49920,N_49565,N_49630);
nor U49921 (N_49921,N_49563,N_49648);
and U49922 (N_49922,N_49612,N_49702);
nand U49923 (N_49923,N_49588,N_49512);
or U49924 (N_49924,N_49694,N_49551);
and U49925 (N_49925,N_49506,N_49528);
and U49926 (N_49926,N_49611,N_49606);
nor U49927 (N_49927,N_49721,N_49728);
or U49928 (N_49928,N_49704,N_49676);
or U49929 (N_49929,N_49524,N_49683);
nand U49930 (N_49930,N_49611,N_49563);
xor U49931 (N_49931,N_49670,N_49641);
or U49932 (N_49932,N_49505,N_49534);
xnor U49933 (N_49933,N_49642,N_49525);
or U49934 (N_49934,N_49662,N_49571);
xor U49935 (N_49935,N_49594,N_49729);
xor U49936 (N_49936,N_49508,N_49603);
and U49937 (N_49937,N_49633,N_49563);
or U49938 (N_49938,N_49545,N_49602);
and U49939 (N_49939,N_49690,N_49501);
and U49940 (N_49940,N_49557,N_49592);
and U49941 (N_49941,N_49656,N_49521);
nand U49942 (N_49942,N_49617,N_49591);
and U49943 (N_49943,N_49740,N_49628);
or U49944 (N_49944,N_49614,N_49619);
or U49945 (N_49945,N_49652,N_49509);
nor U49946 (N_49946,N_49744,N_49632);
nand U49947 (N_49947,N_49637,N_49552);
or U49948 (N_49948,N_49523,N_49747);
and U49949 (N_49949,N_49621,N_49652);
nor U49950 (N_49950,N_49684,N_49547);
or U49951 (N_49951,N_49556,N_49519);
nor U49952 (N_49952,N_49666,N_49621);
or U49953 (N_49953,N_49556,N_49547);
nor U49954 (N_49954,N_49728,N_49540);
and U49955 (N_49955,N_49528,N_49684);
nand U49956 (N_49956,N_49507,N_49715);
or U49957 (N_49957,N_49654,N_49689);
nor U49958 (N_49958,N_49655,N_49726);
and U49959 (N_49959,N_49540,N_49685);
nor U49960 (N_49960,N_49614,N_49570);
and U49961 (N_49961,N_49537,N_49553);
nor U49962 (N_49962,N_49535,N_49572);
xor U49963 (N_49963,N_49725,N_49512);
xnor U49964 (N_49964,N_49668,N_49659);
nor U49965 (N_49965,N_49657,N_49516);
or U49966 (N_49966,N_49539,N_49683);
nand U49967 (N_49967,N_49717,N_49528);
nand U49968 (N_49968,N_49737,N_49587);
nor U49969 (N_49969,N_49709,N_49718);
and U49970 (N_49970,N_49515,N_49617);
and U49971 (N_49971,N_49500,N_49674);
nand U49972 (N_49972,N_49720,N_49661);
nor U49973 (N_49973,N_49695,N_49654);
or U49974 (N_49974,N_49717,N_49598);
and U49975 (N_49975,N_49650,N_49541);
and U49976 (N_49976,N_49541,N_49733);
xor U49977 (N_49977,N_49745,N_49705);
xnor U49978 (N_49978,N_49557,N_49702);
xnor U49979 (N_49979,N_49536,N_49529);
nand U49980 (N_49980,N_49638,N_49564);
nand U49981 (N_49981,N_49573,N_49713);
or U49982 (N_49982,N_49552,N_49535);
or U49983 (N_49983,N_49664,N_49594);
or U49984 (N_49984,N_49723,N_49564);
and U49985 (N_49985,N_49604,N_49723);
nand U49986 (N_49986,N_49524,N_49695);
nand U49987 (N_49987,N_49649,N_49585);
and U49988 (N_49988,N_49589,N_49567);
xor U49989 (N_49989,N_49663,N_49687);
nand U49990 (N_49990,N_49749,N_49658);
xnor U49991 (N_49991,N_49535,N_49555);
or U49992 (N_49992,N_49727,N_49566);
xor U49993 (N_49993,N_49660,N_49522);
nand U49994 (N_49994,N_49695,N_49661);
xnor U49995 (N_49995,N_49674,N_49709);
xnor U49996 (N_49996,N_49721,N_49589);
nand U49997 (N_49997,N_49551,N_49593);
nor U49998 (N_49998,N_49664,N_49675);
and U49999 (N_49999,N_49636,N_49700);
nand UO_0 (O_0,N_49990,N_49839);
xor UO_1 (O_1,N_49797,N_49964);
nor UO_2 (O_2,N_49836,N_49965);
xor UO_3 (O_3,N_49763,N_49943);
nand UO_4 (O_4,N_49944,N_49800);
nor UO_5 (O_5,N_49981,N_49808);
nand UO_6 (O_6,N_49805,N_49818);
or UO_7 (O_7,N_49774,N_49766);
nand UO_8 (O_8,N_49760,N_49927);
xnor UO_9 (O_9,N_49933,N_49866);
nor UO_10 (O_10,N_49863,N_49849);
xnor UO_11 (O_11,N_49779,N_49916);
nand UO_12 (O_12,N_49857,N_49770);
and UO_13 (O_13,N_49977,N_49974);
nand UO_14 (O_14,N_49895,N_49903);
and UO_15 (O_15,N_49949,N_49835);
nor UO_16 (O_16,N_49906,N_49784);
nor UO_17 (O_17,N_49987,N_49781);
or UO_18 (O_18,N_49907,N_49796);
nor UO_19 (O_19,N_49850,N_49798);
and UO_20 (O_20,N_49844,N_49862);
nor UO_21 (O_21,N_49956,N_49861);
nor UO_22 (O_22,N_49997,N_49832);
or UO_23 (O_23,N_49958,N_49915);
and UO_24 (O_24,N_49864,N_49820);
xor UO_25 (O_25,N_49950,N_49754);
or UO_26 (O_26,N_49834,N_49919);
xor UO_27 (O_27,N_49829,N_49999);
or UO_28 (O_28,N_49817,N_49790);
or UO_29 (O_29,N_49822,N_49802);
nand UO_30 (O_30,N_49904,N_49752);
and UO_31 (O_31,N_49924,N_49876);
nand UO_32 (O_32,N_49967,N_49815);
nor UO_33 (O_33,N_49942,N_49828);
xnor UO_34 (O_34,N_49898,N_49940);
or UO_35 (O_35,N_49966,N_49877);
or UO_36 (O_36,N_49914,N_49750);
xor UO_37 (O_37,N_49890,N_49871);
nor UO_38 (O_38,N_49778,N_49755);
or UO_39 (O_39,N_49757,N_49908);
and UO_40 (O_40,N_49994,N_49762);
xor UO_41 (O_41,N_49892,N_49771);
xor UO_42 (O_42,N_49992,N_49773);
nor UO_43 (O_43,N_49792,N_49955);
xnor UO_44 (O_44,N_49780,N_49759);
nand UO_45 (O_45,N_49772,N_49957);
and UO_46 (O_46,N_49920,N_49970);
nor UO_47 (O_47,N_49851,N_49870);
nor UO_48 (O_48,N_49941,N_49925);
nand UO_49 (O_49,N_49803,N_49806);
nor UO_50 (O_50,N_49804,N_49969);
and UO_51 (O_51,N_49991,N_49926);
nor UO_52 (O_52,N_49913,N_49872);
and UO_53 (O_53,N_49810,N_49888);
or UO_54 (O_54,N_49910,N_49900);
or UO_55 (O_55,N_49794,N_49945);
xnor UO_56 (O_56,N_49935,N_49983);
and UO_57 (O_57,N_49859,N_49911);
nand UO_58 (O_58,N_49962,N_49909);
and UO_59 (O_59,N_49756,N_49824);
nand UO_60 (O_60,N_49972,N_49886);
nor UO_61 (O_61,N_49827,N_49880);
nor UO_62 (O_62,N_49936,N_49881);
or UO_63 (O_63,N_49833,N_49782);
nand UO_64 (O_64,N_49947,N_49982);
nor UO_65 (O_65,N_49894,N_49858);
nand UO_66 (O_66,N_49998,N_49793);
and UO_67 (O_67,N_49865,N_49874);
or UO_68 (O_68,N_49901,N_49812);
nor UO_69 (O_69,N_49801,N_49985);
or UO_70 (O_70,N_49786,N_49830);
nor UO_71 (O_71,N_49954,N_49795);
xor UO_72 (O_72,N_49825,N_49845);
xor UO_73 (O_73,N_49893,N_49768);
nand UO_74 (O_74,N_49921,N_49873);
or UO_75 (O_75,N_49897,N_49867);
nand UO_76 (O_76,N_49842,N_49847);
xnor UO_77 (O_77,N_49975,N_49878);
or UO_78 (O_78,N_49889,N_49785);
and UO_79 (O_79,N_49860,N_49930);
xor UO_80 (O_80,N_49996,N_49995);
or UO_81 (O_81,N_49971,N_49918);
and UO_82 (O_82,N_49751,N_49789);
or UO_83 (O_83,N_49929,N_49846);
and UO_84 (O_84,N_49978,N_49905);
or UO_85 (O_85,N_49765,N_49776);
or UO_86 (O_86,N_49869,N_49960);
nand UO_87 (O_87,N_49896,N_49788);
or UO_88 (O_88,N_49952,N_49931);
and UO_89 (O_89,N_49767,N_49988);
or UO_90 (O_90,N_49753,N_49769);
or UO_91 (O_91,N_49807,N_49912);
or UO_92 (O_92,N_49986,N_49875);
nor UO_93 (O_93,N_49814,N_49917);
and UO_94 (O_94,N_49813,N_49946);
xor UO_95 (O_95,N_49973,N_49843);
xor UO_96 (O_96,N_49968,N_49882);
nor UO_97 (O_97,N_49791,N_49938);
xnor UO_98 (O_98,N_49821,N_49826);
nor UO_99 (O_99,N_49979,N_49984);
or UO_100 (O_100,N_49887,N_49959);
nand UO_101 (O_101,N_49838,N_49848);
and UO_102 (O_102,N_49799,N_49856);
xnor UO_103 (O_103,N_49932,N_49823);
and UO_104 (O_104,N_49922,N_49923);
nand UO_105 (O_105,N_49837,N_49855);
and UO_106 (O_106,N_49840,N_49891);
nor UO_107 (O_107,N_49899,N_49775);
and UO_108 (O_108,N_49761,N_49811);
nand UO_109 (O_109,N_49853,N_49883);
xnor UO_110 (O_110,N_49854,N_49777);
nor UO_111 (O_111,N_49963,N_49758);
xor UO_112 (O_112,N_49939,N_49809);
xor UO_113 (O_113,N_49783,N_49764);
or UO_114 (O_114,N_49868,N_49879);
and UO_115 (O_115,N_49787,N_49819);
nand UO_116 (O_116,N_49928,N_49989);
or UO_117 (O_117,N_49852,N_49816);
and UO_118 (O_118,N_49831,N_49841);
and UO_119 (O_119,N_49902,N_49885);
xnor UO_120 (O_120,N_49980,N_49976);
or UO_121 (O_121,N_49948,N_49951);
nor UO_122 (O_122,N_49993,N_49961);
or UO_123 (O_123,N_49934,N_49937);
xnor UO_124 (O_124,N_49884,N_49953);
or UO_125 (O_125,N_49759,N_49837);
xor UO_126 (O_126,N_49836,N_49899);
xnor UO_127 (O_127,N_49943,N_49836);
xor UO_128 (O_128,N_49762,N_49920);
nand UO_129 (O_129,N_49983,N_49817);
xor UO_130 (O_130,N_49812,N_49987);
nand UO_131 (O_131,N_49809,N_49874);
nor UO_132 (O_132,N_49975,N_49877);
nor UO_133 (O_133,N_49957,N_49972);
nand UO_134 (O_134,N_49836,N_49801);
nor UO_135 (O_135,N_49964,N_49840);
nor UO_136 (O_136,N_49880,N_49956);
nand UO_137 (O_137,N_49846,N_49821);
and UO_138 (O_138,N_49811,N_49950);
xnor UO_139 (O_139,N_49923,N_49887);
nand UO_140 (O_140,N_49854,N_49856);
and UO_141 (O_141,N_49813,N_49907);
and UO_142 (O_142,N_49879,N_49796);
nand UO_143 (O_143,N_49760,N_49922);
and UO_144 (O_144,N_49990,N_49841);
xor UO_145 (O_145,N_49933,N_49952);
xnor UO_146 (O_146,N_49787,N_49926);
nor UO_147 (O_147,N_49750,N_49926);
nand UO_148 (O_148,N_49868,N_49825);
or UO_149 (O_149,N_49899,N_49975);
and UO_150 (O_150,N_49945,N_49820);
or UO_151 (O_151,N_49801,N_49768);
nand UO_152 (O_152,N_49932,N_49892);
xor UO_153 (O_153,N_49862,N_49923);
and UO_154 (O_154,N_49927,N_49775);
xor UO_155 (O_155,N_49786,N_49875);
or UO_156 (O_156,N_49887,N_49956);
nand UO_157 (O_157,N_49984,N_49915);
xnor UO_158 (O_158,N_49768,N_49958);
and UO_159 (O_159,N_49887,N_49908);
or UO_160 (O_160,N_49788,N_49943);
xor UO_161 (O_161,N_49819,N_49803);
nor UO_162 (O_162,N_49836,N_49837);
or UO_163 (O_163,N_49927,N_49751);
nor UO_164 (O_164,N_49801,N_49773);
xor UO_165 (O_165,N_49890,N_49879);
or UO_166 (O_166,N_49918,N_49805);
or UO_167 (O_167,N_49786,N_49758);
nand UO_168 (O_168,N_49937,N_49814);
and UO_169 (O_169,N_49973,N_49956);
nor UO_170 (O_170,N_49934,N_49981);
and UO_171 (O_171,N_49858,N_49841);
xnor UO_172 (O_172,N_49880,N_49800);
and UO_173 (O_173,N_49973,N_49923);
or UO_174 (O_174,N_49914,N_49889);
xor UO_175 (O_175,N_49909,N_49832);
nand UO_176 (O_176,N_49793,N_49778);
xor UO_177 (O_177,N_49843,N_49981);
nand UO_178 (O_178,N_49850,N_49928);
xnor UO_179 (O_179,N_49914,N_49882);
or UO_180 (O_180,N_49838,N_49907);
nor UO_181 (O_181,N_49854,N_49969);
and UO_182 (O_182,N_49815,N_49951);
nor UO_183 (O_183,N_49801,N_49907);
nand UO_184 (O_184,N_49801,N_49812);
nand UO_185 (O_185,N_49795,N_49875);
nand UO_186 (O_186,N_49897,N_49777);
and UO_187 (O_187,N_49852,N_49968);
or UO_188 (O_188,N_49773,N_49795);
nor UO_189 (O_189,N_49944,N_49796);
nor UO_190 (O_190,N_49821,N_49903);
and UO_191 (O_191,N_49796,N_49904);
nand UO_192 (O_192,N_49954,N_49832);
nor UO_193 (O_193,N_49880,N_49913);
or UO_194 (O_194,N_49969,N_49750);
or UO_195 (O_195,N_49902,N_49765);
and UO_196 (O_196,N_49924,N_49921);
nand UO_197 (O_197,N_49765,N_49804);
or UO_198 (O_198,N_49889,N_49942);
and UO_199 (O_199,N_49794,N_49985);
xnor UO_200 (O_200,N_49999,N_49779);
xnor UO_201 (O_201,N_49845,N_49925);
xor UO_202 (O_202,N_49970,N_49864);
or UO_203 (O_203,N_49806,N_49994);
nor UO_204 (O_204,N_49964,N_49938);
nand UO_205 (O_205,N_49840,N_49753);
nor UO_206 (O_206,N_49797,N_49963);
nor UO_207 (O_207,N_49991,N_49920);
nand UO_208 (O_208,N_49817,N_49885);
nor UO_209 (O_209,N_49992,N_49793);
and UO_210 (O_210,N_49946,N_49913);
nor UO_211 (O_211,N_49974,N_49971);
or UO_212 (O_212,N_49914,N_49843);
and UO_213 (O_213,N_49851,N_49892);
or UO_214 (O_214,N_49952,N_49867);
and UO_215 (O_215,N_49955,N_49989);
or UO_216 (O_216,N_49825,N_49765);
and UO_217 (O_217,N_49922,N_49988);
xnor UO_218 (O_218,N_49844,N_49916);
nand UO_219 (O_219,N_49792,N_49825);
or UO_220 (O_220,N_49965,N_49824);
and UO_221 (O_221,N_49765,N_49958);
nand UO_222 (O_222,N_49929,N_49756);
or UO_223 (O_223,N_49972,N_49880);
or UO_224 (O_224,N_49900,N_49932);
xor UO_225 (O_225,N_49978,N_49849);
nand UO_226 (O_226,N_49787,N_49760);
and UO_227 (O_227,N_49846,N_49801);
nand UO_228 (O_228,N_49777,N_49903);
nand UO_229 (O_229,N_49906,N_49957);
xor UO_230 (O_230,N_49952,N_49871);
xnor UO_231 (O_231,N_49899,N_49831);
or UO_232 (O_232,N_49787,N_49907);
and UO_233 (O_233,N_49754,N_49886);
nand UO_234 (O_234,N_49944,N_49770);
xor UO_235 (O_235,N_49790,N_49967);
nand UO_236 (O_236,N_49762,N_49915);
and UO_237 (O_237,N_49916,N_49848);
nand UO_238 (O_238,N_49971,N_49832);
nor UO_239 (O_239,N_49957,N_49895);
and UO_240 (O_240,N_49789,N_49775);
xnor UO_241 (O_241,N_49918,N_49843);
or UO_242 (O_242,N_49911,N_49814);
and UO_243 (O_243,N_49857,N_49755);
and UO_244 (O_244,N_49846,N_49862);
or UO_245 (O_245,N_49967,N_49831);
nor UO_246 (O_246,N_49869,N_49761);
xnor UO_247 (O_247,N_49949,N_49951);
nand UO_248 (O_248,N_49792,N_49790);
and UO_249 (O_249,N_49832,N_49836);
xnor UO_250 (O_250,N_49942,N_49832);
nor UO_251 (O_251,N_49869,N_49931);
xnor UO_252 (O_252,N_49993,N_49955);
or UO_253 (O_253,N_49864,N_49765);
nand UO_254 (O_254,N_49755,N_49833);
xnor UO_255 (O_255,N_49894,N_49769);
xor UO_256 (O_256,N_49899,N_49825);
xnor UO_257 (O_257,N_49957,N_49841);
nor UO_258 (O_258,N_49950,N_49931);
and UO_259 (O_259,N_49853,N_49838);
or UO_260 (O_260,N_49945,N_49911);
xnor UO_261 (O_261,N_49910,N_49895);
xnor UO_262 (O_262,N_49947,N_49852);
nor UO_263 (O_263,N_49765,N_49900);
and UO_264 (O_264,N_49758,N_49959);
xor UO_265 (O_265,N_49840,N_49755);
nor UO_266 (O_266,N_49761,N_49801);
or UO_267 (O_267,N_49758,N_49890);
and UO_268 (O_268,N_49767,N_49964);
nor UO_269 (O_269,N_49799,N_49891);
nand UO_270 (O_270,N_49867,N_49811);
and UO_271 (O_271,N_49972,N_49799);
nand UO_272 (O_272,N_49856,N_49858);
xor UO_273 (O_273,N_49809,N_49908);
and UO_274 (O_274,N_49895,N_49822);
and UO_275 (O_275,N_49832,N_49899);
or UO_276 (O_276,N_49918,N_49974);
xnor UO_277 (O_277,N_49951,N_49820);
xor UO_278 (O_278,N_49976,N_49755);
or UO_279 (O_279,N_49837,N_49999);
nand UO_280 (O_280,N_49778,N_49978);
or UO_281 (O_281,N_49859,N_49933);
nor UO_282 (O_282,N_49827,N_49925);
or UO_283 (O_283,N_49821,N_49768);
or UO_284 (O_284,N_49761,N_49954);
or UO_285 (O_285,N_49770,N_49902);
nor UO_286 (O_286,N_49867,N_49762);
and UO_287 (O_287,N_49796,N_49752);
or UO_288 (O_288,N_49962,N_49983);
nand UO_289 (O_289,N_49831,N_49881);
xor UO_290 (O_290,N_49804,N_49919);
or UO_291 (O_291,N_49955,N_49908);
or UO_292 (O_292,N_49984,N_49823);
and UO_293 (O_293,N_49944,N_49858);
xnor UO_294 (O_294,N_49824,N_49964);
xnor UO_295 (O_295,N_49857,N_49939);
and UO_296 (O_296,N_49762,N_49871);
xnor UO_297 (O_297,N_49809,N_49853);
nand UO_298 (O_298,N_49933,N_49794);
or UO_299 (O_299,N_49886,N_49955);
and UO_300 (O_300,N_49808,N_49885);
xor UO_301 (O_301,N_49770,N_49941);
nand UO_302 (O_302,N_49908,N_49976);
or UO_303 (O_303,N_49992,N_49809);
nor UO_304 (O_304,N_49753,N_49812);
nand UO_305 (O_305,N_49973,N_49821);
nor UO_306 (O_306,N_49856,N_49826);
and UO_307 (O_307,N_49920,N_49921);
nand UO_308 (O_308,N_49798,N_49877);
nand UO_309 (O_309,N_49762,N_49887);
nor UO_310 (O_310,N_49932,N_49972);
and UO_311 (O_311,N_49955,N_49761);
xnor UO_312 (O_312,N_49780,N_49977);
xor UO_313 (O_313,N_49935,N_49840);
or UO_314 (O_314,N_49962,N_49844);
or UO_315 (O_315,N_49989,N_49915);
or UO_316 (O_316,N_49802,N_49933);
xor UO_317 (O_317,N_49870,N_49774);
and UO_318 (O_318,N_49825,N_49943);
xnor UO_319 (O_319,N_49890,N_49969);
nand UO_320 (O_320,N_49915,N_49751);
nand UO_321 (O_321,N_49889,N_49946);
nand UO_322 (O_322,N_49821,N_49850);
or UO_323 (O_323,N_49768,N_49875);
xnor UO_324 (O_324,N_49986,N_49833);
or UO_325 (O_325,N_49793,N_49957);
or UO_326 (O_326,N_49808,N_49907);
nor UO_327 (O_327,N_49849,N_49835);
or UO_328 (O_328,N_49905,N_49771);
nand UO_329 (O_329,N_49827,N_49765);
nor UO_330 (O_330,N_49976,N_49786);
and UO_331 (O_331,N_49828,N_49892);
and UO_332 (O_332,N_49825,N_49770);
xnor UO_333 (O_333,N_49937,N_49819);
or UO_334 (O_334,N_49774,N_49960);
or UO_335 (O_335,N_49891,N_49923);
and UO_336 (O_336,N_49901,N_49972);
nand UO_337 (O_337,N_49755,N_49979);
nand UO_338 (O_338,N_49917,N_49900);
nor UO_339 (O_339,N_49991,N_49827);
nor UO_340 (O_340,N_49902,N_49976);
xor UO_341 (O_341,N_49852,N_49905);
nor UO_342 (O_342,N_49849,N_49932);
or UO_343 (O_343,N_49770,N_49923);
or UO_344 (O_344,N_49935,N_49850);
nor UO_345 (O_345,N_49955,N_49921);
or UO_346 (O_346,N_49876,N_49975);
nand UO_347 (O_347,N_49969,N_49928);
xnor UO_348 (O_348,N_49893,N_49940);
nor UO_349 (O_349,N_49949,N_49937);
and UO_350 (O_350,N_49801,N_49854);
nand UO_351 (O_351,N_49955,N_49944);
xnor UO_352 (O_352,N_49880,N_49873);
nand UO_353 (O_353,N_49899,N_49751);
and UO_354 (O_354,N_49771,N_49847);
xnor UO_355 (O_355,N_49777,N_49992);
nor UO_356 (O_356,N_49797,N_49800);
xor UO_357 (O_357,N_49974,N_49885);
xnor UO_358 (O_358,N_49769,N_49933);
or UO_359 (O_359,N_49978,N_49892);
and UO_360 (O_360,N_49954,N_49874);
and UO_361 (O_361,N_49964,N_49855);
nand UO_362 (O_362,N_49903,N_49761);
and UO_363 (O_363,N_49772,N_49846);
xor UO_364 (O_364,N_49997,N_49965);
nor UO_365 (O_365,N_49963,N_49970);
xnor UO_366 (O_366,N_49965,N_49809);
xnor UO_367 (O_367,N_49873,N_49987);
nor UO_368 (O_368,N_49920,N_49807);
nor UO_369 (O_369,N_49959,N_49997);
xnor UO_370 (O_370,N_49861,N_49960);
xnor UO_371 (O_371,N_49893,N_49788);
nor UO_372 (O_372,N_49858,N_49754);
and UO_373 (O_373,N_49802,N_49994);
or UO_374 (O_374,N_49945,N_49782);
or UO_375 (O_375,N_49862,N_49886);
or UO_376 (O_376,N_49966,N_49894);
or UO_377 (O_377,N_49939,N_49782);
nor UO_378 (O_378,N_49885,N_49884);
and UO_379 (O_379,N_49990,N_49837);
or UO_380 (O_380,N_49750,N_49779);
or UO_381 (O_381,N_49929,N_49779);
and UO_382 (O_382,N_49991,N_49768);
nor UO_383 (O_383,N_49909,N_49878);
xnor UO_384 (O_384,N_49766,N_49906);
and UO_385 (O_385,N_49854,N_49830);
nand UO_386 (O_386,N_49789,N_49903);
nand UO_387 (O_387,N_49963,N_49813);
and UO_388 (O_388,N_49878,N_49898);
nand UO_389 (O_389,N_49782,N_49845);
nand UO_390 (O_390,N_49800,N_49911);
nand UO_391 (O_391,N_49778,N_49806);
nor UO_392 (O_392,N_49929,N_49863);
nand UO_393 (O_393,N_49884,N_49813);
nor UO_394 (O_394,N_49760,N_49955);
or UO_395 (O_395,N_49856,N_49999);
xor UO_396 (O_396,N_49969,N_49829);
or UO_397 (O_397,N_49918,N_49921);
xor UO_398 (O_398,N_49985,N_49966);
nand UO_399 (O_399,N_49838,N_49904);
nor UO_400 (O_400,N_49782,N_49907);
nand UO_401 (O_401,N_49777,N_49913);
nand UO_402 (O_402,N_49931,N_49777);
or UO_403 (O_403,N_49937,N_49932);
and UO_404 (O_404,N_49757,N_49942);
xor UO_405 (O_405,N_49841,N_49755);
nand UO_406 (O_406,N_49868,N_49917);
nor UO_407 (O_407,N_49777,N_49809);
xnor UO_408 (O_408,N_49920,N_49851);
nand UO_409 (O_409,N_49915,N_49966);
and UO_410 (O_410,N_49815,N_49968);
nand UO_411 (O_411,N_49887,N_49820);
and UO_412 (O_412,N_49790,N_49753);
or UO_413 (O_413,N_49818,N_49897);
and UO_414 (O_414,N_49822,N_49987);
xnor UO_415 (O_415,N_49876,N_49902);
nor UO_416 (O_416,N_49844,N_49832);
or UO_417 (O_417,N_49926,N_49890);
and UO_418 (O_418,N_49841,N_49770);
xor UO_419 (O_419,N_49858,N_49778);
nand UO_420 (O_420,N_49852,N_49932);
nand UO_421 (O_421,N_49803,N_49915);
or UO_422 (O_422,N_49995,N_49846);
and UO_423 (O_423,N_49877,N_49937);
nor UO_424 (O_424,N_49932,N_49778);
or UO_425 (O_425,N_49789,N_49871);
or UO_426 (O_426,N_49911,N_49903);
xor UO_427 (O_427,N_49796,N_49998);
nor UO_428 (O_428,N_49772,N_49834);
nor UO_429 (O_429,N_49896,N_49923);
nor UO_430 (O_430,N_49879,N_49909);
and UO_431 (O_431,N_49755,N_49860);
nand UO_432 (O_432,N_49756,N_49857);
or UO_433 (O_433,N_49966,N_49831);
or UO_434 (O_434,N_49800,N_49764);
nand UO_435 (O_435,N_49797,N_49973);
xor UO_436 (O_436,N_49774,N_49781);
or UO_437 (O_437,N_49880,N_49754);
or UO_438 (O_438,N_49961,N_49990);
or UO_439 (O_439,N_49942,N_49950);
or UO_440 (O_440,N_49880,N_49916);
nand UO_441 (O_441,N_49788,N_49780);
and UO_442 (O_442,N_49855,N_49873);
xnor UO_443 (O_443,N_49977,N_49773);
xor UO_444 (O_444,N_49895,N_49939);
and UO_445 (O_445,N_49964,N_49801);
or UO_446 (O_446,N_49764,N_49796);
and UO_447 (O_447,N_49839,N_49820);
nand UO_448 (O_448,N_49888,N_49980);
and UO_449 (O_449,N_49919,N_49987);
nand UO_450 (O_450,N_49838,N_49770);
xor UO_451 (O_451,N_49963,N_49883);
nand UO_452 (O_452,N_49863,N_49945);
xor UO_453 (O_453,N_49986,N_49893);
nand UO_454 (O_454,N_49799,N_49826);
nand UO_455 (O_455,N_49804,N_49898);
or UO_456 (O_456,N_49809,N_49882);
nand UO_457 (O_457,N_49913,N_49766);
xor UO_458 (O_458,N_49762,N_49939);
or UO_459 (O_459,N_49782,N_49813);
xor UO_460 (O_460,N_49859,N_49754);
nor UO_461 (O_461,N_49753,N_49943);
or UO_462 (O_462,N_49821,N_49757);
or UO_463 (O_463,N_49808,N_49752);
or UO_464 (O_464,N_49884,N_49868);
and UO_465 (O_465,N_49784,N_49863);
nand UO_466 (O_466,N_49802,N_49824);
nand UO_467 (O_467,N_49758,N_49987);
xor UO_468 (O_468,N_49906,N_49810);
nor UO_469 (O_469,N_49958,N_49964);
and UO_470 (O_470,N_49807,N_49830);
or UO_471 (O_471,N_49958,N_49922);
nor UO_472 (O_472,N_49831,N_49806);
xnor UO_473 (O_473,N_49948,N_49795);
and UO_474 (O_474,N_49836,N_49858);
or UO_475 (O_475,N_49854,N_49908);
xnor UO_476 (O_476,N_49750,N_49909);
or UO_477 (O_477,N_49967,N_49945);
nor UO_478 (O_478,N_49752,N_49972);
nor UO_479 (O_479,N_49984,N_49849);
xnor UO_480 (O_480,N_49825,N_49932);
xnor UO_481 (O_481,N_49791,N_49931);
nor UO_482 (O_482,N_49908,N_49775);
and UO_483 (O_483,N_49784,N_49831);
nor UO_484 (O_484,N_49781,N_49855);
or UO_485 (O_485,N_49812,N_49975);
and UO_486 (O_486,N_49959,N_49788);
and UO_487 (O_487,N_49893,N_49914);
xnor UO_488 (O_488,N_49943,N_49973);
xor UO_489 (O_489,N_49993,N_49757);
nand UO_490 (O_490,N_49824,N_49768);
xor UO_491 (O_491,N_49854,N_49941);
xor UO_492 (O_492,N_49978,N_49855);
nor UO_493 (O_493,N_49906,N_49856);
and UO_494 (O_494,N_49754,N_49785);
or UO_495 (O_495,N_49874,N_49970);
and UO_496 (O_496,N_49821,N_49946);
nand UO_497 (O_497,N_49896,N_49849);
or UO_498 (O_498,N_49813,N_49868);
xnor UO_499 (O_499,N_49756,N_49773);
xor UO_500 (O_500,N_49878,N_49955);
and UO_501 (O_501,N_49753,N_49820);
nor UO_502 (O_502,N_49909,N_49969);
nand UO_503 (O_503,N_49782,N_49859);
nor UO_504 (O_504,N_49818,N_49951);
nand UO_505 (O_505,N_49997,N_49870);
nor UO_506 (O_506,N_49959,N_49933);
and UO_507 (O_507,N_49806,N_49779);
xor UO_508 (O_508,N_49888,N_49772);
and UO_509 (O_509,N_49835,N_49974);
xor UO_510 (O_510,N_49905,N_49846);
or UO_511 (O_511,N_49873,N_49928);
nand UO_512 (O_512,N_49877,N_49971);
or UO_513 (O_513,N_49957,N_49932);
or UO_514 (O_514,N_49851,N_49865);
or UO_515 (O_515,N_49918,N_49801);
and UO_516 (O_516,N_49975,N_49843);
or UO_517 (O_517,N_49888,N_49896);
and UO_518 (O_518,N_49758,N_49914);
or UO_519 (O_519,N_49986,N_49926);
nand UO_520 (O_520,N_49854,N_49860);
nand UO_521 (O_521,N_49907,N_49803);
nor UO_522 (O_522,N_49908,N_49769);
and UO_523 (O_523,N_49945,N_49807);
xnor UO_524 (O_524,N_49999,N_49835);
nand UO_525 (O_525,N_49796,N_49833);
and UO_526 (O_526,N_49854,N_49880);
xnor UO_527 (O_527,N_49769,N_49831);
or UO_528 (O_528,N_49967,N_49920);
and UO_529 (O_529,N_49939,N_49768);
nand UO_530 (O_530,N_49946,N_49866);
nand UO_531 (O_531,N_49944,N_49886);
xnor UO_532 (O_532,N_49973,N_49773);
xnor UO_533 (O_533,N_49883,N_49828);
xor UO_534 (O_534,N_49996,N_49889);
or UO_535 (O_535,N_49922,N_49938);
and UO_536 (O_536,N_49790,N_49974);
nand UO_537 (O_537,N_49833,N_49985);
nand UO_538 (O_538,N_49967,N_49821);
xor UO_539 (O_539,N_49956,N_49954);
nand UO_540 (O_540,N_49854,N_49815);
xnor UO_541 (O_541,N_49825,N_49865);
and UO_542 (O_542,N_49987,N_49907);
nor UO_543 (O_543,N_49844,N_49923);
xnor UO_544 (O_544,N_49967,N_49980);
nand UO_545 (O_545,N_49831,N_49906);
nand UO_546 (O_546,N_49789,N_49999);
xnor UO_547 (O_547,N_49758,N_49927);
nand UO_548 (O_548,N_49775,N_49895);
nor UO_549 (O_549,N_49969,N_49761);
nor UO_550 (O_550,N_49839,N_49966);
nand UO_551 (O_551,N_49767,N_49983);
or UO_552 (O_552,N_49938,N_49801);
xnor UO_553 (O_553,N_49876,N_49814);
nor UO_554 (O_554,N_49912,N_49889);
nor UO_555 (O_555,N_49995,N_49812);
nor UO_556 (O_556,N_49826,N_49911);
xnor UO_557 (O_557,N_49957,N_49836);
nor UO_558 (O_558,N_49844,N_49824);
or UO_559 (O_559,N_49847,N_49888);
or UO_560 (O_560,N_49826,N_49959);
and UO_561 (O_561,N_49777,N_49794);
or UO_562 (O_562,N_49851,N_49825);
or UO_563 (O_563,N_49898,N_49858);
or UO_564 (O_564,N_49773,N_49888);
nand UO_565 (O_565,N_49875,N_49805);
and UO_566 (O_566,N_49802,N_49942);
or UO_567 (O_567,N_49817,N_49947);
xor UO_568 (O_568,N_49972,N_49971);
nor UO_569 (O_569,N_49759,N_49917);
xnor UO_570 (O_570,N_49927,N_49785);
nor UO_571 (O_571,N_49855,N_49989);
xor UO_572 (O_572,N_49910,N_49867);
or UO_573 (O_573,N_49959,N_49767);
or UO_574 (O_574,N_49918,N_49965);
nor UO_575 (O_575,N_49940,N_49766);
nor UO_576 (O_576,N_49831,N_49888);
xor UO_577 (O_577,N_49753,N_49819);
nor UO_578 (O_578,N_49827,N_49804);
and UO_579 (O_579,N_49893,N_49795);
or UO_580 (O_580,N_49910,N_49773);
nor UO_581 (O_581,N_49816,N_49875);
nand UO_582 (O_582,N_49767,N_49873);
nor UO_583 (O_583,N_49834,N_49953);
xor UO_584 (O_584,N_49833,N_49801);
nor UO_585 (O_585,N_49753,N_49940);
xor UO_586 (O_586,N_49783,N_49961);
or UO_587 (O_587,N_49920,N_49802);
nor UO_588 (O_588,N_49938,N_49850);
nor UO_589 (O_589,N_49956,N_49939);
xnor UO_590 (O_590,N_49828,N_49777);
and UO_591 (O_591,N_49767,N_49984);
nor UO_592 (O_592,N_49864,N_49771);
nor UO_593 (O_593,N_49985,N_49953);
xor UO_594 (O_594,N_49861,N_49920);
nor UO_595 (O_595,N_49995,N_49839);
and UO_596 (O_596,N_49880,N_49926);
nor UO_597 (O_597,N_49825,N_49832);
nand UO_598 (O_598,N_49785,N_49867);
or UO_599 (O_599,N_49773,N_49884);
and UO_600 (O_600,N_49962,N_49992);
or UO_601 (O_601,N_49993,N_49766);
xor UO_602 (O_602,N_49884,N_49798);
nor UO_603 (O_603,N_49768,N_49861);
nor UO_604 (O_604,N_49759,N_49914);
and UO_605 (O_605,N_49784,N_49920);
or UO_606 (O_606,N_49772,N_49985);
or UO_607 (O_607,N_49838,N_49965);
nor UO_608 (O_608,N_49873,N_49936);
xor UO_609 (O_609,N_49961,N_49788);
or UO_610 (O_610,N_49805,N_49831);
or UO_611 (O_611,N_49900,N_49827);
xor UO_612 (O_612,N_49828,N_49907);
or UO_613 (O_613,N_49885,N_49861);
nor UO_614 (O_614,N_49769,N_49989);
and UO_615 (O_615,N_49967,N_49808);
nand UO_616 (O_616,N_49937,N_49817);
or UO_617 (O_617,N_49964,N_49930);
or UO_618 (O_618,N_49995,N_49955);
xnor UO_619 (O_619,N_49788,N_49771);
xor UO_620 (O_620,N_49968,N_49767);
or UO_621 (O_621,N_49750,N_49828);
nor UO_622 (O_622,N_49826,N_49925);
xnor UO_623 (O_623,N_49980,N_49890);
or UO_624 (O_624,N_49937,N_49927);
or UO_625 (O_625,N_49999,N_49772);
or UO_626 (O_626,N_49928,N_49764);
nand UO_627 (O_627,N_49904,N_49864);
nand UO_628 (O_628,N_49756,N_49779);
nor UO_629 (O_629,N_49858,N_49873);
nand UO_630 (O_630,N_49995,N_49931);
nand UO_631 (O_631,N_49870,N_49962);
xor UO_632 (O_632,N_49966,N_49760);
nand UO_633 (O_633,N_49844,N_49764);
and UO_634 (O_634,N_49840,N_49867);
and UO_635 (O_635,N_49869,N_49815);
nand UO_636 (O_636,N_49952,N_49767);
nand UO_637 (O_637,N_49902,N_49960);
nand UO_638 (O_638,N_49805,N_49842);
or UO_639 (O_639,N_49961,N_49897);
xnor UO_640 (O_640,N_49802,N_49898);
or UO_641 (O_641,N_49990,N_49777);
and UO_642 (O_642,N_49893,N_49813);
nand UO_643 (O_643,N_49945,N_49763);
or UO_644 (O_644,N_49802,N_49879);
nor UO_645 (O_645,N_49830,N_49923);
nor UO_646 (O_646,N_49980,N_49763);
or UO_647 (O_647,N_49985,N_49919);
xor UO_648 (O_648,N_49794,N_49813);
xnor UO_649 (O_649,N_49792,N_49937);
nand UO_650 (O_650,N_49969,N_49795);
nor UO_651 (O_651,N_49921,N_49911);
or UO_652 (O_652,N_49936,N_49937);
nor UO_653 (O_653,N_49943,N_49804);
xnor UO_654 (O_654,N_49891,N_49939);
xnor UO_655 (O_655,N_49835,N_49799);
or UO_656 (O_656,N_49803,N_49791);
nor UO_657 (O_657,N_49791,N_49883);
nand UO_658 (O_658,N_49968,N_49869);
nor UO_659 (O_659,N_49934,N_49889);
xor UO_660 (O_660,N_49894,N_49960);
nand UO_661 (O_661,N_49894,N_49759);
nor UO_662 (O_662,N_49857,N_49820);
xnor UO_663 (O_663,N_49895,N_49835);
and UO_664 (O_664,N_49756,N_49941);
xnor UO_665 (O_665,N_49969,N_49929);
or UO_666 (O_666,N_49897,N_49753);
or UO_667 (O_667,N_49939,N_49853);
nor UO_668 (O_668,N_49888,N_49956);
or UO_669 (O_669,N_49812,N_49977);
and UO_670 (O_670,N_49763,N_49982);
nor UO_671 (O_671,N_49832,N_49990);
nand UO_672 (O_672,N_49924,N_49875);
or UO_673 (O_673,N_49815,N_49875);
or UO_674 (O_674,N_49981,N_49897);
nand UO_675 (O_675,N_49795,N_49894);
or UO_676 (O_676,N_49839,N_49913);
nor UO_677 (O_677,N_49982,N_49785);
or UO_678 (O_678,N_49895,N_49857);
xor UO_679 (O_679,N_49975,N_49964);
xnor UO_680 (O_680,N_49839,N_49815);
nor UO_681 (O_681,N_49888,N_49862);
xnor UO_682 (O_682,N_49853,N_49931);
and UO_683 (O_683,N_49811,N_49957);
or UO_684 (O_684,N_49790,N_49868);
xor UO_685 (O_685,N_49900,N_49792);
nor UO_686 (O_686,N_49953,N_49771);
nand UO_687 (O_687,N_49846,N_49861);
nor UO_688 (O_688,N_49999,N_49840);
and UO_689 (O_689,N_49847,N_49993);
and UO_690 (O_690,N_49765,N_49848);
or UO_691 (O_691,N_49922,N_49862);
nand UO_692 (O_692,N_49927,N_49842);
and UO_693 (O_693,N_49911,N_49986);
or UO_694 (O_694,N_49905,N_49770);
xor UO_695 (O_695,N_49900,N_49960);
nor UO_696 (O_696,N_49957,N_49825);
and UO_697 (O_697,N_49808,N_49923);
xnor UO_698 (O_698,N_49869,N_49752);
xnor UO_699 (O_699,N_49778,N_49777);
nor UO_700 (O_700,N_49923,N_49956);
xnor UO_701 (O_701,N_49893,N_49882);
and UO_702 (O_702,N_49958,N_49769);
nor UO_703 (O_703,N_49838,N_49852);
xnor UO_704 (O_704,N_49863,N_49861);
nand UO_705 (O_705,N_49766,N_49850);
and UO_706 (O_706,N_49881,N_49781);
xnor UO_707 (O_707,N_49839,N_49925);
nor UO_708 (O_708,N_49779,N_49876);
nand UO_709 (O_709,N_49972,N_49920);
or UO_710 (O_710,N_49989,N_49898);
nand UO_711 (O_711,N_49962,N_49856);
xor UO_712 (O_712,N_49757,N_49923);
xor UO_713 (O_713,N_49909,N_49761);
or UO_714 (O_714,N_49869,N_49864);
or UO_715 (O_715,N_49944,N_49843);
and UO_716 (O_716,N_49806,N_49932);
nor UO_717 (O_717,N_49772,N_49791);
nand UO_718 (O_718,N_49846,N_49850);
nand UO_719 (O_719,N_49857,N_49995);
and UO_720 (O_720,N_49868,N_49883);
xnor UO_721 (O_721,N_49966,N_49936);
or UO_722 (O_722,N_49954,N_49911);
nand UO_723 (O_723,N_49754,N_49901);
xor UO_724 (O_724,N_49980,N_49954);
nand UO_725 (O_725,N_49916,N_49902);
nand UO_726 (O_726,N_49824,N_49987);
or UO_727 (O_727,N_49791,N_49879);
and UO_728 (O_728,N_49927,N_49852);
and UO_729 (O_729,N_49863,N_49956);
nor UO_730 (O_730,N_49809,N_49986);
nand UO_731 (O_731,N_49765,N_49935);
nor UO_732 (O_732,N_49752,N_49971);
nor UO_733 (O_733,N_49779,N_49990);
nand UO_734 (O_734,N_49868,N_49801);
xnor UO_735 (O_735,N_49754,N_49998);
nand UO_736 (O_736,N_49851,N_49797);
nand UO_737 (O_737,N_49972,N_49982);
or UO_738 (O_738,N_49945,N_49985);
nor UO_739 (O_739,N_49800,N_49882);
or UO_740 (O_740,N_49866,N_49805);
nor UO_741 (O_741,N_49980,N_49767);
nand UO_742 (O_742,N_49810,N_49919);
and UO_743 (O_743,N_49821,N_49753);
nor UO_744 (O_744,N_49765,N_49845);
xnor UO_745 (O_745,N_49861,N_49915);
and UO_746 (O_746,N_49993,N_49856);
and UO_747 (O_747,N_49947,N_49851);
nor UO_748 (O_748,N_49802,N_49860);
and UO_749 (O_749,N_49801,N_49988);
or UO_750 (O_750,N_49862,N_49867);
nor UO_751 (O_751,N_49992,N_49833);
nand UO_752 (O_752,N_49838,N_49861);
nand UO_753 (O_753,N_49769,N_49925);
or UO_754 (O_754,N_49773,N_49893);
xnor UO_755 (O_755,N_49986,N_49920);
nand UO_756 (O_756,N_49836,N_49797);
nand UO_757 (O_757,N_49853,N_49850);
nor UO_758 (O_758,N_49810,N_49875);
or UO_759 (O_759,N_49949,N_49821);
nand UO_760 (O_760,N_49806,N_49889);
xnor UO_761 (O_761,N_49921,N_49865);
nor UO_762 (O_762,N_49771,N_49997);
and UO_763 (O_763,N_49871,N_49863);
xnor UO_764 (O_764,N_49922,N_49802);
and UO_765 (O_765,N_49919,N_49833);
and UO_766 (O_766,N_49755,N_49891);
and UO_767 (O_767,N_49973,N_49767);
nor UO_768 (O_768,N_49778,N_49980);
and UO_769 (O_769,N_49995,N_49921);
nand UO_770 (O_770,N_49868,N_49788);
nand UO_771 (O_771,N_49797,N_49983);
and UO_772 (O_772,N_49765,N_49830);
xor UO_773 (O_773,N_49918,N_49913);
xor UO_774 (O_774,N_49805,N_49949);
or UO_775 (O_775,N_49866,N_49787);
or UO_776 (O_776,N_49815,N_49781);
and UO_777 (O_777,N_49755,N_49988);
xor UO_778 (O_778,N_49976,N_49817);
and UO_779 (O_779,N_49891,N_49915);
xnor UO_780 (O_780,N_49801,N_49862);
and UO_781 (O_781,N_49801,N_49957);
or UO_782 (O_782,N_49882,N_49947);
and UO_783 (O_783,N_49801,N_49879);
and UO_784 (O_784,N_49969,N_49965);
xnor UO_785 (O_785,N_49770,N_49751);
xor UO_786 (O_786,N_49804,N_49986);
nor UO_787 (O_787,N_49927,N_49990);
nand UO_788 (O_788,N_49766,N_49754);
nand UO_789 (O_789,N_49884,N_49888);
or UO_790 (O_790,N_49948,N_49895);
or UO_791 (O_791,N_49851,N_49857);
xnor UO_792 (O_792,N_49812,N_49998);
xnor UO_793 (O_793,N_49803,N_49763);
nor UO_794 (O_794,N_49824,N_49870);
and UO_795 (O_795,N_49755,N_49998);
xor UO_796 (O_796,N_49840,N_49926);
nor UO_797 (O_797,N_49940,N_49985);
xnor UO_798 (O_798,N_49798,N_49925);
or UO_799 (O_799,N_49948,N_49790);
xnor UO_800 (O_800,N_49902,N_49872);
nor UO_801 (O_801,N_49844,N_49855);
nand UO_802 (O_802,N_49853,N_49772);
nand UO_803 (O_803,N_49871,N_49810);
nand UO_804 (O_804,N_49969,N_49783);
xor UO_805 (O_805,N_49872,N_49955);
nor UO_806 (O_806,N_49983,N_49857);
and UO_807 (O_807,N_49945,N_49914);
nand UO_808 (O_808,N_49782,N_49896);
xnor UO_809 (O_809,N_49781,N_49810);
and UO_810 (O_810,N_49919,N_49803);
nor UO_811 (O_811,N_49922,N_49796);
and UO_812 (O_812,N_49762,N_49849);
or UO_813 (O_813,N_49870,N_49814);
or UO_814 (O_814,N_49912,N_49779);
and UO_815 (O_815,N_49928,N_49816);
and UO_816 (O_816,N_49884,N_49980);
xnor UO_817 (O_817,N_49970,N_49771);
nor UO_818 (O_818,N_49941,N_49908);
xor UO_819 (O_819,N_49909,N_49966);
and UO_820 (O_820,N_49913,N_49770);
or UO_821 (O_821,N_49876,N_49911);
nand UO_822 (O_822,N_49790,N_49926);
nand UO_823 (O_823,N_49898,N_49880);
nor UO_824 (O_824,N_49966,N_49762);
nand UO_825 (O_825,N_49765,N_49829);
xnor UO_826 (O_826,N_49940,N_49975);
nand UO_827 (O_827,N_49909,N_49949);
xor UO_828 (O_828,N_49826,N_49809);
nor UO_829 (O_829,N_49818,N_49975);
xnor UO_830 (O_830,N_49934,N_49762);
nand UO_831 (O_831,N_49847,N_49778);
or UO_832 (O_832,N_49846,N_49879);
nor UO_833 (O_833,N_49970,N_49959);
xor UO_834 (O_834,N_49785,N_49883);
and UO_835 (O_835,N_49924,N_49974);
or UO_836 (O_836,N_49903,N_49926);
xnor UO_837 (O_837,N_49956,N_49756);
or UO_838 (O_838,N_49855,N_49758);
or UO_839 (O_839,N_49925,N_49776);
nor UO_840 (O_840,N_49928,N_49808);
xnor UO_841 (O_841,N_49764,N_49761);
nor UO_842 (O_842,N_49784,N_49854);
or UO_843 (O_843,N_49831,N_49882);
xnor UO_844 (O_844,N_49887,N_49814);
and UO_845 (O_845,N_49926,N_49866);
nor UO_846 (O_846,N_49955,N_49991);
and UO_847 (O_847,N_49878,N_49779);
and UO_848 (O_848,N_49761,N_49994);
xnor UO_849 (O_849,N_49781,N_49769);
and UO_850 (O_850,N_49985,N_49751);
nor UO_851 (O_851,N_49835,N_49936);
and UO_852 (O_852,N_49811,N_49949);
or UO_853 (O_853,N_49821,N_49882);
nor UO_854 (O_854,N_49750,N_49992);
nand UO_855 (O_855,N_49760,N_49815);
xor UO_856 (O_856,N_49811,N_49926);
xor UO_857 (O_857,N_49858,N_49875);
and UO_858 (O_858,N_49945,N_49759);
and UO_859 (O_859,N_49834,N_49935);
or UO_860 (O_860,N_49774,N_49933);
nand UO_861 (O_861,N_49999,N_49932);
nor UO_862 (O_862,N_49832,N_49939);
and UO_863 (O_863,N_49797,N_49780);
nor UO_864 (O_864,N_49946,N_49812);
xnor UO_865 (O_865,N_49981,N_49862);
nor UO_866 (O_866,N_49859,N_49993);
and UO_867 (O_867,N_49819,N_49755);
or UO_868 (O_868,N_49892,N_49936);
nand UO_869 (O_869,N_49859,N_49752);
xor UO_870 (O_870,N_49811,N_49985);
and UO_871 (O_871,N_49903,N_49976);
or UO_872 (O_872,N_49921,N_49907);
nor UO_873 (O_873,N_49880,N_49961);
and UO_874 (O_874,N_49804,N_49805);
xnor UO_875 (O_875,N_49787,N_49967);
or UO_876 (O_876,N_49893,N_49835);
and UO_877 (O_877,N_49813,N_49769);
nand UO_878 (O_878,N_49785,N_49897);
nor UO_879 (O_879,N_49772,N_49983);
or UO_880 (O_880,N_49982,N_49910);
or UO_881 (O_881,N_49835,N_49916);
and UO_882 (O_882,N_49842,N_49851);
nor UO_883 (O_883,N_49877,N_49834);
xor UO_884 (O_884,N_49967,N_49960);
or UO_885 (O_885,N_49937,N_49829);
nand UO_886 (O_886,N_49940,N_49778);
nor UO_887 (O_887,N_49954,N_49787);
xnor UO_888 (O_888,N_49986,N_49970);
and UO_889 (O_889,N_49882,N_49994);
and UO_890 (O_890,N_49998,N_49807);
and UO_891 (O_891,N_49794,N_49928);
xor UO_892 (O_892,N_49880,N_49838);
or UO_893 (O_893,N_49885,N_49759);
xor UO_894 (O_894,N_49757,N_49973);
and UO_895 (O_895,N_49851,N_49909);
xor UO_896 (O_896,N_49847,N_49956);
nand UO_897 (O_897,N_49983,N_49888);
xor UO_898 (O_898,N_49899,N_49781);
or UO_899 (O_899,N_49780,N_49898);
xor UO_900 (O_900,N_49950,N_49989);
or UO_901 (O_901,N_49791,N_49932);
nor UO_902 (O_902,N_49812,N_49775);
xnor UO_903 (O_903,N_49847,N_49995);
xor UO_904 (O_904,N_49822,N_49821);
nor UO_905 (O_905,N_49756,N_49863);
nand UO_906 (O_906,N_49808,N_49817);
nor UO_907 (O_907,N_49925,N_49805);
or UO_908 (O_908,N_49888,N_49928);
nor UO_909 (O_909,N_49853,N_49768);
and UO_910 (O_910,N_49801,N_49881);
or UO_911 (O_911,N_49973,N_49905);
or UO_912 (O_912,N_49921,N_49896);
xnor UO_913 (O_913,N_49798,N_49764);
and UO_914 (O_914,N_49815,N_49751);
nor UO_915 (O_915,N_49835,N_49846);
xnor UO_916 (O_916,N_49766,N_49878);
nor UO_917 (O_917,N_49777,N_49792);
nand UO_918 (O_918,N_49851,N_49813);
xor UO_919 (O_919,N_49769,N_49890);
nor UO_920 (O_920,N_49936,N_49926);
nand UO_921 (O_921,N_49862,N_49781);
and UO_922 (O_922,N_49760,N_49798);
nand UO_923 (O_923,N_49784,N_49968);
nor UO_924 (O_924,N_49772,N_49920);
xnor UO_925 (O_925,N_49795,N_49982);
nand UO_926 (O_926,N_49938,N_49815);
nor UO_927 (O_927,N_49963,N_49834);
nor UO_928 (O_928,N_49859,N_49904);
or UO_929 (O_929,N_49902,N_49962);
nand UO_930 (O_930,N_49901,N_49839);
nor UO_931 (O_931,N_49845,N_49915);
xnor UO_932 (O_932,N_49786,N_49797);
or UO_933 (O_933,N_49756,N_49989);
or UO_934 (O_934,N_49890,N_49812);
nand UO_935 (O_935,N_49897,N_49979);
xnor UO_936 (O_936,N_49871,N_49959);
nand UO_937 (O_937,N_49750,N_49768);
nand UO_938 (O_938,N_49983,N_49945);
nand UO_939 (O_939,N_49931,N_49997);
or UO_940 (O_940,N_49995,N_49852);
nor UO_941 (O_941,N_49811,N_49755);
xnor UO_942 (O_942,N_49802,N_49797);
xnor UO_943 (O_943,N_49974,N_49897);
nand UO_944 (O_944,N_49777,N_49799);
and UO_945 (O_945,N_49889,N_49902);
nor UO_946 (O_946,N_49817,N_49952);
nand UO_947 (O_947,N_49828,N_49958);
nor UO_948 (O_948,N_49802,N_49875);
xor UO_949 (O_949,N_49938,N_49770);
nor UO_950 (O_950,N_49963,N_49811);
xor UO_951 (O_951,N_49828,N_49977);
xor UO_952 (O_952,N_49868,N_49806);
nand UO_953 (O_953,N_49899,N_49930);
nor UO_954 (O_954,N_49819,N_49969);
or UO_955 (O_955,N_49904,N_49875);
xor UO_956 (O_956,N_49855,N_49838);
nor UO_957 (O_957,N_49836,N_49802);
nor UO_958 (O_958,N_49938,N_49826);
or UO_959 (O_959,N_49942,N_49846);
nor UO_960 (O_960,N_49934,N_49849);
nand UO_961 (O_961,N_49985,N_49955);
xnor UO_962 (O_962,N_49859,N_49837);
nor UO_963 (O_963,N_49877,N_49904);
xor UO_964 (O_964,N_49812,N_49842);
or UO_965 (O_965,N_49971,N_49766);
xnor UO_966 (O_966,N_49814,N_49776);
nor UO_967 (O_967,N_49904,N_49919);
xor UO_968 (O_968,N_49795,N_49986);
nand UO_969 (O_969,N_49794,N_49981);
xor UO_970 (O_970,N_49939,N_49984);
nor UO_971 (O_971,N_49915,N_49790);
xor UO_972 (O_972,N_49925,N_49754);
or UO_973 (O_973,N_49795,N_49930);
nor UO_974 (O_974,N_49863,N_49873);
and UO_975 (O_975,N_49845,N_49995);
nand UO_976 (O_976,N_49821,N_49783);
nand UO_977 (O_977,N_49939,N_49927);
nor UO_978 (O_978,N_49960,N_49924);
nor UO_979 (O_979,N_49933,N_49922);
or UO_980 (O_980,N_49762,N_49752);
xnor UO_981 (O_981,N_49807,N_49911);
or UO_982 (O_982,N_49996,N_49797);
or UO_983 (O_983,N_49992,N_49857);
xnor UO_984 (O_984,N_49887,N_49819);
or UO_985 (O_985,N_49948,N_49857);
nor UO_986 (O_986,N_49956,N_49850);
nand UO_987 (O_987,N_49953,N_49920);
nor UO_988 (O_988,N_49765,N_49824);
nand UO_989 (O_989,N_49904,N_49773);
and UO_990 (O_990,N_49907,N_49850);
or UO_991 (O_991,N_49908,N_49931);
nand UO_992 (O_992,N_49761,N_49989);
or UO_993 (O_993,N_49812,N_49892);
and UO_994 (O_994,N_49932,N_49912);
xnor UO_995 (O_995,N_49819,N_49825);
or UO_996 (O_996,N_49808,N_49819);
nand UO_997 (O_997,N_49801,N_49844);
xnor UO_998 (O_998,N_49924,N_49797);
nor UO_999 (O_999,N_49906,N_49800);
xnor UO_1000 (O_1000,N_49771,N_49785);
or UO_1001 (O_1001,N_49911,N_49953);
xnor UO_1002 (O_1002,N_49883,N_49995);
nand UO_1003 (O_1003,N_49972,N_49975);
xor UO_1004 (O_1004,N_49798,N_49771);
nor UO_1005 (O_1005,N_49988,N_49944);
nand UO_1006 (O_1006,N_49849,N_49880);
xor UO_1007 (O_1007,N_49902,N_49798);
or UO_1008 (O_1008,N_49771,N_49758);
or UO_1009 (O_1009,N_49768,N_49914);
or UO_1010 (O_1010,N_49950,N_49804);
nor UO_1011 (O_1011,N_49876,N_49827);
nand UO_1012 (O_1012,N_49790,N_49998);
nand UO_1013 (O_1013,N_49980,N_49784);
xor UO_1014 (O_1014,N_49899,N_49969);
nor UO_1015 (O_1015,N_49980,N_49819);
or UO_1016 (O_1016,N_49857,N_49799);
nand UO_1017 (O_1017,N_49991,N_49822);
and UO_1018 (O_1018,N_49779,N_49905);
nand UO_1019 (O_1019,N_49774,N_49847);
and UO_1020 (O_1020,N_49948,N_49990);
xor UO_1021 (O_1021,N_49839,N_49768);
nor UO_1022 (O_1022,N_49961,N_49817);
or UO_1023 (O_1023,N_49830,N_49867);
xor UO_1024 (O_1024,N_49909,N_49814);
and UO_1025 (O_1025,N_49971,N_49879);
nand UO_1026 (O_1026,N_49854,N_49928);
xor UO_1027 (O_1027,N_49955,N_49804);
xor UO_1028 (O_1028,N_49793,N_49886);
nor UO_1029 (O_1029,N_49849,N_49829);
or UO_1030 (O_1030,N_49862,N_49830);
nor UO_1031 (O_1031,N_49962,N_49793);
nand UO_1032 (O_1032,N_49759,N_49887);
nand UO_1033 (O_1033,N_49891,N_49914);
nand UO_1034 (O_1034,N_49967,N_49941);
nor UO_1035 (O_1035,N_49753,N_49973);
nand UO_1036 (O_1036,N_49805,N_49850);
xor UO_1037 (O_1037,N_49768,N_49804);
nor UO_1038 (O_1038,N_49971,N_49990);
and UO_1039 (O_1039,N_49983,N_49955);
nor UO_1040 (O_1040,N_49968,N_49772);
xnor UO_1041 (O_1041,N_49917,N_49841);
nand UO_1042 (O_1042,N_49874,N_49853);
xnor UO_1043 (O_1043,N_49940,N_49756);
or UO_1044 (O_1044,N_49906,N_49943);
xor UO_1045 (O_1045,N_49754,N_49827);
and UO_1046 (O_1046,N_49786,N_49835);
nand UO_1047 (O_1047,N_49996,N_49917);
and UO_1048 (O_1048,N_49808,N_49926);
or UO_1049 (O_1049,N_49911,N_49900);
nand UO_1050 (O_1050,N_49832,N_49993);
and UO_1051 (O_1051,N_49782,N_49969);
xor UO_1052 (O_1052,N_49890,N_49932);
or UO_1053 (O_1053,N_49814,N_49886);
nand UO_1054 (O_1054,N_49837,N_49860);
and UO_1055 (O_1055,N_49936,N_49999);
or UO_1056 (O_1056,N_49844,N_49853);
xor UO_1057 (O_1057,N_49916,N_49893);
nand UO_1058 (O_1058,N_49939,N_49997);
and UO_1059 (O_1059,N_49868,N_49755);
or UO_1060 (O_1060,N_49920,N_49833);
and UO_1061 (O_1061,N_49915,N_49902);
nor UO_1062 (O_1062,N_49990,N_49883);
xor UO_1063 (O_1063,N_49771,N_49961);
nand UO_1064 (O_1064,N_49854,N_49907);
and UO_1065 (O_1065,N_49756,N_49992);
nor UO_1066 (O_1066,N_49811,N_49972);
nand UO_1067 (O_1067,N_49761,N_49796);
or UO_1068 (O_1068,N_49893,N_49967);
or UO_1069 (O_1069,N_49880,N_49903);
nand UO_1070 (O_1070,N_49779,N_49755);
nand UO_1071 (O_1071,N_49891,N_49921);
or UO_1072 (O_1072,N_49920,N_49842);
and UO_1073 (O_1073,N_49800,N_49866);
and UO_1074 (O_1074,N_49751,N_49943);
and UO_1075 (O_1075,N_49877,N_49911);
nand UO_1076 (O_1076,N_49892,N_49847);
or UO_1077 (O_1077,N_49955,N_49819);
and UO_1078 (O_1078,N_49984,N_49848);
nand UO_1079 (O_1079,N_49824,N_49901);
nor UO_1080 (O_1080,N_49753,N_49978);
xor UO_1081 (O_1081,N_49988,N_49887);
or UO_1082 (O_1082,N_49915,N_49886);
or UO_1083 (O_1083,N_49920,N_49817);
nor UO_1084 (O_1084,N_49973,N_49912);
nor UO_1085 (O_1085,N_49840,N_49947);
and UO_1086 (O_1086,N_49898,N_49822);
or UO_1087 (O_1087,N_49912,N_49776);
nand UO_1088 (O_1088,N_49946,N_49951);
nand UO_1089 (O_1089,N_49889,N_49900);
and UO_1090 (O_1090,N_49869,N_49804);
or UO_1091 (O_1091,N_49827,N_49884);
xnor UO_1092 (O_1092,N_49770,N_49883);
or UO_1093 (O_1093,N_49791,N_49979);
xor UO_1094 (O_1094,N_49777,N_49972);
nor UO_1095 (O_1095,N_49757,N_49964);
nand UO_1096 (O_1096,N_49969,N_49866);
nor UO_1097 (O_1097,N_49872,N_49998);
nor UO_1098 (O_1098,N_49909,N_49801);
nand UO_1099 (O_1099,N_49906,N_49792);
nor UO_1100 (O_1100,N_49867,N_49978);
xnor UO_1101 (O_1101,N_49927,N_49764);
xnor UO_1102 (O_1102,N_49805,N_49868);
xor UO_1103 (O_1103,N_49875,N_49780);
and UO_1104 (O_1104,N_49888,N_49762);
nor UO_1105 (O_1105,N_49999,N_49871);
xnor UO_1106 (O_1106,N_49875,N_49880);
xnor UO_1107 (O_1107,N_49867,N_49802);
xor UO_1108 (O_1108,N_49784,N_49801);
and UO_1109 (O_1109,N_49895,N_49872);
nand UO_1110 (O_1110,N_49803,N_49813);
nand UO_1111 (O_1111,N_49842,N_49809);
nor UO_1112 (O_1112,N_49863,N_49814);
nor UO_1113 (O_1113,N_49866,N_49857);
nor UO_1114 (O_1114,N_49802,N_49990);
or UO_1115 (O_1115,N_49961,N_49970);
or UO_1116 (O_1116,N_49796,N_49853);
xor UO_1117 (O_1117,N_49924,N_49789);
or UO_1118 (O_1118,N_49823,N_49796);
nor UO_1119 (O_1119,N_49948,N_49900);
nor UO_1120 (O_1120,N_49800,N_49968);
nor UO_1121 (O_1121,N_49803,N_49868);
xnor UO_1122 (O_1122,N_49837,N_49975);
and UO_1123 (O_1123,N_49859,N_49923);
and UO_1124 (O_1124,N_49835,N_49874);
nor UO_1125 (O_1125,N_49763,N_49848);
and UO_1126 (O_1126,N_49991,N_49783);
or UO_1127 (O_1127,N_49915,N_49867);
nor UO_1128 (O_1128,N_49989,N_49755);
xnor UO_1129 (O_1129,N_49981,N_49914);
or UO_1130 (O_1130,N_49760,N_49988);
xor UO_1131 (O_1131,N_49847,N_49795);
nand UO_1132 (O_1132,N_49977,N_49795);
nand UO_1133 (O_1133,N_49917,N_49915);
or UO_1134 (O_1134,N_49783,N_49928);
or UO_1135 (O_1135,N_49943,N_49948);
or UO_1136 (O_1136,N_49801,N_49823);
and UO_1137 (O_1137,N_49786,N_49876);
nand UO_1138 (O_1138,N_49840,N_49978);
or UO_1139 (O_1139,N_49812,N_49990);
nand UO_1140 (O_1140,N_49786,N_49780);
nor UO_1141 (O_1141,N_49999,N_49760);
or UO_1142 (O_1142,N_49769,N_49991);
nor UO_1143 (O_1143,N_49813,N_49752);
or UO_1144 (O_1144,N_49804,N_49829);
xor UO_1145 (O_1145,N_49856,N_49903);
and UO_1146 (O_1146,N_49986,N_49789);
nor UO_1147 (O_1147,N_49911,N_49848);
or UO_1148 (O_1148,N_49990,N_49813);
or UO_1149 (O_1149,N_49856,N_49913);
and UO_1150 (O_1150,N_49948,N_49901);
xnor UO_1151 (O_1151,N_49777,N_49986);
xor UO_1152 (O_1152,N_49928,N_49948);
nand UO_1153 (O_1153,N_49764,N_49991);
xor UO_1154 (O_1154,N_49759,N_49988);
or UO_1155 (O_1155,N_49843,N_49893);
or UO_1156 (O_1156,N_49834,N_49868);
nor UO_1157 (O_1157,N_49904,N_49891);
xnor UO_1158 (O_1158,N_49906,N_49833);
xnor UO_1159 (O_1159,N_49944,N_49840);
or UO_1160 (O_1160,N_49810,N_49877);
nor UO_1161 (O_1161,N_49820,N_49870);
nand UO_1162 (O_1162,N_49805,N_49874);
or UO_1163 (O_1163,N_49981,N_49782);
nand UO_1164 (O_1164,N_49956,N_49872);
xor UO_1165 (O_1165,N_49919,N_49893);
and UO_1166 (O_1166,N_49789,N_49876);
or UO_1167 (O_1167,N_49810,N_49912);
or UO_1168 (O_1168,N_49966,N_49904);
or UO_1169 (O_1169,N_49758,N_49906);
xnor UO_1170 (O_1170,N_49930,N_49788);
nand UO_1171 (O_1171,N_49783,N_49831);
nor UO_1172 (O_1172,N_49861,N_49978);
nor UO_1173 (O_1173,N_49953,N_49873);
nor UO_1174 (O_1174,N_49993,N_49852);
and UO_1175 (O_1175,N_49883,N_49893);
nor UO_1176 (O_1176,N_49915,N_49999);
or UO_1177 (O_1177,N_49968,N_49994);
or UO_1178 (O_1178,N_49926,N_49923);
xnor UO_1179 (O_1179,N_49912,N_49802);
xnor UO_1180 (O_1180,N_49829,N_49813);
nor UO_1181 (O_1181,N_49876,N_49905);
xnor UO_1182 (O_1182,N_49885,N_49813);
and UO_1183 (O_1183,N_49891,N_49842);
nand UO_1184 (O_1184,N_49856,N_49862);
xnor UO_1185 (O_1185,N_49981,N_49952);
and UO_1186 (O_1186,N_49981,N_49902);
nand UO_1187 (O_1187,N_49940,N_49962);
or UO_1188 (O_1188,N_49914,N_49810);
nand UO_1189 (O_1189,N_49757,N_49774);
xor UO_1190 (O_1190,N_49833,N_49787);
nor UO_1191 (O_1191,N_49845,N_49768);
xnor UO_1192 (O_1192,N_49969,N_49930);
nor UO_1193 (O_1193,N_49858,N_49948);
and UO_1194 (O_1194,N_49750,N_49771);
nor UO_1195 (O_1195,N_49927,N_49805);
nand UO_1196 (O_1196,N_49916,N_49778);
nor UO_1197 (O_1197,N_49788,N_49812);
xor UO_1198 (O_1198,N_49770,N_49966);
and UO_1199 (O_1199,N_49888,N_49910);
and UO_1200 (O_1200,N_49769,N_49988);
nor UO_1201 (O_1201,N_49970,N_49891);
and UO_1202 (O_1202,N_49868,N_49840);
nand UO_1203 (O_1203,N_49788,N_49770);
nor UO_1204 (O_1204,N_49818,N_49870);
nor UO_1205 (O_1205,N_49886,N_49952);
and UO_1206 (O_1206,N_49855,N_49819);
or UO_1207 (O_1207,N_49752,N_49769);
or UO_1208 (O_1208,N_49750,N_49967);
and UO_1209 (O_1209,N_49824,N_49951);
or UO_1210 (O_1210,N_49764,N_49930);
nor UO_1211 (O_1211,N_49902,N_49781);
or UO_1212 (O_1212,N_49926,N_49765);
nand UO_1213 (O_1213,N_49979,N_49895);
xnor UO_1214 (O_1214,N_49928,N_49774);
nand UO_1215 (O_1215,N_49821,N_49945);
nand UO_1216 (O_1216,N_49852,N_49954);
nand UO_1217 (O_1217,N_49867,N_49875);
and UO_1218 (O_1218,N_49975,N_49855);
xnor UO_1219 (O_1219,N_49918,N_49842);
and UO_1220 (O_1220,N_49811,N_49787);
and UO_1221 (O_1221,N_49975,N_49785);
nor UO_1222 (O_1222,N_49904,N_49994);
nand UO_1223 (O_1223,N_49892,N_49909);
or UO_1224 (O_1224,N_49858,N_49933);
nand UO_1225 (O_1225,N_49956,N_49874);
xor UO_1226 (O_1226,N_49857,N_49818);
nand UO_1227 (O_1227,N_49921,N_49942);
or UO_1228 (O_1228,N_49767,N_49809);
or UO_1229 (O_1229,N_49859,N_49879);
nand UO_1230 (O_1230,N_49800,N_49757);
nand UO_1231 (O_1231,N_49979,N_49869);
nand UO_1232 (O_1232,N_49918,N_49937);
xor UO_1233 (O_1233,N_49919,N_49869);
or UO_1234 (O_1234,N_49751,N_49922);
or UO_1235 (O_1235,N_49765,N_49898);
nor UO_1236 (O_1236,N_49841,N_49860);
xor UO_1237 (O_1237,N_49941,N_49876);
or UO_1238 (O_1238,N_49910,N_49980);
or UO_1239 (O_1239,N_49898,N_49844);
and UO_1240 (O_1240,N_49994,N_49929);
and UO_1241 (O_1241,N_49791,N_49777);
and UO_1242 (O_1242,N_49859,N_49915);
or UO_1243 (O_1243,N_49931,N_49771);
nor UO_1244 (O_1244,N_49959,N_49995);
nand UO_1245 (O_1245,N_49942,N_49870);
nand UO_1246 (O_1246,N_49996,N_49818);
or UO_1247 (O_1247,N_49858,N_49830);
nand UO_1248 (O_1248,N_49803,N_49962);
or UO_1249 (O_1249,N_49978,N_49844);
or UO_1250 (O_1250,N_49889,N_49924);
xnor UO_1251 (O_1251,N_49941,N_49921);
and UO_1252 (O_1252,N_49782,N_49751);
xnor UO_1253 (O_1253,N_49772,N_49945);
and UO_1254 (O_1254,N_49796,N_49815);
or UO_1255 (O_1255,N_49836,N_49789);
nand UO_1256 (O_1256,N_49928,N_49925);
xnor UO_1257 (O_1257,N_49962,N_49995);
and UO_1258 (O_1258,N_49925,N_49868);
or UO_1259 (O_1259,N_49983,N_49932);
or UO_1260 (O_1260,N_49847,N_49800);
nor UO_1261 (O_1261,N_49833,N_49947);
or UO_1262 (O_1262,N_49954,N_49938);
nand UO_1263 (O_1263,N_49905,N_49821);
and UO_1264 (O_1264,N_49870,N_49909);
nor UO_1265 (O_1265,N_49883,N_49762);
xnor UO_1266 (O_1266,N_49756,N_49785);
nor UO_1267 (O_1267,N_49951,N_49831);
xor UO_1268 (O_1268,N_49893,N_49905);
nor UO_1269 (O_1269,N_49931,N_49837);
and UO_1270 (O_1270,N_49887,N_49799);
and UO_1271 (O_1271,N_49946,N_49773);
or UO_1272 (O_1272,N_49755,N_49983);
or UO_1273 (O_1273,N_49842,N_49981);
xnor UO_1274 (O_1274,N_49890,N_49976);
nor UO_1275 (O_1275,N_49918,N_49997);
nor UO_1276 (O_1276,N_49883,N_49887);
nor UO_1277 (O_1277,N_49883,N_49886);
and UO_1278 (O_1278,N_49840,N_49847);
nor UO_1279 (O_1279,N_49999,N_49788);
nand UO_1280 (O_1280,N_49955,N_49754);
xnor UO_1281 (O_1281,N_49908,N_49883);
xor UO_1282 (O_1282,N_49929,N_49990);
xor UO_1283 (O_1283,N_49983,N_49867);
nand UO_1284 (O_1284,N_49863,N_49760);
nor UO_1285 (O_1285,N_49894,N_49983);
nand UO_1286 (O_1286,N_49960,N_49886);
nor UO_1287 (O_1287,N_49846,N_49784);
xor UO_1288 (O_1288,N_49761,N_49824);
nand UO_1289 (O_1289,N_49995,N_49808);
nand UO_1290 (O_1290,N_49982,N_49758);
nand UO_1291 (O_1291,N_49916,N_49983);
or UO_1292 (O_1292,N_49954,N_49755);
nor UO_1293 (O_1293,N_49756,N_49887);
nand UO_1294 (O_1294,N_49771,N_49782);
or UO_1295 (O_1295,N_49814,N_49869);
nand UO_1296 (O_1296,N_49869,N_49800);
nor UO_1297 (O_1297,N_49913,N_49998);
nor UO_1298 (O_1298,N_49786,N_49791);
or UO_1299 (O_1299,N_49993,N_49986);
nand UO_1300 (O_1300,N_49757,N_49998);
nor UO_1301 (O_1301,N_49765,N_49883);
or UO_1302 (O_1302,N_49807,N_49821);
nor UO_1303 (O_1303,N_49784,N_49813);
nor UO_1304 (O_1304,N_49835,N_49892);
and UO_1305 (O_1305,N_49770,N_49996);
or UO_1306 (O_1306,N_49833,N_49934);
nor UO_1307 (O_1307,N_49772,N_49813);
or UO_1308 (O_1308,N_49881,N_49786);
or UO_1309 (O_1309,N_49858,N_49813);
nor UO_1310 (O_1310,N_49911,N_49778);
nor UO_1311 (O_1311,N_49978,N_49832);
or UO_1312 (O_1312,N_49892,N_49753);
nand UO_1313 (O_1313,N_49874,N_49761);
xor UO_1314 (O_1314,N_49803,N_49765);
nor UO_1315 (O_1315,N_49989,N_49798);
xnor UO_1316 (O_1316,N_49758,N_49800);
xor UO_1317 (O_1317,N_49868,N_49811);
and UO_1318 (O_1318,N_49950,N_49988);
or UO_1319 (O_1319,N_49971,N_49781);
or UO_1320 (O_1320,N_49882,N_49923);
and UO_1321 (O_1321,N_49985,N_49761);
xor UO_1322 (O_1322,N_49904,N_49979);
nor UO_1323 (O_1323,N_49847,N_49945);
nor UO_1324 (O_1324,N_49769,N_49782);
or UO_1325 (O_1325,N_49980,N_49878);
nor UO_1326 (O_1326,N_49861,N_49810);
nand UO_1327 (O_1327,N_49884,N_49857);
nand UO_1328 (O_1328,N_49906,N_49979);
nand UO_1329 (O_1329,N_49821,N_49791);
or UO_1330 (O_1330,N_49841,N_49764);
nor UO_1331 (O_1331,N_49820,N_49846);
or UO_1332 (O_1332,N_49974,N_49814);
and UO_1333 (O_1333,N_49752,N_49888);
nand UO_1334 (O_1334,N_49809,N_49752);
nor UO_1335 (O_1335,N_49877,N_49913);
and UO_1336 (O_1336,N_49970,N_49884);
or UO_1337 (O_1337,N_49773,N_49764);
and UO_1338 (O_1338,N_49788,N_49998);
or UO_1339 (O_1339,N_49959,N_49856);
nand UO_1340 (O_1340,N_49780,N_49830);
nor UO_1341 (O_1341,N_49958,N_49894);
nor UO_1342 (O_1342,N_49913,N_49876);
and UO_1343 (O_1343,N_49852,N_49990);
nand UO_1344 (O_1344,N_49935,N_49833);
nor UO_1345 (O_1345,N_49793,N_49954);
xnor UO_1346 (O_1346,N_49854,N_49820);
and UO_1347 (O_1347,N_49875,N_49836);
xor UO_1348 (O_1348,N_49929,N_49819);
or UO_1349 (O_1349,N_49867,N_49925);
or UO_1350 (O_1350,N_49944,N_49787);
nor UO_1351 (O_1351,N_49885,N_49830);
or UO_1352 (O_1352,N_49945,N_49986);
nor UO_1353 (O_1353,N_49954,N_49953);
nor UO_1354 (O_1354,N_49808,N_49753);
nor UO_1355 (O_1355,N_49932,N_49987);
and UO_1356 (O_1356,N_49996,N_49840);
or UO_1357 (O_1357,N_49891,N_49944);
or UO_1358 (O_1358,N_49839,N_49868);
and UO_1359 (O_1359,N_49844,N_49925);
xor UO_1360 (O_1360,N_49943,N_49911);
nor UO_1361 (O_1361,N_49813,N_49787);
nand UO_1362 (O_1362,N_49796,N_49891);
nor UO_1363 (O_1363,N_49844,N_49930);
nor UO_1364 (O_1364,N_49840,N_49766);
nand UO_1365 (O_1365,N_49827,N_49973);
nor UO_1366 (O_1366,N_49814,N_49868);
nor UO_1367 (O_1367,N_49966,N_49843);
nor UO_1368 (O_1368,N_49825,N_49953);
xnor UO_1369 (O_1369,N_49807,N_49917);
and UO_1370 (O_1370,N_49961,N_49926);
or UO_1371 (O_1371,N_49761,N_49795);
and UO_1372 (O_1372,N_49780,N_49965);
nor UO_1373 (O_1373,N_49879,N_49906);
or UO_1374 (O_1374,N_49814,N_49884);
and UO_1375 (O_1375,N_49951,N_49967);
and UO_1376 (O_1376,N_49866,N_49925);
and UO_1377 (O_1377,N_49992,N_49795);
or UO_1378 (O_1378,N_49925,N_49892);
nor UO_1379 (O_1379,N_49783,N_49972);
or UO_1380 (O_1380,N_49940,N_49801);
or UO_1381 (O_1381,N_49786,N_49968);
and UO_1382 (O_1382,N_49918,N_49973);
nand UO_1383 (O_1383,N_49767,N_49907);
and UO_1384 (O_1384,N_49977,N_49846);
nand UO_1385 (O_1385,N_49988,N_49852);
nor UO_1386 (O_1386,N_49941,N_49946);
and UO_1387 (O_1387,N_49787,N_49789);
or UO_1388 (O_1388,N_49846,N_49803);
nor UO_1389 (O_1389,N_49885,N_49846);
xor UO_1390 (O_1390,N_49798,N_49918);
and UO_1391 (O_1391,N_49775,N_49905);
or UO_1392 (O_1392,N_49937,N_49933);
or UO_1393 (O_1393,N_49853,N_49756);
xnor UO_1394 (O_1394,N_49767,N_49888);
and UO_1395 (O_1395,N_49912,N_49825);
nor UO_1396 (O_1396,N_49955,N_49810);
or UO_1397 (O_1397,N_49857,N_49870);
nand UO_1398 (O_1398,N_49833,N_49909);
nor UO_1399 (O_1399,N_49853,N_49810);
nor UO_1400 (O_1400,N_49914,N_49780);
and UO_1401 (O_1401,N_49894,N_49796);
and UO_1402 (O_1402,N_49973,N_49879);
nor UO_1403 (O_1403,N_49803,N_49867);
xnor UO_1404 (O_1404,N_49839,N_49986);
or UO_1405 (O_1405,N_49814,N_49800);
or UO_1406 (O_1406,N_49804,N_49790);
nor UO_1407 (O_1407,N_49906,N_49844);
nand UO_1408 (O_1408,N_49881,N_49852);
xnor UO_1409 (O_1409,N_49919,N_49931);
xnor UO_1410 (O_1410,N_49945,N_49797);
nor UO_1411 (O_1411,N_49903,N_49935);
nand UO_1412 (O_1412,N_49802,N_49851);
or UO_1413 (O_1413,N_49874,N_49833);
nor UO_1414 (O_1414,N_49890,N_49790);
xor UO_1415 (O_1415,N_49758,N_49924);
or UO_1416 (O_1416,N_49961,N_49809);
nand UO_1417 (O_1417,N_49992,N_49884);
or UO_1418 (O_1418,N_49946,N_49806);
nor UO_1419 (O_1419,N_49790,N_49882);
or UO_1420 (O_1420,N_49942,N_49808);
nor UO_1421 (O_1421,N_49994,N_49835);
or UO_1422 (O_1422,N_49938,N_49886);
and UO_1423 (O_1423,N_49981,N_49804);
xnor UO_1424 (O_1424,N_49877,N_49941);
nand UO_1425 (O_1425,N_49943,N_49996);
xnor UO_1426 (O_1426,N_49791,N_49957);
nand UO_1427 (O_1427,N_49928,N_49904);
nand UO_1428 (O_1428,N_49922,N_49916);
and UO_1429 (O_1429,N_49841,N_49929);
or UO_1430 (O_1430,N_49869,N_49779);
nand UO_1431 (O_1431,N_49821,N_49955);
or UO_1432 (O_1432,N_49818,N_49782);
nor UO_1433 (O_1433,N_49816,N_49926);
nor UO_1434 (O_1434,N_49904,N_49787);
nand UO_1435 (O_1435,N_49940,N_49755);
or UO_1436 (O_1436,N_49840,N_49986);
and UO_1437 (O_1437,N_49765,N_49901);
xnor UO_1438 (O_1438,N_49960,N_49994);
nor UO_1439 (O_1439,N_49824,N_49857);
nand UO_1440 (O_1440,N_49861,N_49793);
or UO_1441 (O_1441,N_49883,N_49960);
nand UO_1442 (O_1442,N_49775,N_49790);
and UO_1443 (O_1443,N_49975,N_49946);
xnor UO_1444 (O_1444,N_49801,N_49841);
nand UO_1445 (O_1445,N_49842,N_49811);
xnor UO_1446 (O_1446,N_49758,N_49994);
xnor UO_1447 (O_1447,N_49838,N_49867);
nor UO_1448 (O_1448,N_49839,N_49811);
and UO_1449 (O_1449,N_49797,N_49840);
nor UO_1450 (O_1450,N_49755,N_49977);
xor UO_1451 (O_1451,N_49933,N_49877);
xnor UO_1452 (O_1452,N_49899,N_49877);
or UO_1453 (O_1453,N_49838,N_49893);
nor UO_1454 (O_1454,N_49760,N_49918);
or UO_1455 (O_1455,N_49865,N_49966);
and UO_1456 (O_1456,N_49967,N_49925);
or UO_1457 (O_1457,N_49799,N_49792);
or UO_1458 (O_1458,N_49958,N_49794);
or UO_1459 (O_1459,N_49773,N_49945);
xnor UO_1460 (O_1460,N_49927,N_49899);
nand UO_1461 (O_1461,N_49859,N_49826);
and UO_1462 (O_1462,N_49826,N_49823);
nand UO_1463 (O_1463,N_49939,N_49985);
or UO_1464 (O_1464,N_49997,N_49864);
or UO_1465 (O_1465,N_49951,N_49932);
xnor UO_1466 (O_1466,N_49853,N_49953);
xnor UO_1467 (O_1467,N_49851,N_49938);
nor UO_1468 (O_1468,N_49854,N_49944);
or UO_1469 (O_1469,N_49899,N_49995);
nor UO_1470 (O_1470,N_49762,N_49880);
nand UO_1471 (O_1471,N_49895,N_49819);
or UO_1472 (O_1472,N_49826,N_49751);
xor UO_1473 (O_1473,N_49919,N_49896);
and UO_1474 (O_1474,N_49967,N_49952);
or UO_1475 (O_1475,N_49888,N_49778);
or UO_1476 (O_1476,N_49991,N_49809);
xnor UO_1477 (O_1477,N_49935,N_49805);
nand UO_1478 (O_1478,N_49854,N_49892);
nand UO_1479 (O_1479,N_49942,N_49750);
or UO_1480 (O_1480,N_49829,N_49904);
and UO_1481 (O_1481,N_49759,N_49989);
nand UO_1482 (O_1482,N_49914,N_49888);
nor UO_1483 (O_1483,N_49787,N_49903);
nand UO_1484 (O_1484,N_49913,N_49899);
nor UO_1485 (O_1485,N_49896,N_49781);
nand UO_1486 (O_1486,N_49782,N_49977);
nand UO_1487 (O_1487,N_49993,N_49799);
or UO_1488 (O_1488,N_49846,N_49869);
xnor UO_1489 (O_1489,N_49948,N_49888);
nand UO_1490 (O_1490,N_49868,N_49841);
xnor UO_1491 (O_1491,N_49997,N_49820);
xor UO_1492 (O_1492,N_49920,N_49993);
nand UO_1493 (O_1493,N_49828,N_49778);
nor UO_1494 (O_1494,N_49833,N_49870);
or UO_1495 (O_1495,N_49970,N_49822);
and UO_1496 (O_1496,N_49950,N_49987);
nand UO_1497 (O_1497,N_49856,N_49865);
xor UO_1498 (O_1498,N_49835,N_49956);
xor UO_1499 (O_1499,N_49868,N_49915);
nand UO_1500 (O_1500,N_49951,N_49842);
xnor UO_1501 (O_1501,N_49768,N_49941);
or UO_1502 (O_1502,N_49820,N_49924);
nor UO_1503 (O_1503,N_49873,N_49824);
nand UO_1504 (O_1504,N_49820,N_49984);
nor UO_1505 (O_1505,N_49888,N_49859);
xor UO_1506 (O_1506,N_49938,N_49946);
nor UO_1507 (O_1507,N_49936,N_49947);
xnor UO_1508 (O_1508,N_49957,N_49936);
nand UO_1509 (O_1509,N_49972,N_49913);
nor UO_1510 (O_1510,N_49782,N_49999);
or UO_1511 (O_1511,N_49943,N_49918);
nand UO_1512 (O_1512,N_49761,N_49902);
nor UO_1513 (O_1513,N_49837,N_49789);
or UO_1514 (O_1514,N_49868,N_49791);
and UO_1515 (O_1515,N_49880,N_49863);
xnor UO_1516 (O_1516,N_49848,N_49863);
nand UO_1517 (O_1517,N_49931,N_49814);
or UO_1518 (O_1518,N_49889,N_49876);
nand UO_1519 (O_1519,N_49894,N_49772);
nor UO_1520 (O_1520,N_49995,N_49775);
and UO_1521 (O_1521,N_49877,N_49962);
nand UO_1522 (O_1522,N_49795,N_49784);
xnor UO_1523 (O_1523,N_49940,N_49775);
or UO_1524 (O_1524,N_49794,N_49965);
and UO_1525 (O_1525,N_49876,N_49936);
or UO_1526 (O_1526,N_49926,N_49900);
xor UO_1527 (O_1527,N_49938,N_49834);
nand UO_1528 (O_1528,N_49769,N_49842);
or UO_1529 (O_1529,N_49913,N_49871);
or UO_1530 (O_1530,N_49938,N_49943);
nand UO_1531 (O_1531,N_49826,N_49989);
nor UO_1532 (O_1532,N_49768,N_49798);
nor UO_1533 (O_1533,N_49765,N_49960);
nor UO_1534 (O_1534,N_49935,N_49844);
nand UO_1535 (O_1535,N_49822,N_49838);
nor UO_1536 (O_1536,N_49952,N_49822);
nand UO_1537 (O_1537,N_49796,N_49765);
nor UO_1538 (O_1538,N_49874,N_49814);
nand UO_1539 (O_1539,N_49937,N_49779);
and UO_1540 (O_1540,N_49853,N_49998);
xor UO_1541 (O_1541,N_49917,N_49805);
nand UO_1542 (O_1542,N_49781,N_49764);
nand UO_1543 (O_1543,N_49908,N_49944);
or UO_1544 (O_1544,N_49832,N_49834);
and UO_1545 (O_1545,N_49784,N_49979);
and UO_1546 (O_1546,N_49944,N_49882);
nor UO_1547 (O_1547,N_49890,N_49813);
nand UO_1548 (O_1548,N_49989,N_49817);
and UO_1549 (O_1549,N_49989,N_49881);
or UO_1550 (O_1550,N_49903,N_49871);
or UO_1551 (O_1551,N_49881,N_49782);
and UO_1552 (O_1552,N_49893,N_49845);
nor UO_1553 (O_1553,N_49950,N_49796);
xnor UO_1554 (O_1554,N_49907,N_49837);
or UO_1555 (O_1555,N_49990,N_49858);
nor UO_1556 (O_1556,N_49823,N_49850);
and UO_1557 (O_1557,N_49795,N_49783);
xnor UO_1558 (O_1558,N_49946,N_49842);
and UO_1559 (O_1559,N_49855,N_49958);
and UO_1560 (O_1560,N_49891,N_49811);
nor UO_1561 (O_1561,N_49751,N_49812);
nand UO_1562 (O_1562,N_49804,N_49916);
or UO_1563 (O_1563,N_49950,N_49760);
or UO_1564 (O_1564,N_49836,N_49778);
nor UO_1565 (O_1565,N_49891,N_49812);
and UO_1566 (O_1566,N_49901,N_49917);
nand UO_1567 (O_1567,N_49839,N_49759);
or UO_1568 (O_1568,N_49891,N_49870);
nor UO_1569 (O_1569,N_49855,N_49935);
and UO_1570 (O_1570,N_49991,N_49954);
and UO_1571 (O_1571,N_49901,N_49925);
nor UO_1572 (O_1572,N_49970,N_49971);
or UO_1573 (O_1573,N_49973,N_49937);
nor UO_1574 (O_1574,N_49785,N_49872);
and UO_1575 (O_1575,N_49962,N_49766);
nor UO_1576 (O_1576,N_49976,N_49990);
nand UO_1577 (O_1577,N_49946,N_49846);
and UO_1578 (O_1578,N_49944,N_49790);
nor UO_1579 (O_1579,N_49944,N_49976);
xor UO_1580 (O_1580,N_49804,N_49832);
and UO_1581 (O_1581,N_49966,N_49955);
and UO_1582 (O_1582,N_49920,N_49796);
and UO_1583 (O_1583,N_49890,N_49974);
and UO_1584 (O_1584,N_49768,N_49906);
or UO_1585 (O_1585,N_49780,N_49767);
or UO_1586 (O_1586,N_49947,N_49827);
or UO_1587 (O_1587,N_49881,N_49990);
nor UO_1588 (O_1588,N_49759,N_49905);
nand UO_1589 (O_1589,N_49851,N_49875);
nor UO_1590 (O_1590,N_49943,N_49819);
nor UO_1591 (O_1591,N_49833,N_49965);
and UO_1592 (O_1592,N_49779,N_49868);
xor UO_1593 (O_1593,N_49960,N_49840);
xor UO_1594 (O_1594,N_49802,N_49962);
or UO_1595 (O_1595,N_49884,N_49895);
or UO_1596 (O_1596,N_49859,N_49922);
nor UO_1597 (O_1597,N_49916,N_49978);
or UO_1598 (O_1598,N_49963,N_49901);
or UO_1599 (O_1599,N_49798,N_49824);
nor UO_1600 (O_1600,N_49802,N_49826);
xnor UO_1601 (O_1601,N_49961,N_49779);
and UO_1602 (O_1602,N_49929,N_49948);
and UO_1603 (O_1603,N_49965,N_49919);
or UO_1604 (O_1604,N_49754,N_49967);
and UO_1605 (O_1605,N_49875,N_49782);
and UO_1606 (O_1606,N_49833,N_49849);
xor UO_1607 (O_1607,N_49761,N_49837);
nand UO_1608 (O_1608,N_49822,N_49775);
xnor UO_1609 (O_1609,N_49843,N_49999);
nand UO_1610 (O_1610,N_49921,N_49753);
nand UO_1611 (O_1611,N_49979,N_49816);
nor UO_1612 (O_1612,N_49917,N_49788);
nor UO_1613 (O_1613,N_49816,N_49975);
and UO_1614 (O_1614,N_49805,N_49813);
and UO_1615 (O_1615,N_49823,N_49860);
nor UO_1616 (O_1616,N_49912,N_49788);
or UO_1617 (O_1617,N_49961,N_49992);
or UO_1618 (O_1618,N_49795,N_49854);
nand UO_1619 (O_1619,N_49786,N_49892);
nand UO_1620 (O_1620,N_49906,N_49971);
xor UO_1621 (O_1621,N_49982,N_49829);
xor UO_1622 (O_1622,N_49760,N_49791);
and UO_1623 (O_1623,N_49893,N_49975);
or UO_1624 (O_1624,N_49779,N_49765);
or UO_1625 (O_1625,N_49988,N_49943);
nor UO_1626 (O_1626,N_49970,N_49782);
nand UO_1627 (O_1627,N_49787,N_49798);
and UO_1628 (O_1628,N_49830,N_49958);
or UO_1629 (O_1629,N_49857,N_49766);
or UO_1630 (O_1630,N_49824,N_49797);
nand UO_1631 (O_1631,N_49959,N_49945);
or UO_1632 (O_1632,N_49995,N_49767);
and UO_1633 (O_1633,N_49871,N_49837);
or UO_1634 (O_1634,N_49933,N_49873);
nand UO_1635 (O_1635,N_49947,N_49924);
and UO_1636 (O_1636,N_49755,N_49927);
or UO_1637 (O_1637,N_49766,N_49957);
or UO_1638 (O_1638,N_49861,N_49941);
and UO_1639 (O_1639,N_49758,N_49901);
or UO_1640 (O_1640,N_49811,N_49887);
nand UO_1641 (O_1641,N_49948,N_49870);
or UO_1642 (O_1642,N_49898,N_49814);
nand UO_1643 (O_1643,N_49810,N_49796);
nand UO_1644 (O_1644,N_49979,N_49819);
nor UO_1645 (O_1645,N_49768,N_49857);
or UO_1646 (O_1646,N_49986,N_49933);
nand UO_1647 (O_1647,N_49873,N_49973);
xor UO_1648 (O_1648,N_49919,N_49755);
nand UO_1649 (O_1649,N_49941,N_49926);
xnor UO_1650 (O_1650,N_49873,N_49877);
nor UO_1651 (O_1651,N_49946,N_49800);
xor UO_1652 (O_1652,N_49920,N_49873);
nor UO_1653 (O_1653,N_49981,N_49944);
nor UO_1654 (O_1654,N_49969,N_49790);
and UO_1655 (O_1655,N_49901,N_49955);
nand UO_1656 (O_1656,N_49766,N_49939);
nand UO_1657 (O_1657,N_49917,N_49947);
xnor UO_1658 (O_1658,N_49769,N_49873);
nor UO_1659 (O_1659,N_49992,N_49780);
and UO_1660 (O_1660,N_49973,N_49857);
xnor UO_1661 (O_1661,N_49959,N_49848);
or UO_1662 (O_1662,N_49992,N_49958);
nand UO_1663 (O_1663,N_49968,N_49976);
or UO_1664 (O_1664,N_49911,N_49831);
and UO_1665 (O_1665,N_49872,N_49854);
and UO_1666 (O_1666,N_49793,N_49750);
xor UO_1667 (O_1667,N_49920,N_49771);
and UO_1668 (O_1668,N_49973,N_49855);
nor UO_1669 (O_1669,N_49966,N_49792);
nand UO_1670 (O_1670,N_49822,N_49989);
nor UO_1671 (O_1671,N_49776,N_49955);
xor UO_1672 (O_1672,N_49801,N_49820);
nor UO_1673 (O_1673,N_49751,N_49901);
and UO_1674 (O_1674,N_49755,N_49936);
and UO_1675 (O_1675,N_49814,N_49809);
and UO_1676 (O_1676,N_49984,N_49819);
xor UO_1677 (O_1677,N_49896,N_49995);
xnor UO_1678 (O_1678,N_49990,N_49909);
nand UO_1679 (O_1679,N_49775,N_49911);
or UO_1680 (O_1680,N_49898,N_49997);
and UO_1681 (O_1681,N_49877,N_49851);
or UO_1682 (O_1682,N_49871,N_49902);
or UO_1683 (O_1683,N_49939,N_49946);
nand UO_1684 (O_1684,N_49902,N_49945);
and UO_1685 (O_1685,N_49768,N_49786);
and UO_1686 (O_1686,N_49904,N_49835);
and UO_1687 (O_1687,N_49761,N_49895);
or UO_1688 (O_1688,N_49939,N_49805);
nor UO_1689 (O_1689,N_49919,N_49882);
nand UO_1690 (O_1690,N_49980,N_49917);
nand UO_1691 (O_1691,N_49859,N_49968);
nand UO_1692 (O_1692,N_49896,N_49951);
nor UO_1693 (O_1693,N_49875,N_49945);
or UO_1694 (O_1694,N_49875,N_49883);
and UO_1695 (O_1695,N_49803,N_49927);
xnor UO_1696 (O_1696,N_49794,N_49917);
xor UO_1697 (O_1697,N_49770,N_49878);
nand UO_1698 (O_1698,N_49956,N_49869);
nand UO_1699 (O_1699,N_49918,N_49905);
and UO_1700 (O_1700,N_49934,N_49888);
and UO_1701 (O_1701,N_49796,N_49751);
or UO_1702 (O_1702,N_49820,N_49813);
or UO_1703 (O_1703,N_49832,N_49986);
or UO_1704 (O_1704,N_49857,N_49900);
xnor UO_1705 (O_1705,N_49779,N_49962);
nand UO_1706 (O_1706,N_49809,N_49922);
nor UO_1707 (O_1707,N_49983,N_49982);
and UO_1708 (O_1708,N_49770,N_49785);
xor UO_1709 (O_1709,N_49994,N_49896);
xor UO_1710 (O_1710,N_49761,N_49866);
xor UO_1711 (O_1711,N_49868,N_49908);
or UO_1712 (O_1712,N_49934,N_49921);
or UO_1713 (O_1713,N_49962,N_49780);
nand UO_1714 (O_1714,N_49813,N_49843);
and UO_1715 (O_1715,N_49907,N_49911);
and UO_1716 (O_1716,N_49952,N_49922);
nand UO_1717 (O_1717,N_49946,N_49810);
nor UO_1718 (O_1718,N_49797,N_49769);
nor UO_1719 (O_1719,N_49750,N_49773);
nand UO_1720 (O_1720,N_49838,N_49890);
xnor UO_1721 (O_1721,N_49861,N_49812);
nor UO_1722 (O_1722,N_49813,N_49818);
or UO_1723 (O_1723,N_49776,N_49759);
and UO_1724 (O_1724,N_49875,N_49847);
xnor UO_1725 (O_1725,N_49936,N_49824);
and UO_1726 (O_1726,N_49980,N_49995);
nand UO_1727 (O_1727,N_49972,N_49828);
xnor UO_1728 (O_1728,N_49828,N_49919);
and UO_1729 (O_1729,N_49972,N_49812);
xor UO_1730 (O_1730,N_49768,N_49800);
or UO_1731 (O_1731,N_49767,N_49992);
nand UO_1732 (O_1732,N_49913,N_49785);
nand UO_1733 (O_1733,N_49984,N_49989);
and UO_1734 (O_1734,N_49948,N_49998);
nand UO_1735 (O_1735,N_49917,N_49967);
nand UO_1736 (O_1736,N_49833,N_49770);
nor UO_1737 (O_1737,N_49811,N_49903);
xor UO_1738 (O_1738,N_49819,N_49807);
and UO_1739 (O_1739,N_49838,N_49899);
or UO_1740 (O_1740,N_49996,N_49845);
or UO_1741 (O_1741,N_49868,N_49918);
xor UO_1742 (O_1742,N_49823,N_49885);
and UO_1743 (O_1743,N_49867,N_49784);
xor UO_1744 (O_1744,N_49958,N_49951);
nor UO_1745 (O_1745,N_49846,N_49756);
nor UO_1746 (O_1746,N_49874,N_49847);
or UO_1747 (O_1747,N_49853,N_49857);
nor UO_1748 (O_1748,N_49942,N_49751);
xnor UO_1749 (O_1749,N_49792,N_49912);
and UO_1750 (O_1750,N_49770,N_49939);
or UO_1751 (O_1751,N_49900,N_49871);
and UO_1752 (O_1752,N_49769,N_49869);
xor UO_1753 (O_1753,N_49773,N_49860);
nor UO_1754 (O_1754,N_49914,N_49877);
and UO_1755 (O_1755,N_49807,N_49798);
xnor UO_1756 (O_1756,N_49804,N_49991);
xor UO_1757 (O_1757,N_49916,N_49763);
nand UO_1758 (O_1758,N_49773,N_49852);
nor UO_1759 (O_1759,N_49848,N_49822);
and UO_1760 (O_1760,N_49871,N_49846);
nand UO_1761 (O_1761,N_49782,N_49893);
nor UO_1762 (O_1762,N_49852,N_49824);
xnor UO_1763 (O_1763,N_49872,N_49973);
and UO_1764 (O_1764,N_49833,N_49851);
nor UO_1765 (O_1765,N_49763,N_49934);
nand UO_1766 (O_1766,N_49917,N_49772);
nand UO_1767 (O_1767,N_49807,N_49862);
or UO_1768 (O_1768,N_49933,N_49957);
nand UO_1769 (O_1769,N_49808,N_49924);
xor UO_1770 (O_1770,N_49946,N_49973);
nand UO_1771 (O_1771,N_49933,N_49921);
and UO_1772 (O_1772,N_49955,N_49856);
and UO_1773 (O_1773,N_49788,N_49833);
nor UO_1774 (O_1774,N_49929,N_49896);
or UO_1775 (O_1775,N_49869,N_49909);
or UO_1776 (O_1776,N_49826,N_49909);
nor UO_1777 (O_1777,N_49845,N_49954);
or UO_1778 (O_1778,N_49790,N_49875);
nand UO_1779 (O_1779,N_49866,N_49899);
and UO_1780 (O_1780,N_49843,N_49859);
or UO_1781 (O_1781,N_49851,N_49953);
and UO_1782 (O_1782,N_49817,N_49921);
xor UO_1783 (O_1783,N_49870,N_49929);
and UO_1784 (O_1784,N_49976,N_49821);
or UO_1785 (O_1785,N_49959,N_49972);
and UO_1786 (O_1786,N_49771,N_49948);
nand UO_1787 (O_1787,N_49983,N_49850);
nor UO_1788 (O_1788,N_49843,N_49970);
nor UO_1789 (O_1789,N_49971,N_49939);
and UO_1790 (O_1790,N_49752,N_49884);
or UO_1791 (O_1791,N_49770,N_49921);
and UO_1792 (O_1792,N_49772,N_49912);
nand UO_1793 (O_1793,N_49814,N_49810);
xor UO_1794 (O_1794,N_49916,N_49982);
xor UO_1795 (O_1795,N_49903,N_49908);
nand UO_1796 (O_1796,N_49849,N_49781);
or UO_1797 (O_1797,N_49764,N_49782);
and UO_1798 (O_1798,N_49777,N_49915);
and UO_1799 (O_1799,N_49844,N_49997);
and UO_1800 (O_1800,N_49983,N_49929);
and UO_1801 (O_1801,N_49897,N_49756);
nor UO_1802 (O_1802,N_49891,N_49889);
nand UO_1803 (O_1803,N_49818,N_49772);
nand UO_1804 (O_1804,N_49751,N_49846);
xor UO_1805 (O_1805,N_49865,N_49945);
and UO_1806 (O_1806,N_49920,N_49819);
or UO_1807 (O_1807,N_49819,N_49963);
xnor UO_1808 (O_1808,N_49782,N_49984);
nand UO_1809 (O_1809,N_49760,N_49771);
or UO_1810 (O_1810,N_49891,N_49873);
nor UO_1811 (O_1811,N_49959,N_49941);
or UO_1812 (O_1812,N_49963,N_49936);
nand UO_1813 (O_1813,N_49945,N_49855);
xor UO_1814 (O_1814,N_49939,N_49867);
xnor UO_1815 (O_1815,N_49779,N_49974);
xor UO_1816 (O_1816,N_49811,N_49786);
nor UO_1817 (O_1817,N_49793,N_49876);
nand UO_1818 (O_1818,N_49939,N_49848);
nand UO_1819 (O_1819,N_49756,N_49962);
xor UO_1820 (O_1820,N_49902,N_49908);
xnor UO_1821 (O_1821,N_49889,N_49894);
xor UO_1822 (O_1822,N_49750,N_49843);
or UO_1823 (O_1823,N_49843,N_49766);
nand UO_1824 (O_1824,N_49848,N_49769);
or UO_1825 (O_1825,N_49994,N_49873);
xnor UO_1826 (O_1826,N_49795,N_49896);
or UO_1827 (O_1827,N_49798,N_49779);
nand UO_1828 (O_1828,N_49942,N_49869);
or UO_1829 (O_1829,N_49818,N_49768);
or UO_1830 (O_1830,N_49845,N_49990);
and UO_1831 (O_1831,N_49763,N_49938);
or UO_1832 (O_1832,N_49799,N_49907);
or UO_1833 (O_1833,N_49969,N_49779);
or UO_1834 (O_1834,N_49755,N_49782);
nand UO_1835 (O_1835,N_49901,N_49820);
nand UO_1836 (O_1836,N_49809,N_49896);
nand UO_1837 (O_1837,N_49944,N_49943);
nand UO_1838 (O_1838,N_49856,N_49860);
nor UO_1839 (O_1839,N_49815,N_49911);
and UO_1840 (O_1840,N_49925,N_49948);
xor UO_1841 (O_1841,N_49945,N_49952);
or UO_1842 (O_1842,N_49889,N_49878);
nor UO_1843 (O_1843,N_49918,N_49934);
and UO_1844 (O_1844,N_49961,N_49805);
nand UO_1845 (O_1845,N_49750,N_49869);
nand UO_1846 (O_1846,N_49893,N_49828);
and UO_1847 (O_1847,N_49849,N_49909);
nor UO_1848 (O_1848,N_49972,N_49902);
and UO_1849 (O_1849,N_49805,N_49947);
and UO_1850 (O_1850,N_49935,N_49900);
xor UO_1851 (O_1851,N_49967,N_49973);
and UO_1852 (O_1852,N_49937,N_49872);
or UO_1853 (O_1853,N_49752,N_49885);
xor UO_1854 (O_1854,N_49800,N_49786);
nor UO_1855 (O_1855,N_49963,N_49877);
xnor UO_1856 (O_1856,N_49826,N_49816);
and UO_1857 (O_1857,N_49883,N_49846);
nand UO_1858 (O_1858,N_49899,N_49978);
xnor UO_1859 (O_1859,N_49991,N_49844);
xor UO_1860 (O_1860,N_49778,N_49831);
nor UO_1861 (O_1861,N_49966,N_49834);
nand UO_1862 (O_1862,N_49892,N_49823);
xnor UO_1863 (O_1863,N_49997,N_49750);
or UO_1864 (O_1864,N_49888,N_49814);
and UO_1865 (O_1865,N_49903,N_49815);
or UO_1866 (O_1866,N_49955,N_49939);
xnor UO_1867 (O_1867,N_49788,N_49981);
and UO_1868 (O_1868,N_49973,N_49770);
xnor UO_1869 (O_1869,N_49959,N_49827);
nor UO_1870 (O_1870,N_49953,N_49955);
and UO_1871 (O_1871,N_49949,N_49831);
nand UO_1872 (O_1872,N_49870,N_49970);
and UO_1873 (O_1873,N_49959,N_49948);
nor UO_1874 (O_1874,N_49812,N_49782);
nand UO_1875 (O_1875,N_49873,N_49911);
nor UO_1876 (O_1876,N_49825,N_49789);
nor UO_1877 (O_1877,N_49968,N_49818);
and UO_1878 (O_1878,N_49893,N_49911);
xnor UO_1879 (O_1879,N_49965,N_49900);
nor UO_1880 (O_1880,N_49925,N_49907);
nor UO_1881 (O_1881,N_49876,N_49912);
nor UO_1882 (O_1882,N_49914,N_49781);
or UO_1883 (O_1883,N_49882,N_49814);
and UO_1884 (O_1884,N_49844,N_49890);
nand UO_1885 (O_1885,N_49876,N_49970);
nand UO_1886 (O_1886,N_49862,N_49934);
and UO_1887 (O_1887,N_49933,N_49887);
nor UO_1888 (O_1888,N_49959,N_49902);
and UO_1889 (O_1889,N_49844,N_49785);
nor UO_1890 (O_1890,N_49900,N_49764);
and UO_1891 (O_1891,N_49868,N_49913);
xnor UO_1892 (O_1892,N_49801,N_49892);
nor UO_1893 (O_1893,N_49867,N_49884);
and UO_1894 (O_1894,N_49920,N_49893);
nand UO_1895 (O_1895,N_49757,N_49889);
nand UO_1896 (O_1896,N_49982,N_49874);
nand UO_1897 (O_1897,N_49892,N_49783);
and UO_1898 (O_1898,N_49962,N_49837);
nand UO_1899 (O_1899,N_49910,N_49859);
and UO_1900 (O_1900,N_49772,N_49756);
or UO_1901 (O_1901,N_49808,N_49997);
and UO_1902 (O_1902,N_49873,N_49813);
nand UO_1903 (O_1903,N_49900,N_49996);
nor UO_1904 (O_1904,N_49775,N_49751);
and UO_1905 (O_1905,N_49783,N_49999);
nor UO_1906 (O_1906,N_49992,N_49753);
xor UO_1907 (O_1907,N_49789,N_49998);
nor UO_1908 (O_1908,N_49988,N_49808);
xor UO_1909 (O_1909,N_49964,N_49897);
or UO_1910 (O_1910,N_49959,N_49973);
and UO_1911 (O_1911,N_49921,N_49800);
nor UO_1912 (O_1912,N_49874,N_49875);
or UO_1913 (O_1913,N_49763,N_49964);
nand UO_1914 (O_1914,N_49872,N_49993);
nor UO_1915 (O_1915,N_49818,N_49955);
xor UO_1916 (O_1916,N_49841,N_49819);
and UO_1917 (O_1917,N_49777,N_49951);
nand UO_1918 (O_1918,N_49955,N_49860);
nand UO_1919 (O_1919,N_49754,N_49933);
xor UO_1920 (O_1920,N_49901,N_49959);
nor UO_1921 (O_1921,N_49932,N_49878);
or UO_1922 (O_1922,N_49942,N_49909);
xnor UO_1923 (O_1923,N_49751,N_49874);
and UO_1924 (O_1924,N_49893,N_49944);
nor UO_1925 (O_1925,N_49953,N_49866);
and UO_1926 (O_1926,N_49880,N_49795);
nand UO_1927 (O_1927,N_49929,N_49808);
nor UO_1928 (O_1928,N_49941,N_49750);
nand UO_1929 (O_1929,N_49989,N_49772);
or UO_1930 (O_1930,N_49784,N_49826);
and UO_1931 (O_1931,N_49902,N_49993);
or UO_1932 (O_1932,N_49763,N_49842);
nand UO_1933 (O_1933,N_49924,N_49870);
and UO_1934 (O_1934,N_49955,N_49949);
or UO_1935 (O_1935,N_49760,N_49807);
or UO_1936 (O_1936,N_49921,N_49990);
and UO_1937 (O_1937,N_49863,N_49761);
nor UO_1938 (O_1938,N_49792,N_49902);
nor UO_1939 (O_1939,N_49907,N_49821);
nor UO_1940 (O_1940,N_49895,N_49894);
xor UO_1941 (O_1941,N_49983,N_49988);
nand UO_1942 (O_1942,N_49869,N_49862);
nor UO_1943 (O_1943,N_49969,N_49832);
nor UO_1944 (O_1944,N_49901,N_49840);
or UO_1945 (O_1945,N_49877,N_49776);
xor UO_1946 (O_1946,N_49834,N_49751);
nand UO_1947 (O_1947,N_49983,N_49889);
nor UO_1948 (O_1948,N_49851,N_49889);
nand UO_1949 (O_1949,N_49897,N_49855);
or UO_1950 (O_1950,N_49930,N_49839);
and UO_1951 (O_1951,N_49860,N_49904);
nand UO_1952 (O_1952,N_49991,N_49812);
nand UO_1953 (O_1953,N_49925,N_49988);
or UO_1954 (O_1954,N_49779,N_49841);
or UO_1955 (O_1955,N_49928,N_49929);
nor UO_1956 (O_1956,N_49819,N_49968);
nand UO_1957 (O_1957,N_49940,N_49884);
or UO_1958 (O_1958,N_49985,N_49982);
and UO_1959 (O_1959,N_49798,N_49966);
nand UO_1960 (O_1960,N_49961,N_49831);
nand UO_1961 (O_1961,N_49830,N_49800);
nand UO_1962 (O_1962,N_49846,N_49884);
or UO_1963 (O_1963,N_49810,N_49797);
and UO_1964 (O_1964,N_49788,N_49794);
and UO_1965 (O_1965,N_49994,N_49812);
and UO_1966 (O_1966,N_49937,N_49898);
and UO_1967 (O_1967,N_49795,N_49842);
or UO_1968 (O_1968,N_49925,N_49890);
xor UO_1969 (O_1969,N_49913,N_49975);
and UO_1970 (O_1970,N_49844,N_49850);
nand UO_1971 (O_1971,N_49783,N_49762);
nand UO_1972 (O_1972,N_49983,N_49822);
nor UO_1973 (O_1973,N_49849,N_49968);
or UO_1974 (O_1974,N_49953,N_49767);
xnor UO_1975 (O_1975,N_49950,N_49802);
or UO_1976 (O_1976,N_49975,N_49926);
nand UO_1977 (O_1977,N_49819,N_49836);
or UO_1978 (O_1978,N_49784,N_49962);
nor UO_1979 (O_1979,N_49923,N_49910);
nand UO_1980 (O_1980,N_49980,N_49926);
nor UO_1981 (O_1981,N_49901,N_49971);
nor UO_1982 (O_1982,N_49867,N_49945);
nand UO_1983 (O_1983,N_49824,N_49788);
or UO_1984 (O_1984,N_49977,N_49897);
and UO_1985 (O_1985,N_49970,N_49777);
or UO_1986 (O_1986,N_49820,N_49856);
nand UO_1987 (O_1987,N_49998,N_49882);
nor UO_1988 (O_1988,N_49997,N_49838);
or UO_1989 (O_1989,N_49813,N_49786);
nor UO_1990 (O_1990,N_49939,N_49763);
nor UO_1991 (O_1991,N_49755,N_49831);
and UO_1992 (O_1992,N_49936,N_49866);
nor UO_1993 (O_1993,N_49778,N_49815);
and UO_1994 (O_1994,N_49795,N_49868);
and UO_1995 (O_1995,N_49867,N_49947);
xnor UO_1996 (O_1996,N_49866,N_49837);
nand UO_1997 (O_1997,N_49886,N_49828);
or UO_1998 (O_1998,N_49886,N_49843);
and UO_1999 (O_1999,N_49906,N_49933);
xnor UO_2000 (O_2000,N_49954,N_49839);
and UO_2001 (O_2001,N_49879,N_49790);
and UO_2002 (O_2002,N_49960,N_49847);
nor UO_2003 (O_2003,N_49807,N_49846);
and UO_2004 (O_2004,N_49980,N_49894);
nor UO_2005 (O_2005,N_49812,N_49874);
xor UO_2006 (O_2006,N_49868,N_49902);
nor UO_2007 (O_2007,N_49889,N_49812);
or UO_2008 (O_2008,N_49751,N_49839);
and UO_2009 (O_2009,N_49931,N_49824);
xnor UO_2010 (O_2010,N_49779,N_49888);
nand UO_2011 (O_2011,N_49802,N_49808);
nand UO_2012 (O_2012,N_49789,N_49898);
nor UO_2013 (O_2013,N_49795,N_49858);
xnor UO_2014 (O_2014,N_49904,N_49764);
and UO_2015 (O_2015,N_49833,N_49817);
nand UO_2016 (O_2016,N_49880,N_49813);
or UO_2017 (O_2017,N_49879,N_49922);
or UO_2018 (O_2018,N_49992,N_49910);
xor UO_2019 (O_2019,N_49916,N_49957);
nand UO_2020 (O_2020,N_49831,N_49821);
nand UO_2021 (O_2021,N_49926,N_49945);
or UO_2022 (O_2022,N_49882,N_49916);
or UO_2023 (O_2023,N_49924,N_49864);
and UO_2024 (O_2024,N_49984,N_49922);
nand UO_2025 (O_2025,N_49806,N_49772);
nor UO_2026 (O_2026,N_49802,N_49781);
or UO_2027 (O_2027,N_49881,N_49895);
xnor UO_2028 (O_2028,N_49757,N_49868);
and UO_2029 (O_2029,N_49814,N_49945);
nor UO_2030 (O_2030,N_49784,N_49786);
and UO_2031 (O_2031,N_49834,N_49784);
nand UO_2032 (O_2032,N_49919,N_49897);
nor UO_2033 (O_2033,N_49814,N_49979);
nand UO_2034 (O_2034,N_49979,N_49916);
and UO_2035 (O_2035,N_49772,N_49954);
xnor UO_2036 (O_2036,N_49904,N_49767);
and UO_2037 (O_2037,N_49928,N_49974);
or UO_2038 (O_2038,N_49903,N_49832);
and UO_2039 (O_2039,N_49771,N_49858);
nor UO_2040 (O_2040,N_49915,N_49986);
and UO_2041 (O_2041,N_49799,N_49936);
xnor UO_2042 (O_2042,N_49860,N_49899);
nand UO_2043 (O_2043,N_49883,N_49773);
xor UO_2044 (O_2044,N_49986,N_49923);
and UO_2045 (O_2045,N_49826,N_49903);
or UO_2046 (O_2046,N_49986,N_49811);
and UO_2047 (O_2047,N_49803,N_49764);
and UO_2048 (O_2048,N_49778,N_49848);
or UO_2049 (O_2049,N_49797,N_49978);
nand UO_2050 (O_2050,N_49862,N_49849);
nand UO_2051 (O_2051,N_49926,N_49785);
nand UO_2052 (O_2052,N_49943,N_49975);
and UO_2053 (O_2053,N_49985,N_49861);
and UO_2054 (O_2054,N_49808,N_49991);
nor UO_2055 (O_2055,N_49994,N_49765);
and UO_2056 (O_2056,N_49898,N_49925);
and UO_2057 (O_2057,N_49963,N_49959);
xnor UO_2058 (O_2058,N_49839,N_49993);
nor UO_2059 (O_2059,N_49948,N_49884);
nand UO_2060 (O_2060,N_49829,N_49996);
xnor UO_2061 (O_2061,N_49979,N_49856);
nor UO_2062 (O_2062,N_49824,N_49928);
nor UO_2063 (O_2063,N_49894,N_49972);
and UO_2064 (O_2064,N_49834,N_49969);
nand UO_2065 (O_2065,N_49869,N_49817);
nor UO_2066 (O_2066,N_49770,N_49958);
nand UO_2067 (O_2067,N_49754,N_49821);
nor UO_2068 (O_2068,N_49873,N_49910);
nand UO_2069 (O_2069,N_49912,N_49904);
nor UO_2070 (O_2070,N_49938,N_49765);
xnor UO_2071 (O_2071,N_49825,N_49918);
xnor UO_2072 (O_2072,N_49901,N_49767);
or UO_2073 (O_2073,N_49765,N_49851);
nor UO_2074 (O_2074,N_49818,N_49972);
xor UO_2075 (O_2075,N_49785,N_49757);
nand UO_2076 (O_2076,N_49816,N_49794);
and UO_2077 (O_2077,N_49986,N_49966);
and UO_2078 (O_2078,N_49827,N_49843);
and UO_2079 (O_2079,N_49826,N_49796);
and UO_2080 (O_2080,N_49849,N_49977);
nand UO_2081 (O_2081,N_49947,N_49888);
or UO_2082 (O_2082,N_49993,N_49999);
nor UO_2083 (O_2083,N_49784,N_49840);
and UO_2084 (O_2084,N_49765,N_49840);
and UO_2085 (O_2085,N_49782,N_49828);
or UO_2086 (O_2086,N_49763,N_49767);
xnor UO_2087 (O_2087,N_49895,N_49867);
or UO_2088 (O_2088,N_49936,N_49812);
nor UO_2089 (O_2089,N_49986,N_49823);
nand UO_2090 (O_2090,N_49985,N_49936);
nor UO_2091 (O_2091,N_49793,N_49770);
xnor UO_2092 (O_2092,N_49890,N_49961);
nor UO_2093 (O_2093,N_49849,N_49987);
and UO_2094 (O_2094,N_49846,N_49949);
nand UO_2095 (O_2095,N_49993,N_49774);
or UO_2096 (O_2096,N_49918,N_49849);
nand UO_2097 (O_2097,N_49932,N_49914);
xnor UO_2098 (O_2098,N_49819,N_49831);
nand UO_2099 (O_2099,N_49796,N_49762);
nand UO_2100 (O_2100,N_49821,N_49876);
and UO_2101 (O_2101,N_49985,N_49954);
nor UO_2102 (O_2102,N_49842,N_49961);
xnor UO_2103 (O_2103,N_49834,N_49968);
or UO_2104 (O_2104,N_49814,N_49824);
xnor UO_2105 (O_2105,N_49987,N_49811);
and UO_2106 (O_2106,N_49853,N_49898);
nand UO_2107 (O_2107,N_49852,N_49760);
nand UO_2108 (O_2108,N_49855,N_49895);
or UO_2109 (O_2109,N_49778,N_49803);
nor UO_2110 (O_2110,N_49794,N_49885);
or UO_2111 (O_2111,N_49872,N_49886);
nand UO_2112 (O_2112,N_49894,N_49908);
and UO_2113 (O_2113,N_49980,N_49948);
nor UO_2114 (O_2114,N_49896,N_49796);
and UO_2115 (O_2115,N_49993,N_49825);
nand UO_2116 (O_2116,N_49933,N_49763);
nand UO_2117 (O_2117,N_49940,N_49791);
nor UO_2118 (O_2118,N_49934,N_49825);
or UO_2119 (O_2119,N_49949,N_49988);
and UO_2120 (O_2120,N_49896,N_49878);
or UO_2121 (O_2121,N_49914,N_49987);
and UO_2122 (O_2122,N_49954,N_49995);
xnor UO_2123 (O_2123,N_49915,N_49770);
xor UO_2124 (O_2124,N_49836,N_49835);
xor UO_2125 (O_2125,N_49902,N_49862);
nand UO_2126 (O_2126,N_49885,N_49932);
and UO_2127 (O_2127,N_49881,N_49978);
nor UO_2128 (O_2128,N_49989,N_49793);
or UO_2129 (O_2129,N_49776,N_49798);
or UO_2130 (O_2130,N_49962,N_49773);
nor UO_2131 (O_2131,N_49822,N_49780);
nor UO_2132 (O_2132,N_49850,N_49974);
xor UO_2133 (O_2133,N_49877,N_49993);
and UO_2134 (O_2134,N_49752,N_49974);
and UO_2135 (O_2135,N_49891,N_49929);
nand UO_2136 (O_2136,N_49990,N_49856);
and UO_2137 (O_2137,N_49903,N_49802);
or UO_2138 (O_2138,N_49786,N_49974);
nand UO_2139 (O_2139,N_49816,N_49833);
xnor UO_2140 (O_2140,N_49819,N_49872);
nand UO_2141 (O_2141,N_49809,N_49831);
nand UO_2142 (O_2142,N_49808,N_49920);
and UO_2143 (O_2143,N_49872,N_49756);
and UO_2144 (O_2144,N_49806,N_49995);
and UO_2145 (O_2145,N_49981,N_49877);
or UO_2146 (O_2146,N_49949,N_49899);
and UO_2147 (O_2147,N_49916,N_49872);
or UO_2148 (O_2148,N_49915,N_49882);
xnor UO_2149 (O_2149,N_49866,N_49797);
and UO_2150 (O_2150,N_49837,N_49800);
xnor UO_2151 (O_2151,N_49806,N_49804);
and UO_2152 (O_2152,N_49869,N_49763);
nor UO_2153 (O_2153,N_49836,N_49928);
nand UO_2154 (O_2154,N_49919,N_49868);
nor UO_2155 (O_2155,N_49927,N_49884);
or UO_2156 (O_2156,N_49828,N_49788);
nand UO_2157 (O_2157,N_49913,N_49760);
xor UO_2158 (O_2158,N_49806,N_49989);
and UO_2159 (O_2159,N_49972,N_49969);
nand UO_2160 (O_2160,N_49957,N_49774);
and UO_2161 (O_2161,N_49827,N_49857);
nor UO_2162 (O_2162,N_49939,N_49903);
and UO_2163 (O_2163,N_49756,N_49867);
or UO_2164 (O_2164,N_49885,N_49816);
or UO_2165 (O_2165,N_49873,N_49934);
xnor UO_2166 (O_2166,N_49778,N_49861);
nor UO_2167 (O_2167,N_49781,N_49834);
nand UO_2168 (O_2168,N_49997,N_49929);
or UO_2169 (O_2169,N_49759,N_49899);
xor UO_2170 (O_2170,N_49915,N_49802);
nand UO_2171 (O_2171,N_49955,N_49787);
and UO_2172 (O_2172,N_49762,N_49804);
nor UO_2173 (O_2173,N_49755,N_49911);
nor UO_2174 (O_2174,N_49932,N_49969);
nand UO_2175 (O_2175,N_49921,N_49979);
nand UO_2176 (O_2176,N_49859,N_49825);
nand UO_2177 (O_2177,N_49994,N_49888);
nor UO_2178 (O_2178,N_49991,N_49852);
xnor UO_2179 (O_2179,N_49944,N_49867);
xnor UO_2180 (O_2180,N_49880,N_49929);
xnor UO_2181 (O_2181,N_49835,N_49811);
nor UO_2182 (O_2182,N_49789,N_49993);
xnor UO_2183 (O_2183,N_49869,N_49967);
and UO_2184 (O_2184,N_49966,N_49971);
or UO_2185 (O_2185,N_49811,N_49871);
nand UO_2186 (O_2186,N_49892,N_49898);
nand UO_2187 (O_2187,N_49946,N_49841);
and UO_2188 (O_2188,N_49943,N_49766);
and UO_2189 (O_2189,N_49838,N_49923);
nor UO_2190 (O_2190,N_49949,N_49902);
and UO_2191 (O_2191,N_49939,N_49816);
nor UO_2192 (O_2192,N_49835,N_49917);
or UO_2193 (O_2193,N_49895,N_49774);
nor UO_2194 (O_2194,N_49787,N_49936);
nand UO_2195 (O_2195,N_49806,N_49836);
and UO_2196 (O_2196,N_49948,N_49949);
or UO_2197 (O_2197,N_49882,N_49908);
nor UO_2198 (O_2198,N_49964,N_49923);
nor UO_2199 (O_2199,N_49928,N_49803);
or UO_2200 (O_2200,N_49775,N_49896);
or UO_2201 (O_2201,N_49945,N_49921);
nor UO_2202 (O_2202,N_49878,N_49780);
and UO_2203 (O_2203,N_49832,N_49917);
and UO_2204 (O_2204,N_49771,N_49854);
xor UO_2205 (O_2205,N_49788,N_49800);
nor UO_2206 (O_2206,N_49962,N_49994);
nor UO_2207 (O_2207,N_49801,N_49843);
nor UO_2208 (O_2208,N_49855,N_49959);
xor UO_2209 (O_2209,N_49822,N_49924);
nand UO_2210 (O_2210,N_49836,N_49902);
and UO_2211 (O_2211,N_49818,N_49854);
nand UO_2212 (O_2212,N_49908,N_49926);
or UO_2213 (O_2213,N_49805,N_49797);
nand UO_2214 (O_2214,N_49811,N_49827);
nand UO_2215 (O_2215,N_49778,N_49867);
or UO_2216 (O_2216,N_49807,N_49786);
and UO_2217 (O_2217,N_49844,N_49984);
or UO_2218 (O_2218,N_49831,N_49915);
nand UO_2219 (O_2219,N_49991,N_49870);
xor UO_2220 (O_2220,N_49878,N_49977);
and UO_2221 (O_2221,N_49985,N_49780);
and UO_2222 (O_2222,N_49858,N_49922);
nor UO_2223 (O_2223,N_49983,N_49816);
nand UO_2224 (O_2224,N_49906,N_49779);
and UO_2225 (O_2225,N_49989,N_49792);
and UO_2226 (O_2226,N_49790,N_49857);
xnor UO_2227 (O_2227,N_49878,N_49888);
and UO_2228 (O_2228,N_49849,N_49780);
xor UO_2229 (O_2229,N_49899,N_49870);
or UO_2230 (O_2230,N_49860,N_49943);
or UO_2231 (O_2231,N_49837,N_49765);
or UO_2232 (O_2232,N_49994,N_49958);
or UO_2233 (O_2233,N_49962,N_49966);
xor UO_2234 (O_2234,N_49817,N_49805);
nor UO_2235 (O_2235,N_49830,N_49810);
or UO_2236 (O_2236,N_49907,N_49882);
and UO_2237 (O_2237,N_49994,N_49990);
and UO_2238 (O_2238,N_49791,N_49892);
or UO_2239 (O_2239,N_49899,N_49878);
nand UO_2240 (O_2240,N_49991,N_49871);
or UO_2241 (O_2241,N_49926,N_49758);
nand UO_2242 (O_2242,N_49963,N_49826);
xnor UO_2243 (O_2243,N_49753,N_49845);
and UO_2244 (O_2244,N_49836,N_49863);
nand UO_2245 (O_2245,N_49874,N_49802);
or UO_2246 (O_2246,N_49989,N_49874);
and UO_2247 (O_2247,N_49822,N_49834);
nand UO_2248 (O_2248,N_49962,N_49892);
nor UO_2249 (O_2249,N_49980,N_49867);
xor UO_2250 (O_2250,N_49796,N_49906);
and UO_2251 (O_2251,N_49751,N_49771);
xor UO_2252 (O_2252,N_49869,N_49932);
and UO_2253 (O_2253,N_49778,N_49851);
nand UO_2254 (O_2254,N_49774,N_49858);
xor UO_2255 (O_2255,N_49798,N_49844);
nor UO_2256 (O_2256,N_49999,N_49802);
or UO_2257 (O_2257,N_49876,N_49795);
or UO_2258 (O_2258,N_49760,N_49829);
nand UO_2259 (O_2259,N_49861,N_49981);
or UO_2260 (O_2260,N_49975,N_49952);
xor UO_2261 (O_2261,N_49887,N_49823);
nor UO_2262 (O_2262,N_49770,N_49801);
and UO_2263 (O_2263,N_49937,N_49874);
xnor UO_2264 (O_2264,N_49992,N_49755);
nand UO_2265 (O_2265,N_49998,N_49902);
xnor UO_2266 (O_2266,N_49906,N_49955);
or UO_2267 (O_2267,N_49994,N_49979);
and UO_2268 (O_2268,N_49927,N_49942);
xor UO_2269 (O_2269,N_49765,N_49828);
nor UO_2270 (O_2270,N_49832,N_49759);
xor UO_2271 (O_2271,N_49993,N_49868);
nand UO_2272 (O_2272,N_49993,N_49917);
or UO_2273 (O_2273,N_49989,N_49809);
and UO_2274 (O_2274,N_49899,N_49757);
nor UO_2275 (O_2275,N_49828,N_49799);
and UO_2276 (O_2276,N_49764,N_49847);
xnor UO_2277 (O_2277,N_49869,N_49877);
xnor UO_2278 (O_2278,N_49870,N_49939);
or UO_2279 (O_2279,N_49839,N_49848);
or UO_2280 (O_2280,N_49941,N_49760);
xnor UO_2281 (O_2281,N_49792,N_49819);
nor UO_2282 (O_2282,N_49891,N_49753);
and UO_2283 (O_2283,N_49812,N_49802);
xnor UO_2284 (O_2284,N_49791,N_49847);
and UO_2285 (O_2285,N_49849,N_49875);
or UO_2286 (O_2286,N_49865,N_49985);
and UO_2287 (O_2287,N_49842,N_49934);
xnor UO_2288 (O_2288,N_49811,N_49886);
xor UO_2289 (O_2289,N_49861,N_49963);
nor UO_2290 (O_2290,N_49933,N_49799);
and UO_2291 (O_2291,N_49810,N_49845);
xnor UO_2292 (O_2292,N_49922,N_49823);
xor UO_2293 (O_2293,N_49794,N_49983);
nor UO_2294 (O_2294,N_49997,N_49869);
nor UO_2295 (O_2295,N_49947,N_49789);
xnor UO_2296 (O_2296,N_49914,N_49971);
and UO_2297 (O_2297,N_49988,N_49930);
nor UO_2298 (O_2298,N_49890,N_49936);
nor UO_2299 (O_2299,N_49980,N_49970);
or UO_2300 (O_2300,N_49981,N_49958);
xor UO_2301 (O_2301,N_49986,N_49848);
nor UO_2302 (O_2302,N_49943,N_49952);
or UO_2303 (O_2303,N_49778,N_49750);
nor UO_2304 (O_2304,N_49898,N_49955);
nand UO_2305 (O_2305,N_49865,N_49829);
xor UO_2306 (O_2306,N_49954,N_49987);
or UO_2307 (O_2307,N_49876,N_49834);
nand UO_2308 (O_2308,N_49975,N_49974);
and UO_2309 (O_2309,N_49997,N_49792);
nor UO_2310 (O_2310,N_49950,N_49869);
nand UO_2311 (O_2311,N_49993,N_49760);
xor UO_2312 (O_2312,N_49919,N_49870);
nand UO_2313 (O_2313,N_49920,N_49897);
or UO_2314 (O_2314,N_49873,N_49816);
nor UO_2315 (O_2315,N_49974,N_49900);
or UO_2316 (O_2316,N_49913,N_49807);
nand UO_2317 (O_2317,N_49908,N_49992);
xnor UO_2318 (O_2318,N_49803,N_49755);
nor UO_2319 (O_2319,N_49766,N_49936);
or UO_2320 (O_2320,N_49883,N_49980);
xnor UO_2321 (O_2321,N_49770,N_49844);
or UO_2322 (O_2322,N_49820,N_49847);
and UO_2323 (O_2323,N_49792,N_49959);
or UO_2324 (O_2324,N_49933,N_49843);
nand UO_2325 (O_2325,N_49924,N_49884);
or UO_2326 (O_2326,N_49767,N_49898);
and UO_2327 (O_2327,N_49992,N_49776);
nand UO_2328 (O_2328,N_49836,N_49936);
nor UO_2329 (O_2329,N_49787,N_49937);
and UO_2330 (O_2330,N_49875,N_49990);
nand UO_2331 (O_2331,N_49963,N_49920);
xor UO_2332 (O_2332,N_49976,N_49945);
nand UO_2333 (O_2333,N_49765,N_49774);
nor UO_2334 (O_2334,N_49978,N_49798);
xnor UO_2335 (O_2335,N_49839,N_49864);
and UO_2336 (O_2336,N_49907,N_49810);
or UO_2337 (O_2337,N_49899,N_49850);
nand UO_2338 (O_2338,N_49845,N_49881);
and UO_2339 (O_2339,N_49801,N_49973);
nand UO_2340 (O_2340,N_49900,N_49775);
xnor UO_2341 (O_2341,N_49751,N_49913);
and UO_2342 (O_2342,N_49852,N_49759);
nor UO_2343 (O_2343,N_49926,N_49887);
or UO_2344 (O_2344,N_49794,N_49963);
nor UO_2345 (O_2345,N_49755,N_49890);
and UO_2346 (O_2346,N_49843,N_49810);
or UO_2347 (O_2347,N_49795,N_49972);
xnor UO_2348 (O_2348,N_49846,N_49792);
or UO_2349 (O_2349,N_49823,N_49839);
nand UO_2350 (O_2350,N_49784,N_49961);
and UO_2351 (O_2351,N_49977,N_49850);
nand UO_2352 (O_2352,N_49784,N_49841);
nand UO_2353 (O_2353,N_49930,N_49934);
nand UO_2354 (O_2354,N_49785,N_49783);
or UO_2355 (O_2355,N_49764,N_49988);
nand UO_2356 (O_2356,N_49778,N_49857);
or UO_2357 (O_2357,N_49894,N_49882);
nand UO_2358 (O_2358,N_49778,N_49817);
nor UO_2359 (O_2359,N_49958,N_49767);
xnor UO_2360 (O_2360,N_49846,N_49838);
nand UO_2361 (O_2361,N_49901,N_49860);
or UO_2362 (O_2362,N_49794,N_49801);
xor UO_2363 (O_2363,N_49999,N_49767);
and UO_2364 (O_2364,N_49851,N_49827);
or UO_2365 (O_2365,N_49813,N_49996);
and UO_2366 (O_2366,N_49881,N_49790);
and UO_2367 (O_2367,N_49910,N_49842);
xnor UO_2368 (O_2368,N_49843,N_49852);
nor UO_2369 (O_2369,N_49957,N_49939);
and UO_2370 (O_2370,N_49830,N_49888);
and UO_2371 (O_2371,N_49924,N_49968);
or UO_2372 (O_2372,N_49894,N_49830);
or UO_2373 (O_2373,N_49937,N_49843);
and UO_2374 (O_2374,N_49892,N_49958);
or UO_2375 (O_2375,N_49846,N_49911);
or UO_2376 (O_2376,N_49870,N_49796);
nand UO_2377 (O_2377,N_49909,N_49974);
or UO_2378 (O_2378,N_49854,N_49767);
xor UO_2379 (O_2379,N_49795,N_49819);
or UO_2380 (O_2380,N_49790,N_49832);
nand UO_2381 (O_2381,N_49982,N_49912);
nor UO_2382 (O_2382,N_49752,N_49824);
nor UO_2383 (O_2383,N_49947,N_49771);
xor UO_2384 (O_2384,N_49941,N_49938);
nand UO_2385 (O_2385,N_49852,N_49918);
or UO_2386 (O_2386,N_49783,N_49889);
nand UO_2387 (O_2387,N_49824,N_49864);
nor UO_2388 (O_2388,N_49885,N_49915);
nor UO_2389 (O_2389,N_49954,N_49779);
nor UO_2390 (O_2390,N_49792,N_49914);
nand UO_2391 (O_2391,N_49892,N_49838);
or UO_2392 (O_2392,N_49928,N_49844);
and UO_2393 (O_2393,N_49777,N_49932);
xor UO_2394 (O_2394,N_49789,N_49980);
or UO_2395 (O_2395,N_49900,N_49851);
or UO_2396 (O_2396,N_49789,N_49857);
and UO_2397 (O_2397,N_49961,N_49764);
and UO_2398 (O_2398,N_49788,N_49950);
nor UO_2399 (O_2399,N_49775,N_49886);
nand UO_2400 (O_2400,N_49869,N_49853);
nand UO_2401 (O_2401,N_49898,N_49908);
nor UO_2402 (O_2402,N_49996,N_49796);
nor UO_2403 (O_2403,N_49940,N_49960);
nand UO_2404 (O_2404,N_49803,N_49931);
or UO_2405 (O_2405,N_49945,N_49972);
or UO_2406 (O_2406,N_49949,N_49867);
or UO_2407 (O_2407,N_49751,N_49768);
nor UO_2408 (O_2408,N_49770,N_49894);
nand UO_2409 (O_2409,N_49883,N_49817);
or UO_2410 (O_2410,N_49883,N_49936);
and UO_2411 (O_2411,N_49775,N_49792);
xnor UO_2412 (O_2412,N_49790,N_49873);
or UO_2413 (O_2413,N_49862,N_49766);
or UO_2414 (O_2414,N_49811,N_49778);
nand UO_2415 (O_2415,N_49766,N_49764);
or UO_2416 (O_2416,N_49816,N_49897);
or UO_2417 (O_2417,N_49971,N_49861);
and UO_2418 (O_2418,N_49781,N_49965);
or UO_2419 (O_2419,N_49997,N_49816);
nor UO_2420 (O_2420,N_49792,N_49768);
and UO_2421 (O_2421,N_49883,N_49903);
and UO_2422 (O_2422,N_49780,N_49854);
xor UO_2423 (O_2423,N_49949,N_49910);
xnor UO_2424 (O_2424,N_49761,N_49860);
nor UO_2425 (O_2425,N_49887,N_49946);
and UO_2426 (O_2426,N_49762,N_49870);
or UO_2427 (O_2427,N_49911,N_49932);
nand UO_2428 (O_2428,N_49787,N_49897);
and UO_2429 (O_2429,N_49868,N_49753);
nor UO_2430 (O_2430,N_49777,N_49963);
or UO_2431 (O_2431,N_49949,N_49885);
or UO_2432 (O_2432,N_49907,N_49761);
or UO_2433 (O_2433,N_49777,N_49941);
xor UO_2434 (O_2434,N_49832,N_49787);
and UO_2435 (O_2435,N_49890,N_49800);
or UO_2436 (O_2436,N_49846,N_49915);
nand UO_2437 (O_2437,N_49790,N_49973);
or UO_2438 (O_2438,N_49908,N_49797);
xnor UO_2439 (O_2439,N_49804,N_49789);
nand UO_2440 (O_2440,N_49758,N_49897);
xnor UO_2441 (O_2441,N_49833,N_49914);
nand UO_2442 (O_2442,N_49758,N_49757);
or UO_2443 (O_2443,N_49936,N_49784);
and UO_2444 (O_2444,N_49774,N_49949);
and UO_2445 (O_2445,N_49874,N_49825);
nand UO_2446 (O_2446,N_49812,N_49984);
and UO_2447 (O_2447,N_49799,N_49923);
or UO_2448 (O_2448,N_49809,N_49793);
nor UO_2449 (O_2449,N_49775,N_49979);
nor UO_2450 (O_2450,N_49753,N_49949);
nand UO_2451 (O_2451,N_49883,N_49857);
xor UO_2452 (O_2452,N_49934,N_49983);
nor UO_2453 (O_2453,N_49826,N_49942);
xnor UO_2454 (O_2454,N_49991,N_49923);
or UO_2455 (O_2455,N_49840,N_49754);
nor UO_2456 (O_2456,N_49849,N_49985);
xor UO_2457 (O_2457,N_49794,N_49807);
nor UO_2458 (O_2458,N_49844,N_49967);
nor UO_2459 (O_2459,N_49894,N_49927);
or UO_2460 (O_2460,N_49936,N_49864);
and UO_2461 (O_2461,N_49908,N_49978);
and UO_2462 (O_2462,N_49954,N_49913);
nor UO_2463 (O_2463,N_49932,N_49988);
or UO_2464 (O_2464,N_49873,N_49917);
nor UO_2465 (O_2465,N_49939,N_49783);
or UO_2466 (O_2466,N_49973,N_49812);
or UO_2467 (O_2467,N_49837,N_49787);
or UO_2468 (O_2468,N_49831,N_49941);
and UO_2469 (O_2469,N_49883,N_49924);
nand UO_2470 (O_2470,N_49899,N_49911);
and UO_2471 (O_2471,N_49843,N_49791);
nor UO_2472 (O_2472,N_49854,N_49930);
nand UO_2473 (O_2473,N_49929,N_49778);
or UO_2474 (O_2474,N_49834,N_49915);
nor UO_2475 (O_2475,N_49869,N_49772);
xnor UO_2476 (O_2476,N_49880,N_49780);
nand UO_2477 (O_2477,N_49824,N_49998);
and UO_2478 (O_2478,N_49913,N_49908);
nand UO_2479 (O_2479,N_49848,N_49896);
and UO_2480 (O_2480,N_49859,N_49811);
nand UO_2481 (O_2481,N_49755,N_49939);
xnor UO_2482 (O_2482,N_49821,N_49909);
or UO_2483 (O_2483,N_49901,N_49939);
or UO_2484 (O_2484,N_49911,N_49854);
or UO_2485 (O_2485,N_49963,N_49908);
and UO_2486 (O_2486,N_49758,N_49940);
xnor UO_2487 (O_2487,N_49808,N_49902);
or UO_2488 (O_2488,N_49954,N_49957);
and UO_2489 (O_2489,N_49793,N_49764);
nor UO_2490 (O_2490,N_49838,N_49842);
xnor UO_2491 (O_2491,N_49878,N_49777);
xnor UO_2492 (O_2492,N_49904,N_49984);
and UO_2493 (O_2493,N_49828,N_49944);
and UO_2494 (O_2494,N_49884,N_49804);
nand UO_2495 (O_2495,N_49960,N_49957);
or UO_2496 (O_2496,N_49768,N_49843);
and UO_2497 (O_2497,N_49791,N_49758);
xor UO_2498 (O_2498,N_49788,N_49906);
xor UO_2499 (O_2499,N_49879,N_49951);
and UO_2500 (O_2500,N_49852,N_49959);
xnor UO_2501 (O_2501,N_49773,N_49811);
and UO_2502 (O_2502,N_49977,N_49991);
and UO_2503 (O_2503,N_49870,N_49920);
and UO_2504 (O_2504,N_49933,N_49816);
nor UO_2505 (O_2505,N_49891,N_49802);
or UO_2506 (O_2506,N_49958,N_49912);
xor UO_2507 (O_2507,N_49800,N_49977);
nor UO_2508 (O_2508,N_49794,N_49861);
or UO_2509 (O_2509,N_49823,N_49998);
nor UO_2510 (O_2510,N_49848,N_49893);
or UO_2511 (O_2511,N_49924,N_49940);
xnor UO_2512 (O_2512,N_49848,N_49789);
nor UO_2513 (O_2513,N_49881,N_49802);
or UO_2514 (O_2514,N_49928,N_49886);
and UO_2515 (O_2515,N_49842,N_49885);
and UO_2516 (O_2516,N_49866,N_49863);
nor UO_2517 (O_2517,N_49977,N_49771);
and UO_2518 (O_2518,N_49797,N_49796);
xor UO_2519 (O_2519,N_49791,N_49907);
nand UO_2520 (O_2520,N_49971,N_49988);
or UO_2521 (O_2521,N_49902,N_49923);
nand UO_2522 (O_2522,N_49833,N_49754);
xnor UO_2523 (O_2523,N_49981,N_49964);
xnor UO_2524 (O_2524,N_49950,N_49813);
nand UO_2525 (O_2525,N_49751,N_49830);
nor UO_2526 (O_2526,N_49874,N_49938);
or UO_2527 (O_2527,N_49833,N_49786);
and UO_2528 (O_2528,N_49956,N_49779);
and UO_2529 (O_2529,N_49911,N_49769);
nand UO_2530 (O_2530,N_49754,N_49964);
or UO_2531 (O_2531,N_49805,N_49950);
xor UO_2532 (O_2532,N_49932,N_49882);
nor UO_2533 (O_2533,N_49997,N_49794);
and UO_2534 (O_2534,N_49946,N_49912);
and UO_2535 (O_2535,N_49846,N_49865);
nand UO_2536 (O_2536,N_49788,N_49940);
xor UO_2537 (O_2537,N_49989,N_49750);
or UO_2538 (O_2538,N_49768,N_49887);
nand UO_2539 (O_2539,N_49869,N_49786);
nand UO_2540 (O_2540,N_49784,N_49852);
xnor UO_2541 (O_2541,N_49969,N_49875);
nand UO_2542 (O_2542,N_49795,N_49918);
nand UO_2543 (O_2543,N_49836,N_49999);
nor UO_2544 (O_2544,N_49788,N_49979);
nor UO_2545 (O_2545,N_49804,N_49951);
nand UO_2546 (O_2546,N_49927,N_49943);
nor UO_2547 (O_2547,N_49982,N_49940);
and UO_2548 (O_2548,N_49759,N_49934);
nor UO_2549 (O_2549,N_49826,N_49974);
and UO_2550 (O_2550,N_49884,N_49772);
or UO_2551 (O_2551,N_49974,N_49945);
nor UO_2552 (O_2552,N_49893,N_49817);
nor UO_2553 (O_2553,N_49830,N_49760);
or UO_2554 (O_2554,N_49890,N_49856);
or UO_2555 (O_2555,N_49830,N_49891);
nor UO_2556 (O_2556,N_49930,N_49970);
or UO_2557 (O_2557,N_49759,N_49869);
nor UO_2558 (O_2558,N_49977,N_49790);
xor UO_2559 (O_2559,N_49774,N_49924);
xor UO_2560 (O_2560,N_49924,N_49777);
xor UO_2561 (O_2561,N_49825,N_49917);
and UO_2562 (O_2562,N_49777,N_49989);
and UO_2563 (O_2563,N_49877,N_49930);
or UO_2564 (O_2564,N_49829,N_49939);
or UO_2565 (O_2565,N_49807,N_49988);
xor UO_2566 (O_2566,N_49799,N_49812);
xor UO_2567 (O_2567,N_49888,N_49824);
nand UO_2568 (O_2568,N_49995,N_49819);
and UO_2569 (O_2569,N_49844,N_49791);
and UO_2570 (O_2570,N_49849,N_49830);
or UO_2571 (O_2571,N_49870,N_49905);
nor UO_2572 (O_2572,N_49965,N_49896);
nand UO_2573 (O_2573,N_49969,N_49967);
nand UO_2574 (O_2574,N_49757,N_49986);
nand UO_2575 (O_2575,N_49946,N_49929);
nor UO_2576 (O_2576,N_49786,N_49994);
or UO_2577 (O_2577,N_49990,N_49964);
nand UO_2578 (O_2578,N_49758,N_49882);
or UO_2579 (O_2579,N_49853,N_49988);
nor UO_2580 (O_2580,N_49967,N_49995);
nand UO_2581 (O_2581,N_49828,N_49906);
nand UO_2582 (O_2582,N_49802,N_49857);
and UO_2583 (O_2583,N_49757,N_49990);
xor UO_2584 (O_2584,N_49801,N_49927);
or UO_2585 (O_2585,N_49761,N_49830);
or UO_2586 (O_2586,N_49813,N_49799);
nand UO_2587 (O_2587,N_49853,N_49817);
nand UO_2588 (O_2588,N_49767,N_49858);
xnor UO_2589 (O_2589,N_49851,N_49773);
nor UO_2590 (O_2590,N_49862,N_49914);
nand UO_2591 (O_2591,N_49796,N_49862);
xnor UO_2592 (O_2592,N_49944,N_49821);
and UO_2593 (O_2593,N_49943,N_49892);
nand UO_2594 (O_2594,N_49954,N_49947);
nor UO_2595 (O_2595,N_49884,N_49796);
nand UO_2596 (O_2596,N_49830,N_49998);
nor UO_2597 (O_2597,N_49799,N_49969);
and UO_2598 (O_2598,N_49757,N_49979);
and UO_2599 (O_2599,N_49842,N_49817);
nor UO_2600 (O_2600,N_49814,N_49912);
nand UO_2601 (O_2601,N_49857,N_49806);
or UO_2602 (O_2602,N_49979,N_49849);
nand UO_2603 (O_2603,N_49805,N_49946);
nor UO_2604 (O_2604,N_49846,N_49918);
xor UO_2605 (O_2605,N_49768,N_49920);
nand UO_2606 (O_2606,N_49844,N_49794);
or UO_2607 (O_2607,N_49756,N_49826);
and UO_2608 (O_2608,N_49965,N_49766);
and UO_2609 (O_2609,N_49881,N_49922);
nor UO_2610 (O_2610,N_49840,N_49758);
nor UO_2611 (O_2611,N_49966,N_49972);
and UO_2612 (O_2612,N_49944,N_49989);
and UO_2613 (O_2613,N_49757,N_49938);
or UO_2614 (O_2614,N_49779,N_49988);
nor UO_2615 (O_2615,N_49856,N_49755);
or UO_2616 (O_2616,N_49921,N_49929);
and UO_2617 (O_2617,N_49976,N_49785);
nor UO_2618 (O_2618,N_49760,N_49827);
xor UO_2619 (O_2619,N_49812,N_49941);
or UO_2620 (O_2620,N_49917,N_49817);
and UO_2621 (O_2621,N_49796,N_49872);
nor UO_2622 (O_2622,N_49856,N_49767);
nand UO_2623 (O_2623,N_49822,N_49906);
nor UO_2624 (O_2624,N_49750,N_49966);
or UO_2625 (O_2625,N_49889,N_49810);
and UO_2626 (O_2626,N_49996,N_49977);
xnor UO_2627 (O_2627,N_49823,N_49849);
and UO_2628 (O_2628,N_49966,N_49793);
nand UO_2629 (O_2629,N_49937,N_49882);
and UO_2630 (O_2630,N_49962,N_49926);
nand UO_2631 (O_2631,N_49993,N_49829);
xor UO_2632 (O_2632,N_49794,N_49786);
nand UO_2633 (O_2633,N_49793,N_49810);
nand UO_2634 (O_2634,N_49810,N_49865);
and UO_2635 (O_2635,N_49818,N_49843);
and UO_2636 (O_2636,N_49799,N_49769);
and UO_2637 (O_2637,N_49906,N_49801);
or UO_2638 (O_2638,N_49836,N_49791);
xnor UO_2639 (O_2639,N_49964,N_49898);
and UO_2640 (O_2640,N_49870,N_49843);
xor UO_2641 (O_2641,N_49830,N_49813);
or UO_2642 (O_2642,N_49928,N_49782);
or UO_2643 (O_2643,N_49919,N_49937);
and UO_2644 (O_2644,N_49781,N_49839);
xor UO_2645 (O_2645,N_49923,N_49791);
xnor UO_2646 (O_2646,N_49870,N_49889);
nand UO_2647 (O_2647,N_49963,N_49887);
or UO_2648 (O_2648,N_49875,N_49911);
nand UO_2649 (O_2649,N_49933,N_49764);
nor UO_2650 (O_2650,N_49885,N_49826);
xnor UO_2651 (O_2651,N_49753,N_49865);
nand UO_2652 (O_2652,N_49806,N_49876);
nand UO_2653 (O_2653,N_49998,N_49857);
or UO_2654 (O_2654,N_49754,N_49844);
and UO_2655 (O_2655,N_49778,N_49988);
or UO_2656 (O_2656,N_49999,N_49780);
nor UO_2657 (O_2657,N_49829,N_49781);
nor UO_2658 (O_2658,N_49872,N_49894);
and UO_2659 (O_2659,N_49995,N_49870);
nand UO_2660 (O_2660,N_49892,N_49764);
nand UO_2661 (O_2661,N_49889,N_49880);
xnor UO_2662 (O_2662,N_49771,N_49936);
and UO_2663 (O_2663,N_49769,N_49804);
xor UO_2664 (O_2664,N_49883,N_49869);
nand UO_2665 (O_2665,N_49980,N_49914);
or UO_2666 (O_2666,N_49933,N_49893);
nand UO_2667 (O_2667,N_49859,N_49955);
nand UO_2668 (O_2668,N_49768,N_49764);
nor UO_2669 (O_2669,N_49767,N_49786);
and UO_2670 (O_2670,N_49841,N_49901);
and UO_2671 (O_2671,N_49755,N_49839);
nor UO_2672 (O_2672,N_49841,N_49975);
or UO_2673 (O_2673,N_49821,N_49800);
and UO_2674 (O_2674,N_49857,N_49852);
nand UO_2675 (O_2675,N_49917,N_49961);
nand UO_2676 (O_2676,N_49976,N_49862);
nand UO_2677 (O_2677,N_49923,N_49833);
or UO_2678 (O_2678,N_49849,N_49922);
and UO_2679 (O_2679,N_49818,N_49994);
nand UO_2680 (O_2680,N_49958,N_49990);
xor UO_2681 (O_2681,N_49914,N_49876);
nand UO_2682 (O_2682,N_49751,N_49902);
or UO_2683 (O_2683,N_49954,N_49753);
nor UO_2684 (O_2684,N_49953,N_49872);
nand UO_2685 (O_2685,N_49777,N_49860);
and UO_2686 (O_2686,N_49959,N_49878);
xor UO_2687 (O_2687,N_49874,N_49902);
nand UO_2688 (O_2688,N_49986,N_49854);
nand UO_2689 (O_2689,N_49774,N_49982);
xor UO_2690 (O_2690,N_49976,N_49787);
nand UO_2691 (O_2691,N_49912,N_49887);
or UO_2692 (O_2692,N_49808,N_49896);
nor UO_2693 (O_2693,N_49839,N_49929);
or UO_2694 (O_2694,N_49894,N_49925);
xor UO_2695 (O_2695,N_49951,N_49989);
or UO_2696 (O_2696,N_49809,N_49879);
nand UO_2697 (O_2697,N_49750,N_49984);
xnor UO_2698 (O_2698,N_49790,N_49860);
nor UO_2699 (O_2699,N_49970,N_49805);
and UO_2700 (O_2700,N_49779,N_49824);
xor UO_2701 (O_2701,N_49992,N_49835);
nor UO_2702 (O_2702,N_49898,N_49906);
nand UO_2703 (O_2703,N_49900,N_49928);
xor UO_2704 (O_2704,N_49781,N_49760);
nand UO_2705 (O_2705,N_49990,N_49768);
nand UO_2706 (O_2706,N_49932,N_49860);
or UO_2707 (O_2707,N_49845,N_49797);
xor UO_2708 (O_2708,N_49900,N_49826);
nand UO_2709 (O_2709,N_49871,N_49861);
nand UO_2710 (O_2710,N_49774,N_49921);
xnor UO_2711 (O_2711,N_49799,N_49808);
xor UO_2712 (O_2712,N_49846,N_49878);
xor UO_2713 (O_2713,N_49766,N_49920);
or UO_2714 (O_2714,N_49912,N_49962);
nand UO_2715 (O_2715,N_49997,N_49936);
xor UO_2716 (O_2716,N_49789,N_49923);
nor UO_2717 (O_2717,N_49808,N_49795);
or UO_2718 (O_2718,N_49787,N_49919);
and UO_2719 (O_2719,N_49966,N_49885);
xor UO_2720 (O_2720,N_49998,N_49952);
and UO_2721 (O_2721,N_49818,N_49929);
nor UO_2722 (O_2722,N_49769,N_49820);
nand UO_2723 (O_2723,N_49872,N_49965);
or UO_2724 (O_2724,N_49988,N_49907);
or UO_2725 (O_2725,N_49889,N_49786);
and UO_2726 (O_2726,N_49940,N_49977);
nand UO_2727 (O_2727,N_49960,N_49879);
or UO_2728 (O_2728,N_49800,N_49804);
or UO_2729 (O_2729,N_49973,N_49940);
and UO_2730 (O_2730,N_49842,N_49899);
and UO_2731 (O_2731,N_49870,N_49765);
nand UO_2732 (O_2732,N_49841,N_49811);
and UO_2733 (O_2733,N_49847,N_49949);
or UO_2734 (O_2734,N_49933,N_49798);
or UO_2735 (O_2735,N_49902,N_49788);
nand UO_2736 (O_2736,N_49878,N_49864);
and UO_2737 (O_2737,N_49760,N_49770);
or UO_2738 (O_2738,N_49900,N_49893);
nor UO_2739 (O_2739,N_49795,N_49763);
and UO_2740 (O_2740,N_49859,N_49902);
nand UO_2741 (O_2741,N_49927,N_49818);
xor UO_2742 (O_2742,N_49758,N_49850);
and UO_2743 (O_2743,N_49800,N_49917);
nor UO_2744 (O_2744,N_49885,N_49912);
or UO_2745 (O_2745,N_49897,N_49864);
xor UO_2746 (O_2746,N_49778,N_49801);
nor UO_2747 (O_2747,N_49829,N_49761);
nand UO_2748 (O_2748,N_49958,N_49856);
or UO_2749 (O_2749,N_49907,N_49950);
nor UO_2750 (O_2750,N_49783,N_49891);
or UO_2751 (O_2751,N_49755,N_49897);
or UO_2752 (O_2752,N_49793,N_49836);
xnor UO_2753 (O_2753,N_49834,N_49913);
nor UO_2754 (O_2754,N_49753,N_49913);
nor UO_2755 (O_2755,N_49924,N_49850);
or UO_2756 (O_2756,N_49820,N_49985);
xor UO_2757 (O_2757,N_49767,N_49966);
or UO_2758 (O_2758,N_49788,N_49904);
nor UO_2759 (O_2759,N_49861,N_49943);
and UO_2760 (O_2760,N_49895,N_49798);
and UO_2761 (O_2761,N_49895,N_49968);
nand UO_2762 (O_2762,N_49844,N_49860);
nor UO_2763 (O_2763,N_49892,N_49897);
nand UO_2764 (O_2764,N_49896,N_49862);
or UO_2765 (O_2765,N_49881,N_49767);
nor UO_2766 (O_2766,N_49821,N_49993);
and UO_2767 (O_2767,N_49846,N_49964);
xnor UO_2768 (O_2768,N_49804,N_49971);
nor UO_2769 (O_2769,N_49896,N_49916);
nand UO_2770 (O_2770,N_49803,N_49924);
or UO_2771 (O_2771,N_49804,N_49825);
nor UO_2772 (O_2772,N_49950,N_49953);
nor UO_2773 (O_2773,N_49956,N_49845);
or UO_2774 (O_2774,N_49782,N_49967);
nor UO_2775 (O_2775,N_49881,N_49809);
xnor UO_2776 (O_2776,N_49986,N_49827);
xnor UO_2777 (O_2777,N_49913,N_49851);
and UO_2778 (O_2778,N_49807,N_49753);
and UO_2779 (O_2779,N_49821,N_49942);
nor UO_2780 (O_2780,N_49884,N_49968);
xor UO_2781 (O_2781,N_49857,N_49967);
and UO_2782 (O_2782,N_49904,N_49944);
nor UO_2783 (O_2783,N_49817,N_49999);
nor UO_2784 (O_2784,N_49785,N_49843);
xor UO_2785 (O_2785,N_49990,N_49885);
xnor UO_2786 (O_2786,N_49933,N_49987);
nand UO_2787 (O_2787,N_49930,N_49823);
or UO_2788 (O_2788,N_49972,N_49911);
or UO_2789 (O_2789,N_49938,N_49820);
xnor UO_2790 (O_2790,N_49968,N_49877);
nor UO_2791 (O_2791,N_49834,N_49778);
and UO_2792 (O_2792,N_49917,N_49787);
xnor UO_2793 (O_2793,N_49946,N_49967);
nand UO_2794 (O_2794,N_49760,N_49796);
and UO_2795 (O_2795,N_49831,N_49907);
nor UO_2796 (O_2796,N_49834,N_49859);
nor UO_2797 (O_2797,N_49819,N_49790);
nand UO_2798 (O_2798,N_49914,N_49928);
or UO_2799 (O_2799,N_49983,N_49784);
nor UO_2800 (O_2800,N_49974,N_49846);
and UO_2801 (O_2801,N_49757,N_49893);
xor UO_2802 (O_2802,N_49930,N_49910);
or UO_2803 (O_2803,N_49793,N_49990);
xor UO_2804 (O_2804,N_49855,N_49809);
xor UO_2805 (O_2805,N_49966,N_49937);
xnor UO_2806 (O_2806,N_49890,N_49905);
and UO_2807 (O_2807,N_49968,N_49845);
xnor UO_2808 (O_2808,N_49918,N_49824);
and UO_2809 (O_2809,N_49804,N_49828);
and UO_2810 (O_2810,N_49803,N_49993);
xor UO_2811 (O_2811,N_49840,N_49863);
nor UO_2812 (O_2812,N_49766,N_49859);
or UO_2813 (O_2813,N_49767,N_49899);
nor UO_2814 (O_2814,N_49807,N_49761);
xnor UO_2815 (O_2815,N_49871,N_49836);
or UO_2816 (O_2816,N_49784,N_49773);
and UO_2817 (O_2817,N_49850,N_49910);
nand UO_2818 (O_2818,N_49887,N_49875);
nor UO_2819 (O_2819,N_49957,N_49812);
xor UO_2820 (O_2820,N_49770,N_49994);
or UO_2821 (O_2821,N_49886,N_49978);
nor UO_2822 (O_2822,N_49774,N_49775);
nand UO_2823 (O_2823,N_49903,N_49899);
nand UO_2824 (O_2824,N_49833,N_49831);
nor UO_2825 (O_2825,N_49990,N_49980);
nand UO_2826 (O_2826,N_49897,N_49762);
xnor UO_2827 (O_2827,N_49980,N_49856);
or UO_2828 (O_2828,N_49816,N_49999);
nand UO_2829 (O_2829,N_49881,N_49750);
xor UO_2830 (O_2830,N_49902,N_49849);
and UO_2831 (O_2831,N_49993,N_49998);
xnor UO_2832 (O_2832,N_49829,N_49880);
and UO_2833 (O_2833,N_49798,N_49810);
or UO_2834 (O_2834,N_49826,N_49825);
and UO_2835 (O_2835,N_49987,N_49830);
xor UO_2836 (O_2836,N_49786,N_49905);
and UO_2837 (O_2837,N_49837,N_49960);
and UO_2838 (O_2838,N_49839,N_49859);
nor UO_2839 (O_2839,N_49815,N_49756);
xor UO_2840 (O_2840,N_49816,N_49792);
nor UO_2841 (O_2841,N_49848,N_49809);
nor UO_2842 (O_2842,N_49953,N_49978);
xnor UO_2843 (O_2843,N_49752,N_49994);
and UO_2844 (O_2844,N_49912,N_49859);
nor UO_2845 (O_2845,N_49772,N_49814);
nor UO_2846 (O_2846,N_49883,N_49977);
xnor UO_2847 (O_2847,N_49895,N_49781);
or UO_2848 (O_2848,N_49861,N_49821);
nand UO_2849 (O_2849,N_49856,N_49759);
and UO_2850 (O_2850,N_49997,N_49961);
and UO_2851 (O_2851,N_49972,N_49771);
and UO_2852 (O_2852,N_49855,N_49793);
xnor UO_2853 (O_2853,N_49965,N_49762);
and UO_2854 (O_2854,N_49973,N_49811);
or UO_2855 (O_2855,N_49837,N_49779);
and UO_2856 (O_2856,N_49945,N_49817);
or UO_2857 (O_2857,N_49854,N_49868);
nand UO_2858 (O_2858,N_49870,N_49964);
nand UO_2859 (O_2859,N_49845,N_49799);
nand UO_2860 (O_2860,N_49902,N_49919);
xnor UO_2861 (O_2861,N_49815,N_49948);
or UO_2862 (O_2862,N_49904,N_49970);
or UO_2863 (O_2863,N_49969,N_49992);
xnor UO_2864 (O_2864,N_49803,N_49800);
nor UO_2865 (O_2865,N_49756,N_49890);
nor UO_2866 (O_2866,N_49818,N_49865);
nor UO_2867 (O_2867,N_49945,N_49996);
or UO_2868 (O_2868,N_49799,N_49889);
or UO_2869 (O_2869,N_49756,N_49988);
or UO_2870 (O_2870,N_49768,N_49936);
nor UO_2871 (O_2871,N_49759,N_49855);
nor UO_2872 (O_2872,N_49896,N_49752);
or UO_2873 (O_2873,N_49950,N_49845);
and UO_2874 (O_2874,N_49849,N_49886);
or UO_2875 (O_2875,N_49902,N_49760);
nand UO_2876 (O_2876,N_49993,N_49806);
xor UO_2877 (O_2877,N_49842,N_49767);
nor UO_2878 (O_2878,N_49789,N_49879);
xor UO_2879 (O_2879,N_49984,N_49810);
or UO_2880 (O_2880,N_49974,N_49774);
xnor UO_2881 (O_2881,N_49971,N_49870);
or UO_2882 (O_2882,N_49929,N_49963);
nand UO_2883 (O_2883,N_49992,N_49917);
xnor UO_2884 (O_2884,N_49972,N_49766);
xnor UO_2885 (O_2885,N_49844,N_49982);
xor UO_2886 (O_2886,N_49788,N_49986);
or UO_2887 (O_2887,N_49978,N_49894);
nor UO_2888 (O_2888,N_49866,N_49876);
nand UO_2889 (O_2889,N_49931,N_49966);
and UO_2890 (O_2890,N_49800,N_49820);
or UO_2891 (O_2891,N_49974,N_49803);
xor UO_2892 (O_2892,N_49914,N_49847);
nor UO_2893 (O_2893,N_49989,N_49918);
nand UO_2894 (O_2894,N_49882,N_49886);
xnor UO_2895 (O_2895,N_49933,N_49894);
nor UO_2896 (O_2896,N_49955,N_49871);
xnor UO_2897 (O_2897,N_49928,N_49877);
and UO_2898 (O_2898,N_49806,N_49866);
nand UO_2899 (O_2899,N_49813,N_49971);
nand UO_2900 (O_2900,N_49921,N_49870);
nor UO_2901 (O_2901,N_49940,N_49900);
or UO_2902 (O_2902,N_49823,N_49841);
xnor UO_2903 (O_2903,N_49996,N_49875);
and UO_2904 (O_2904,N_49832,N_49913);
nor UO_2905 (O_2905,N_49873,N_49806);
nand UO_2906 (O_2906,N_49940,N_49945);
nand UO_2907 (O_2907,N_49941,N_49947);
and UO_2908 (O_2908,N_49846,N_49941);
nor UO_2909 (O_2909,N_49978,N_49903);
nor UO_2910 (O_2910,N_49801,N_49946);
nand UO_2911 (O_2911,N_49989,N_49859);
or UO_2912 (O_2912,N_49772,N_49799);
xnor UO_2913 (O_2913,N_49840,N_49757);
nand UO_2914 (O_2914,N_49755,N_49806);
and UO_2915 (O_2915,N_49846,N_49927);
or UO_2916 (O_2916,N_49758,N_49849);
and UO_2917 (O_2917,N_49926,N_49776);
nand UO_2918 (O_2918,N_49861,N_49973);
nand UO_2919 (O_2919,N_49853,N_49812);
or UO_2920 (O_2920,N_49870,N_49838);
nor UO_2921 (O_2921,N_49801,N_49888);
xnor UO_2922 (O_2922,N_49999,N_49982);
or UO_2923 (O_2923,N_49889,N_49973);
xnor UO_2924 (O_2924,N_49797,N_49948);
nand UO_2925 (O_2925,N_49945,N_49790);
nor UO_2926 (O_2926,N_49981,N_49836);
nand UO_2927 (O_2927,N_49912,N_49898);
nor UO_2928 (O_2928,N_49933,N_49938);
nand UO_2929 (O_2929,N_49838,N_49882);
nand UO_2930 (O_2930,N_49976,N_49844);
nor UO_2931 (O_2931,N_49994,N_49887);
or UO_2932 (O_2932,N_49825,N_49879);
and UO_2933 (O_2933,N_49780,N_49944);
and UO_2934 (O_2934,N_49995,N_49988);
or UO_2935 (O_2935,N_49854,N_49913);
nand UO_2936 (O_2936,N_49872,N_49880);
xnor UO_2937 (O_2937,N_49941,N_49781);
nor UO_2938 (O_2938,N_49936,N_49830);
nor UO_2939 (O_2939,N_49911,N_49777);
or UO_2940 (O_2940,N_49853,N_49763);
nor UO_2941 (O_2941,N_49818,N_49786);
or UO_2942 (O_2942,N_49873,N_49907);
nor UO_2943 (O_2943,N_49815,N_49769);
or UO_2944 (O_2944,N_49821,N_49956);
nor UO_2945 (O_2945,N_49855,N_49997);
nor UO_2946 (O_2946,N_49922,N_49811);
and UO_2947 (O_2947,N_49993,N_49780);
and UO_2948 (O_2948,N_49885,N_49972);
xnor UO_2949 (O_2949,N_49788,N_49818);
nand UO_2950 (O_2950,N_49823,N_49939);
and UO_2951 (O_2951,N_49850,N_49764);
nand UO_2952 (O_2952,N_49766,N_49868);
and UO_2953 (O_2953,N_49935,N_49885);
xnor UO_2954 (O_2954,N_49899,N_49982);
and UO_2955 (O_2955,N_49906,N_49907);
or UO_2956 (O_2956,N_49907,N_49775);
xor UO_2957 (O_2957,N_49932,N_49877);
and UO_2958 (O_2958,N_49925,N_49803);
xor UO_2959 (O_2959,N_49917,N_49957);
nand UO_2960 (O_2960,N_49961,N_49758);
xor UO_2961 (O_2961,N_49805,N_49826);
or UO_2962 (O_2962,N_49867,N_49873);
xnor UO_2963 (O_2963,N_49961,N_49989);
nor UO_2964 (O_2964,N_49862,N_49977);
xnor UO_2965 (O_2965,N_49979,N_49866);
nand UO_2966 (O_2966,N_49790,N_49904);
or UO_2967 (O_2967,N_49977,N_49866);
xor UO_2968 (O_2968,N_49923,N_49847);
nor UO_2969 (O_2969,N_49953,N_49943);
nand UO_2970 (O_2970,N_49962,N_49928);
xor UO_2971 (O_2971,N_49862,N_49785);
and UO_2972 (O_2972,N_49949,N_49827);
nor UO_2973 (O_2973,N_49806,N_49758);
nand UO_2974 (O_2974,N_49806,N_49845);
and UO_2975 (O_2975,N_49851,N_49973);
or UO_2976 (O_2976,N_49997,N_49994);
or UO_2977 (O_2977,N_49813,N_49826);
nand UO_2978 (O_2978,N_49910,N_49781);
nand UO_2979 (O_2979,N_49924,N_49817);
or UO_2980 (O_2980,N_49788,N_49878);
nor UO_2981 (O_2981,N_49868,N_49780);
nor UO_2982 (O_2982,N_49935,N_49800);
xor UO_2983 (O_2983,N_49865,N_49885);
nand UO_2984 (O_2984,N_49951,N_49904);
and UO_2985 (O_2985,N_49953,N_49968);
and UO_2986 (O_2986,N_49905,N_49793);
and UO_2987 (O_2987,N_49904,N_49882);
and UO_2988 (O_2988,N_49847,N_49877);
or UO_2989 (O_2989,N_49878,N_49919);
nand UO_2990 (O_2990,N_49827,N_49753);
and UO_2991 (O_2991,N_49863,N_49947);
nand UO_2992 (O_2992,N_49957,N_49792);
nor UO_2993 (O_2993,N_49829,N_49863);
and UO_2994 (O_2994,N_49753,N_49786);
or UO_2995 (O_2995,N_49879,N_49937);
or UO_2996 (O_2996,N_49951,N_49846);
or UO_2997 (O_2997,N_49989,N_49878);
xor UO_2998 (O_2998,N_49940,N_49929);
and UO_2999 (O_2999,N_49825,N_49897);
and UO_3000 (O_3000,N_49980,N_49943);
and UO_3001 (O_3001,N_49790,N_49869);
nand UO_3002 (O_3002,N_49905,N_49935);
or UO_3003 (O_3003,N_49992,N_49822);
nor UO_3004 (O_3004,N_49790,N_49830);
xor UO_3005 (O_3005,N_49799,N_49927);
nor UO_3006 (O_3006,N_49828,N_49998);
and UO_3007 (O_3007,N_49937,N_49755);
or UO_3008 (O_3008,N_49835,N_49995);
or UO_3009 (O_3009,N_49896,N_49762);
or UO_3010 (O_3010,N_49759,N_49806);
nand UO_3011 (O_3011,N_49898,N_49939);
xnor UO_3012 (O_3012,N_49810,N_49801);
xnor UO_3013 (O_3013,N_49949,N_49751);
or UO_3014 (O_3014,N_49824,N_49995);
xnor UO_3015 (O_3015,N_49970,N_49998);
nor UO_3016 (O_3016,N_49943,N_49907);
nand UO_3017 (O_3017,N_49785,N_49985);
nor UO_3018 (O_3018,N_49940,N_49850);
xor UO_3019 (O_3019,N_49794,N_49827);
xnor UO_3020 (O_3020,N_49907,N_49773);
xor UO_3021 (O_3021,N_49863,N_49802);
nand UO_3022 (O_3022,N_49786,N_49954);
nor UO_3023 (O_3023,N_49834,N_49900);
nor UO_3024 (O_3024,N_49796,N_49893);
and UO_3025 (O_3025,N_49963,N_49796);
nor UO_3026 (O_3026,N_49890,N_49857);
xor UO_3027 (O_3027,N_49974,N_49976);
nor UO_3028 (O_3028,N_49898,N_49781);
and UO_3029 (O_3029,N_49819,N_49922);
and UO_3030 (O_3030,N_49945,N_49850);
and UO_3031 (O_3031,N_49949,N_49837);
xnor UO_3032 (O_3032,N_49960,N_49827);
nand UO_3033 (O_3033,N_49837,N_49892);
or UO_3034 (O_3034,N_49807,N_49969);
nand UO_3035 (O_3035,N_49895,N_49811);
xor UO_3036 (O_3036,N_49994,N_49824);
and UO_3037 (O_3037,N_49947,N_49971);
xnor UO_3038 (O_3038,N_49840,N_49830);
nand UO_3039 (O_3039,N_49936,N_49809);
nor UO_3040 (O_3040,N_49811,N_49925);
xor UO_3041 (O_3041,N_49875,N_49779);
or UO_3042 (O_3042,N_49761,N_49818);
nand UO_3043 (O_3043,N_49838,N_49951);
nor UO_3044 (O_3044,N_49852,N_49799);
and UO_3045 (O_3045,N_49794,N_49839);
xnor UO_3046 (O_3046,N_49858,N_49992);
nand UO_3047 (O_3047,N_49773,N_49971);
xnor UO_3048 (O_3048,N_49788,N_49772);
or UO_3049 (O_3049,N_49825,N_49984);
xnor UO_3050 (O_3050,N_49782,N_49821);
nor UO_3051 (O_3051,N_49926,N_49982);
xor UO_3052 (O_3052,N_49789,N_49773);
or UO_3053 (O_3053,N_49768,N_49823);
and UO_3054 (O_3054,N_49936,N_49811);
or UO_3055 (O_3055,N_49976,N_49842);
xnor UO_3056 (O_3056,N_49876,N_49816);
and UO_3057 (O_3057,N_49825,N_49889);
nand UO_3058 (O_3058,N_49964,N_49902);
nand UO_3059 (O_3059,N_49922,N_49753);
or UO_3060 (O_3060,N_49822,N_49893);
or UO_3061 (O_3061,N_49752,N_49931);
and UO_3062 (O_3062,N_49988,N_49878);
xnor UO_3063 (O_3063,N_49975,N_49970);
or UO_3064 (O_3064,N_49834,N_49950);
and UO_3065 (O_3065,N_49815,N_49929);
nor UO_3066 (O_3066,N_49803,N_49876);
nor UO_3067 (O_3067,N_49758,N_49976);
and UO_3068 (O_3068,N_49819,N_49764);
nand UO_3069 (O_3069,N_49827,N_49983);
and UO_3070 (O_3070,N_49775,N_49956);
nor UO_3071 (O_3071,N_49885,N_49844);
xnor UO_3072 (O_3072,N_49979,N_49892);
xnor UO_3073 (O_3073,N_49809,N_49875);
and UO_3074 (O_3074,N_49777,N_49824);
and UO_3075 (O_3075,N_49842,N_49813);
or UO_3076 (O_3076,N_49897,N_49766);
nor UO_3077 (O_3077,N_49800,N_49841);
and UO_3078 (O_3078,N_49889,N_49935);
and UO_3079 (O_3079,N_49939,N_49773);
and UO_3080 (O_3080,N_49840,N_49934);
xor UO_3081 (O_3081,N_49880,N_49917);
xor UO_3082 (O_3082,N_49851,N_49868);
nand UO_3083 (O_3083,N_49765,N_49757);
nor UO_3084 (O_3084,N_49982,N_49901);
xor UO_3085 (O_3085,N_49847,N_49839);
xor UO_3086 (O_3086,N_49802,N_49815);
nor UO_3087 (O_3087,N_49863,N_49925);
and UO_3088 (O_3088,N_49992,N_49885);
nor UO_3089 (O_3089,N_49804,N_49814);
nor UO_3090 (O_3090,N_49891,N_49885);
or UO_3091 (O_3091,N_49776,N_49821);
nand UO_3092 (O_3092,N_49815,N_49855);
nand UO_3093 (O_3093,N_49818,N_49998);
nor UO_3094 (O_3094,N_49910,N_49911);
nand UO_3095 (O_3095,N_49877,N_49817);
xnor UO_3096 (O_3096,N_49829,N_49858);
and UO_3097 (O_3097,N_49795,N_49848);
or UO_3098 (O_3098,N_49781,N_49933);
xnor UO_3099 (O_3099,N_49962,N_49985);
and UO_3100 (O_3100,N_49895,N_49981);
nor UO_3101 (O_3101,N_49999,N_49811);
and UO_3102 (O_3102,N_49991,N_49756);
nand UO_3103 (O_3103,N_49764,N_49975);
nand UO_3104 (O_3104,N_49806,N_49945);
and UO_3105 (O_3105,N_49861,N_49996);
and UO_3106 (O_3106,N_49845,N_49844);
or UO_3107 (O_3107,N_49909,N_49891);
nand UO_3108 (O_3108,N_49896,N_49935);
and UO_3109 (O_3109,N_49908,N_49816);
or UO_3110 (O_3110,N_49762,N_49919);
and UO_3111 (O_3111,N_49949,N_49863);
or UO_3112 (O_3112,N_49887,N_49903);
and UO_3113 (O_3113,N_49786,N_49894);
and UO_3114 (O_3114,N_49798,N_49755);
and UO_3115 (O_3115,N_49999,N_49896);
and UO_3116 (O_3116,N_49906,N_49928);
and UO_3117 (O_3117,N_49787,N_49835);
nor UO_3118 (O_3118,N_49852,N_49914);
xnor UO_3119 (O_3119,N_49773,N_49982);
nand UO_3120 (O_3120,N_49968,N_49754);
or UO_3121 (O_3121,N_49834,N_49807);
xor UO_3122 (O_3122,N_49765,N_49770);
or UO_3123 (O_3123,N_49947,N_49850);
and UO_3124 (O_3124,N_49801,N_49875);
nand UO_3125 (O_3125,N_49854,N_49787);
and UO_3126 (O_3126,N_49851,N_49834);
or UO_3127 (O_3127,N_49944,N_49906);
nor UO_3128 (O_3128,N_49801,N_49878);
or UO_3129 (O_3129,N_49885,N_49857);
and UO_3130 (O_3130,N_49935,N_49959);
and UO_3131 (O_3131,N_49880,N_49823);
or UO_3132 (O_3132,N_49768,N_49868);
nand UO_3133 (O_3133,N_49908,N_49861);
xnor UO_3134 (O_3134,N_49999,N_49917);
nand UO_3135 (O_3135,N_49790,N_49845);
or UO_3136 (O_3136,N_49757,N_49807);
nor UO_3137 (O_3137,N_49943,N_49878);
or UO_3138 (O_3138,N_49863,N_49875);
xnor UO_3139 (O_3139,N_49830,N_49839);
xnor UO_3140 (O_3140,N_49966,N_49833);
and UO_3141 (O_3141,N_49864,N_49829);
xnor UO_3142 (O_3142,N_49786,N_49886);
xnor UO_3143 (O_3143,N_49923,N_49754);
nor UO_3144 (O_3144,N_49957,N_49803);
xnor UO_3145 (O_3145,N_49826,N_49781);
or UO_3146 (O_3146,N_49771,N_49789);
or UO_3147 (O_3147,N_49936,N_49891);
or UO_3148 (O_3148,N_49930,N_49758);
nor UO_3149 (O_3149,N_49879,N_49761);
and UO_3150 (O_3150,N_49896,N_49822);
xnor UO_3151 (O_3151,N_49893,N_49760);
and UO_3152 (O_3152,N_49823,N_49914);
xnor UO_3153 (O_3153,N_49776,N_49928);
and UO_3154 (O_3154,N_49751,N_49962);
and UO_3155 (O_3155,N_49850,N_49813);
or UO_3156 (O_3156,N_49880,N_49884);
nor UO_3157 (O_3157,N_49887,N_49797);
nand UO_3158 (O_3158,N_49899,N_49977);
nor UO_3159 (O_3159,N_49916,N_49877);
xnor UO_3160 (O_3160,N_49868,N_49903);
xor UO_3161 (O_3161,N_49939,N_49998);
xor UO_3162 (O_3162,N_49989,N_49827);
or UO_3163 (O_3163,N_49981,N_49820);
nor UO_3164 (O_3164,N_49964,N_49871);
xnor UO_3165 (O_3165,N_49988,N_49786);
nor UO_3166 (O_3166,N_49978,N_49981);
nor UO_3167 (O_3167,N_49851,N_49963);
and UO_3168 (O_3168,N_49941,N_49787);
or UO_3169 (O_3169,N_49935,N_49908);
or UO_3170 (O_3170,N_49825,N_49927);
or UO_3171 (O_3171,N_49752,N_49819);
nor UO_3172 (O_3172,N_49870,N_49896);
nor UO_3173 (O_3173,N_49818,N_49915);
xnor UO_3174 (O_3174,N_49966,N_49921);
and UO_3175 (O_3175,N_49886,N_49776);
nor UO_3176 (O_3176,N_49761,N_49805);
xnor UO_3177 (O_3177,N_49988,N_49828);
xor UO_3178 (O_3178,N_49839,N_49985);
nor UO_3179 (O_3179,N_49765,N_49967);
or UO_3180 (O_3180,N_49981,N_49791);
nor UO_3181 (O_3181,N_49844,N_49773);
nand UO_3182 (O_3182,N_49935,N_49893);
and UO_3183 (O_3183,N_49954,N_49784);
or UO_3184 (O_3184,N_49822,N_49791);
nand UO_3185 (O_3185,N_49913,N_49900);
or UO_3186 (O_3186,N_49962,N_49808);
xnor UO_3187 (O_3187,N_49971,N_49999);
nand UO_3188 (O_3188,N_49776,N_49863);
xor UO_3189 (O_3189,N_49769,N_49973);
or UO_3190 (O_3190,N_49840,N_49759);
and UO_3191 (O_3191,N_49992,N_49911);
and UO_3192 (O_3192,N_49904,N_49813);
and UO_3193 (O_3193,N_49889,N_49966);
or UO_3194 (O_3194,N_49905,N_49947);
nor UO_3195 (O_3195,N_49978,N_49785);
nand UO_3196 (O_3196,N_49894,N_49781);
nand UO_3197 (O_3197,N_49989,N_49766);
or UO_3198 (O_3198,N_49792,N_49929);
and UO_3199 (O_3199,N_49977,N_49805);
and UO_3200 (O_3200,N_49820,N_49786);
nor UO_3201 (O_3201,N_49798,N_49881);
or UO_3202 (O_3202,N_49792,N_49907);
and UO_3203 (O_3203,N_49840,N_49973);
or UO_3204 (O_3204,N_49880,N_49790);
xnor UO_3205 (O_3205,N_49915,N_49822);
nor UO_3206 (O_3206,N_49931,N_49987);
and UO_3207 (O_3207,N_49765,N_49965);
xnor UO_3208 (O_3208,N_49769,N_49896);
nand UO_3209 (O_3209,N_49845,N_49795);
nand UO_3210 (O_3210,N_49868,N_49954);
or UO_3211 (O_3211,N_49817,N_49770);
and UO_3212 (O_3212,N_49785,N_49967);
nor UO_3213 (O_3213,N_49833,N_49777);
and UO_3214 (O_3214,N_49774,N_49942);
nand UO_3215 (O_3215,N_49808,N_49914);
nor UO_3216 (O_3216,N_49991,N_49798);
xor UO_3217 (O_3217,N_49761,N_49753);
and UO_3218 (O_3218,N_49766,N_49772);
xnor UO_3219 (O_3219,N_49814,N_49791);
nand UO_3220 (O_3220,N_49789,N_49961);
nor UO_3221 (O_3221,N_49916,N_49899);
xnor UO_3222 (O_3222,N_49955,N_49789);
xnor UO_3223 (O_3223,N_49924,N_49823);
nor UO_3224 (O_3224,N_49811,N_49824);
nand UO_3225 (O_3225,N_49754,N_49966);
or UO_3226 (O_3226,N_49911,N_49810);
or UO_3227 (O_3227,N_49761,N_49928);
nor UO_3228 (O_3228,N_49930,N_49993);
or UO_3229 (O_3229,N_49802,N_49887);
or UO_3230 (O_3230,N_49966,N_49822);
nand UO_3231 (O_3231,N_49991,N_49840);
xor UO_3232 (O_3232,N_49922,N_49889);
xor UO_3233 (O_3233,N_49877,N_49980);
or UO_3234 (O_3234,N_49860,N_49989);
nor UO_3235 (O_3235,N_49923,N_49790);
xor UO_3236 (O_3236,N_49916,N_49803);
or UO_3237 (O_3237,N_49921,N_49787);
and UO_3238 (O_3238,N_49808,N_49977);
and UO_3239 (O_3239,N_49942,N_49895);
xnor UO_3240 (O_3240,N_49825,N_49951);
xnor UO_3241 (O_3241,N_49751,N_49982);
and UO_3242 (O_3242,N_49955,N_49779);
or UO_3243 (O_3243,N_49840,N_49819);
nor UO_3244 (O_3244,N_49807,N_49840);
and UO_3245 (O_3245,N_49763,N_49802);
nor UO_3246 (O_3246,N_49975,N_49803);
nor UO_3247 (O_3247,N_49841,N_49883);
nand UO_3248 (O_3248,N_49928,N_49955);
and UO_3249 (O_3249,N_49980,N_49780);
and UO_3250 (O_3250,N_49840,N_49839);
xor UO_3251 (O_3251,N_49892,N_49931);
nand UO_3252 (O_3252,N_49809,N_49802);
nor UO_3253 (O_3253,N_49814,N_49893);
or UO_3254 (O_3254,N_49754,N_49784);
and UO_3255 (O_3255,N_49847,N_49905);
or UO_3256 (O_3256,N_49998,N_49855);
and UO_3257 (O_3257,N_49955,N_49831);
xnor UO_3258 (O_3258,N_49873,N_49841);
or UO_3259 (O_3259,N_49952,N_49996);
or UO_3260 (O_3260,N_49960,N_49832);
nand UO_3261 (O_3261,N_49962,N_49829);
or UO_3262 (O_3262,N_49774,N_49752);
nor UO_3263 (O_3263,N_49892,N_49994);
xnor UO_3264 (O_3264,N_49808,N_49964);
or UO_3265 (O_3265,N_49944,N_49979);
xnor UO_3266 (O_3266,N_49977,N_49970);
nand UO_3267 (O_3267,N_49783,N_49815);
xor UO_3268 (O_3268,N_49887,N_49940);
xor UO_3269 (O_3269,N_49926,N_49990);
xor UO_3270 (O_3270,N_49892,N_49908);
xor UO_3271 (O_3271,N_49916,N_49860);
nand UO_3272 (O_3272,N_49963,N_49772);
and UO_3273 (O_3273,N_49901,N_49933);
xor UO_3274 (O_3274,N_49865,N_49984);
xor UO_3275 (O_3275,N_49852,N_49888);
nor UO_3276 (O_3276,N_49930,N_49906);
nor UO_3277 (O_3277,N_49833,N_49837);
and UO_3278 (O_3278,N_49985,N_49969);
and UO_3279 (O_3279,N_49777,N_49967);
xnor UO_3280 (O_3280,N_49948,N_49843);
or UO_3281 (O_3281,N_49968,N_49780);
nand UO_3282 (O_3282,N_49770,N_49814);
nor UO_3283 (O_3283,N_49914,N_49972);
nor UO_3284 (O_3284,N_49814,N_49798);
nor UO_3285 (O_3285,N_49964,N_49953);
and UO_3286 (O_3286,N_49828,N_49986);
nand UO_3287 (O_3287,N_49947,N_49763);
xor UO_3288 (O_3288,N_49929,N_49904);
and UO_3289 (O_3289,N_49781,N_49970);
or UO_3290 (O_3290,N_49916,N_49856);
or UO_3291 (O_3291,N_49785,N_49859);
nand UO_3292 (O_3292,N_49784,N_49950);
nand UO_3293 (O_3293,N_49785,N_49989);
or UO_3294 (O_3294,N_49976,N_49819);
and UO_3295 (O_3295,N_49957,N_49999);
nor UO_3296 (O_3296,N_49920,N_49894);
or UO_3297 (O_3297,N_49962,N_49851);
or UO_3298 (O_3298,N_49858,N_49761);
and UO_3299 (O_3299,N_49775,N_49946);
and UO_3300 (O_3300,N_49971,N_49838);
xor UO_3301 (O_3301,N_49833,N_49921);
xor UO_3302 (O_3302,N_49940,N_49928);
and UO_3303 (O_3303,N_49790,N_49878);
nor UO_3304 (O_3304,N_49811,N_49805);
or UO_3305 (O_3305,N_49813,N_49789);
xnor UO_3306 (O_3306,N_49923,N_49919);
xor UO_3307 (O_3307,N_49788,N_49787);
or UO_3308 (O_3308,N_49981,N_49887);
nand UO_3309 (O_3309,N_49871,N_49998);
xnor UO_3310 (O_3310,N_49940,N_49826);
and UO_3311 (O_3311,N_49846,N_49844);
nor UO_3312 (O_3312,N_49966,N_49997);
and UO_3313 (O_3313,N_49919,N_49943);
nor UO_3314 (O_3314,N_49973,N_49791);
xor UO_3315 (O_3315,N_49865,N_49834);
nor UO_3316 (O_3316,N_49901,N_49809);
nand UO_3317 (O_3317,N_49952,N_49773);
nor UO_3318 (O_3318,N_49923,N_49852);
and UO_3319 (O_3319,N_49896,N_49806);
and UO_3320 (O_3320,N_49927,N_49772);
or UO_3321 (O_3321,N_49862,N_49798);
nor UO_3322 (O_3322,N_49976,N_49849);
nand UO_3323 (O_3323,N_49922,N_49945);
nand UO_3324 (O_3324,N_49880,N_49991);
or UO_3325 (O_3325,N_49956,N_49857);
or UO_3326 (O_3326,N_49917,N_49920);
and UO_3327 (O_3327,N_49971,N_49843);
nand UO_3328 (O_3328,N_49827,N_49762);
nor UO_3329 (O_3329,N_49884,N_49808);
or UO_3330 (O_3330,N_49802,N_49993);
nor UO_3331 (O_3331,N_49925,N_49832);
xor UO_3332 (O_3332,N_49835,N_49789);
nand UO_3333 (O_3333,N_49829,N_49968);
or UO_3334 (O_3334,N_49904,N_49794);
nand UO_3335 (O_3335,N_49814,N_49996);
nor UO_3336 (O_3336,N_49774,N_49853);
or UO_3337 (O_3337,N_49852,N_49830);
or UO_3338 (O_3338,N_49763,N_49854);
xor UO_3339 (O_3339,N_49960,N_49797);
or UO_3340 (O_3340,N_49837,N_49841);
or UO_3341 (O_3341,N_49757,N_49850);
or UO_3342 (O_3342,N_49867,N_49971);
nor UO_3343 (O_3343,N_49900,N_49761);
xor UO_3344 (O_3344,N_49936,N_49870);
xor UO_3345 (O_3345,N_49818,N_49906);
and UO_3346 (O_3346,N_49752,N_49849);
nand UO_3347 (O_3347,N_49858,N_49806);
nor UO_3348 (O_3348,N_49888,N_49981);
nor UO_3349 (O_3349,N_49863,N_49788);
and UO_3350 (O_3350,N_49863,N_49809);
or UO_3351 (O_3351,N_49968,N_49861);
or UO_3352 (O_3352,N_49758,N_49775);
xor UO_3353 (O_3353,N_49888,N_49829);
xnor UO_3354 (O_3354,N_49765,N_49920);
nor UO_3355 (O_3355,N_49844,N_49893);
nand UO_3356 (O_3356,N_49797,N_49944);
or UO_3357 (O_3357,N_49771,N_49882);
nand UO_3358 (O_3358,N_49776,N_49847);
and UO_3359 (O_3359,N_49838,N_49789);
and UO_3360 (O_3360,N_49851,N_49824);
nor UO_3361 (O_3361,N_49884,N_49866);
nand UO_3362 (O_3362,N_49895,N_49961);
or UO_3363 (O_3363,N_49782,N_49964);
and UO_3364 (O_3364,N_49974,N_49961);
xor UO_3365 (O_3365,N_49911,N_49789);
xor UO_3366 (O_3366,N_49840,N_49968);
or UO_3367 (O_3367,N_49768,N_49900);
nor UO_3368 (O_3368,N_49969,N_49820);
or UO_3369 (O_3369,N_49751,N_49947);
or UO_3370 (O_3370,N_49816,N_49754);
nor UO_3371 (O_3371,N_49828,N_49967);
or UO_3372 (O_3372,N_49764,N_49865);
xor UO_3373 (O_3373,N_49955,N_49988);
nand UO_3374 (O_3374,N_49925,N_49986);
nand UO_3375 (O_3375,N_49981,N_49972);
xor UO_3376 (O_3376,N_49832,N_49843);
nor UO_3377 (O_3377,N_49915,N_49914);
nor UO_3378 (O_3378,N_49833,N_49860);
nand UO_3379 (O_3379,N_49860,N_49784);
or UO_3380 (O_3380,N_49791,N_49769);
nor UO_3381 (O_3381,N_49754,N_49826);
nand UO_3382 (O_3382,N_49864,N_49837);
nand UO_3383 (O_3383,N_49770,N_49830);
or UO_3384 (O_3384,N_49760,N_49764);
or UO_3385 (O_3385,N_49920,N_49853);
nor UO_3386 (O_3386,N_49859,N_49853);
nor UO_3387 (O_3387,N_49993,N_49842);
nand UO_3388 (O_3388,N_49963,N_49756);
nor UO_3389 (O_3389,N_49976,N_49933);
nand UO_3390 (O_3390,N_49755,N_49996);
nor UO_3391 (O_3391,N_49869,N_49854);
and UO_3392 (O_3392,N_49909,N_49889);
nor UO_3393 (O_3393,N_49921,N_49786);
nand UO_3394 (O_3394,N_49937,N_49930);
xor UO_3395 (O_3395,N_49914,N_49807);
nor UO_3396 (O_3396,N_49925,N_49995);
nor UO_3397 (O_3397,N_49892,N_49906);
or UO_3398 (O_3398,N_49806,N_49839);
xor UO_3399 (O_3399,N_49926,N_49801);
nand UO_3400 (O_3400,N_49999,N_49970);
nor UO_3401 (O_3401,N_49822,N_49965);
or UO_3402 (O_3402,N_49916,N_49881);
xor UO_3403 (O_3403,N_49792,N_49880);
nand UO_3404 (O_3404,N_49758,N_49832);
nand UO_3405 (O_3405,N_49970,N_49966);
nor UO_3406 (O_3406,N_49752,N_49848);
or UO_3407 (O_3407,N_49785,N_49751);
nand UO_3408 (O_3408,N_49873,N_49852);
nor UO_3409 (O_3409,N_49896,N_49798);
or UO_3410 (O_3410,N_49979,N_49872);
nor UO_3411 (O_3411,N_49760,N_49816);
xor UO_3412 (O_3412,N_49952,N_49963);
nand UO_3413 (O_3413,N_49932,N_49826);
nor UO_3414 (O_3414,N_49939,N_49974);
and UO_3415 (O_3415,N_49820,N_49778);
or UO_3416 (O_3416,N_49885,N_49940);
and UO_3417 (O_3417,N_49950,N_49926);
xnor UO_3418 (O_3418,N_49973,N_49806);
nand UO_3419 (O_3419,N_49855,N_49750);
and UO_3420 (O_3420,N_49967,N_49816);
and UO_3421 (O_3421,N_49790,N_49993);
or UO_3422 (O_3422,N_49790,N_49984);
nand UO_3423 (O_3423,N_49756,N_49881);
xor UO_3424 (O_3424,N_49982,N_49838);
nand UO_3425 (O_3425,N_49913,N_49997);
xor UO_3426 (O_3426,N_49950,N_49896);
and UO_3427 (O_3427,N_49821,N_49814);
nor UO_3428 (O_3428,N_49881,N_49862);
or UO_3429 (O_3429,N_49893,N_49800);
xnor UO_3430 (O_3430,N_49961,N_49871);
nor UO_3431 (O_3431,N_49826,N_49830);
nor UO_3432 (O_3432,N_49910,N_49892);
and UO_3433 (O_3433,N_49916,N_49766);
nand UO_3434 (O_3434,N_49841,N_49832);
nand UO_3435 (O_3435,N_49954,N_49886);
xor UO_3436 (O_3436,N_49997,N_49826);
and UO_3437 (O_3437,N_49917,N_49770);
or UO_3438 (O_3438,N_49791,N_49867);
xnor UO_3439 (O_3439,N_49939,N_49781);
nand UO_3440 (O_3440,N_49949,N_49771);
or UO_3441 (O_3441,N_49754,N_49798);
or UO_3442 (O_3442,N_49815,N_49945);
or UO_3443 (O_3443,N_49934,N_49844);
nor UO_3444 (O_3444,N_49964,N_49827);
or UO_3445 (O_3445,N_49852,N_49987);
xor UO_3446 (O_3446,N_49784,N_49779);
nor UO_3447 (O_3447,N_49926,N_49882);
and UO_3448 (O_3448,N_49762,N_49978);
nand UO_3449 (O_3449,N_49783,N_49943);
or UO_3450 (O_3450,N_49921,N_49961);
nor UO_3451 (O_3451,N_49840,N_49954);
or UO_3452 (O_3452,N_49945,N_49877);
nor UO_3453 (O_3453,N_49846,N_49754);
xnor UO_3454 (O_3454,N_49870,N_49990);
nand UO_3455 (O_3455,N_49988,N_49916);
xor UO_3456 (O_3456,N_49948,N_49761);
nor UO_3457 (O_3457,N_49828,N_49785);
or UO_3458 (O_3458,N_49935,N_49902);
nor UO_3459 (O_3459,N_49848,N_49818);
nor UO_3460 (O_3460,N_49956,N_49906);
nand UO_3461 (O_3461,N_49837,N_49899);
or UO_3462 (O_3462,N_49892,N_49924);
xnor UO_3463 (O_3463,N_49890,N_49782);
and UO_3464 (O_3464,N_49988,N_49851);
nand UO_3465 (O_3465,N_49901,N_49848);
nor UO_3466 (O_3466,N_49975,N_49962);
nand UO_3467 (O_3467,N_49903,N_49840);
or UO_3468 (O_3468,N_49861,N_49984);
or UO_3469 (O_3469,N_49757,N_49978);
or UO_3470 (O_3470,N_49914,N_49969);
or UO_3471 (O_3471,N_49945,N_49934);
xnor UO_3472 (O_3472,N_49846,N_49901);
nand UO_3473 (O_3473,N_49906,N_49984);
nand UO_3474 (O_3474,N_49789,N_49893);
or UO_3475 (O_3475,N_49913,N_49805);
nand UO_3476 (O_3476,N_49994,N_49985);
and UO_3477 (O_3477,N_49964,N_49971);
nor UO_3478 (O_3478,N_49789,N_49942);
and UO_3479 (O_3479,N_49759,N_49823);
xor UO_3480 (O_3480,N_49800,N_49851);
or UO_3481 (O_3481,N_49870,N_49846);
and UO_3482 (O_3482,N_49961,N_49818);
or UO_3483 (O_3483,N_49773,N_49881);
xor UO_3484 (O_3484,N_49772,N_49760);
nand UO_3485 (O_3485,N_49778,N_49873);
xnor UO_3486 (O_3486,N_49858,N_49828);
xor UO_3487 (O_3487,N_49880,N_49767);
nor UO_3488 (O_3488,N_49819,N_49834);
or UO_3489 (O_3489,N_49862,N_49790);
or UO_3490 (O_3490,N_49753,N_49914);
nor UO_3491 (O_3491,N_49803,N_49779);
and UO_3492 (O_3492,N_49948,N_49832);
or UO_3493 (O_3493,N_49826,N_49777);
and UO_3494 (O_3494,N_49930,N_49974);
nor UO_3495 (O_3495,N_49757,N_49857);
or UO_3496 (O_3496,N_49856,N_49885);
xor UO_3497 (O_3497,N_49838,N_49963);
or UO_3498 (O_3498,N_49966,N_49924);
nor UO_3499 (O_3499,N_49855,N_49936);
or UO_3500 (O_3500,N_49907,N_49867);
xor UO_3501 (O_3501,N_49991,N_49933);
and UO_3502 (O_3502,N_49813,N_49841);
or UO_3503 (O_3503,N_49933,N_49751);
xnor UO_3504 (O_3504,N_49885,N_49870);
xnor UO_3505 (O_3505,N_49942,N_49831);
and UO_3506 (O_3506,N_49945,N_49838);
nand UO_3507 (O_3507,N_49761,N_49981);
and UO_3508 (O_3508,N_49896,N_49789);
nand UO_3509 (O_3509,N_49918,N_49763);
or UO_3510 (O_3510,N_49787,N_49769);
or UO_3511 (O_3511,N_49942,N_49859);
xnor UO_3512 (O_3512,N_49967,N_49861);
or UO_3513 (O_3513,N_49857,N_49829);
xor UO_3514 (O_3514,N_49927,N_49993);
or UO_3515 (O_3515,N_49965,N_49998);
or UO_3516 (O_3516,N_49755,N_49991);
and UO_3517 (O_3517,N_49813,N_49895);
nand UO_3518 (O_3518,N_49976,N_49948);
nand UO_3519 (O_3519,N_49942,N_49795);
xnor UO_3520 (O_3520,N_49796,N_49863);
nor UO_3521 (O_3521,N_49943,N_49990);
nor UO_3522 (O_3522,N_49880,N_49770);
or UO_3523 (O_3523,N_49767,N_49830);
nand UO_3524 (O_3524,N_49779,N_49997);
nor UO_3525 (O_3525,N_49849,N_49965);
xnor UO_3526 (O_3526,N_49921,N_49931);
nand UO_3527 (O_3527,N_49834,N_49779);
xor UO_3528 (O_3528,N_49805,N_49902);
nand UO_3529 (O_3529,N_49993,N_49954);
nor UO_3530 (O_3530,N_49928,N_49883);
nand UO_3531 (O_3531,N_49970,N_49945);
nand UO_3532 (O_3532,N_49777,N_49856);
xnor UO_3533 (O_3533,N_49753,N_49926);
and UO_3534 (O_3534,N_49762,N_49924);
nor UO_3535 (O_3535,N_49922,N_49795);
or UO_3536 (O_3536,N_49796,N_49948);
and UO_3537 (O_3537,N_49892,N_49948);
xnor UO_3538 (O_3538,N_49958,N_49862);
xnor UO_3539 (O_3539,N_49854,N_49888);
or UO_3540 (O_3540,N_49915,N_49923);
xnor UO_3541 (O_3541,N_49980,N_49861);
nand UO_3542 (O_3542,N_49917,N_49776);
or UO_3543 (O_3543,N_49829,N_49955);
nor UO_3544 (O_3544,N_49844,N_49974);
nand UO_3545 (O_3545,N_49759,N_49867);
and UO_3546 (O_3546,N_49925,N_49780);
nor UO_3547 (O_3547,N_49977,N_49916);
nor UO_3548 (O_3548,N_49912,N_49758);
nor UO_3549 (O_3549,N_49803,N_49797);
xor UO_3550 (O_3550,N_49771,N_49848);
nand UO_3551 (O_3551,N_49851,N_49815);
and UO_3552 (O_3552,N_49880,N_49874);
nor UO_3553 (O_3553,N_49800,N_49792);
and UO_3554 (O_3554,N_49769,N_49852);
or UO_3555 (O_3555,N_49797,N_49752);
nand UO_3556 (O_3556,N_49897,N_49990);
nand UO_3557 (O_3557,N_49952,N_49898);
xnor UO_3558 (O_3558,N_49933,N_49982);
nand UO_3559 (O_3559,N_49802,N_49773);
or UO_3560 (O_3560,N_49950,N_49892);
or UO_3561 (O_3561,N_49773,N_49956);
and UO_3562 (O_3562,N_49967,N_49909);
nor UO_3563 (O_3563,N_49805,N_49784);
xnor UO_3564 (O_3564,N_49778,N_49950);
or UO_3565 (O_3565,N_49894,N_49870);
xnor UO_3566 (O_3566,N_49905,N_49997);
or UO_3567 (O_3567,N_49882,N_49782);
and UO_3568 (O_3568,N_49795,N_49841);
and UO_3569 (O_3569,N_49973,N_49816);
and UO_3570 (O_3570,N_49760,N_49851);
xor UO_3571 (O_3571,N_49847,N_49837);
nor UO_3572 (O_3572,N_49929,N_49981);
nand UO_3573 (O_3573,N_49844,N_49833);
or UO_3574 (O_3574,N_49869,N_49991);
or UO_3575 (O_3575,N_49985,N_49829);
nor UO_3576 (O_3576,N_49955,N_49877);
xor UO_3577 (O_3577,N_49886,N_49783);
or UO_3578 (O_3578,N_49971,N_49982);
nor UO_3579 (O_3579,N_49883,N_49952);
xor UO_3580 (O_3580,N_49932,N_49982);
and UO_3581 (O_3581,N_49936,N_49897);
nand UO_3582 (O_3582,N_49969,N_49851);
or UO_3583 (O_3583,N_49908,N_49792);
or UO_3584 (O_3584,N_49751,N_49996);
and UO_3585 (O_3585,N_49979,N_49772);
nand UO_3586 (O_3586,N_49751,N_49822);
nand UO_3587 (O_3587,N_49934,N_49986);
or UO_3588 (O_3588,N_49889,N_49823);
xor UO_3589 (O_3589,N_49765,N_49794);
xor UO_3590 (O_3590,N_49853,N_49839);
nor UO_3591 (O_3591,N_49785,N_49979);
xor UO_3592 (O_3592,N_49932,N_49984);
nor UO_3593 (O_3593,N_49881,N_49776);
xor UO_3594 (O_3594,N_49822,N_49900);
or UO_3595 (O_3595,N_49758,N_49809);
and UO_3596 (O_3596,N_49878,N_49830);
nor UO_3597 (O_3597,N_49865,N_49911);
xnor UO_3598 (O_3598,N_49999,N_49758);
or UO_3599 (O_3599,N_49915,N_49988);
and UO_3600 (O_3600,N_49753,N_49948);
and UO_3601 (O_3601,N_49989,N_49962);
xnor UO_3602 (O_3602,N_49979,N_49977);
nor UO_3603 (O_3603,N_49978,N_49818);
xnor UO_3604 (O_3604,N_49886,N_49855);
and UO_3605 (O_3605,N_49795,N_49917);
nand UO_3606 (O_3606,N_49751,N_49854);
nand UO_3607 (O_3607,N_49951,N_49939);
nand UO_3608 (O_3608,N_49834,N_49816);
xnor UO_3609 (O_3609,N_49801,N_49970);
nand UO_3610 (O_3610,N_49775,N_49898);
nand UO_3611 (O_3611,N_49949,N_49976);
and UO_3612 (O_3612,N_49909,N_49895);
nor UO_3613 (O_3613,N_49972,N_49841);
or UO_3614 (O_3614,N_49757,N_49756);
and UO_3615 (O_3615,N_49812,N_49778);
nor UO_3616 (O_3616,N_49865,N_49904);
and UO_3617 (O_3617,N_49776,N_49977);
and UO_3618 (O_3618,N_49796,N_49803);
nor UO_3619 (O_3619,N_49911,N_49917);
and UO_3620 (O_3620,N_49781,N_49878);
nor UO_3621 (O_3621,N_49783,N_49847);
nand UO_3622 (O_3622,N_49970,N_49878);
nor UO_3623 (O_3623,N_49931,N_49847);
or UO_3624 (O_3624,N_49916,N_49788);
or UO_3625 (O_3625,N_49859,N_49849);
xor UO_3626 (O_3626,N_49823,N_49871);
and UO_3627 (O_3627,N_49846,N_49752);
xor UO_3628 (O_3628,N_49976,N_49966);
nor UO_3629 (O_3629,N_49801,N_49849);
and UO_3630 (O_3630,N_49875,N_49769);
and UO_3631 (O_3631,N_49847,N_49770);
nand UO_3632 (O_3632,N_49791,N_49888);
nand UO_3633 (O_3633,N_49892,N_49880);
or UO_3634 (O_3634,N_49750,N_49765);
and UO_3635 (O_3635,N_49860,N_49984);
or UO_3636 (O_3636,N_49971,N_49977);
nand UO_3637 (O_3637,N_49934,N_49809);
or UO_3638 (O_3638,N_49765,N_49871);
nor UO_3639 (O_3639,N_49859,N_49909);
nand UO_3640 (O_3640,N_49820,N_49930);
nor UO_3641 (O_3641,N_49766,N_49969);
or UO_3642 (O_3642,N_49970,N_49753);
and UO_3643 (O_3643,N_49990,N_49825);
nor UO_3644 (O_3644,N_49772,N_49845);
nand UO_3645 (O_3645,N_49922,N_49976);
nand UO_3646 (O_3646,N_49968,N_49847);
nor UO_3647 (O_3647,N_49973,N_49875);
nand UO_3648 (O_3648,N_49896,N_49947);
or UO_3649 (O_3649,N_49771,N_49896);
nor UO_3650 (O_3650,N_49916,N_49898);
or UO_3651 (O_3651,N_49906,N_49799);
or UO_3652 (O_3652,N_49892,N_49907);
and UO_3653 (O_3653,N_49877,N_49797);
nand UO_3654 (O_3654,N_49852,N_49820);
or UO_3655 (O_3655,N_49957,N_49881);
nor UO_3656 (O_3656,N_49872,N_49762);
and UO_3657 (O_3657,N_49878,N_49820);
nor UO_3658 (O_3658,N_49839,N_49915);
nand UO_3659 (O_3659,N_49770,N_49935);
or UO_3660 (O_3660,N_49992,N_49995);
or UO_3661 (O_3661,N_49845,N_49820);
nand UO_3662 (O_3662,N_49987,N_49968);
nand UO_3663 (O_3663,N_49965,N_49887);
nand UO_3664 (O_3664,N_49867,N_49761);
or UO_3665 (O_3665,N_49900,N_49755);
and UO_3666 (O_3666,N_49869,N_49771);
xor UO_3667 (O_3667,N_49997,N_49795);
and UO_3668 (O_3668,N_49890,N_49897);
nor UO_3669 (O_3669,N_49792,N_49813);
or UO_3670 (O_3670,N_49762,N_49843);
nand UO_3671 (O_3671,N_49864,N_49858);
or UO_3672 (O_3672,N_49864,N_49757);
nand UO_3673 (O_3673,N_49798,N_49990);
and UO_3674 (O_3674,N_49875,N_49761);
or UO_3675 (O_3675,N_49988,N_49772);
and UO_3676 (O_3676,N_49963,N_49793);
and UO_3677 (O_3677,N_49987,N_49757);
nand UO_3678 (O_3678,N_49955,N_49981);
nor UO_3679 (O_3679,N_49956,N_49925);
nor UO_3680 (O_3680,N_49957,N_49986);
and UO_3681 (O_3681,N_49882,N_49996);
nand UO_3682 (O_3682,N_49841,N_49991);
xor UO_3683 (O_3683,N_49856,N_49932);
and UO_3684 (O_3684,N_49953,N_49855);
or UO_3685 (O_3685,N_49864,N_49852);
and UO_3686 (O_3686,N_49998,N_49895);
or UO_3687 (O_3687,N_49803,N_49902);
nor UO_3688 (O_3688,N_49780,N_49834);
nor UO_3689 (O_3689,N_49823,N_49879);
nor UO_3690 (O_3690,N_49769,N_49891);
and UO_3691 (O_3691,N_49820,N_49889);
and UO_3692 (O_3692,N_49907,N_49967);
or UO_3693 (O_3693,N_49751,N_49781);
nand UO_3694 (O_3694,N_49927,N_49774);
nor UO_3695 (O_3695,N_49984,N_49987);
nor UO_3696 (O_3696,N_49837,N_49959);
or UO_3697 (O_3697,N_49975,N_49917);
or UO_3698 (O_3698,N_49916,N_49756);
or UO_3699 (O_3699,N_49987,N_49842);
and UO_3700 (O_3700,N_49865,N_49786);
xor UO_3701 (O_3701,N_49789,N_49796);
xnor UO_3702 (O_3702,N_49981,N_49787);
and UO_3703 (O_3703,N_49776,N_49849);
nor UO_3704 (O_3704,N_49918,N_49990);
nand UO_3705 (O_3705,N_49899,N_49844);
nor UO_3706 (O_3706,N_49767,N_49785);
nand UO_3707 (O_3707,N_49814,N_49873);
or UO_3708 (O_3708,N_49796,N_49827);
nor UO_3709 (O_3709,N_49973,N_49828);
or UO_3710 (O_3710,N_49759,N_49819);
xor UO_3711 (O_3711,N_49864,N_49870);
nor UO_3712 (O_3712,N_49835,N_49938);
and UO_3713 (O_3713,N_49974,N_49836);
xor UO_3714 (O_3714,N_49942,N_49845);
and UO_3715 (O_3715,N_49840,N_49880);
xor UO_3716 (O_3716,N_49890,N_49829);
and UO_3717 (O_3717,N_49771,N_49933);
xnor UO_3718 (O_3718,N_49851,N_49864);
xor UO_3719 (O_3719,N_49844,N_49822);
and UO_3720 (O_3720,N_49852,N_49889);
nand UO_3721 (O_3721,N_49961,N_49751);
xnor UO_3722 (O_3722,N_49928,N_49957);
xnor UO_3723 (O_3723,N_49945,N_49788);
and UO_3724 (O_3724,N_49800,N_49886);
nor UO_3725 (O_3725,N_49794,N_49778);
nand UO_3726 (O_3726,N_49957,N_49776);
and UO_3727 (O_3727,N_49950,N_49863);
and UO_3728 (O_3728,N_49950,N_49944);
xnor UO_3729 (O_3729,N_49810,N_49870);
and UO_3730 (O_3730,N_49874,N_49905);
nand UO_3731 (O_3731,N_49837,N_49804);
nand UO_3732 (O_3732,N_49980,N_49826);
nor UO_3733 (O_3733,N_49833,N_49990);
xor UO_3734 (O_3734,N_49869,N_49936);
and UO_3735 (O_3735,N_49942,N_49945);
nand UO_3736 (O_3736,N_49983,N_49985);
and UO_3737 (O_3737,N_49930,N_49966);
nand UO_3738 (O_3738,N_49853,N_49916);
nand UO_3739 (O_3739,N_49874,N_49907);
xor UO_3740 (O_3740,N_49789,N_49991);
xnor UO_3741 (O_3741,N_49902,N_49855);
nor UO_3742 (O_3742,N_49756,N_49767);
nor UO_3743 (O_3743,N_49764,N_49846);
nor UO_3744 (O_3744,N_49814,N_49771);
or UO_3745 (O_3745,N_49864,N_49860);
nand UO_3746 (O_3746,N_49845,N_49783);
nor UO_3747 (O_3747,N_49936,N_49874);
or UO_3748 (O_3748,N_49873,N_49937);
nand UO_3749 (O_3749,N_49906,N_49785);
nand UO_3750 (O_3750,N_49939,N_49921);
xor UO_3751 (O_3751,N_49888,N_49915);
nand UO_3752 (O_3752,N_49764,N_49816);
nor UO_3753 (O_3753,N_49910,N_49831);
and UO_3754 (O_3754,N_49946,N_49875);
xor UO_3755 (O_3755,N_49780,N_49940);
nand UO_3756 (O_3756,N_49821,N_49912);
xor UO_3757 (O_3757,N_49874,N_49788);
nor UO_3758 (O_3758,N_49766,N_49938);
and UO_3759 (O_3759,N_49830,N_49956);
nand UO_3760 (O_3760,N_49941,N_49913);
or UO_3761 (O_3761,N_49895,N_49806);
xor UO_3762 (O_3762,N_49865,N_49767);
nand UO_3763 (O_3763,N_49994,N_49947);
nand UO_3764 (O_3764,N_49754,N_49885);
and UO_3765 (O_3765,N_49959,N_49862);
and UO_3766 (O_3766,N_49780,N_49983);
nor UO_3767 (O_3767,N_49901,N_49803);
or UO_3768 (O_3768,N_49981,N_49765);
nand UO_3769 (O_3769,N_49823,N_49935);
or UO_3770 (O_3770,N_49870,N_49884);
or UO_3771 (O_3771,N_49797,N_49934);
or UO_3772 (O_3772,N_49917,N_49820);
nand UO_3773 (O_3773,N_49822,N_49810);
xor UO_3774 (O_3774,N_49912,N_49869);
nor UO_3775 (O_3775,N_49807,N_49766);
nor UO_3776 (O_3776,N_49809,N_49782);
nor UO_3777 (O_3777,N_49859,N_49936);
or UO_3778 (O_3778,N_49922,N_49960);
nor UO_3779 (O_3779,N_49809,N_49792);
nor UO_3780 (O_3780,N_49975,N_49887);
and UO_3781 (O_3781,N_49967,N_49970);
and UO_3782 (O_3782,N_49939,N_49902);
nor UO_3783 (O_3783,N_49931,N_49808);
or UO_3784 (O_3784,N_49969,N_49785);
nor UO_3785 (O_3785,N_49974,N_49862);
xnor UO_3786 (O_3786,N_49869,N_49843);
xor UO_3787 (O_3787,N_49831,N_49892);
nand UO_3788 (O_3788,N_49814,N_49857);
and UO_3789 (O_3789,N_49938,N_49905);
or UO_3790 (O_3790,N_49922,N_49759);
and UO_3791 (O_3791,N_49976,N_49909);
xnor UO_3792 (O_3792,N_49873,N_49905);
nor UO_3793 (O_3793,N_49821,N_49883);
xnor UO_3794 (O_3794,N_49773,N_49866);
nor UO_3795 (O_3795,N_49832,N_49881);
and UO_3796 (O_3796,N_49837,N_49880);
or UO_3797 (O_3797,N_49994,N_49961);
nor UO_3798 (O_3798,N_49904,N_49802);
nand UO_3799 (O_3799,N_49765,N_49976);
nand UO_3800 (O_3800,N_49781,N_49977);
nand UO_3801 (O_3801,N_49886,N_49926);
xor UO_3802 (O_3802,N_49953,N_49979);
or UO_3803 (O_3803,N_49769,N_49966);
nor UO_3804 (O_3804,N_49867,N_49795);
nand UO_3805 (O_3805,N_49791,N_49905);
and UO_3806 (O_3806,N_49865,N_49891);
or UO_3807 (O_3807,N_49943,N_49757);
and UO_3808 (O_3808,N_49835,N_49927);
or UO_3809 (O_3809,N_49787,N_49810);
and UO_3810 (O_3810,N_49821,N_49769);
and UO_3811 (O_3811,N_49853,N_49954);
nand UO_3812 (O_3812,N_49890,N_49939);
or UO_3813 (O_3813,N_49846,N_49953);
and UO_3814 (O_3814,N_49946,N_49870);
nand UO_3815 (O_3815,N_49763,N_49777);
xnor UO_3816 (O_3816,N_49912,N_49989);
nor UO_3817 (O_3817,N_49935,N_49864);
nand UO_3818 (O_3818,N_49771,N_49849);
or UO_3819 (O_3819,N_49750,N_49797);
xor UO_3820 (O_3820,N_49813,N_49961);
or UO_3821 (O_3821,N_49917,N_49837);
and UO_3822 (O_3822,N_49919,N_49826);
and UO_3823 (O_3823,N_49778,N_49943);
nor UO_3824 (O_3824,N_49818,N_49976);
nor UO_3825 (O_3825,N_49913,N_49796);
or UO_3826 (O_3826,N_49915,N_49945);
nor UO_3827 (O_3827,N_49781,N_49918);
nor UO_3828 (O_3828,N_49783,N_49813);
nor UO_3829 (O_3829,N_49997,N_49996);
and UO_3830 (O_3830,N_49765,N_49915);
or UO_3831 (O_3831,N_49850,N_49904);
nor UO_3832 (O_3832,N_49799,N_49781);
xor UO_3833 (O_3833,N_49984,N_49976);
nand UO_3834 (O_3834,N_49934,N_49977);
xnor UO_3835 (O_3835,N_49878,N_49854);
and UO_3836 (O_3836,N_49882,N_49794);
xnor UO_3837 (O_3837,N_49863,N_49799);
nor UO_3838 (O_3838,N_49863,N_49775);
nand UO_3839 (O_3839,N_49979,N_49813);
or UO_3840 (O_3840,N_49997,N_49868);
or UO_3841 (O_3841,N_49967,N_49843);
or UO_3842 (O_3842,N_49811,N_49791);
and UO_3843 (O_3843,N_49968,N_49947);
nor UO_3844 (O_3844,N_49771,N_49780);
xor UO_3845 (O_3845,N_49949,N_49959);
and UO_3846 (O_3846,N_49935,N_49863);
nand UO_3847 (O_3847,N_49883,N_49790);
or UO_3848 (O_3848,N_49918,N_49812);
nor UO_3849 (O_3849,N_49870,N_49959);
and UO_3850 (O_3850,N_49946,N_49958);
xor UO_3851 (O_3851,N_49844,N_49970);
xnor UO_3852 (O_3852,N_49819,N_49871);
and UO_3853 (O_3853,N_49960,N_49937);
nor UO_3854 (O_3854,N_49911,N_49762);
nand UO_3855 (O_3855,N_49798,N_49956);
xor UO_3856 (O_3856,N_49817,N_49822);
nand UO_3857 (O_3857,N_49939,N_49780);
nor UO_3858 (O_3858,N_49892,N_49760);
xnor UO_3859 (O_3859,N_49900,N_49914);
and UO_3860 (O_3860,N_49859,N_49763);
nor UO_3861 (O_3861,N_49925,N_49985);
or UO_3862 (O_3862,N_49800,N_49793);
nand UO_3863 (O_3863,N_49901,N_49874);
xnor UO_3864 (O_3864,N_49772,N_49850);
nor UO_3865 (O_3865,N_49990,N_49912);
xnor UO_3866 (O_3866,N_49803,N_49849);
and UO_3867 (O_3867,N_49916,N_49777);
xnor UO_3868 (O_3868,N_49939,N_49968);
nor UO_3869 (O_3869,N_49969,N_49976);
and UO_3870 (O_3870,N_49800,N_49997);
and UO_3871 (O_3871,N_49862,N_49840);
and UO_3872 (O_3872,N_49853,N_49995);
nor UO_3873 (O_3873,N_49912,N_49828);
and UO_3874 (O_3874,N_49856,N_49880);
or UO_3875 (O_3875,N_49805,N_49930);
xor UO_3876 (O_3876,N_49803,N_49909);
nand UO_3877 (O_3877,N_49950,N_49840);
nand UO_3878 (O_3878,N_49865,N_49861);
nand UO_3879 (O_3879,N_49847,N_49910);
and UO_3880 (O_3880,N_49879,N_49787);
nand UO_3881 (O_3881,N_49945,N_49963);
xnor UO_3882 (O_3882,N_49830,N_49953);
and UO_3883 (O_3883,N_49995,N_49981);
and UO_3884 (O_3884,N_49886,N_49831);
nor UO_3885 (O_3885,N_49824,N_49879);
or UO_3886 (O_3886,N_49797,N_49993);
nor UO_3887 (O_3887,N_49786,N_49906);
and UO_3888 (O_3888,N_49845,N_49788);
or UO_3889 (O_3889,N_49764,N_49926);
and UO_3890 (O_3890,N_49856,N_49982);
nand UO_3891 (O_3891,N_49908,N_49793);
nand UO_3892 (O_3892,N_49861,N_49849);
nor UO_3893 (O_3893,N_49844,N_49983);
nor UO_3894 (O_3894,N_49882,N_49824);
xnor UO_3895 (O_3895,N_49816,N_49962);
nor UO_3896 (O_3896,N_49875,N_49752);
xor UO_3897 (O_3897,N_49911,N_49984);
xor UO_3898 (O_3898,N_49800,N_49894);
nor UO_3899 (O_3899,N_49977,N_49768);
xor UO_3900 (O_3900,N_49978,N_49792);
and UO_3901 (O_3901,N_49812,N_49898);
nor UO_3902 (O_3902,N_49803,N_49989);
or UO_3903 (O_3903,N_49881,N_49785);
nand UO_3904 (O_3904,N_49907,N_49944);
or UO_3905 (O_3905,N_49877,N_49840);
xor UO_3906 (O_3906,N_49989,N_49825);
or UO_3907 (O_3907,N_49927,N_49954);
xnor UO_3908 (O_3908,N_49817,N_49841);
and UO_3909 (O_3909,N_49782,N_49868);
xnor UO_3910 (O_3910,N_49756,N_49873);
and UO_3911 (O_3911,N_49987,N_49787);
xor UO_3912 (O_3912,N_49957,N_49959);
or UO_3913 (O_3913,N_49981,N_49954);
nand UO_3914 (O_3914,N_49843,N_49764);
or UO_3915 (O_3915,N_49856,N_49987);
nand UO_3916 (O_3916,N_49796,N_49770);
or UO_3917 (O_3917,N_49882,N_49775);
xnor UO_3918 (O_3918,N_49929,N_49809);
nor UO_3919 (O_3919,N_49893,N_49957);
and UO_3920 (O_3920,N_49994,N_49866);
nand UO_3921 (O_3921,N_49802,N_49816);
xnor UO_3922 (O_3922,N_49970,N_49754);
or UO_3923 (O_3923,N_49811,N_49940);
nand UO_3924 (O_3924,N_49954,N_49767);
and UO_3925 (O_3925,N_49920,N_49787);
xor UO_3926 (O_3926,N_49891,N_49955);
xnor UO_3927 (O_3927,N_49857,N_49970);
nand UO_3928 (O_3928,N_49907,N_49884);
or UO_3929 (O_3929,N_49978,N_49930);
nand UO_3930 (O_3930,N_49758,N_49848);
or UO_3931 (O_3931,N_49856,N_49950);
nor UO_3932 (O_3932,N_49753,N_49904);
or UO_3933 (O_3933,N_49826,N_49782);
and UO_3934 (O_3934,N_49811,N_49877);
xnor UO_3935 (O_3935,N_49783,N_49802);
xor UO_3936 (O_3936,N_49943,N_49999);
or UO_3937 (O_3937,N_49899,N_49900);
xor UO_3938 (O_3938,N_49868,N_49865);
and UO_3939 (O_3939,N_49927,N_49780);
xor UO_3940 (O_3940,N_49799,N_49973);
and UO_3941 (O_3941,N_49776,N_49993);
nor UO_3942 (O_3942,N_49873,N_49836);
nand UO_3943 (O_3943,N_49892,N_49826);
nand UO_3944 (O_3944,N_49817,N_49773);
nand UO_3945 (O_3945,N_49855,N_49806);
nand UO_3946 (O_3946,N_49853,N_49902);
and UO_3947 (O_3947,N_49898,N_49969);
or UO_3948 (O_3948,N_49964,N_49768);
xnor UO_3949 (O_3949,N_49993,N_49823);
and UO_3950 (O_3950,N_49912,N_49777);
xnor UO_3951 (O_3951,N_49998,N_49838);
xnor UO_3952 (O_3952,N_49868,N_49781);
nor UO_3953 (O_3953,N_49804,N_49975);
and UO_3954 (O_3954,N_49772,N_49932);
xnor UO_3955 (O_3955,N_49897,N_49883);
nor UO_3956 (O_3956,N_49758,N_49900);
and UO_3957 (O_3957,N_49802,N_49913);
nor UO_3958 (O_3958,N_49867,N_49804);
xnor UO_3959 (O_3959,N_49789,N_49969);
nand UO_3960 (O_3960,N_49812,N_49951);
xnor UO_3961 (O_3961,N_49972,N_49754);
nor UO_3962 (O_3962,N_49754,N_49934);
and UO_3963 (O_3963,N_49870,N_49782);
and UO_3964 (O_3964,N_49918,N_49878);
xnor UO_3965 (O_3965,N_49848,N_49857);
and UO_3966 (O_3966,N_49850,N_49881);
or UO_3967 (O_3967,N_49816,N_49922);
and UO_3968 (O_3968,N_49877,N_49908);
xor UO_3969 (O_3969,N_49917,N_49848);
or UO_3970 (O_3970,N_49750,N_49922);
and UO_3971 (O_3971,N_49996,N_49990);
nor UO_3972 (O_3972,N_49818,N_49829);
nor UO_3973 (O_3973,N_49965,N_49790);
or UO_3974 (O_3974,N_49970,N_49846);
or UO_3975 (O_3975,N_49808,N_49940);
xor UO_3976 (O_3976,N_49831,N_49868);
nand UO_3977 (O_3977,N_49794,N_49782);
or UO_3978 (O_3978,N_49785,N_49958);
xor UO_3979 (O_3979,N_49787,N_49871);
and UO_3980 (O_3980,N_49963,N_49969);
xor UO_3981 (O_3981,N_49983,N_49936);
nand UO_3982 (O_3982,N_49899,N_49758);
xnor UO_3983 (O_3983,N_49862,N_49861);
nand UO_3984 (O_3984,N_49802,N_49859);
xnor UO_3985 (O_3985,N_49970,N_49758);
xnor UO_3986 (O_3986,N_49969,N_49865);
xnor UO_3987 (O_3987,N_49818,N_49824);
nor UO_3988 (O_3988,N_49873,N_49844);
or UO_3989 (O_3989,N_49827,N_49950);
and UO_3990 (O_3990,N_49802,N_49894);
xor UO_3991 (O_3991,N_49834,N_49771);
nor UO_3992 (O_3992,N_49775,N_49843);
nand UO_3993 (O_3993,N_49774,N_49903);
nor UO_3994 (O_3994,N_49859,N_49798);
or UO_3995 (O_3995,N_49833,N_49901);
or UO_3996 (O_3996,N_49916,N_49828);
xnor UO_3997 (O_3997,N_49782,N_49962);
nand UO_3998 (O_3998,N_49975,N_49790);
nand UO_3999 (O_3999,N_49801,N_49930);
nor UO_4000 (O_4000,N_49765,N_49942);
and UO_4001 (O_4001,N_49988,N_49857);
or UO_4002 (O_4002,N_49869,N_49849);
xor UO_4003 (O_4003,N_49990,N_49864);
and UO_4004 (O_4004,N_49848,N_49897);
xor UO_4005 (O_4005,N_49854,N_49758);
nor UO_4006 (O_4006,N_49889,N_49831);
nand UO_4007 (O_4007,N_49943,N_49870);
and UO_4008 (O_4008,N_49779,N_49932);
or UO_4009 (O_4009,N_49852,N_49936);
nor UO_4010 (O_4010,N_49899,N_49891);
nor UO_4011 (O_4011,N_49974,N_49817);
or UO_4012 (O_4012,N_49887,N_49931);
nor UO_4013 (O_4013,N_49924,N_49835);
or UO_4014 (O_4014,N_49902,N_49821);
nand UO_4015 (O_4015,N_49754,N_49788);
and UO_4016 (O_4016,N_49775,N_49972);
nand UO_4017 (O_4017,N_49952,N_49861);
xnor UO_4018 (O_4018,N_49938,N_49935);
nand UO_4019 (O_4019,N_49864,N_49950);
nor UO_4020 (O_4020,N_49862,N_49863);
and UO_4021 (O_4021,N_49968,N_49949);
nand UO_4022 (O_4022,N_49891,N_49945);
xnor UO_4023 (O_4023,N_49838,N_49874);
xor UO_4024 (O_4024,N_49930,N_49779);
nor UO_4025 (O_4025,N_49897,N_49944);
nor UO_4026 (O_4026,N_49781,N_49844);
nand UO_4027 (O_4027,N_49830,N_49929);
nand UO_4028 (O_4028,N_49831,N_49828);
nand UO_4029 (O_4029,N_49784,N_49750);
or UO_4030 (O_4030,N_49821,N_49996);
and UO_4031 (O_4031,N_49804,N_49851);
and UO_4032 (O_4032,N_49793,N_49779);
xnor UO_4033 (O_4033,N_49784,N_49948);
and UO_4034 (O_4034,N_49904,N_49751);
nand UO_4035 (O_4035,N_49808,N_49840);
and UO_4036 (O_4036,N_49859,N_49842);
nand UO_4037 (O_4037,N_49879,N_49888);
nor UO_4038 (O_4038,N_49978,N_49964);
xnor UO_4039 (O_4039,N_49948,N_49940);
or UO_4040 (O_4040,N_49942,N_49830);
or UO_4041 (O_4041,N_49947,N_49799);
and UO_4042 (O_4042,N_49875,N_49936);
or UO_4043 (O_4043,N_49922,N_49959);
or UO_4044 (O_4044,N_49948,N_49826);
or UO_4045 (O_4045,N_49818,N_49885);
xor UO_4046 (O_4046,N_49841,N_49870);
nand UO_4047 (O_4047,N_49902,N_49822);
and UO_4048 (O_4048,N_49938,N_49923);
and UO_4049 (O_4049,N_49987,N_49868);
xnor UO_4050 (O_4050,N_49869,N_49845);
nor UO_4051 (O_4051,N_49892,N_49927);
nand UO_4052 (O_4052,N_49993,N_49794);
and UO_4053 (O_4053,N_49873,N_49909);
or UO_4054 (O_4054,N_49867,N_49976);
nor UO_4055 (O_4055,N_49754,N_49843);
or UO_4056 (O_4056,N_49927,N_49779);
xnor UO_4057 (O_4057,N_49776,N_49812);
nand UO_4058 (O_4058,N_49910,N_49819);
xor UO_4059 (O_4059,N_49797,N_49991);
xnor UO_4060 (O_4060,N_49938,N_49853);
xnor UO_4061 (O_4061,N_49971,N_49875);
nand UO_4062 (O_4062,N_49955,N_49943);
nand UO_4063 (O_4063,N_49951,N_49857);
or UO_4064 (O_4064,N_49854,N_49785);
or UO_4065 (O_4065,N_49863,N_49854);
and UO_4066 (O_4066,N_49774,N_49922);
and UO_4067 (O_4067,N_49932,N_49832);
nor UO_4068 (O_4068,N_49968,N_49856);
xnor UO_4069 (O_4069,N_49758,N_49921);
xnor UO_4070 (O_4070,N_49940,N_49927);
nand UO_4071 (O_4071,N_49893,N_49853);
nor UO_4072 (O_4072,N_49766,N_49909);
or UO_4073 (O_4073,N_49983,N_49799);
nand UO_4074 (O_4074,N_49751,N_49906);
xor UO_4075 (O_4075,N_49880,N_49993);
and UO_4076 (O_4076,N_49790,N_49777);
and UO_4077 (O_4077,N_49922,N_49786);
xor UO_4078 (O_4078,N_49847,N_49813);
and UO_4079 (O_4079,N_49797,N_49853);
nand UO_4080 (O_4080,N_49876,N_49768);
xor UO_4081 (O_4081,N_49753,N_49806);
nand UO_4082 (O_4082,N_49972,N_49898);
and UO_4083 (O_4083,N_49819,N_49992);
nand UO_4084 (O_4084,N_49864,N_49796);
xor UO_4085 (O_4085,N_49937,N_49863);
and UO_4086 (O_4086,N_49792,N_49807);
xor UO_4087 (O_4087,N_49975,N_49896);
and UO_4088 (O_4088,N_49964,N_49764);
nand UO_4089 (O_4089,N_49976,N_49877);
and UO_4090 (O_4090,N_49802,N_49754);
nor UO_4091 (O_4091,N_49828,N_49766);
xor UO_4092 (O_4092,N_49939,N_49989);
nor UO_4093 (O_4093,N_49877,N_49942);
xor UO_4094 (O_4094,N_49847,N_49860);
or UO_4095 (O_4095,N_49911,N_49791);
or UO_4096 (O_4096,N_49858,N_49909);
nor UO_4097 (O_4097,N_49779,N_49863);
nor UO_4098 (O_4098,N_49773,N_49969);
nand UO_4099 (O_4099,N_49774,N_49929);
or UO_4100 (O_4100,N_49937,N_49772);
nand UO_4101 (O_4101,N_49761,N_49932);
and UO_4102 (O_4102,N_49784,N_49869);
nor UO_4103 (O_4103,N_49892,N_49821);
and UO_4104 (O_4104,N_49921,N_49808);
nand UO_4105 (O_4105,N_49828,N_49819);
or UO_4106 (O_4106,N_49772,N_49757);
nor UO_4107 (O_4107,N_49972,N_49784);
xnor UO_4108 (O_4108,N_49782,N_49902);
and UO_4109 (O_4109,N_49931,N_49929);
nand UO_4110 (O_4110,N_49996,N_49805);
nor UO_4111 (O_4111,N_49790,N_49961);
xor UO_4112 (O_4112,N_49863,N_49908);
nor UO_4113 (O_4113,N_49795,N_49794);
or UO_4114 (O_4114,N_49986,N_49822);
nand UO_4115 (O_4115,N_49848,N_49988);
nand UO_4116 (O_4116,N_49853,N_49818);
nor UO_4117 (O_4117,N_49931,N_49982);
and UO_4118 (O_4118,N_49782,N_49892);
nor UO_4119 (O_4119,N_49873,N_49893);
or UO_4120 (O_4120,N_49860,N_49936);
nand UO_4121 (O_4121,N_49876,N_49797);
nand UO_4122 (O_4122,N_49977,N_49983);
xor UO_4123 (O_4123,N_49769,N_49893);
nand UO_4124 (O_4124,N_49840,N_49932);
xnor UO_4125 (O_4125,N_49896,N_49812);
nor UO_4126 (O_4126,N_49883,N_49809);
and UO_4127 (O_4127,N_49925,N_49779);
or UO_4128 (O_4128,N_49776,N_49893);
nand UO_4129 (O_4129,N_49759,N_49936);
and UO_4130 (O_4130,N_49954,N_49842);
xnor UO_4131 (O_4131,N_49814,N_49830);
xor UO_4132 (O_4132,N_49783,N_49890);
or UO_4133 (O_4133,N_49763,N_49805);
nor UO_4134 (O_4134,N_49947,N_49974);
nor UO_4135 (O_4135,N_49874,N_49987);
nor UO_4136 (O_4136,N_49863,N_49797);
xnor UO_4137 (O_4137,N_49937,N_49826);
xor UO_4138 (O_4138,N_49805,N_49859);
and UO_4139 (O_4139,N_49821,N_49796);
nand UO_4140 (O_4140,N_49842,N_49931);
nand UO_4141 (O_4141,N_49997,N_49823);
xor UO_4142 (O_4142,N_49804,N_49810);
or UO_4143 (O_4143,N_49965,N_49966);
nand UO_4144 (O_4144,N_49792,N_49988);
nand UO_4145 (O_4145,N_49987,N_49876);
or UO_4146 (O_4146,N_49753,N_49929);
nor UO_4147 (O_4147,N_49891,N_49813);
and UO_4148 (O_4148,N_49990,N_49988);
nor UO_4149 (O_4149,N_49968,N_49959);
nand UO_4150 (O_4150,N_49762,N_49910);
and UO_4151 (O_4151,N_49771,N_49755);
and UO_4152 (O_4152,N_49964,N_49952);
nand UO_4153 (O_4153,N_49822,N_49934);
or UO_4154 (O_4154,N_49826,N_49962);
xnor UO_4155 (O_4155,N_49900,N_49961);
nand UO_4156 (O_4156,N_49898,N_49907);
or UO_4157 (O_4157,N_49763,N_49756);
xor UO_4158 (O_4158,N_49953,N_49932);
xor UO_4159 (O_4159,N_49901,N_49887);
nor UO_4160 (O_4160,N_49879,N_49931);
nand UO_4161 (O_4161,N_49824,N_49922);
and UO_4162 (O_4162,N_49911,N_49824);
nand UO_4163 (O_4163,N_49892,N_49773);
or UO_4164 (O_4164,N_49993,N_49855);
nor UO_4165 (O_4165,N_49805,N_49768);
xor UO_4166 (O_4166,N_49762,N_49818);
xnor UO_4167 (O_4167,N_49928,N_49897);
and UO_4168 (O_4168,N_49971,N_49894);
nor UO_4169 (O_4169,N_49943,N_49966);
and UO_4170 (O_4170,N_49945,N_49868);
and UO_4171 (O_4171,N_49991,N_49835);
or UO_4172 (O_4172,N_49888,N_49939);
nand UO_4173 (O_4173,N_49965,N_49891);
or UO_4174 (O_4174,N_49923,N_49993);
nor UO_4175 (O_4175,N_49829,N_49924);
or UO_4176 (O_4176,N_49848,N_49788);
nor UO_4177 (O_4177,N_49999,N_49784);
nor UO_4178 (O_4178,N_49874,N_49852);
and UO_4179 (O_4179,N_49823,N_49775);
and UO_4180 (O_4180,N_49773,N_49848);
and UO_4181 (O_4181,N_49945,N_49948);
and UO_4182 (O_4182,N_49917,N_49831);
or UO_4183 (O_4183,N_49945,N_49764);
nor UO_4184 (O_4184,N_49961,N_49787);
nand UO_4185 (O_4185,N_49851,N_49781);
and UO_4186 (O_4186,N_49920,N_49955);
and UO_4187 (O_4187,N_49886,N_49951);
nand UO_4188 (O_4188,N_49762,N_49813);
nand UO_4189 (O_4189,N_49872,N_49869);
xor UO_4190 (O_4190,N_49795,N_49957);
xor UO_4191 (O_4191,N_49985,N_49813);
xnor UO_4192 (O_4192,N_49833,N_49998);
and UO_4193 (O_4193,N_49934,N_49908);
nand UO_4194 (O_4194,N_49987,N_49833);
nand UO_4195 (O_4195,N_49963,N_49991);
or UO_4196 (O_4196,N_49814,N_49949);
xnor UO_4197 (O_4197,N_49897,N_49987);
nand UO_4198 (O_4198,N_49903,N_49918);
nor UO_4199 (O_4199,N_49931,N_49786);
nand UO_4200 (O_4200,N_49817,N_49882);
nor UO_4201 (O_4201,N_49962,N_49786);
or UO_4202 (O_4202,N_49875,N_49814);
or UO_4203 (O_4203,N_49759,N_49871);
and UO_4204 (O_4204,N_49845,N_49840);
xnor UO_4205 (O_4205,N_49770,N_49842);
nor UO_4206 (O_4206,N_49892,N_49774);
nor UO_4207 (O_4207,N_49886,N_49984);
nand UO_4208 (O_4208,N_49806,N_49921);
nand UO_4209 (O_4209,N_49923,N_49924);
and UO_4210 (O_4210,N_49865,N_49981);
and UO_4211 (O_4211,N_49947,N_49908);
xnor UO_4212 (O_4212,N_49961,N_49860);
and UO_4213 (O_4213,N_49793,N_49932);
nor UO_4214 (O_4214,N_49990,N_49855);
or UO_4215 (O_4215,N_49755,N_49813);
and UO_4216 (O_4216,N_49950,N_49898);
xnor UO_4217 (O_4217,N_49778,N_49934);
nor UO_4218 (O_4218,N_49807,N_49828);
nand UO_4219 (O_4219,N_49788,N_49969);
or UO_4220 (O_4220,N_49965,N_49825);
or UO_4221 (O_4221,N_49945,N_49981);
xor UO_4222 (O_4222,N_49966,N_49949);
nand UO_4223 (O_4223,N_49949,N_49828);
nand UO_4224 (O_4224,N_49807,N_49903);
and UO_4225 (O_4225,N_49851,N_49978);
nand UO_4226 (O_4226,N_49904,N_49768);
or UO_4227 (O_4227,N_49799,N_49757);
xnor UO_4228 (O_4228,N_49850,N_49979);
and UO_4229 (O_4229,N_49861,N_49914);
nor UO_4230 (O_4230,N_49925,N_49982);
or UO_4231 (O_4231,N_49770,N_49779);
or UO_4232 (O_4232,N_49985,N_49750);
xor UO_4233 (O_4233,N_49769,N_49971);
nand UO_4234 (O_4234,N_49751,N_49753);
xor UO_4235 (O_4235,N_49845,N_49754);
nand UO_4236 (O_4236,N_49869,N_49980);
nand UO_4237 (O_4237,N_49999,N_49766);
nor UO_4238 (O_4238,N_49792,N_49833);
nor UO_4239 (O_4239,N_49785,N_49865);
or UO_4240 (O_4240,N_49941,N_49931);
xor UO_4241 (O_4241,N_49774,N_49769);
xor UO_4242 (O_4242,N_49847,N_49869);
nor UO_4243 (O_4243,N_49828,N_49956);
xnor UO_4244 (O_4244,N_49882,N_49776);
nor UO_4245 (O_4245,N_49830,N_49815);
xnor UO_4246 (O_4246,N_49869,N_49916);
and UO_4247 (O_4247,N_49856,N_49758);
and UO_4248 (O_4248,N_49782,N_49836);
nor UO_4249 (O_4249,N_49903,N_49931);
and UO_4250 (O_4250,N_49858,N_49854);
xor UO_4251 (O_4251,N_49953,N_49859);
or UO_4252 (O_4252,N_49981,N_49858);
xnor UO_4253 (O_4253,N_49859,N_49949);
xnor UO_4254 (O_4254,N_49996,N_49774);
nand UO_4255 (O_4255,N_49945,N_49880);
and UO_4256 (O_4256,N_49803,N_49768);
xnor UO_4257 (O_4257,N_49774,N_49877);
and UO_4258 (O_4258,N_49974,N_49860);
xnor UO_4259 (O_4259,N_49859,N_49821);
nand UO_4260 (O_4260,N_49881,N_49927);
xnor UO_4261 (O_4261,N_49847,N_49768);
xnor UO_4262 (O_4262,N_49947,N_49754);
xor UO_4263 (O_4263,N_49869,N_49898);
nand UO_4264 (O_4264,N_49883,N_49843);
and UO_4265 (O_4265,N_49906,N_49850);
nor UO_4266 (O_4266,N_49863,N_49780);
or UO_4267 (O_4267,N_49786,N_49911);
or UO_4268 (O_4268,N_49959,N_49854);
nand UO_4269 (O_4269,N_49793,N_49751);
nor UO_4270 (O_4270,N_49979,N_49875);
nand UO_4271 (O_4271,N_49907,N_49919);
and UO_4272 (O_4272,N_49906,N_49894);
or UO_4273 (O_4273,N_49932,N_49756);
nand UO_4274 (O_4274,N_49884,N_49889);
xor UO_4275 (O_4275,N_49967,N_49939);
and UO_4276 (O_4276,N_49935,N_49990);
nand UO_4277 (O_4277,N_49853,N_49980);
xor UO_4278 (O_4278,N_49925,N_49833);
xnor UO_4279 (O_4279,N_49820,N_49779);
nor UO_4280 (O_4280,N_49919,N_49858);
and UO_4281 (O_4281,N_49809,N_49865);
nor UO_4282 (O_4282,N_49942,N_49820);
nor UO_4283 (O_4283,N_49970,N_49950);
nand UO_4284 (O_4284,N_49779,N_49850);
or UO_4285 (O_4285,N_49870,N_49766);
or UO_4286 (O_4286,N_49841,N_49781);
nand UO_4287 (O_4287,N_49763,N_49864);
nor UO_4288 (O_4288,N_49819,N_49865);
or UO_4289 (O_4289,N_49937,N_49967);
xnor UO_4290 (O_4290,N_49975,N_49908);
and UO_4291 (O_4291,N_49873,N_49810);
nor UO_4292 (O_4292,N_49901,N_49821);
or UO_4293 (O_4293,N_49814,N_49819);
xnor UO_4294 (O_4294,N_49857,N_49843);
nand UO_4295 (O_4295,N_49990,N_49949);
nor UO_4296 (O_4296,N_49932,N_49758);
nand UO_4297 (O_4297,N_49926,N_49818);
xor UO_4298 (O_4298,N_49793,N_49923);
xnor UO_4299 (O_4299,N_49812,N_49899);
and UO_4300 (O_4300,N_49818,N_49954);
xor UO_4301 (O_4301,N_49822,N_49940);
or UO_4302 (O_4302,N_49835,N_49905);
and UO_4303 (O_4303,N_49882,N_49784);
nor UO_4304 (O_4304,N_49812,N_49880);
or UO_4305 (O_4305,N_49817,N_49936);
or UO_4306 (O_4306,N_49777,N_49886);
and UO_4307 (O_4307,N_49889,N_49791);
xor UO_4308 (O_4308,N_49861,N_49879);
nor UO_4309 (O_4309,N_49932,N_49965);
nand UO_4310 (O_4310,N_49801,N_49937);
nor UO_4311 (O_4311,N_49833,N_49940);
xnor UO_4312 (O_4312,N_49895,N_49773);
and UO_4313 (O_4313,N_49901,N_49890);
nor UO_4314 (O_4314,N_49965,N_49945);
and UO_4315 (O_4315,N_49785,N_49891);
and UO_4316 (O_4316,N_49879,N_49842);
xor UO_4317 (O_4317,N_49888,N_49839);
xnor UO_4318 (O_4318,N_49915,N_49775);
xnor UO_4319 (O_4319,N_49987,N_49992);
or UO_4320 (O_4320,N_49849,N_49810);
or UO_4321 (O_4321,N_49986,N_49954);
or UO_4322 (O_4322,N_49921,N_49866);
xor UO_4323 (O_4323,N_49854,N_49786);
and UO_4324 (O_4324,N_49860,N_49909);
nand UO_4325 (O_4325,N_49925,N_49802);
nor UO_4326 (O_4326,N_49799,N_49866);
or UO_4327 (O_4327,N_49818,N_49775);
nand UO_4328 (O_4328,N_49837,N_49920);
nor UO_4329 (O_4329,N_49882,N_49920);
and UO_4330 (O_4330,N_49782,N_49797);
xor UO_4331 (O_4331,N_49991,N_49912);
nor UO_4332 (O_4332,N_49844,N_49979);
and UO_4333 (O_4333,N_49859,N_49815);
and UO_4334 (O_4334,N_49932,N_49795);
xor UO_4335 (O_4335,N_49898,N_49927);
nand UO_4336 (O_4336,N_49792,N_49893);
xor UO_4337 (O_4337,N_49825,N_49903);
and UO_4338 (O_4338,N_49927,N_49908);
nor UO_4339 (O_4339,N_49965,N_49883);
nor UO_4340 (O_4340,N_49783,N_49959);
or UO_4341 (O_4341,N_49870,N_49972);
nand UO_4342 (O_4342,N_49850,N_49972);
nor UO_4343 (O_4343,N_49965,N_49938);
xor UO_4344 (O_4344,N_49861,N_49830);
or UO_4345 (O_4345,N_49951,N_49768);
or UO_4346 (O_4346,N_49772,N_49959);
nand UO_4347 (O_4347,N_49890,N_49954);
and UO_4348 (O_4348,N_49902,N_49843);
xnor UO_4349 (O_4349,N_49802,N_49833);
or UO_4350 (O_4350,N_49824,N_49991);
or UO_4351 (O_4351,N_49793,N_49955);
or UO_4352 (O_4352,N_49915,N_49898);
nor UO_4353 (O_4353,N_49884,N_49954);
xnor UO_4354 (O_4354,N_49956,N_49921);
nand UO_4355 (O_4355,N_49750,N_49915);
nand UO_4356 (O_4356,N_49911,N_49975);
or UO_4357 (O_4357,N_49756,N_49806);
nor UO_4358 (O_4358,N_49784,N_49851);
and UO_4359 (O_4359,N_49805,N_49898);
and UO_4360 (O_4360,N_49772,N_49796);
xor UO_4361 (O_4361,N_49933,N_49953);
and UO_4362 (O_4362,N_49912,N_49857);
nand UO_4363 (O_4363,N_49991,N_49894);
or UO_4364 (O_4364,N_49823,N_49803);
nand UO_4365 (O_4365,N_49999,N_49764);
xor UO_4366 (O_4366,N_49933,N_49977);
nand UO_4367 (O_4367,N_49980,N_49973);
or UO_4368 (O_4368,N_49799,N_49764);
xor UO_4369 (O_4369,N_49893,N_49833);
nand UO_4370 (O_4370,N_49753,N_49917);
nand UO_4371 (O_4371,N_49831,N_49832);
or UO_4372 (O_4372,N_49844,N_49868);
nand UO_4373 (O_4373,N_49920,N_49804);
and UO_4374 (O_4374,N_49839,N_49780);
nor UO_4375 (O_4375,N_49875,N_49987);
and UO_4376 (O_4376,N_49803,N_49827);
nor UO_4377 (O_4377,N_49809,N_49830);
nor UO_4378 (O_4378,N_49915,N_49890);
and UO_4379 (O_4379,N_49807,N_49983);
or UO_4380 (O_4380,N_49917,N_49762);
xor UO_4381 (O_4381,N_49944,N_49833);
nor UO_4382 (O_4382,N_49883,N_49775);
or UO_4383 (O_4383,N_49917,N_49869);
nor UO_4384 (O_4384,N_49928,N_49759);
and UO_4385 (O_4385,N_49752,N_49828);
nor UO_4386 (O_4386,N_49828,N_49820);
or UO_4387 (O_4387,N_49884,N_49774);
nand UO_4388 (O_4388,N_49757,N_49833);
or UO_4389 (O_4389,N_49958,N_49948);
nand UO_4390 (O_4390,N_49833,N_49768);
and UO_4391 (O_4391,N_49819,N_49774);
nor UO_4392 (O_4392,N_49773,N_49935);
nor UO_4393 (O_4393,N_49840,N_49760);
nand UO_4394 (O_4394,N_49923,N_49979);
and UO_4395 (O_4395,N_49775,N_49990);
nor UO_4396 (O_4396,N_49928,N_49935);
xor UO_4397 (O_4397,N_49961,N_49948);
or UO_4398 (O_4398,N_49846,N_49822);
xnor UO_4399 (O_4399,N_49933,N_49861);
nor UO_4400 (O_4400,N_49872,N_49822);
or UO_4401 (O_4401,N_49810,N_49891);
nor UO_4402 (O_4402,N_49948,N_49977);
nor UO_4403 (O_4403,N_49922,N_49970);
and UO_4404 (O_4404,N_49851,N_49923);
nand UO_4405 (O_4405,N_49763,N_49784);
xnor UO_4406 (O_4406,N_49772,N_49934);
nand UO_4407 (O_4407,N_49906,N_49960);
nand UO_4408 (O_4408,N_49921,N_49796);
nand UO_4409 (O_4409,N_49836,N_49912);
and UO_4410 (O_4410,N_49883,N_49764);
xnor UO_4411 (O_4411,N_49856,N_49994);
xor UO_4412 (O_4412,N_49810,N_49904);
nand UO_4413 (O_4413,N_49759,N_49795);
or UO_4414 (O_4414,N_49959,N_49766);
xnor UO_4415 (O_4415,N_49977,N_49975);
or UO_4416 (O_4416,N_49900,N_49879);
and UO_4417 (O_4417,N_49959,N_49967);
and UO_4418 (O_4418,N_49905,N_49895);
nand UO_4419 (O_4419,N_49800,N_49816);
or UO_4420 (O_4420,N_49864,N_49941);
nand UO_4421 (O_4421,N_49966,N_49999);
or UO_4422 (O_4422,N_49975,N_49920);
or UO_4423 (O_4423,N_49871,N_49937);
and UO_4424 (O_4424,N_49917,N_49971);
nor UO_4425 (O_4425,N_49929,N_49909);
xnor UO_4426 (O_4426,N_49935,N_49837);
and UO_4427 (O_4427,N_49905,N_49843);
nor UO_4428 (O_4428,N_49967,N_49791);
and UO_4429 (O_4429,N_49850,N_49874);
nor UO_4430 (O_4430,N_49852,N_49831);
nor UO_4431 (O_4431,N_49882,N_49880);
or UO_4432 (O_4432,N_49765,N_49978);
nand UO_4433 (O_4433,N_49932,N_49815);
nand UO_4434 (O_4434,N_49843,N_49949);
nand UO_4435 (O_4435,N_49977,N_49937);
and UO_4436 (O_4436,N_49802,N_49927);
or UO_4437 (O_4437,N_49758,N_49846);
nor UO_4438 (O_4438,N_49861,N_49775);
or UO_4439 (O_4439,N_49910,N_49972);
xnor UO_4440 (O_4440,N_49847,N_49846);
and UO_4441 (O_4441,N_49965,N_49956);
or UO_4442 (O_4442,N_49960,N_49849);
nand UO_4443 (O_4443,N_49836,N_49772);
xnor UO_4444 (O_4444,N_49843,N_49853);
xor UO_4445 (O_4445,N_49915,N_49979);
xor UO_4446 (O_4446,N_49755,N_49933);
nand UO_4447 (O_4447,N_49909,N_49908);
nand UO_4448 (O_4448,N_49952,N_49766);
nor UO_4449 (O_4449,N_49859,N_49901);
nor UO_4450 (O_4450,N_49796,N_49878);
and UO_4451 (O_4451,N_49870,N_49822);
or UO_4452 (O_4452,N_49924,N_49936);
nand UO_4453 (O_4453,N_49811,N_49955);
or UO_4454 (O_4454,N_49878,N_49843);
nor UO_4455 (O_4455,N_49854,N_49995);
and UO_4456 (O_4456,N_49976,N_49752);
nand UO_4457 (O_4457,N_49864,N_49995);
xor UO_4458 (O_4458,N_49873,N_49866);
and UO_4459 (O_4459,N_49787,N_49914);
xnor UO_4460 (O_4460,N_49928,N_49796);
nor UO_4461 (O_4461,N_49830,N_49962);
or UO_4462 (O_4462,N_49800,N_49763);
nor UO_4463 (O_4463,N_49868,N_49897);
xor UO_4464 (O_4464,N_49933,N_49948);
nor UO_4465 (O_4465,N_49786,N_49789);
xnor UO_4466 (O_4466,N_49836,N_49966);
nor UO_4467 (O_4467,N_49852,N_49765);
xnor UO_4468 (O_4468,N_49943,N_49877);
or UO_4469 (O_4469,N_49751,N_49844);
nand UO_4470 (O_4470,N_49950,N_49874);
xor UO_4471 (O_4471,N_49810,N_49857);
nand UO_4472 (O_4472,N_49793,N_49922);
and UO_4473 (O_4473,N_49881,N_49827);
and UO_4474 (O_4474,N_49908,N_49996);
or UO_4475 (O_4475,N_49965,N_49909);
xor UO_4476 (O_4476,N_49781,N_49805);
or UO_4477 (O_4477,N_49775,N_49914);
nand UO_4478 (O_4478,N_49916,N_49970);
and UO_4479 (O_4479,N_49992,N_49875);
or UO_4480 (O_4480,N_49940,N_49797);
nand UO_4481 (O_4481,N_49769,N_49868);
or UO_4482 (O_4482,N_49759,N_49980);
nor UO_4483 (O_4483,N_49822,N_49835);
xor UO_4484 (O_4484,N_49956,N_49788);
xor UO_4485 (O_4485,N_49932,N_49899);
xor UO_4486 (O_4486,N_49846,N_49826);
or UO_4487 (O_4487,N_49763,N_49970);
nor UO_4488 (O_4488,N_49796,N_49890);
nor UO_4489 (O_4489,N_49805,N_49991);
and UO_4490 (O_4490,N_49839,N_49950);
nand UO_4491 (O_4491,N_49752,N_49952);
or UO_4492 (O_4492,N_49847,N_49921);
and UO_4493 (O_4493,N_49994,N_49788);
xnor UO_4494 (O_4494,N_49877,N_49894);
xor UO_4495 (O_4495,N_49825,N_49847);
or UO_4496 (O_4496,N_49900,N_49979);
nand UO_4497 (O_4497,N_49890,N_49768);
xor UO_4498 (O_4498,N_49795,N_49908);
xnor UO_4499 (O_4499,N_49787,N_49756);
nor UO_4500 (O_4500,N_49923,N_49971);
nand UO_4501 (O_4501,N_49932,N_49783);
or UO_4502 (O_4502,N_49841,N_49881);
and UO_4503 (O_4503,N_49901,N_49889);
nand UO_4504 (O_4504,N_49860,N_49981);
and UO_4505 (O_4505,N_49843,N_49831);
xor UO_4506 (O_4506,N_49794,N_49960);
xnor UO_4507 (O_4507,N_49863,N_49852);
xnor UO_4508 (O_4508,N_49824,N_49948);
or UO_4509 (O_4509,N_49774,N_49843);
nor UO_4510 (O_4510,N_49851,N_49997);
nor UO_4511 (O_4511,N_49894,N_49962);
or UO_4512 (O_4512,N_49872,N_49968);
xor UO_4513 (O_4513,N_49966,N_49887);
or UO_4514 (O_4514,N_49834,N_49782);
and UO_4515 (O_4515,N_49791,N_49966);
or UO_4516 (O_4516,N_49984,N_49818);
nand UO_4517 (O_4517,N_49991,N_49795);
or UO_4518 (O_4518,N_49962,N_49997);
or UO_4519 (O_4519,N_49853,N_49944);
nand UO_4520 (O_4520,N_49758,N_49851);
or UO_4521 (O_4521,N_49811,N_49797);
xnor UO_4522 (O_4522,N_49889,N_49842);
and UO_4523 (O_4523,N_49888,N_49944);
xnor UO_4524 (O_4524,N_49777,N_49880);
nand UO_4525 (O_4525,N_49999,N_49933);
or UO_4526 (O_4526,N_49972,N_49788);
and UO_4527 (O_4527,N_49945,N_49834);
or UO_4528 (O_4528,N_49938,N_49949);
nor UO_4529 (O_4529,N_49803,N_49851);
or UO_4530 (O_4530,N_49815,N_49837);
nor UO_4531 (O_4531,N_49754,N_49786);
nor UO_4532 (O_4532,N_49996,N_49976);
or UO_4533 (O_4533,N_49896,N_49993);
xnor UO_4534 (O_4534,N_49812,N_49767);
or UO_4535 (O_4535,N_49881,N_49945);
nor UO_4536 (O_4536,N_49803,N_49923);
or UO_4537 (O_4537,N_49800,N_49902);
nand UO_4538 (O_4538,N_49988,N_49909);
nor UO_4539 (O_4539,N_49979,N_49888);
nor UO_4540 (O_4540,N_49863,N_49785);
and UO_4541 (O_4541,N_49827,N_49937);
nor UO_4542 (O_4542,N_49861,N_49901);
or UO_4543 (O_4543,N_49983,N_49795);
nand UO_4544 (O_4544,N_49886,N_49940);
or UO_4545 (O_4545,N_49782,N_49867);
nand UO_4546 (O_4546,N_49898,N_49882);
nand UO_4547 (O_4547,N_49920,N_49940);
nor UO_4548 (O_4548,N_49914,N_49827);
or UO_4549 (O_4549,N_49788,N_49914);
and UO_4550 (O_4550,N_49955,N_49794);
and UO_4551 (O_4551,N_49984,N_49972);
nor UO_4552 (O_4552,N_49856,N_49952);
xnor UO_4553 (O_4553,N_49769,N_49755);
nor UO_4554 (O_4554,N_49960,N_49993);
and UO_4555 (O_4555,N_49935,N_49925);
nand UO_4556 (O_4556,N_49775,N_49921);
xor UO_4557 (O_4557,N_49835,N_49800);
or UO_4558 (O_4558,N_49808,N_49985);
xnor UO_4559 (O_4559,N_49937,N_49993);
nand UO_4560 (O_4560,N_49761,N_49873);
xnor UO_4561 (O_4561,N_49781,N_49776);
or UO_4562 (O_4562,N_49793,N_49806);
nor UO_4563 (O_4563,N_49784,N_49776);
or UO_4564 (O_4564,N_49865,N_49922);
nor UO_4565 (O_4565,N_49879,N_49852);
or UO_4566 (O_4566,N_49888,N_49919);
or UO_4567 (O_4567,N_49919,N_49922);
or UO_4568 (O_4568,N_49900,N_49896);
and UO_4569 (O_4569,N_49914,N_49902);
xor UO_4570 (O_4570,N_49939,N_49978);
and UO_4571 (O_4571,N_49967,N_49854);
or UO_4572 (O_4572,N_49825,N_49835);
nand UO_4573 (O_4573,N_49964,N_49841);
nor UO_4574 (O_4574,N_49963,N_49812);
nor UO_4575 (O_4575,N_49806,N_49892);
or UO_4576 (O_4576,N_49755,N_49861);
or UO_4577 (O_4577,N_49908,N_49842);
nand UO_4578 (O_4578,N_49937,N_49854);
nor UO_4579 (O_4579,N_49791,N_49835);
or UO_4580 (O_4580,N_49950,N_49919);
nand UO_4581 (O_4581,N_49901,N_49753);
or UO_4582 (O_4582,N_49750,N_49959);
nor UO_4583 (O_4583,N_49842,N_49929);
nor UO_4584 (O_4584,N_49953,N_49798);
and UO_4585 (O_4585,N_49948,N_49786);
or UO_4586 (O_4586,N_49850,N_49804);
or UO_4587 (O_4587,N_49863,N_49790);
or UO_4588 (O_4588,N_49999,N_49948);
xnor UO_4589 (O_4589,N_49833,N_49794);
xor UO_4590 (O_4590,N_49999,N_49904);
or UO_4591 (O_4591,N_49913,N_49896);
or UO_4592 (O_4592,N_49758,N_49947);
and UO_4593 (O_4593,N_49791,N_49983);
or UO_4594 (O_4594,N_49805,N_49920);
nand UO_4595 (O_4595,N_49809,N_49791);
nand UO_4596 (O_4596,N_49887,N_49958);
xor UO_4597 (O_4597,N_49805,N_49936);
nor UO_4598 (O_4598,N_49873,N_49753);
or UO_4599 (O_4599,N_49858,N_49978);
xor UO_4600 (O_4600,N_49864,N_49972);
and UO_4601 (O_4601,N_49769,N_49913);
and UO_4602 (O_4602,N_49910,N_49789);
or UO_4603 (O_4603,N_49985,N_49790);
or UO_4604 (O_4604,N_49951,N_49991);
xor UO_4605 (O_4605,N_49972,N_49861);
or UO_4606 (O_4606,N_49975,N_49756);
xnor UO_4607 (O_4607,N_49841,N_49910);
nor UO_4608 (O_4608,N_49785,N_49957);
and UO_4609 (O_4609,N_49876,N_49765);
and UO_4610 (O_4610,N_49905,N_49977);
nand UO_4611 (O_4611,N_49845,N_49876);
xor UO_4612 (O_4612,N_49772,N_49759);
nand UO_4613 (O_4613,N_49904,N_49977);
nor UO_4614 (O_4614,N_49804,N_49802);
or UO_4615 (O_4615,N_49765,N_49916);
nand UO_4616 (O_4616,N_49884,N_49891);
nand UO_4617 (O_4617,N_49768,N_49932);
xor UO_4618 (O_4618,N_49757,N_49956);
or UO_4619 (O_4619,N_49947,N_49909);
nor UO_4620 (O_4620,N_49845,N_49912);
xor UO_4621 (O_4621,N_49901,N_49868);
nand UO_4622 (O_4622,N_49874,N_49924);
xor UO_4623 (O_4623,N_49763,N_49794);
and UO_4624 (O_4624,N_49851,N_49752);
nand UO_4625 (O_4625,N_49901,N_49999);
or UO_4626 (O_4626,N_49841,N_49847);
or UO_4627 (O_4627,N_49994,N_49776);
and UO_4628 (O_4628,N_49909,N_49985);
or UO_4629 (O_4629,N_49828,N_49834);
or UO_4630 (O_4630,N_49760,N_49938);
nand UO_4631 (O_4631,N_49993,N_49952);
and UO_4632 (O_4632,N_49905,N_49796);
nand UO_4633 (O_4633,N_49843,N_49913);
and UO_4634 (O_4634,N_49848,N_49801);
or UO_4635 (O_4635,N_49761,N_49968);
nor UO_4636 (O_4636,N_49864,N_49783);
and UO_4637 (O_4637,N_49768,N_49880);
nor UO_4638 (O_4638,N_49758,N_49980);
or UO_4639 (O_4639,N_49845,N_49952);
nor UO_4640 (O_4640,N_49802,N_49787);
nor UO_4641 (O_4641,N_49822,N_49792);
xor UO_4642 (O_4642,N_49869,N_49802);
xnor UO_4643 (O_4643,N_49949,N_49801);
nand UO_4644 (O_4644,N_49833,N_49877);
nand UO_4645 (O_4645,N_49889,N_49795);
or UO_4646 (O_4646,N_49809,N_49904);
and UO_4647 (O_4647,N_49796,N_49987);
xnor UO_4648 (O_4648,N_49780,N_49919);
nand UO_4649 (O_4649,N_49816,N_49947);
xnor UO_4650 (O_4650,N_49891,N_49856);
and UO_4651 (O_4651,N_49950,N_49923);
nor UO_4652 (O_4652,N_49826,N_49761);
xnor UO_4653 (O_4653,N_49894,N_49930);
nand UO_4654 (O_4654,N_49925,N_49957);
nor UO_4655 (O_4655,N_49773,N_49986);
nor UO_4656 (O_4656,N_49790,N_49963);
xor UO_4657 (O_4657,N_49796,N_49780);
nor UO_4658 (O_4658,N_49855,N_49929);
or UO_4659 (O_4659,N_49783,N_49947);
nand UO_4660 (O_4660,N_49953,N_49836);
nand UO_4661 (O_4661,N_49949,N_49892);
nand UO_4662 (O_4662,N_49790,N_49761);
or UO_4663 (O_4663,N_49808,N_49888);
nand UO_4664 (O_4664,N_49773,N_49984);
xor UO_4665 (O_4665,N_49939,N_49843);
nand UO_4666 (O_4666,N_49818,N_49776);
xnor UO_4667 (O_4667,N_49905,N_49768);
or UO_4668 (O_4668,N_49976,N_49904);
nand UO_4669 (O_4669,N_49884,N_49835);
xor UO_4670 (O_4670,N_49829,N_49801);
nor UO_4671 (O_4671,N_49992,N_49883);
or UO_4672 (O_4672,N_49894,N_49753);
and UO_4673 (O_4673,N_49798,N_49841);
nand UO_4674 (O_4674,N_49974,N_49979);
or UO_4675 (O_4675,N_49963,N_49873);
nor UO_4676 (O_4676,N_49968,N_49962);
xnor UO_4677 (O_4677,N_49938,N_49902);
nand UO_4678 (O_4678,N_49860,N_49782);
xor UO_4679 (O_4679,N_49862,N_49756);
xor UO_4680 (O_4680,N_49994,N_49798);
or UO_4681 (O_4681,N_49999,N_49832);
nor UO_4682 (O_4682,N_49947,N_49913);
xnor UO_4683 (O_4683,N_49919,N_49860);
or UO_4684 (O_4684,N_49757,N_49967);
or UO_4685 (O_4685,N_49847,N_49961);
and UO_4686 (O_4686,N_49960,N_49751);
and UO_4687 (O_4687,N_49857,N_49923);
nor UO_4688 (O_4688,N_49848,N_49981);
or UO_4689 (O_4689,N_49756,N_49849);
xor UO_4690 (O_4690,N_49996,N_49822);
nand UO_4691 (O_4691,N_49955,N_49851);
or UO_4692 (O_4692,N_49750,N_49920);
xnor UO_4693 (O_4693,N_49945,N_49775);
xnor UO_4694 (O_4694,N_49904,N_49890);
xnor UO_4695 (O_4695,N_49844,N_49805);
nand UO_4696 (O_4696,N_49921,N_49814);
nand UO_4697 (O_4697,N_49762,N_49992);
nor UO_4698 (O_4698,N_49946,N_49915);
nand UO_4699 (O_4699,N_49892,N_49891);
or UO_4700 (O_4700,N_49870,N_49985);
nor UO_4701 (O_4701,N_49877,N_49996);
nor UO_4702 (O_4702,N_49804,N_49839);
and UO_4703 (O_4703,N_49971,N_49887);
xor UO_4704 (O_4704,N_49757,N_49896);
nand UO_4705 (O_4705,N_49920,N_49822);
and UO_4706 (O_4706,N_49791,N_49815);
and UO_4707 (O_4707,N_49970,N_49972);
xor UO_4708 (O_4708,N_49924,N_49964);
or UO_4709 (O_4709,N_49911,N_49867);
xnor UO_4710 (O_4710,N_49966,N_49916);
nand UO_4711 (O_4711,N_49750,N_49976);
and UO_4712 (O_4712,N_49998,N_49936);
xnor UO_4713 (O_4713,N_49826,N_49999);
or UO_4714 (O_4714,N_49928,N_49799);
or UO_4715 (O_4715,N_49881,N_49962);
nand UO_4716 (O_4716,N_49856,N_49996);
and UO_4717 (O_4717,N_49765,N_49999);
nor UO_4718 (O_4718,N_49858,N_49906);
or UO_4719 (O_4719,N_49787,N_49779);
and UO_4720 (O_4720,N_49833,N_49820);
nand UO_4721 (O_4721,N_49803,N_49900);
nor UO_4722 (O_4722,N_49917,N_49923);
and UO_4723 (O_4723,N_49847,N_49928);
or UO_4724 (O_4724,N_49862,N_49780);
nand UO_4725 (O_4725,N_49840,N_49974);
and UO_4726 (O_4726,N_49808,N_49950);
and UO_4727 (O_4727,N_49940,N_49825);
and UO_4728 (O_4728,N_49811,N_49889);
or UO_4729 (O_4729,N_49792,N_49783);
or UO_4730 (O_4730,N_49813,N_49976);
or UO_4731 (O_4731,N_49949,N_49980);
and UO_4732 (O_4732,N_49752,N_49778);
nor UO_4733 (O_4733,N_49973,N_49936);
and UO_4734 (O_4734,N_49983,N_49879);
nand UO_4735 (O_4735,N_49898,N_49982);
xnor UO_4736 (O_4736,N_49761,N_49825);
nor UO_4737 (O_4737,N_49838,N_49941);
nor UO_4738 (O_4738,N_49963,N_49781);
xor UO_4739 (O_4739,N_49899,N_49901);
nand UO_4740 (O_4740,N_49757,N_49842);
or UO_4741 (O_4741,N_49965,N_49846);
xor UO_4742 (O_4742,N_49827,N_49963);
xnor UO_4743 (O_4743,N_49871,N_49850);
or UO_4744 (O_4744,N_49910,N_49904);
nand UO_4745 (O_4745,N_49864,N_49966);
or UO_4746 (O_4746,N_49920,N_49760);
and UO_4747 (O_4747,N_49835,N_49851);
nand UO_4748 (O_4748,N_49792,N_49887);
nor UO_4749 (O_4749,N_49905,N_49845);
nand UO_4750 (O_4750,N_49856,N_49926);
nand UO_4751 (O_4751,N_49822,N_49889);
nand UO_4752 (O_4752,N_49932,N_49939);
nand UO_4753 (O_4753,N_49945,N_49755);
or UO_4754 (O_4754,N_49945,N_49978);
xnor UO_4755 (O_4755,N_49982,N_49849);
and UO_4756 (O_4756,N_49956,N_49866);
nand UO_4757 (O_4757,N_49920,N_49839);
nor UO_4758 (O_4758,N_49946,N_49982);
and UO_4759 (O_4759,N_49850,N_49794);
and UO_4760 (O_4760,N_49946,N_49876);
or UO_4761 (O_4761,N_49850,N_49802);
xor UO_4762 (O_4762,N_49931,N_49763);
nand UO_4763 (O_4763,N_49848,N_49977);
or UO_4764 (O_4764,N_49960,N_49805);
or UO_4765 (O_4765,N_49913,N_49779);
nor UO_4766 (O_4766,N_49999,N_49862);
nand UO_4767 (O_4767,N_49923,N_49940);
xor UO_4768 (O_4768,N_49856,N_49902);
nand UO_4769 (O_4769,N_49759,N_49831);
or UO_4770 (O_4770,N_49781,N_49961);
xor UO_4771 (O_4771,N_49948,N_49780);
nor UO_4772 (O_4772,N_49993,N_49777);
nand UO_4773 (O_4773,N_49909,N_49922);
or UO_4774 (O_4774,N_49880,N_49773);
nand UO_4775 (O_4775,N_49921,N_49912);
nand UO_4776 (O_4776,N_49775,N_49804);
nor UO_4777 (O_4777,N_49974,N_49931);
nor UO_4778 (O_4778,N_49771,N_49986);
or UO_4779 (O_4779,N_49806,N_49853);
or UO_4780 (O_4780,N_49915,N_49794);
xor UO_4781 (O_4781,N_49920,N_49982);
and UO_4782 (O_4782,N_49750,N_49856);
nor UO_4783 (O_4783,N_49866,N_49791);
nand UO_4784 (O_4784,N_49981,N_49864);
nand UO_4785 (O_4785,N_49994,N_49803);
or UO_4786 (O_4786,N_49808,N_49969);
and UO_4787 (O_4787,N_49825,N_49970);
or UO_4788 (O_4788,N_49969,N_49765);
xnor UO_4789 (O_4789,N_49887,N_49924);
nor UO_4790 (O_4790,N_49844,N_49808);
or UO_4791 (O_4791,N_49787,N_49874);
nand UO_4792 (O_4792,N_49895,N_49817);
nor UO_4793 (O_4793,N_49767,N_49903);
and UO_4794 (O_4794,N_49881,N_49983);
xnor UO_4795 (O_4795,N_49936,N_49914);
or UO_4796 (O_4796,N_49989,N_49937);
nand UO_4797 (O_4797,N_49762,N_49985);
or UO_4798 (O_4798,N_49920,N_49965);
nand UO_4799 (O_4799,N_49960,N_49775);
nor UO_4800 (O_4800,N_49819,N_49959);
and UO_4801 (O_4801,N_49900,N_49841);
nor UO_4802 (O_4802,N_49768,N_49917);
nor UO_4803 (O_4803,N_49808,N_49801);
nor UO_4804 (O_4804,N_49940,N_49914);
and UO_4805 (O_4805,N_49995,N_49956);
and UO_4806 (O_4806,N_49933,N_49761);
nand UO_4807 (O_4807,N_49916,N_49950);
nor UO_4808 (O_4808,N_49995,N_49843);
xor UO_4809 (O_4809,N_49819,N_49810);
nor UO_4810 (O_4810,N_49978,N_49796);
xnor UO_4811 (O_4811,N_49952,N_49937);
and UO_4812 (O_4812,N_49754,N_49792);
or UO_4813 (O_4813,N_49763,N_49816);
nor UO_4814 (O_4814,N_49962,N_49833);
or UO_4815 (O_4815,N_49774,N_49999);
and UO_4816 (O_4816,N_49832,N_49849);
nor UO_4817 (O_4817,N_49793,N_49974);
nand UO_4818 (O_4818,N_49801,N_49950);
xor UO_4819 (O_4819,N_49954,N_49861);
or UO_4820 (O_4820,N_49855,N_49968);
and UO_4821 (O_4821,N_49895,N_49880);
nand UO_4822 (O_4822,N_49857,N_49772);
or UO_4823 (O_4823,N_49812,N_49908);
nand UO_4824 (O_4824,N_49932,N_49960);
nor UO_4825 (O_4825,N_49787,N_49929);
and UO_4826 (O_4826,N_49875,N_49948);
or UO_4827 (O_4827,N_49812,N_49784);
and UO_4828 (O_4828,N_49883,N_49926);
xor UO_4829 (O_4829,N_49989,N_49789);
or UO_4830 (O_4830,N_49924,N_49873);
and UO_4831 (O_4831,N_49973,N_49822);
or UO_4832 (O_4832,N_49790,N_49976);
and UO_4833 (O_4833,N_49980,N_49935);
nand UO_4834 (O_4834,N_49841,N_49842);
and UO_4835 (O_4835,N_49828,N_49981);
nand UO_4836 (O_4836,N_49812,N_49976);
xor UO_4837 (O_4837,N_49947,N_49752);
xnor UO_4838 (O_4838,N_49903,N_49820);
nand UO_4839 (O_4839,N_49818,N_49909);
and UO_4840 (O_4840,N_49984,N_49846);
and UO_4841 (O_4841,N_49868,N_49770);
nand UO_4842 (O_4842,N_49857,N_49984);
or UO_4843 (O_4843,N_49915,N_49925);
xor UO_4844 (O_4844,N_49932,N_49945);
nor UO_4845 (O_4845,N_49826,N_49898);
xor UO_4846 (O_4846,N_49891,N_49913);
and UO_4847 (O_4847,N_49944,N_49980);
xor UO_4848 (O_4848,N_49833,N_49830);
nand UO_4849 (O_4849,N_49989,N_49757);
and UO_4850 (O_4850,N_49813,N_49867);
nand UO_4851 (O_4851,N_49809,N_49926);
nor UO_4852 (O_4852,N_49970,N_49933);
or UO_4853 (O_4853,N_49942,N_49987);
nor UO_4854 (O_4854,N_49802,N_49975);
nor UO_4855 (O_4855,N_49895,N_49951);
nand UO_4856 (O_4856,N_49853,N_49917);
or UO_4857 (O_4857,N_49801,N_49980);
nand UO_4858 (O_4858,N_49991,N_49832);
xor UO_4859 (O_4859,N_49940,N_49902);
or UO_4860 (O_4860,N_49994,N_49923);
and UO_4861 (O_4861,N_49930,N_49872);
and UO_4862 (O_4862,N_49910,N_49915);
nor UO_4863 (O_4863,N_49901,N_49837);
or UO_4864 (O_4864,N_49879,N_49867);
or UO_4865 (O_4865,N_49997,N_49914);
nand UO_4866 (O_4866,N_49769,N_49794);
or UO_4867 (O_4867,N_49793,N_49915);
or UO_4868 (O_4868,N_49892,N_49794);
nor UO_4869 (O_4869,N_49816,N_49998);
nor UO_4870 (O_4870,N_49898,N_49835);
nand UO_4871 (O_4871,N_49865,N_49859);
or UO_4872 (O_4872,N_49916,N_49866);
nor UO_4873 (O_4873,N_49889,N_49919);
and UO_4874 (O_4874,N_49869,N_49832);
or UO_4875 (O_4875,N_49817,N_49775);
and UO_4876 (O_4876,N_49769,N_49796);
or UO_4877 (O_4877,N_49834,N_49869);
xor UO_4878 (O_4878,N_49807,N_49810);
xor UO_4879 (O_4879,N_49827,N_49976);
nor UO_4880 (O_4880,N_49893,N_49821);
or UO_4881 (O_4881,N_49954,N_49781);
or UO_4882 (O_4882,N_49950,N_49924);
nand UO_4883 (O_4883,N_49839,N_49809);
or UO_4884 (O_4884,N_49990,N_49944);
nor UO_4885 (O_4885,N_49780,N_49790);
nand UO_4886 (O_4886,N_49856,N_49819);
nor UO_4887 (O_4887,N_49844,N_49894);
nand UO_4888 (O_4888,N_49854,N_49886);
nor UO_4889 (O_4889,N_49878,N_49992);
or UO_4890 (O_4890,N_49787,N_49888);
xor UO_4891 (O_4891,N_49930,N_49819);
xnor UO_4892 (O_4892,N_49781,N_49904);
nor UO_4893 (O_4893,N_49863,N_49820);
xnor UO_4894 (O_4894,N_49943,N_49923);
and UO_4895 (O_4895,N_49880,N_49815);
or UO_4896 (O_4896,N_49861,N_49910);
xnor UO_4897 (O_4897,N_49935,N_49810);
and UO_4898 (O_4898,N_49862,N_49924);
and UO_4899 (O_4899,N_49764,N_49818);
nor UO_4900 (O_4900,N_49940,N_49802);
nor UO_4901 (O_4901,N_49781,N_49836);
xnor UO_4902 (O_4902,N_49814,N_49854);
nand UO_4903 (O_4903,N_49981,N_49891);
and UO_4904 (O_4904,N_49841,N_49768);
and UO_4905 (O_4905,N_49791,N_49788);
or UO_4906 (O_4906,N_49919,N_49955);
nand UO_4907 (O_4907,N_49883,N_49901);
or UO_4908 (O_4908,N_49847,N_49796);
nor UO_4909 (O_4909,N_49881,N_49834);
or UO_4910 (O_4910,N_49850,N_49793);
nand UO_4911 (O_4911,N_49774,N_49856);
or UO_4912 (O_4912,N_49751,N_49990);
nand UO_4913 (O_4913,N_49773,N_49810);
nand UO_4914 (O_4914,N_49756,N_49842);
nor UO_4915 (O_4915,N_49970,N_49952);
xor UO_4916 (O_4916,N_49971,N_49755);
nor UO_4917 (O_4917,N_49892,N_49973);
xnor UO_4918 (O_4918,N_49834,N_49804);
xor UO_4919 (O_4919,N_49999,N_49921);
or UO_4920 (O_4920,N_49925,N_49854);
nor UO_4921 (O_4921,N_49992,N_49769);
or UO_4922 (O_4922,N_49791,N_49869);
nand UO_4923 (O_4923,N_49803,N_49986);
nor UO_4924 (O_4924,N_49882,N_49950);
nor UO_4925 (O_4925,N_49800,N_49833);
or UO_4926 (O_4926,N_49949,N_49808);
or UO_4927 (O_4927,N_49911,N_49837);
nor UO_4928 (O_4928,N_49880,N_49920);
nor UO_4929 (O_4929,N_49823,N_49817);
and UO_4930 (O_4930,N_49901,N_49816);
nor UO_4931 (O_4931,N_49766,N_49982);
nand UO_4932 (O_4932,N_49987,N_49861);
xnor UO_4933 (O_4933,N_49806,N_49883);
and UO_4934 (O_4934,N_49936,N_49841);
nand UO_4935 (O_4935,N_49893,N_49926);
nor UO_4936 (O_4936,N_49872,N_49833);
nor UO_4937 (O_4937,N_49826,N_49957);
or UO_4938 (O_4938,N_49925,N_49778);
xor UO_4939 (O_4939,N_49998,N_49961);
or UO_4940 (O_4940,N_49938,N_49897);
and UO_4941 (O_4941,N_49839,N_49969);
and UO_4942 (O_4942,N_49898,N_49944);
nand UO_4943 (O_4943,N_49825,N_49808);
nor UO_4944 (O_4944,N_49750,N_49878);
or UO_4945 (O_4945,N_49796,N_49866);
nand UO_4946 (O_4946,N_49994,N_49847);
nand UO_4947 (O_4947,N_49787,N_49780);
nand UO_4948 (O_4948,N_49991,N_49750);
nand UO_4949 (O_4949,N_49913,N_49792);
or UO_4950 (O_4950,N_49829,N_49755);
nor UO_4951 (O_4951,N_49897,N_49893);
xor UO_4952 (O_4952,N_49811,N_49916);
and UO_4953 (O_4953,N_49837,N_49824);
or UO_4954 (O_4954,N_49854,N_49852);
and UO_4955 (O_4955,N_49892,N_49761);
or UO_4956 (O_4956,N_49858,N_49888);
or UO_4957 (O_4957,N_49963,N_49967);
xor UO_4958 (O_4958,N_49869,N_49774);
nand UO_4959 (O_4959,N_49976,N_49942);
nand UO_4960 (O_4960,N_49881,N_49797);
or UO_4961 (O_4961,N_49805,N_49998);
nor UO_4962 (O_4962,N_49779,N_49796);
xnor UO_4963 (O_4963,N_49933,N_49800);
nor UO_4964 (O_4964,N_49902,N_49842);
xor UO_4965 (O_4965,N_49975,N_49807);
or UO_4966 (O_4966,N_49758,N_49853);
nand UO_4967 (O_4967,N_49847,N_49867);
nor UO_4968 (O_4968,N_49828,N_49784);
nor UO_4969 (O_4969,N_49936,N_49984);
or UO_4970 (O_4970,N_49939,N_49769);
xnor UO_4971 (O_4971,N_49966,N_49897);
xnor UO_4972 (O_4972,N_49906,N_49851);
nor UO_4973 (O_4973,N_49770,N_49986);
and UO_4974 (O_4974,N_49960,N_49766);
and UO_4975 (O_4975,N_49754,N_49852);
or UO_4976 (O_4976,N_49902,N_49826);
nand UO_4977 (O_4977,N_49907,N_49869);
xor UO_4978 (O_4978,N_49940,N_49846);
xor UO_4979 (O_4979,N_49882,N_49910);
nor UO_4980 (O_4980,N_49886,N_49899);
nand UO_4981 (O_4981,N_49925,N_49913);
and UO_4982 (O_4982,N_49775,N_49810);
or UO_4983 (O_4983,N_49994,N_49922);
xnor UO_4984 (O_4984,N_49763,N_49882);
and UO_4985 (O_4985,N_49881,N_49926);
and UO_4986 (O_4986,N_49992,N_49971);
nor UO_4987 (O_4987,N_49890,N_49801);
and UO_4988 (O_4988,N_49787,N_49885);
xnor UO_4989 (O_4989,N_49887,N_49804);
and UO_4990 (O_4990,N_49760,N_49981);
xor UO_4991 (O_4991,N_49954,N_49994);
xor UO_4992 (O_4992,N_49936,N_49756);
or UO_4993 (O_4993,N_49868,N_49800);
or UO_4994 (O_4994,N_49901,N_49774);
nand UO_4995 (O_4995,N_49987,N_49845);
nor UO_4996 (O_4996,N_49896,N_49986);
and UO_4997 (O_4997,N_49964,N_49970);
nor UO_4998 (O_4998,N_49753,N_49933);
or UO_4999 (O_4999,N_49777,N_49768);
endmodule