module basic_1500_15000_2000_3_levels_10xor_3(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10012,N_10013,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10030,N_10031,N_10032,N_10034,N_10035,N_10036,N_10037,N_10038,N_10040,N_10041,N_10042,N_10043,N_10045,N_10046,N_10047,N_10049,N_10050,N_10051,N_10052,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10070,N_10076,N_10077,N_10078,N_10079,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10093,N_10095,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10105,N_10106,N_10107,N_10108,N_10110,N_10111,N_10112,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10137,N_10138,N_10140,N_10144,N_10145,N_10146,N_10148,N_10149,N_10150,N_10151,N_10154,N_10155,N_10156,N_10157,N_10159,N_10160,N_10161,N_10163,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10180,N_10181,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10193,N_10194,N_10195,N_10196,N_10197,N_10199,N_10201,N_10202,N_10203,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10234,N_10235,N_10236,N_10238,N_10240,N_10241,N_10242,N_10244,N_10245,N_10247,N_10248,N_10249,N_10250,N_10251,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10281,N_10282,N_10284,N_10285,N_10286,N_10287,N_10288,N_10290,N_10291,N_10293,N_10294,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10304,N_10305,N_10306,N_10307,N_10309,N_10310,N_10311,N_10313,N_10316,N_10317,N_10318,N_10319,N_10320,N_10322,N_10323,N_10324,N_10325,N_10326,N_10328,N_10329,N_10330,N_10332,N_10333,N_10334,N_10337,N_10338,N_10339,N_10340,N_10342,N_10344,N_10345,N_10347,N_10348,N_10349,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10376,N_10377,N_10378,N_10379,N_10381,N_10384,N_10388,N_10389,N_10390,N_10391,N_10392,N_10394,N_10395,N_10396,N_10397,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10410,N_10411,N_10412,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10429,N_10431,N_10432,N_10433,N_10434,N_10435,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10462,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10483,N_10484,N_10486,N_10488,N_10489,N_10490,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10508,N_10509,N_10510,N_10511,N_10512,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10523,N_10524,N_10526,N_10527,N_10528,N_10529,N_10530,N_10533,N_10534,N_10535,N_10536,N_10538,N_10540,N_10541,N_10542,N_10543,N_10544,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10557,N_10558,N_10560,N_10563,N_10564,N_10565,N_10567,N_10568,N_10569,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10580,N_10581,N_10582,N_10583,N_10584,N_10587,N_10588,N_10589,N_10591,N_10592,N_10593,N_10594,N_10596,N_10598,N_10599,N_10601,N_10603,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10617,N_10618,N_10619,N_10620,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10633,N_10634,N_10635,N_10636,N_10637,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10668,N_10669,N_10670,N_10672,N_10674,N_10675,N_10676,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10685,N_10687,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10698,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10723,N_10724,N_10725,N_10726,N_10727,N_10729,N_10730,N_10732,N_10734,N_10735,N_10736,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10761,N_10762,N_10763,N_10764,N_10765,N_10768,N_10769,N_10770,N_10771,N_10772,N_10775,N_10776,N_10777,N_10778,N_10779,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10793,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10835,N_10836,N_10837,N_10838,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10853,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10871,N_10872,N_10873,N_10874,N_10876,N_10877,N_10878,N_10882,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10891,N_10892,N_10893,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10930,N_10931,N_10932,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10954,N_10955,N_10957,N_10958,N_10960,N_10961,N_10962,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10986,N_10987,N_10989,N_10990,N_10991,N_10992,N_10993,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11026,N_11027,N_11028,N_11029,N_11031,N_11032,N_11033,N_11035,N_11036,N_11037,N_11038,N_11039,N_11041,N_11042,N_11043,N_11044,N_11045,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11075,N_11077,N_11078,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11088,N_11089,N_11091,N_11093,N_11094,N_11095,N_11097,N_11098,N_11099,N_11101,N_11102,N_11104,N_11105,N_11106,N_11107,N_11108,N_11110,N_11111,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11132,N_11133,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11145,N_11146,N_11147,N_11151,N_11152,N_11153,N_11154,N_11155,N_11157,N_11158,N_11159,N_11160,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11173,N_11174,N_11176,N_11178,N_11179,N_11180,N_11181,N_11182,N_11187,N_11189,N_11190,N_11191,N_11193,N_11194,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11211,N_11213,N_11214,N_11215,N_11217,N_11218,N_11219,N_11220,N_11222,N_11223,N_11224,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11233,N_11234,N_11235,N_11236,N_11238,N_11239,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11272,N_11273,N_11274,N_11276,N_11277,N_11278,N_11279,N_11280,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11295,N_11296,N_11297,N_11299,N_11300,N_11302,N_11303,N_11306,N_11307,N_11308,N_11309,N_11310,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11341,N_11343,N_11344,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11353,N_11355,N_11357,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11376,N_11378,N_11379,N_11381,N_11382,N_11383,N_11386,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11397,N_11398,N_11403,N_11404,N_11405,N_11407,N_11408,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11420,N_11422,N_11423,N_11424,N_11427,N_11428,N_11429,N_11430,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11444,N_11445,N_11446,N_11447,N_11449,N_11450,N_11451,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11471,N_11473,N_11475,N_11476,N_11477,N_11479,N_11480,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11493,N_11494,N_11495,N_11496,N_11503,N_11504,N_11506,N_11507,N_11509,N_11510,N_11511,N_11512,N_11514,N_11515,N_11517,N_11519,N_11521,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11534,N_11535,N_11537,N_11538,N_11539,N_11541,N_11542,N_11543,N_11544,N_11546,N_11547,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11571,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11593,N_11594,N_11595,N_11596,N_11599,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11613,N_11614,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11627,N_11628,N_11629,N_11631,N_11632,N_11633,N_11634,N_11635,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11652,N_11653,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11677,N_11679,N_11680,N_11682,N_11683,N_11684,N_11685,N_11686,N_11688,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11698,N_11699,N_11701,N_11702,N_11703,N_11704,N_11707,N_11708,N_11709,N_11710,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11721,N_11722,N_11723,N_11724,N_11727,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11743,N_11744,N_11745,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11767,N_11768,N_11769,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11784,N_11785,N_11786,N_11787,N_11788,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11806,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11820,N_11822,N_11823,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11841,N_11842,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11852,N_11853,N_11854,N_11856,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11888,N_11889,N_11890,N_11891,N_11892,N_11894,N_11896,N_11898,N_11899,N_11900,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11915,N_11916,N_11917,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11939,N_11940,N_11942,N_11943,N_11944,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11954,N_11955,N_11957,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11969,N_11970,N_11971,N_11972,N_11973,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12010,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12019,N_12021,N_12022,N_12023,N_12024,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12039,N_12040,N_12041,N_12044,N_12045,N_12046,N_12047,N_12049,N_12052,N_12053,N_12054,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12066,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12079,N_12082,N_12083,N_12084,N_12085,N_12086,N_12088,N_12089,N_12090,N_12091,N_12093,N_12094,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12105,N_12106,N_12107,N_12109,N_12110,N_12112,N_12113,N_12114,N_12115,N_12116,N_12118,N_12119,N_12120,N_12121,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12139,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12153,N_12154,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12185,N_12186,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12212,N_12213,N_12214,N_12215,N_12216,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12227,N_12228,N_12230,N_12231,N_12232,N_12233,N_12235,N_12236,N_12237,N_12239,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12250,N_12251,N_12252,N_12253,N_12254,N_12257,N_12258,N_12259,N_12260,N_12262,N_12263,N_12264,N_12266,N_12267,N_12268,N_12269,N_12271,N_12274,N_12275,N_12276,N_12277,N_12278,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12362,N_12363,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12372,N_12373,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12388,N_12389,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12399,N_12400,N_12401,N_12403,N_12405,N_12406,N_12407,N_12408,N_12409,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12426,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12439,N_12441,N_12443,N_12445,N_12446,N_12447,N_12449,N_12450,N_12451,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12473,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12485,N_12486,N_12487,N_12489,N_12490,N_12491,N_12492,N_12493,N_12495,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12504,N_12506,N_12508,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12524,N_12525,N_12526,N_12527,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12573,N_12575,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12584,N_12585,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12604,N_12605,N_12607,N_12609,N_12610,N_12612,N_12613,N_12614,N_12616,N_12618,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12639,N_12642,N_12643,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12666,N_12667,N_12668,N_12669,N_12670,N_12672,N_12673,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12697,N_12700,N_12701,N_12702,N_12704,N_12705,N_12706,N_12707,N_12708,N_12710,N_12711,N_12712,N_12714,N_12715,N_12716,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12734,N_12735,N_12737,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12755,N_12756,N_12758,N_12759,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12774,N_12777,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12795,N_12798,N_12799,N_12802,N_12803,N_12804,N_12805,N_12807,N_12808,N_12810,N_12811,N_12812,N_12813,N_12814,N_12816,N_12817,N_12818,N_12819,N_12821,N_12823,N_12824,N_12825,N_12826,N_12828,N_12829,N_12830,N_12831,N_12833,N_12834,N_12835,N_12836,N_12838,N_12840,N_12842,N_12843,N_12844,N_12846,N_12849,N_12850,N_12851,N_12853,N_12858,N_12859,N_12860,N_12861,N_12862,N_12865,N_12866,N_12867,N_12868,N_12869,N_12871,N_12872,N_12874,N_12877,N_12878,N_12879,N_12881,N_12882,N_12883,N_12884,N_12885,N_12887,N_12890,N_12892,N_12893,N_12897,N_12899,N_12900,N_12901,N_12902,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12913,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12924,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12935,N_12936,N_12937,N_12939,N_12940,N_12941,N_12943,N_12945,N_12946,N_12947,N_12948,N_12949,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12968,N_12969,N_12970,N_12971,N_12974,N_12975,N_12976,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13006,N_13007,N_13010,N_13012,N_13013,N_13014,N_13015,N_13017,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13038,N_13039,N_13040,N_13041,N_13043,N_13045,N_13048,N_13049,N_13054,N_13055,N_13056,N_13058,N_13060,N_13061,N_13062,N_13063,N_13065,N_13066,N_13067,N_13070,N_13071,N_13073,N_13075,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13085,N_13087,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13110,N_13111,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13148,N_13149,N_13150,N_13152,N_13153,N_13154,N_13155,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13176,N_13178,N_13179,N_13181,N_13182,N_13184,N_13185,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13209,N_13210,N_13211,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13223,N_13225,N_13226,N_13227,N_13228,N_13230,N_13231,N_13234,N_13235,N_13236,N_13237,N_13238,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13249,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13330,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13357,N_13358,N_13360,N_13361,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13379,N_13380,N_13381,N_13382,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13400,N_13401,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13418,N_13419,N_13420,N_13421,N_13422,N_13424,N_13425,N_13426,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13435,N_13436,N_13437,N_13438,N_13439,N_13443,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13458,N_13459,N_13460,N_13461,N_13463,N_13464,N_13465,N_13466,N_13468,N_13469,N_13470,N_13471,N_13472,N_13474,N_13475,N_13476,N_13478,N_13479,N_13480,N_13481,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13517,N_13518,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13531,N_13533,N_13534,N_13535,N_13536,N_13537,N_13539,N_13540,N_13542,N_13543,N_13544,N_13545,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13557,N_13558,N_13559,N_13560,N_13561,N_13563,N_13564,N_13567,N_13569,N_13570,N_13571,N_13573,N_13575,N_13576,N_13579,N_13580,N_13581,N_13582,N_13584,N_13586,N_13587,N_13588,N_13589,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13601,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13632,N_13633,N_13634,N_13635,N_13637,N_13638,N_13639,N_13640,N_13641,N_13644,N_13645,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13668,N_13669,N_13670,N_13671,N_13672,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13683,N_13684,N_13685,N_13686,N_13687,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13699,N_13701,N_13704,N_13705,N_13708,N_13709,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13730,N_13731,N_13732,N_13736,N_13739,N_13740,N_13741,N_13743,N_13744,N_13745,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13767,N_13768,N_13770,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13806,N_13808,N_13809,N_13811,N_13812,N_13813,N_13815,N_13816,N_13817,N_13819,N_13820,N_13821,N_13822,N_13823,N_13825,N_13826,N_13827,N_13828,N_13831,N_13832,N_13834,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13863,N_13864,N_13865,N_13867,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13904,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13915,N_13916,N_13917,N_13918,N_13919,N_13921,N_13922,N_13923,N_13924,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13938,N_13939,N_13940,N_13941,N_13943,N_13944,N_13945,N_13947,N_13948,N_13949,N_13950,N_13951,N_13953,N_13954,N_13955,N_13956,N_13957,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13983,N_13984,N_13985,N_13986,N_13988,N_13989,N_13991,N_13992,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14018,N_14020,N_14021,N_14022,N_14024,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14038,N_14039,N_14040,N_14042,N_14043,N_14045,N_14046,N_14047,N_14048,N_14049,N_14051,N_14054,N_14056,N_14057,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14070,N_14071,N_14072,N_14074,N_14075,N_14076,N_14077,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14099,N_14100,N_14101,N_14103,N_14104,N_14105,N_14106,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14120,N_14121,N_14122,N_14123,N_14124,N_14126,N_14127,N_14129,N_14130,N_14131,N_14132,N_14133,N_14135,N_14136,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14145,N_14146,N_14147,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14160,N_14161,N_14162,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14195,N_14198,N_14199,N_14200,N_14201,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14213,N_14215,N_14216,N_14217,N_14218,N_14219,N_14221,N_14222,N_14225,N_14226,N_14227,N_14228,N_14230,N_14232,N_14233,N_14234,N_14235,N_14236,N_14238,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14264,N_14265,N_14266,N_14267,N_14268,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14284,N_14286,N_14287,N_14288,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14309,N_14311,N_14312,N_14313,N_14314,N_14316,N_14317,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14330,N_14331,N_14332,N_14333,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14351,N_14352,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14367,N_14368,N_14370,N_14371,N_14372,N_14373,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14395,N_14396,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14407,N_14409,N_14410,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14422,N_14424,N_14425,N_14426,N_14427,N_14429,N_14431,N_14432,N_14433,N_14435,N_14438,N_14440,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14459,N_14460,N_14464,N_14465,N_14467,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14485,N_14486,N_14487,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14497,N_14498,N_14499,N_14500,N_14501,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14516,N_14518,N_14519,N_14520,N_14523,N_14525,N_14527,N_14528,N_14530,N_14531,N_14532,N_14533,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14582,N_14583,N_14584,N_14585,N_14587,N_14588,N_14589,N_14590,N_14591,N_14594,N_14595,N_14596,N_14597,N_14598,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14618,N_14619,N_14620,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14634,N_14635,N_14636,N_14638,N_14639,N_14640,N_14642,N_14643,N_14646,N_14648,N_14649,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14661,N_14663,N_14664,N_14665,N_14666,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14690,N_14691,N_14694,N_14695,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14708,N_14709,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14746,N_14747,N_14748,N_14751,N_14753,N_14754,N_14755,N_14759,N_14760,N_14761,N_14762,N_14764,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14778,N_14779,N_14780,N_14782,N_14783,N_14784,N_14785,N_14786,N_14788,N_14789,N_14790,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14804,N_14805,N_14807,N_14808,N_14811,N_14812,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14860,N_14861,N_14863,N_14864,N_14865,N_14866,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14877,N_14879,N_14880,N_14881,N_14882,N_14884,N_14885,N_14886,N_14889,N_14890,N_14891,N_14892,N_14894,N_14895,N_14896,N_14897,N_14898,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14908,N_14910,N_14911,N_14912,N_14915,N_14917,N_14918,N_14920,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14931,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14948,N_14949,N_14955,N_14956,N_14958,N_14960,N_14962,N_14963,N_14965,N_14966,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14985,N_14986,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14995,N_14996,N_14997,N_14998,N_14999;
nor U0 (N_0,In_1029,In_933);
nand U1 (N_1,In_1133,In_532);
and U2 (N_2,In_1083,In_574);
xor U3 (N_3,In_937,In_18);
xnor U4 (N_4,In_122,In_1086);
xor U5 (N_5,In_1400,In_768);
nor U6 (N_6,In_1257,In_877);
and U7 (N_7,In_582,In_668);
and U8 (N_8,In_921,In_647);
nor U9 (N_9,In_896,In_539);
and U10 (N_10,In_562,In_792);
xor U11 (N_11,In_607,In_22);
nor U12 (N_12,In_451,In_1119);
nor U13 (N_13,In_1420,In_375);
or U14 (N_14,In_34,In_711);
or U15 (N_15,In_1055,In_1235);
xnor U16 (N_16,In_153,In_518);
and U17 (N_17,In_300,In_371);
xnor U18 (N_18,In_643,In_84);
xor U19 (N_19,In_201,In_1042);
and U20 (N_20,In_411,In_435);
or U21 (N_21,In_1246,In_5);
nor U22 (N_22,In_839,In_906);
or U23 (N_23,In_732,In_360);
xnor U24 (N_24,In_97,In_1025);
nor U25 (N_25,In_853,In_769);
nor U26 (N_26,In_525,In_900);
xnor U27 (N_27,In_1310,In_616);
or U28 (N_28,In_347,In_0);
and U29 (N_29,In_1388,In_764);
nor U30 (N_30,In_1241,In_850);
xor U31 (N_31,In_7,In_954);
or U32 (N_32,In_901,In_237);
xnor U33 (N_33,In_962,In_425);
xor U34 (N_34,In_366,In_265);
nand U35 (N_35,In_756,In_317);
nor U36 (N_36,In_899,In_698);
nor U37 (N_37,In_581,In_880);
nor U38 (N_38,In_571,In_564);
or U39 (N_39,In_830,In_71);
or U40 (N_40,In_1239,In_489);
xor U41 (N_41,In_154,In_87);
or U42 (N_42,In_1339,In_444);
or U43 (N_43,In_148,In_1250);
xor U44 (N_44,In_775,In_1305);
and U45 (N_45,In_1410,In_1084);
or U46 (N_46,In_1456,In_1249);
or U47 (N_47,In_1403,In_1460);
and U48 (N_48,In_939,In_433);
and U49 (N_49,In_1152,In_251);
and U50 (N_50,In_348,In_398);
xor U51 (N_51,In_471,In_117);
nand U52 (N_52,In_1346,In_859);
xor U53 (N_53,In_608,In_1028);
nand U54 (N_54,In_1040,In_553);
and U55 (N_55,In_514,In_1099);
nor U56 (N_56,In_78,In_273);
or U57 (N_57,In_1402,In_697);
nor U58 (N_58,In_1004,In_187);
nor U59 (N_59,In_79,In_150);
or U60 (N_60,In_579,In_660);
nand U61 (N_61,In_865,In_794);
or U62 (N_62,In_816,In_1205);
nand U63 (N_63,In_889,In_29);
and U64 (N_64,In_909,In_973);
nor U65 (N_65,In_980,In_1491);
xor U66 (N_66,In_531,In_842);
and U67 (N_67,In_1343,In_924);
xor U68 (N_68,In_923,In_207);
nor U69 (N_69,In_1315,In_17);
nor U70 (N_70,In_1313,In_1077);
or U71 (N_71,In_715,In_1110);
nand U72 (N_72,In_202,In_881);
nand U73 (N_73,In_191,In_767);
and U74 (N_74,In_524,In_641);
nand U75 (N_75,In_548,In_1476);
or U76 (N_76,In_964,In_86);
nand U77 (N_77,In_740,In_1264);
and U78 (N_78,In_834,In_1211);
nor U79 (N_79,In_892,In_1244);
nor U80 (N_80,In_1461,In_802);
and U81 (N_81,In_1416,In_384);
xnor U82 (N_82,In_165,In_984);
nor U83 (N_83,In_1181,In_640);
xor U84 (N_84,In_1306,In_103);
nand U85 (N_85,In_1340,In_426);
and U86 (N_86,In_1018,In_227);
or U87 (N_87,In_389,In_1115);
nor U88 (N_88,In_837,In_1465);
or U89 (N_89,In_1330,In_293);
nand U90 (N_90,In_599,In_602);
nand U91 (N_91,In_1143,In_350);
nand U92 (N_92,In_1300,In_573);
nand U93 (N_93,In_415,In_1356);
or U94 (N_94,In_314,In_345);
nor U95 (N_95,In_1467,In_864);
nand U96 (N_96,In_594,In_898);
or U97 (N_97,In_10,In_129);
nand U98 (N_98,In_456,In_593);
xnor U99 (N_99,In_142,In_1058);
xnor U100 (N_100,In_603,In_195);
nor U101 (N_101,In_1136,In_441);
and U102 (N_102,In_311,In_1167);
xnor U103 (N_103,In_1213,In_59);
and U104 (N_104,In_982,In_346);
nand U105 (N_105,In_367,In_811);
and U106 (N_106,In_379,In_497);
and U107 (N_107,In_945,In_1071);
or U108 (N_108,In_744,In_989);
nand U109 (N_109,In_509,In_793);
nand U110 (N_110,In_556,In_1030);
nor U111 (N_111,In_1422,In_663);
xnor U112 (N_112,In_1,In_1159);
and U113 (N_113,In_790,In_835);
nor U114 (N_114,In_484,In_1328);
nand U115 (N_115,In_1389,In_479);
and U116 (N_116,In_1064,In_94);
or U117 (N_117,In_519,In_1049);
and U118 (N_118,In_1434,In_667);
xnor U119 (N_119,In_753,In_85);
xor U120 (N_120,In_240,In_799);
and U121 (N_121,In_507,In_520);
nor U122 (N_122,In_143,In_1118);
xnor U123 (N_123,In_1166,In_496);
xor U124 (N_124,In_320,In_417);
nand U125 (N_125,In_1015,In_1147);
nand U126 (N_126,In_797,In_961);
and U127 (N_127,In_1254,In_1351);
nor U128 (N_128,In_726,In_866);
and U129 (N_129,In_693,In_828);
or U130 (N_130,In_1425,In_259);
xor U131 (N_131,In_88,In_105);
xor U132 (N_132,In_1394,In_1171);
or U133 (N_133,In_1163,In_179);
and U134 (N_134,In_437,In_1296);
xor U135 (N_135,In_51,In_529);
xnor U136 (N_136,In_890,In_781);
and U137 (N_137,In_501,In_37);
xor U138 (N_138,In_1242,In_874);
nand U139 (N_139,In_316,In_1121);
or U140 (N_140,In_772,In_469);
nor U141 (N_141,In_851,In_952);
or U142 (N_142,In_1318,In_356);
nand U143 (N_143,In_470,In_999);
nand U144 (N_144,In_804,In_1453);
and U145 (N_145,In_645,In_1124);
nand U146 (N_146,In_681,In_115);
nor U147 (N_147,In_355,In_592);
or U148 (N_148,In_1303,In_138);
and U149 (N_149,In_1063,In_729);
xnor U150 (N_150,In_1195,In_189);
and U151 (N_151,In_763,In_622);
xor U152 (N_152,In_157,In_869);
nand U153 (N_153,In_109,In_95);
xnor U154 (N_154,In_1485,In_1386);
nor U155 (N_155,In_26,In_1041);
nand U156 (N_156,In_272,In_1010);
and U157 (N_157,In_1353,In_528);
nand U158 (N_158,In_450,In_1347);
or U159 (N_159,In_826,In_1367);
or U160 (N_160,In_770,In_15);
nor U161 (N_161,In_601,In_1428);
nand U162 (N_162,In_803,In_1319);
xor U163 (N_163,In_161,In_610);
and U164 (N_164,In_502,In_281);
nor U165 (N_165,In_738,In_27);
xnor U166 (N_166,In_1126,In_1038);
and U167 (N_167,In_577,In_819);
and U168 (N_168,In_1379,In_1003);
or U169 (N_169,In_158,In_440);
nand U170 (N_170,In_266,In_1258);
nand U171 (N_171,In_1317,In_760);
and U172 (N_172,In_1415,In_1093);
xor U173 (N_173,In_624,In_1228);
nand U174 (N_174,In_654,In_878);
xnor U175 (N_175,In_919,In_175);
and U176 (N_176,In_757,In_387);
or U177 (N_177,In_140,In_1285);
nor U178 (N_178,In_1380,In_810);
and U179 (N_179,In_1139,In_670);
nor U180 (N_180,In_337,In_914);
or U181 (N_181,In_65,In_1269);
nand U182 (N_182,In_1260,In_332);
xnor U183 (N_183,In_98,In_749);
nand U184 (N_184,In_1382,In_1290);
or U185 (N_185,In_506,In_787);
nand U186 (N_186,In_132,In_1350);
and U187 (N_187,In_269,In_1160);
xnor U188 (N_188,In_541,In_1463);
and U189 (N_189,In_118,In_1407);
or U190 (N_190,In_1019,In_1373);
xnor U191 (N_191,In_1482,In_1455);
nor U192 (N_192,In_1162,In_75);
and U193 (N_193,In_766,In_222);
xnor U194 (N_194,In_62,In_1131);
or U195 (N_195,In_133,In_883);
nor U196 (N_196,In_588,In_453);
or U197 (N_197,In_100,In_45);
nor U198 (N_198,In_414,In_746);
nor U199 (N_199,In_959,In_578);
xor U200 (N_200,In_253,In_170);
nor U201 (N_201,In_570,In_305);
xnor U202 (N_202,In_1108,In_907);
nand U203 (N_203,In_723,In_801);
nor U204 (N_204,In_891,In_242);
or U205 (N_205,In_1366,In_183);
nand U206 (N_206,In_1332,In_644);
nor U207 (N_207,In_1277,In_515);
nor U208 (N_208,In_257,In_778);
or U209 (N_209,In_478,In_691);
and U210 (N_210,In_1096,In_701);
and U211 (N_211,In_167,In_1059);
xnor U212 (N_212,In_1387,In_333);
and U213 (N_213,In_743,In_68);
or U214 (N_214,In_261,In_653);
and U215 (N_215,In_213,In_1026);
xor U216 (N_216,In_1497,In_1419);
nand U217 (N_217,In_223,In_1472);
nor U218 (N_218,In_975,In_405);
or U219 (N_219,In_545,In_141);
nand U220 (N_220,In_427,In_632);
xnor U221 (N_221,In_1289,In_1448);
nand U222 (N_222,In_893,In_1033);
xor U223 (N_223,In_217,In_682);
xor U224 (N_224,In_1128,In_586);
nor U225 (N_225,In_537,In_407);
xnor U226 (N_226,In_689,In_872);
and U227 (N_227,In_1390,In_784);
nor U228 (N_228,In_220,In_894);
nand U229 (N_229,In_1145,In_1088);
and U230 (N_230,In_580,In_720);
nand U231 (N_231,In_193,In_651);
and U232 (N_232,In_1374,In_284);
nor U233 (N_233,In_1335,In_996);
and U234 (N_234,In_761,In_294);
or U235 (N_235,In_719,In_1035);
or U236 (N_236,In_985,In_981);
nor U237 (N_237,In_1188,In_80);
or U238 (N_238,In_1481,In_1091);
or U239 (N_239,In_549,In_1056);
nand U240 (N_240,In_1252,In_1298);
nor U241 (N_241,In_800,In_1344);
nand U242 (N_242,In_1120,In_1438);
nor U243 (N_243,In_1457,In_752);
nand U244 (N_244,In_307,In_447);
or U245 (N_245,In_256,In_243);
nor U246 (N_246,In_1368,In_1469);
nor U247 (N_247,In_9,In_558);
xor U248 (N_248,In_671,In_1288);
and U249 (N_249,In_90,In_14);
xnor U250 (N_250,In_1095,In_554);
or U251 (N_251,In_146,In_61);
nand U252 (N_252,In_1102,In_920);
nor U253 (N_253,In_1174,In_331);
and U254 (N_254,In_67,In_882);
nand U255 (N_255,In_416,In_847);
and U256 (N_256,In_1376,In_385);
or U257 (N_257,In_759,In_124);
or U258 (N_258,In_788,In_915);
or U259 (N_259,In_1262,In_1433);
and U260 (N_260,In_1138,In_1224);
nand U261 (N_261,In_268,In_718);
or U262 (N_262,In_302,In_480);
or U263 (N_263,In_822,In_1069);
or U264 (N_264,In_1279,In_1232);
or U265 (N_265,In_675,In_1381);
nor U266 (N_266,In_156,In_20);
and U267 (N_267,In_762,In_870);
nor U268 (N_268,In_1348,In_1117);
or U269 (N_269,In_633,In_377);
nor U270 (N_270,In_596,In_833);
or U271 (N_271,In_637,In_1436);
xnor U272 (N_272,In_1284,In_134);
nand U273 (N_273,In_412,In_1474);
or U274 (N_274,In_796,In_813);
xor U275 (N_275,In_508,In_838);
and U276 (N_276,In_1414,In_638);
or U277 (N_277,In_182,In_987);
or U278 (N_278,In_364,In_617);
nand U279 (N_279,In_352,In_465);
nor U280 (N_280,In_1243,In_276);
nor U281 (N_281,In_1293,In_33);
nand U282 (N_282,In_1230,In_848);
and U283 (N_283,In_461,In_184);
xor U284 (N_284,In_448,In_733);
nand U285 (N_285,In_1203,In_957);
nor U286 (N_286,In_1342,In_953);
or U287 (N_287,In_1067,In_319);
nor U288 (N_288,In_475,In_127);
nor U289 (N_289,In_32,In_938);
nor U290 (N_290,In_1238,In_946);
or U291 (N_291,In_128,In_655);
nand U292 (N_292,In_1359,In_409);
or U293 (N_293,In_338,In_1255);
or U294 (N_294,In_997,In_664);
or U295 (N_295,In_990,In_685);
nand U296 (N_296,In_849,In_4);
nand U297 (N_297,In_551,In_1154);
xor U298 (N_298,In_606,In_649);
or U299 (N_299,In_41,In_485);
nand U300 (N_300,In_438,In_126);
and U301 (N_301,In_406,In_821);
xnor U302 (N_302,In_249,In_73);
and U303 (N_303,In_735,In_1307);
and U304 (N_304,In_383,In_852);
nand U305 (N_305,In_500,In_1215);
or U306 (N_306,In_292,In_754);
nand U307 (N_307,In_93,In_1274);
and U308 (N_308,In_1046,In_1473);
and U309 (N_309,In_1259,In_751);
nor U310 (N_310,In_1354,In_1053);
nand U311 (N_311,In_198,In_1459);
xor U312 (N_312,In_330,In_477);
or U313 (N_313,In_1349,In_1236);
xor U314 (N_314,In_680,In_69);
nor U315 (N_315,In_464,In_679);
and U316 (N_316,In_993,In_844);
nor U317 (N_317,In_1125,In_1404);
nor U318 (N_318,In_618,In_374);
xor U319 (N_319,In_30,In_1068);
xor U320 (N_320,In_1198,In_1323);
nor U321 (N_321,In_306,In_258);
or U322 (N_322,In_466,In_1357);
or U323 (N_323,In_178,In_785);
nand U324 (N_324,In_998,In_1142);
nor U325 (N_325,In_1146,In_176);
and U326 (N_326,In_1111,In_1101);
xor U327 (N_327,In_160,In_1287);
nand U328 (N_328,In_399,In_327);
nand U329 (N_329,In_544,In_1047);
nand U330 (N_330,In_807,In_1207);
or U331 (N_331,In_63,In_977);
nand U332 (N_332,In_626,In_1247);
or U333 (N_333,In_543,In_559);
and U334 (N_334,In_404,In_871);
xnor U335 (N_335,In_370,In_634);
nor U336 (N_336,In_1226,In_340);
or U337 (N_337,In_1273,In_748);
or U338 (N_338,In_436,In_716);
or U339 (N_339,In_221,In_1312);
nor U340 (N_340,In_605,In_123);
xnor U341 (N_341,In_1470,In_858);
nor U342 (N_342,In_277,In_530);
nand U343 (N_343,In_1202,In_394);
xnor U344 (N_344,In_349,In_16);
xnor U345 (N_345,In_861,In_561);
xnor U346 (N_346,In_1192,In_534);
nand U347 (N_347,In_1446,In_212);
nand U348 (N_348,In_820,In_1294);
xnor U349 (N_349,In_111,In_846);
nand U350 (N_350,In_1322,In_522);
nand U351 (N_351,In_776,In_1377);
nor U352 (N_352,In_1429,In_361);
and U353 (N_353,In_773,In_646);
xor U354 (N_354,In_390,In_125);
xnor U355 (N_355,In_730,In_1383);
or U356 (N_356,In_1218,In_144);
xnor U357 (N_357,In_72,In_504);
or U358 (N_358,In_628,In_1237);
nand U359 (N_359,In_970,In_232);
nand U360 (N_360,In_488,In_1275);
or U361 (N_361,In_1089,In_755);
nand U362 (N_362,In_995,In_1370);
nor U363 (N_363,In_600,In_1081);
or U364 (N_364,In_1098,In_1362);
and U365 (N_365,In_625,In_911);
or U366 (N_366,In_343,In_92);
or U367 (N_367,In_1130,In_270);
or U368 (N_368,In_782,In_494);
nand U369 (N_369,In_876,In_991);
or U370 (N_370,In_354,In_468);
or U371 (N_371,In_408,In_1027);
and U372 (N_372,In_296,In_166);
nor U373 (N_373,In_521,In_827);
and U374 (N_374,In_1338,In_1008);
nand U375 (N_375,In_1043,In_326);
and U376 (N_376,In_282,In_935);
xnor U377 (N_377,In_1057,In_557);
nand U378 (N_378,In_1179,In_3);
nand U379 (N_379,In_1196,In_597);
nor U380 (N_380,In_325,In_54);
and U381 (N_381,In_1375,In_339);
nor U382 (N_382,In_503,In_1129);
and U383 (N_383,In_245,In_1426);
and U384 (N_384,In_721,In_493);
nand U385 (N_385,In_1184,In_555);
and U386 (N_386,In_585,In_380);
or U387 (N_387,In_462,In_1176);
and U388 (N_388,In_114,In_1087);
nor U389 (N_389,In_925,In_1051);
nand U390 (N_390,In_590,In_1173);
xnor U391 (N_391,In_1219,In_1170);
nand U392 (N_392,In_1141,In_1304);
xnor U393 (N_393,In_863,In_1392);
nor U394 (N_394,In_897,In_895);
nand U395 (N_395,In_452,In_280);
and U396 (N_396,In_728,In_1169);
nand U397 (N_397,In_423,In_208);
xnor U398 (N_398,In_1271,In_1090);
or U399 (N_399,In_1107,In_190);
nor U400 (N_400,In_252,In_1144);
and U401 (N_401,In_421,In_758);
and U402 (N_402,In_1331,In_49);
nor U403 (N_403,In_724,In_236);
or U404 (N_404,In_1291,In_376);
or U405 (N_405,In_854,In_395);
nor U406 (N_406,In_771,In_677);
nor U407 (N_407,In_974,In_712);
and U408 (N_408,In_1158,In_1187);
nand U409 (N_409,In_650,In_809);
xor U410 (N_410,In_702,In_587);
nand U411 (N_411,In_976,In_1079);
nor U412 (N_412,In_152,In_779);
xnor U413 (N_413,In_1085,In_917);
nand U414 (N_414,In_1080,In_495);
nand U415 (N_415,In_589,In_944);
or U416 (N_416,In_536,In_53);
xor U417 (N_417,In_1417,In_1214);
nand U418 (N_418,In_1208,In_298);
and U419 (N_419,In_196,In_1217);
and U420 (N_420,In_583,In_174);
and U421 (N_421,In_439,In_420);
xor U422 (N_422,In_145,In_1037);
nand U423 (N_423,In_513,In_1127);
nor U424 (N_424,In_902,In_843);
or U425 (N_425,In_1123,In_1175);
or U426 (N_426,In_473,In_986);
nand U427 (N_427,In_224,In_565);
xnor U428 (N_428,In_1484,In_1045);
nor U429 (N_429,In_540,In_2);
or U430 (N_430,In_89,In_1292);
nand U431 (N_431,In_1248,In_1148);
and U432 (N_432,In_547,In_614);
or U433 (N_433,In_392,In_322);
nor U434 (N_434,In_745,In_566);
nor U435 (N_435,In_1480,In_1371);
nor U436 (N_436,In_867,In_840);
nor U437 (N_437,In_1430,In_1253);
or U438 (N_438,In_215,In_1075);
and U439 (N_439,In_455,In_686);
nand U440 (N_440,In_487,In_6);
and U441 (N_441,In_91,In_1233);
nand U442 (N_442,In_584,In_699);
xnor U443 (N_443,In_278,In_1193);
xor U444 (N_444,In_1462,In_185);
nand U445 (N_445,In_1190,In_1398);
nor U446 (N_446,In_1231,In_786);
and U447 (N_447,In_572,In_777);
and U448 (N_448,In_1200,In_798);
nand U449 (N_449,In_727,In_696);
and U450 (N_450,In_538,In_910);
or U451 (N_451,In_552,In_381);
nand U452 (N_452,In_527,In_359);
nor U453 (N_453,In_235,In_1464);
xnor U454 (N_454,In_206,In_458);
and U455 (N_455,In_472,In_110);
and U456 (N_456,In_868,In_965);
or U457 (N_457,In_620,In_533);
nand U458 (N_458,In_397,In_1490);
and U459 (N_459,In_1440,In_824);
or U460 (N_460,In_931,In_1223);
nor U461 (N_461,In_430,In_130);
nor U462 (N_462,In_40,In_928);
or U463 (N_463,In_1212,In_1391);
or U464 (N_464,In_1444,In_1393);
and U465 (N_465,In_1337,In_814);
nand U466 (N_466,In_1024,In_1256);
nor U467 (N_467,In_1189,In_1281);
xnor U468 (N_468,In_1321,In_612);
nand U469 (N_469,In_683,In_669);
or U470 (N_470,In_279,In_363);
nor U471 (N_471,In_308,In_658);
xor U472 (N_472,In_318,In_1406);
nand U473 (N_473,In_1437,In_1445);
or U474 (N_474,In_855,In_806);
xor U475 (N_475,In_1452,In_1116);
or U476 (N_476,In_836,In_181);
and U477 (N_477,In_930,In_887);
xor U478 (N_478,In_81,In_1266);
and U479 (N_479,In_947,In_1135);
nand U480 (N_480,In_665,In_76);
xnor U481 (N_481,In_563,In_369);
nor U482 (N_482,In_1150,In_1283);
nor U483 (N_483,In_832,In_1418);
nor U484 (N_484,In_818,In_1012);
nand U485 (N_485,In_862,In_1194);
or U486 (N_486,In_1395,In_24);
nor U487 (N_487,In_831,In_1454);
and U488 (N_488,In_512,In_490);
xnor U489 (N_489,In_1113,In_948);
nor U490 (N_490,In_905,In_1061);
xor U491 (N_491,In_1122,In_285);
and U492 (N_492,In_1034,In_283);
and U493 (N_493,In_1031,In_13);
nand U494 (N_494,In_841,In_676);
and U495 (N_495,In_613,In_1432);
xor U496 (N_496,In_432,In_1106);
nand U497 (N_497,In_323,In_1065);
and U498 (N_498,In_1329,In_1109);
or U499 (N_499,In_267,In_825);
and U500 (N_500,In_731,In_12);
xor U501 (N_501,In_312,In_1487);
nand U502 (N_502,In_1450,In_401);
xnor U503 (N_503,In_690,In_290);
nor U504 (N_504,In_904,In_234);
and U505 (N_505,In_1039,In_1021);
xor U506 (N_506,In_1316,In_260);
and U507 (N_507,In_1066,In_1278);
xnor U508 (N_508,In_805,In_1206);
or U509 (N_509,In_1302,In_1334);
or U510 (N_510,In_1427,In_511);
or U511 (N_511,In_297,In_860);
and U512 (N_512,In_1411,In_926);
nand U513 (N_513,In_873,In_1409);
xnor U514 (N_514,In_913,In_783);
and U515 (N_515,In_200,In_888);
xnor U516 (N_516,In_1000,In_301);
and U517 (N_517,In_216,In_943);
and U518 (N_518,In_474,In_1282);
and U519 (N_519,In_64,In_966);
nand U520 (N_520,In_1225,In_1220);
or U521 (N_521,In_60,In_886);
and U522 (N_522,In_113,In_1489);
or U523 (N_523,In_713,In_373);
nor U524 (N_524,In_324,In_591);
nand U525 (N_525,In_774,In_789);
nand U526 (N_526,In_546,In_1009);
and U527 (N_527,In_172,In_979);
and U528 (N_528,In_102,In_598);
or U529 (N_529,In_1265,In_684);
nand U530 (N_530,In_304,In_418);
nor U531 (N_531,In_1165,In_99);
nor U532 (N_532,In_250,In_1222);
or U533 (N_533,In_459,In_845);
nor U534 (N_534,In_1201,In_1022);
nand U535 (N_535,In_823,In_1365);
or U536 (N_536,In_362,In_1092);
xor U537 (N_537,In_568,In_949);
xor U538 (N_538,In_1105,In_674);
and U539 (N_539,In_321,In_169);
nor U540 (N_540,In_710,In_1451);
and U541 (N_541,In_1155,In_687);
or U542 (N_542,In_358,In_922);
xnor U543 (N_543,In_210,In_988);
nand U544 (N_544,In_334,In_1272);
nand U545 (N_545,In_1361,In_255);
xnor U546 (N_546,In_666,In_659);
nand U547 (N_547,In_535,In_1276);
nor U548 (N_548,In_615,In_1499);
xnor U549 (N_549,In_936,In_747);
nand U550 (N_550,In_177,In_1486);
and U551 (N_551,In_972,In_1050);
or U552 (N_552,In_58,In_1336);
nand U553 (N_553,In_107,In_523);
xnor U554 (N_554,In_275,In_1369);
xnor U555 (N_555,In_47,In_328);
xnor U556 (N_556,In_627,In_765);
xnor U557 (N_557,In_1245,In_96);
xor U558 (N_558,In_310,In_817);
and U559 (N_559,In_192,In_274);
nand U560 (N_560,In_454,In_288);
nand U561 (N_561,In_1327,In_742);
or U562 (N_562,In_446,In_291);
xnor U563 (N_563,In_510,In_1094);
or U564 (N_564,In_378,In_23);
nor U565 (N_565,In_424,In_233);
nand U566 (N_566,In_431,In_1384);
nor U567 (N_567,In_569,In_725);
nand U568 (N_568,In_526,In_28);
nand U569 (N_569,In_1197,In_21);
nor U570 (N_570,In_595,In_386);
xor U571 (N_571,In_163,In_74);
nand U572 (N_572,In_11,In_885);
nand U573 (N_573,In_1270,In_1435);
xor U574 (N_574,In_1421,In_630);
nand U575 (N_575,In_211,In_629);
nand U576 (N_576,In_1014,In_119);
and U577 (N_577,In_44,In_101);
or U578 (N_578,In_1424,In_42);
nand U579 (N_579,In_429,In_286);
and U580 (N_580,In_203,In_621);
and U581 (N_581,In_661,In_576);
nand U582 (N_582,In_1052,In_1060);
nor U583 (N_583,In_159,In_131);
or U584 (N_584,In_1449,In_135);
or U585 (N_585,In_657,In_542);
nor U586 (N_586,In_1044,In_457);
and U587 (N_587,In_400,In_1020);
or U588 (N_588,In_1132,In_1185);
nor U589 (N_589,In_978,In_1324);
nand U590 (N_590,In_351,In_25);
nor U591 (N_591,In_1140,In_1413);
nand U592 (N_592,In_106,In_499);
or U593 (N_593,In_1070,In_705);
and U594 (N_594,In_31,In_1227);
xor U595 (N_595,In_717,In_1358);
nand U596 (N_596,In_1308,In_1396);
or U597 (N_597,In_967,In_1210);
and U598 (N_598,In_516,In_1234);
nor U599 (N_599,In_1471,In_1498);
nand U600 (N_600,In_491,In_1263);
and U601 (N_601,In_197,In_739);
xor U602 (N_602,In_8,In_1011);
xor U603 (N_603,In_353,In_1177);
or U604 (N_604,In_498,In_271);
xnor U605 (N_605,In_992,In_136);
or U606 (N_606,In_631,In_884);
nand U607 (N_607,In_1333,In_1002);
nor U608 (N_608,In_104,In_460);
nor U609 (N_609,In_1180,In_151);
nor U610 (N_610,In_734,In_1468);
or U611 (N_611,In_956,In_1054);
or U612 (N_612,In_1431,In_1005);
xor U613 (N_613,In_1355,In_205);
nor U614 (N_614,In_449,In_619);
and U615 (N_615,In_1443,In_1072);
or U616 (N_616,In_1267,In_56);
nor U617 (N_617,In_875,In_1408);
or U618 (N_618,In_1100,In_1299);
nor U619 (N_619,In_402,In_70);
nand U620 (N_620,In_1017,In_635);
and U621 (N_621,In_1442,In_1082);
nand U622 (N_622,In_149,In_1164);
and U623 (N_623,In_228,In_492);
xnor U624 (N_624,In_929,In_1397);
or U625 (N_625,In_248,In_1360);
nor U626 (N_626,In_1151,In_942);
xor U627 (N_627,In_428,In_77);
nor U628 (N_628,In_1494,In_442);
nand U629 (N_629,In_48,In_1104);
nand U630 (N_630,In_329,In_112);
or U631 (N_631,In_1495,In_1001);
or U632 (N_632,In_1309,In_171);
nor U633 (N_633,In_1412,In_1149);
xor U634 (N_634,In_1114,In_1295);
and U635 (N_635,In_121,In_1492);
and U636 (N_636,In_238,In_1153);
nand U637 (N_637,In_289,In_422);
nor U638 (N_638,In_299,In_219);
nor U639 (N_639,In_108,In_391);
xnor U640 (N_640,In_1466,In_116);
nand U641 (N_641,In_609,In_264);
nand U642 (N_642,In_186,In_1191);
and U643 (N_643,In_927,In_1023);
nor U644 (N_644,In_648,In_313);
nor U645 (N_645,In_209,In_1157);
xnor U646 (N_646,In_1013,In_636);
or U647 (N_647,In_38,In_517);
and U648 (N_648,In_780,In_372);
or U649 (N_649,In_180,In_188);
xor U650 (N_650,In_737,In_955);
nor U651 (N_651,In_1280,In_262);
xnor U652 (N_652,In_969,In_704);
nand U653 (N_653,In_382,In_365);
xnor U654 (N_654,In_692,In_1372);
and U655 (N_655,In_1341,In_1204);
or U656 (N_656,In_918,In_560);
and U657 (N_657,In_410,In_341);
nor U658 (N_658,In_443,In_120);
xor U659 (N_659,In_1240,In_1073);
nor U660 (N_660,In_1182,In_1137);
or U661 (N_661,In_403,In_194);
nor U662 (N_662,In_1326,In_204);
nor U663 (N_663,In_342,In_19);
or U664 (N_664,In_1172,In_714);
or U665 (N_665,In_1199,In_1297);
or U666 (N_666,In_1161,In_57);
nand U667 (N_667,In_1475,In_36);
xor U668 (N_668,In_168,In_52);
nand U669 (N_669,In_1007,In_218);
xnor U670 (N_670,In_396,In_812);
nor U671 (N_671,In_709,In_950);
nand U672 (N_672,In_295,In_1447);
and U673 (N_673,In_940,In_795);
or U674 (N_674,In_155,In_963);
nor U675 (N_675,In_736,In_445);
or U676 (N_676,In_1006,In_137);
and U677 (N_677,In_1405,In_1103);
xnor U678 (N_678,In_971,In_173);
and U679 (N_679,In_1062,In_1479);
and U680 (N_680,In_1423,In_388);
xor U681 (N_681,In_476,In_467);
nand U682 (N_682,In_857,In_1178);
xor U683 (N_683,In_879,In_1183);
or U684 (N_684,In_43,In_815);
nor U685 (N_685,In_662,In_912);
and U686 (N_686,In_1320,In_707);
or U687 (N_687,In_694,In_309);
and U688 (N_688,In_50,In_1352);
and U689 (N_689,In_856,In_623);
nor U690 (N_690,In_1261,In_1478);
and U691 (N_691,In_246,In_336);
and U692 (N_692,In_434,In_567);
nand U693 (N_693,In_226,In_1378);
nor U694 (N_694,In_934,In_1477);
xor U695 (N_695,In_903,In_199);
nor U696 (N_696,In_263,In_673);
nor U697 (N_697,In_483,In_1074);
nand U698 (N_698,In_656,In_968);
or U699 (N_699,In_1112,In_230);
nor U700 (N_700,In_82,In_1401);
and U701 (N_701,In_1439,In_239);
or U702 (N_702,In_1097,In_1268);
or U703 (N_703,In_1483,In_164);
xor U704 (N_704,In_486,In_672);
nand U705 (N_705,In_1345,In_700);
or U706 (N_706,In_66,In_1325);
xor U707 (N_707,In_225,In_413);
and U708 (N_708,In_1311,In_419);
and U709 (N_709,In_39,In_994);
or U710 (N_710,In_722,In_575);
nor U711 (N_711,In_703,In_231);
nor U712 (N_712,In_247,In_932);
or U713 (N_713,In_611,In_941);
and U714 (N_714,In_829,In_708);
or U715 (N_715,In_335,In_1032);
xnor U716 (N_716,In_791,In_1364);
and U717 (N_717,In_254,In_1314);
and U718 (N_718,In_214,In_139);
or U719 (N_719,In_1385,In_1016);
and U720 (N_720,In_229,In_1048);
and U721 (N_721,In_1251,In_1488);
or U722 (N_722,In_706,In_1076);
nand U723 (N_723,In_652,In_1134);
nor U724 (N_724,In_241,In_344);
xnor U725 (N_725,In_162,In_916);
and U726 (N_726,In_1301,In_463);
nor U727 (N_727,In_695,In_1216);
and U728 (N_728,In_639,In_642);
xnor U729 (N_729,In_35,In_368);
xnor U730 (N_730,In_315,In_303);
xnor U731 (N_731,In_951,In_1186);
xor U732 (N_732,In_1399,In_1441);
or U733 (N_733,In_55,In_357);
nor U734 (N_734,In_1229,In_147);
and U735 (N_735,In_83,In_958);
nor U736 (N_736,In_1286,In_1036);
xnor U737 (N_737,In_1363,In_1221);
and U738 (N_738,In_983,In_1493);
xnor U739 (N_739,In_1156,In_393);
xor U740 (N_740,In_1458,In_1496);
nor U741 (N_741,In_244,In_550);
nor U742 (N_742,In_604,In_505);
nor U743 (N_743,In_960,In_287);
or U744 (N_744,In_1168,In_481);
nand U745 (N_745,In_678,In_688);
or U746 (N_746,In_46,In_482);
nand U747 (N_747,In_808,In_741);
and U748 (N_748,In_750,In_1078);
xor U749 (N_749,In_1209,In_908);
xnor U750 (N_750,In_1166,In_820);
or U751 (N_751,In_936,In_89);
xor U752 (N_752,In_456,In_801);
or U753 (N_753,In_389,In_466);
nand U754 (N_754,In_1214,In_390);
nor U755 (N_755,In_306,In_1311);
or U756 (N_756,In_353,In_473);
nand U757 (N_757,In_723,In_1221);
and U758 (N_758,In_393,In_1037);
or U759 (N_759,In_343,In_494);
nor U760 (N_760,In_725,In_73);
and U761 (N_761,In_297,In_169);
or U762 (N_762,In_673,In_172);
nor U763 (N_763,In_471,In_1472);
nor U764 (N_764,In_514,In_341);
nor U765 (N_765,In_1000,In_392);
xor U766 (N_766,In_1103,In_424);
nor U767 (N_767,In_1497,In_649);
nand U768 (N_768,In_931,In_336);
nand U769 (N_769,In_1401,In_970);
nand U770 (N_770,In_600,In_1210);
nor U771 (N_771,In_244,In_616);
xnor U772 (N_772,In_1046,In_591);
nand U773 (N_773,In_833,In_669);
and U774 (N_774,In_1260,In_810);
or U775 (N_775,In_1103,In_382);
nor U776 (N_776,In_303,In_131);
and U777 (N_777,In_440,In_29);
xor U778 (N_778,In_590,In_363);
and U779 (N_779,In_259,In_283);
xor U780 (N_780,In_503,In_858);
nor U781 (N_781,In_1377,In_9);
nor U782 (N_782,In_829,In_1159);
nand U783 (N_783,In_462,In_581);
or U784 (N_784,In_272,In_892);
nand U785 (N_785,In_1425,In_734);
xnor U786 (N_786,In_147,In_397);
and U787 (N_787,In_1155,In_1241);
or U788 (N_788,In_1230,In_779);
nor U789 (N_789,In_346,In_1032);
nor U790 (N_790,In_1113,In_518);
xor U791 (N_791,In_904,In_875);
nor U792 (N_792,In_901,In_908);
or U793 (N_793,In_52,In_1437);
xnor U794 (N_794,In_894,In_1287);
nand U795 (N_795,In_470,In_1437);
or U796 (N_796,In_549,In_284);
and U797 (N_797,In_56,In_40);
and U798 (N_798,In_1169,In_784);
or U799 (N_799,In_708,In_891);
xnor U800 (N_800,In_308,In_1196);
nand U801 (N_801,In_603,In_987);
xor U802 (N_802,In_1182,In_15);
xnor U803 (N_803,In_1137,In_636);
or U804 (N_804,In_6,In_1054);
and U805 (N_805,In_557,In_1327);
xor U806 (N_806,In_13,In_410);
or U807 (N_807,In_788,In_745);
or U808 (N_808,In_1046,In_481);
xor U809 (N_809,In_281,In_313);
or U810 (N_810,In_229,In_963);
nand U811 (N_811,In_1451,In_1050);
nand U812 (N_812,In_1319,In_694);
and U813 (N_813,In_117,In_285);
and U814 (N_814,In_1375,In_241);
nor U815 (N_815,In_1372,In_894);
nand U816 (N_816,In_500,In_645);
xnor U817 (N_817,In_799,In_1476);
nand U818 (N_818,In_971,In_112);
and U819 (N_819,In_1344,In_324);
or U820 (N_820,In_1413,In_137);
or U821 (N_821,In_166,In_1419);
nor U822 (N_822,In_1359,In_368);
or U823 (N_823,In_525,In_930);
nor U824 (N_824,In_792,In_1389);
nand U825 (N_825,In_283,In_1264);
or U826 (N_826,In_1243,In_790);
nand U827 (N_827,In_239,In_1298);
nor U828 (N_828,In_1394,In_372);
or U829 (N_829,In_1116,In_958);
or U830 (N_830,In_1112,In_190);
xor U831 (N_831,In_1377,In_349);
xor U832 (N_832,In_84,In_558);
nor U833 (N_833,In_669,In_1150);
or U834 (N_834,In_100,In_1321);
xor U835 (N_835,In_1285,In_536);
nand U836 (N_836,In_344,In_398);
xnor U837 (N_837,In_1308,In_1474);
nor U838 (N_838,In_474,In_115);
and U839 (N_839,In_547,In_1306);
xnor U840 (N_840,In_897,In_323);
or U841 (N_841,In_49,In_170);
nor U842 (N_842,In_942,In_491);
nand U843 (N_843,In_14,In_820);
or U844 (N_844,In_963,In_1407);
and U845 (N_845,In_890,In_661);
nand U846 (N_846,In_1075,In_1162);
nor U847 (N_847,In_896,In_495);
or U848 (N_848,In_592,In_1026);
and U849 (N_849,In_1040,In_1415);
xor U850 (N_850,In_1395,In_255);
nor U851 (N_851,In_1055,In_168);
xnor U852 (N_852,In_857,In_729);
xor U853 (N_853,In_710,In_521);
or U854 (N_854,In_576,In_14);
xnor U855 (N_855,In_1125,In_293);
nand U856 (N_856,In_1278,In_1294);
nor U857 (N_857,In_491,In_108);
nand U858 (N_858,In_900,In_1251);
nor U859 (N_859,In_0,In_62);
or U860 (N_860,In_505,In_493);
or U861 (N_861,In_495,In_1302);
nor U862 (N_862,In_226,In_389);
nor U863 (N_863,In_576,In_485);
or U864 (N_864,In_264,In_1095);
nand U865 (N_865,In_845,In_657);
and U866 (N_866,In_1312,In_348);
nand U867 (N_867,In_200,In_931);
nor U868 (N_868,In_960,In_938);
xnor U869 (N_869,In_971,In_1032);
nand U870 (N_870,In_981,In_276);
nand U871 (N_871,In_609,In_295);
xor U872 (N_872,In_354,In_1096);
and U873 (N_873,In_118,In_61);
or U874 (N_874,In_304,In_196);
and U875 (N_875,In_186,In_1329);
and U876 (N_876,In_134,In_1261);
nor U877 (N_877,In_172,In_757);
nor U878 (N_878,In_122,In_1015);
nand U879 (N_879,In_1428,In_1313);
nor U880 (N_880,In_184,In_1013);
nand U881 (N_881,In_1067,In_887);
nand U882 (N_882,In_934,In_1492);
nand U883 (N_883,In_352,In_1379);
nor U884 (N_884,In_1392,In_802);
nand U885 (N_885,In_266,In_1213);
or U886 (N_886,In_956,In_734);
nand U887 (N_887,In_356,In_1315);
and U888 (N_888,In_838,In_1171);
nor U889 (N_889,In_1199,In_687);
and U890 (N_890,In_62,In_163);
xnor U891 (N_891,In_600,In_967);
xnor U892 (N_892,In_1201,In_1021);
and U893 (N_893,In_255,In_1077);
and U894 (N_894,In_512,In_742);
and U895 (N_895,In_1218,In_810);
nand U896 (N_896,In_761,In_88);
nor U897 (N_897,In_931,In_118);
xnor U898 (N_898,In_353,In_1102);
nand U899 (N_899,In_1390,In_580);
xnor U900 (N_900,In_974,In_983);
nor U901 (N_901,In_1025,In_1210);
xor U902 (N_902,In_1297,In_840);
xnor U903 (N_903,In_372,In_1039);
xnor U904 (N_904,In_422,In_1279);
or U905 (N_905,In_1438,In_1105);
and U906 (N_906,In_480,In_1138);
nor U907 (N_907,In_513,In_1490);
nor U908 (N_908,In_1126,In_1180);
xnor U909 (N_909,In_872,In_778);
nor U910 (N_910,In_278,In_547);
and U911 (N_911,In_835,In_408);
xnor U912 (N_912,In_731,In_1480);
nor U913 (N_913,In_964,In_1026);
and U914 (N_914,In_128,In_176);
nor U915 (N_915,In_1178,In_157);
nor U916 (N_916,In_783,In_1035);
nor U917 (N_917,In_766,In_1298);
and U918 (N_918,In_160,In_484);
xor U919 (N_919,In_767,In_1469);
nand U920 (N_920,In_797,In_1109);
nand U921 (N_921,In_140,In_704);
xor U922 (N_922,In_1039,In_833);
nor U923 (N_923,In_362,In_1006);
or U924 (N_924,In_506,In_953);
or U925 (N_925,In_1291,In_764);
nand U926 (N_926,In_1011,In_1005);
or U927 (N_927,In_1296,In_635);
nand U928 (N_928,In_1457,In_210);
and U929 (N_929,In_741,In_1341);
nand U930 (N_930,In_1193,In_252);
nor U931 (N_931,In_1270,In_390);
or U932 (N_932,In_1330,In_1354);
nor U933 (N_933,In_1371,In_1460);
xnor U934 (N_934,In_6,In_595);
xnor U935 (N_935,In_1085,In_245);
or U936 (N_936,In_476,In_732);
nand U937 (N_937,In_1414,In_1494);
and U938 (N_938,In_496,In_553);
xnor U939 (N_939,In_1192,In_395);
and U940 (N_940,In_424,In_825);
and U941 (N_941,In_622,In_1123);
or U942 (N_942,In_1129,In_1030);
nand U943 (N_943,In_922,In_1031);
and U944 (N_944,In_260,In_1312);
xnor U945 (N_945,In_1215,In_1492);
nor U946 (N_946,In_92,In_1456);
xor U947 (N_947,In_758,In_1223);
nor U948 (N_948,In_958,In_182);
nor U949 (N_949,In_271,In_41);
nor U950 (N_950,In_843,In_1406);
nand U951 (N_951,In_273,In_1479);
and U952 (N_952,In_332,In_384);
nand U953 (N_953,In_181,In_358);
or U954 (N_954,In_715,In_1038);
nand U955 (N_955,In_1382,In_126);
xnor U956 (N_956,In_502,In_39);
nor U957 (N_957,In_443,In_256);
xnor U958 (N_958,In_1337,In_24);
or U959 (N_959,In_875,In_416);
xor U960 (N_960,In_1026,In_1464);
nand U961 (N_961,In_577,In_573);
and U962 (N_962,In_1237,In_1486);
or U963 (N_963,In_52,In_1146);
xnor U964 (N_964,In_297,In_888);
xnor U965 (N_965,In_1222,In_353);
nor U966 (N_966,In_725,In_439);
nor U967 (N_967,In_1105,In_1239);
nor U968 (N_968,In_1032,In_1389);
or U969 (N_969,In_156,In_786);
nand U970 (N_970,In_515,In_247);
and U971 (N_971,In_919,In_57);
xor U972 (N_972,In_360,In_1091);
and U973 (N_973,In_855,In_956);
and U974 (N_974,In_294,In_648);
and U975 (N_975,In_88,In_1472);
or U976 (N_976,In_362,In_1336);
nand U977 (N_977,In_996,In_991);
and U978 (N_978,In_500,In_432);
and U979 (N_979,In_716,In_836);
nor U980 (N_980,In_485,In_1285);
xor U981 (N_981,In_579,In_29);
or U982 (N_982,In_126,In_327);
and U983 (N_983,In_46,In_115);
nand U984 (N_984,In_1358,In_309);
nand U985 (N_985,In_753,In_1064);
and U986 (N_986,In_979,In_1438);
and U987 (N_987,In_465,In_666);
or U988 (N_988,In_257,In_694);
nor U989 (N_989,In_935,In_614);
xor U990 (N_990,In_374,In_182);
xor U991 (N_991,In_1107,In_619);
or U992 (N_992,In_1120,In_1010);
and U993 (N_993,In_137,In_211);
or U994 (N_994,In_257,In_1131);
or U995 (N_995,In_233,In_409);
xor U996 (N_996,In_976,In_1080);
and U997 (N_997,In_1025,In_145);
nor U998 (N_998,In_1194,In_1297);
nand U999 (N_999,In_1239,In_1492);
nand U1000 (N_1000,In_32,In_1396);
nand U1001 (N_1001,In_41,In_1038);
or U1002 (N_1002,In_644,In_1151);
or U1003 (N_1003,In_561,In_1440);
nor U1004 (N_1004,In_1077,In_694);
and U1005 (N_1005,In_1499,In_1005);
nand U1006 (N_1006,In_1235,In_1187);
or U1007 (N_1007,In_1339,In_978);
xor U1008 (N_1008,In_107,In_259);
and U1009 (N_1009,In_1173,In_9);
xor U1010 (N_1010,In_92,In_1395);
and U1011 (N_1011,In_175,In_239);
and U1012 (N_1012,In_313,In_1433);
and U1013 (N_1013,In_327,In_647);
nor U1014 (N_1014,In_717,In_711);
and U1015 (N_1015,In_432,In_1466);
xnor U1016 (N_1016,In_617,In_1253);
nor U1017 (N_1017,In_411,In_975);
nor U1018 (N_1018,In_154,In_569);
nand U1019 (N_1019,In_875,In_1106);
nor U1020 (N_1020,In_325,In_976);
xor U1021 (N_1021,In_1485,In_1444);
nand U1022 (N_1022,In_1459,In_917);
xnor U1023 (N_1023,In_1232,In_987);
or U1024 (N_1024,In_450,In_969);
or U1025 (N_1025,In_312,In_240);
nand U1026 (N_1026,In_1043,In_914);
nor U1027 (N_1027,In_105,In_78);
xnor U1028 (N_1028,In_306,In_712);
nor U1029 (N_1029,In_218,In_106);
nand U1030 (N_1030,In_1025,In_824);
nand U1031 (N_1031,In_307,In_1344);
and U1032 (N_1032,In_511,In_913);
and U1033 (N_1033,In_703,In_1294);
nor U1034 (N_1034,In_672,In_556);
and U1035 (N_1035,In_296,In_792);
nand U1036 (N_1036,In_567,In_11);
xor U1037 (N_1037,In_831,In_1247);
or U1038 (N_1038,In_1405,In_1492);
nand U1039 (N_1039,In_70,In_1035);
and U1040 (N_1040,In_445,In_1057);
nor U1041 (N_1041,In_1271,In_854);
or U1042 (N_1042,In_338,In_451);
or U1043 (N_1043,In_561,In_566);
or U1044 (N_1044,In_261,In_744);
nand U1045 (N_1045,In_417,In_440);
or U1046 (N_1046,In_244,In_822);
or U1047 (N_1047,In_1300,In_186);
xor U1048 (N_1048,In_807,In_892);
and U1049 (N_1049,In_400,In_379);
nor U1050 (N_1050,In_365,In_1206);
and U1051 (N_1051,In_1261,In_530);
and U1052 (N_1052,In_539,In_1317);
or U1053 (N_1053,In_1275,In_292);
nor U1054 (N_1054,In_1181,In_994);
and U1055 (N_1055,In_1352,In_231);
and U1056 (N_1056,In_329,In_138);
nor U1057 (N_1057,In_199,In_1257);
nor U1058 (N_1058,In_191,In_532);
or U1059 (N_1059,In_698,In_851);
xnor U1060 (N_1060,In_950,In_1307);
or U1061 (N_1061,In_262,In_279);
nor U1062 (N_1062,In_1311,In_1435);
nand U1063 (N_1063,In_560,In_802);
nand U1064 (N_1064,In_58,In_1095);
nor U1065 (N_1065,In_45,In_1016);
nand U1066 (N_1066,In_448,In_80);
and U1067 (N_1067,In_961,In_555);
or U1068 (N_1068,In_1137,In_1286);
nand U1069 (N_1069,In_1239,In_14);
nor U1070 (N_1070,In_155,In_1186);
nor U1071 (N_1071,In_574,In_839);
nand U1072 (N_1072,In_958,In_1344);
xor U1073 (N_1073,In_361,In_1469);
nand U1074 (N_1074,In_1430,In_712);
nor U1075 (N_1075,In_235,In_1270);
nand U1076 (N_1076,In_443,In_532);
and U1077 (N_1077,In_1300,In_614);
or U1078 (N_1078,In_896,In_376);
xor U1079 (N_1079,In_1086,In_918);
nand U1080 (N_1080,In_1380,In_746);
nor U1081 (N_1081,In_683,In_1076);
nand U1082 (N_1082,In_616,In_121);
or U1083 (N_1083,In_916,In_732);
and U1084 (N_1084,In_1489,In_1321);
or U1085 (N_1085,In_506,In_1034);
nor U1086 (N_1086,In_641,In_1462);
nor U1087 (N_1087,In_277,In_1382);
xnor U1088 (N_1088,In_488,In_178);
nand U1089 (N_1089,In_1072,In_765);
xor U1090 (N_1090,In_1323,In_1039);
nand U1091 (N_1091,In_262,In_694);
xnor U1092 (N_1092,In_698,In_1103);
nand U1093 (N_1093,In_1378,In_1000);
nor U1094 (N_1094,In_482,In_644);
or U1095 (N_1095,In_420,In_318);
nand U1096 (N_1096,In_185,In_732);
or U1097 (N_1097,In_267,In_274);
nor U1098 (N_1098,In_193,In_859);
nand U1099 (N_1099,In_853,In_1234);
nand U1100 (N_1100,In_316,In_1432);
and U1101 (N_1101,In_299,In_697);
and U1102 (N_1102,In_505,In_731);
or U1103 (N_1103,In_1390,In_38);
xor U1104 (N_1104,In_1320,In_792);
nor U1105 (N_1105,In_1452,In_35);
xnor U1106 (N_1106,In_766,In_916);
xor U1107 (N_1107,In_1162,In_171);
xnor U1108 (N_1108,In_506,In_1023);
or U1109 (N_1109,In_179,In_1307);
nand U1110 (N_1110,In_926,In_20);
or U1111 (N_1111,In_1078,In_1323);
and U1112 (N_1112,In_448,In_259);
nor U1113 (N_1113,In_1213,In_1211);
or U1114 (N_1114,In_1339,In_763);
or U1115 (N_1115,In_515,In_1114);
and U1116 (N_1116,In_415,In_22);
nand U1117 (N_1117,In_943,In_1418);
nor U1118 (N_1118,In_1419,In_1130);
xor U1119 (N_1119,In_829,In_923);
xnor U1120 (N_1120,In_505,In_633);
xor U1121 (N_1121,In_325,In_728);
or U1122 (N_1122,In_1152,In_1117);
or U1123 (N_1123,In_954,In_1195);
or U1124 (N_1124,In_791,In_1211);
nand U1125 (N_1125,In_1427,In_1225);
nor U1126 (N_1126,In_994,In_699);
xor U1127 (N_1127,In_291,In_715);
nor U1128 (N_1128,In_898,In_139);
nand U1129 (N_1129,In_738,In_75);
nand U1130 (N_1130,In_351,In_575);
and U1131 (N_1131,In_323,In_1113);
or U1132 (N_1132,In_487,In_737);
nor U1133 (N_1133,In_39,In_1352);
and U1134 (N_1134,In_87,In_1339);
nand U1135 (N_1135,In_1130,In_931);
nand U1136 (N_1136,In_1306,In_170);
xnor U1137 (N_1137,In_576,In_1102);
and U1138 (N_1138,In_849,In_555);
xnor U1139 (N_1139,In_594,In_1351);
and U1140 (N_1140,In_729,In_1105);
or U1141 (N_1141,In_864,In_1325);
nand U1142 (N_1142,In_143,In_239);
xnor U1143 (N_1143,In_413,In_951);
xnor U1144 (N_1144,In_127,In_1381);
or U1145 (N_1145,In_618,In_884);
nor U1146 (N_1146,In_751,In_215);
and U1147 (N_1147,In_35,In_1479);
and U1148 (N_1148,In_1059,In_1297);
and U1149 (N_1149,In_1205,In_906);
and U1150 (N_1150,In_124,In_1324);
nor U1151 (N_1151,In_632,In_566);
or U1152 (N_1152,In_157,In_259);
nor U1153 (N_1153,In_35,In_110);
nor U1154 (N_1154,In_650,In_118);
xnor U1155 (N_1155,In_493,In_679);
and U1156 (N_1156,In_1402,In_180);
xor U1157 (N_1157,In_1003,In_451);
xor U1158 (N_1158,In_561,In_85);
and U1159 (N_1159,In_1074,In_32);
xor U1160 (N_1160,In_1065,In_438);
and U1161 (N_1161,In_248,In_1243);
nor U1162 (N_1162,In_829,In_557);
xnor U1163 (N_1163,In_28,In_520);
nand U1164 (N_1164,In_1008,In_5);
or U1165 (N_1165,In_985,In_25);
xnor U1166 (N_1166,In_41,In_1041);
and U1167 (N_1167,In_1041,In_136);
and U1168 (N_1168,In_983,In_232);
xnor U1169 (N_1169,In_1016,In_552);
xnor U1170 (N_1170,In_1304,In_1467);
nor U1171 (N_1171,In_691,In_1210);
nor U1172 (N_1172,In_955,In_1027);
xnor U1173 (N_1173,In_1224,In_110);
nor U1174 (N_1174,In_952,In_435);
or U1175 (N_1175,In_199,In_148);
xnor U1176 (N_1176,In_188,In_1452);
nor U1177 (N_1177,In_573,In_746);
xnor U1178 (N_1178,In_940,In_1460);
nand U1179 (N_1179,In_885,In_784);
and U1180 (N_1180,In_594,In_895);
nand U1181 (N_1181,In_655,In_347);
xnor U1182 (N_1182,In_1451,In_243);
nor U1183 (N_1183,In_81,In_902);
xnor U1184 (N_1184,In_262,In_268);
nor U1185 (N_1185,In_1420,In_636);
or U1186 (N_1186,In_1146,In_1199);
and U1187 (N_1187,In_1433,In_987);
xnor U1188 (N_1188,In_211,In_185);
or U1189 (N_1189,In_267,In_432);
and U1190 (N_1190,In_230,In_329);
nor U1191 (N_1191,In_204,In_700);
or U1192 (N_1192,In_1099,In_486);
nand U1193 (N_1193,In_643,In_783);
nand U1194 (N_1194,In_942,In_750);
nand U1195 (N_1195,In_1083,In_983);
or U1196 (N_1196,In_1304,In_290);
or U1197 (N_1197,In_668,In_1319);
xnor U1198 (N_1198,In_138,In_1064);
and U1199 (N_1199,In_565,In_171);
and U1200 (N_1200,In_92,In_139);
or U1201 (N_1201,In_313,In_798);
nor U1202 (N_1202,In_1431,In_10);
nor U1203 (N_1203,In_454,In_780);
or U1204 (N_1204,In_582,In_1127);
nand U1205 (N_1205,In_1020,In_603);
nor U1206 (N_1206,In_619,In_570);
nor U1207 (N_1207,In_202,In_1058);
or U1208 (N_1208,In_473,In_312);
xor U1209 (N_1209,In_1299,In_1129);
and U1210 (N_1210,In_169,In_869);
and U1211 (N_1211,In_653,In_792);
xnor U1212 (N_1212,In_1382,In_142);
xor U1213 (N_1213,In_840,In_1144);
xnor U1214 (N_1214,In_1318,In_39);
or U1215 (N_1215,In_857,In_616);
nor U1216 (N_1216,In_805,In_914);
and U1217 (N_1217,In_1323,In_198);
xnor U1218 (N_1218,In_565,In_984);
nor U1219 (N_1219,In_390,In_1326);
or U1220 (N_1220,In_355,In_1378);
or U1221 (N_1221,In_753,In_685);
and U1222 (N_1222,In_714,In_447);
and U1223 (N_1223,In_1260,In_856);
xnor U1224 (N_1224,In_171,In_256);
nor U1225 (N_1225,In_1494,In_1452);
nor U1226 (N_1226,In_300,In_1274);
xor U1227 (N_1227,In_424,In_1438);
nand U1228 (N_1228,In_524,In_789);
xor U1229 (N_1229,In_231,In_758);
nand U1230 (N_1230,In_989,In_1120);
and U1231 (N_1231,In_289,In_612);
nand U1232 (N_1232,In_444,In_458);
or U1233 (N_1233,In_419,In_668);
and U1234 (N_1234,In_1469,In_831);
nand U1235 (N_1235,In_1344,In_832);
nor U1236 (N_1236,In_330,In_395);
xor U1237 (N_1237,In_1455,In_1195);
and U1238 (N_1238,In_1203,In_1003);
or U1239 (N_1239,In_528,In_60);
or U1240 (N_1240,In_88,In_3);
or U1241 (N_1241,In_102,In_239);
and U1242 (N_1242,In_393,In_700);
nor U1243 (N_1243,In_931,In_65);
xor U1244 (N_1244,In_751,In_1068);
or U1245 (N_1245,In_1364,In_1376);
xor U1246 (N_1246,In_1492,In_1085);
or U1247 (N_1247,In_216,In_123);
nand U1248 (N_1248,In_1410,In_958);
nor U1249 (N_1249,In_216,In_752);
nor U1250 (N_1250,In_64,In_155);
nand U1251 (N_1251,In_1402,In_415);
nand U1252 (N_1252,In_1417,In_320);
or U1253 (N_1253,In_679,In_584);
nor U1254 (N_1254,In_271,In_1070);
xor U1255 (N_1255,In_787,In_399);
and U1256 (N_1256,In_939,In_1140);
xnor U1257 (N_1257,In_743,In_60);
nand U1258 (N_1258,In_1054,In_505);
or U1259 (N_1259,In_674,In_1176);
or U1260 (N_1260,In_1016,In_150);
and U1261 (N_1261,In_198,In_1107);
xnor U1262 (N_1262,In_486,In_1137);
xnor U1263 (N_1263,In_482,In_794);
nand U1264 (N_1264,In_297,In_187);
and U1265 (N_1265,In_1218,In_1214);
nor U1266 (N_1266,In_1211,In_589);
nand U1267 (N_1267,In_1007,In_1326);
nand U1268 (N_1268,In_439,In_161);
nor U1269 (N_1269,In_718,In_1373);
xnor U1270 (N_1270,In_225,In_978);
xor U1271 (N_1271,In_1044,In_21);
nor U1272 (N_1272,In_580,In_747);
and U1273 (N_1273,In_322,In_1305);
xor U1274 (N_1274,In_851,In_1236);
or U1275 (N_1275,In_468,In_358);
and U1276 (N_1276,In_84,In_522);
and U1277 (N_1277,In_725,In_291);
or U1278 (N_1278,In_1031,In_1351);
or U1279 (N_1279,In_354,In_815);
xor U1280 (N_1280,In_870,In_660);
or U1281 (N_1281,In_858,In_96);
and U1282 (N_1282,In_217,In_526);
nand U1283 (N_1283,In_94,In_1143);
nor U1284 (N_1284,In_1349,In_547);
nor U1285 (N_1285,In_1388,In_13);
xnor U1286 (N_1286,In_628,In_415);
xnor U1287 (N_1287,In_874,In_605);
xnor U1288 (N_1288,In_586,In_302);
or U1289 (N_1289,In_1193,In_1157);
nand U1290 (N_1290,In_711,In_529);
nand U1291 (N_1291,In_1381,In_872);
nand U1292 (N_1292,In_1000,In_269);
or U1293 (N_1293,In_1496,In_1414);
and U1294 (N_1294,In_290,In_166);
xnor U1295 (N_1295,In_509,In_725);
and U1296 (N_1296,In_889,In_1402);
and U1297 (N_1297,In_335,In_697);
and U1298 (N_1298,In_554,In_418);
and U1299 (N_1299,In_529,In_574);
and U1300 (N_1300,In_241,In_839);
or U1301 (N_1301,In_503,In_742);
xor U1302 (N_1302,In_923,In_1390);
or U1303 (N_1303,In_1257,In_280);
or U1304 (N_1304,In_1489,In_1171);
or U1305 (N_1305,In_1257,In_1497);
nand U1306 (N_1306,In_638,In_530);
xnor U1307 (N_1307,In_760,In_840);
nor U1308 (N_1308,In_1095,In_623);
nor U1309 (N_1309,In_309,In_980);
nand U1310 (N_1310,In_173,In_1077);
nor U1311 (N_1311,In_197,In_1497);
or U1312 (N_1312,In_1217,In_619);
or U1313 (N_1313,In_309,In_319);
and U1314 (N_1314,In_1176,In_463);
nand U1315 (N_1315,In_349,In_398);
nand U1316 (N_1316,In_748,In_1200);
nand U1317 (N_1317,In_1232,In_1479);
nand U1318 (N_1318,In_220,In_998);
xnor U1319 (N_1319,In_1414,In_64);
xnor U1320 (N_1320,In_1259,In_781);
and U1321 (N_1321,In_1363,In_1007);
nor U1322 (N_1322,In_687,In_566);
and U1323 (N_1323,In_1353,In_825);
nand U1324 (N_1324,In_646,In_141);
and U1325 (N_1325,In_275,In_1400);
xor U1326 (N_1326,In_1340,In_1333);
xor U1327 (N_1327,In_588,In_758);
and U1328 (N_1328,In_1224,In_180);
xnor U1329 (N_1329,In_1249,In_730);
and U1330 (N_1330,In_454,In_593);
or U1331 (N_1331,In_457,In_1484);
xor U1332 (N_1332,In_381,In_658);
nor U1333 (N_1333,In_100,In_1035);
nand U1334 (N_1334,In_202,In_1475);
xor U1335 (N_1335,In_1363,In_683);
nand U1336 (N_1336,In_292,In_324);
nor U1337 (N_1337,In_236,In_1371);
xnor U1338 (N_1338,In_2,In_723);
or U1339 (N_1339,In_127,In_10);
xor U1340 (N_1340,In_327,In_1045);
or U1341 (N_1341,In_1246,In_978);
xor U1342 (N_1342,In_1077,In_1263);
or U1343 (N_1343,In_379,In_526);
or U1344 (N_1344,In_1383,In_334);
nand U1345 (N_1345,In_141,In_1425);
and U1346 (N_1346,In_724,In_341);
and U1347 (N_1347,In_49,In_1275);
or U1348 (N_1348,In_415,In_435);
xnor U1349 (N_1349,In_1231,In_1191);
and U1350 (N_1350,In_218,In_469);
and U1351 (N_1351,In_677,In_482);
and U1352 (N_1352,In_1373,In_1258);
and U1353 (N_1353,In_93,In_903);
nand U1354 (N_1354,In_485,In_1058);
and U1355 (N_1355,In_910,In_892);
nor U1356 (N_1356,In_284,In_986);
or U1357 (N_1357,In_954,In_563);
xor U1358 (N_1358,In_415,In_266);
nand U1359 (N_1359,In_106,In_774);
nand U1360 (N_1360,In_453,In_1350);
nor U1361 (N_1361,In_860,In_1333);
or U1362 (N_1362,In_1055,In_1343);
or U1363 (N_1363,In_340,In_1022);
nor U1364 (N_1364,In_976,In_224);
nand U1365 (N_1365,In_1117,In_1086);
nand U1366 (N_1366,In_185,In_523);
and U1367 (N_1367,In_624,In_334);
nor U1368 (N_1368,In_693,In_40);
xnor U1369 (N_1369,In_1286,In_1475);
nand U1370 (N_1370,In_1104,In_1442);
or U1371 (N_1371,In_963,In_1398);
nor U1372 (N_1372,In_452,In_206);
xnor U1373 (N_1373,In_829,In_754);
nand U1374 (N_1374,In_1163,In_1248);
nand U1375 (N_1375,In_227,In_207);
or U1376 (N_1376,In_1121,In_1303);
nand U1377 (N_1377,In_494,In_1250);
nand U1378 (N_1378,In_1298,In_1466);
and U1379 (N_1379,In_825,In_1412);
nand U1380 (N_1380,In_1409,In_839);
or U1381 (N_1381,In_531,In_933);
xor U1382 (N_1382,In_1107,In_118);
xnor U1383 (N_1383,In_72,In_990);
and U1384 (N_1384,In_1209,In_980);
nor U1385 (N_1385,In_807,In_187);
or U1386 (N_1386,In_672,In_285);
and U1387 (N_1387,In_873,In_1351);
nand U1388 (N_1388,In_913,In_100);
and U1389 (N_1389,In_1033,In_54);
and U1390 (N_1390,In_430,In_730);
nor U1391 (N_1391,In_1203,In_649);
or U1392 (N_1392,In_196,In_775);
xnor U1393 (N_1393,In_659,In_253);
nand U1394 (N_1394,In_161,In_1117);
nand U1395 (N_1395,In_974,In_458);
nor U1396 (N_1396,In_1296,In_547);
nor U1397 (N_1397,In_1074,In_754);
nand U1398 (N_1398,In_336,In_830);
nor U1399 (N_1399,In_685,In_221);
nand U1400 (N_1400,In_19,In_1286);
or U1401 (N_1401,In_242,In_1412);
and U1402 (N_1402,In_123,In_727);
nor U1403 (N_1403,In_1234,In_1435);
nor U1404 (N_1404,In_105,In_833);
nor U1405 (N_1405,In_39,In_928);
xnor U1406 (N_1406,In_1161,In_1072);
and U1407 (N_1407,In_1030,In_704);
xnor U1408 (N_1408,In_1351,In_1280);
nor U1409 (N_1409,In_75,In_439);
and U1410 (N_1410,In_818,In_1388);
and U1411 (N_1411,In_313,In_920);
nor U1412 (N_1412,In_723,In_141);
and U1413 (N_1413,In_327,In_1391);
and U1414 (N_1414,In_1207,In_287);
nor U1415 (N_1415,In_262,In_1268);
nand U1416 (N_1416,In_397,In_1082);
and U1417 (N_1417,In_785,In_598);
xnor U1418 (N_1418,In_584,In_1373);
nand U1419 (N_1419,In_895,In_696);
or U1420 (N_1420,In_334,In_812);
and U1421 (N_1421,In_645,In_1368);
nor U1422 (N_1422,In_955,In_1454);
or U1423 (N_1423,In_1131,In_1386);
nand U1424 (N_1424,In_444,In_1409);
xor U1425 (N_1425,In_954,In_1227);
or U1426 (N_1426,In_373,In_1418);
or U1427 (N_1427,In_343,In_1214);
nor U1428 (N_1428,In_237,In_954);
nand U1429 (N_1429,In_661,In_1082);
nand U1430 (N_1430,In_751,In_1263);
nor U1431 (N_1431,In_944,In_700);
nand U1432 (N_1432,In_309,In_1492);
and U1433 (N_1433,In_553,In_270);
nor U1434 (N_1434,In_83,In_1070);
nand U1435 (N_1435,In_420,In_25);
or U1436 (N_1436,In_520,In_1088);
nand U1437 (N_1437,In_1371,In_1433);
and U1438 (N_1438,In_15,In_148);
and U1439 (N_1439,In_1174,In_387);
xnor U1440 (N_1440,In_798,In_1287);
nand U1441 (N_1441,In_902,In_421);
xnor U1442 (N_1442,In_84,In_193);
nor U1443 (N_1443,In_670,In_570);
and U1444 (N_1444,In_640,In_715);
or U1445 (N_1445,In_1401,In_177);
or U1446 (N_1446,In_365,In_1134);
xor U1447 (N_1447,In_711,In_1478);
and U1448 (N_1448,In_484,In_21);
and U1449 (N_1449,In_112,In_1326);
and U1450 (N_1450,In_119,In_913);
and U1451 (N_1451,In_774,In_175);
and U1452 (N_1452,In_1338,In_1076);
nand U1453 (N_1453,In_1381,In_282);
or U1454 (N_1454,In_1454,In_642);
nand U1455 (N_1455,In_998,In_926);
or U1456 (N_1456,In_1149,In_867);
and U1457 (N_1457,In_1168,In_726);
or U1458 (N_1458,In_287,In_603);
nand U1459 (N_1459,In_22,In_440);
nand U1460 (N_1460,In_751,In_978);
nor U1461 (N_1461,In_128,In_1315);
and U1462 (N_1462,In_115,In_1447);
xor U1463 (N_1463,In_555,In_626);
nor U1464 (N_1464,In_1313,In_788);
or U1465 (N_1465,In_441,In_1286);
nand U1466 (N_1466,In_221,In_302);
or U1467 (N_1467,In_446,In_300);
or U1468 (N_1468,In_375,In_1348);
nor U1469 (N_1469,In_136,In_236);
nand U1470 (N_1470,In_74,In_116);
nand U1471 (N_1471,In_303,In_1442);
nand U1472 (N_1472,In_1142,In_150);
or U1473 (N_1473,In_821,In_1170);
nor U1474 (N_1474,In_1245,In_1323);
xnor U1475 (N_1475,In_375,In_649);
nor U1476 (N_1476,In_1459,In_66);
nand U1477 (N_1477,In_181,In_1304);
nor U1478 (N_1478,In_1124,In_1119);
xnor U1479 (N_1479,In_449,In_188);
or U1480 (N_1480,In_1291,In_8);
nand U1481 (N_1481,In_830,In_280);
and U1482 (N_1482,In_965,In_1454);
and U1483 (N_1483,In_376,In_991);
nor U1484 (N_1484,In_299,In_867);
xor U1485 (N_1485,In_382,In_818);
nor U1486 (N_1486,In_73,In_167);
or U1487 (N_1487,In_154,In_957);
and U1488 (N_1488,In_414,In_1121);
or U1489 (N_1489,In_1226,In_1168);
nor U1490 (N_1490,In_1275,In_829);
xor U1491 (N_1491,In_1020,In_1243);
xor U1492 (N_1492,In_1415,In_342);
xor U1493 (N_1493,In_922,In_564);
nor U1494 (N_1494,In_1055,In_628);
nor U1495 (N_1495,In_1121,In_597);
nand U1496 (N_1496,In_973,In_537);
and U1497 (N_1497,In_1325,In_654);
or U1498 (N_1498,In_1351,In_1187);
or U1499 (N_1499,In_318,In_718);
nor U1500 (N_1500,In_1418,In_37);
and U1501 (N_1501,In_501,In_1217);
and U1502 (N_1502,In_366,In_87);
xor U1503 (N_1503,In_1314,In_219);
nor U1504 (N_1504,In_13,In_779);
and U1505 (N_1505,In_199,In_1385);
nor U1506 (N_1506,In_1202,In_1048);
nand U1507 (N_1507,In_709,In_168);
nand U1508 (N_1508,In_1475,In_990);
nor U1509 (N_1509,In_296,In_19);
or U1510 (N_1510,In_593,In_966);
nand U1511 (N_1511,In_874,In_1100);
nand U1512 (N_1512,In_448,In_626);
or U1513 (N_1513,In_419,In_595);
nand U1514 (N_1514,In_682,In_506);
nor U1515 (N_1515,In_1228,In_959);
nor U1516 (N_1516,In_192,In_996);
xor U1517 (N_1517,In_1092,In_365);
or U1518 (N_1518,In_181,In_477);
xnor U1519 (N_1519,In_612,In_357);
and U1520 (N_1520,In_713,In_398);
or U1521 (N_1521,In_310,In_17);
and U1522 (N_1522,In_284,In_1107);
nand U1523 (N_1523,In_1250,In_760);
nand U1524 (N_1524,In_1194,In_1376);
or U1525 (N_1525,In_707,In_762);
nor U1526 (N_1526,In_763,In_1377);
or U1527 (N_1527,In_453,In_953);
nand U1528 (N_1528,In_561,In_14);
nor U1529 (N_1529,In_1243,In_1212);
nand U1530 (N_1530,In_1181,In_396);
and U1531 (N_1531,In_74,In_419);
nor U1532 (N_1532,In_763,In_1234);
nand U1533 (N_1533,In_688,In_1318);
nand U1534 (N_1534,In_425,In_1321);
and U1535 (N_1535,In_200,In_1089);
nor U1536 (N_1536,In_537,In_822);
or U1537 (N_1537,In_1483,In_771);
nand U1538 (N_1538,In_1253,In_801);
xnor U1539 (N_1539,In_924,In_1074);
xnor U1540 (N_1540,In_555,In_1331);
nand U1541 (N_1541,In_1041,In_635);
or U1542 (N_1542,In_678,In_563);
nor U1543 (N_1543,In_901,In_1457);
nand U1544 (N_1544,In_600,In_216);
or U1545 (N_1545,In_900,In_1328);
or U1546 (N_1546,In_433,In_782);
nand U1547 (N_1547,In_1238,In_1051);
nor U1548 (N_1548,In_1282,In_1146);
or U1549 (N_1549,In_672,In_107);
xnor U1550 (N_1550,In_258,In_331);
or U1551 (N_1551,In_746,In_797);
nor U1552 (N_1552,In_1420,In_452);
and U1553 (N_1553,In_553,In_1221);
and U1554 (N_1554,In_35,In_750);
nand U1555 (N_1555,In_489,In_1223);
and U1556 (N_1556,In_1138,In_530);
nor U1557 (N_1557,In_149,In_499);
nor U1558 (N_1558,In_582,In_537);
and U1559 (N_1559,In_279,In_407);
nand U1560 (N_1560,In_700,In_51);
nand U1561 (N_1561,In_235,In_1067);
or U1562 (N_1562,In_418,In_47);
and U1563 (N_1563,In_55,In_937);
nand U1564 (N_1564,In_289,In_398);
xnor U1565 (N_1565,In_209,In_1473);
or U1566 (N_1566,In_184,In_185);
nand U1567 (N_1567,In_688,In_910);
nand U1568 (N_1568,In_857,In_667);
or U1569 (N_1569,In_581,In_550);
or U1570 (N_1570,In_611,In_209);
nor U1571 (N_1571,In_334,In_1398);
nor U1572 (N_1572,In_1184,In_199);
nand U1573 (N_1573,In_521,In_1031);
and U1574 (N_1574,In_226,In_1493);
nand U1575 (N_1575,In_1037,In_240);
or U1576 (N_1576,In_978,In_916);
nand U1577 (N_1577,In_2,In_27);
and U1578 (N_1578,In_702,In_548);
or U1579 (N_1579,In_325,In_186);
xnor U1580 (N_1580,In_428,In_708);
nand U1581 (N_1581,In_310,In_902);
nor U1582 (N_1582,In_753,In_191);
or U1583 (N_1583,In_1447,In_166);
or U1584 (N_1584,In_323,In_1266);
nor U1585 (N_1585,In_411,In_213);
xnor U1586 (N_1586,In_757,In_408);
nand U1587 (N_1587,In_561,In_952);
nor U1588 (N_1588,In_296,In_793);
nand U1589 (N_1589,In_6,In_758);
or U1590 (N_1590,In_1289,In_1409);
nand U1591 (N_1591,In_1446,In_1018);
nand U1592 (N_1592,In_1276,In_182);
and U1593 (N_1593,In_887,In_820);
nor U1594 (N_1594,In_373,In_437);
nand U1595 (N_1595,In_505,In_1009);
nor U1596 (N_1596,In_783,In_1228);
xnor U1597 (N_1597,In_1242,In_1186);
nand U1598 (N_1598,In_1046,In_1055);
and U1599 (N_1599,In_416,In_809);
and U1600 (N_1600,In_943,In_475);
and U1601 (N_1601,In_197,In_12);
xor U1602 (N_1602,In_1098,In_45);
and U1603 (N_1603,In_1104,In_853);
or U1604 (N_1604,In_597,In_256);
nor U1605 (N_1605,In_858,In_725);
or U1606 (N_1606,In_259,In_944);
nor U1607 (N_1607,In_247,In_1451);
or U1608 (N_1608,In_1240,In_454);
or U1609 (N_1609,In_1379,In_662);
nand U1610 (N_1610,In_1215,In_738);
nand U1611 (N_1611,In_1413,In_820);
nand U1612 (N_1612,In_559,In_936);
xnor U1613 (N_1613,In_1123,In_403);
xor U1614 (N_1614,In_839,In_421);
or U1615 (N_1615,In_630,In_881);
nand U1616 (N_1616,In_1208,In_524);
xor U1617 (N_1617,In_167,In_377);
or U1618 (N_1618,In_593,In_101);
or U1619 (N_1619,In_1200,In_566);
nor U1620 (N_1620,In_507,In_132);
nand U1621 (N_1621,In_952,In_641);
or U1622 (N_1622,In_369,In_42);
or U1623 (N_1623,In_630,In_489);
or U1624 (N_1624,In_855,In_1078);
nor U1625 (N_1625,In_711,In_321);
nand U1626 (N_1626,In_1475,In_1091);
and U1627 (N_1627,In_690,In_1367);
nor U1628 (N_1628,In_19,In_944);
xnor U1629 (N_1629,In_669,In_300);
nor U1630 (N_1630,In_233,In_1072);
nand U1631 (N_1631,In_844,In_81);
and U1632 (N_1632,In_176,In_1301);
xnor U1633 (N_1633,In_573,In_1461);
nand U1634 (N_1634,In_1497,In_467);
nand U1635 (N_1635,In_375,In_885);
and U1636 (N_1636,In_647,In_622);
xnor U1637 (N_1637,In_1201,In_670);
and U1638 (N_1638,In_733,In_999);
or U1639 (N_1639,In_85,In_1317);
xor U1640 (N_1640,In_1317,In_372);
nand U1641 (N_1641,In_942,In_351);
or U1642 (N_1642,In_698,In_1105);
xnor U1643 (N_1643,In_593,In_779);
nor U1644 (N_1644,In_1285,In_284);
and U1645 (N_1645,In_432,In_561);
xnor U1646 (N_1646,In_1157,In_406);
nor U1647 (N_1647,In_5,In_649);
xor U1648 (N_1648,In_303,In_566);
xor U1649 (N_1649,In_1463,In_144);
nand U1650 (N_1650,In_613,In_1308);
nor U1651 (N_1651,In_822,In_317);
xnor U1652 (N_1652,In_1316,In_232);
nand U1653 (N_1653,In_1213,In_1018);
nor U1654 (N_1654,In_188,In_1420);
xnor U1655 (N_1655,In_1172,In_1342);
xor U1656 (N_1656,In_1065,In_1153);
or U1657 (N_1657,In_1010,In_546);
nor U1658 (N_1658,In_882,In_1235);
xnor U1659 (N_1659,In_1429,In_1354);
nand U1660 (N_1660,In_931,In_510);
xor U1661 (N_1661,In_1185,In_546);
or U1662 (N_1662,In_662,In_581);
xnor U1663 (N_1663,In_241,In_534);
xnor U1664 (N_1664,In_1227,In_84);
xnor U1665 (N_1665,In_1439,In_30);
nand U1666 (N_1666,In_459,In_375);
nand U1667 (N_1667,In_469,In_1113);
xnor U1668 (N_1668,In_204,In_1491);
nand U1669 (N_1669,In_1286,In_333);
or U1670 (N_1670,In_607,In_984);
nor U1671 (N_1671,In_388,In_693);
nor U1672 (N_1672,In_1105,In_514);
or U1673 (N_1673,In_1043,In_324);
and U1674 (N_1674,In_922,In_850);
nor U1675 (N_1675,In_862,In_105);
and U1676 (N_1676,In_158,In_643);
or U1677 (N_1677,In_1426,In_176);
and U1678 (N_1678,In_1307,In_812);
and U1679 (N_1679,In_57,In_642);
nand U1680 (N_1680,In_297,In_554);
nand U1681 (N_1681,In_367,In_257);
and U1682 (N_1682,In_297,In_125);
and U1683 (N_1683,In_58,In_767);
or U1684 (N_1684,In_453,In_648);
nor U1685 (N_1685,In_13,In_1013);
xnor U1686 (N_1686,In_1404,In_1266);
or U1687 (N_1687,In_741,In_947);
nand U1688 (N_1688,In_92,In_1383);
or U1689 (N_1689,In_578,In_960);
xor U1690 (N_1690,In_163,In_437);
nor U1691 (N_1691,In_1061,In_639);
nor U1692 (N_1692,In_1368,In_721);
or U1693 (N_1693,In_1436,In_1294);
nor U1694 (N_1694,In_1254,In_420);
or U1695 (N_1695,In_677,In_455);
or U1696 (N_1696,In_128,In_578);
nor U1697 (N_1697,In_369,In_1324);
xnor U1698 (N_1698,In_69,In_1036);
or U1699 (N_1699,In_1128,In_997);
nor U1700 (N_1700,In_732,In_471);
and U1701 (N_1701,In_605,In_1127);
nand U1702 (N_1702,In_150,In_67);
nand U1703 (N_1703,In_64,In_435);
or U1704 (N_1704,In_1210,In_46);
nand U1705 (N_1705,In_1228,In_1219);
xor U1706 (N_1706,In_721,In_306);
nand U1707 (N_1707,In_1034,In_975);
and U1708 (N_1708,In_512,In_503);
xnor U1709 (N_1709,In_724,In_243);
nand U1710 (N_1710,In_520,In_83);
xnor U1711 (N_1711,In_1167,In_574);
xnor U1712 (N_1712,In_126,In_1295);
and U1713 (N_1713,In_1184,In_48);
and U1714 (N_1714,In_1493,In_1165);
or U1715 (N_1715,In_1264,In_536);
nand U1716 (N_1716,In_473,In_860);
and U1717 (N_1717,In_136,In_798);
nand U1718 (N_1718,In_1038,In_777);
nor U1719 (N_1719,In_1041,In_1221);
nor U1720 (N_1720,In_649,In_1486);
and U1721 (N_1721,In_645,In_1233);
and U1722 (N_1722,In_1327,In_108);
nand U1723 (N_1723,In_1278,In_1420);
and U1724 (N_1724,In_1147,In_1145);
nor U1725 (N_1725,In_358,In_39);
or U1726 (N_1726,In_311,In_1078);
nor U1727 (N_1727,In_1257,In_457);
nor U1728 (N_1728,In_600,In_582);
nor U1729 (N_1729,In_1336,In_646);
and U1730 (N_1730,In_762,In_1363);
nand U1731 (N_1731,In_523,In_1240);
xor U1732 (N_1732,In_273,In_329);
and U1733 (N_1733,In_1459,In_1129);
xnor U1734 (N_1734,In_1148,In_531);
xnor U1735 (N_1735,In_1073,In_1167);
or U1736 (N_1736,In_188,In_95);
nand U1737 (N_1737,In_1448,In_125);
xor U1738 (N_1738,In_376,In_943);
nor U1739 (N_1739,In_329,In_588);
nand U1740 (N_1740,In_291,In_997);
nor U1741 (N_1741,In_309,In_67);
or U1742 (N_1742,In_601,In_1236);
nand U1743 (N_1743,In_1240,In_637);
and U1744 (N_1744,In_1331,In_965);
nand U1745 (N_1745,In_174,In_1473);
xnor U1746 (N_1746,In_476,In_758);
and U1747 (N_1747,In_1209,In_135);
xor U1748 (N_1748,In_790,In_1084);
nand U1749 (N_1749,In_572,In_407);
or U1750 (N_1750,In_187,In_1015);
or U1751 (N_1751,In_182,In_87);
or U1752 (N_1752,In_1001,In_838);
nor U1753 (N_1753,In_866,In_711);
or U1754 (N_1754,In_909,In_620);
and U1755 (N_1755,In_91,In_453);
nor U1756 (N_1756,In_1244,In_920);
xnor U1757 (N_1757,In_826,In_403);
xor U1758 (N_1758,In_708,In_541);
nand U1759 (N_1759,In_347,In_68);
or U1760 (N_1760,In_921,In_297);
nand U1761 (N_1761,In_823,In_452);
nand U1762 (N_1762,In_286,In_122);
xnor U1763 (N_1763,In_1043,In_764);
or U1764 (N_1764,In_1411,In_941);
nand U1765 (N_1765,In_817,In_439);
nor U1766 (N_1766,In_304,In_594);
and U1767 (N_1767,In_1066,In_453);
xnor U1768 (N_1768,In_5,In_341);
and U1769 (N_1769,In_1119,In_1489);
xnor U1770 (N_1770,In_1054,In_1123);
xnor U1771 (N_1771,In_1407,In_1448);
nor U1772 (N_1772,In_750,In_1421);
and U1773 (N_1773,In_240,In_851);
xor U1774 (N_1774,In_1336,In_330);
xor U1775 (N_1775,In_1475,In_319);
or U1776 (N_1776,In_363,In_468);
or U1777 (N_1777,In_1109,In_1116);
and U1778 (N_1778,In_398,In_485);
nor U1779 (N_1779,In_1098,In_973);
and U1780 (N_1780,In_663,In_34);
nand U1781 (N_1781,In_1129,In_780);
and U1782 (N_1782,In_363,In_857);
xnor U1783 (N_1783,In_1189,In_624);
xor U1784 (N_1784,In_1378,In_523);
nor U1785 (N_1785,In_82,In_844);
and U1786 (N_1786,In_551,In_1369);
xor U1787 (N_1787,In_534,In_22);
nand U1788 (N_1788,In_390,In_1484);
xor U1789 (N_1789,In_44,In_1145);
xnor U1790 (N_1790,In_592,In_61);
nor U1791 (N_1791,In_325,In_10);
nand U1792 (N_1792,In_666,In_66);
xnor U1793 (N_1793,In_653,In_128);
and U1794 (N_1794,In_698,In_1331);
and U1795 (N_1795,In_1189,In_1296);
nor U1796 (N_1796,In_1101,In_1268);
or U1797 (N_1797,In_1135,In_287);
xor U1798 (N_1798,In_32,In_204);
or U1799 (N_1799,In_401,In_247);
and U1800 (N_1800,In_721,In_496);
nor U1801 (N_1801,In_748,In_723);
and U1802 (N_1802,In_1244,In_463);
nand U1803 (N_1803,In_968,In_841);
nand U1804 (N_1804,In_484,In_959);
nor U1805 (N_1805,In_1019,In_1421);
or U1806 (N_1806,In_1253,In_1059);
or U1807 (N_1807,In_1065,In_1096);
and U1808 (N_1808,In_1305,In_178);
nor U1809 (N_1809,In_1192,In_1169);
nand U1810 (N_1810,In_112,In_716);
nor U1811 (N_1811,In_668,In_1095);
or U1812 (N_1812,In_1397,In_1239);
and U1813 (N_1813,In_286,In_170);
nor U1814 (N_1814,In_548,In_1289);
and U1815 (N_1815,In_517,In_109);
or U1816 (N_1816,In_1345,In_1426);
and U1817 (N_1817,In_778,In_1295);
or U1818 (N_1818,In_1060,In_804);
nand U1819 (N_1819,In_561,In_902);
or U1820 (N_1820,In_811,In_71);
nor U1821 (N_1821,In_972,In_1223);
and U1822 (N_1822,In_247,In_802);
xor U1823 (N_1823,In_562,In_1093);
and U1824 (N_1824,In_1080,In_36);
and U1825 (N_1825,In_335,In_962);
and U1826 (N_1826,In_1491,In_697);
nor U1827 (N_1827,In_480,In_687);
or U1828 (N_1828,In_682,In_895);
nor U1829 (N_1829,In_41,In_662);
and U1830 (N_1830,In_1047,In_1111);
nor U1831 (N_1831,In_906,In_360);
nand U1832 (N_1832,In_30,In_892);
nor U1833 (N_1833,In_1261,In_1144);
nand U1834 (N_1834,In_642,In_554);
nor U1835 (N_1835,In_1421,In_152);
and U1836 (N_1836,In_1278,In_199);
nand U1837 (N_1837,In_797,In_127);
or U1838 (N_1838,In_580,In_162);
or U1839 (N_1839,In_1126,In_590);
and U1840 (N_1840,In_1274,In_741);
or U1841 (N_1841,In_1216,In_680);
nand U1842 (N_1842,In_1071,In_1410);
and U1843 (N_1843,In_1337,In_774);
nand U1844 (N_1844,In_993,In_1408);
or U1845 (N_1845,In_56,In_48);
or U1846 (N_1846,In_1289,In_1149);
xor U1847 (N_1847,In_31,In_1477);
and U1848 (N_1848,In_1262,In_1175);
nor U1849 (N_1849,In_511,In_497);
nor U1850 (N_1850,In_979,In_127);
nand U1851 (N_1851,In_568,In_1135);
xor U1852 (N_1852,In_1472,In_524);
nor U1853 (N_1853,In_634,In_859);
nor U1854 (N_1854,In_668,In_1189);
nand U1855 (N_1855,In_140,In_1278);
nor U1856 (N_1856,In_50,In_773);
or U1857 (N_1857,In_127,In_219);
nand U1858 (N_1858,In_811,In_1086);
nor U1859 (N_1859,In_427,In_245);
and U1860 (N_1860,In_917,In_36);
or U1861 (N_1861,In_578,In_1166);
and U1862 (N_1862,In_140,In_756);
xor U1863 (N_1863,In_135,In_858);
or U1864 (N_1864,In_1170,In_725);
or U1865 (N_1865,In_444,In_89);
or U1866 (N_1866,In_207,In_1030);
nor U1867 (N_1867,In_1273,In_1026);
nand U1868 (N_1868,In_531,In_151);
nor U1869 (N_1869,In_755,In_900);
and U1870 (N_1870,In_778,In_378);
and U1871 (N_1871,In_838,In_953);
nor U1872 (N_1872,In_309,In_141);
and U1873 (N_1873,In_1438,In_287);
and U1874 (N_1874,In_328,In_935);
xnor U1875 (N_1875,In_58,In_1225);
xor U1876 (N_1876,In_1152,In_1356);
and U1877 (N_1877,In_438,In_205);
and U1878 (N_1878,In_189,In_945);
or U1879 (N_1879,In_292,In_25);
or U1880 (N_1880,In_748,In_279);
nor U1881 (N_1881,In_1102,In_499);
or U1882 (N_1882,In_1354,In_1441);
xor U1883 (N_1883,In_1318,In_931);
xnor U1884 (N_1884,In_1053,In_641);
or U1885 (N_1885,In_318,In_1485);
and U1886 (N_1886,In_613,In_1405);
and U1887 (N_1887,In_1399,In_1201);
nand U1888 (N_1888,In_284,In_1168);
or U1889 (N_1889,In_1102,In_201);
nor U1890 (N_1890,In_1307,In_1193);
or U1891 (N_1891,In_228,In_761);
or U1892 (N_1892,In_1011,In_21);
nand U1893 (N_1893,In_364,In_564);
xnor U1894 (N_1894,In_1410,In_1188);
xnor U1895 (N_1895,In_1496,In_237);
and U1896 (N_1896,In_1309,In_32);
or U1897 (N_1897,In_598,In_742);
nor U1898 (N_1898,In_479,In_795);
or U1899 (N_1899,In_25,In_680);
or U1900 (N_1900,In_807,In_610);
and U1901 (N_1901,In_246,In_847);
or U1902 (N_1902,In_934,In_326);
nor U1903 (N_1903,In_1309,In_1040);
nor U1904 (N_1904,In_276,In_1471);
or U1905 (N_1905,In_1401,In_150);
and U1906 (N_1906,In_980,In_1257);
nand U1907 (N_1907,In_950,In_1301);
and U1908 (N_1908,In_374,In_198);
nor U1909 (N_1909,In_665,In_107);
nand U1910 (N_1910,In_1379,In_453);
xnor U1911 (N_1911,In_1298,In_1013);
xor U1912 (N_1912,In_284,In_548);
nor U1913 (N_1913,In_108,In_900);
xnor U1914 (N_1914,In_336,In_275);
xor U1915 (N_1915,In_1367,In_350);
nand U1916 (N_1916,In_196,In_120);
and U1917 (N_1917,In_57,In_167);
xnor U1918 (N_1918,In_791,In_1467);
nand U1919 (N_1919,In_1453,In_302);
or U1920 (N_1920,In_1350,In_1485);
nor U1921 (N_1921,In_513,In_168);
nor U1922 (N_1922,In_243,In_902);
xnor U1923 (N_1923,In_49,In_847);
nand U1924 (N_1924,In_369,In_515);
or U1925 (N_1925,In_735,In_643);
or U1926 (N_1926,In_1406,In_788);
or U1927 (N_1927,In_571,In_384);
nor U1928 (N_1928,In_1130,In_1448);
nand U1929 (N_1929,In_723,In_429);
nand U1930 (N_1930,In_414,In_1212);
nor U1931 (N_1931,In_624,In_1081);
xnor U1932 (N_1932,In_766,In_974);
nor U1933 (N_1933,In_390,In_693);
or U1934 (N_1934,In_1107,In_1022);
or U1935 (N_1935,In_1366,In_1217);
and U1936 (N_1936,In_522,In_58);
and U1937 (N_1937,In_665,In_756);
and U1938 (N_1938,In_679,In_1146);
nor U1939 (N_1939,In_647,In_621);
or U1940 (N_1940,In_1013,In_938);
xor U1941 (N_1941,In_811,In_1056);
and U1942 (N_1942,In_394,In_929);
and U1943 (N_1943,In_192,In_1427);
and U1944 (N_1944,In_441,In_1133);
xor U1945 (N_1945,In_266,In_158);
nand U1946 (N_1946,In_1140,In_117);
nor U1947 (N_1947,In_627,In_932);
nor U1948 (N_1948,In_825,In_538);
nor U1949 (N_1949,In_421,In_1335);
or U1950 (N_1950,In_421,In_959);
and U1951 (N_1951,In_192,In_91);
nand U1952 (N_1952,In_243,In_987);
xnor U1953 (N_1953,In_1312,In_1092);
nor U1954 (N_1954,In_1455,In_63);
xor U1955 (N_1955,In_701,In_104);
nor U1956 (N_1956,In_900,In_474);
or U1957 (N_1957,In_1435,In_313);
and U1958 (N_1958,In_918,In_1174);
nor U1959 (N_1959,In_395,In_1477);
xor U1960 (N_1960,In_433,In_312);
nor U1961 (N_1961,In_873,In_745);
xor U1962 (N_1962,In_917,In_1358);
and U1963 (N_1963,In_1002,In_287);
nand U1964 (N_1964,In_1009,In_1408);
nor U1965 (N_1965,In_1467,In_570);
xnor U1966 (N_1966,In_527,In_410);
or U1967 (N_1967,In_19,In_124);
xor U1968 (N_1968,In_678,In_56);
and U1969 (N_1969,In_701,In_201);
nand U1970 (N_1970,In_141,In_1419);
and U1971 (N_1971,In_762,In_358);
nor U1972 (N_1972,In_58,In_1021);
or U1973 (N_1973,In_1169,In_217);
nand U1974 (N_1974,In_1270,In_831);
xnor U1975 (N_1975,In_473,In_105);
xnor U1976 (N_1976,In_985,In_43);
or U1977 (N_1977,In_1226,In_1320);
or U1978 (N_1978,In_1458,In_407);
xnor U1979 (N_1979,In_1433,In_805);
or U1980 (N_1980,In_344,In_731);
and U1981 (N_1981,In_776,In_425);
nor U1982 (N_1982,In_891,In_1310);
and U1983 (N_1983,In_822,In_1284);
or U1984 (N_1984,In_776,In_90);
and U1985 (N_1985,In_964,In_770);
nor U1986 (N_1986,In_262,In_918);
and U1987 (N_1987,In_272,In_436);
xor U1988 (N_1988,In_779,In_1313);
nor U1989 (N_1989,In_825,In_332);
and U1990 (N_1990,In_395,In_1098);
and U1991 (N_1991,In_1281,In_1080);
xnor U1992 (N_1992,In_1313,In_1408);
nand U1993 (N_1993,In_1334,In_1057);
nor U1994 (N_1994,In_238,In_921);
and U1995 (N_1995,In_1391,In_526);
nand U1996 (N_1996,In_1262,In_1365);
or U1997 (N_1997,In_1336,In_831);
nor U1998 (N_1998,In_9,In_81);
xnor U1999 (N_1999,In_807,In_804);
nand U2000 (N_2000,In_527,In_621);
and U2001 (N_2001,In_616,In_394);
or U2002 (N_2002,In_720,In_1124);
nand U2003 (N_2003,In_1454,In_134);
and U2004 (N_2004,In_789,In_885);
xnor U2005 (N_2005,In_1206,In_899);
nor U2006 (N_2006,In_722,In_602);
or U2007 (N_2007,In_893,In_499);
or U2008 (N_2008,In_1169,In_1251);
and U2009 (N_2009,In_775,In_379);
xor U2010 (N_2010,In_413,In_509);
xor U2011 (N_2011,In_600,In_1412);
nand U2012 (N_2012,In_1445,In_1035);
nor U2013 (N_2013,In_1405,In_511);
and U2014 (N_2014,In_27,In_142);
nor U2015 (N_2015,In_864,In_930);
and U2016 (N_2016,In_1305,In_1457);
or U2017 (N_2017,In_441,In_1313);
nand U2018 (N_2018,In_1015,In_510);
nor U2019 (N_2019,In_1420,In_448);
nand U2020 (N_2020,In_1456,In_1495);
or U2021 (N_2021,In_157,In_1037);
nand U2022 (N_2022,In_105,In_1046);
and U2023 (N_2023,In_774,In_1037);
or U2024 (N_2024,In_389,In_445);
or U2025 (N_2025,In_1435,In_1439);
nor U2026 (N_2026,In_385,In_929);
and U2027 (N_2027,In_1113,In_286);
nand U2028 (N_2028,In_1248,In_539);
xor U2029 (N_2029,In_909,In_1204);
or U2030 (N_2030,In_1477,In_398);
nand U2031 (N_2031,In_1132,In_95);
nand U2032 (N_2032,In_272,In_370);
xor U2033 (N_2033,In_129,In_1421);
or U2034 (N_2034,In_827,In_984);
nor U2035 (N_2035,In_474,In_962);
nor U2036 (N_2036,In_505,In_608);
nand U2037 (N_2037,In_870,In_993);
xor U2038 (N_2038,In_983,In_268);
nand U2039 (N_2039,In_277,In_306);
xnor U2040 (N_2040,In_635,In_1156);
nand U2041 (N_2041,In_221,In_900);
and U2042 (N_2042,In_1195,In_852);
nand U2043 (N_2043,In_47,In_107);
nor U2044 (N_2044,In_1233,In_1218);
nand U2045 (N_2045,In_568,In_346);
xnor U2046 (N_2046,In_284,In_716);
nor U2047 (N_2047,In_1107,In_1117);
xnor U2048 (N_2048,In_92,In_1177);
nand U2049 (N_2049,In_219,In_1108);
xnor U2050 (N_2050,In_92,In_1037);
and U2051 (N_2051,In_955,In_747);
and U2052 (N_2052,In_785,In_1183);
xnor U2053 (N_2053,In_291,In_395);
nand U2054 (N_2054,In_1166,In_487);
or U2055 (N_2055,In_693,In_727);
xnor U2056 (N_2056,In_508,In_755);
or U2057 (N_2057,In_718,In_821);
nor U2058 (N_2058,In_1229,In_541);
and U2059 (N_2059,In_286,In_15);
and U2060 (N_2060,In_321,In_1381);
nand U2061 (N_2061,In_458,In_383);
nand U2062 (N_2062,In_887,In_1463);
nor U2063 (N_2063,In_1209,In_1084);
nor U2064 (N_2064,In_193,In_1253);
and U2065 (N_2065,In_612,In_538);
or U2066 (N_2066,In_759,In_423);
nand U2067 (N_2067,In_439,In_47);
and U2068 (N_2068,In_627,In_563);
nor U2069 (N_2069,In_862,In_258);
nand U2070 (N_2070,In_1333,In_794);
nor U2071 (N_2071,In_36,In_1465);
and U2072 (N_2072,In_285,In_384);
nand U2073 (N_2073,In_1018,In_803);
nand U2074 (N_2074,In_265,In_738);
and U2075 (N_2075,In_75,In_1118);
and U2076 (N_2076,In_1451,In_201);
and U2077 (N_2077,In_346,In_1338);
and U2078 (N_2078,In_276,In_879);
or U2079 (N_2079,In_1094,In_899);
xor U2080 (N_2080,In_1305,In_1194);
or U2081 (N_2081,In_3,In_1451);
or U2082 (N_2082,In_1273,In_25);
xor U2083 (N_2083,In_617,In_522);
or U2084 (N_2084,In_300,In_116);
and U2085 (N_2085,In_1240,In_1482);
nand U2086 (N_2086,In_528,In_523);
or U2087 (N_2087,In_783,In_8);
nor U2088 (N_2088,In_663,In_526);
and U2089 (N_2089,In_627,In_1279);
and U2090 (N_2090,In_1352,In_1484);
nor U2091 (N_2091,In_657,In_907);
nor U2092 (N_2092,In_698,In_430);
nand U2093 (N_2093,In_600,In_957);
nor U2094 (N_2094,In_850,In_1050);
nor U2095 (N_2095,In_398,In_361);
xor U2096 (N_2096,In_288,In_224);
or U2097 (N_2097,In_807,In_206);
xnor U2098 (N_2098,In_871,In_77);
and U2099 (N_2099,In_1420,In_145);
nor U2100 (N_2100,In_463,In_1236);
xor U2101 (N_2101,In_667,In_1253);
nand U2102 (N_2102,In_1201,In_401);
or U2103 (N_2103,In_931,In_1237);
xnor U2104 (N_2104,In_431,In_1475);
or U2105 (N_2105,In_476,In_607);
xnor U2106 (N_2106,In_1397,In_91);
nor U2107 (N_2107,In_912,In_1024);
and U2108 (N_2108,In_323,In_79);
nor U2109 (N_2109,In_1319,In_591);
xor U2110 (N_2110,In_796,In_135);
and U2111 (N_2111,In_1384,In_598);
xor U2112 (N_2112,In_1162,In_995);
nor U2113 (N_2113,In_1176,In_778);
or U2114 (N_2114,In_658,In_1304);
or U2115 (N_2115,In_1229,In_969);
xnor U2116 (N_2116,In_542,In_1295);
nand U2117 (N_2117,In_1443,In_592);
nor U2118 (N_2118,In_84,In_561);
nand U2119 (N_2119,In_1146,In_789);
nand U2120 (N_2120,In_860,In_374);
or U2121 (N_2121,In_1390,In_176);
nand U2122 (N_2122,In_168,In_1179);
nor U2123 (N_2123,In_1408,In_61);
nor U2124 (N_2124,In_443,In_960);
nor U2125 (N_2125,In_1236,In_444);
nor U2126 (N_2126,In_641,In_1455);
or U2127 (N_2127,In_213,In_282);
or U2128 (N_2128,In_1101,In_720);
xnor U2129 (N_2129,In_1396,In_1180);
nor U2130 (N_2130,In_80,In_1213);
nand U2131 (N_2131,In_355,In_652);
nand U2132 (N_2132,In_262,In_920);
nor U2133 (N_2133,In_1184,In_429);
or U2134 (N_2134,In_111,In_892);
xnor U2135 (N_2135,In_1038,In_614);
or U2136 (N_2136,In_1216,In_264);
nor U2137 (N_2137,In_121,In_853);
xor U2138 (N_2138,In_1079,In_1278);
nand U2139 (N_2139,In_1286,In_856);
xor U2140 (N_2140,In_1435,In_1091);
nand U2141 (N_2141,In_178,In_992);
nor U2142 (N_2142,In_1229,In_1475);
xnor U2143 (N_2143,In_311,In_1089);
and U2144 (N_2144,In_1006,In_354);
xnor U2145 (N_2145,In_910,In_989);
and U2146 (N_2146,In_934,In_1372);
nand U2147 (N_2147,In_77,In_535);
nand U2148 (N_2148,In_581,In_190);
or U2149 (N_2149,In_418,In_336);
nand U2150 (N_2150,In_760,In_583);
or U2151 (N_2151,In_1260,In_1031);
xnor U2152 (N_2152,In_888,In_1388);
xnor U2153 (N_2153,In_1410,In_751);
or U2154 (N_2154,In_984,In_184);
nor U2155 (N_2155,In_798,In_1433);
or U2156 (N_2156,In_1080,In_140);
and U2157 (N_2157,In_268,In_1078);
and U2158 (N_2158,In_287,In_854);
nor U2159 (N_2159,In_1454,In_1290);
and U2160 (N_2160,In_436,In_1248);
xor U2161 (N_2161,In_328,In_832);
and U2162 (N_2162,In_221,In_91);
nand U2163 (N_2163,In_1092,In_816);
xnor U2164 (N_2164,In_652,In_356);
and U2165 (N_2165,In_29,In_515);
or U2166 (N_2166,In_429,In_385);
nand U2167 (N_2167,In_456,In_177);
nand U2168 (N_2168,In_359,In_1392);
nor U2169 (N_2169,In_421,In_417);
or U2170 (N_2170,In_959,In_365);
and U2171 (N_2171,In_374,In_1290);
and U2172 (N_2172,In_0,In_82);
and U2173 (N_2173,In_1333,In_91);
and U2174 (N_2174,In_612,In_977);
xnor U2175 (N_2175,In_814,In_1232);
nand U2176 (N_2176,In_889,In_318);
or U2177 (N_2177,In_431,In_1006);
or U2178 (N_2178,In_383,In_179);
xor U2179 (N_2179,In_406,In_897);
and U2180 (N_2180,In_253,In_1167);
nor U2181 (N_2181,In_1068,In_1098);
and U2182 (N_2182,In_1433,In_683);
nor U2183 (N_2183,In_242,In_162);
xnor U2184 (N_2184,In_445,In_10);
or U2185 (N_2185,In_823,In_1006);
and U2186 (N_2186,In_1215,In_906);
and U2187 (N_2187,In_555,In_907);
nand U2188 (N_2188,In_255,In_1424);
and U2189 (N_2189,In_500,In_928);
xnor U2190 (N_2190,In_1237,In_969);
xor U2191 (N_2191,In_648,In_658);
or U2192 (N_2192,In_271,In_152);
and U2193 (N_2193,In_20,In_560);
nand U2194 (N_2194,In_953,In_302);
xnor U2195 (N_2195,In_843,In_371);
and U2196 (N_2196,In_1324,In_374);
or U2197 (N_2197,In_111,In_951);
or U2198 (N_2198,In_1112,In_737);
and U2199 (N_2199,In_459,In_1132);
nor U2200 (N_2200,In_514,In_19);
nand U2201 (N_2201,In_748,In_173);
or U2202 (N_2202,In_1220,In_908);
or U2203 (N_2203,In_911,In_1384);
or U2204 (N_2204,In_1448,In_476);
nor U2205 (N_2205,In_812,In_1303);
nand U2206 (N_2206,In_1236,In_777);
nand U2207 (N_2207,In_430,In_806);
xnor U2208 (N_2208,In_213,In_1076);
xor U2209 (N_2209,In_902,In_1037);
or U2210 (N_2210,In_763,In_1068);
xnor U2211 (N_2211,In_173,In_1320);
nand U2212 (N_2212,In_138,In_496);
nand U2213 (N_2213,In_630,In_1299);
nor U2214 (N_2214,In_1421,In_1415);
or U2215 (N_2215,In_1485,In_1058);
xnor U2216 (N_2216,In_628,In_1286);
and U2217 (N_2217,In_681,In_1429);
nor U2218 (N_2218,In_0,In_141);
nor U2219 (N_2219,In_1314,In_177);
and U2220 (N_2220,In_1318,In_902);
and U2221 (N_2221,In_643,In_1017);
or U2222 (N_2222,In_636,In_238);
or U2223 (N_2223,In_349,In_546);
and U2224 (N_2224,In_598,In_164);
nor U2225 (N_2225,In_949,In_272);
and U2226 (N_2226,In_852,In_49);
nand U2227 (N_2227,In_414,In_332);
nor U2228 (N_2228,In_378,In_197);
nor U2229 (N_2229,In_1032,In_1484);
nand U2230 (N_2230,In_30,In_455);
nor U2231 (N_2231,In_1416,In_787);
xnor U2232 (N_2232,In_429,In_1255);
nand U2233 (N_2233,In_325,In_287);
xor U2234 (N_2234,In_1400,In_1231);
or U2235 (N_2235,In_571,In_255);
or U2236 (N_2236,In_963,In_250);
nand U2237 (N_2237,In_207,In_590);
nand U2238 (N_2238,In_887,In_383);
nand U2239 (N_2239,In_22,In_806);
and U2240 (N_2240,In_61,In_1477);
xnor U2241 (N_2241,In_1100,In_350);
or U2242 (N_2242,In_435,In_183);
nand U2243 (N_2243,In_109,In_802);
nand U2244 (N_2244,In_455,In_988);
nand U2245 (N_2245,In_828,In_1071);
xnor U2246 (N_2246,In_45,In_1121);
and U2247 (N_2247,In_817,In_1116);
nand U2248 (N_2248,In_170,In_1076);
nor U2249 (N_2249,In_911,In_99);
and U2250 (N_2250,In_212,In_130);
nor U2251 (N_2251,In_437,In_376);
nand U2252 (N_2252,In_905,In_1407);
nor U2253 (N_2253,In_1469,In_651);
or U2254 (N_2254,In_399,In_246);
or U2255 (N_2255,In_973,In_829);
nand U2256 (N_2256,In_531,In_1105);
nand U2257 (N_2257,In_516,In_1391);
nand U2258 (N_2258,In_608,In_103);
or U2259 (N_2259,In_226,In_866);
and U2260 (N_2260,In_189,In_1146);
or U2261 (N_2261,In_740,In_343);
or U2262 (N_2262,In_223,In_619);
and U2263 (N_2263,In_232,In_1278);
or U2264 (N_2264,In_280,In_1140);
nor U2265 (N_2265,In_1006,In_1178);
or U2266 (N_2266,In_534,In_1119);
and U2267 (N_2267,In_553,In_1412);
nand U2268 (N_2268,In_1049,In_963);
or U2269 (N_2269,In_46,In_669);
and U2270 (N_2270,In_351,In_505);
or U2271 (N_2271,In_671,In_1131);
nor U2272 (N_2272,In_734,In_586);
xor U2273 (N_2273,In_1419,In_160);
or U2274 (N_2274,In_100,In_803);
nand U2275 (N_2275,In_352,In_1046);
xor U2276 (N_2276,In_1372,In_557);
and U2277 (N_2277,In_1052,In_85);
and U2278 (N_2278,In_466,In_443);
and U2279 (N_2279,In_489,In_268);
nand U2280 (N_2280,In_546,In_1275);
nand U2281 (N_2281,In_1241,In_841);
and U2282 (N_2282,In_276,In_17);
xnor U2283 (N_2283,In_119,In_1462);
nor U2284 (N_2284,In_912,In_611);
xnor U2285 (N_2285,In_1054,In_950);
xnor U2286 (N_2286,In_976,In_58);
and U2287 (N_2287,In_1031,In_542);
xnor U2288 (N_2288,In_5,In_1315);
nand U2289 (N_2289,In_555,In_4);
and U2290 (N_2290,In_230,In_1143);
and U2291 (N_2291,In_51,In_392);
or U2292 (N_2292,In_713,In_199);
or U2293 (N_2293,In_271,In_897);
and U2294 (N_2294,In_956,In_101);
xor U2295 (N_2295,In_1277,In_1041);
nor U2296 (N_2296,In_874,In_284);
nand U2297 (N_2297,In_83,In_183);
or U2298 (N_2298,In_787,In_411);
xor U2299 (N_2299,In_1008,In_1481);
nor U2300 (N_2300,In_497,In_389);
and U2301 (N_2301,In_493,In_1366);
or U2302 (N_2302,In_413,In_466);
nor U2303 (N_2303,In_793,In_1140);
xor U2304 (N_2304,In_34,In_689);
and U2305 (N_2305,In_36,In_894);
and U2306 (N_2306,In_1280,In_1385);
nand U2307 (N_2307,In_775,In_788);
nor U2308 (N_2308,In_1377,In_1348);
xor U2309 (N_2309,In_1290,In_119);
xor U2310 (N_2310,In_1253,In_777);
nand U2311 (N_2311,In_235,In_1188);
nor U2312 (N_2312,In_607,In_466);
and U2313 (N_2313,In_1398,In_81);
nor U2314 (N_2314,In_1324,In_400);
nor U2315 (N_2315,In_1392,In_797);
xnor U2316 (N_2316,In_1461,In_781);
xnor U2317 (N_2317,In_681,In_405);
nor U2318 (N_2318,In_569,In_492);
nor U2319 (N_2319,In_262,In_632);
xnor U2320 (N_2320,In_94,In_817);
nor U2321 (N_2321,In_931,In_168);
xnor U2322 (N_2322,In_453,In_612);
nor U2323 (N_2323,In_17,In_288);
and U2324 (N_2324,In_471,In_444);
nand U2325 (N_2325,In_788,In_1276);
or U2326 (N_2326,In_1264,In_1266);
nor U2327 (N_2327,In_189,In_403);
xor U2328 (N_2328,In_412,In_799);
nor U2329 (N_2329,In_1023,In_1231);
nand U2330 (N_2330,In_1123,In_770);
and U2331 (N_2331,In_1028,In_250);
or U2332 (N_2332,In_844,In_1299);
xor U2333 (N_2333,In_1256,In_344);
xor U2334 (N_2334,In_1263,In_506);
xnor U2335 (N_2335,In_1277,In_645);
nor U2336 (N_2336,In_640,In_1029);
or U2337 (N_2337,In_112,In_1207);
nand U2338 (N_2338,In_909,In_272);
and U2339 (N_2339,In_1214,In_481);
nand U2340 (N_2340,In_92,In_1163);
nand U2341 (N_2341,In_275,In_1262);
nand U2342 (N_2342,In_346,In_1320);
xnor U2343 (N_2343,In_1116,In_720);
nor U2344 (N_2344,In_538,In_1004);
or U2345 (N_2345,In_709,In_901);
nor U2346 (N_2346,In_1448,In_637);
nand U2347 (N_2347,In_1218,In_1024);
and U2348 (N_2348,In_1407,In_201);
or U2349 (N_2349,In_1012,In_1230);
xor U2350 (N_2350,In_613,In_1346);
nand U2351 (N_2351,In_996,In_38);
xnor U2352 (N_2352,In_1382,In_524);
and U2353 (N_2353,In_429,In_624);
nand U2354 (N_2354,In_462,In_762);
nand U2355 (N_2355,In_705,In_1318);
xor U2356 (N_2356,In_261,In_1497);
or U2357 (N_2357,In_827,In_816);
xnor U2358 (N_2358,In_1130,In_477);
nand U2359 (N_2359,In_77,In_1252);
nand U2360 (N_2360,In_1259,In_640);
xnor U2361 (N_2361,In_1246,In_391);
xnor U2362 (N_2362,In_553,In_656);
and U2363 (N_2363,In_224,In_1344);
nor U2364 (N_2364,In_404,In_470);
nand U2365 (N_2365,In_765,In_1377);
and U2366 (N_2366,In_49,In_914);
nand U2367 (N_2367,In_742,In_1344);
xor U2368 (N_2368,In_428,In_733);
nor U2369 (N_2369,In_1233,In_1440);
and U2370 (N_2370,In_1499,In_1239);
nand U2371 (N_2371,In_640,In_838);
xor U2372 (N_2372,In_57,In_1388);
or U2373 (N_2373,In_1353,In_968);
and U2374 (N_2374,In_869,In_102);
xor U2375 (N_2375,In_555,In_180);
nor U2376 (N_2376,In_910,In_890);
xnor U2377 (N_2377,In_1342,In_1457);
nor U2378 (N_2378,In_49,In_605);
and U2379 (N_2379,In_602,In_281);
nor U2380 (N_2380,In_1064,In_367);
nor U2381 (N_2381,In_1094,In_1424);
nor U2382 (N_2382,In_569,In_548);
xnor U2383 (N_2383,In_42,In_188);
and U2384 (N_2384,In_1352,In_1345);
and U2385 (N_2385,In_798,In_945);
xnor U2386 (N_2386,In_877,In_1090);
nor U2387 (N_2387,In_545,In_336);
or U2388 (N_2388,In_731,In_734);
nor U2389 (N_2389,In_174,In_1055);
xnor U2390 (N_2390,In_1,In_1060);
nor U2391 (N_2391,In_1273,In_503);
nand U2392 (N_2392,In_78,In_180);
and U2393 (N_2393,In_445,In_1170);
xnor U2394 (N_2394,In_444,In_466);
and U2395 (N_2395,In_1471,In_183);
or U2396 (N_2396,In_1384,In_1045);
and U2397 (N_2397,In_209,In_90);
or U2398 (N_2398,In_1277,In_243);
xor U2399 (N_2399,In_983,In_1424);
xor U2400 (N_2400,In_676,In_184);
and U2401 (N_2401,In_370,In_119);
or U2402 (N_2402,In_1441,In_1167);
nor U2403 (N_2403,In_562,In_146);
nor U2404 (N_2404,In_1006,In_786);
and U2405 (N_2405,In_628,In_489);
or U2406 (N_2406,In_1027,In_308);
nand U2407 (N_2407,In_460,In_637);
or U2408 (N_2408,In_177,In_666);
nand U2409 (N_2409,In_1330,In_493);
xor U2410 (N_2410,In_788,In_708);
nand U2411 (N_2411,In_724,In_79);
xnor U2412 (N_2412,In_1010,In_1190);
xor U2413 (N_2413,In_1459,In_761);
or U2414 (N_2414,In_260,In_237);
nor U2415 (N_2415,In_1319,In_926);
xnor U2416 (N_2416,In_1271,In_557);
nor U2417 (N_2417,In_1051,In_1081);
nor U2418 (N_2418,In_755,In_109);
nor U2419 (N_2419,In_446,In_524);
nor U2420 (N_2420,In_7,In_943);
or U2421 (N_2421,In_763,In_393);
and U2422 (N_2422,In_1353,In_752);
nand U2423 (N_2423,In_896,In_437);
xnor U2424 (N_2424,In_997,In_467);
nand U2425 (N_2425,In_784,In_450);
xor U2426 (N_2426,In_402,In_771);
and U2427 (N_2427,In_1069,In_373);
and U2428 (N_2428,In_1454,In_573);
nor U2429 (N_2429,In_892,In_458);
xnor U2430 (N_2430,In_1307,In_688);
nand U2431 (N_2431,In_534,In_805);
xor U2432 (N_2432,In_1165,In_14);
or U2433 (N_2433,In_367,In_137);
or U2434 (N_2434,In_93,In_223);
nor U2435 (N_2435,In_41,In_324);
nand U2436 (N_2436,In_927,In_1321);
nor U2437 (N_2437,In_1456,In_1006);
xnor U2438 (N_2438,In_616,In_900);
nor U2439 (N_2439,In_1390,In_833);
xnor U2440 (N_2440,In_604,In_242);
xnor U2441 (N_2441,In_1461,In_1117);
xor U2442 (N_2442,In_890,In_449);
nand U2443 (N_2443,In_314,In_778);
xor U2444 (N_2444,In_697,In_1123);
nor U2445 (N_2445,In_1213,In_1152);
and U2446 (N_2446,In_827,In_1107);
nor U2447 (N_2447,In_893,In_1105);
and U2448 (N_2448,In_903,In_292);
nor U2449 (N_2449,In_329,In_590);
nor U2450 (N_2450,In_697,In_325);
nand U2451 (N_2451,In_1141,In_747);
xor U2452 (N_2452,In_461,In_880);
nand U2453 (N_2453,In_813,In_140);
xor U2454 (N_2454,In_1078,In_889);
xor U2455 (N_2455,In_622,In_299);
or U2456 (N_2456,In_11,In_273);
nor U2457 (N_2457,In_135,In_724);
and U2458 (N_2458,In_850,In_1389);
nor U2459 (N_2459,In_527,In_104);
and U2460 (N_2460,In_27,In_419);
and U2461 (N_2461,In_1026,In_324);
nor U2462 (N_2462,In_972,In_211);
nor U2463 (N_2463,In_1241,In_580);
xnor U2464 (N_2464,In_549,In_190);
or U2465 (N_2465,In_1453,In_1099);
and U2466 (N_2466,In_1255,In_770);
nor U2467 (N_2467,In_567,In_471);
nand U2468 (N_2468,In_13,In_1429);
nor U2469 (N_2469,In_873,In_1332);
nand U2470 (N_2470,In_513,In_416);
and U2471 (N_2471,In_483,In_1431);
nand U2472 (N_2472,In_1301,In_689);
nor U2473 (N_2473,In_522,In_3);
and U2474 (N_2474,In_1120,In_43);
or U2475 (N_2475,In_264,In_1382);
and U2476 (N_2476,In_1021,In_422);
nor U2477 (N_2477,In_529,In_682);
nand U2478 (N_2478,In_207,In_1373);
nand U2479 (N_2479,In_1124,In_1464);
and U2480 (N_2480,In_1226,In_505);
and U2481 (N_2481,In_480,In_643);
xor U2482 (N_2482,In_909,In_6);
or U2483 (N_2483,In_58,In_647);
nor U2484 (N_2484,In_31,In_218);
nand U2485 (N_2485,In_119,In_373);
and U2486 (N_2486,In_731,In_1105);
and U2487 (N_2487,In_1239,In_98);
xnor U2488 (N_2488,In_983,In_81);
or U2489 (N_2489,In_867,In_37);
xor U2490 (N_2490,In_497,In_919);
nand U2491 (N_2491,In_1332,In_417);
and U2492 (N_2492,In_19,In_1021);
xor U2493 (N_2493,In_606,In_973);
nand U2494 (N_2494,In_153,In_1437);
and U2495 (N_2495,In_759,In_374);
and U2496 (N_2496,In_1300,In_869);
xor U2497 (N_2497,In_913,In_455);
or U2498 (N_2498,In_524,In_387);
and U2499 (N_2499,In_325,In_34);
or U2500 (N_2500,In_612,In_1263);
or U2501 (N_2501,In_786,In_1014);
or U2502 (N_2502,In_663,In_307);
or U2503 (N_2503,In_223,In_240);
xor U2504 (N_2504,In_288,In_1396);
or U2505 (N_2505,In_258,In_1114);
or U2506 (N_2506,In_1014,In_835);
nand U2507 (N_2507,In_916,In_444);
or U2508 (N_2508,In_675,In_307);
xnor U2509 (N_2509,In_157,In_1230);
nand U2510 (N_2510,In_968,In_793);
nand U2511 (N_2511,In_24,In_1183);
nor U2512 (N_2512,In_688,In_928);
or U2513 (N_2513,In_908,In_938);
or U2514 (N_2514,In_395,In_1023);
nor U2515 (N_2515,In_210,In_1124);
nand U2516 (N_2516,In_212,In_538);
or U2517 (N_2517,In_545,In_52);
nor U2518 (N_2518,In_136,In_37);
nor U2519 (N_2519,In_635,In_273);
nand U2520 (N_2520,In_112,In_632);
nor U2521 (N_2521,In_270,In_1137);
and U2522 (N_2522,In_474,In_279);
xor U2523 (N_2523,In_1148,In_434);
nor U2524 (N_2524,In_353,In_1065);
or U2525 (N_2525,In_1111,In_111);
xor U2526 (N_2526,In_301,In_1037);
xnor U2527 (N_2527,In_1321,In_80);
nor U2528 (N_2528,In_944,In_950);
nand U2529 (N_2529,In_112,In_1287);
or U2530 (N_2530,In_972,In_672);
xnor U2531 (N_2531,In_865,In_1335);
nand U2532 (N_2532,In_1010,In_29);
or U2533 (N_2533,In_714,In_1142);
xnor U2534 (N_2534,In_887,In_704);
or U2535 (N_2535,In_1243,In_475);
nor U2536 (N_2536,In_103,In_1444);
xnor U2537 (N_2537,In_150,In_1342);
or U2538 (N_2538,In_418,In_362);
nor U2539 (N_2539,In_182,In_1200);
nor U2540 (N_2540,In_307,In_1113);
nor U2541 (N_2541,In_173,In_906);
and U2542 (N_2542,In_28,In_265);
nand U2543 (N_2543,In_452,In_444);
nor U2544 (N_2544,In_996,In_1034);
and U2545 (N_2545,In_900,In_808);
nor U2546 (N_2546,In_334,In_1104);
and U2547 (N_2547,In_214,In_954);
or U2548 (N_2548,In_562,In_11);
nand U2549 (N_2549,In_289,In_933);
and U2550 (N_2550,In_1016,In_1162);
xor U2551 (N_2551,In_1009,In_816);
or U2552 (N_2552,In_1190,In_729);
and U2553 (N_2553,In_310,In_629);
or U2554 (N_2554,In_635,In_242);
or U2555 (N_2555,In_1497,In_666);
or U2556 (N_2556,In_1216,In_487);
nor U2557 (N_2557,In_449,In_581);
xor U2558 (N_2558,In_1349,In_780);
and U2559 (N_2559,In_380,In_229);
nor U2560 (N_2560,In_174,In_1224);
and U2561 (N_2561,In_1421,In_1109);
or U2562 (N_2562,In_0,In_476);
nor U2563 (N_2563,In_831,In_1445);
nor U2564 (N_2564,In_961,In_163);
xnor U2565 (N_2565,In_1180,In_393);
or U2566 (N_2566,In_885,In_430);
xor U2567 (N_2567,In_309,In_1250);
and U2568 (N_2568,In_424,In_625);
nor U2569 (N_2569,In_1147,In_323);
nand U2570 (N_2570,In_715,In_1250);
and U2571 (N_2571,In_1273,In_67);
nor U2572 (N_2572,In_773,In_316);
nand U2573 (N_2573,In_614,In_879);
and U2574 (N_2574,In_1094,In_659);
xor U2575 (N_2575,In_339,In_1210);
xor U2576 (N_2576,In_41,In_125);
xnor U2577 (N_2577,In_327,In_294);
and U2578 (N_2578,In_714,In_474);
nor U2579 (N_2579,In_141,In_1169);
xor U2580 (N_2580,In_1356,In_419);
xnor U2581 (N_2581,In_514,In_971);
or U2582 (N_2582,In_879,In_179);
nand U2583 (N_2583,In_620,In_636);
or U2584 (N_2584,In_316,In_1196);
or U2585 (N_2585,In_878,In_925);
xor U2586 (N_2586,In_483,In_1276);
nor U2587 (N_2587,In_205,In_1147);
and U2588 (N_2588,In_560,In_85);
nand U2589 (N_2589,In_1475,In_1411);
nor U2590 (N_2590,In_1307,In_169);
xnor U2591 (N_2591,In_156,In_586);
nand U2592 (N_2592,In_1426,In_1124);
or U2593 (N_2593,In_776,In_460);
nor U2594 (N_2594,In_1114,In_837);
nor U2595 (N_2595,In_1388,In_829);
nand U2596 (N_2596,In_758,In_603);
nand U2597 (N_2597,In_657,In_1365);
nand U2598 (N_2598,In_627,In_647);
nand U2599 (N_2599,In_185,In_942);
nor U2600 (N_2600,In_6,In_194);
nor U2601 (N_2601,In_587,In_892);
and U2602 (N_2602,In_1150,In_1142);
and U2603 (N_2603,In_687,In_356);
nor U2604 (N_2604,In_592,In_196);
and U2605 (N_2605,In_1277,In_412);
or U2606 (N_2606,In_1125,In_1255);
or U2607 (N_2607,In_1135,In_1415);
xnor U2608 (N_2608,In_405,In_36);
xnor U2609 (N_2609,In_56,In_364);
xnor U2610 (N_2610,In_477,In_172);
or U2611 (N_2611,In_1037,In_1387);
xnor U2612 (N_2612,In_58,In_771);
nand U2613 (N_2613,In_681,In_975);
xnor U2614 (N_2614,In_259,In_1232);
and U2615 (N_2615,In_842,In_1422);
or U2616 (N_2616,In_695,In_510);
xor U2617 (N_2617,In_365,In_685);
or U2618 (N_2618,In_788,In_913);
nand U2619 (N_2619,In_832,In_1444);
and U2620 (N_2620,In_1070,In_1218);
xnor U2621 (N_2621,In_1211,In_1023);
nor U2622 (N_2622,In_451,In_1204);
xor U2623 (N_2623,In_627,In_1110);
or U2624 (N_2624,In_747,In_82);
or U2625 (N_2625,In_1332,In_275);
nor U2626 (N_2626,In_719,In_1164);
nand U2627 (N_2627,In_1276,In_694);
nand U2628 (N_2628,In_1405,In_546);
xor U2629 (N_2629,In_337,In_547);
xor U2630 (N_2630,In_1444,In_930);
or U2631 (N_2631,In_207,In_70);
nor U2632 (N_2632,In_1495,In_79);
nor U2633 (N_2633,In_249,In_538);
nand U2634 (N_2634,In_436,In_404);
nand U2635 (N_2635,In_21,In_493);
xnor U2636 (N_2636,In_797,In_562);
nor U2637 (N_2637,In_1414,In_1245);
or U2638 (N_2638,In_1482,In_1170);
xnor U2639 (N_2639,In_1478,In_241);
nand U2640 (N_2640,In_978,In_1277);
nor U2641 (N_2641,In_905,In_1216);
or U2642 (N_2642,In_318,In_1216);
nor U2643 (N_2643,In_371,In_1407);
nand U2644 (N_2644,In_1242,In_159);
and U2645 (N_2645,In_1221,In_998);
nand U2646 (N_2646,In_874,In_207);
and U2647 (N_2647,In_928,In_610);
xnor U2648 (N_2648,In_589,In_1340);
or U2649 (N_2649,In_383,In_573);
or U2650 (N_2650,In_919,In_54);
xor U2651 (N_2651,In_164,In_471);
and U2652 (N_2652,In_462,In_1076);
or U2653 (N_2653,In_1334,In_928);
nor U2654 (N_2654,In_1108,In_314);
nand U2655 (N_2655,In_1344,In_631);
nand U2656 (N_2656,In_530,In_278);
xnor U2657 (N_2657,In_1123,In_1044);
nand U2658 (N_2658,In_1177,In_446);
xnor U2659 (N_2659,In_1144,In_83);
nor U2660 (N_2660,In_407,In_1427);
xnor U2661 (N_2661,In_1026,In_247);
or U2662 (N_2662,In_966,In_1249);
xnor U2663 (N_2663,In_277,In_1478);
or U2664 (N_2664,In_233,In_1452);
or U2665 (N_2665,In_632,In_1057);
and U2666 (N_2666,In_1422,In_1359);
nor U2667 (N_2667,In_1323,In_288);
or U2668 (N_2668,In_55,In_934);
or U2669 (N_2669,In_1077,In_808);
nor U2670 (N_2670,In_1239,In_708);
nor U2671 (N_2671,In_207,In_727);
xor U2672 (N_2672,In_265,In_1484);
xor U2673 (N_2673,In_1375,In_104);
xor U2674 (N_2674,In_179,In_719);
or U2675 (N_2675,In_133,In_484);
xnor U2676 (N_2676,In_1129,In_405);
nor U2677 (N_2677,In_1424,In_187);
xor U2678 (N_2678,In_1201,In_933);
nand U2679 (N_2679,In_1318,In_1412);
and U2680 (N_2680,In_130,In_819);
nor U2681 (N_2681,In_305,In_1183);
or U2682 (N_2682,In_626,In_522);
or U2683 (N_2683,In_1394,In_450);
or U2684 (N_2684,In_143,In_200);
xor U2685 (N_2685,In_210,In_885);
or U2686 (N_2686,In_591,In_800);
or U2687 (N_2687,In_252,In_882);
xor U2688 (N_2688,In_159,In_1033);
and U2689 (N_2689,In_622,In_1041);
and U2690 (N_2690,In_1304,In_459);
nand U2691 (N_2691,In_982,In_1076);
and U2692 (N_2692,In_1338,In_1321);
xor U2693 (N_2693,In_453,In_1495);
or U2694 (N_2694,In_329,In_1210);
nand U2695 (N_2695,In_1369,In_1105);
nand U2696 (N_2696,In_452,In_67);
nor U2697 (N_2697,In_152,In_669);
nor U2698 (N_2698,In_568,In_1354);
or U2699 (N_2699,In_836,In_805);
nor U2700 (N_2700,In_290,In_392);
xor U2701 (N_2701,In_922,In_1496);
or U2702 (N_2702,In_1365,In_761);
nand U2703 (N_2703,In_1177,In_1298);
xor U2704 (N_2704,In_1356,In_477);
and U2705 (N_2705,In_818,In_856);
xor U2706 (N_2706,In_852,In_221);
and U2707 (N_2707,In_50,In_237);
nor U2708 (N_2708,In_1403,In_361);
nand U2709 (N_2709,In_205,In_430);
xor U2710 (N_2710,In_17,In_355);
nor U2711 (N_2711,In_521,In_117);
xor U2712 (N_2712,In_760,In_1393);
and U2713 (N_2713,In_697,In_438);
nand U2714 (N_2714,In_496,In_63);
nand U2715 (N_2715,In_1326,In_1409);
or U2716 (N_2716,In_121,In_881);
and U2717 (N_2717,In_131,In_529);
and U2718 (N_2718,In_763,In_646);
and U2719 (N_2719,In_110,In_1326);
nor U2720 (N_2720,In_1363,In_969);
nor U2721 (N_2721,In_495,In_92);
xor U2722 (N_2722,In_1004,In_407);
xor U2723 (N_2723,In_1326,In_968);
xnor U2724 (N_2724,In_1111,In_1377);
or U2725 (N_2725,In_241,In_1156);
xnor U2726 (N_2726,In_520,In_1421);
or U2727 (N_2727,In_924,In_1162);
xor U2728 (N_2728,In_920,In_747);
xnor U2729 (N_2729,In_244,In_356);
or U2730 (N_2730,In_628,In_1302);
xnor U2731 (N_2731,In_1097,In_546);
nand U2732 (N_2732,In_1101,In_1370);
or U2733 (N_2733,In_1393,In_840);
nand U2734 (N_2734,In_997,In_1097);
xor U2735 (N_2735,In_1383,In_655);
or U2736 (N_2736,In_490,In_78);
and U2737 (N_2737,In_163,In_575);
nor U2738 (N_2738,In_514,In_1284);
or U2739 (N_2739,In_1004,In_1226);
nor U2740 (N_2740,In_1234,In_1008);
xnor U2741 (N_2741,In_1021,In_674);
nor U2742 (N_2742,In_1361,In_480);
or U2743 (N_2743,In_376,In_491);
and U2744 (N_2744,In_689,In_979);
nand U2745 (N_2745,In_616,In_268);
xor U2746 (N_2746,In_1138,In_395);
or U2747 (N_2747,In_158,In_384);
and U2748 (N_2748,In_719,In_364);
or U2749 (N_2749,In_878,In_1245);
or U2750 (N_2750,In_996,In_1046);
xor U2751 (N_2751,In_932,In_1047);
nor U2752 (N_2752,In_1225,In_777);
xor U2753 (N_2753,In_570,In_912);
xor U2754 (N_2754,In_236,In_821);
nor U2755 (N_2755,In_379,In_957);
and U2756 (N_2756,In_325,In_261);
nand U2757 (N_2757,In_154,In_1453);
nor U2758 (N_2758,In_1229,In_96);
nand U2759 (N_2759,In_1474,In_437);
and U2760 (N_2760,In_1037,In_413);
xor U2761 (N_2761,In_1475,In_98);
or U2762 (N_2762,In_941,In_850);
and U2763 (N_2763,In_4,In_726);
nand U2764 (N_2764,In_243,In_75);
or U2765 (N_2765,In_1018,In_929);
nand U2766 (N_2766,In_1265,In_1313);
or U2767 (N_2767,In_774,In_1451);
nand U2768 (N_2768,In_256,In_179);
and U2769 (N_2769,In_815,In_1057);
and U2770 (N_2770,In_1075,In_1467);
xor U2771 (N_2771,In_690,In_305);
nor U2772 (N_2772,In_1135,In_1398);
xnor U2773 (N_2773,In_167,In_317);
and U2774 (N_2774,In_774,In_469);
and U2775 (N_2775,In_335,In_1295);
xnor U2776 (N_2776,In_1269,In_1391);
nand U2777 (N_2777,In_586,In_816);
nand U2778 (N_2778,In_522,In_893);
xor U2779 (N_2779,In_334,In_294);
nor U2780 (N_2780,In_114,In_1043);
nand U2781 (N_2781,In_1473,In_1491);
xor U2782 (N_2782,In_1413,In_749);
nand U2783 (N_2783,In_796,In_639);
or U2784 (N_2784,In_1212,In_1248);
nor U2785 (N_2785,In_486,In_942);
nand U2786 (N_2786,In_383,In_1196);
or U2787 (N_2787,In_415,In_1072);
and U2788 (N_2788,In_236,In_1314);
nand U2789 (N_2789,In_58,In_1338);
nand U2790 (N_2790,In_528,In_1379);
and U2791 (N_2791,In_216,In_329);
or U2792 (N_2792,In_31,In_383);
or U2793 (N_2793,In_1048,In_1169);
and U2794 (N_2794,In_499,In_906);
nor U2795 (N_2795,In_541,In_1465);
nand U2796 (N_2796,In_576,In_1166);
or U2797 (N_2797,In_1398,In_741);
and U2798 (N_2798,In_1349,In_960);
nand U2799 (N_2799,In_1261,In_952);
nor U2800 (N_2800,In_401,In_122);
nand U2801 (N_2801,In_1388,In_1039);
xnor U2802 (N_2802,In_371,In_4);
nand U2803 (N_2803,In_1058,In_1395);
nor U2804 (N_2804,In_1297,In_158);
nor U2805 (N_2805,In_107,In_1122);
nand U2806 (N_2806,In_432,In_836);
nand U2807 (N_2807,In_479,In_1273);
or U2808 (N_2808,In_1132,In_102);
xnor U2809 (N_2809,In_981,In_290);
nor U2810 (N_2810,In_222,In_1375);
xnor U2811 (N_2811,In_510,In_666);
nor U2812 (N_2812,In_1265,In_1495);
xnor U2813 (N_2813,In_983,In_513);
and U2814 (N_2814,In_201,In_1117);
nor U2815 (N_2815,In_498,In_293);
and U2816 (N_2816,In_958,In_1126);
or U2817 (N_2817,In_475,In_105);
and U2818 (N_2818,In_1375,In_577);
or U2819 (N_2819,In_1482,In_1140);
and U2820 (N_2820,In_1349,In_159);
xnor U2821 (N_2821,In_392,In_149);
or U2822 (N_2822,In_77,In_754);
or U2823 (N_2823,In_435,In_510);
or U2824 (N_2824,In_1074,In_1236);
and U2825 (N_2825,In_326,In_819);
nor U2826 (N_2826,In_1438,In_26);
xnor U2827 (N_2827,In_230,In_775);
and U2828 (N_2828,In_236,In_1093);
nor U2829 (N_2829,In_469,In_93);
or U2830 (N_2830,In_865,In_174);
or U2831 (N_2831,In_712,In_81);
nor U2832 (N_2832,In_1018,In_896);
xor U2833 (N_2833,In_1066,In_1210);
or U2834 (N_2834,In_248,In_1120);
and U2835 (N_2835,In_1150,In_211);
nand U2836 (N_2836,In_37,In_733);
nor U2837 (N_2837,In_314,In_720);
nand U2838 (N_2838,In_1466,In_459);
or U2839 (N_2839,In_902,In_394);
nor U2840 (N_2840,In_246,In_353);
or U2841 (N_2841,In_1110,In_474);
and U2842 (N_2842,In_1346,In_1273);
and U2843 (N_2843,In_418,In_1333);
or U2844 (N_2844,In_1360,In_1144);
nor U2845 (N_2845,In_754,In_63);
nor U2846 (N_2846,In_184,In_499);
nand U2847 (N_2847,In_680,In_1034);
and U2848 (N_2848,In_646,In_180);
and U2849 (N_2849,In_66,In_1290);
nand U2850 (N_2850,In_17,In_618);
nand U2851 (N_2851,In_875,In_61);
nand U2852 (N_2852,In_260,In_238);
xnor U2853 (N_2853,In_1175,In_1151);
nor U2854 (N_2854,In_1128,In_1468);
nand U2855 (N_2855,In_672,In_907);
and U2856 (N_2856,In_1324,In_1308);
nor U2857 (N_2857,In_368,In_775);
nand U2858 (N_2858,In_557,In_396);
xor U2859 (N_2859,In_1002,In_732);
or U2860 (N_2860,In_1285,In_1064);
nand U2861 (N_2861,In_1399,In_213);
and U2862 (N_2862,In_329,In_774);
xnor U2863 (N_2863,In_1109,In_1032);
xor U2864 (N_2864,In_1346,In_183);
nand U2865 (N_2865,In_571,In_110);
xor U2866 (N_2866,In_1066,In_1125);
or U2867 (N_2867,In_976,In_195);
and U2868 (N_2868,In_973,In_687);
or U2869 (N_2869,In_123,In_848);
xor U2870 (N_2870,In_1471,In_441);
or U2871 (N_2871,In_67,In_1352);
or U2872 (N_2872,In_1226,In_1384);
and U2873 (N_2873,In_707,In_972);
and U2874 (N_2874,In_808,In_1332);
or U2875 (N_2875,In_1298,In_1441);
nor U2876 (N_2876,In_874,In_382);
or U2877 (N_2877,In_1307,In_1013);
nand U2878 (N_2878,In_697,In_47);
or U2879 (N_2879,In_1073,In_1249);
and U2880 (N_2880,In_699,In_1474);
nand U2881 (N_2881,In_949,In_69);
xor U2882 (N_2882,In_995,In_612);
xor U2883 (N_2883,In_785,In_1471);
nand U2884 (N_2884,In_928,In_136);
xor U2885 (N_2885,In_666,In_1188);
nand U2886 (N_2886,In_1301,In_727);
or U2887 (N_2887,In_1081,In_1222);
nor U2888 (N_2888,In_752,In_491);
nor U2889 (N_2889,In_937,In_599);
or U2890 (N_2890,In_264,In_923);
nor U2891 (N_2891,In_1498,In_296);
or U2892 (N_2892,In_115,In_1204);
xnor U2893 (N_2893,In_611,In_980);
xnor U2894 (N_2894,In_404,In_19);
and U2895 (N_2895,In_537,In_1192);
nand U2896 (N_2896,In_80,In_758);
xor U2897 (N_2897,In_1301,In_350);
or U2898 (N_2898,In_679,In_964);
nand U2899 (N_2899,In_168,In_152);
nor U2900 (N_2900,In_1242,In_1234);
and U2901 (N_2901,In_705,In_270);
nor U2902 (N_2902,In_268,In_94);
or U2903 (N_2903,In_1442,In_326);
and U2904 (N_2904,In_671,In_711);
and U2905 (N_2905,In_678,In_1022);
xnor U2906 (N_2906,In_330,In_406);
xor U2907 (N_2907,In_499,In_1090);
and U2908 (N_2908,In_577,In_1231);
xor U2909 (N_2909,In_222,In_1394);
xnor U2910 (N_2910,In_813,In_45);
xnor U2911 (N_2911,In_1150,In_638);
xor U2912 (N_2912,In_888,In_371);
nor U2913 (N_2913,In_1424,In_483);
xnor U2914 (N_2914,In_501,In_330);
or U2915 (N_2915,In_890,In_870);
nand U2916 (N_2916,In_635,In_927);
nand U2917 (N_2917,In_645,In_981);
xor U2918 (N_2918,In_834,In_559);
nor U2919 (N_2919,In_1052,In_232);
nand U2920 (N_2920,In_827,In_754);
nor U2921 (N_2921,In_1197,In_256);
xnor U2922 (N_2922,In_20,In_584);
nand U2923 (N_2923,In_535,In_1198);
and U2924 (N_2924,In_502,In_4);
xnor U2925 (N_2925,In_715,In_86);
and U2926 (N_2926,In_1087,In_1221);
xnor U2927 (N_2927,In_1233,In_511);
and U2928 (N_2928,In_1004,In_526);
nand U2929 (N_2929,In_869,In_1266);
nand U2930 (N_2930,In_223,In_615);
xnor U2931 (N_2931,In_213,In_1179);
and U2932 (N_2932,In_366,In_1053);
xnor U2933 (N_2933,In_663,In_372);
or U2934 (N_2934,In_1333,In_1089);
xor U2935 (N_2935,In_764,In_484);
nand U2936 (N_2936,In_1380,In_1428);
xor U2937 (N_2937,In_1220,In_958);
nor U2938 (N_2938,In_74,In_182);
nor U2939 (N_2939,In_334,In_1001);
and U2940 (N_2940,In_1430,In_867);
nor U2941 (N_2941,In_1085,In_1285);
and U2942 (N_2942,In_926,In_866);
nand U2943 (N_2943,In_1086,In_1271);
nor U2944 (N_2944,In_596,In_1018);
nor U2945 (N_2945,In_889,In_290);
xnor U2946 (N_2946,In_703,In_121);
xnor U2947 (N_2947,In_889,In_106);
nand U2948 (N_2948,In_699,In_1095);
xnor U2949 (N_2949,In_1065,In_149);
xnor U2950 (N_2950,In_1000,In_39);
or U2951 (N_2951,In_1391,In_708);
nor U2952 (N_2952,In_799,In_435);
or U2953 (N_2953,In_865,In_100);
or U2954 (N_2954,In_732,In_1436);
and U2955 (N_2955,In_909,In_1207);
or U2956 (N_2956,In_584,In_254);
or U2957 (N_2957,In_4,In_355);
nand U2958 (N_2958,In_1327,In_724);
nor U2959 (N_2959,In_1343,In_784);
or U2960 (N_2960,In_1361,In_601);
or U2961 (N_2961,In_597,In_1037);
nor U2962 (N_2962,In_519,In_1172);
nand U2963 (N_2963,In_245,In_670);
or U2964 (N_2964,In_57,In_736);
xor U2965 (N_2965,In_1422,In_11);
or U2966 (N_2966,In_876,In_1023);
nor U2967 (N_2967,In_438,In_1212);
xor U2968 (N_2968,In_194,In_9);
xor U2969 (N_2969,In_910,In_1077);
xnor U2970 (N_2970,In_522,In_955);
nand U2971 (N_2971,In_1220,In_297);
nor U2972 (N_2972,In_1019,In_1148);
nor U2973 (N_2973,In_766,In_1333);
nand U2974 (N_2974,In_1223,In_1116);
nor U2975 (N_2975,In_1001,In_736);
xor U2976 (N_2976,In_70,In_382);
xnor U2977 (N_2977,In_632,In_1243);
nor U2978 (N_2978,In_1334,In_578);
nor U2979 (N_2979,In_795,In_1175);
xnor U2980 (N_2980,In_102,In_910);
nor U2981 (N_2981,In_1495,In_1065);
or U2982 (N_2982,In_1011,In_38);
or U2983 (N_2983,In_1485,In_356);
xnor U2984 (N_2984,In_972,In_1097);
or U2985 (N_2985,In_234,In_1063);
nand U2986 (N_2986,In_2,In_756);
nand U2987 (N_2987,In_1178,In_880);
xor U2988 (N_2988,In_620,In_915);
xor U2989 (N_2989,In_644,In_1012);
or U2990 (N_2990,In_454,In_74);
xnor U2991 (N_2991,In_1263,In_1310);
xor U2992 (N_2992,In_1381,In_1016);
nor U2993 (N_2993,In_1445,In_19);
xnor U2994 (N_2994,In_944,In_544);
nand U2995 (N_2995,In_521,In_166);
nand U2996 (N_2996,In_55,In_802);
or U2997 (N_2997,In_67,In_17);
nor U2998 (N_2998,In_108,In_1036);
xor U2999 (N_2999,In_1436,In_929);
or U3000 (N_3000,In_1059,In_478);
or U3001 (N_3001,In_768,In_1121);
and U3002 (N_3002,In_839,In_1001);
nor U3003 (N_3003,In_921,In_1226);
xnor U3004 (N_3004,In_1478,In_340);
or U3005 (N_3005,In_772,In_1180);
nand U3006 (N_3006,In_1033,In_858);
and U3007 (N_3007,In_995,In_948);
nand U3008 (N_3008,In_1386,In_863);
xor U3009 (N_3009,In_39,In_442);
xnor U3010 (N_3010,In_698,In_125);
nand U3011 (N_3011,In_951,In_1238);
nand U3012 (N_3012,In_1491,In_1298);
nor U3013 (N_3013,In_277,In_573);
or U3014 (N_3014,In_926,In_357);
or U3015 (N_3015,In_426,In_407);
nor U3016 (N_3016,In_1234,In_172);
or U3017 (N_3017,In_998,In_1433);
or U3018 (N_3018,In_1029,In_956);
nor U3019 (N_3019,In_947,In_37);
nand U3020 (N_3020,In_1479,In_1306);
and U3021 (N_3021,In_994,In_440);
nand U3022 (N_3022,In_59,In_541);
or U3023 (N_3023,In_1179,In_429);
and U3024 (N_3024,In_407,In_77);
nand U3025 (N_3025,In_1246,In_887);
or U3026 (N_3026,In_1448,In_510);
or U3027 (N_3027,In_1092,In_910);
xor U3028 (N_3028,In_584,In_1458);
xnor U3029 (N_3029,In_1348,In_1422);
nor U3030 (N_3030,In_382,In_508);
and U3031 (N_3031,In_58,In_436);
xnor U3032 (N_3032,In_349,In_611);
xnor U3033 (N_3033,In_334,In_451);
and U3034 (N_3034,In_1308,In_212);
or U3035 (N_3035,In_1245,In_331);
xor U3036 (N_3036,In_326,In_532);
nor U3037 (N_3037,In_78,In_422);
nand U3038 (N_3038,In_554,In_261);
nor U3039 (N_3039,In_665,In_1214);
xnor U3040 (N_3040,In_1113,In_396);
or U3041 (N_3041,In_80,In_1143);
or U3042 (N_3042,In_158,In_924);
and U3043 (N_3043,In_387,In_345);
and U3044 (N_3044,In_1078,In_744);
nor U3045 (N_3045,In_1429,In_1445);
nor U3046 (N_3046,In_659,In_1277);
and U3047 (N_3047,In_77,In_653);
and U3048 (N_3048,In_772,In_259);
nand U3049 (N_3049,In_792,In_1218);
and U3050 (N_3050,In_91,In_599);
nor U3051 (N_3051,In_631,In_333);
nand U3052 (N_3052,In_432,In_973);
or U3053 (N_3053,In_1001,In_888);
and U3054 (N_3054,In_750,In_858);
nor U3055 (N_3055,In_607,In_1403);
and U3056 (N_3056,In_560,In_903);
and U3057 (N_3057,In_921,In_111);
nand U3058 (N_3058,In_1094,In_1427);
and U3059 (N_3059,In_935,In_430);
xnor U3060 (N_3060,In_762,In_784);
and U3061 (N_3061,In_375,In_1453);
nand U3062 (N_3062,In_345,In_49);
nand U3063 (N_3063,In_107,In_1475);
nand U3064 (N_3064,In_151,In_620);
and U3065 (N_3065,In_1304,In_962);
or U3066 (N_3066,In_1305,In_406);
nor U3067 (N_3067,In_239,In_1423);
or U3068 (N_3068,In_367,In_154);
and U3069 (N_3069,In_274,In_367);
or U3070 (N_3070,In_1004,In_205);
and U3071 (N_3071,In_70,In_407);
and U3072 (N_3072,In_637,In_205);
nand U3073 (N_3073,In_330,In_850);
nand U3074 (N_3074,In_418,In_1072);
nand U3075 (N_3075,In_476,In_627);
nand U3076 (N_3076,In_1091,In_248);
xor U3077 (N_3077,In_17,In_411);
xnor U3078 (N_3078,In_897,In_1212);
or U3079 (N_3079,In_1355,In_1318);
nand U3080 (N_3080,In_659,In_265);
and U3081 (N_3081,In_1187,In_224);
nand U3082 (N_3082,In_712,In_385);
nor U3083 (N_3083,In_1267,In_1455);
xor U3084 (N_3084,In_623,In_1239);
xnor U3085 (N_3085,In_740,In_21);
xnor U3086 (N_3086,In_1051,In_356);
and U3087 (N_3087,In_744,In_1021);
and U3088 (N_3088,In_503,In_720);
nand U3089 (N_3089,In_110,In_1255);
or U3090 (N_3090,In_367,In_1468);
nand U3091 (N_3091,In_1242,In_684);
or U3092 (N_3092,In_1067,In_855);
or U3093 (N_3093,In_1104,In_1217);
nand U3094 (N_3094,In_421,In_208);
nor U3095 (N_3095,In_445,In_173);
or U3096 (N_3096,In_1463,In_1217);
xor U3097 (N_3097,In_298,In_642);
xnor U3098 (N_3098,In_998,In_674);
nand U3099 (N_3099,In_1474,In_877);
xor U3100 (N_3100,In_1414,In_1010);
xor U3101 (N_3101,In_1338,In_1043);
and U3102 (N_3102,In_729,In_11);
and U3103 (N_3103,In_539,In_664);
or U3104 (N_3104,In_489,In_664);
nor U3105 (N_3105,In_766,In_215);
or U3106 (N_3106,In_185,In_1333);
nand U3107 (N_3107,In_529,In_728);
and U3108 (N_3108,In_388,In_339);
or U3109 (N_3109,In_293,In_735);
and U3110 (N_3110,In_1001,In_1150);
and U3111 (N_3111,In_443,In_1386);
nand U3112 (N_3112,In_147,In_819);
nor U3113 (N_3113,In_86,In_592);
or U3114 (N_3114,In_456,In_130);
and U3115 (N_3115,In_257,In_731);
or U3116 (N_3116,In_854,In_293);
and U3117 (N_3117,In_52,In_375);
nor U3118 (N_3118,In_1164,In_707);
xor U3119 (N_3119,In_1432,In_187);
and U3120 (N_3120,In_72,In_979);
and U3121 (N_3121,In_893,In_646);
xor U3122 (N_3122,In_1036,In_1313);
nor U3123 (N_3123,In_1323,In_225);
nand U3124 (N_3124,In_488,In_929);
and U3125 (N_3125,In_1165,In_906);
nand U3126 (N_3126,In_1356,In_855);
nor U3127 (N_3127,In_668,In_669);
or U3128 (N_3128,In_617,In_183);
or U3129 (N_3129,In_568,In_363);
xor U3130 (N_3130,In_201,In_736);
and U3131 (N_3131,In_797,In_456);
nor U3132 (N_3132,In_534,In_839);
or U3133 (N_3133,In_1307,In_417);
nand U3134 (N_3134,In_519,In_567);
or U3135 (N_3135,In_342,In_153);
nand U3136 (N_3136,In_313,In_776);
nor U3137 (N_3137,In_143,In_858);
nand U3138 (N_3138,In_220,In_955);
nand U3139 (N_3139,In_363,In_245);
nor U3140 (N_3140,In_1144,In_866);
and U3141 (N_3141,In_6,In_49);
and U3142 (N_3142,In_671,In_899);
nor U3143 (N_3143,In_14,In_462);
and U3144 (N_3144,In_532,In_747);
nand U3145 (N_3145,In_931,In_38);
nor U3146 (N_3146,In_268,In_639);
and U3147 (N_3147,In_983,In_1274);
or U3148 (N_3148,In_165,In_548);
or U3149 (N_3149,In_1411,In_895);
xnor U3150 (N_3150,In_119,In_150);
nand U3151 (N_3151,In_248,In_567);
nor U3152 (N_3152,In_483,In_510);
nand U3153 (N_3153,In_632,In_1375);
or U3154 (N_3154,In_1447,In_996);
or U3155 (N_3155,In_1353,In_480);
nor U3156 (N_3156,In_653,In_513);
nor U3157 (N_3157,In_1460,In_65);
and U3158 (N_3158,In_1119,In_170);
or U3159 (N_3159,In_1036,In_1271);
nor U3160 (N_3160,In_986,In_951);
nor U3161 (N_3161,In_770,In_1444);
or U3162 (N_3162,In_1286,In_879);
and U3163 (N_3163,In_1075,In_315);
nor U3164 (N_3164,In_1487,In_806);
nor U3165 (N_3165,In_841,In_748);
nand U3166 (N_3166,In_1131,In_458);
nand U3167 (N_3167,In_693,In_1423);
and U3168 (N_3168,In_12,In_952);
nor U3169 (N_3169,In_330,In_1165);
and U3170 (N_3170,In_832,In_558);
nor U3171 (N_3171,In_1329,In_11);
and U3172 (N_3172,In_557,In_230);
and U3173 (N_3173,In_874,In_637);
and U3174 (N_3174,In_1319,In_950);
xor U3175 (N_3175,In_975,In_250);
and U3176 (N_3176,In_989,In_181);
xnor U3177 (N_3177,In_215,In_787);
or U3178 (N_3178,In_683,In_1213);
or U3179 (N_3179,In_808,In_49);
xor U3180 (N_3180,In_1298,In_719);
nor U3181 (N_3181,In_1061,In_1403);
and U3182 (N_3182,In_495,In_206);
nor U3183 (N_3183,In_873,In_411);
and U3184 (N_3184,In_361,In_357);
xor U3185 (N_3185,In_233,In_208);
nor U3186 (N_3186,In_1385,In_14);
or U3187 (N_3187,In_827,In_1257);
nor U3188 (N_3188,In_1487,In_964);
and U3189 (N_3189,In_1053,In_1314);
xor U3190 (N_3190,In_657,In_867);
and U3191 (N_3191,In_681,In_1117);
or U3192 (N_3192,In_1482,In_300);
or U3193 (N_3193,In_136,In_1000);
nor U3194 (N_3194,In_1120,In_1048);
or U3195 (N_3195,In_1278,In_683);
or U3196 (N_3196,In_726,In_1403);
or U3197 (N_3197,In_1426,In_562);
nand U3198 (N_3198,In_947,In_1229);
nand U3199 (N_3199,In_793,In_1111);
nor U3200 (N_3200,In_753,In_1027);
xnor U3201 (N_3201,In_159,In_425);
xor U3202 (N_3202,In_477,In_940);
nor U3203 (N_3203,In_528,In_237);
or U3204 (N_3204,In_655,In_973);
xnor U3205 (N_3205,In_1391,In_1089);
nand U3206 (N_3206,In_46,In_618);
nand U3207 (N_3207,In_494,In_1181);
and U3208 (N_3208,In_41,In_404);
nor U3209 (N_3209,In_703,In_1225);
nor U3210 (N_3210,In_899,In_947);
nand U3211 (N_3211,In_1115,In_1276);
nand U3212 (N_3212,In_1106,In_1452);
nor U3213 (N_3213,In_1299,In_1244);
or U3214 (N_3214,In_842,In_1070);
xor U3215 (N_3215,In_1443,In_709);
and U3216 (N_3216,In_1086,In_560);
nand U3217 (N_3217,In_766,In_109);
nor U3218 (N_3218,In_1046,In_2);
and U3219 (N_3219,In_1334,In_1142);
nor U3220 (N_3220,In_1472,In_116);
xnor U3221 (N_3221,In_8,In_1250);
and U3222 (N_3222,In_188,In_1366);
or U3223 (N_3223,In_426,In_1003);
and U3224 (N_3224,In_1421,In_909);
xnor U3225 (N_3225,In_740,In_196);
nand U3226 (N_3226,In_987,In_919);
and U3227 (N_3227,In_574,In_504);
and U3228 (N_3228,In_1294,In_1313);
nor U3229 (N_3229,In_773,In_151);
xor U3230 (N_3230,In_579,In_1049);
nor U3231 (N_3231,In_268,In_1421);
and U3232 (N_3232,In_1488,In_1082);
xnor U3233 (N_3233,In_1390,In_639);
and U3234 (N_3234,In_469,In_163);
nor U3235 (N_3235,In_148,In_142);
or U3236 (N_3236,In_616,In_445);
xnor U3237 (N_3237,In_1395,In_397);
nor U3238 (N_3238,In_976,In_887);
nor U3239 (N_3239,In_810,In_269);
nand U3240 (N_3240,In_119,In_33);
nand U3241 (N_3241,In_206,In_1399);
and U3242 (N_3242,In_206,In_1448);
nor U3243 (N_3243,In_1333,In_812);
xnor U3244 (N_3244,In_969,In_1210);
or U3245 (N_3245,In_1271,In_872);
nor U3246 (N_3246,In_322,In_1342);
xnor U3247 (N_3247,In_858,In_1411);
and U3248 (N_3248,In_1419,In_148);
nand U3249 (N_3249,In_885,In_1143);
nand U3250 (N_3250,In_142,In_1362);
xor U3251 (N_3251,In_852,In_1332);
nor U3252 (N_3252,In_1265,In_213);
nor U3253 (N_3253,In_1474,In_561);
and U3254 (N_3254,In_1414,In_969);
xnor U3255 (N_3255,In_273,In_1465);
nand U3256 (N_3256,In_955,In_374);
or U3257 (N_3257,In_209,In_866);
nor U3258 (N_3258,In_840,In_1213);
nor U3259 (N_3259,In_477,In_95);
xnor U3260 (N_3260,In_1117,In_1297);
or U3261 (N_3261,In_1282,In_281);
or U3262 (N_3262,In_415,In_23);
xnor U3263 (N_3263,In_13,In_739);
xor U3264 (N_3264,In_783,In_647);
and U3265 (N_3265,In_1229,In_1117);
or U3266 (N_3266,In_1019,In_1314);
nor U3267 (N_3267,In_960,In_34);
and U3268 (N_3268,In_702,In_773);
and U3269 (N_3269,In_1315,In_314);
nor U3270 (N_3270,In_419,In_253);
nand U3271 (N_3271,In_429,In_682);
xor U3272 (N_3272,In_571,In_1044);
or U3273 (N_3273,In_1426,In_4);
nor U3274 (N_3274,In_1405,In_394);
or U3275 (N_3275,In_1304,In_1035);
and U3276 (N_3276,In_246,In_1060);
nand U3277 (N_3277,In_1054,In_1452);
xor U3278 (N_3278,In_284,In_1265);
or U3279 (N_3279,In_1459,In_174);
xor U3280 (N_3280,In_1468,In_612);
nand U3281 (N_3281,In_139,In_235);
nand U3282 (N_3282,In_409,In_13);
nor U3283 (N_3283,In_275,In_871);
or U3284 (N_3284,In_825,In_1027);
xor U3285 (N_3285,In_224,In_1474);
or U3286 (N_3286,In_1040,In_1144);
nand U3287 (N_3287,In_1394,In_772);
nor U3288 (N_3288,In_176,In_738);
xor U3289 (N_3289,In_1277,In_1324);
nor U3290 (N_3290,In_1083,In_994);
nand U3291 (N_3291,In_620,In_1453);
nor U3292 (N_3292,In_613,In_1062);
or U3293 (N_3293,In_688,In_1194);
or U3294 (N_3294,In_128,In_1347);
xnor U3295 (N_3295,In_1048,In_1488);
or U3296 (N_3296,In_840,In_489);
nor U3297 (N_3297,In_1279,In_309);
or U3298 (N_3298,In_142,In_661);
or U3299 (N_3299,In_633,In_1424);
xor U3300 (N_3300,In_1407,In_307);
or U3301 (N_3301,In_579,In_517);
nor U3302 (N_3302,In_687,In_1252);
xor U3303 (N_3303,In_1476,In_479);
nor U3304 (N_3304,In_522,In_777);
nand U3305 (N_3305,In_1148,In_1013);
or U3306 (N_3306,In_334,In_745);
xor U3307 (N_3307,In_163,In_1293);
nor U3308 (N_3308,In_462,In_1393);
and U3309 (N_3309,In_1055,In_60);
nor U3310 (N_3310,In_715,In_335);
and U3311 (N_3311,In_1431,In_638);
nand U3312 (N_3312,In_1492,In_1400);
nor U3313 (N_3313,In_814,In_834);
xnor U3314 (N_3314,In_130,In_393);
nor U3315 (N_3315,In_616,In_279);
or U3316 (N_3316,In_161,In_1214);
or U3317 (N_3317,In_1227,In_884);
or U3318 (N_3318,In_802,In_724);
and U3319 (N_3319,In_474,In_269);
and U3320 (N_3320,In_1298,In_1254);
nor U3321 (N_3321,In_536,In_648);
or U3322 (N_3322,In_720,In_1477);
and U3323 (N_3323,In_183,In_46);
nand U3324 (N_3324,In_363,In_1240);
xor U3325 (N_3325,In_148,In_1178);
nor U3326 (N_3326,In_931,In_514);
and U3327 (N_3327,In_1052,In_691);
nand U3328 (N_3328,In_712,In_165);
or U3329 (N_3329,In_155,In_1223);
nand U3330 (N_3330,In_1320,In_136);
or U3331 (N_3331,In_301,In_615);
xnor U3332 (N_3332,In_1361,In_1459);
and U3333 (N_3333,In_1408,In_572);
and U3334 (N_3334,In_770,In_1378);
or U3335 (N_3335,In_761,In_478);
xnor U3336 (N_3336,In_738,In_1039);
or U3337 (N_3337,In_1245,In_178);
xnor U3338 (N_3338,In_379,In_485);
or U3339 (N_3339,In_1471,In_104);
xnor U3340 (N_3340,In_1202,In_874);
or U3341 (N_3341,In_1131,In_1317);
or U3342 (N_3342,In_271,In_898);
xor U3343 (N_3343,In_213,In_713);
and U3344 (N_3344,In_1274,In_107);
or U3345 (N_3345,In_1182,In_280);
nand U3346 (N_3346,In_6,In_774);
and U3347 (N_3347,In_925,In_1428);
nand U3348 (N_3348,In_1199,In_1078);
or U3349 (N_3349,In_1062,In_32);
or U3350 (N_3350,In_1054,In_474);
or U3351 (N_3351,In_789,In_1338);
xnor U3352 (N_3352,In_932,In_117);
nand U3353 (N_3353,In_1038,In_1309);
or U3354 (N_3354,In_632,In_339);
xnor U3355 (N_3355,In_110,In_872);
nor U3356 (N_3356,In_260,In_340);
xor U3357 (N_3357,In_922,In_1473);
and U3358 (N_3358,In_446,In_748);
and U3359 (N_3359,In_880,In_126);
and U3360 (N_3360,In_1260,In_643);
or U3361 (N_3361,In_154,In_748);
xnor U3362 (N_3362,In_129,In_275);
xnor U3363 (N_3363,In_977,In_1009);
and U3364 (N_3364,In_66,In_884);
nor U3365 (N_3365,In_846,In_600);
or U3366 (N_3366,In_425,In_206);
nor U3367 (N_3367,In_72,In_1418);
and U3368 (N_3368,In_587,In_1119);
or U3369 (N_3369,In_957,In_1026);
or U3370 (N_3370,In_297,In_774);
and U3371 (N_3371,In_382,In_32);
or U3372 (N_3372,In_1447,In_1410);
and U3373 (N_3373,In_412,In_445);
xnor U3374 (N_3374,In_1395,In_1118);
xor U3375 (N_3375,In_903,In_24);
xor U3376 (N_3376,In_67,In_522);
nor U3377 (N_3377,In_524,In_1075);
nor U3378 (N_3378,In_1325,In_1234);
and U3379 (N_3379,In_994,In_639);
nor U3380 (N_3380,In_815,In_1364);
nor U3381 (N_3381,In_1187,In_275);
xor U3382 (N_3382,In_127,In_1128);
or U3383 (N_3383,In_1237,In_352);
nor U3384 (N_3384,In_1253,In_174);
and U3385 (N_3385,In_1386,In_576);
nand U3386 (N_3386,In_719,In_769);
nand U3387 (N_3387,In_1245,In_1150);
nand U3388 (N_3388,In_848,In_1482);
or U3389 (N_3389,In_1483,In_1149);
nand U3390 (N_3390,In_566,In_1421);
and U3391 (N_3391,In_811,In_1272);
nand U3392 (N_3392,In_175,In_727);
or U3393 (N_3393,In_440,In_724);
xnor U3394 (N_3394,In_1302,In_174);
nand U3395 (N_3395,In_501,In_512);
nand U3396 (N_3396,In_535,In_858);
or U3397 (N_3397,In_911,In_360);
nand U3398 (N_3398,In_1169,In_181);
nor U3399 (N_3399,In_569,In_265);
nor U3400 (N_3400,In_1029,In_1471);
nand U3401 (N_3401,In_311,In_651);
and U3402 (N_3402,In_1008,In_990);
nor U3403 (N_3403,In_40,In_1178);
nand U3404 (N_3404,In_183,In_549);
and U3405 (N_3405,In_109,In_718);
nor U3406 (N_3406,In_143,In_1447);
nand U3407 (N_3407,In_1150,In_402);
or U3408 (N_3408,In_979,In_347);
xnor U3409 (N_3409,In_1086,In_155);
nand U3410 (N_3410,In_178,In_1319);
nand U3411 (N_3411,In_904,In_1316);
nand U3412 (N_3412,In_1491,In_1079);
nand U3413 (N_3413,In_49,In_174);
nand U3414 (N_3414,In_943,In_371);
nand U3415 (N_3415,In_1472,In_1368);
and U3416 (N_3416,In_263,In_999);
or U3417 (N_3417,In_681,In_1200);
nor U3418 (N_3418,In_479,In_66);
xor U3419 (N_3419,In_879,In_131);
xnor U3420 (N_3420,In_1020,In_1424);
or U3421 (N_3421,In_512,In_172);
xnor U3422 (N_3422,In_48,In_1116);
and U3423 (N_3423,In_360,In_1333);
xor U3424 (N_3424,In_1491,In_652);
xor U3425 (N_3425,In_155,In_874);
xnor U3426 (N_3426,In_1294,In_992);
nand U3427 (N_3427,In_716,In_1103);
nor U3428 (N_3428,In_1058,In_869);
nor U3429 (N_3429,In_1300,In_1279);
nor U3430 (N_3430,In_1374,In_1181);
nor U3431 (N_3431,In_791,In_947);
nand U3432 (N_3432,In_81,In_133);
nor U3433 (N_3433,In_1136,In_757);
and U3434 (N_3434,In_1018,In_1071);
nand U3435 (N_3435,In_842,In_651);
or U3436 (N_3436,In_355,In_312);
nand U3437 (N_3437,In_199,In_1413);
xor U3438 (N_3438,In_1116,In_142);
nor U3439 (N_3439,In_1401,In_906);
and U3440 (N_3440,In_547,In_1013);
and U3441 (N_3441,In_103,In_647);
nor U3442 (N_3442,In_951,In_125);
nor U3443 (N_3443,In_1213,In_83);
or U3444 (N_3444,In_252,In_1394);
xor U3445 (N_3445,In_82,In_437);
nand U3446 (N_3446,In_1383,In_31);
and U3447 (N_3447,In_1294,In_102);
nand U3448 (N_3448,In_688,In_1016);
nand U3449 (N_3449,In_733,In_968);
nand U3450 (N_3450,In_849,In_737);
nor U3451 (N_3451,In_140,In_1449);
or U3452 (N_3452,In_295,In_1399);
xnor U3453 (N_3453,In_1366,In_1167);
nor U3454 (N_3454,In_1326,In_421);
or U3455 (N_3455,In_1070,In_473);
nor U3456 (N_3456,In_373,In_692);
xor U3457 (N_3457,In_1086,In_814);
or U3458 (N_3458,In_655,In_656);
or U3459 (N_3459,In_289,In_678);
and U3460 (N_3460,In_612,In_410);
or U3461 (N_3461,In_1113,In_528);
nor U3462 (N_3462,In_1347,In_910);
nor U3463 (N_3463,In_125,In_87);
and U3464 (N_3464,In_1325,In_1449);
nor U3465 (N_3465,In_352,In_396);
nor U3466 (N_3466,In_1065,In_1164);
or U3467 (N_3467,In_788,In_1119);
nor U3468 (N_3468,In_67,In_27);
and U3469 (N_3469,In_382,In_1021);
and U3470 (N_3470,In_154,In_135);
xor U3471 (N_3471,In_385,In_172);
xnor U3472 (N_3472,In_1142,In_641);
nor U3473 (N_3473,In_313,In_833);
or U3474 (N_3474,In_596,In_1129);
and U3475 (N_3475,In_154,In_709);
nor U3476 (N_3476,In_169,In_925);
nor U3477 (N_3477,In_1095,In_485);
or U3478 (N_3478,In_1405,In_106);
and U3479 (N_3479,In_431,In_1480);
and U3480 (N_3480,In_1059,In_73);
nand U3481 (N_3481,In_726,In_420);
nand U3482 (N_3482,In_177,In_948);
and U3483 (N_3483,In_854,In_187);
xnor U3484 (N_3484,In_538,In_1431);
nor U3485 (N_3485,In_1394,In_1041);
nor U3486 (N_3486,In_963,In_504);
nand U3487 (N_3487,In_671,In_452);
or U3488 (N_3488,In_53,In_83);
nor U3489 (N_3489,In_1368,In_584);
and U3490 (N_3490,In_369,In_425);
nand U3491 (N_3491,In_502,In_1467);
and U3492 (N_3492,In_293,In_1238);
or U3493 (N_3493,In_1475,In_1132);
and U3494 (N_3494,In_289,In_1334);
xor U3495 (N_3495,In_1479,In_493);
or U3496 (N_3496,In_1045,In_1244);
and U3497 (N_3497,In_326,In_868);
and U3498 (N_3498,In_1403,In_120);
nand U3499 (N_3499,In_1292,In_822);
and U3500 (N_3500,In_744,In_140);
nand U3501 (N_3501,In_466,In_1410);
nand U3502 (N_3502,In_1248,In_707);
xor U3503 (N_3503,In_419,In_614);
or U3504 (N_3504,In_1360,In_132);
nor U3505 (N_3505,In_547,In_133);
nor U3506 (N_3506,In_436,In_1174);
and U3507 (N_3507,In_474,In_1051);
nand U3508 (N_3508,In_493,In_79);
xor U3509 (N_3509,In_671,In_813);
nor U3510 (N_3510,In_158,In_962);
xnor U3511 (N_3511,In_432,In_55);
or U3512 (N_3512,In_830,In_1294);
nand U3513 (N_3513,In_339,In_1455);
xor U3514 (N_3514,In_1189,In_405);
xor U3515 (N_3515,In_741,In_571);
or U3516 (N_3516,In_279,In_1438);
nand U3517 (N_3517,In_129,In_1212);
nand U3518 (N_3518,In_1386,In_806);
nor U3519 (N_3519,In_798,In_534);
and U3520 (N_3520,In_548,In_1359);
nand U3521 (N_3521,In_1200,In_1026);
nor U3522 (N_3522,In_486,In_1340);
nand U3523 (N_3523,In_1331,In_1117);
or U3524 (N_3524,In_250,In_115);
nor U3525 (N_3525,In_632,In_814);
xnor U3526 (N_3526,In_320,In_1161);
or U3527 (N_3527,In_1255,In_84);
xnor U3528 (N_3528,In_356,In_779);
and U3529 (N_3529,In_770,In_829);
and U3530 (N_3530,In_1252,In_67);
and U3531 (N_3531,In_1313,In_807);
nand U3532 (N_3532,In_418,In_1205);
nand U3533 (N_3533,In_353,In_623);
nand U3534 (N_3534,In_357,In_968);
or U3535 (N_3535,In_56,In_479);
nor U3536 (N_3536,In_214,In_1496);
and U3537 (N_3537,In_720,In_1481);
and U3538 (N_3538,In_268,In_1400);
xor U3539 (N_3539,In_17,In_898);
or U3540 (N_3540,In_1429,In_357);
nand U3541 (N_3541,In_177,In_494);
or U3542 (N_3542,In_1390,In_1081);
and U3543 (N_3543,In_1257,In_784);
xor U3544 (N_3544,In_1110,In_253);
nor U3545 (N_3545,In_1070,In_910);
nand U3546 (N_3546,In_377,In_964);
and U3547 (N_3547,In_1485,In_646);
nand U3548 (N_3548,In_1112,In_91);
or U3549 (N_3549,In_65,In_489);
or U3550 (N_3550,In_1448,In_99);
or U3551 (N_3551,In_1045,In_1145);
nand U3552 (N_3552,In_907,In_196);
and U3553 (N_3553,In_716,In_1150);
and U3554 (N_3554,In_1393,In_1092);
and U3555 (N_3555,In_735,In_221);
xor U3556 (N_3556,In_954,In_327);
and U3557 (N_3557,In_1393,In_826);
nand U3558 (N_3558,In_338,In_737);
xnor U3559 (N_3559,In_1435,In_541);
or U3560 (N_3560,In_621,In_291);
and U3561 (N_3561,In_471,In_907);
and U3562 (N_3562,In_1245,In_511);
and U3563 (N_3563,In_524,In_545);
nand U3564 (N_3564,In_1144,In_575);
xor U3565 (N_3565,In_352,In_1083);
xor U3566 (N_3566,In_225,In_7);
nand U3567 (N_3567,In_1165,In_633);
xnor U3568 (N_3568,In_1201,In_557);
nor U3569 (N_3569,In_1023,In_900);
nand U3570 (N_3570,In_335,In_640);
and U3571 (N_3571,In_1286,In_480);
or U3572 (N_3572,In_146,In_3);
nor U3573 (N_3573,In_129,In_1258);
nor U3574 (N_3574,In_337,In_1048);
nand U3575 (N_3575,In_895,In_1363);
or U3576 (N_3576,In_287,In_795);
and U3577 (N_3577,In_440,In_1388);
xnor U3578 (N_3578,In_521,In_258);
and U3579 (N_3579,In_968,In_227);
or U3580 (N_3580,In_92,In_1146);
and U3581 (N_3581,In_1461,In_596);
or U3582 (N_3582,In_187,In_990);
nand U3583 (N_3583,In_1168,In_1114);
or U3584 (N_3584,In_1486,In_472);
and U3585 (N_3585,In_871,In_288);
nand U3586 (N_3586,In_1319,In_929);
nor U3587 (N_3587,In_334,In_1232);
nor U3588 (N_3588,In_1293,In_213);
or U3589 (N_3589,In_603,In_408);
nand U3590 (N_3590,In_1459,In_85);
xnor U3591 (N_3591,In_227,In_1462);
or U3592 (N_3592,In_1211,In_1020);
nor U3593 (N_3593,In_309,In_1475);
and U3594 (N_3594,In_625,In_1454);
xnor U3595 (N_3595,In_1341,In_488);
and U3596 (N_3596,In_509,In_337);
and U3597 (N_3597,In_1299,In_26);
and U3598 (N_3598,In_176,In_1107);
nand U3599 (N_3599,In_953,In_1320);
nor U3600 (N_3600,In_552,In_369);
xor U3601 (N_3601,In_515,In_143);
and U3602 (N_3602,In_149,In_888);
or U3603 (N_3603,In_571,In_451);
xnor U3604 (N_3604,In_1275,In_529);
nand U3605 (N_3605,In_679,In_391);
nand U3606 (N_3606,In_1293,In_254);
nand U3607 (N_3607,In_1357,In_1154);
and U3608 (N_3608,In_1203,In_968);
or U3609 (N_3609,In_647,In_1018);
nor U3610 (N_3610,In_147,In_588);
nand U3611 (N_3611,In_1027,In_544);
and U3612 (N_3612,In_1093,In_1300);
nand U3613 (N_3613,In_494,In_31);
or U3614 (N_3614,In_1019,In_160);
nor U3615 (N_3615,In_833,In_1366);
nand U3616 (N_3616,In_417,In_376);
nand U3617 (N_3617,In_863,In_210);
nor U3618 (N_3618,In_878,In_787);
or U3619 (N_3619,In_774,In_1288);
xnor U3620 (N_3620,In_723,In_597);
nor U3621 (N_3621,In_998,In_1206);
nand U3622 (N_3622,In_424,In_225);
nand U3623 (N_3623,In_1166,In_1101);
nand U3624 (N_3624,In_994,In_171);
nor U3625 (N_3625,In_590,In_170);
nand U3626 (N_3626,In_1419,In_610);
or U3627 (N_3627,In_617,In_439);
nor U3628 (N_3628,In_1399,In_1362);
xor U3629 (N_3629,In_761,In_1242);
xnor U3630 (N_3630,In_1236,In_1271);
xor U3631 (N_3631,In_1182,In_597);
or U3632 (N_3632,In_1021,In_678);
nand U3633 (N_3633,In_589,In_1219);
and U3634 (N_3634,In_703,In_1034);
or U3635 (N_3635,In_198,In_442);
and U3636 (N_3636,In_994,In_667);
nor U3637 (N_3637,In_1030,In_583);
or U3638 (N_3638,In_876,In_364);
nor U3639 (N_3639,In_547,In_1234);
nor U3640 (N_3640,In_502,In_979);
nor U3641 (N_3641,In_904,In_800);
and U3642 (N_3642,In_1490,In_1268);
nand U3643 (N_3643,In_879,In_761);
xor U3644 (N_3644,In_76,In_1149);
xor U3645 (N_3645,In_616,In_271);
nor U3646 (N_3646,In_317,In_1019);
xnor U3647 (N_3647,In_1074,In_216);
and U3648 (N_3648,In_1090,In_214);
and U3649 (N_3649,In_316,In_672);
nor U3650 (N_3650,In_1012,In_421);
or U3651 (N_3651,In_844,In_611);
xnor U3652 (N_3652,In_267,In_685);
and U3653 (N_3653,In_764,In_613);
or U3654 (N_3654,In_1474,In_135);
or U3655 (N_3655,In_371,In_704);
or U3656 (N_3656,In_803,In_669);
and U3657 (N_3657,In_405,In_458);
nor U3658 (N_3658,In_894,In_599);
and U3659 (N_3659,In_1020,In_996);
or U3660 (N_3660,In_208,In_115);
nor U3661 (N_3661,In_1151,In_1368);
and U3662 (N_3662,In_340,In_454);
xor U3663 (N_3663,In_592,In_353);
nor U3664 (N_3664,In_1423,In_1439);
nand U3665 (N_3665,In_303,In_1122);
nor U3666 (N_3666,In_791,In_904);
xnor U3667 (N_3667,In_387,In_316);
or U3668 (N_3668,In_114,In_1499);
nor U3669 (N_3669,In_682,In_659);
xor U3670 (N_3670,In_892,In_432);
or U3671 (N_3671,In_798,In_892);
nand U3672 (N_3672,In_922,In_350);
xor U3673 (N_3673,In_264,In_513);
nor U3674 (N_3674,In_1252,In_57);
nor U3675 (N_3675,In_1196,In_747);
nor U3676 (N_3676,In_958,In_674);
xor U3677 (N_3677,In_18,In_1313);
nor U3678 (N_3678,In_295,In_421);
nor U3679 (N_3679,In_462,In_560);
nor U3680 (N_3680,In_286,In_105);
nor U3681 (N_3681,In_1024,In_21);
or U3682 (N_3682,In_1364,In_1037);
xor U3683 (N_3683,In_1228,In_273);
or U3684 (N_3684,In_1434,In_1121);
or U3685 (N_3685,In_1161,In_1403);
and U3686 (N_3686,In_233,In_253);
or U3687 (N_3687,In_177,In_1105);
and U3688 (N_3688,In_799,In_243);
nand U3689 (N_3689,In_924,In_61);
nand U3690 (N_3690,In_1386,In_487);
xor U3691 (N_3691,In_637,In_108);
nand U3692 (N_3692,In_843,In_62);
nor U3693 (N_3693,In_1374,In_73);
or U3694 (N_3694,In_880,In_854);
or U3695 (N_3695,In_146,In_62);
and U3696 (N_3696,In_140,In_1212);
nand U3697 (N_3697,In_1051,In_801);
nor U3698 (N_3698,In_258,In_910);
or U3699 (N_3699,In_229,In_982);
and U3700 (N_3700,In_926,In_1418);
or U3701 (N_3701,In_1049,In_787);
nor U3702 (N_3702,In_1463,In_601);
nand U3703 (N_3703,In_233,In_696);
xor U3704 (N_3704,In_497,In_426);
nand U3705 (N_3705,In_586,In_1184);
xnor U3706 (N_3706,In_726,In_1124);
nor U3707 (N_3707,In_554,In_908);
nand U3708 (N_3708,In_974,In_228);
nor U3709 (N_3709,In_204,In_1104);
or U3710 (N_3710,In_684,In_671);
nand U3711 (N_3711,In_597,In_528);
nand U3712 (N_3712,In_386,In_1391);
nor U3713 (N_3713,In_245,In_799);
and U3714 (N_3714,In_147,In_10);
nand U3715 (N_3715,In_404,In_604);
or U3716 (N_3716,In_329,In_301);
nor U3717 (N_3717,In_897,In_1248);
and U3718 (N_3718,In_436,In_802);
and U3719 (N_3719,In_730,In_963);
nor U3720 (N_3720,In_550,In_1335);
xor U3721 (N_3721,In_1334,In_842);
and U3722 (N_3722,In_1215,In_518);
xor U3723 (N_3723,In_805,In_741);
nor U3724 (N_3724,In_1019,In_1237);
nand U3725 (N_3725,In_926,In_945);
or U3726 (N_3726,In_284,In_323);
or U3727 (N_3727,In_1024,In_378);
xnor U3728 (N_3728,In_1110,In_1375);
and U3729 (N_3729,In_851,In_1393);
and U3730 (N_3730,In_473,In_783);
or U3731 (N_3731,In_947,In_31);
or U3732 (N_3732,In_1184,In_846);
and U3733 (N_3733,In_639,In_656);
nand U3734 (N_3734,In_322,In_785);
nand U3735 (N_3735,In_1174,In_986);
or U3736 (N_3736,In_901,In_1015);
xnor U3737 (N_3737,In_1165,In_155);
nor U3738 (N_3738,In_336,In_299);
xor U3739 (N_3739,In_537,In_860);
and U3740 (N_3740,In_25,In_893);
or U3741 (N_3741,In_422,In_25);
xor U3742 (N_3742,In_836,In_613);
nor U3743 (N_3743,In_77,In_468);
nand U3744 (N_3744,In_284,In_307);
nand U3745 (N_3745,In_400,In_722);
nand U3746 (N_3746,In_883,In_10);
and U3747 (N_3747,In_1408,In_306);
nor U3748 (N_3748,In_766,In_473);
and U3749 (N_3749,In_563,In_91);
nor U3750 (N_3750,In_1030,In_611);
and U3751 (N_3751,In_875,In_1187);
xnor U3752 (N_3752,In_110,In_873);
xnor U3753 (N_3753,In_195,In_491);
or U3754 (N_3754,In_213,In_118);
and U3755 (N_3755,In_1168,In_497);
or U3756 (N_3756,In_78,In_911);
or U3757 (N_3757,In_1487,In_1302);
xor U3758 (N_3758,In_1015,In_91);
or U3759 (N_3759,In_1348,In_365);
and U3760 (N_3760,In_289,In_1017);
and U3761 (N_3761,In_1186,In_232);
nand U3762 (N_3762,In_1342,In_1034);
nor U3763 (N_3763,In_973,In_81);
nand U3764 (N_3764,In_196,In_1417);
nor U3765 (N_3765,In_631,In_1375);
and U3766 (N_3766,In_1177,In_143);
nor U3767 (N_3767,In_1268,In_988);
or U3768 (N_3768,In_1381,In_210);
or U3769 (N_3769,In_541,In_459);
xor U3770 (N_3770,In_1497,In_1090);
nor U3771 (N_3771,In_992,In_886);
or U3772 (N_3772,In_83,In_1192);
and U3773 (N_3773,In_1108,In_632);
and U3774 (N_3774,In_823,In_884);
xor U3775 (N_3775,In_323,In_151);
nor U3776 (N_3776,In_961,In_147);
or U3777 (N_3777,In_1490,In_42);
nor U3778 (N_3778,In_644,In_857);
nand U3779 (N_3779,In_802,In_1279);
nand U3780 (N_3780,In_762,In_549);
nor U3781 (N_3781,In_17,In_1334);
nand U3782 (N_3782,In_1229,In_133);
nand U3783 (N_3783,In_908,In_1238);
or U3784 (N_3784,In_561,In_135);
nor U3785 (N_3785,In_535,In_784);
or U3786 (N_3786,In_541,In_1225);
or U3787 (N_3787,In_922,In_472);
xnor U3788 (N_3788,In_1117,In_1398);
or U3789 (N_3789,In_869,In_952);
and U3790 (N_3790,In_222,In_851);
xor U3791 (N_3791,In_943,In_1282);
or U3792 (N_3792,In_593,In_895);
nand U3793 (N_3793,In_1006,In_873);
nor U3794 (N_3794,In_881,In_578);
and U3795 (N_3795,In_784,In_191);
nand U3796 (N_3796,In_809,In_753);
nand U3797 (N_3797,In_780,In_1375);
xnor U3798 (N_3798,In_390,In_1006);
xor U3799 (N_3799,In_1036,In_1290);
or U3800 (N_3800,In_582,In_700);
nand U3801 (N_3801,In_317,In_80);
nand U3802 (N_3802,In_279,In_418);
xor U3803 (N_3803,In_933,In_1196);
or U3804 (N_3804,In_750,In_1205);
or U3805 (N_3805,In_447,In_459);
xor U3806 (N_3806,In_1180,In_701);
xnor U3807 (N_3807,In_413,In_1314);
nor U3808 (N_3808,In_1374,In_674);
nand U3809 (N_3809,In_54,In_259);
nand U3810 (N_3810,In_1258,In_571);
or U3811 (N_3811,In_428,In_1293);
and U3812 (N_3812,In_62,In_1207);
or U3813 (N_3813,In_913,In_1436);
xnor U3814 (N_3814,In_83,In_17);
nand U3815 (N_3815,In_1138,In_238);
and U3816 (N_3816,In_916,In_647);
nand U3817 (N_3817,In_534,In_575);
xnor U3818 (N_3818,In_1224,In_360);
and U3819 (N_3819,In_115,In_1365);
nor U3820 (N_3820,In_746,In_58);
or U3821 (N_3821,In_645,In_846);
xnor U3822 (N_3822,In_174,In_665);
nor U3823 (N_3823,In_1105,In_591);
nor U3824 (N_3824,In_473,In_776);
and U3825 (N_3825,In_104,In_1314);
xor U3826 (N_3826,In_295,In_1314);
nand U3827 (N_3827,In_629,In_1461);
nand U3828 (N_3828,In_258,In_1469);
xor U3829 (N_3829,In_777,In_675);
xnor U3830 (N_3830,In_383,In_909);
and U3831 (N_3831,In_920,In_497);
and U3832 (N_3832,In_729,In_306);
nor U3833 (N_3833,In_1353,In_648);
and U3834 (N_3834,In_420,In_444);
nor U3835 (N_3835,In_215,In_47);
or U3836 (N_3836,In_698,In_1261);
nand U3837 (N_3837,In_594,In_1130);
nand U3838 (N_3838,In_382,In_1463);
xnor U3839 (N_3839,In_615,In_178);
nor U3840 (N_3840,In_575,In_564);
nand U3841 (N_3841,In_1283,In_1083);
nor U3842 (N_3842,In_323,In_929);
xnor U3843 (N_3843,In_618,In_175);
nor U3844 (N_3844,In_1170,In_577);
nor U3845 (N_3845,In_1091,In_434);
nor U3846 (N_3846,In_472,In_825);
or U3847 (N_3847,In_811,In_709);
or U3848 (N_3848,In_160,In_940);
xor U3849 (N_3849,In_877,In_1132);
nand U3850 (N_3850,In_245,In_626);
nor U3851 (N_3851,In_104,In_1293);
xor U3852 (N_3852,In_1312,In_847);
and U3853 (N_3853,In_170,In_235);
or U3854 (N_3854,In_600,In_1261);
nand U3855 (N_3855,In_1351,In_1159);
nor U3856 (N_3856,In_1320,In_128);
xnor U3857 (N_3857,In_1111,In_1189);
xor U3858 (N_3858,In_1264,In_1464);
nor U3859 (N_3859,In_760,In_832);
xor U3860 (N_3860,In_969,In_3);
nand U3861 (N_3861,In_1089,In_153);
and U3862 (N_3862,In_555,In_505);
nand U3863 (N_3863,In_537,In_411);
and U3864 (N_3864,In_149,In_3);
nor U3865 (N_3865,In_1243,In_612);
nor U3866 (N_3866,In_298,In_899);
and U3867 (N_3867,In_235,In_413);
nor U3868 (N_3868,In_591,In_559);
xor U3869 (N_3869,In_890,In_604);
nand U3870 (N_3870,In_45,In_200);
xor U3871 (N_3871,In_186,In_1102);
nor U3872 (N_3872,In_1314,In_1311);
nor U3873 (N_3873,In_530,In_241);
and U3874 (N_3874,In_12,In_1454);
nand U3875 (N_3875,In_352,In_1040);
and U3876 (N_3876,In_750,In_1348);
xnor U3877 (N_3877,In_1364,In_1114);
or U3878 (N_3878,In_1336,In_1280);
nor U3879 (N_3879,In_1105,In_80);
nand U3880 (N_3880,In_217,In_1364);
and U3881 (N_3881,In_1275,In_749);
and U3882 (N_3882,In_722,In_191);
xnor U3883 (N_3883,In_1347,In_711);
or U3884 (N_3884,In_458,In_445);
and U3885 (N_3885,In_806,In_1078);
or U3886 (N_3886,In_1237,In_981);
xnor U3887 (N_3887,In_940,In_1361);
xor U3888 (N_3888,In_622,In_3);
xnor U3889 (N_3889,In_1253,In_1294);
nor U3890 (N_3890,In_137,In_162);
xnor U3891 (N_3891,In_1429,In_1055);
nor U3892 (N_3892,In_678,In_274);
nand U3893 (N_3893,In_1457,In_924);
xnor U3894 (N_3894,In_1145,In_75);
nor U3895 (N_3895,In_334,In_1470);
or U3896 (N_3896,In_464,In_700);
nand U3897 (N_3897,In_450,In_197);
and U3898 (N_3898,In_1006,In_1477);
nand U3899 (N_3899,In_966,In_213);
and U3900 (N_3900,In_782,In_929);
or U3901 (N_3901,In_1232,In_819);
and U3902 (N_3902,In_56,In_427);
or U3903 (N_3903,In_781,In_685);
nor U3904 (N_3904,In_1192,In_264);
nor U3905 (N_3905,In_1008,In_166);
nand U3906 (N_3906,In_448,In_536);
nor U3907 (N_3907,In_889,In_1450);
xor U3908 (N_3908,In_22,In_1249);
nand U3909 (N_3909,In_179,In_212);
nor U3910 (N_3910,In_7,In_460);
and U3911 (N_3911,In_789,In_63);
xor U3912 (N_3912,In_626,In_259);
nor U3913 (N_3913,In_1359,In_712);
nor U3914 (N_3914,In_1235,In_1467);
and U3915 (N_3915,In_49,In_1469);
nand U3916 (N_3916,In_1383,In_678);
nand U3917 (N_3917,In_268,In_1378);
or U3918 (N_3918,In_983,In_441);
nand U3919 (N_3919,In_597,In_982);
and U3920 (N_3920,In_221,In_955);
xor U3921 (N_3921,In_194,In_72);
and U3922 (N_3922,In_1140,In_59);
or U3923 (N_3923,In_201,In_970);
and U3924 (N_3924,In_1062,In_1476);
nor U3925 (N_3925,In_1031,In_848);
nor U3926 (N_3926,In_1198,In_1151);
or U3927 (N_3927,In_1148,In_906);
or U3928 (N_3928,In_597,In_128);
xor U3929 (N_3929,In_391,In_1323);
nand U3930 (N_3930,In_1362,In_504);
or U3931 (N_3931,In_1043,In_66);
xnor U3932 (N_3932,In_1117,In_46);
nand U3933 (N_3933,In_187,In_542);
nor U3934 (N_3934,In_1208,In_11);
nand U3935 (N_3935,In_1407,In_1014);
nor U3936 (N_3936,In_1360,In_21);
and U3937 (N_3937,In_993,In_379);
nand U3938 (N_3938,In_137,In_1226);
xor U3939 (N_3939,In_474,In_1289);
nor U3940 (N_3940,In_1315,In_880);
and U3941 (N_3941,In_1247,In_951);
or U3942 (N_3942,In_1168,In_763);
nand U3943 (N_3943,In_21,In_246);
and U3944 (N_3944,In_890,In_1226);
nand U3945 (N_3945,In_1218,In_708);
nor U3946 (N_3946,In_364,In_140);
nor U3947 (N_3947,In_22,In_815);
or U3948 (N_3948,In_1359,In_615);
xnor U3949 (N_3949,In_44,In_1278);
or U3950 (N_3950,In_371,In_304);
nor U3951 (N_3951,In_1168,In_827);
xor U3952 (N_3952,In_860,In_897);
and U3953 (N_3953,In_1147,In_161);
nor U3954 (N_3954,In_97,In_1033);
and U3955 (N_3955,In_1175,In_1092);
and U3956 (N_3956,In_144,In_1349);
nor U3957 (N_3957,In_1442,In_448);
nor U3958 (N_3958,In_193,In_1325);
or U3959 (N_3959,In_273,In_278);
nand U3960 (N_3960,In_284,In_26);
and U3961 (N_3961,In_1398,In_611);
xnor U3962 (N_3962,In_519,In_1348);
nor U3963 (N_3963,In_1335,In_606);
xnor U3964 (N_3964,In_239,In_1192);
and U3965 (N_3965,In_1097,In_1363);
or U3966 (N_3966,In_357,In_123);
nor U3967 (N_3967,In_821,In_867);
nand U3968 (N_3968,In_80,In_176);
xor U3969 (N_3969,In_907,In_381);
xnor U3970 (N_3970,In_1100,In_1261);
xor U3971 (N_3971,In_403,In_978);
nand U3972 (N_3972,In_39,In_389);
xnor U3973 (N_3973,In_383,In_77);
nor U3974 (N_3974,In_415,In_1480);
nor U3975 (N_3975,In_831,In_83);
or U3976 (N_3976,In_1377,In_137);
xnor U3977 (N_3977,In_785,In_508);
or U3978 (N_3978,In_661,In_1069);
xnor U3979 (N_3979,In_1455,In_1272);
xor U3980 (N_3980,In_60,In_892);
nand U3981 (N_3981,In_1216,In_1414);
and U3982 (N_3982,In_1248,In_113);
nand U3983 (N_3983,In_1394,In_301);
xor U3984 (N_3984,In_357,In_559);
nand U3985 (N_3985,In_248,In_436);
or U3986 (N_3986,In_331,In_1111);
and U3987 (N_3987,In_1337,In_233);
or U3988 (N_3988,In_195,In_1255);
nand U3989 (N_3989,In_257,In_1237);
xor U3990 (N_3990,In_4,In_89);
or U3991 (N_3991,In_1259,In_1458);
nor U3992 (N_3992,In_1064,In_828);
nor U3993 (N_3993,In_1494,In_959);
nor U3994 (N_3994,In_99,In_517);
or U3995 (N_3995,In_61,In_642);
xor U3996 (N_3996,In_310,In_1213);
nand U3997 (N_3997,In_742,In_183);
xor U3998 (N_3998,In_910,In_765);
nand U3999 (N_3999,In_509,In_1171);
and U4000 (N_4000,In_1020,In_1188);
and U4001 (N_4001,In_262,In_90);
and U4002 (N_4002,In_1434,In_968);
nor U4003 (N_4003,In_211,In_681);
nand U4004 (N_4004,In_422,In_42);
nand U4005 (N_4005,In_916,In_1154);
nand U4006 (N_4006,In_389,In_1473);
nor U4007 (N_4007,In_653,In_511);
nand U4008 (N_4008,In_324,In_230);
xnor U4009 (N_4009,In_907,In_366);
nor U4010 (N_4010,In_588,In_780);
xnor U4011 (N_4011,In_255,In_496);
and U4012 (N_4012,In_210,In_1438);
or U4013 (N_4013,In_1331,In_619);
nand U4014 (N_4014,In_11,In_158);
xnor U4015 (N_4015,In_921,In_273);
nand U4016 (N_4016,In_1400,In_266);
xor U4017 (N_4017,In_1439,In_330);
xnor U4018 (N_4018,In_602,In_1381);
xnor U4019 (N_4019,In_187,In_397);
nand U4020 (N_4020,In_795,In_980);
xor U4021 (N_4021,In_812,In_968);
or U4022 (N_4022,In_556,In_1495);
and U4023 (N_4023,In_529,In_215);
nand U4024 (N_4024,In_524,In_295);
and U4025 (N_4025,In_471,In_1290);
xnor U4026 (N_4026,In_68,In_1023);
xnor U4027 (N_4027,In_1333,In_1075);
nand U4028 (N_4028,In_232,In_943);
and U4029 (N_4029,In_1218,In_1481);
or U4030 (N_4030,In_1471,In_349);
nand U4031 (N_4031,In_10,In_933);
or U4032 (N_4032,In_150,In_1353);
xor U4033 (N_4033,In_936,In_990);
xor U4034 (N_4034,In_857,In_1257);
and U4035 (N_4035,In_718,In_1328);
xor U4036 (N_4036,In_777,In_778);
and U4037 (N_4037,In_359,In_904);
nor U4038 (N_4038,In_878,In_232);
xor U4039 (N_4039,In_842,In_1326);
and U4040 (N_4040,In_439,In_660);
and U4041 (N_4041,In_1220,In_1208);
nand U4042 (N_4042,In_610,In_617);
and U4043 (N_4043,In_671,In_542);
xor U4044 (N_4044,In_1182,In_1407);
nand U4045 (N_4045,In_589,In_322);
xnor U4046 (N_4046,In_953,In_1054);
nand U4047 (N_4047,In_1271,In_1429);
and U4048 (N_4048,In_685,In_1246);
xor U4049 (N_4049,In_927,In_804);
nand U4050 (N_4050,In_1166,In_817);
nand U4051 (N_4051,In_159,In_508);
or U4052 (N_4052,In_514,In_1444);
and U4053 (N_4053,In_673,In_1228);
and U4054 (N_4054,In_141,In_1271);
or U4055 (N_4055,In_365,In_1217);
or U4056 (N_4056,In_243,In_1428);
xnor U4057 (N_4057,In_1147,In_1283);
nor U4058 (N_4058,In_313,In_1176);
nor U4059 (N_4059,In_716,In_1098);
nor U4060 (N_4060,In_618,In_635);
xnor U4061 (N_4061,In_1393,In_296);
and U4062 (N_4062,In_962,In_1111);
and U4063 (N_4063,In_902,In_1002);
xor U4064 (N_4064,In_1045,In_1156);
xor U4065 (N_4065,In_553,In_62);
and U4066 (N_4066,In_1421,In_1258);
xor U4067 (N_4067,In_53,In_508);
nor U4068 (N_4068,In_1165,In_96);
and U4069 (N_4069,In_34,In_1143);
nor U4070 (N_4070,In_535,In_733);
nor U4071 (N_4071,In_964,In_131);
nand U4072 (N_4072,In_591,In_1457);
or U4073 (N_4073,In_906,In_1314);
xnor U4074 (N_4074,In_955,In_1480);
xor U4075 (N_4075,In_940,In_364);
or U4076 (N_4076,In_907,In_553);
and U4077 (N_4077,In_919,In_8);
nand U4078 (N_4078,In_86,In_338);
or U4079 (N_4079,In_194,In_814);
xnor U4080 (N_4080,In_1129,In_1499);
nor U4081 (N_4081,In_730,In_1158);
nor U4082 (N_4082,In_293,In_420);
or U4083 (N_4083,In_1433,In_1268);
and U4084 (N_4084,In_1112,In_1177);
or U4085 (N_4085,In_114,In_1477);
xor U4086 (N_4086,In_518,In_1361);
nand U4087 (N_4087,In_966,In_1145);
xnor U4088 (N_4088,In_569,In_167);
nor U4089 (N_4089,In_306,In_1151);
or U4090 (N_4090,In_480,In_772);
or U4091 (N_4091,In_754,In_474);
xor U4092 (N_4092,In_1234,In_394);
xor U4093 (N_4093,In_1227,In_390);
nor U4094 (N_4094,In_1404,In_35);
nand U4095 (N_4095,In_304,In_1310);
nor U4096 (N_4096,In_523,In_376);
xor U4097 (N_4097,In_676,In_1192);
nand U4098 (N_4098,In_1225,In_1470);
nand U4099 (N_4099,In_348,In_992);
nand U4100 (N_4100,In_414,In_717);
nor U4101 (N_4101,In_1444,In_1452);
nand U4102 (N_4102,In_812,In_667);
nand U4103 (N_4103,In_867,In_1323);
xnor U4104 (N_4104,In_720,In_903);
nor U4105 (N_4105,In_1312,In_1378);
nor U4106 (N_4106,In_562,In_1046);
and U4107 (N_4107,In_944,In_1407);
or U4108 (N_4108,In_846,In_437);
and U4109 (N_4109,In_449,In_127);
xnor U4110 (N_4110,In_738,In_365);
nand U4111 (N_4111,In_840,In_1059);
xor U4112 (N_4112,In_1143,In_402);
xnor U4113 (N_4113,In_190,In_889);
and U4114 (N_4114,In_860,In_932);
and U4115 (N_4115,In_851,In_463);
and U4116 (N_4116,In_159,In_977);
nand U4117 (N_4117,In_1364,In_100);
and U4118 (N_4118,In_1183,In_1052);
or U4119 (N_4119,In_285,In_211);
or U4120 (N_4120,In_665,In_1144);
nor U4121 (N_4121,In_923,In_1153);
nor U4122 (N_4122,In_461,In_1188);
nand U4123 (N_4123,In_452,In_64);
nor U4124 (N_4124,In_1403,In_800);
or U4125 (N_4125,In_1279,In_1059);
nand U4126 (N_4126,In_196,In_237);
nand U4127 (N_4127,In_423,In_508);
or U4128 (N_4128,In_478,In_607);
and U4129 (N_4129,In_1230,In_101);
and U4130 (N_4130,In_500,In_882);
nor U4131 (N_4131,In_544,In_149);
nor U4132 (N_4132,In_604,In_1293);
nand U4133 (N_4133,In_530,In_997);
and U4134 (N_4134,In_980,In_95);
xnor U4135 (N_4135,In_978,In_120);
and U4136 (N_4136,In_126,In_765);
nor U4137 (N_4137,In_686,In_802);
nand U4138 (N_4138,In_1488,In_387);
nand U4139 (N_4139,In_368,In_841);
xor U4140 (N_4140,In_1198,In_1156);
and U4141 (N_4141,In_1428,In_1382);
nand U4142 (N_4142,In_1478,In_1243);
or U4143 (N_4143,In_255,In_451);
nand U4144 (N_4144,In_337,In_915);
and U4145 (N_4145,In_513,In_940);
or U4146 (N_4146,In_477,In_111);
nand U4147 (N_4147,In_1141,In_846);
xnor U4148 (N_4148,In_305,In_534);
and U4149 (N_4149,In_1370,In_1408);
xor U4150 (N_4150,In_453,In_935);
and U4151 (N_4151,In_1481,In_936);
xnor U4152 (N_4152,In_1228,In_473);
nand U4153 (N_4153,In_739,In_1409);
and U4154 (N_4154,In_440,In_770);
nand U4155 (N_4155,In_80,In_1084);
nor U4156 (N_4156,In_1172,In_891);
nor U4157 (N_4157,In_1111,In_666);
nand U4158 (N_4158,In_512,In_1065);
xnor U4159 (N_4159,In_1422,In_642);
nand U4160 (N_4160,In_722,In_769);
nor U4161 (N_4161,In_303,In_1237);
or U4162 (N_4162,In_1487,In_541);
nor U4163 (N_4163,In_1267,In_872);
xnor U4164 (N_4164,In_368,In_1209);
nand U4165 (N_4165,In_1106,In_739);
nor U4166 (N_4166,In_605,In_928);
xor U4167 (N_4167,In_247,In_297);
nor U4168 (N_4168,In_1434,In_315);
nand U4169 (N_4169,In_978,In_926);
nand U4170 (N_4170,In_956,In_408);
xnor U4171 (N_4171,In_93,In_594);
or U4172 (N_4172,In_1030,In_57);
or U4173 (N_4173,In_392,In_764);
or U4174 (N_4174,In_1478,In_920);
and U4175 (N_4175,In_1153,In_1324);
xnor U4176 (N_4176,In_413,In_155);
and U4177 (N_4177,In_997,In_1286);
xor U4178 (N_4178,In_1208,In_521);
and U4179 (N_4179,In_798,In_771);
and U4180 (N_4180,In_20,In_162);
or U4181 (N_4181,In_215,In_1398);
or U4182 (N_4182,In_1354,In_125);
nor U4183 (N_4183,In_976,In_1006);
nor U4184 (N_4184,In_1101,In_1470);
and U4185 (N_4185,In_586,In_107);
nand U4186 (N_4186,In_202,In_623);
or U4187 (N_4187,In_47,In_915);
and U4188 (N_4188,In_1316,In_795);
or U4189 (N_4189,In_353,In_821);
or U4190 (N_4190,In_1126,In_1283);
xnor U4191 (N_4191,In_979,In_297);
or U4192 (N_4192,In_952,In_1088);
or U4193 (N_4193,In_71,In_139);
and U4194 (N_4194,In_1340,In_74);
and U4195 (N_4195,In_924,In_966);
and U4196 (N_4196,In_43,In_1419);
or U4197 (N_4197,In_414,In_441);
xnor U4198 (N_4198,In_633,In_770);
nand U4199 (N_4199,In_1303,In_58);
nor U4200 (N_4200,In_196,In_970);
nand U4201 (N_4201,In_532,In_701);
nand U4202 (N_4202,In_61,In_1069);
nand U4203 (N_4203,In_600,In_920);
xor U4204 (N_4204,In_0,In_326);
nand U4205 (N_4205,In_1086,In_347);
nand U4206 (N_4206,In_1155,In_1013);
and U4207 (N_4207,In_153,In_901);
or U4208 (N_4208,In_1281,In_1208);
and U4209 (N_4209,In_1493,In_323);
or U4210 (N_4210,In_164,In_670);
or U4211 (N_4211,In_1055,In_125);
and U4212 (N_4212,In_811,In_91);
nand U4213 (N_4213,In_944,In_386);
nor U4214 (N_4214,In_157,In_915);
nand U4215 (N_4215,In_79,In_1324);
nand U4216 (N_4216,In_1429,In_162);
nor U4217 (N_4217,In_1059,In_1146);
xor U4218 (N_4218,In_840,In_1040);
or U4219 (N_4219,In_368,In_844);
nand U4220 (N_4220,In_564,In_1105);
nand U4221 (N_4221,In_1118,In_1080);
and U4222 (N_4222,In_1165,In_1154);
nor U4223 (N_4223,In_229,In_71);
or U4224 (N_4224,In_455,In_412);
nor U4225 (N_4225,In_362,In_515);
or U4226 (N_4226,In_1454,In_345);
xor U4227 (N_4227,In_1195,In_1465);
nor U4228 (N_4228,In_1003,In_317);
or U4229 (N_4229,In_314,In_160);
or U4230 (N_4230,In_1054,In_1052);
or U4231 (N_4231,In_184,In_1062);
and U4232 (N_4232,In_802,In_90);
nor U4233 (N_4233,In_208,In_1288);
nand U4234 (N_4234,In_1022,In_909);
nor U4235 (N_4235,In_421,In_201);
nand U4236 (N_4236,In_419,In_1441);
or U4237 (N_4237,In_1133,In_611);
xor U4238 (N_4238,In_60,In_755);
and U4239 (N_4239,In_471,In_1211);
and U4240 (N_4240,In_854,In_532);
nor U4241 (N_4241,In_973,In_6);
or U4242 (N_4242,In_1311,In_273);
xnor U4243 (N_4243,In_958,In_188);
and U4244 (N_4244,In_1183,In_984);
nor U4245 (N_4245,In_252,In_965);
xor U4246 (N_4246,In_826,In_1312);
xnor U4247 (N_4247,In_743,In_603);
nand U4248 (N_4248,In_838,In_583);
nand U4249 (N_4249,In_462,In_872);
or U4250 (N_4250,In_460,In_946);
and U4251 (N_4251,In_856,In_457);
nand U4252 (N_4252,In_1365,In_155);
and U4253 (N_4253,In_525,In_828);
xor U4254 (N_4254,In_1158,In_86);
xor U4255 (N_4255,In_1172,In_25);
nor U4256 (N_4256,In_1014,In_837);
and U4257 (N_4257,In_701,In_1364);
nand U4258 (N_4258,In_974,In_93);
nand U4259 (N_4259,In_746,In_1240);
nor U4260 (N_4260,In_457,In_1171);
or U4261 (N_4261,In_764,In_277);
nand U4262 (N_4262,In_417,In_1413);
nor U4263 (N_4263,In_625,In_443);
or U4264 (N_4264,In_623,In_919);
nor U4265 (N_4265,In_433,In_44);
xor U4266 (N_4266,In_1177,In_634);
xor U4267 (N_4267,In_1064,In_268);
nor U4268 (N_4268,In_404,In_627);
or U4269 (N_4269,In_1,In_623);
nand U4270 (N_4270,In_1351,In_1006);
and U4271 (N_4271,In_586,In_138);
xor U4272 (N_4272,In_1439,In_1044);
nor U4273 (N_4273,In_1093,In_1481);
nor U4274 (N_4274,In_1091,In_1105);
nor U4275 (N_4275,In_43,In_1366);
and U4276 (N_4276,In_1394,In_400);
nand U4277 (N_4277,In_486,In_1163);
and U4278 (N_4278,In_588,In_135);
nor U4279 (N_4279,In_1222,In_1045);
xor U4280 (N_4280,In_1222,In_1047);
or U4281 (N_4281,In_1129,In_268);
xor U4282 (N_4282,In_1414,In_1214);
nand U4283 (N_4283,In_944,In_197);
nand U4284 (N_4284,In_816,In_1420);
and U4285 (N_4285,In_16,In_655);
and U4286 (N_4286,In_746,In_1261);
or U4287 (N_4287,In_1471,In_492);
or U4288 (N_4288,In_126,In_1308);
or U4289 (N_4289,In_1070,In_1066);
or U4290 (N_4290,In_121,In_379);
nor U4291 (N_4291,In_359,In_1004);
or U4292 (N_4292,In_1140,In_285);
nor U4293 (N_4293,In_674,In_355);
nand U4294 (N_4294,In_1109,In_937);
nor U4295 (N_4295,In_691,In_936);
or U4296 (N_4296,In_1174,In_1182);
nor U4297 (N_4297,In_389,In_891);
or U4298 (N_4298,In_1055,In_1127);
xor U4299 (N_4299,In_476,In_1247);
nor U4300 (N_4300,In_265,In_1459);
xor U4301 (N_4301,In_895,In_714);
xor U4302 (N_4302,In_1133,In_1023);
nand U4303 (N_4303,In_0,In_936);
xnor U4304 (N_4304,In_847,In_1113);
nor U4305 (N_4305,In_19,In_1208);
xnor U4306 (N_4306,In_352,In_956);
nand U4307 (N_4307,In_1487,In_0);
or U4308 (N_4308,In_299,In_343);
and U4309 (N_4309,In_299,In_86);
nand U4310 (N_4310,In_185,In_765);
nand U4311 (N_4311,In_687,In_1416);
nand U4312 (N_4312,In_765,In_73);
nand U4313 (N_4313,In_644,In_938);
nor U4314 (N_4314,In_354,In_902);
and U4315 (N_4315,In_357,In_108);
or U4316 (N_4316,In_1212,In_153);
xor U4317 (N_4317,In_147,In_109);
and U4318 (N_4318,In_18,In_1332);
nand U4319 (N_4319,In_965,In_1320);
nor U4320 (N_4320,In_1053,In_450);
and U4321 (N_4321,In_21,In_1077);
xnor U4322 (N_4322,In_1469,In_1348);
xor U4323 (N_4323,In_93,In_869);
nand U4324 (N_4324,In_1254,In_294);
nor U4325 (N_4325,In_638,In_1342);
and U4326 (N_4326,In_1051,In_309);
and U4327 (N_4327,In_928,In_106);
nand U4328 (N_4328,In_1357,In_495);
and U4329 (N_4329,In_585,In_1190);
or U4330 (N_4330,In_109,In_40);
xor U4331 (N_4331,In_1319,In_7);
nor U4332 (N_4332,In_202,In_534);
xnor U4333 (N_4333,In_581,In_1192);
nor U4334 (N_4334,In_1110,In_579);
or U4335 (N_4335,In_1440,In_1277);
nor U4336 (N_4336,In_378,In_1092);
nor U4337 (N_4337,In_630,In_443);
nand U4338 (N_4338,In_51,In_1305);
or U4339 (N_4339,In_1363,In_230);
or U4340 (N_4340,In_475,In_1477);
nand U4341 (N_4341,In_25,In_802);
nand U4342 (N_4342,In_424,In_1243);
and U4343 (N_4343,In_1177,In_1498);
xor U4344 (N_4344,In_123,In_363);
nand U4345 (N_4345,In_256,In_1478);
nor U4346 (N_4346,In_173,In_741);
nor U4347 (N_4347,In_431,In_566);
xnor U4348 (N_4348,In_989,In_1080);
xor U4349 (N_4349,In_650,In_447);
or U4350 (N_4350,In_205,In_773);
nor U4351 (N_4351,In_587,In_811);
xnor U4352 (N_4352,In_834,In_443);
xor U4353 (N_4353,In_1314,In_248);
and U4354 (N_4354,In_901,In_1386);
nor U4355 (N_4355,In_969,In_302);
or U4356 (N_4356,In_237,In_404);
nor U4357 (N_4357,In_615,In_1121);
and U4358 (N_4358,In_905,In_247);
nor U4359 (N_4359,In_511,In_1334);
or U4360 (N_4360,In_955,In_710);
xnor U4361 (N_4361,In_881,In_521);
and U4362 (N_4362,In_774,In_644);
nand U4363 (N_4363,In_1476,In_390);
and U4364 (N_4364,In_1050,In_690);
nand U4365 (N_4365,In_382,In_458);
and U4366 (N_4366,In_437,In_990);
and U4367 (N_4367,In_671,In_885);
and U4368 (N_4368,In_398,In_1032);
nand U4369 (N_4369,In_1358,In_506);
xor U4370 (N_4370,In_903,In_1453);
nor U4371 (N_4371,In_897,In_1103);
xnor U4372 (N_4372,In_850,In_856);
xnor U4373 (N_4373,In_447,In_916);
xnor U4374 (N_4374,In_1162,In_313);
nand U4375 (N_4375,In_1293,In_439);
nor U4376 (N_4376,In_334,In_894);
nand U4377 (N_4377,In_173,In_1293);
or U4378 (N_4378,In_513,In_320);
nor U4379 (N_4379,In_403,In_111);
nand U4380 (N_4380,In_1445,In_861);
or U4381 (N_4381,In_1382,In_295);
and U4382 (N_4382,In_201,In_472);
xor U4383 (N_4383,In_1107,In_627);
nand U4384 (N_4384,In_559,In_1305);
nor U4385 (N_4385,In_1331,In_1384);
nor U4386 (N_4386,In_497,In_164);
xor U4387 (N_4387,In_97,In_1149);
xor U4388 (N_4388,In_281,In_1284);
nand U4389 (N_4389,In_1147,In_9);
xor U4390 (N_4390,In_324,In_75);
nor U4391 (N_4391,In_544,In_1162);
and U4392 (N_4392,In_744,In_1200);
xnor U4393 (N_4393,In_118,In_393);
xor U4394 (N_4394,In_887,In_981);
or U4395 (N_4395,In_1086,In_927);
and U4396 (N_4396,In_61,In_825);
and U4397 (N_4397,In_1386,In_1159);
nor U4398 (N_4398,In_1186,In_673);
xnor U4399 (N_4399,In_1191,In_822);
and U4400 (N_4400,In_514,In_22);
xor U4401 (N_4401,In_1464,In_1396);
or U4402 (N_4402,In_1238,In_342);
nor U4403 (N_4403,In_1466,In_356);
and U4404 (N_4404,In_1155,In_635);
and U4405 (N_4405,In_1374,In_273);
or U4406 (N_4406,In_495,In_777);
and U4407 (N_4407,In_1008,In_467);
or U4408 (N_4408,In_648,In_1156);
xnor U4409 (N_4409,In_91,In_695);
and U4410 (N_4410,In_1483,In_977);
or U4411 (N_4411,In_349,In_941);
xor U4412 (N_4412,In_1039,In_894);
nor U4413 (N_4413,In_758,In_935);
nor U4414 (N_4414,In_1385,In_1101);
nand U4415 (N_4415,In_654,In_393);
xor U4416 (N_4416,In_413,In_813);
xnor U4417 (N_4417,In_424,In_1169);
or U4418 (N_4418,In_351,In_116);
nand U4419 (N_4419,In_597,In_11);
nand U4420 (N_4420,In_727,In_229);
nand U4421 (N_4421,In_640,In_389);
or U4422 (N_4422,In_266,In_186);
or U4423 (N_4423,In_297,In_410);
nand U4424 (N_4424,In_260,In_1185);
or U4425 (N_4425,In_1424,In_770);
and U4426 (N_4426,In_506,In_802);
xnor U4427 (N_4427,In_33,In_923);
xor U4428 (N_4428,In_979,In_807);
and U4429 (N_4429,In_933,In_1258);
or U4430 (N_4430,In_241,In_730);
or U4431 (N_4431,In_1239,In_767);
nand U4432 (N_4432,In_1378,In_358);
and U4433 (N_4433,In_21,In_521);
nand U4434 (N_4434,In_186,In_1360);
and U4435 (N_4435,In_465,In_1198);
or U4436 (N_4436,In_655,In_521);
xor U4437 (N_4437,In_138,In_1388);
nor U4438 (N_4438,In_929,In_1499);
or U4439 (N_4439,In_691,In_28);
xnor U4440 (N_4440,In_1036,In_261);
or U4441 (N_4441,In_543,In_695);
nor U4442 (N_4442,In_40,In_1171);
xnor U4443 (N_4443,In_703,In_865);
nor U4444 (N_4444,In_143,In_1078);
nand U4445 (N_4445,In_992,In_546);
and U4446 (N_4446,In_1145,In_1402);
nand U4447 (N_4447,In_1251,In_1297);
nand U4448 (N_4448,In_1158,In_1033);
xnor U4449 (N_4449,In_121,In_1328);
nand U4450 (N_4450,In_1402,In_645);
and U4451 (N_4451,In_1305,In_552);
and U4452 (N_4452,In_1400,In_318);
nand U4453 (N_4453,In_1114,In_859);
nand U4454 (N_4454,In_81,In_1074);
or U4455 (N_4455,In_673,In_1064);
nand U4456 (N_4456,In_244,In_485);
or U4457 (N_4457,In_716,In_537);
nor U4458 (N_4458,In_577,In_90);
or U4459 (N_4459,In_1357,In_541);
nand U4460 (N_4460,In_1010,In_1225);
or U4461 (N_4461,In_1268,In_1350);
nor U4462 (N_4462,In_730,In_381);
nor U4463 (N_4463,In_503,In_645);
nor U4464 (N_4464,In_35,In_1116);
xor U4465 (N_4465,In_455,In_1225);
or U4466 (N_4466,In_486,In_631);
nand U4467 (N_4467,In_317,In_1448);
xor U4468 (N_4468,In_1494,In_135);
xor U4469 (N_4469,In_1170,In_148);
xor U4470 (N_4470,In_1239,In_1273);
or U4471 (N_4471,In_256,In_299);
xnor U4472 (N_4472,In_653,In_286);
xor U4473 (N_4473,In_1053,In_813);
and U4474 (N_4474,In_630,In_1487);
and U4475 (N_4475,In_625,In_806);
nand U4476 (N_4476,In_155,In_806);
xnor U4477 (N_4477,In_1062,In_382);
or U4478 (N_4478,In_392,In_601);
xor U4479 (N_4479,In_1043,In_471);
and U4480 (N_4480,In_558,In_755);
nor U4481 (N_4481,In_171,In_594);
or U4482 (N_4482,In_1415,In_191);
nor U4483 (N_4483,In_945,In_646);
nor U4484 (N_4484,In_648,In_1320);
or U4485 (N_4485,In_1144,In_1233);
or U4486 (N_4486,In_1422,In_129);
or U4487 (N_4487,In_862,In_1104);
nand U4488 (N_4488,In_879,In_342);
nor U4489 (N_4489,In_106,In_1219);
and U4490 (N_4490,In_37,In_1167);
and U4491 (N_4491,In_879,In_941);
nor U4492 (N_4492,In_693,In_233);
nand U4493 (N_4493,In_272,In_893);
xnor U4494 (N_4494,In_101,In_1215);
nand U4495 (N_4495,In_406,In_1071);
xnor U4496 (N_4496,In_812,In_244);
and U4497 (N_4497,In_31,In_973);
nor U4498 (N_4498,In_1226,In_1041);
nand U4499 (N_4499,In_492,In_943);
nor U4500 (N_4500,In_650,In_109);
xnor U4501 (N_4501,In_19,In_810);
and U4502 (N_4502,In_626,In_1066);
xnor U4503 (N_4503,In_821,In_1145);
nor U4504 (N_4504,In_726,In_90);
xor U4505 (N_4505,In_263,In_385);
nand U4506 (N_4506,In_1426,In_491);
xnor U4507 (N_4507,In_46,In_1464);
or U4508 (N_4508,In_523,In_717);
nand U4509 (N_4509,In_595,In_110);
nand U4510 (N_4510,In_1085,In_793);
nor U4511 (N_4511,In_1074,In_899);
nand U4512 (N_4512,In_924,In_68);
and U4513 (N_4513,In_472,In_870);
and U4514 (N_4514,In_570,In_923);
or U4515 (N_4515,In_223,In_1094);
and U4516 (N_4516,In_112,In_344);
or U4517 (N_4517,In_1300,In_526);
and U4518 (N_4518,In_819,In_116);
xor U4519 (N_4519,In_960,In_1381);
nand U4520 (N_4520,In_99,In_334);
xor U4521 (N_4521,In_789,In_1143);
and U4522 (N_4522,In_152,In_575);
nand U4523 (N_4523,In_131,In_931);
or U4524 (N_4524,In_1121,In_215);
nand U4525 (N_4525,In_548,In_1384);
and U4526 (N_4526,In_219,In_335);
and U4527 (N_4527,In_344,In_905);
nand U4528 (N_4528,In_637,In_624);
or U4529 (N_4529,In_791,In_1455);
or U4530 (N_4530,In_1195,In_289);
xor U4531 (N_4531,In_1312,In_595);
and U4532 (N_4532,In_831,In_819);
nand U4533 (N_4533,In_801,In_1167);
xor U4534 (N_4534,In_1092,In_592);
nor U4535 (N_4535,In_1244,In_589);
xor U4536 (N_4536,In_654,In_1016);
and U4537 (N_4537,In_1022,In_236);
nand U4538 (N_4538,In_197,In_194);
nand U4539 (N_4539,In_1484,In_156);
nor U4540 (N_4540,In_0,In_663);
and U4541 (N_4541,In_844,In_167);
and U4542 (N_4542,In_1132,In_570);
nand U4543 (N_4543,In_1405,In_288);
or U4544 (N_4544,In_918,In_1029);
or U4545 (N_4545,In_25,In_785);
or U4546 (N_4546,In_415,In_808);
nand U4547 (N_4547,In_385,In_606);
and U4548 (N_4548,In_581,In_84);
nor U4549 (N_4549,In_946,In_848);
nor U4550 (N_4550,In_595,In_520);
or U4551 (N_4551,In_778,In_1323);
nor U4552 (N_4552,In_463,In_469);
or U4553 (N_4553,In_1338,In_804);
nand U4554 (N_4554,In_530,In_1039);
xnor U4555 (N_4555,In_960,In_1384);
nand U4556 (N_4556,In_916,In_1423);
xnor U4557 (N_4557,In_1194,In_261);
xor U4558 (N_4558,In_33,In_997);
or U4559 (N_4559,In_1126,In_1077);
nor U4560 (N_4560,In_980,In_1351);
and U4561 (N_4561,In_328,In_1102);
xor U4562 (N_4562,In_438,In_967);
or U4563 (N_4563,In_1391,In_1115);
or U4564 (N_4564,In_1484,In_627);
or U4565 (N_4565,In_633,In_718);
xnor U4566 (N_4566,In_434,In_777);
or U4567 (N_4567,In_607,In_968);
or U4568 (N_4568,In_184,In_990);
or U4569 (N_4569,In_1462,In_726);
and U4570 (N_4570,In_701,In_616);
or U4571 (N_4571,In_1464,In_680);
or U4572 (N_4572,In_388,In_925);
or U4573 (N_4573,In_229,In_335);
or U4574 (N_4574,In_1028,In_841);
or U4575 (N_4575,In_905,In_926);
xor U4576 (N_4576,In_392,In_1276);
nand U4577 (N_4577,In_554,In_669);
nor U4578 (N_4578,In_136,In_578);
nor U4579 (N_4579,In_1090,In_961);
nand U4580 (N_4580,In_708,In_199);
nand U4581 (N_4581,In_345,In_1369);
nand U4582 (N_4582,In_468,In_946);
nor U4583 (N_4583,In_550,In_1341);
nor U4584 (N_4584,In_1007,In_99);
nand U4585 (N_4585,In_198,In_68);
nand U4586 (N_4586,In_215,In_1234);
nand U4587 (N_4587,In_551,In_1484);
and U4588 (N_4588,In_470,In_568);
or U4589 (N_4589,In_137,In_653);
nand U4590 (N_4590,In_1140,In_1244);
nor U4591 (N_4591,In_738,In_241);
or U4592 (N_4592,In_1188,In_252);
xor U4593 (N_4593,In_1381,In_80);
and U4594 (N_4594,In_1302,In_1224);
xor U4595 (N_4595,In_1335,In_0);
xor U4596 (N_4596,In_462,In_1376);
xnor U4597 (N_4597,In_284,In_887);
xnor U4598 (N_4598,In_1339,In_1468);
nor U4599 (N_4599,In_1159,In_780);
xnor U4600 (N_4600,In_997,In_417);
or U4601 (N_4601,In_1117,In_429);
xnor U4602 (N_4602,In_1095,In_487);
and U4603 (N_4603,In_1407,In_1225);
xnor U4604 (N_4604,In_1180,In_524);
and U4605 (N_4605,In_1369,In_1465);
xor U4606 (N_4606,In_1430,In_1095);
nor U4607 (N_4607,In_139,In_1453);
or U4608 (N_4608,In_224,In_308);
nand U4609 (N_4609,In_1208,In_664);
or U4610 (N_4610,In_387,In_982);
nand U4611 (N_4611,In_803,In_1344);
xnor U4612 (N_4612,In_734,In_1321);
nand U4613 (N_4613,In_1215,In_1255);
or U4614 (N_4614,In_738,In_1235);
xor U4615 (N_4615,In_202,In_644);
and U4616 (N_4616,In_849,In_878);
xor U4617 (N_4617,In_915,In_797);
or U4618 (N_4618,In_1325,In_886);
or U4619 (N_4619,In_294,In_487);
xnor U4620 (N_4620,In_675,In_1348);
xnor U4621 (N_4621,In_778,In_1100);
nand U4622 (N_4622,In_1143,In_768);
and U4623 (N_4623,In_489,In_777);
and U4624 (N_4624,In_423,In_1008);
nor U4625 (N_4625,In_1350,In_640);
and U4626 (N_4626,In_722,In_676);
nand U4627 (N_4627,In_444,In_290);
xor U4628 (N_4628,In_890,In_1170);
nand U4629 (N_4629,In_879,In_1379);
nor U4630 (N_4630,In_1071,In_234);
and U4631 (N_4631,In_1209,In_822);
or U4632 (N_4632,In_1379,In_1386);
xnor U4633 (N_4633,In_127,In_455);
and U4634 (N_4634,In_1408,In_866);
nand U4635 (N_4635,In_745,In_843);
and U4636 (N_4636,In_800,In_680);
and U4637 (N_4637,In_1051,In_407);
nand U4638 (N_4638,In_1288,In_965);
and U4639 (N_4639,In_1388,In_1485);
or U4640 (N_4640,In_804,In_1359);
nor U4641 (N_4641,In_199,In_576);
xor U4642 (N_4642,In_294,In_1262);
or U4643 (N_4643,In_566,In_333);
xor U4644 (N_4644,In_868,In_1243);
nand U4645 (N_4645,In_459,In_928);
nand U4646 (N_4646,In_1214,In_668);
or U4647 (N_4647,In_30,In_929);
and U4648 (N_4648,In_211,In_529);
xor U4649 (N_4649,In_179,In_1369);
and U4650 (N_4650,In_701,In_516);
xor U4651 (N_4651,In_558,In_124);
and U4652 (N_4652,In_1188,In_717);
xor U4653 (N_4653,In_1298,In_794);
and U4654 (N_4654,In_1383,In_173);
nor U4655 (N_4655,In_1200,In_908);
xor U4656 (N_4656,In_822,In_1278);
nand U4657 (N_4657,In_475,In_281);
xnor U4658 (N_4658,In_408,In_1477);
or U4659 (N_4659,In_580,In_976);
xor U4660 (N_4660,In_1355,In_1099);
nand U4661 (N_4661,In_323,In_221);
and U4662 (N_4662,In_486,In_893);
nor U4663 (N_4663,In_1298,In_635);
and U4664 (N_4664,In_556,In_660);
nand U4665 (N_4665,In_209,In_585);
or U4666 (N_4666,In_30,In_554);
xnor U4667 (N_4667,In_590,In_1452);
or U4668 (N_4668,In_812,In_750);
nor U4669 (N_4669,In_817,In_1360);
nor U4670 (N_4670,In_383,In_497);
nor U4671 (N_4671,In_72,In_1035);
and U4672 (N_4672,In_1241,In_371);
nand U4673 (N_4673,In_905,In_1230);
and U4674 (N_4674,In_1368,In_686);
nor U4675 (N_4675,In_242,In_591);
nand U4676 (N_4676,In_464,In_446);
nand U4677 (N_4677,In_185,In_229);
or U4678 (N_4678,In_492,In_236);
or U4679 (N_4679,In_954,In_180);
and U4680 (N_4680,In_1279,In_1313);
and U4681 (N_4681,In_66,In_612);
and U4682 (N_4682,In_1328,In_1113);
xnor U4683 (N_4683,In_797,In_663);
nor U4684 (N_4684,In_192,In_756);
and U4685 (N_4685,In_1361,In_709);
nand U4686 (N_4686,In_482,In_795);
nand U4687 (N_4687,In_1111,In_144);
or U4688 (N_4688,In_447,In_800);
xnor U4689 (N_4689,In_1114,In_49);
nand U4690 (N_4690,In_1456,In_342);
and U4691 (N_4691,In_1492,In_836);
nor U4692 (N_4692,In_180,In_824);
nand U4693 (N_4693,In_1205,In_70);
xnor U4694 (N_4694,In_137,In_70);
nor U4695 (N_4695,In_229,In_1269);
nor U4696 (N_4696,In_1325,In_984);
and U4697 (N_4697,In_71,In_982);
nor U4698 (N_4698,In_546,In_628);
and U4699 (N_4699,In_1329,In_1074);
nor U4700 (N_4700,In_807,In_930);
nand U4701 (N_4701,In_396,In_1231);
nand U4702 (N_4702,In_102,In_1156);
xnor U4703 (N_4703,In_1320,In_521);
nand U4704 (N_4704,In_829,In_183);
xor U4705 (N_4705,In_740,In_518);
nand U4706 (N_4706,In_587,In_1313);
nor U4707 (N_4707,In_1389,In_794);
and U4708 (N_4708,In_1220,In_888);
or U4709 (N_4709,In_1226,In_599);
nand U4710 (N_4710,In_1487,In_1470);
nor U4711 (N_4711,In_670,In_1468);
and U4712 (N_4712,In_871,In_642);
nor U4713 (N_4713,In_85,In_641);
or U4714 (N_4714,In_99,In_1163);
and U4715 (N_4715,In_1196,In_829);
and U4716 (N_4716,In_1181,In_155);
nor U4717 (N_4717,In_713,In_19);
nor U4718 (N_4718,In_704,In_512);
or U4719 (N_4719,In_1321,In_928);
and U4720 (N_4720,In_55,In_212);
nor U4721 (N_4721,In_1157,In_969);
xnor U4722 (N_4722,In_984,In_818);
nand U4723 (N_4723,In_37,In_518);
or U4724 (N_4724,In_1214,In_1287);
xor U4725 (N_4725,In_124,In_1084);
or U4726 (N_4726,In_358,In_48);
or U4727 (N_4727,In_1202,In_599);
xor U4728 (N_4728,In_1423,In_7);
or U4729 (N_4729,In_188,In_1271);
xnor U4730 (N_4730,In_4,In_757);
xnor U4731 (N_4731,In_1185,In_1400);
nand U4732 (N_4732,In_483,In_1209);
or U4733 (N_4733,In_638,In_712);
nand U4734 (N_4734,In_86,In_1092);
nand U4735 (N_4735,In_121,In_994);
and U4736 (N_4736,In_852,In_1419);
or U4737 (N_4737,In_748,In_125);
xnor U4738 (N_4738,In_1322,In_1400);
xnor U4739 (N_4739,In_776,In_1059);
nand U4740 (N_4740,In_1257,In_700);
nor U4741 (N_4741,In_1233,In_723);
and U4742 (N_4742,In_1297,In_225);
nor U4743 (N_4743,In_835,In_1285);
xnor U4744 (N_4744,In_737,In_885);
or U4745 (N_4745,In_810,In_159);
nor U4746 (N_4746,In_540,In_909);
xor U4747 (N_4747,In_624,In_1147);
nand U4748 (N_4748,In_516,In_51);
or U4749 (N_4749,In_568,In_1324);
nand U4750 (N_4750,In_194,In_1115);
nand U4751 (N_4751,In_230,In_331);
nand U4752 (N_4752,In_1026,In_91);
xnor U4753 (N_4753,In_319,In_1330);
and U4754 (N_4754,In_1449,In_1271);
nor U4755 (N_4755,In_910,In_885);
and U4756 (N_4756,In_1445,In_578);
or U4757 (N_4757,In_1280,In_477);
nor U4758 (N_4758,In_545,In_1125);
and U4759 (N_4759,In_1170,In_1194);
xnor U4760 (N_4760,In_1264,In_389);
xnor U4761 (N_4761,In_277,In_801);
xnor U4762 (N_4762,In_967,In_280);
nand U4763 (N_4763,In_914,In_1019);
and U4764 (N_4764,In_955,In_1086);
nand U4765 (N_4765,In_1144,In_1068);
and U4766 (N_4766,In_651,In_415);
nand U4767 (N_4767,In_617,In_299);
xnor U4768 (N_4768,In_887,In_166);
or U4769 (N_4769,In_725,In_336);
xor U4770 (N_4770,In_1449,In_1461);
nand U4771 (N_4771,In_1020,In_106);
xnor U4772 (N_4772,In_58,In_925);
and U4773 (N_4773,In_513,In_41);
or U4774 (N_4774,In_412,In_235);
or U4775 (N_4775,In_285,In_26);
xnor U4776 (N_4776,In_775,In_610);
and U4777 (N_4777,In_250,In_827);
xor U4778 (N_4778,In_1198,In_475);
nor U4779 (N_4779,In_1037,In_248);
nor U4780 (N_4780,In_605,In_345);
or U4781 (N_4781,In_1127,In_576);
or U4782 (N_4782,In_1256,In_1057);
nor U4783 (N_4783,In_784,In_841);
xor U4784 (N_4784,In_271,In_618);
nand U4785 (N_4785,In_1161,In_408);
xor U4786 (N_4786,In_237,In_1168);
nand U4787 (N_4787,In_15,In_1085);
nor U4788 (N_4788,In_864,In_503);
nand U4789 (N_4789,In_320,In_587);
or U4790 (N_4790,In_23,In_91);
and U4791 (N_4791,In_924,In_579);
nand U4792 (N_4792,In_1096,In_261);
nor U4793 (N_4793,In_809,In_193);
nand U4794 (N_4794,In_257,In_1207);
nand U4795 (N_4795,In_328,In_1317);
xnor U4796 (N_4796,In_1450,In_1056);
nor U4797 (N_4797,In_1068,In_921);
nor U4798 (N_4798,In_1120,In_1472);
and U4799 (N_4799,In_242,In_79);
xor U4800 (N_4800,In_162,In_223);
nand U4801 (N_4801,In_764,In_381);
nand U4802 (N_4802,In_617,In_336);
xnor U4803 (N_4803,In_915,In_268);
nor U4804 (N_4804,In_1278,In_696);
or U4805 (N_4805,In_549,In_710);
nand U4806 (N_4806,In_880,In_469);
nor U4807 (N_4807,In_197,In_107);
and U4808 (N_4808,In_545,In_825);
or U4809 (N_4809,In_496,In_677);
or U4810 (N_4810,In_745,In_288);
and U4811 (N_4811,In_21,In_1411);
or U4812 (N_4812,In_195,In_1167);
nand U4813 (N_4813,In_1203,In_744);
nand U4814 (N_4814,In_233,In_603);
nand U4815 (N_4815,In_191,In_706);
xor U4816 (N_4816,In_553,In_1477);
xor U4817 (N_4817,In_720,In_939);
or U4818 (N_4818,In_655,In_1390);
xor U4819 (N_4819,In_1122,In_782);
nor U4820 (N_4820,In_616,In_426);
nor U4821 (N_4821,In_353,In_1024);
xnor U4822 (N_4822,In_874,In_62);
nor U4823 (N_4823,In_492,In_520);
nand U4824 (N_4824,In_512,In_271);
nand U4825 (N_4825,In_1328,In_1141);
or U4826 (N_4826,In_1394,In_511);
and U4827 (N_4827,In_571,In_1321);
nor U4828 (N_4828,In_676,In_767);
and U4829 (N_4829,In_119,In_1492);
or U4830 (N_4830,In_727,In_1079);
or U4831 (N_4831,In_563,In_1200);
nand U4832 (N_4832,In_1184,In_520);
nand U4833 (N_4833,In_725,In_942);
xnor U4834 (N_4834,In_1141,In_589);
and U4835 (N_4835,In_490,In_513);
or U4836 (N_4836,In_955,In_461);
nor U4837 (N_4837,In_827,In_477);
nor U4838 (N_4838,In_1167,In_1477);
nand U4839 (N_4839,In_1078,In_468);
nor U4840 (N_4840,In_288,In_1022);
xnor U4841 (N_4841,In_906,In_830);
and U4842 (N_4842,In_384,In_1025);
xnor U4843 (N_4843,In_731,In_97);
nand U4844 (N_4844,In_32,In_422);
xor U4845 (N_4845,In_158,In_885);
and U4846 (N_4846,In_1422,In_1335);
xor U4847 (N_4847,In_947,In_1128);
and U4848 (N_4848,In_1440,In_740);
xnor U4849 (N_4849,In_784,In_1389);
nand U4850 (N_4850,In_1146,In_1491);
xor U4851 (N_4851,In_1154,In_1039);
nor U4852 (N_4852,In_1394,In_61);
nand U4853 (N_4853,In_61,In_164);
nand U4854 (N_4854,In_210,In_883);
xor U4855 (N_4855,In_817,In_1410);
or U4856 (N_4856,In_113,In_956);
nand U4857 (N_4857,In_273,In_1220);
nor U4858 (N_4858,In_1249,In_561);
and U4859 (N_4859,In_1201,In_729);
nand U4860 (N_4860,In_934,In_1110);
and U4861 (N_4861,In_1468,In_1497);
xor U4862 (N_4862,In_1383,In_614);
or U4863 (N_4863,In_665,In_1125);
nand U4864 (N_4864,In_995,In_1422);
nand U4865 (N_4865,In_511,In_727);
or U4866 (N_4866,In_1223,In_7);
or U4867 (N_4867,In_413,In_229);
and U4868 (N_4868,In_471,In_719);
nor U4869 (N_4869,In_762,In_945);
nand U4870 (N_4870,In_545,In_72);
xor U4871 (N_4871,In_1090,In_918);
nand U4872 (N_4872,In_291,In_226);
nand U4873 (N_4873,In_412,In_913);
or U4874 (N_4874,In_171,In_1391);
or U4875 (N_4875,In_110,In_855);
or U4876 (N_4876,In_673,In_537);
nand U4877 (N_4877,In_524,In_495);
or U4878 (N_4878,In_221,In_1075);
nand U4879 (N_4879,In_23,In_430);
and U4880 (N_4880,In_1301,In_716);
nand U4881 (N_4881,In_847,In_472);
xor U4882 (N_4882,In_304,In_1059);
nand U4883 (N_4883,In_577,In_314);
nor U4884 (N_4884,In_1163,In_439);
nor U4885 (N_4885,In_966,In_539);
nand U4886 (N_4886,In_1421,In_60);
and U4887 (N_4887,In_838,In_259);
or U4888 (N_4888,In_645,In_1270);
xor U4889 (N_4889,In_844,In_804);
or U4890 (N_4890,In_108,In_837);
and U4891 (N_4891,In_646,In_321);
or U4892 (N_4892,In_917,In_488);
and U4893 (N_4893,In_804,In_321);
and U4894 (N_4894,In_451,In_1277);
nor U4895 (N_4895,In_1326,In_570);
nand U4896 (N_4896,In_324,In_101);
xnor U4897 (N_4897,In_1470,In_836);
nor U4898 (N_4898,In_1327,In_279);
xor U4899 (N_4899,In_934,In_1150);
nand U4900 (N_4900,In_727,In_1451);
nor U4901 (N_4901,In_818,In_1266);
nand U4902 (N_4902,In_778,In_205);
nand U4903 (N_4903,In_1259,In_1216);
or U4904 (N_4904,In_929,In_148);
nand U4905 (N_4905,In_1190,In_1149);
xor U4906 (N_4906,In_647,In_546);
nand U4907 (N_4907,In_919,In_1194);
and U4908 (N_4908,In_538,In_762);
or U4909 (N_4909,In_1446,In_1266);
xnor U4910 (N_4910,In_1009,In_361);
xor U4911 (N_4911,In_587,In_1443);
nand U4912 (N_4912,In_1361,In_1250);
xor U4913 (N_4913,In_917,In_616);
or U4914 (N_4914,In_942,In_229);
or U4915 (N_4915,In_1303,In_361);
xor U4916 (N_4916,In_366,In_851);
xor U4917 (N_4917,In_767,In_1326);
or U4918 (N_4918,In_1372,In_1295);
or U4919 (N_4919,In_208,In_1075);
nand U4920 (N_4920,In_1038,In_832);
nor U4921 (N_4921,In_430,In_1457);
or U4922 (N_4922,In_56,In_563);
or U4923 (N_4923,In_1398,In_870);
or U4924 (N_4924,In_836,In_1098);
and U4925 (N_4925,In_766,In_956);
nand U4926 (N_4926,In_335,In_972);
xor U4927 (N_4927,In_1389,In_703);
and U4928 (N_4928,In_1018,In_714);
nor U4929 (N_4929,In_1005,In_119);
nor U4930 (N_4930,In_1435,In_233);
or U4931 (N_4931,In_1422,In_22);
and U4932 (N_4932,In_734,In_1153);
or U4933 (N_4933,In_507,In_415);
nor U4934 (N_4934,In_901,In_461);
nor U4935 (N_4935,In_1109,In_347);
nand U4936 (N_4936,In_642,In_1075);
or U4937 (N_4937,In_1274,In_653);
xnor U4938 (N_4938,In_776,In_1298);
and U4939 (N_4939,In_53,In_403);
and U4940 (N_4940,In_135,In_784);
nor U4941 (N_4941,In_314,In_237);
nor U4942 (N_4942,In_518,In_102);
nand U4943 (N_4943,In_974,In_1114);
nor U4944 (N_4944,In_1362,In_1255);
xor U4945 (N_4945,In_1121,In_855);
nand U4946 (N_4946,In_539,In_1220);
or U4947 (N_4947,In_1186,In_248);
or U4948 (N_4948,In_998,In_823);
or U4949 (N_4949,In_47,In_541);
and U4950 (N_4950,In_259,In_798);
nand U4951 (N_4951,In_232,In_1185);
nor U4952 (N_4952,In_929,In_1033);
or U4953 (N_4953,In_206,In_670);
xor U4954 (N_4954,In_531,In_922);
or U4955 (N_4955,In_1035,In_762);
nor U4956 (N_4956,In_846,In_660);
nand U4957 (N_4957,In_1059,In_607);
or U4958 (N_4958,In_1275,In_184);
nor U4959 (N_4959,In_782,In_198);
nand U4960 (N_4960,In_667,In_1182);
and U4961 (N_4961,In_1047,In_620);
and U4962 (N_4962,In_108,In_98);
nand U4963 (N_4963,In_57,In_646);
nand U4964 (N_4964,In_91,In_1336);
xnor U4965 (N_4965,In_1032,In_1486);
or U4966 (N_4966,In_1125,In_952);
or U4967 (N_4967,In_971,In_1165);
and U4968 (N_4968,In_1112,In_11);
or U4969 (N_4969,In_1097,In_1371);
nor U4970 (N_4970,In_331,In_1303);
and U4971 (N_4971,In_468,In_62);
and U4972 (N_4972,In_1024,In_1290);
xor U4973 (N_4973,In_705,In_615);
xnor U4974 (N_4974,In_209,In_63);
nor U4975 (N_4975,In_850,In_44);
xor U4976 (N_4976,In_1180,In_181);
and U4977 (N_4977,In_604,In_1012);
nand U4978 (N_4978,In_316,In_718);
or U4979 (N_4979,In_775,In_61);
nor U4980 (N_4980,In_1136,In_968);
nand U4981 (N_4981,In_1089,In_1428);
nor U4982 (N_4982,In_295,In_509);
nand U4983 (N_4983,In_78,In_74);
nor U4984 (N_4984,In_928,In_924);
xnor U4985 (N_4985,In_1372,In_930);
xnor U4986 (N_4986,In_911,In_1168);
nand U4987 (N_4987,In_1471,In_721);
and U4988 (N_4988,In_14,In_1424);
or U4989 (N_4989,In_1214,In_720);
or U4990 (N_4990,In_1356,In_858);
nor U4991 (N_4991,In_442,In_378);
xor U4992 (N_4992,In_968,In_1413);
or U4993 (N_4993,In_1463,In_641);
nor U4994 (N_4994,In_1028,In_668);
and U4995 (N_4995,In_1100,In_1455);
nor U4996 (N_4996,In_447,In_371);
nand U4997 (N_4997,In_385,In_768);
and U4998 (N_4998,In_81,In_260);
and U4999 (N_4999,In_1338,In_196);
nand U5000 (N_5000,N_2509,N_931);
nand U5001 (N_5001,N_4271,N_3656);
xor U5002 (N_5002,N_540,N_1521);
nor U5003 (N_5003,N_130,N_3456);
xnor U5004 (N_5004,N_2405,N_3706);
xnor U5005 (N_5005,N_4987,N_1162);
xnor U5006 (N_5006,N_1371,N_2733);
nand U5007 (N_5007,N_24,N_4554);
and U5008 (N_5008,N_3079,N_1463);
and U5009 (N_5009,N_4153,N_1026);
and U5010 (N_5010,N_4031,N_418);
nor U5011 (N_5011,N_1193,N_2673);
nor U5012 (N_5012,N_3904,N_4482);
xor U5013 (N_5013,N_2348,N_3486);
nor U5014 (N_5014,N_3325,N_4771);
xor U5015 (N_5015,N_2598,N_4546);
and U5016 (N_5016,N_1070,N_1042);
xnor U5017 (N_5017,N_3741,N_3749);
or U5018 (N_5018,N_684,N_1221);
and U5019 (N_5019,N_909,N_1702);
nor U5020 (N_5020,N_338,N_4532);
or U5021 (N_5021,N_2525,N_4872);
or U5022 (N_5022,N_18,N_1054);
and U5023 (N_5023,N_3849,N_4486);
nor U5024 (N_5024,N_4113,N_3568);
nand U5025 (N_5025,N_3435,N_4230);
xor U5026 (N_5026,N_373,N_2634);
and U5027 (N_5027,N_4093,N_1027);
and U5028 (N_5028,N_1700,N_502);
and U5029 (N_5029,N_3681,N_2165);
and U5030 (N_5030,N_1100,N_3990);
or U5031 (N_5031,N_431,N_1148);
nand U5032 (N_5032,N_4525,N_4212);
nand U5033 (N_5033,N_720,N_3474);
xor U5034 (N_5034,N_4604,N_2421);
nand U5035 (N_5035,N_1134,N_366);
or U5036 (N_5036,N_3023,N_3705);
or U5037 (N_5037,N_3738,N_1562);
and U5038 (N_5038,N_2178,N_22);
nor U5039 (N_5039,N_2305,N_942);
or U5040 (N_5040,N_3016,N_499);
and U5041 (N_5041,N_648,N_4178);
nand U5042 (N_5042,N_1681,N_2296);
nor U5043 (N_5043,N_3508,N_2869);
and U5044 (N_5044,N_1331,N_126);
or U5045 (N_5045,N_4477,N_4308);
xor U5046 (N_5046,N_2859,N_2020);
xor U5047 (N_5047,N_1428,N_3610);
nor U5048 (N_5048,N_3215,N_2422);
or U5049 (N_5049,N_2795,N_1970);
nor U5050 (N_5050,N_2280,N_2460);
and U5051 (N_5051,N_3346,N_328);
and U5052 (N_5052,N_4009,N_4294);
and U5053 (N_5053,N_63,N_4639);
nand U5054 (N_5054,N_3751,N_2491);
nor U5055 (N_5055,N_4876,N_281);
nand U5056 (N_5056,N_1957,N_2454);
and U5057 (N_5057,N_1672,N_2394);
nor U5058 (N_5058,N_2785,N_602);
and U5059 (N_5059,N_3658,N_3034);
xnor U5060 (N_5060,N_1487,N_4171);
and U5061 (N_5061,N_2988,N_1457);
nand U5062 (N_5062,N_3226,N_204);
or U5063 (N_5063,N_3632,N_2094);
or U5064 (N_5064,N_4255,N_1788);
nor U5065 (N_5065,N_2116,N_4471);
nand U5066 (N_5066,N_4084,N_457);
and U5067 (N_5067,N_3512,N_2319);
and U5068 (N_5068,N_3283,N_2963);
nand U5069 (N_5069,N_3947,N_640);
and U5070 (N_5070,N_1746,N_2860);
or U5071 (N_5071,N_1663,N_159);
xnor U5072 (N_5072,N_4493,N_456);
or U5073 (N_5073,N_2936,N_2419);
or U5074 (N_5074,N_1769,N_3671);
or U5075 (N_5075,N_4997,N_521);
xnor U5076 (N_5076,N_320,N_899);
or U5077 (N_5077,N_1912,N_3551);
and U5078 (N_5078,N_1418,N_3110);
nand U5079 (N_5079,N_3184,N_3822);
xnor U5080 (N_5080,N_1851,N_1359);
and U5081 (N_5081,N_2397,N_1108);
and U5082 (N_5082,N_4431,N_4733);
xor U5083 (N_5083,N_4908,N_3376);
xor U5084 (N_5084,N_3466,N_4354);
xor U5085 (N_5085,N_3121,N_1741);
nand U5086 (N_5086,N_210,N_2373);
and U5087 (N_5087,N_1955,N_1842);
nand U5088 (N_5088,N_4231,N_1282);
and U5089 (N_5089,N_738,N_1308);
nand U5090 (N_5090,N_544,N_2360);
xor U5091 (N_5091,N_4242,N_2058);
and U5092 (N_5092,N_2036,N_3020);
nand U5093 (N_5093,N_3928,N_3434);
xnor U5094 (N_5094,N_3878,N_2645);
or U5095 (N_5095,N_4557,N_3061);
or U5096 (N_5096,N_3120,N_1831);
nor U5097 (N_5097,N_3044,N_3267);
nor U5098 (N_5098,N_4207,N_2226);
nor U5099 (N_5099,N_2221,N_4626);
nand U5100 (N_5100,N_2725,N_4960);
and U5101 (N_5101,N_2299,N_400);
or U5102 (N_5102,N_1061,N_688);
xor U5103 (N_5103,N_2736,N_2528);
xor U5104 (N_5104,N_3560,N_788);
or U5105 (N_5105,N_3567,N_4819);
nor U5106 (N_5106,N_4569,N_1944);
or U5107 (N_5107,N_3861,N_1640);
nor U5108 (N_5108,N_3549,N_2462);
or U5109 (N_5109,N_2483,N_1563);
or U5110 (N_5110,N_1569,N_1805);
or U5111 (N_5111,N_1478,N_2463);
nand U5112 (N_5112,N_3497,N_1347);
nand U5113 (N_5113,N_923,N_1911);
nor U5114 (N_5114,N_4511,N_472);
nor U5115 (N_5115,N_3850,N_62);
nand U5116 (N_5116,N_1990,N_113);
or U5117 (N_5117,N_4364,N_4622);
nand U5118 (N_5118,N_1548,N_2225);
and U5119 (N_5119,N_3894,N_2987);
or U5120 (N_5120,N_1315,N_1650);
and U5121 (N_5121,N_3098,N_1690);
nor U5122 (N_5122,N_858,N_2119);
nand U5123 (N_5123,N_4918,N_298);
xor U5124 (N_5124,N_2335,N_3882);
xor U5125 (N_5125,N_4362,N_187);
xnor U5126 (N_5126,N_3031,N_1033);
nand U5127 (N_5127,N_1713,N_928);
nand U5128 (N_5128,N_4609,N_1124);
or U5129 (N_5129,N_3926,N_2030);
xnor U5130 (N_5130,N_2264,N_331);
and U5131 (N_5131,N_741,N_636);
and U5132 (N_5132,N_3889,N_987);
xnor U5133 (N_5133,N_1089,N_1709);
xor U5134 (N_5134,N_940,N_624);
nand U5135 (N_5135,N_2189,N_4046);
nand U5136 (N_5136,N_360,N_322);
xnor U5137 (N_5137,N_3745,N_4290);
or U5138 (N_5138,N_1183,N_1489);
xor U5139 (N_5139,N_2130,N_4528);
nand U5140 (N_5140,N_2612,N_1517);
nor U5141 (N_5141,N_3866,N_1723);
and U5142 (N_5142,N_4959,N_4065);
nand U5143 (N_5143,N_888,N_3320);
nand U5144 (N_5144,N_2793,N_2105);
or U5145 (N_5145,N_4864,N_4766);
nor U5146 (N_5146,N_4110,N_3423);
or U5147 (N_5147,N_3627,N_2787);
or U5148 (N_5148,N_223,N_2018);
or U5149 (N_5149,N_3930,N_4284);
nand U5150 (N_5150,N_4800,N_3351);
xnor U5151 (N_5151,N_1960,N_3363);
nor U5152 (N_5152,N_3246,N_2025);
and U5153 (N_5153,N_96,N_3495);
or U5154 (N_5154,N_69,N_737);
or U5155 (N_5155,N_1157,N_3287);
nor U5156 (N_5156,N_1461,N_4785);
nor U5157 (N_5157,N_496,N_2633);
nor U5158 (N_5158,N_736,N_4000);
nor U5159 (N_5159,N_983,N_3471);
nand U5160 (N_5160,N_4323,N_1223);
or U5161 (N_5161,N_2039,N_4698);
nor U5162 (N_5162,N_3250,N_616);
or U5163 (N_5163,N_1513,N_3694);
nand U5164 (N_5164,N_3914,N_1365);
or U5165 (N_5165,N_2705,N_2540);
nand U5166 (N_5166,N_3304,N_3714);
or U5167 (N_5167,N_763,N_3203);
xor U5168 (N_5168,N_3692,N_2206);
nor U5169 (N_5169,N_4878,N_1734);
and U5170 (N_5170,N_1730,N_406);
or U5171 (N_5171,N_1085,N_1274);
and U5172 (N_5172,N_2726,N_866);
nand U5173 (N_5173,N_3931,N_2470);
nor U5174 (N_5174,N_1310,N_2970);
and U5175 (N_5175,N_4372,N_1067);
and U5176 (N_5176,N_1506,N_3643);
or U5177 (N_5177,N_4795,N_2340);
or U5178 (N_5178,N_108,N_219);
and U5179 (N_5179,N_4317,N_4285);
nand U5180 (N_5180,N_3564,N_4253);
and U5181 (N_5181,N_2666,N_1235);
and U5182 (N_5182,N_415,N_395);
nor U5183 (N_5183,N_1825,N_82);
and U5184 (N_5184,N_4907,N_149);
and U5185 (N_5185,N_4923,N_1128);
nand U5186 (N_5186,N_343,N_1847);
or U5187 (N_5187,N_559,N_1916);
nand U5188 (N_5188,N_2883,N_1450);
or U5189 (N_5189,N_2583,N_686);
nand U5190 (N_5190,N_4660,N_32);
or U5191 (N_5191,N_4168,N_1080);
nor U5192 (N_5192,N_355,N_2717);
nor U5193 (N_5193,N_629,N_1322);
xor U5194 (N_5194,N_1777,N_3265);
nor U5195 (N_5195,N_1592,N_1856);
nor U5196 (N_5196,N_4512,N_3485);
xnor U5197 (N_5197,N_614,N_1287);
xnor U5198 (N_5198,N_4999,N_4919);
or U5199 (N_5199,N_454,N_3397);
or U5200 (N_5200,N_1895,N_482);
nor U5201 (N_5201,N_2064,N_1989);
nor U5202 (N_5202,N_1049,N_3489);
nor U5203 (N_5203,N_1948,N_574);
and U5204 (N_5204,N_1606,N_3594);
and U5205 (N_5205,N_3177,N_347);
or U5206 (N_5206,N_2383,N_4088);
and U5207 (N_5207,N_3446,N_2060);
nor U5208 (N_5208,N_1707,N_2448);
nor U5209 (N_5209,N_3377,N_2721);
and U5210 (N_5210,N_3647,N_1171);
xor U5211 (N_5211,N_4547,N_2144);
and U5212 (N_5212,N_4881,N_630);
nor U5213 (N_5213,N_893,N_3836);
xor U5214 (N_5214,N_4183,N_1139);
or U5215 (N_5215,N_631,N_2196);
xnor U5216 (N_5216,N_2620,N_2849);
and U5217 (N_5217,N_2567,N_285);
or U5218 (N_5218,N_878,N_4325);
nand U5219 (N_5219,N_1285,N_970);
and U5220 (N_5220,N_1182,N_2112);
nand U5221 (N_5221,N_2866,N_4472);
nand U5222 (N_5222,N_770,N_3359);
or U5223 (N_5223,N_2701,N_4984);
and U5224 (N_5224,N_4076,N_958);
or U5225 (N_5225,N_3787,N_4976);
nor U5226 (N_5226,N_817,N_4107);
or U5227 (N_5227,N_1991,N_4479);
nor U5228 (N_5228,N_3401,N_3187);
nand U5229 (N_5229,N_4192,N_4464);
nand U5230 (N_5230,N_1036,N_4939);
or U5231 (N_5231,N_3905,N_4992);
xnor U5232 (N_5232,N_3422,N_2820);
and U5233 (N_5233,N_4659,N_259);
nor U5234 (N_5234,N_1999,N_2902);
nand U5235 (N_5235,N_3729,N_3007);
and U5236 (N_5236,N_417,N_696);
or U5237 (N_5237,N_284,N_4086);
nand U5238 (N_5238,N_74,N_447);
nor U5239 (N_5239,N_3747,N_261);
nor U5240 (N_5240,N_1732,N_2152);
nand U5241 (N_5241,N_3563,N_701);
xor U5242 (N_5242,N_2602,N_4135);
and U5243 (N_5243,N_765,N_2950);
xor U5244 (N_5244,N_1488,N_3504);
xor U5245 (N_5245,N_638,N_613);
and U5246 (N_5246,N_4637,N_4896);
and U5247 (N_5247,N_2535,N_2);
xor U5248 (N_5248,N_811,N_4565);
and U5249 (N_5249,N_4322,N_3342);
or U5250 (N_5250,N_1336,N_428);
xnor U5251 (N_5251,N_2723,N_4498);
nor U5252 (N_5252,N_843,N_4829);
and U5253 (N_5253,N_19,N_795);
and U5254 (N_5254,N_4357,N_304);
xnor U5255 (N_5255,N_804,N_4397);
xnor U5256 (N_5256,N_3319,N_898);
nand U5257 (N_5257,N_1023,N_1740);
nand U5258 (N_5258,N_517,N_356);
nand U5259 (N_5259,N_4151,N_97);
and U5260 (N_5260,N_3072,N_666);
nand U5261 (N_5261,N_730,N_1971);
or U5262 (N_5262,N_1430,N_1753);
nand U5263 (N_5263,N_3676,N_2745);
xor U5264 (N_5264,N_4851,N_4188);
nor U5265 (N_5265,N_3232,N_4758);
nand U5266 (N_5266,N_323,N_4309);
nand U5267 (N_5267,N_3938,N_2870);
nand U5268 (N_5268,N_3666,N_3049);
or U5269 (N_5269,N_4899,N_2054);
nor U5270 (N_5270,N_2026,N_2381);
or U5271 (N_5271,N_3212,N_2449);
and U5272 (N_5272,N_4,N_867);
nand U5273 (N_5273,N_2435,N_4710);
nor U5274 (N_5274,N_1077,N_4406);
xor U5275 (N_5275,N_1214,N_3989);
or U5276 (N_5276,N_4782,N_2316);
nor U5277 (N_5277,N_586,N_2364);
xnor U5278 (N_5278,N_4662,N_4399);
and U5279 (N_5279,N_2984,N_2814);
xor U5280 (N_5280,N_218,N_1622);
or U5281 (N_5281,N_2131,N_4166);
xnor U5282 (N_5282,N_4366,N_3825);
nand U5283 (N_5283,N_1051,N_50);
or U5284 (N_5284,N_3924,N_3565);
nand U5285 (N_5285,N_4582,N_3244);
nor U5286 (N_5286,N_4156,N_1063);
and U5287 (N_5287,N_2012,N_1008);
and U5288 (N_5288,N_3988,N_3799);
nor U5289 (N_5289,N_292,N_2545);
nand U5290 (N_5290,N_1243,N_3827);
or U5291 (N_5291,N_3355,N_1815);
xor U5292 (N_5292,N_4543,N_633);
or U5293 (N_5293,N_4892,N_4011);
nor U5294 (N_5294,N_4529,N_1385);
nand U5295 (N_5295,N_2948,N_514);
or U5296 (N_5296,N_3831,N_3982);
or U5297 (N_5297,N_2711,N_2103);
and U5298 (N_5298,N_810,N_3657);
and U5299 (N_5299,N_354,N_3022);
nor U5300 (N_5300,N_709,N_4213);
or U5301 (N_5301,N_4602,N_985);
nand U5302 (N_5302,N_1111,N_998);
and U5303 (N_5303,N_3733,N_365);
and U5304 (N_5304,N_1328,N_4684);
nand U5305 (N_5305,N_1192,N_4664);
nor U5306 (N_5306,N_3161,N_538);
or U5307 (N_5307,N_2589,N_4560);
and U5308 (N_5308,N_244,N_4839);
xnor U5309 (N_5309,N_3211,N_3717);
xnor U5310 (N_5310,N_708,N_567);
nor U5311 (N_5311,N_4342,N_2256);
nand U5312 (N_5312,N_4601,N_1693);
nand U5313 (N_5313,N_4937,N_1863);
and U5314 (N_5314,N_4013,N_1742);
nand U5315 (N_5315,N_254,N_556);
nand U5316 (N_5316,N_3027,N_1407);
nor U5317 (N_5317,N_3256,N_3992);
and U5318 (N_5318,N_3893,N_656);
xor U5319 (N_5319,N_4097,N_4169);
or U5320 (N_5320,N_2160,N_2926);
and U5321 (N_5321,N_4927,N_4778);
xor U5322 (N_5322,N_3472,N_4217);
nand U5323 (N_5323,N_110,N_4579);
xnor U5324 (N_5324,N_917,N_2811);
nand U5325 (N_5325,N_1780,N_1495);
or U5326 (N_5326,N_3750,N_1229);
or U5327 (N_5327,N_834,N_125);
xnor U5328 (N_5328,N_1520,N_2300);
nand U5329 (N_5329,N_4624,N_2111);
and U5330 (N_5330,N_1617,N_1539);
xnor U5331 (N_5331,N_4860,N_3686);
and U5332 (N_5332,N_1006,N_3393);
and U5333 (N_5333,N_2230,N_520);
nor U5334 (N_5334,N_2268,N_492);
nand U5335 (N_5335,N_584,N_3711);
xor U5336 (N_5336,N_4327,N_4863);
nand U5337 (N_5337,N_753,N_4541);
and U5338 (N_5338,N_3726,N_644);
and U5339 (N_5339,N_2217,N_1394);
xnor U5340 (N_5340,N_1284,N_785);
nand U5341 (N_5341,N_2120,N_570);
nor U5342 (N_5342,N_3442,N_516);
xor U5343 (N_5343,N_3307,N_3769);
xor U5344 (N_5344,N_3114,N_3170);
nor U5345 (N_5345,N_3865,N_1390);
nand U5346 (N_5346,N_4005,N_195);
or U5347 (N_5347,N_2901,N_2081);
nor U5348 (N_5348,N_267,N_4905);
nor U5349 (N_5349,N_3619,N_4934);
and U5350 (N_5350,N_776,N_1422);
xnor U5351 (N_5351,N_3655,N_727);
xor U5352 (N_5352,N_1572,N_2287);
xor U5353 (N_5353,N_2716,N_3502);
nor U5354 (N_5354,N_4690,N_3190);
nor U5355 (N_5355,N_3185,N_3891);
and U5356 (N_5356,N_4643,N_839);
and U5357 (N_5357,N_301,N_2377);
xnor U5358 (N_5358,N_4935,N_2402);
xnor U5359 (N_5359,N_2762,N_1174);
xor U5360 (N_5360,N_2563,N_249);
nor U5361 (N_5361,N_3997,N_2657);
xor U5362 (N_5362,N_3102,N_3392);
nor U5363 (N_5363,N_1695,N_4817);
or U5364 (N_5364,N_4897,N_3217);
xor U5365 (N_5365,N_3235,N_6);
and U5366 (N_5366,N_335,N_1245);
and U5367 (N_5367,N_1503,N_4515);
or U5368 (N_5368,N_3862,N_161);
and U5369 (N_5369,N_3182,N_3562);
nor U5370 (N_5370,N_1518,N_4359);
and U5371 (N_5371,N_3654,N_919);
xor U5372 (N_5372,N_4400,N_697);
or U5373 (N_5373,N_3449,N_132);
nor U5374 (N_5374,N_2106,N_4124);
and U5375 (N_5375,N_1885,N_1072);
xor U5376 (N_5376,N_1620,N_1968);
nand U5377 (N_5377,N_2067,N_3765);
xnor U5378 (N_5378,N_3592,N_1158);
or U5379 (N_5379,N_2115,N_2908);
nand U5380 (N_5380,N_394,N_2191);
nand U5381 (N_5381,N_3948,N_4268);
or U5382 (N_5382,N_699,N_1280);
nor U5383 (N_5383,N_2617,N_1232);
or U5384 (N_5384,N_1393,N_501);
xnor U5385 (N_5385,N_3275,N_4351);
or U5386 (N_5386,N_2514,N_3888);
nor U5387 (N_5387,N_2822,N_276);
and U5388 (N_5388,N_3224,N_140);
or U5389 (N_5389,N_216,N_2239);
and U5390 (N_5390,N_4734,N_2019);
nand U5391 (N_5391,N_2411,N_3732);
nand U5392 (N_5392,N_3361,N_90);
nor U5393 (N_5393,N_2806,N_857);
xor U5394 (N_5394,N_330,N_4832);
nand U5395 (N_5395,N_1890,N_3242);
and U5396 (N_5396,N_4034,N_4506);
or U5397 (N_5397,N_4405,N_627);
nand U5398 (N_5398,N_1002,N_3354);
and U5399 (N_5399,N_1845,N_3500);
nand U5400 (N_5400,N_321,N_1380);
nor U5401 (N_5401,N_767,N_313);
xnor U5402 (N_5402,N_1903,N_2027);
xor U5403 (N_5403,N_2237,N_4078);
nand U5404 (N_5404,N_1798,N_2747);
nand U5405 (N_5405,N_2539,N_3236);
nor U5406 (N_5406,N_3649,N_2065);
nand U5407 (N_5407,N_639,N_924);
xor U5408 (N_5408,N_4804,N_883);
and U5409 (N_5409,N_180,N_768);
xor U5410 (N_5410,N_4380,N_557);
xnor U5411 (N_5411,N_3720,N_2033);
nor U5412 (N_5412,N_446,N_2578);
xor U5413 (N_5413,N_3478,N_2838);
nor U5414 (N_5414,N_4451,N_246);
or U5415 (N_5415,N_2861,N_4779);
nor U5416 (N_5416,N_611,N_2210);
xor U5417 (N_5417,N_4681,N_2248);
nor U5418 (N_5418,N_3383,N_1932);
xor U5419 (N_5419,N_1482,N_55);
xnor U5420 (N_5420,N_1743,N_3756);
or U5421 (N_5421,N_2609,N_3651);
nor U5422 (N_5422,N_3807,N_2604);
nand U5423 (N_5423,N_4002,N_2444);
and U5424 (N_5424,N_4336,N_179);
or U5425 (N_5425,N_2660,N_2088);
or U5426 (N_5426,N_2149,N_4634);
and U5427 (N_5427,N_4016,N_2552);
and U5428 (N_5428,N_2288,N_332);
nor U5429 (N_5429,N_2326,N_2181);
nor U5430 (N_5430,N_4033,N_4735);
xnor U5431 (N_5431,N_4886,N_3927);
or U5432 (N_5432,N_3356,N_3712);
xnor U5433 (N_5433,N_2185,N_758);
nand U5434 (N_5434,N_937,N_3757);
nor U5435 (N_5435,N_4221,N_3477);
xor U5436 (N_5436,N_3641,N_4211);
nor U5437 (N_5437,N_2694,N_2342);
and U5438 (N_5438,N_3123,N_726);
nor U5439 (N_5439,N_3585,N_4942);
or U5440 (N_5440,N_2114,N_2391);
and U5441 (N_5441,N_3279,N_2864);
xor U5442 (N_5442,N_3680,N_2681);
and U5443 (N_5443,N_1455,N_2775);
xor U5444 (N_5444,N_4835,N_816);
or U5445 (N_5445,N_390,N_2555);
or U5446 (N_5446,N_1161,N_553);
and U5447 (N_5447,N_1588,N_4458);
nand U5448 (N_5448,N_4555,N_3852);
and U5449 (N_5449,N_4115,N_173);
and U5450 (N_5450,N_1103,N_4657);
xnor U5451 (N_5451,N_4588,N_4446);
nor U5452 (N_5452,N_3042,N_1047);
xnor U5453 (N_5453,N_1848,N_3199);
nor U5454 (N_5454,N_635,N_1490);
nand U5455 (N_5455,N_473,N_2972);
nor U5456 (N_5456,N_2265,N_980);
or U5457 (N_5457,N_1819,N_2179);
nor U5458 (N_5458,N_4225,N_3445);
nor U5459 (N_5459,N_1424,N_3962);
or U5460 (N_5460,N_4006,N_1281);
nand U5461 (N_5461,N_3727,N_3009);
xor U5462 (N_5462,N_712,N_2479);
and U5463 (N_5463,N_3830,N_2016);
and U5464 (N_5464,N_3548,N_4286);
xor U5465 (N_5465,N_4567,N_3605);
nor U5466 (N_5466,N_3367,N_3682);
and U5467 (N_5467,N_3977,N_563);
and U5468 (N_5468,N_2765,N_3333);
nand U5469 (N_5469,N_2993,N_4334);
xnor U5470 (N_5470,N_3026,N_197);
nand U5471 (N_5471,N_4875,N_475);
xnor U5472 (N_5472,N_383,N_4702);
nor U5473 (N_5473,N_4858,N_2174);
nand U5474 (N_5474,N_3458,N_4012);
xnor U5475 (N_5475,N_4092,N_801);
or U5476 (N_5476,N_1748,N_163);
and U5477 (N_5477,N_36,N_3532);
xor U5478 (N_5478,N_1528,N_4813);
nor U5479 (N_5479,N_3105,N_1486);
and U5480 (N_5480,N_2341,N_830);
and U5481 (N_5481,N_4254,N_3119);
nand U5482 (N_5482,N_2164,N_1614);
nand U5483 (N_5483,N_2443,N_2109);
nand U5484 (N_5484,N_1557,N_2709);
nor U5485 (N_5485,N_3191,N_936);
and U5486 (N_5486,N_812,N_4149);
or U5487 (N_5487,N_4335,N_4859);
xnor U5488 (N_5488,N_3536,N_1833);
nor U5489 (N_5489,N_2318,N_2580);
nand U5490 (N_5490,N_1053,N_932);
nor U5491 (N_5491,N_2575,N_2622);
or U5492 (N_5492,N_2241,N_4954);
xnor U5493 (N_5493,N_524,N_2925);
or U5494 (N_5494,N_1983,N_3909);
nor U5495 (N_5495,N_2302,N_4131);
or U5496 (N_5496,N_2032,N_68);
or U5497 (N_5497,N_2706,N_1934);
and U5498 (N_5498,N_2974,N_4514);
or U5499 (N_5499,N_3863,N_3127);
xnor U5500 (N_5500,N_3625,N_1318);
nand U5501 (N_5501,N_220,N_3484);
nand U5502 (N_5502,N_1443,N_3364);
nor U5503 (N_5503,N_4676,N_2631);
nand U5504 (N_5504,N_4014,N_2504);
xor U5505 (N_5505,N_3076,N_4754);
xor U5506 (N_5506,N_4552,N_1603);
xor U5507 (N_5507,N_2325,N_1629);
nand U5508 (N_5508,N_2590,N_1758);
nand U5509 (N_5509,N_2978,N_3368);
nor U5510 (N_5510,N_3517,N_3172);
nor U5511 (N_5511,N_3764,N_1410);
or U5512 (N_5512,N_3837,N_670);
xor U5513 (N_5513,N_4879,N_1254);
or U5514 (N_5514,N_646,N_4067);
nand U5515 (N_5515,N_4390,N_3648);
nand U5516 (N_5516,N_4931,N_1074);
or U5517 (N_5517,N_3803,N_1196);
and U5518 (N_5518,N_2147,N_1019);
nand U5519 (N_5519,N_2654,N_3229);
nand U5520 (N_5520,N_511,N_881);
or U5521 (N_5521,N_3308,N_549);
xnor U5522 (N_5522,N_3949,N_3986);
or U5523 (N_5523,N_1278,N_1209);
nand U5524 (N_5524,N_4398,N_3010);
nor U5525 (N_5525,N_2766,N_2267);
and U5526 (N_5526,N_3160,N_680);
and U5527 (N_5527,N_2068,N_3703);
and U5528 (N_5528,N_2388,N_781);
nor U5529 (N_5529,N_162,N_325);
or U5530 (N_5530,N_3886,N_2526);
nand U5531 (N_5531,N_3394,N_240);
nor U5532 (N_5532,N_2442,N_1190);
or U5533 (N_5533,N_178,N_4689);
nor U5534 (N_5534,N_2289,N_1947);
and U5535 (N_5535,N_3510,N_2072);
nand U5536 (N_5536,N_1222,N_1706);
or U5537 (N_5537,N_1391,N_1649);
xnor U5538 (N_5538,N_884,N_3778);
xor U5539 (N_5539,N_1295,N_3598);
xnor U5540 (N_5540,N_815,N_4094);
nand U5541 (N_5541,N_3038,N_2450);
nor U5542 (N_5542,N_1453,N_643);
xnor U5543 (N_5543,N_1154,N_4620);
nor U5544 (N_5544,N_1810,N_3073);
xor U5545 (N_5545,N_2371,N_4027);
and U5546 (N_5546,N_2899,N_2625);
and U5547 (N_5547,N_1066,N_116);
nor U5548 (N_5548,N_3074,N_35);
xor U5549 (N_5549,N_3652,N_345);
nand U5550 (N_5550,N_92,N_4220);
xnor U5551 (N_5551,N_297,N_2805);
or U5552 (N_5552,N_326,N_1406);
xor U5553 (N_5553,N_4724,N_1471);
nor U5554 (N_5554,N_2843,N_3834);
nor U5555 (N_5555,N_1686,N_463);
nor U5556 (N_5556,N_1782,N_4669);
xnor U5557 (N_5557,N_2549,N_3314);
xnor U5558 (N_5558,N_1388,N_4307);
and U5559 (N_5559,N_840,N_808);
nand U5560 (N_5560,N_4667,N_2414);
and U5561 (N_5561,N_488,N_4053);
nand U5562 (N_5562,N_2461,N_1972);
xnor U5563 (N_5563,N_539,N_4263);
xor U5564 (N_5564,N_3833,N_407);
or U5565 (N_5565,N_3595,N_1936);
nor U5566 (N_5566,N_2190,N_4200);
or U5567 (N_5567,N_1112,N_3227);
and U5568 (N_5568,N_2516,N_405);
nand U5569 (N_5569,N_4150,N_182);
nand U5570 (N_5570,N_1420,N_1717);
nor U5571 (N_5571,N_1073,N_1203);
or U5572 (N_5572,N_2254,N_3855);
or U5573 (N_5573,N_2997,N_3137);
xnor U5574 (N_5574,N_3142,N_1037);
nand U5575 (N_5575,N_692,N_2324);
nor U5576 (N_5576,N_713,N_4982);
xnor U5577 (N_5577,N_2593,N_2066);
nor U5578 (N_5578,N_3180,N_637);
nor U5579 (N_5579,N_3328,N_3708);
or U5580 (N_5580,N_2886,N_4952);
nor U5581 (N_5581,N_3677,N_1338);
nor U5582 (N_5582,N_4060,N_2133);
xor U5583 (N_5583,N_4729,N_537);
nand U5584 (N_5584,N_2393,N_308);
nand U5585 (N_5585,N_4069,N_3231);
xor U5586 (N_5586,N_3468,N_587);
and U5587 (N_5587,N_814,N_4701);
nand U5588 (N_5588,N_892,N_2837);
and U5589 (N_5589,N_3976,N_4535);
nand U5590 (N_5590,N_1197,N_2720);
or U5591 (N_5591,N_2712,N_963);
nand U5592 (N_5592,N_2955,N_363);
and U5593 (N_5593,N_4452,N_3511);
or U5594 (N_5594,N_1007,N_2197);
nor U5595 (N_5595,N_2070,N_1212);
nand U5596 (N_5596,N_1220,N_641);
and U5597 (N_5597,N_3507,N_2703);
xor U5598 (N_5598,N_2854,N_1060);
nand U5599 (N_5599,N_734,N_1754);
nor U5600 (N_5600,N_4226,N_3631);
nand U5601 (N_5601,N_1299,N_2476);
and U5602 (N_5602,N_4834,N_4861);
and U5603 (N_5603,N_2798,N_1660);
nor U5604 (N_5604,N_3746,N_4404);
xnor U5605 (N_5605,N_4513,N_3981);
xnor U5606 (N_5606,N_2472,N_136);
and U5607 (N_5607,N_3252,N_3668);
or U5608 (N_5608,N_2829,N_4563);
nand U5609 (N_5609,N_1577,N_300);
and U5610 (N_5610,N_4439,N_4642);
xor U5611 (N_5611,N_2494,N_3097);
nor U5612 (N_5612,N_2322,N_4129);
nor U5613 (N_5613,N_3513,N_4048);
xnor U5614 (N_5614,N_3601,N_1744);
nor U5615 (N_5615,N_494,N_619);
nor U5616 (N_5616,N_280,N_590);
and U5617 (N_5617,N_237,N_2004);
nor U5618 (N_5618,N_2788,N_4744);
or U5619 (N_5619,N_2098,N_2235);
nor U5620 (N_5620,N_2420,N_3552);
nor U5621 (N_5621,N_3636,N_3306);
or U5622 (N_5622,N_2942,N_3183);
or U5623 (N_5623,N_4244,N_4668);
xnor U5624 (N_5624,N_3853,N_1963);
xnor U5625 (N_5625,N_2281,N_4035);
nand U5626 (N_5626,N_1868,N_3338);
nor U5627 (N_5627,N_992,N_547);
and U5628 (N_5628,N_1638,N_4182);
or U5629 (N_5629,N_4059,N_4723);
xor U5630 (N_5630,N_3885,N_3154);
xor U5631 (N_5631,N_2734,N_2292);
nand U5632 (N_5632,N_2357,N_973);
nor U5633 (N_5633,N_1522,N_2917);
nand U5634 (N_5634,N_4103,N_1998);
and U5635 (N_5635,N_2495,N_2808);
and U5636 (N_5636,N_1163,N_2406);
or U5637 (N_5637,N_3277,N_1529);
or U5638 (N_5638,N_486,N_3533);
nand U5639 (N_5639,N_3626,N_1218);
and U5640 (N_5640,N_3752,N_1883);
and U5641 (N_5641,N_1186,N_3494);
or U5642 (N_5642,N_3104,N_1710);
xor U5643 (N_5643,N_2658,N_1779);
and U5644 (N_5644,N_1584,N_4559);
nor U5645 (N_5645,N_4416,N_2676);
and U5646 (N_5646,N_1068,N_2317);
nor U5647 (N_5647,N_3133,N_2770);
or U5648 (N_5648,N_1821,N_4889);
or U5649 (N_5649,N_4450,N_3200);
nand U5650 (N_5650,N_4007,N_142);
or U5651 (N_5651,N_4728,N_3080);
and U5652 (N_5652,N_2485,N_3847);
nor U5653 (N_5653,N_4134,N_2274);
or U5654 (N_5654,N_860,N_3993);
nor U5655 (N_5655,N_1558,N_2148);
nand U5656 (N_5656,N_4343,N_617);
and U5657 (N_5657,N_3664,N_435);
and U5658 (N_5658,N_399,N_634);
or U5659 (N_5659,N_52,N_3587);
nor U5660 (N_5660,N_483,N_3932);
nor U5661 (N_5661,N_1014,N_2566);
and U5662 (N_5662,N_4981,N_1914);
nor U5663 (N_5663,N_724,N_1994);
and U5664 (N_5664,N_3578,N_1316);
nand U5665 (N_5665,N_3840,N_1747);
nand U5666 (N_5666,N_621,N_4594);
nand U5667 (N_5667,N_1987,N_2989);
or U5668 (N_5668,N_3412,N_2177);
and U5669 (N_5669,N_1130,N_2176);
and U5670 (N_5670,N_3247,N_2467);
and U5671 (N_5671,N_2986,N_4587);
and U5672 (N_5672,N_2212,N_2015);
nand U5673 (N_5673,N_531,N_4696);
or U5674 (N_5674,N_4970,N_796);
or U5675 (N_5675,N_379,N_1680);
xor U5676 (N_5676,N_3348,N_2113);
nor U5677 (N_5677,N_3254,N_2892);
and U5678 (N_5678,N_2192,N_3432);
nor U5679 (N_5679,N_1206,N_2363);
xor U5680 (N_5680,N_4630,N_3295);
and U5681 (N_5681,N_902,N_913);
nor U5682 (N_5682,N_4098,N_3047);
nand U5683 (N_5683,N_1088,N_3763);
and U5684 (N_5684,N_303,N_995);
or U5685 (N_5685,N_1515,N_4712);
nor U5686 (N_5686,N_4841,N_2315);
and U5687 (N_5687,N_3448,N_2832);
and U5688 (N_5688,N_2474,N_2964);
nand U5689 (N_5689,N_2487,N_231);
nor U5690 (N_5690,N_1590,N_947);
nor U5691 (N_5691,N_2746,N_3334);
nand U5692 (N_5692,N_124,N_4962);
nand U5693 (N_5693,N_4108,N_4877);
nor U5694 (N_5694,N_4019,N_4441);
nand U5695 (N_5695,N_702,N_2652);
and U5696 (N_5696,N_4163,N_3417);
nor U5697 (N_5697,N_4277,N_3857);
and U5698 (N_5698,N_850,N_779);
nand U5699 (N_5699,N_2992,N_498);
or U5700 (N_5700,N_972,N_1731);
or U5701 (N_5701,N_1783,N_1050);
nor U5702 (N_5702,N_1477,N_4544);
or U5703 (N_5703,N_4969,N_257);
nand U5704 (N_5704,N_1613,N_3715);
nand U5705 (N_5705,N_4476,N_119);
or U5706 (N_5706,N_3276,N_2903);
or U5707 (N_5707,N_2799,N_3030);
nor U5708 (N_5708,N_4259,N_4191);
or U5709 (N_5709,N_2758,N_3457);
and U5710 (N_5710,N_2269,N_3091);
nand U5711 (N_5711,N_3858,N_2909);
xnor U5712 (N_5712,N_2082,N_4946);
and U5713 (N_5713,N_3936,N_1735);
nor U5714 (N_5714,N_2477,N_2358);
and U5715 (N_5715,N_4561,N_2534);
xnor U5716 (N_5716,N_4548,N_824);
nand U5717 (N_5717,N_1566,N_1321);
nand U5718 (N_5718,N_4167,N_4492);
xor U5719 (N_5719,N_4592,N_283);
nand U5720 (N_5720,N_3550,N_2678);
or U5721 (N_5721,N_956,N_1290);
nand U5722 (N_5722,N_1345,N_3633);
or U5723 (N_5723,N_4673,N_2900);
or U5724 (N_5724,N_3896,N_3326);
and U5725 (N_5725,N_1526,N_3069);
or U5726 (N_5726,N_4989,N_1995);
or U5727 (N_5727,N_3743,N_91);
or U5728 (N_5728,N_1809,N_4686);
nand U5729 (N_5729,N_783,N_3744);
and U5730 (N_5730,N_2983,N_1750);
or U5731 (N_5731,N_3341,N_1784);
and U5732 (N_5732,N_1715,N_4142);
and U5733 (N_5733,N_1442,N_4425);
xnor U5734 (N_5734,N_3895,N_3476);
xor U5735 (N_5735,N_411,N_2384);
or U5736 (N_5736,N_663,N_1448);
or U5737 (N_5737,N_3390,N_1368);
nand U5738 (N_5738,N_3499,N_2562);
or U5739 (N_5739,N_11,N_3103);
and U5740 (N_5740,N_287,N_131);
and U5741 (N_5741,N_2488,N_1651);
nor U5742 (N_5742,N_2002,N_4840);
nand U5743 (N_5743,N_1257,N_4003);
or U5744 (N_5744,N_1705,N_2952);
nor U5745 (N_5745,N_34,N_3057);
xor U5746 (N_5746,N_3087,N_3111);
xor U5747 (N_5747,N_2781,N_2154);
and U5748 (N_5748,N_2227,N_4716);
and U5749 (N_5749,N_4251,N_3910);
nand U5750 (N_5750,N_403,N_3243);
xor U5751 (N_5751,N_4385,N_3698);
or U5752 (N_5752,N_3722,N_3089);
nand U5753 (N_5753,N_2597,N_589);
xnor U5754 (N_5754,N_4321,N_3218);
nand U5755 (N_5755,N_3399,N_4943);
nand U5756 (N_5756,N_4282,N_3545);
and U5757 (N_5757,N_4765,N_3264);
nor U5758 (N_5758,N_976,N_4845);
nor U5759 (N_5759,N_3475,N_2275);
nand U5760 (N_5760,N_2417,N_1546);
xor U5761 (N_5761,N_3222,N_402);
nand U5762 (N_5762,N_1545,N_1017);
and U5763 (N_5763,N_2272,N_3126);
xor U5764 (N_5764,N_217,N_2836);
xnor U5765 (N_5765,N_4868,N_3795);
xnor U5766 (N_5766,N_9,N_2236);
xnor U5767 (N_5767,N_2924,N_2127);
and U5768 (N_5768,N_3289,N_2270);
nand U5769 (N_5769,N_1867,N_609);
nor U5770 (N_5770,N_3033,N_4320);
and U5771 (N_5771,N_2153,N_2579);
and U5772 (N_5772,N_1858,N_3864);
xor U5773 (N_5773,N_802,N_2965);
xor U5774 (N_5774,N_2865,N_4043);
and U5775 (N_5775,N_2238,N_1301);
and U5776 (N_5776,N_3505,N_3856);
nand U5777 (N_5777,N_4158,N_2202);
xnor U5778 (N_5778,N_4401,N_2671);
xnor U5779 (N_5779,N_143,N_2368);
xnor U5780 (N_5780,N_181,N_4196);
nor U5781 (N_5781,N_2118,N_357);
or U5782 (N_5782,N_3519,N_4485);
xor U5783 (N_5783,N_711,N_3196);
xor U5784 (N_5784,N_2556,N_2430);
nand U5785 (N_5785,N_423,N_3005);
nand U5786 (N_5786,N_4447,N_3249);
and U5787 (N_5787,N_4945,N_2911);
nand U5788 (N_5788,N_4792,N_3115);
and U5789 (N_5789,N_2823,N_288);
or U5790 (N_5790,N_564,N_3122);
or U5791 (N_5791,N_193,N_98);
xnor U5792 (N_5792,N_2544,N_1818);
nand U5793 (N_5793,N_4545,N_4112);
nor U5794 (N_5794,N_1793,N_3055);
xor U5795 (N_5795,N_4075,N_1694);
nand U5796 (N_5796,N_4155,N_200);
nor U5797 (N_5797,N_2513,N_4503);
xor U5798 (N_5798,N_453,N_273);
nor U5799 (N_5799,N_3300,N_127);
and U5800 (N_5800,N_728,N_2323);
and U5801 (N_5801,N_4929,N_1302);
nor U5802 (N_5802,N_1860,N_133);
and U5803 (N_5803,N_4138,N_818);
or U5804 (N_5804,N_3622,N_3943);
xor U5805 (N_5805,N_3979,N_989);
nor U5806 (N_5806,N_2351,N_2410);
or U5807 (N_5807,N_71,N_3593);
or U5808 (N_5808,N_4235,N_2769);
xor U5809 (N_5809,N_452,N_3262);
nand U5810 (N_5810,N_4024,N_4403);
and U5811 (N_5811,N_2350,N_449);
nand U5812 (N_5812,N_1652,N_2372);
nand U5813 (N_5813,N_2614,N_3646);
xnor U5814 (N_5814,N_105,N_1561);
xor U5815 (N_5815,N_2233,N_2459);
and U5816 (N_5816,N_2161,N_43);
nor U5817 (N_5817,N_1724,N_294);
xor U5818 (N_5818,N_1877,N_1967);
xor U5819 (N_5819,N_645,N_3136);
and U5820 (N_5820,N_2457,N_3786);
nand U5821 (N_5821,N_4412,N_4440);
xor U5822 (N_5822,N_2428,N_1946);
nand U5823 (N_5823,N_3425,N_2551);
and U5824 (N_5824,N_20,N_2803);
xor U5825 (N_5825,N_3162,N_3071);
or U5826 (N_5826,N_3620,N_1484);
and U5827 (N_5827,N_1514,N_4793);
nor U5828 (N_5828,N_4311,N_4283);
or U5829 (N_5829,N_2303,N_1565);
nand U5830 (N_5830,N_3282,N_1211);
nand U5831 (N_5831,N_4358,N_64);
nor U5832 (N_5832,N_4481,N_542);
nor U5833 (N_5833,N_2365,N_185);
or U5834 (N_5834,N_4953,N_37);
and U5835 (N_5835,N_4374,N_4300);
nor U5836 (N_5836,N_3309,N_485);
or U5837 (N_5837,N_687,N_1095);
and U5838 (N_5838,N_1440,N_1534);
nor U5839 (N_5839,N_2738,N_4789);
xnor U5840 (N_5840,N_927,N_102);
nand U5841 (N_5841,N_1532,N_2749);
and U5842 (N_5842,N_4232,N_4680);
xor U5843 (N_5843,N_3583,N_2629);
or U5844 (N_5844,N_546,N_4445);
xnor U5845 (N_5845,N_2468,N_3209);
nand U5846 (N_5846,N_2568,N_2186);
or U5847 (N_5847,N_4688,N_3245);
xnor U5848 (N_5848,N_3782,N_4104);
or U5849 (N_5849,N_3173,N_1703);
xnor U5850 (N_5850,N_2353,N_3219);
and U5851 (N_5851,N_455,N_529);
nor U5852 (N_5852,N_3672,N_1122);
xor U5853 (N_5853,N_1175,N_2856);
and U5854 (N_5854,N_2960,N_3461);
and U5855 (N_5855,N_359,N_2742);
nor U5856 (N_5856,N_2507,N_4566);
xnor U5857 (N_5857,N_579,N_2730);
nor U5858 (N_5858,N_2731,N_1403);
and U5859 (N_5859,N_3176,N_4082);
xor U5860 (N_5860,N_882,N_1708);
nor U5861 (N_5861,N_1602,N_3994);
and U5862 (N_5862,N_4944,N_642);
xnor U5863 (N_5863,N_2408,N_1114);
or U5864 (N_5864,N_3131,N_2768);
xor U5865 (N_5865,N_657,N_1346);
nor U5866 (N_5866,N_2713,N_2651);
nor U5867 (N_5867,N_599,N_1512);
or U5868 (N_5868,N_4473,N_3509);
xnor U5869 (N_5869,N_1648,N_2542);
xnor U5870 (N_5870,N_4794,N_3255);
or U5871 (N_5871,N_3608,N_4963);
xnor U5872 (N_5872,N_4365,N_2253);
or U5873 (N_5873,N_2167,N_1458);
nor U5874 (N_5874,N_141,N_2531);
and U5875 (N_5875,N_1927,N_4768);
or U5876 (N_5876,N_2260,N_2234);
and U5877 (N_5877,N_2985,N_793);
nand U5878 (N_5878,N_1684,N_2398);
and U5879 (N_5879,N_4611,N_1749);
nor U5880 (N_5880,N_3572,N_1040);
nor U5881 (N_5881,N_4633,N_4010);
nand U5882 (N_5882,N_3168,N_946);
xor U5883 (N_5883,N_4310,N_4955);
or U5884 (N_5884,N_1035,N_5);
or U5885 (N_5885,N_4392,N_168);
nand U5886 (N_5886,N_4562,N_3788);
nand U5887 (N_5887,N_1020,N_3954);
and U5888 (N_5888,N_4926,N_1141);
or U5889 (N_5889,N_868,N_1801);
or U5890 (N_5890,N_2362,N_1277);
or U5891 (N_5891,N_1504,N_2171);
nor U5892 (N_5892,N_2370,N_2355);
or U5893 (N_5893,N_3000,N_4470);
and U5894 (N_5894,N_2073,N_89);
nand U5895 (N_5895,N_1116,N_4306);
or U5896 (N_5896,N_1436,N_4256);
and U5897 (N_5897,N_1071,N_4760);
nor U5898 (N_5898,N_4363,N_3045);
nand U5899 (N_5899,N_1213,N_3297);
xnor U5900 (N_5900,N_536,N_3441);
and U5901 (N_5901,N_2889,N_1537);
nand U5902 (N_5902,N_4414,N_2201);
or U5903 (N_5903,N_1598,N_623);
xnor U5904 (N_5904,N_4453,N_797);
or U5905 (N_5905,N_3590,N_3335);
nor U5906 (N_5906,N_2518,N_856);
or U5907 (N_5907,N_4972,N_3349);
xnor U5908 (N_5908,N_3753,N_4079);
nand U5909 (N_5909,N_3129,N_2880);
and U5910 (N_5910,N_1836,N_194);
nand U5911 (N_5911,N_2868,N_4130);
xnor U5912 (N_5912,N_1312,N_3639);
nor U5913 (N_5913,N_4621,N_2290);
xnor U5914 (N_5914,N_3251,N_1587);
nand U5915 (N_5915,N_361,N_174);
xnor U5916 (N_5916,N_3826,N_2434);
and U5917 (N_5917,N_2572,N_3140);
and U5918 (N_5918,N_2591,N_3164);
xor U5919 (N_5919,N_820,N_4181);
nand U5920 (N_5920,N_3225,N_1043);
nor U5921 (N_5921,N_150,N_4523);
nor U5922 (N_5922,N_2451,N_1574);
or U5923 (N_5923,N_122,N_4752);
xnor U5924 (N_5924,N_1379,N_2273);
xor U5925 (N_5925,N_4239,N_2043);
and U5926 (N_5926,N_3350,N_1355);
nand U5927 (N_5927,N_2828,N_177);
xnor U5928 (N_5928,N_3285,N_1511);
nand U5929 (N_5929,N_3642,N_3101);
or U5930 (N_5930,N_3774,N_1098);
nor U5931 (N_5931,N_4909,N_3597);
or U5932 (N_5932,N_572,N_1959);
nor U5933 (N_5933,N_842,N_2688);
and U5934 (N_5934,N_1499,N_1645);
nor U5935 (N_5935,N_1283,N_4665);
or U5936 (N_5936,N_3966,N_3066);
and U5937 (N_5937,N_1372,N_3876);
nand U5938 (N_5938,N_3908,N_1882);
xnor U5939 (N_5939,N_2285,N_2146);
or U5940 (N_5940,N_3790,N_4288);
nor U5941 (N_5941,N_750,N_2930);
xnor U5942 (N_5942,N_1752,N_1240);
xnor U5943 (N_5943,N_4597,N_4709);
nor U5944 (N_5944,N_3758,N_2121);
nand U5945 (N_5945,N_886,N_342);
nand U5946 (N_5946,N_337,N_115);
xor U5947 (N_5947,N_145,N_266);
and U5948 (N_5948,N_2510,N_3239);
xnor U5949 (N_5949,N_3035,N_476);
nor U5950 (N_5950,N_2630,N_1908);
nand U5951 (N_5951,N_2390,N_1156);
nor U5952 (N_5952,N_4646,N_853);
and U5953 (N_5953,N_993,N_1913);
nor U5954 (N_5954,N_3838,N_2223);
nand U5955 (N_5955,N_1444,N_2320);
nand U5956 (N_5956,N_1984,N_312);
xnor U5957 (N_5957,N_945,N_2387);
or U5958 (N_5958,N_3952,N_3439);
nand U5959 (N_5959,N_153,N_3371);
or U5960 (N_5960,N_3459,N_4638);
and U5961 (N_5961,N_1449,N_2771);
nor U5962 (N_5962,N_984,N_2521);
or U5963 (N_5963,N_235,N_4674);
nand U5964 (N_5964,N_4313,N_4823);
nor U5965 (N_5965,N_4843,N_1341);
or U5966 (N_5966,N_2458,N_4679);
nor U5967 (N_5967,N_1854,N_3469);
and U5968 (N_5968,N_2220,N_4045);
nor U5969 (N_5969,N_48,N_3735);
nor U5970 (N_5970,N_1432,N_533);
nand U5971 (N_5971,N_1510,N_2929);
xor U5972 (N_5972,N_4391,N_128);
xor U5973 (N_5973,N_2180,N_4193);
nor U5974 (N_5974,N_911,N_1736);
nand U5975 (N_5975,N_3205,N_851);
or U5976 (N_5976,N_3791,N_4056);
nand U5977 (N_5977,N_1721,N_1616);
and U5978 (N_5978,N_1728,N_3824);
nor U5979 (N_5979,N_1524,N_1644);
nor U5980 (N_5980,N_4100,N_2684);
xor U5981 (N_5981,N_1786,N_2090);
and U5982 (N_5982,N_4302,N_2076);
or U5983 (N_5983,N_1554,N_4337);
and U5984 (N_5984,N_1591,N_2776);
or U5985 (N_5985,N_2240,N_2744);
xnor U5986 (N_5986,N_3946,N_756);
or U5987 (N_5987,N_2169,N_2990);
nand U5988 (N_5988,N_2246,N_751);
nand U5989 (N_5989,N_2792,N_1064);
nand U5990 (N_5990,N_2595,N_969);
xor U5991 (N_5991,N_3463,N_1081);
and U5992 (N_5992,N_4435,N_2907);
xor U5993 (N_5993,N_2940,N_4683);
or U5994 (N_5994,N_2392,N_3995);
nand U5995 (N_5995,N_957,N_3148);
or U5996 (N_5996,N_2433,N_2853);
and U5997 (N_5997,N_3796,N_1398);
xnor U5998 (N_5998,N_1427,N_4717);
and U5999 (N_5999,N_3296,N_1412);
nand U6000 (N_6000,N_771,N_2452);
or U6001 (N_6001,N_3996,N_1939);
nor U6002 (N_6002,N_2276,N_1658);
nor U6003 (N_6003,N_2155,N_1409);
nor U6004 (N_6004,N_416,N_3128);
xnor U6005 (N_6005,N_2857,N_4350);
and U6006 (N_6006,N_3284,N_4617);
xnor U6007 (N_6007,N_1013,N_2376);
xor U6008 (N_6008,N_2085,N_466);
nand U6009 (N_6009,N_1459,N_3580);
and U6010 (N_6010,N_2848,N_1142);
or U6011 (N_6011,N_555,N_2339);
xnor U6012 (N_6012,N_1567,N_3382);
and U6013 (N_6013,N_4316,N_1058);
nor U6014 (N_6014,N_471,N_3925);
nor U6015 (N_6015,N_349,N_4052);
and U6016 (N_6016,N_1659,N_2515);
xor U6017 (N_6017,N_3266,N_4170);
and U6018 (N_6018,N_872,N_1635);
or U6019 (N_6019,N_2321,N_4501);
or U6020 (N_6020,N_3387,N_910);
nor U6021 (N_6021,N_695,N_865);
or U6022 (N_6022,N_241,N_4670);
or U6023 (N_6023,N_4199,N_1711);
or U6024 (N_6024,N_1337,N_2162);
or U6025 (N_6025,N_1527,N_3233);
nand U6026 (N_6026,N_2831,N_3524);
and U6027 (N_6027,N_2877,N_1307);
nor U6028 (N_6028,N_828,N_4172);
and U6029 (N_6029,N_170,N_3902);
and U6030 (N_6030,N_2649,N_341);
nand U6031 (N_6031,N_2751,N_4623);
or U6032 (N_6032,N_2530,N_2777);
xnor U6033 (N_6033,N_3268,N_4266);
nor U6034 (N_6034,N_2656,N_2048);
xor U6035 (N_6035,N_1516,N_4619);
xor U6036 (N_6036,N_4777,N_3528);
xor U6037 (N_6037,N_2904,N_3135);
and U6038 (N_6038,N_3670,N_3454);
or U6039 (N_6039,N_222,N_4318);
xnor U6040 (N_6040,N_4928,N_4018);
and U6041 (N_6041,N_2559,N_1624);
nand U6042 (N_6042,N_4095,N_4649);
or U6043 (N_6043,N_157,N_2445);
xnor U6044 (N_6044,N_4836,N_172);
and U6045 (N_6045,N_1224,N_2259);
or U6046 (N_6046,N_2931,N_4227);
nand U6047 (N_6047,N_1384,N_1208);
xnor U6048 (N_6048,N_1507,N_855);
nor U6049 (N_6049,N_4114,N_46);
nor U6050 (N_6050,N_979,N_4165);
nor U6051 (N_6051,N_650,N_260);
nand U6052 (N_6052,N_139,N_2588);
xnor U6053 (N_6053,N_582,N_1136);
nor U6054 (N_6054,N_3198,N_3579);
nor U6055 (N_6055,N_1300,N_3207);
nand U6056 (N_6056,N_1733,N_4978);
and U6057 (N_6057,N_769,N_4159);
or U6058 (N_6058,N_3175,N_674);
and U6059 (N_6059,N_2729,N_165);
and U6060 (N_6060,N_236,N_1344);
nor U6061 (N_6061,N_577,N_3330);
and U6062 (N_6062,N_4504,N_3797);
nor U6063 (N_6063,N_2680,N_3158);
and U6064 (N_6064,N_1767,N_4558);
nor U6065 (N_6065,N_4589,N_2708);
xor U6066 (N_6066,N_1900,N_2361);
or U6067 (N_6067,N_1188,N_3145);
and U6068 (N_6068,N_598,N_2674);
nor U6069 (N_6069,N_3391,N_4924);
nor U6070 (N_6070,N_2041,N_1905);
xor U6071 (N_6071,N_138,N_1878);
and U6072 (N_6072,N_1268,N_4001);
nor U6073 (N_6073,N_2512,N_1585);
xnor U6074 (N_6074,N_1294,N_39);
nor U6075 (N_6075,N_4761,N_1773);
or U6076 (N_6076,N_3898,N_2695);
xor U6077 (N_6077,N_3404,N_1404);
nor U6078 (N_6078,N_4161,N_4995);
xnor U6079 (N_6079,N_4087,N_3453);
nor U6080 (N_6080,N_2134,N_4057);
or U6081 (N_6081,N_2382,N_4345);
or U6082 (N_6082,N_3482,N_3313);
or U6083 (N_6083,N_2619,N_4081);
nor U6084 (N_6084,N_3188,N_4971);
nor U6085 (N_6085,N_3543,N_1004);
xnor U6086 (N_6086,N_1447,N_3234);
xor U6087 (N_6087,N_1123,N_480);
nor U6088 (N_6088,N_1261,N_675);
nand U6089 (N_6089,N_2022,N_4423);
and U6090 (N_6090,N_3014,N_2663);
nand U6091 (N_6091,N_4332,N_2074);
or U6092 (N_6092,N_1918,N_2922);
nand U6093 (N_6093,N_2639,N_847);
nand U6094 (N_6094,N_1204,N_1799);
xor U6095 (N_6095,N_4849,N_2063);
xnor U6096 (N_6096,N_3576,N_1126);
or U6097 (N_6097,N_809,N_14);
nor U6098 (N_6098,N_3843,N_4260);
nor U6099 (N_6099,N_3556,N_1297);
or U6100 (N_6100,N_2750,N_622);
nor U6101 (N_6101,N_4988,N_1022);
nand U6102 (N_6102,N_2819,N_1291);
nor U6103 (N_6103,N_1323,N_1985);
or U6104 (N_6104,N_4616,N_1350);
and U6105 (N_6105,N_968,N_3596);
and U6106 (N_6106,N_3216,N_925);
nor U6107 (N_6107,N_4276,N_2826);
nor U6108 (N_6108,N_3854,N_3967);
xnor U6109 (N_6109,N_2087,N_4739);
and U6110 (N_6110,N_4691,N_4422);
nor U6111 (N_6111,N_3144,N_1897);
and U6112 (N_6112,N_2080,N_1255);
xnor U6113 (N_6113,N_4848,N_2635);
nand U6114 (N_6114,N_3060,N_2136);
nor U6115 (N_6115,N_3372,N_3141);
or U6116 (N_6116,N_4049,N_4706);
and U6117 (N_6117,N_1933,N_4344);
or U6118 (N_6118,N_58,N_3379);
xnor U6119 (N_6119,N_1056,N_3017);
or U6120 (N_6120,N_4958,N_1150);
or U6121 (N_6121,N_798,N_497);
nand U6122 (N_6122,N_3496,N_426);
and U6123 (N_6123,N_1170,N_1997);
nand U6124 (N_6124,N_2484,N_3202);
nor U6125 (N_6125,N_317,N_550);
nand U6126 (N_6126,N_334,N_1250);
or U6127 (N_6127,N_4697,N_4177);
nor U6128 (N_6128,N_3734,N_3075);
xor U6129 (N_6129,N_4838,N_4564);
and U6130 (N_6130,N_56,N_4329);
or U6131 (N_6131,N_3957,N_4719);
and U6132 (N_6132,N_2224,N_3292);
nor U6133 (N_6133,N_4072,N_2897);
nor U6134 (N_6134,N_1419,N_1438);
and U6135 (N_6135,N_4387,N_1993);
xor U6136 (N_6136,N_889,N_714);
nor U6137 (N_6137,N_2401,N_1303);
xnor U6138 (N_6138,N_4162,N_4824);
nor U6139 (N_6139,N_2097,N_3900);
and U6140 (N_6140,N_1674,N_81);
xnor U6141 (N_6141,N_2642,N_4571);
nand U6142 (N_6142,N_371,N_4073);
nor U6143 (N_6143,N_1079,N_2855);
nand U6144 (N_6144,N_3396,N_4096);
nand U6145 (N_6145,N_4647,N_1317);
nand U6146 (N_6146,N_1244,N_4738);
and U6147 (N_6147,N_1107,N_2875);
nand U6148 (N_6148,N_1333,N_2416);
nand U6149 (N_6149,N_1691,N_4123);
or U6150 (N_6150,N_3777,N_3600);
or U6151 (N_6151,N_392,N_3281);
nor U6152 (N_6152,N_775,N_3214);
nand U6153 (N_6153,N_2594,N_2538);
nor U6154 (N_6154,N_353,N_4595);
or U6155 (N_6155,N_4599,N_4483);
nand U6156 (N_6156,N_1151,N_1884);
nor U6157 (N_6157,N_2083,N_4028);
nor U6158 (N_6158,N_2096,N_2577);
nor U6159 (N_6159,N_1582,N_1544);
nor U6160 (N_6160,N_2980,N_1928);
and U6161 (N_6161,N_367,N_2095);
and U6162 (N_6162,N_4855,N_3223);
nand U6163 (N_6163,N_3690,N_967);
nand U6164 (N_6164,N_2928,N_4415);
nand U6165 (N_6165,N_915,N_1024);
nor U6166 (N_6166,N_2399,N_3241);
nand U6167 (N_6167,N_12,N_316);
nor U6168 (N_6168,N_17,N_4903);
xor U6169 (N_6169,N_2021,N_1181);
nand U6170 (N_6170,N_4977,N_3004);
nand U6171 (N_6171,N_344,N_4578);
nand U6172 (N_6172,N_3974,N_933);
xnor U6173 (N_6173,N_921,N_3935);
nand U6174 (N_6174,N_4246,N_4389);
xnor U6175 (N_6175,N_2582,N_2524);
and U6176 (N_6176,N_3537,N_3152);
xor U6177 (N_6177,N_2062,N_1656);
nand U6178 (N_6178,N_3428,N_3872);
nand U6179 (N_6179,N_2093,N_3628);
xor U6180 (N_6180,N_1464,N_4189);
and U6181 (N_6181,N_401,N_571);
or U6182 (N_6182,N_1823,N_4292);
and U6183 (N_6183,N_2464,N_554);
or U6184 (N_6184,N_3693,N_1121);
nand U6185 (N_6185,N_2126,N_4538);
xnor U6186 (N_6186,N_3844,N_3762);
xnor U6187 (N_6187,N_2141,N_3286);
and U6188 (N_6188,N_4154,N_3310);
or U6189 (N_6189,N_3793,N_2425);
nor U6190 (N_6190,N_671,N_513);
or U6191 (N_6191,N_1795,N_774);
xnor U6192 (N_6192,N_4757,N_495);
and U6193 (N_6193,N_4421,N_484);
nand U6194 (N_6194,N_474,N_2207);
nor U6195 (N_6195,N_1553,N_4145);
nand U6196 (N_6196,N_398,N_3613);
nor U6197 (N_6197,N_1293,N_4496);
nand U6198 (N_6198,N_4141,N_3897);
nor U6199 (N_6199,N_3980,N_1469);
nand U6200 (N_6200,N_3929,N_3999);
xor U6201 (N_6201,N_2636,N_3450);
nand U6202 (N_6202,N_2110,N_591);
or U6203 (N_6203,N_3868,N_1766);
nand U6204 (N_6204,N_907,N_1435);
nor U6205 (N_6205,N_2968,N_3875);
nor U6206 (N_6206,N_4216,N_3883);
nand U6207 (N_6207,N_1760,N_3942);
xnor U6208 (N_6208,N_1475,N_121);
and U6209 (N_6209,N_1400,N_4091);
nand U6210 (N_6210,N_2061,N_1177);
xnor U6211 (N_6211,N_1145,N_1697);
nand U6212 (N_6212,N_1353,N_3640);
and U6213 (N_6213,N_971,N_2187);
xor U6214 (N_6214,N_2437,N_1146);
xor U6215 (N_6215,N_4510,N_272);
nand U6216 (N_6216,N_1377,N_2175);
xnor U6217 (N_6217,N_3395,N_1945);
xor U6218 (N_6218,N_1231,N_299);
or U6219 (N_6219,N_3915,N_4865);
and U6220 (N_6220,N_1789,N_1679);
or U6221 (N_6221,N_1816,N_4520);
nand U6222 (N_6222,N_3181,N_2852);
and U6223 (N_6223,N_615,N_3037);
nor U6224 (N_6224,N_608,N_4930);
and U6225 (N_6225,N_1726,N_4692);
or U6226 (N_6226,N_749,N_101);
and U6227 (N_6227,N_3555,N_1147);
nor U6228 (N_6228,N_1201,N_4157);
and U6229 (N_6229,N_4240,N_2205);
nor U6230 (N_6230,N_148,N_772);
nor U6231 (N_6231,N_409,N_4961);
nand U6232 (N_6232,N_4788,N_2415);
xnor U6233 (N_6233,N_2913,N_918);
xor U6234 (N_6234,N_3709,N_1889);
nand U6235 (N_6235,N_3903,N_2941);
or U6236 (N_6236,N_3958,N_4015);
xor U6237 (N_6237,N_1893,N_245);
or U6238 (N_6238,N_2982,N_3018);
nand U6239 (N_6239,N_1830,N_61);
xnor U6240 (N_6240,N_1579,N_1956);
and U6241 (N_6241,N_4627,N_4986);
xor U6242 (N_6242,N_3447,N_3159);
nand U6243 (N_6243,N_4883,N_4711);
and U6244 (N_6244,N_1646,N_93);
and U6245 (N_6245,N_4826,N_3530);
nand U6246 (N_6246,N_4448,N_859);
nand U6247 (N_6247,N_2481,N_2839);
and U6248 (N_6248,N_4828,N_2773);
and U6249 (N_6249,N_247,N_1491);
xor U6250 (N_6250,N_2879,N_1445);
nor U6251 (N_6251,N_1920,N_3816);
and U6252 (N_6252,N_1940,N_2753);
and U6253 (N_6253,N_2117,N_1279);
nand U6254 (N_6254,N_1153,N_1943);
nor U6255 (N_6255,N_44,N_4542);
nor U6256 (N_6256,N_1839,N_3841);
nor U6257 (N_6257,N_4763,N_4042);
nor U6258 (N_6258,N_807,N_4204);
or U6259 (N_6259,N_1466,N_4912);
xnor U6260 (N_6260,N_3659,N_3409);
nor U6261 (N_6261,N_437,N_764);
xnor U6262 (N_6262,N_1325,N_2294);
xor U6263 (N_6263,N_4333,N_1405);
xnor U6264 (N_6264,N_901,N_3036);
xor U6265 (N_6265,N_1386,N_369);
nor U6266 (N_6266,N_4219,N_4648);
xor U6267 (N_6267,N_4811,N_4821);
or U6268 (N_6268,N_3736,N_4382);
nor U6269 (N_6269,N_3899,N_4721);
nand U6270 (N_6270,N_3403,N_4160);
nor U6271 (N_6271,N_2605,N_718);
and U6272 (N_6272,N_3238,N_581);
and U6273 (N_6273,N_4540,N_487);
or U6274 (N_6274,N_1901,N_874);
or U6275 (N_6275,N_4901,N_4265);
nand U6276 (N_6276,N_4722,N_518);
nor U6277 (N_6277,N_336,N_1029);
nor U6278 (N_6278,N_1977,N_4803);
nor U6279 (N_6279,N_3531,N_2932);
nand U6280 (N_6280,N_2541,N_873);
and U6281 (N_6281,N_990,N_676);
nand U6282 (N_6282,N_2168,N_2055);
nand U6283 (N_6283,N_4975,N_1930);
and U6284 (N_6284,N_876,N_4449);
and U6285 (N_6285,N_2810,N_944);
xor U6286 (N_6286,N_2211,N_3470);
or U6287 (N_6287,N_1745,N_3086);
or U6288 (N_6288,N_3937,N_118);
or U6289 (N_6289,N_2571,N_67);
nand U6290 (N_6290,N_4749,N_2885);
xor U6291 (N_6291,N_4644,N_4825);
and U6292 (N_6292,N_607,N_4610);
or U6293 (N_6293,N_4179,N_4491);
nand U6294 (N_6294,N_3721,N_977);
or U6295 (N_6295,N_2867,N_1937);
nand U6296 (N_6296,N_1664,N_4913);
nand U6297 (N_6297,N_4497,N_3385);
xor U6298 (N_6298,N_504,N_1167);
xnor U6299 (N_6299,N_3051,N_4585);
xor U6300 (N_6300,N_4687,N_4762);
xnor U6301 (N_6301,N_2172,N_4812);
xor U6302 (N_6302,N_2182,N_3859);
nor U6303 (N_6303,N_3381,N_1319);
nor U6304 (N_6304,N_3430,N_2737);
or U6305 (N_6305,N_3464,N_192);
xnor U6306 (N_6306,N_413,N_1179);
nand U6307 (N_6307,N_566,N_112);
xnor U6308 (N_6308,N_1807,N_2693);
or U6309 (N_6309,N_4419,N_1626);
or U6310 (N_6310,N_4467,N_73);
and U6311 (N_6311,N_2607,N_26);
or U6312 (N_6312,N_3375,N_3151);
xnor U6313 (N_6313,N_41,N_3065);
nand U6314 (N_6314,N_3077,N_2426);
nor U6315 (N_6315,N_3431,N_4245);
or U6316 (N_6316,N_215,N_1248);
xnor U6317 (N_6317,N_3337,N_224);
nand U6318 (N_6318,N_1580,N_1327);
nor U6319 (N_6319,N_1653,N_391);
and U6320 (N_6320,N_2679,N_760);
nand U6321 (N_6321,N_1952,N_226);
xor U6322 (N_6322,N_3197,N_3718);
or U6323 (N_6323,N_10,N_2301);
or U6324 (N_6324,N_1260,N_2250);
nand U6325 (N_6325,N_2453,N_151);
nand U6326 (N_6326,N_3083,N_135);
nor U6327 (N_6327,N_673,N_3426);
nor U6328 (N_6328,N_3109,N_961);
and U6329 (N_6329,N_4991,N_792);
and U6330 (N_6330,N_94,N_1135);
nand U6331 (N_6331,N_2489,N_745);
nor U6332 (N_6332,N_2816,N_4900);
and U6333 (N_6333,N_2278,N_3194);
xor U6334 (N_6334,N_1973,N_4022);
or U6335 (N_6335,N_875,N_3582);
nor U6336 (N_6336,N_1378,N_4489);
or U6337 (N_6337,N_4388,N_1476);
or U6338 (N_6338,N_678,N_1117);
nand U6339 (N_6339,N_3253,N_4353);
xor U6340 (N_6340,N_3153,N_787);
and U6341 (N_6341,N_2975,N_4424);
and U6342 (N_6342,N_1092,N_4198);
or U6343 (N_6343,N_2047,N_1195);
nand U6344 (N_6344,N_2767,N_4249);
nand U6345 (N_6345,N_4197,N_2374);
xnor U6346 (N_6346,N_1452,N_4645);
or U6347 (N_6347,N_491,N_628);
or U6348 (N_6348,N_2715,N_2994);
nand U6349 (N_6349,N_761,N_2756);
xnor U6350 (N_6350,N_4726,N_302);
nor U6351 (N_6351,N_479,N_4008);
xnor U6352 (N_6352,N_583,N_777);
nor U6353 (N_6353,N_459,N_1589);
nor U6354 (N_6354,N_4287,N_4980);
nand U6355 (N_6355,N_83,N_1110);
nand U6356 (N_6356,N_4274,N_3024);
nor U6357 (N_6357,N_2313,N_4361);
or U6358 (N_6358,N_4586,N_3189);
xor U6359 (N_6359,N_733,N_2204);
nand U6360 (N_6360,N_4164,N_4846);
and U6361 (N_6361,N_4281,N_42);
nand U6362 (N_6362,N_1401,N_1468);
nand U6363 (N_6363,N_3829,N_632);
xnor U6364 (N_6364,N_4796,N_903);
nor U6365 (N_6365,N_393,N_3318);
xnor U6366 (N_6366,N_1467,N_1052);
xor U6367 (N_6367,N_211,N_1465);
nand U6368 (N_6368,N_2214,N_2565);
or U6369 (N_6369,N_3221,N_1414);
and U6370 (N_6370,N_111,N_1120);
xnor U6371 (N_6371,N_3688,N_1164);
nand U6372 (N_6372,N_4815,N_1774);
nor U6373 (N_6373,N_3617,N_4517);
nand U6374 (N_6374,N_3514,N_4583);
xor U6375 (N_6375,N_30,N_4737);
or U6376 (N_6376,N_661,N_1048);
or U6377 (N_6377,N_3070,N_1964);
and U6378 (N_6378,N_1718,N_3890);
and U6379 (N_6379,N_2279,N_2486);
nor U6380 (N_6380,N_3178,N_3945);
or U6381 (N_6381,N_2662,N_314);
xor U6382 (N_6382,N_2840,N_4413);
nand U6383 (N_6383,N_4475,N_1543);
nor U6384 (N_6384,N_4776,N_2077);
and U6385 (N_6385,N_916,N_3301);
nand U6386 (N_6386,N_3046,N_3566);
xnor U6387 (N_6387,N_551,N_3783);
nand U6388 (N_6388,N_2796,N_2418);
and U6389 (N_6389,N_156,N_79);
xnor U6390 (N_6390,N_4488,N_2283);
nor U6391 (N_6391,N_3369,N_3134);
nor U6392 (N_6392,N_3842,N_3880);
or U6393 (N_6393,N_4731,N_470);
and U6394 (N_6394,N_3754,N_2560);
nand U6395 (N_6395,N_4175,N_4654);
nand U6396 (N_6396,N_4898,N_252);
and U6397 (N_6397,N_4973,N_2603);
nor U6398 (N_6398,N_1251,N_1078);
xor U6399 (N_6399,N_4433,N_4536);
nand U6400 (N_6400,N_3606,N_3081);
xor U6401 (N_6401,N_2570,N_4695);
or U6402 (N_6402,N_707,N_3220);
nor U6403 (N_6403,N_350,N_370);
xor U6404 (N_6404,N_95,N_2436);
and U6405 (N_6405,N_1239,N_1492);
or U6406 (N_6406,N_2546,N_3813);
or U6407 (N_6407,N_1979,N_3959);
nand U6408 (N_6408,N_3766,N_268);
nor U6409 (N_6409,N_3169,N_2687);
or U6410 (N_6410,N_4223,N_1906);
or U6411 (N_6411,N_2710,N_4518);
or U6412 (N_6412,N_4635,N_578);
nand U6413 (N_6413,N_420,N_2851);
and U6414 (N_6414,N_844,N_1219);
xnor U6415 (N_6415,N_3408,N_4818);
xnor U6416 (N_6416,N_2520,N_3257);
and U6417 (N_6417,N_3665,N_490);
nand U6418 (N_6418,N_4370,N_4205);
nand U6419 (N_6419,N_3603,N_1907);
and U6420 (N_6420,N_2400,N_3402);
or U6421 (N_6421,N_4755,N_1535);
nand U6422 (N_6422,N_3479,N_3193);
and U6423 (N_6423,N_4064,N_1096);
nand U6424 (N_6424,N_3019,N_3001);
nand U6425 (N_6425,N_2244,N_999);
and U6426 (N_6426,N_2532,N_2439);
or U6427 (N_6427,N_747,N_3518);
nor U6428 (N_6428,N_2328,N_3759);
and U6429 (N_6429,N_1009,N_176);
xor U6430 (N_6430,N_4584,N_1792);
nor U6431 (N_6431,N_3685,N_1547);
nand U6432 (N_6432,N_3146,N_4921);
nand U6433 (N_6433,N_4748,N_3424);
and U6434 (N_6434,N_1028,N_2078);
nand U6435 (N_6435,N_4814,N_595);
xor U6436 (N_6436,N_2668,N_1138);
nand U6437 (N_6437,N_4118,N_4037);
and U6438 (N_6438,N_4500,N_3586);
or U6439 (N_6439,N_1596,N_3695);
nor U6440 (N_6440,N_4270,N_2667);
xnor U6441 (N_6441,N_1314,N_1376);
nand U6442 (N_6442,N_2034,N_4068);
or U6443 (N_6443,N_1701,N_4462);
nand U6444 (N_6444,N_100,N_146);
xor U6445 (N_6445,N_4454,N_265);
xnor U6446 (N_6446,N_1011,N_230);
nand U6447 (N_6447,N_660,N_4436);
and U6448 (N_6448,N_4593,N_2714);
or U6449 (N_6449,N_4998,N_4703);
or U6450 (N_6450,N_1881,N_1238);
xnor U6451 (N_6451,N_4315,N_1309);
xor U6452 (N_6452,N_1502,N_4376);
or U6453 (N_6453,N_408,N_478);
xor U6454 (N_6454,N_4375,N_3015);
xnor U6455 (N_6455,N_2051,N_3621);
nand U6456 (N_6456,N_653,N_106);
nand U6457 (N_6457,N_196,N_207);
or U6458 (N_6458,N_1202,N_385);
and U6459 (N_6459,N_3419,N_3873);
nor U6460 (N_6460,N_4787,N_3918);
nor U6461 (N_6461,N_823,N_4857);
nor U6462 (N_6462,N_2493,N_271);
nand U6463 (N_6463,N_4614,N_4873);
xnor U6464 (N_6464,N_2478,N_1902);
nand U6465 (N_6465,N_4125,N_1055);
and U6466 (N_6466,N_107,N_705);
nand U6467 (N_6467,N_4575,N_2760);
nor U6468 (N_6468,N_2257,N_4074);
nand U6469 (N_6469,N_3108,N_3107);
and U6470 (N_6470,N_685,N_206);
xnor U6471 (N_6471,N_1152,N_894);
or U6472 (N_6472,N_2346,N_3971);
xnor U6473 (N_6473,N_1494,N_2101);
nand U6474 (N_6474,N_1187,N_441);
xnor U6475 (N_6475,N_3323,N_4713);
nor U6476 (N_6476,N_1637,N_1610);
nand U6477 (N_6477,N_4974,N_4705);
nor U6478 (N_6478,N_3780,N_2336);
nor U6479 (N_6479,N_4377,N_3272);
nand U6480 (N_6480,N_4906,N_1904);
xnor U6481 (N_6481,N_1269,N_4017);
nor U6482 (N_6482,N_2774,N_2222);
xnor U6483 (N_6483,N_778,N_1641);
nand U6484 (N_6484,N_3792,N_1304);
and U6485 (N_6485,N_1791,N_2500);
and U6486 (N_6486,N_2277,N_3520);
nand U6487 (N_6487,N_4764,N_1087);
and U6488 (N_6488,N_848,N_2128);
xor U6489 (N_6489,N_4730,N_526);
or U6490 (N_6490,N_4598,N_2890);
xnor U6491 (N_6491,N_3772,N_3630);
and U6492 (N_6492,N_2200,N_3050);
and U6493 (N_6493,N_896,N_3832);
nand U6494 (N_6494,N_4116,N_953);
xnor U6495 (N_6495,N_2884,N_3370);
nand U6496 (N_6496,N_1382,N_2550);
and U6497 (N_6497,N_2404,N_3163);
nand U6498 (N_6498,N_4133,N_3436);
and U6499 (N_6499,N_248,N_1497);
and U6500 (N_6500,N_2252,N_837);
or U6501 (N_6501,N_229,N_2203);
xor U6502 (N_6502,N_1781,N_1673);
xnor U6503 (N_6503,N_3575,N_4732);
nand U6504 (N_6504,N_784,N_4468);
nor U6505 (N_6505,N_601,N_1233);
nand U6506 (N_6506,N_1876,N_1655);
nor U6507 (N_6507,N_2624,N_3616);
nand U6508 (N_6508,N_4085,N_422);
nor U6509 (N_6509,N_2732,N_1039);
or U6510 (N_6510,N_1759,N_4753);
or U6511 (N_6511,N_700,N_2702);
or U6512 (N_6512,N_3638,N_2661);
and U6513 (N_6513,N_4314,N_352);
nand U6514 (N_6514,N_4463,N_2755);
nor U6515 (N_6515,N_1776,N_4993);
or U6516 (N_6516,N_4106,N_3270);
nor U6517 (N_6517,N_4152,N_3673);
nor U6518 (N_6518,N_364,N_277);
nand U6519 (N_6519,N_2412,N_1256);
nor U6520 (N_6520,N_1519,N_905);
and U6521 (N_6521,N_4985,N_3118);
nor U6522 (N_6522,N_3384,N_1762);
xnor U6523 (N_6523,N_2023,N_2311);
or U6524 (N_6524,N_4061,N_752);
or U6525 (N_6525,N_743,N_1429);
nor U6526 (N_6526,N_2050,N_1954);
xor U6527 (N_6527,N_2010,N_3480);
or U6528 (N_6528,N_4184,N_51);
nand U6529 (N_6529,N_387,N_3846);
xnor U6530 (N_6530,N_1041,N_2784);
nor U6531 (N_6531,N_4831,N_1541);
nor U6532 (N_6532,N_3345,N_3794);
nor U6533 (N_6533,N_3473,N_2455);
nand U6534 (N_6534,N_934,N_1632);
and U6535 (N_6535,N_3312,N_954);
and U6536 (N_6536,N_3003,N_1662);
or U6537 (N_6537,N_1144,N_4613);
and U6538 (N_6538,N_3506,N_3802);
xor U6539 (N_6539,N_2102,N_1270);
and U6540 (N_6540,N_1853,N_2896);
and U6541 (N_6541,N_2882,N_404);
nand U6542 (N_6542,N_209,N_4708);
xnor U6543 (N_6543,N_2099,N_664);
xnor U6544 (N_6544,N_3405,N_458);
and U6545 (N_6545,N_3984,N_1803);
nand U6546 (N_6546,N_239,N_1215);
xor U6547 (N_6547,N_445,N_2009);
and U6548 (N_6548,N_2262,N_2529);
xnor U6549 (N_6549,N_243,N_1552);
or U6550 (N_6550,N_2309,N_3805);
and U6551 (N_6551,N_4331,N_4369);
and U6552 (N_6552,N_4324,N_4301);
xnor U6553 (N_6553,N_1375,N_2933);
nor U6554 (N_6554,N_3488,N_2724);
nand U6555 (N_6555,N_3599,N_4264);
and U6556 (N_6556,N_2945,N_278);
nand U6557 (N_6557,N_3515,N_2378);
xor U6558 (N_6558,N_4267,N_4556);
nor U6559 (N_6559,N_1935,N_4772);
or U6560 (N_6560,N_4495,N_1737);
or U6561 (N_6561,N_309,N_1844);
xor U6562 (N_6562,N_424,N_3021);
or U6563 (N_6563,N_3881,N_832);
or U6564 (N_6564,N_465,N_4631);
nor U6565 (N_6565,N_3013,N_2396);
nor U6566 (N_6566,N_262,N_4628);
nor U6567 (N_6567,N_4830,N_1259);
xnor U6568 (N_6568,N_2071,N_597);
nor U6569 (N_6569,N_4021,N_4402);
nand U6570 (N_6570,N_2482,N_3322);
or U6571 (N_6571,N_1575,N_594);
nand U6572 (N_6572,N_4080,N_307);
xor U6573 (N_6573,N_1615,N_4044);
nor U6574 (N_6574,N_3964,N_2163);
or U6575 (N_6575,N_2107,N_4742);
nand U6576 (N_6576,N_1454,N_2573);
xor U6577 (N_6577,N_188,N_87);
or U6578 (N_6578,N_1237,N_3407);
nor U6579 (N_6579,N_4600,N_439);
and U6580 (N_6580,N_1962,N_4341);
nor U6581 (N_6581,N_1576,N_258);
nand U6582 (N_6582,N_4041,N_4950);
nand U6583 (N_6583,N_1012,N_4291);
xnor U6584 (N_6584,N_3570,N_3529);
nor U6585 (N_6585,N_3975,N_926);
nand U6586 (N_6586,N_3884,N_311);
and U6587 (N_6587,N_464,N_4429);
xor U6588 (N_6588,N_2271,N_4209);
and U6589 (N_6589,N_1493,N_1631);
nor U6590 (N_6590,N_938,N_4384);
and U6591 (N_6591,N_1633,N_4516);
nand U6592 (N_6592,N_1800,N_4121);
and U6593 (N_6593,N_3316,N_4465);
xor U6594 (N_6594,N_1437,N_377);
and U6595 (N_6595,N_4853,N_2873);
or U6596 (N_6596,N_1343,N_4666);
nand U6597 (N_6597,N_1460,N_1082);
or U6598 (N_6598,N_1252,N_4808);
and U6599 (N_6599,N_1612,N_2722);
nor U6600 (N_6600,N_2809,N_3143);
or U6601 (N_6601,N_3923,N_4228);
or U6602 (N_6602,N_4039,N_4651);
and U6603 (N_6603,N_800,N_1924);
or U6604 (N_6604,N_3094,N_790);
xor U6605 (N_6605,N_759,N_1892);
xor U6606 (N_6606,N_3303,N_3740);
and U6607 (N_6607,N_80,N_3933);
xor U6608 (N_6608,N_3806,N_4948);
xor U6609 (N_6609,N_2243,N_1824);
xnor U6610 (N_6610,N_396,N_620);
xor U6611 (N_6611,N_826,N_4769);
nor U6612 (N_6612,N_2166,N_2876);
or U6613 (N_6613,N_3819,N_1601);
or U6614 (N_6614,N_561,N_1840);
and U6615 (N_6615,N_293,N_3380);
or U6616 (N_6616,N_4466,N_4273);
xor U6617 (N_6617,N_3667,N_2306);
nor U6618 (N_6618,N_1320,N_672);
and U6619 (N_6619,N_558,N_3358);
xnor U6620 (N_6620,N_214,N_982);
or U6621 (N_6621,N_2561,N_1236);
and U6622 (N_6622,N_1787,N_3269);
nor U6623 (N_6623,N_943,N_2031);
xnor U6624 (N_6624,N_3339,N_4430);
nand U6625 (N_6625,N_1888,N_3058);
or U6626 (N_6626,N_3165,N_2480);
and U6627 (N_6627,N_3336,N_3906);
xor U6628 (N_6628,N_2813,N_1872);
or U6629 (N_6629,N_221,N_1771);
nor U6630 (N_6630,N_1298,N_444);
xor U6631 (N_6631,N_4882,N_386);
or U6632 (N_6632,N_4572,N_3388);
nor U6633 (N_6633,N_2492,N_3809);
nor U6634 (N_6634,N_4111,N_748);
nor U6635 (N_6635,N_4781,N_4694);
or U6636 (N_6636,N_1775,N_4174);
nor U6637 (N_6637,N_3674,N_3106);
and U6638 (N_6638,N_3059,N_250);
xor U6639 (N_6639,N_2844,N_3581);
nor U6640 (N_6640,N_3870,N_1127);
nand U6641 (N_6641,N_3650,N_3554);
nor U6642 (N_6642,N_2407,N_3547);
xor U6643 (N_6643,N_1500,N_3280);
xnor U6644 (N_6644,N_1891,N_3305);
xor U6645 (N_6645,N_1849,N_3008);
xor U6646 (N_6646,N_2006,N_1712);
nor U6647 (N_6647,N_505,N_3612);
xor U6648 (N_6648,N_3315,N_3125);
or U6649 (N_6649,N_2626,N_4940);
nor U6650 (N_6650,N_4801,N_4139);
nand U6651 (N_6651,N_4725,N_4741);
nor U6652 (N_6652,N_255,N_1275);
nand U6653 (N_6653,N_612,N_66);
or U6654 (N_6654,N_1583,N_86);
or U6655 (N_6655,N_1841,N_4293);
and U6656 (N_6656,N_2042,N_3985);
nor U6657 (N_6657,N_744,N_2862);
or U6658 (N_6658,N_4854,N_1996);
xnor U6659 (N_6659,N_3553,N_4920);
nand U6660 (N_6660,N_203,N_4714);
nor U6661 (N_6661,N_1480,N_305);
nand U6662 (N_6662,N_2345,N_1340);
nor U6663 (N_6663,N_2938,N_846);
and U6664 (N_6664,N_4891,N_1249);
or U6665 (N_6665,N_580,N_3779);
and U6666 (N_6666,N_1804,N_2343);
nand U6667 (N_6667,N_2834,N_869);
xor U6668 (N_6668,N_1030,N_1661);
and U6669 (N_6669,N_1417,N_3204);
or U6670 (N_6670,N_2100,N_4964);
nor U6671 (N_6671,N_1751,N_3321);
nand U6672 (N_6672,N_2231,N_4533);
nand U6673 (N_6673,N_625,N_1953);
or U6674 (N_6674,N_3716,N_253);
xnor U6675 (N_6675,N_109,N_3978);
and U6676 (N_6676,N_2014,N_1358);
and U6677 (N_6677,N_1738,N_1896);
xor U6678 (N_6678,N_2718,N_1276);
nor U6679 (N_6679,N_78,N_2409);
nand U6680 (N_6680,N_2685,N_4348);
nor U6681 (N_6681,N_2842,N_3501);
or U6682 (N_6682,N_2914,N_1923);
and U6683 (N_6683,N_3311,N_412);
nand U6684 (N_6684,N_1866,N_2782);
nor U6685 (N_6685,N_780,N_4224);
or U6686 (N_6686,N_410,N_4745);
nand U6687 (N_6687,N_242,N_1194);
or U6688 (N_6688,N_3041,N_2069);
or U6689 (N_6689,N_120,N_3344);
nor U6690 (N_6690,N_2145,N_72);
nor U6691 (N_6691,N_794,N_4596);
and U6692 (N_6692,N_3298,N_1560);
and U6693 (N_6693,N_1796,N_1425);
nor U6694 (N_6694,N_3331,N_2375);
xor U6695 (N_6695,N_4026,N_3012);
and U6696 (N_6696,N_3775,N_1354);
and U6697 (N_6697,N_3635,N_4539);
or U6698 (N_6698,N_279,N_1501);
xnor U6699 (N_6699,N_2366,N_2759);
xor U6700 (N_6700,N_1265,N_950);
xor U6701 (N_6701,N_4894,N_4432);
xnor U6702 (N_6702,N_4756,N_1975);
and U6703 (N_6703,N_4455,N_3139);
xor U6704 (N_6704,N_3302,N_339);
nor U6705 (N_6705,N_2284,N_543);
and U6706 (N_6706,N_1829,N_2035);
nor U6707 (N_6707,N_2707,N_4661);
nand U6708 (N_6708,N_2894,N_681);
nand U6709 (N_6709,N_2800,N_1408);
nor U6710 (N_6710,N_2698,N_669);
nand U6711 (N_6711,N_2427,N_2772);
or U6712 (N_6712,N_4508,N_1980);
and U6713 (N_6713,N_4629,N_264);
xor U6714 (N_6714,N_3467,N_117);
and U6715 (N_6715,N_2044,N_649);
nor U6716 (N_6716,N_2704,N_4299);
or U6717 (N_6717,N_4050,N_2502);
and U6718 (N_6718,N_434,N_2017);
xor U6719 (N_6719,N_4524,N_626);
xor U6720 (N_6720,N_2670,N_789);
nor U6721 (N_6721,N_2386,N_1381);
or U6722 (N_6722,N_2606,N_2523);
nand U6723 (N_6723,N_1678,N_2000);
xnor U6724 (N_6724,N_4411,N_2804);
nor U6725 (N_6725,N_3062,N_1925);
or U6726 (N_6726,N_319,N_183);
nand U6727 (N_6727,N_84,N_1226);
xor U6728 (N_6728,N_4386,N_2628);
and U6729 (N_6729,N_2735,N_2429);
nor U6730 (N_6730,N_158,N_2581);
and U6731 (N_6731,N_1843,N_2332);
nor U6732 (N_6732,N_421,N_2898);
xor U6733 (N_6733,N_4229,N_3433);
nor U6734 (N_6734,N_21,N_3781);
nand U6735 (N_6735,N_841,N_4888);
and U6736 (N_6736,N_1785,N_2440);
or U6737 (N_6737,N_4147,N_2627);
xnor U6738 (N_6738,N_2763,N_2700);
xnor U6739 (N_6739,N_2927,N_3683);
nand U6740 (N_6740,N_2817,N_3812);
nor U6741 (N_6741,N_1573,N_2644);
nor U6742 (N_6742,N_3818,N_2079);
xor U6743 (N_6743,N_99,N_430);
xnor U6744 (N_6744,N_1364,N_129);
or U6745 (N_6745,N_2871,N_929);
xor U6746 (N_6746,N_2490,N_2075);
nor U6747 (N_6747,N_890,N_4770);
xnor U6748 (N_6748,N_4658,N_1305);
and U6749 (N_6749,N_3274,N_951);
nor U6750 (N_6750,N_201,N_4699);
and U6751 (N_6751,N_3602,N_3415);
nor U6752 (N_6752,N_1262,N_879);
nand U6753 (N_6753,N_2611,N_4295);
xnor U6754 (N_6754,N_4373,N_2957);
and U6755 (N_6755,N_1609,N_3724);
xor U6756 (N_6756,N_1670,N_3156);
or U6757 (N_6757,N_552,N_507);
nor U6758 (N_6758,N_1820,N_4933);
and U6759 (N_6759,N_4417,N_1599);
nor U6760 (N_6760,N_2159,N_4606);
nor U6761 (N_6761,N_4444,N_1689);
nand U6762 (N_6762,N_3823,N_4360);
nor U6763 (N_6763,N_822,N_2356);
and U6764 (N_6764,N_4459,N_659);
and U6765 (N_6765,N_3719,N_351);
nor U6766 (N_6766,N_2247,N_682);
or U6767 (N_6767,N_4663,N_3901);
or U6768 (N_6768,N_3483,N_4866);
nor U6769 (N_6769,N_1446,N_85);
xnor U6770 (N_6770,N_1581,N_3357);
xor U6771 (N_6771,N_3689,N_2170);
nor U6772 (N_6772,N_3258,N_2209);
xor U6773 (N_6773,N_1556,N_508);
nand U6774 (N_6774,N_4880,N_2923);
nor U6775 (N_6775,N_493,N_3963);
nand U6776 (N_6776,N_2331,N_4346);
nor U6777 (N_6777,N_1434,N_2140);
and U6778 (N_6778,N_560,N_831);
nor U6779 (N_6779,N_1200,N_3887);
nand U6780 (N_6780,N_233,N_4837);
or U6781 (N_6781,N_166,N_3117);
and U6782 (N_6782,N_1593,N_3678);
nand U6783 (N_6783,N_981,N_1625);
or U6784 (N_6784,N_3725,N_920);
xnor U6785 (N_6785,N_4248,N_3869);
nand U6786 (N_6786,N_3950,N_263);
or U6787 (N_6787,N_2242,N_4871);
nor U6788 (N_6788,N_2613,N_4279);
nor U6789 (N_6789,N_4494,N_1178);
xor U6790 (N_6790,N_1413,N_541);
or U6791 (N_6791,N_4127,N_2937);
nor U6792 (N_6792,N_3288,N_975);
and U6793 (N_6793,N_835,N_1951);
or U6794 (N_6794,N_448,N_380);
or U6795 (N_6795,N_3278,N_0);
xor U6796 (N_6796,N_2219,N_1286);
or U6797 (N_6797,N_2794,N_4427);
xor U6798 (N_6798,N_1415,N_213);
xor U6799 (N_6799,N_1496,N_3039);
xor U6800 (N_6800,N_4750,N_295);
nand U6801 (N_6801,N_4347,N_4258);
nor U6802 (N_6802,N_3006,N_2675);
xnor U6803 (N_6803,N_450,N_4236);
or U6804 (N_6804,N_419,N_715);
nand U6805 (N_6805,N_4983,N_1273);
or U6806 (N_6806,N_4605,N_4298);
nand U6807 (N_6807,N_59,N_3874);
or U6808 (N_6808,N_3248,N_1185);
or U6809 (N_6809,N_1266,N_2508);
and U6810 (N_6810,N_4650,N_4682);
and U6811 (N_6811,N_4089,N_2845);
nand U6812 (N_6812,N_2887,N_1169);
xor U6813 (N_6813,N_1667,N_4237);
nor U6814 (N_6814,N_604,N_3538);
or U6815 (N_6815,N_4727,N_460);
xor U6816 (N_6816,N_782,N_275);
nand U6817 (N_6817,N_2213,N_966);
nand U6818 (N_6818,N_994,N_1199);
or U6819 (N_6819,N_4925,N_2841);
nand U6820 (N_6820,N_2623,N_4409);
nand U6821 (N_6821,N_282,N_4608);
or U6822 (N_6822,N_3970,N_1770);
nand U6823 (N_6823,N_562,N_4895);
xnor U6824 (N_6824,N_2511,N_1360);
or U6825 (N_6825,N_4568,N_786);
nor U6826 (N_6826,N_1922,N_4640);
xor U6827 (N_6827,N_2028,N_891);
nand U6828 (N_6828,N_4786,N_3609);
and U6829 (N_6829,N_3969,N_2664);
or U6830 (N_6830,N_3684,N_3987);
nor U6831 (N_6831,N_1046,N_3879);
or U6832 (N_6832,N_1075,N_154);
nor U6833 (N_6833,N_467,N_4636);
nand U6834 (N_6834,N_1292,N_1003);
nand U6835 (N_6835,N_3998,N_2142);
nor U6836 (N_6836,N_4071,N_568);
nor U6837 (N_6837,N_3029,N_1166);
nand U6838 (N_6838,N_1057,N_368);
or U6839 (N_6839,N_2835,N_1988);
and U6840 (N_6840,N_960,N_1198);
or U6841 (N_6841,N_4185,N_33);
xor U6842 (N_6842,N_1802,N_3491);
nor U6843 (N_6843,N_852,N_4144);
and U6844 (N_6844,N_1966,N_1608);
nand U6845 (N_6845,N_2958,N_2996);
or U6846 (N_6846,N_4783,N_3366);
and U6847 (N_6847,N_4759,N_593);
and U6848 (N_6848,N_2846,N_1826);
nor U6849 (N_6849,N_854,N_2827);
nor U6850 (N_6850,N_4330,N_3653);
or U6851 (N_6851,N_4383,N_4109);
or U6852 (N_6852,N_2789,N_4951);
xnor U6853 (N_6853,N_1363,N_729);
and U6854 (N_6854,N_1369,N_522);
nand U6855 (N_6855,N_4967,N_3584);
and U6856 (N_6856,N_25,N_3814);
and U6857 (N_6857,N_1311,N_429);
nand U6858 (N_6858,N_3527,N_1083);
and U6859 (N_6859,N_2533,N_1772);
nor U6860 (N_6860,N_2517,N_4054);
or U6861 (N_6861,N_3092,N_2665);
nand U6862 (N_6862,N_2690,N_2049);
nor U6863 (N_6863,N_1383,N_1533);
or U6864 (N_6864,N_1814,N_1258);
nand U6865 (N_6865,N_3124,N_4852);
nand U6866 (N_6866,N_1289,N_3052);
nand U6867 (N_6867,N_438,N_1958);
xor U6868 (N_6868,N_2881,N_327);
xnor U6869 (N_6869,N_186,N_1216);
and U6870 (N_6870,N_2920,N_4457);
or U6871 (N_6871,N_4257,N_4773);
nand U6872 (N_6872,N_4296,N_1949);
xnor U6873 (N_6873,N_1871,N_3174);
and U6874 (N_6874,N_2918,N_4367);
or U6875 (N_6875,N_3607,N_2916);
nor U6876 (N_6876,N_651,N_4570);
or U6877 (N_6877,N_2499,N_4979);
nand U6878 (N_6878,N_2173,N_4132);
and U6879 (N_6879,N_1263,N_4136);
and U6880 (N_6880,N_3645,N_2557);
nand U6881 (N_6881,N_155,N_2610);
or U6882 (N_6882,N_4105,N_2779);
and U6883 (N_6883,N_76,N_1184);
nor U6884 (N_6884,N_525,N_2255);
nand U6885 (N_6885,N_2632,N_3100);
xor U6886 (N_6886,N_897,N_4280);
xor U6887 (N_6887,N_1137,N_1431);
xnor U6888 (N_6888,N_1764,N_3452);
xor U6889 (N_6889,N_4303,N_1267);
xor U6890 (N_6890,N_3171,N_2432);
or U6891 (N_6891,N_1395,N_2314);
xor U6892 (N_6892,N_4395,N_2245);
xor U6893 (N_6893,N_2045,N_2232);
nor U6894 (N_6894,N_3820,N_3637);
and U6895 (N_6895,N_1001,N_4434);
nor U6896 (N_6896,N_1109,N_4469);
and U6897 (N_6897,N_1389,N_270);
nor U6898 (N_6898,N_4126,N_4677);
nor U6899 (N_6899,N_2506,N_3941);
nand U6900 (N_6900,N_3462,N_1456);
nand U6901 (N_6901,N_4607,N_523);
xor U6902 (N_6902,N_710,N_1869);
xnor U6903 (N_6903,N_1725,N_606);
xnor U6904 (N_6904,N_175,N_2124);
nand U6905 (N_6905,N_2215,N_4029);
nor U6906 (N_6906,N_3558,N_4063);
xor U6907 (N_6907,N_4740,N_2143);
nor U6908 (N_6908,N_1439,N_3157);
xnor U6909 (N_6909,N_4747,N_3770);
and U6910 (N_6910,N_722,N_4574);
and U6911 (N_6911,N_4025,N_4004);
nand U6912 (N_6912,N_3679,N_4120);
nor U6913 (N_6913,N_3084,N_1909);
or U6914 (N_6914,N_1538,N_3696);
nand U6915 (N_6915,N_2198,N_719);
xor U6916 (N_6916,N_1242,N_1016);
xor U6917 (N_6917,N_4553,N_3811);
or U6918 (N_6918,N_1974,N_827);
and U6919 (N_6919,N_2637,N_123);
xnor U6920 (N_6920,N_959,N_1862);
nor U6921 (N_6921,N_2850,N_1021);
and U6922 (N_6922,N_2863,N_1850);
nand U6923 (N_6923,N_821,N_4537);
xor U6924 (N_6924,N_2024,N_4603);
xor U6925 (N_6925,N_3569,N_15);
xor U6926 (N_6926,N_4122,N_1875);
xor U6927 (N_6927,N_1642,N_1950);
nand U6928 (N_6928,N_4272,N_3411);
or U6929 (N_6929,N_1969,N_4671);
or U6930 (N_6930,N_1763,N_2441);
nor U6931 (N_6931,N_2893,N_4522);
or U6932 (N_6932,N_3589,N_3912);
and U6933 (N_6933,N_2537,N_3147);
or U6934 (N_6934,N_1101,N_4487);
nor U6935 (N_6935,N_3095,N_4672);
nor U6936 (N_6936,N_38,N_1621);
xnor U6937 (N_6937,N_382,N_468);
or U6938 (N_6938,N_3421,N_1462);
or U6939 (N_6939,N_647,N_740);
nor U6940 (N_6940,N_77,N_3324);
nand U6941 (N_6941,N_372,N_4856);
and U6942 (N_6942,N_29,N_4194);
or U6943 (N_6943,N_1246,N_2122);
nor U6944 (N_6944,N_592,N_1812);
nand U6945 (N_6945,N_1634,N_2764);
and U6946 (N_6946,N_1084,N_4550);
nand U6947 (N_6947,N_755,N_4576);
nor U6948 (N_6948,N_2740,N_836);
or U6949 (N_6949,N_4798,N_1160);
xor U6950 (N_6950,N_4675,N_1855);
nand U6951 (N_6951,N_2228,N_1929);
nand U6952 (N_6952,N_2447,N_3700);
and U6953 (N_6953,N_4437,N_1339);
or U6954 (N_6954,N_3487,N_791);
nand U6955 (N_6955,N_4911,N_4577);
nor U6956 (N_6956,N_2961,N_3040);
xor U6957 (N_6957,N_4612,N_3661);
xor U6958 (N_6958,N_2413,N_2125);
nor U6959 (N_6959,N_4847,N_4289);
xor U6960 (N_6960,N_1470,N_3939);
and U6961 (N_6961,N_3561,N_2046);
and U6962 (N_6962,N_2132,N_3293);
nor U6963 (N_6963,N_665,N_374);
or U6964 (N_6964,N_2258,N_199);
or U6965 (N_6965,N_1919,N_1313);
or U6966 (N_6966,N_1714,N_4214);
nand U6967 (N_6967,N_1362,N_4480);
or U6968 (N_6968,N_469,N_2858);
and U6969 (N_6969,N_4102,N_773);
nand U6970 (N_6970,N_4143,N_3913);
xor U6971 (N_6971,N_4947,N_3917);
nor U6972 (N_6972,N_1411,N_152);
and U6973 (N_6973,N_986,N_1654);
and U6974 (N_6974,N_4505,N_4379);
xnor U6975 (N_6975,N_3025,N_4218);
and U6976 (N_6976,N_2304,N_1797);
nor U6977 (N_6977,N_4806,N_4780);
or U6978 (N_6978,N_1692,N_1586);
nor U6979 (N_6979,N_1334,N_2086);
nand U6980 (N_6980,N_49,N_2553);
or U6981 (N_6981,N_2910,N_1761);
or U6982 (N_6982,N_4551,N_1332);
and U6983 (N_6983,N_3090,N_2158);
xnor U6984 (N_6984,N_1032,N_1396);
and U6985 (N_6985,N_4941,N_1118);
xnor U6986 (N_6986,N_2536,N_4243);
xnor U6987 (N_6987,N_2748,N_4410);
or U6988 (N_6988,N_4442,N_3835);
nor U6989 (N_6989,N_519,N_1349);
nor U6990 (N_6990,N_2138,N_2369);
or U6991 (N_6991,N_4822,N_3960);
nor U6992 (N_6992,N_2183,N_4083);
xor U6993 (N_6993,N_530,N_3481);
nand U6994 (N_6994,N_4885,N_4502);
or U6995 (N_6995,N_912,N_4509);
nand U6996 (N_6996,N_4887,N_1044);
and U6997 (N_6997,N_3761,N_3731);
nand U6998 (N_6998,N_4148,N_2295);
or U6999 (N_6999,N_1941,N_184);
or U7000 (N_7000,N_3228,N_2216);
nor U7001 (N_7001,N_4146,N_691);
or U7002 (N_7002,N_4278,N_346);
and U7003 (N_7003,N_4820,N_7);
and U7004 (N_7004,N_1857,N_3099);
xnor U7005 (N_7005,N_191,N_2824);
and U7006 (N_7006,N_3702,N_144);
and U7007 (N_7007,N_4549,N_717);
or U7008 (N_7008,N_4040,N_3525);
and U7009 (N_7009,N_575,N_3465);
and U7010 (N_7010,N_2547,N_3748);
nand U7011 (N_7011,N_2791,N_2921);
or U7012 (N_7012,N_3922,N_4507);
and U7013 (N_7013,N_4070,N_716);
xnor U7014 (N_7014,N_900,N_4250);
nand U7015 (N_7015,N_3440,N_4349);
and U7016 (N_7016,N_1834,N_2659);
and U7017 (N_7017,N_4615,N_4910);
or U7018 (N_7018,N_1264,N_3845);
nor U7019 (N_7019,N_2150,N_527);
nand U7020 (N_7020,N_2878,N_2337);
nor U7021 (N_7021,N_2519,N_251);
nor U7022 (N_7022,N_2334,N_318);
nor U7023 (N_7023,N_4312,N_1525);
nand U7024 (N_7024,N_3414,N_1898);
nor U7025 (N_7025,N_3116,N_376);
or U7026 (N_7026,N_3892,N_1611);
or U7027 (N_7027,N_4490,N_4478);
nor U7028 (N_7028,N_1387,N_3002);
nor U7029 (N_7029,N_2199,N_1090);
xnor U7030 (N_7030,N_4201,N_378);
nor U7031 (N_7031,N_3771,N_3534);
and U7032 (N_7032,N_333,N_4338);
or U7033 (N_7033,N_1034,N_2812);
nand U7034 (N_7034,N_2741,N_3611);
nand U7035 (N_7035,N_2543,N_3618);
xnor U7036 (N_7036,N_2830,N_845);
nand U7037 (N_7037,N_1441,N_1356);
nor U7038 (N_7038,N_2522,N_2354);
and U7039 (N_7039,N_3571,N_3624);
or U7040 (N_7040,N_1272,N_4020);
xor U7041 (N_7041,N_1433,N_1230);
nand U7042 (N_7042,N_605,N_4693);
xnor U7043 (N_7043,N_1342,N_3710);
nand U7044 (N_7044,N_2672,N_1155);
nand U7045 (N_7045,N_952,N_3113);
and U7046 (N_7046,N_1451,N_389);
nand U7047 (N_7047,N_4526,N_1481);
and U7048 (N_7048,N_1861,N_2261);
nor U7049 (N_7049,N_652,N_2643);
nor U7050 (N_7050,N_3427,N_3644);
and U7051 (N_7051,N_545,N_208);
nand U7052 (N_7052,N_3406,N_1910);
or U7053 (N_7053,N_2498,N_3418);
and U7054 (N_7054,N_3261,N_2139);
or U7055 (N_7055,N_2344,N_2156);
nor U7056 (N_7056,N_1508,N_4641);
or U7057 (N_7057,N_4618,N_503);
xnor U7058 (N_7058,N_4707,N_1961);
or U7059 (N_7059,N_1865,N_3043);
and U7060 (N_7060,N_610,N_515);
xor U7061 (N_7061,N_1813,N_1227);
nand U7062 (N_7062,N_2692,N_171);
xor U7063 (N_7063,N_1965,N_433);
nand U7064 (N_7064,N_3867,N_965);
or U7065 (N_7065,N_3290,N_1886);
nand U7066 (N_7066,N_3420,N_2380);
nor U7067 (N_7067,N_358,N_2998);
nand U7068 (N_7068,N_1426,N_1564);
xnor U7069 (N_7069,N_4715,N_3150);
and U7070 (N_7070,N_3574,N_489);
nor U7071 (N_7071,N_2888,N_3944);
xnor U7072 (N_7072,N_2587,N_1873);
xnor U7073 (N_7073,N_813,N_3230);
or U7074 (N_7074,N_3615,N_880);
nand U7075 (N_7075,N_2967,N_2037);
nand U7076 (N_7076,N_3327,N_1076);
nand U7077 (N_7077,N_3730,N_3961);
and U7078 (N_7078,N_3132,N_904);
or U7079 (N_7079,N_3064,N_2188);
and U7080 (N_7080,N_658,N_667);
nand U7081 (N_7081,N_1370,N_1822);
or U7082 (N_7082,N_1296,N_1578);
or U7083 (N_7083,N_3800,N_2689);
nor U7084 (N_7084,N_799,N_4474);
nor U7085 (N_7085,N_3237,N_512);
or U7086 (N_7086,N_3028,N_1542);
nor U7087 (N_7087,N_1335,N_3352);
or U7088 (N_7088,N_1,N_2104);
nor U7089 (N_7089,N_3067,N_1729);
and U7090 (N_7090,N_576,N_2802);
xnor U7091 (N_7091,N_3687,N_1485);
and U7092 (N_7092,N_4581,N_2969);
or U7093 (N_7093,N_432,N_2934);
nand U7094 (N_7094,N_3195,N_2847);
xor U7095 (N_7095,N_2977,N_1132);
nor U7096 (N_7096,N_3544,N_2683);
nand U7097 (N_7097,N_694,N_477);
nor U7098 (N_7098,N_1627,N_2954);
and U7099 (N_7099,N_2263,N_2655);
xnor U7100 (N_7100,N_1675,N_3011);
nor U7101 (N_7101,N_2151,N_3149);
and U7102 (N_7102,N_2752,N_1808);
and U7103 (N_7103,N_703,N_3085);
xor U7104 (N_7104,N_3785,N_2697);
nor U7105 (N_7105,N_4203,N_3557);
nand U7106 (N_7106,N_88,N_1704);
and U7107 (N_7107,N_3416,N_2686);
nor U7108 (N_7108,N_978,N_2991);
and U7109 (N_7109,N_2056,N_60);
or U7110 (N_7110,N_2298,N_147);
xor U7111 (N_7111,N_289,N_1402);
and U7112 (N_7112,N_3413,N_1131);
or U7113 (N_7113,N_3540,N_1811);
or U7114 (N_7114,N_1479,N_462);
nand U7115 (N_7115,N_949,N_2338);
nand U7116 (N_7116,N_4319,N_2333);
xnor U7117 (N_7117,N_1600,N_384);
nand U7118 (N_7118,N_75,N_4807);
xnor U7119 (N_7119,N_914,N_4531);
xor U7120 (N_7120,N_114,N_1696);
nand U7121 (N_7121,N_4038,N_1607);
nand U7122 (N_7122,N_3032,N_4304);
or U7123 (N_7123,N_4902,N_3299);
or U7124 (N_7124,N_3155,N_1978);
nor U7125 (N_7125,N_2291,N_3138);
nor U7126 (N_7126,N_4922,N_4890);
nor U7127 (N_7127,N_3347,N_4206);
or U7128 (N_7128,N_2403,N_1623);
xnor U7129 (N_7129,N_4456,N_2471);
or U7130 (N_7130,N_4805,N_2641);
xor U7131 (N_7131,N_2157,N_1113);
xor U7132 (N_7132,N_4101,N_57);
nor U7133 (N_7133,N_3362,N_1838);
nor U7134 (N_7134,N_3991,N_4140);
xnor U7135 (N_7135,N_3271,N_4355);
nor U7136 (N_7136,N_3192,N_3546);
xor U7137 (N_7137,N_3353,N_2754);
nor U7138 (N_7138,N_3210,N_4996);
and U7139 (N_7139,N_306,N_4904);
nor U7140 (N_7140,N_2218,N_1992);
and U7141 (N_7141,N_4187,N_1149);
xnor U7142 (N_7142,N_1374,N_510);
and U7143 (N_7143,N_2872,N_256);
nor U7144 (N_7144,N_4378,N_1102);
nor U7145 (N_7145,N_2385,N_4833);
nand U7146 (N_7146,N_1630,N_4407);
or U7147 (N_7147,N_2466,N_3713);
xor U7148 (N_7148,N_2089,N_2786);
and U7149 (N_7149,N_588,N_1828);
nor U7150 (N_7150,N_1416,N_3492);
nor U7151 (N_7151,N_4117,N_4215);
and U7152 (N_7152,N_4428,N_1423);
nand U7153 (N_7153,N_535,N_4368);
xor U7154 (N_7154,N_4023,N_3493);
nor U7155 (N_7155,N_2638,N_4238);
nand U7156 (N_7156,N_2251,N_1926);
xnor U7157 (N_7157,N_569,N_1790);
xnor U7158 (N_7158,N_4932,N_1647);
nor U7159 (N_7159,N_2040,N_1104);
and U7160 (N_7160,N_442,N_4990);
and U7161 (N_7161,N_4957,N_935);
or U7162 (N_7162,N_2615,N_2905);
and U7163 (N_7163,N_1756,N_689);
nor U7164 (N_7164,N_4784,N_3660);
xor U7165 (N_7165,N_3983,N_955);
nand U7166 (N_7166,N_3815,N_3801);
and U7167 (N_7167,N_4055,N_2249);
nand U7168 (N_7168,N_3821,N_4058);
or U7169 (N_7169,N_1982,N_3919);
nor U7170 (N_7170,N_3972,N_819);
nand U7171 (N_7171,N_1571,N_47);
xor U7172 (N_7172,N_2956,N_1065);
or U7173 (N_7173,N_2585,N_238);
nand U7174 (N_7174,N_291,N_3166);
nand U7175 (N_7175,N_1846,N_3921);
and U7176 (N_7176,N_654,N_296);
and U7177 (N_7177,N_1720,N_4036);
or U7178 (N_7178,N_2999,N_340);
nand U7179 (N_7179,N_3522,N_4802);
nand U7180 (N_7180,N_2699,N_1619);
nor U7181 (N_7181,N_1643,N_1106);
or U7182 (N_7182,N_3112,N_3839);
nand U7183 (N_7183,N_3707,N_3810);
or U7184 (N_7184,N_3088,N_234);
and U7185 (N_7185,N_1288,N_500);
nor U7186 (N_7186,N_2790,N_1768);
and U7187 (N_7187,N_2743,N_1597);
xor U7188 (N_7188,N_871,N_962);
nor U7189 (N_7189,N_4938,N_4356);
or U7190 (N_7190,N_2308,N_1837);
nor U7191 (N_7191,N_3078,N_189);
nor U7192 (N_7192,N_3591,N_1716);
xor U7193 (N_7193,N_4874,N_1687);
nand U7194 (N_7194,N_4915,N_1399);
and U7195 (N_7195,N_2007,N_690);
nand U7196 (N_7196,N_3206,N_2895);
nor U7197 (N_7197,N_1326,N_1817);
nor U7198 (N_7198,N_3742,N_1550);
nand U7199 (N_7199,N_440,N_706);
or U7200 (N_7200,N_3096,N_1361);
nand U7201 (N_7201,N_198,N_4062);
xor U7202 (N_7202,N_329,N_1367);
xor U7203 (N_7203,N_3629,N_2971);
and U7204 (N_7204,N_2618,N_2564);
xnor U7205 (N_7205,N_4530,N_2719);
or U7206 (N_7206,N_1832,N_1271);
or U7207 (N_7207,N_4790,N_2951);
or U7208 (N_7208,N_3907,N_3535);
nor U7209 (N_7209,N_4746,N_2229);
nand U7210 (N_7210,N_1806,N_2691);
or U7211 (N_7211,N_375,N_2359);
xor U7212 (N_7212,N_974,N_1639);
and U7213 (N_7213,N_2891,N_1119);
nand U7214 (N_7214,N_528,N_31);
and U7215 (N_7215,N_2995,N_735);
and U7216 (N_7216,N_4791,N_4381);
or U7217 (N_7217,N_2833,N_2569);
and U7218 (N_7218,N_3521,N_202);
nand U7219 (N_7219,N_4339,N_4810);
nor U7220 (N_7220,N_1794,N_1366);
nand U7221 (N_7221,N_4850,N_1228);
xnor U7222 (N_7222,N_2807,N_1253);
or U7223 (N_7223,N_1505,N_3240);
nor U7224 (N_7224,N_4484,N_1099);
nor U7225 (N_7225,N_996,N_1205);
nor U7226 (N_7226,N_1536,N_4956);
nor U7227 (N_7227,N_1657,N_4077);
or U7228 (N_7228,N_1683,N_1894);
or U7229 (N_7229,N_2616,N_3054);
and U7230 (N_7230,N_2052,N_1549);
xor U7231 (N_7231,N_4261,N_1921);
nor U7232 (N_7232,N_948,N_4252);
nand U7233 (N_7233,N_65,N_3968);
nand U7234 (N_7234,N_2757,N_1306);
or U7235 (N_7235,N_662,N_3634);
xor U7236 (N_7236,N_3273,N_1140);
xnor U7237 (N_7237,N_2973,N_2797);
or U7238 (N_7238,N_45,N_2456);
nor U7239 (N_7239,N_3443,N_908);
nor U7240 (N_7240,N_2424,N_4869);
nand U7241 (N_7241,N_1677,N_2554);
xnor U7242 (N_7242,N_2728,N_3965);
and U7243 (N_7243,N_2008,N_668);
nor U7244 (N_7244,N_2330,N_1757);
nand U7245 (N_7245,N_4917,N_2137);
xnor U7246 (N_7246,N_2001,N_2505);
xnor U7247 (N_7247,N_4190,N_1942);
or U7248 (N_7248,N_988,N_3451);
nor U7249 (N_7249,N_2446,N_4461);
or U7250 (N_7250,N_3911,N_2584);
nor U7251 (N_7251,N_3953,N_1668);
xor U7252 (N_7252,N_1189,N_655);
nand U7253 (N_7253,N_4186,N_679);
nor U7254 (N_7254,N_3739,N_565);
xnor U7255 (N_7255,N_3332,N_3808);
and U7256 (N_7256,N_4775,N_4867);
or U7257 (N_7257,N_1879,N_274);
or U7258 (N_7258,N_443,N_315);
xnor U7259 (N_7259,N_4653,N_4844);
xnor U7260 (N_7260,N_1172,N_1025);
or U7261 (N_7261,N_1874,N_1685);
xor U7262 (N_7262,N_3526,N_2193);
nand U7263 (N_7263,N_3817,N_4128);
or U7264 (N_7264,N_3294,N_2647);
or U7265 (N_7265,N_4652,N_3378);
nand U7266 (N_7266,N_906,N_3048);
or U7267 (N_7267,N_2469,N_1671);
nand U7268 (N_7268,N_2761,N_2029);
nand U7269 (N_7269,N_3955,N_698);
or U7270 (N_7270,N_2501,N_3386);
and U7271 (N_7271,N_2005,N_3053);
nor U7272 (N_7272,N_3588,N_2548);
nor U7273 (N_7273,N_1086,N_103);
and U7274 (N_7274,N_1105,N_4625);
nor U7275 (N_7275,N_4968,N_1234);
and U7276 (N_7276,N_991,N_4842);
xnor U7277 (N_7277,N_4914,N_1530);
or U7278 (N_7278,N_1698,N_723);
nand U7279 (N_7279,N_862,N_2979);
xnor U7280 (N_7280,N_2286,N_1217);
nand U7281 (N_7281,N_232,N_2347);
or U7282 (N_7282,N_3373,N_739);
nor U7283 (N_7283,N_4949,N_3755);
or U7284 (N_7284,N_4396,N_2677);
nor U7285 (N_7285,N_2329,N_4137);
or U7286 (N_7286,N_362,N_4180);
nor U7287 (N_7287,N_4656,N_2669);
nor U7288 (N_7288,N_3776,N_3460);
and U7289 (N_7289,N_3804,N_3663);
nand U7290 (N_7290,N_1094,N_1031);
nor U7291 (N_7291,N_381,N_4176);
and U7292 (N_7292,N_2266,N_1472);
nor U7293 (N_7293,N_1887,N_4460);
and U7294 (N_7294,N_3956,N_4751);
nor U7295 (N_7295,N_1483,N_2367);
or U7296 (N_7296,N_1324,N_4222);
nor U7297 (N_7297,N_3691,N_3828);
and U7298 (N_7298,N_1045,N_618);
xor U7299 (N_7299,N_1618,N_2682);
and U7300 (N_7300,N_3201,N_2312);
and U7301 (N_7301,N_4340,N_573);
nor U7302 (N_7302,N_1097,N_1595);
or U7303 (N_7303,N_2108,N_1835);
xnor U7304 (N_7304,N_290,N_1722);
and U7305 (N_7305,N_2912,N_4210);
nand U7306 (N_7306,N_3940,N_603);
and U7307 (N_7307,N_4893,N_4767);
xnor U7308 (N_7308,N_4994,N_3082);
and U7309 (N_7309,N_1133,N_2780);
xor U7310 (N_7310,N_4032,N_509);
and U7311 (N_7311,N_3374,N_941);
nand U7312 (N_7312,N_1540,N_861);
nand U7313 (N_7313,N_3699,N_4393);
and U7314 (N_7314,N_2282,N_4685);
and U7315 (N_7315,N_4527,N_1210);
or U7316 (N_7316,N_930,N_1498);
and U7317 (N_7317,N_3789,N_2915);
or U7318 (N_7318,N_2640,N_1665);
xnor U7319 (N_7319,N_3784,N_427);
nand U7320 (N_7320,N_1062,N_3662);
nor U7321 (N_7321,N_1676,N_160);
and U7322 (N_7322,N_451,N_1870);
nor U7323 (N_7323,N_190,N_725);
xor U7324 (N_7324,N_104,N_3848);
and U7325 (N_7325,N_2650,N_1755);
xor U7326 (N_7326,N_746,N_2038);
xor U7327 (N_7327,N_3704,N_2696);
or U7328 (N_7328,N_1159,N_4247);
nand U7329 (N_7329,N_3920,N_3697);
nor U7330 (N_7330,N_3916,N_1555);
or U7331 (N_7331,N_2946,N_1010);
or U7332 (N_7332,N_4884,N_4352);
and U7333 (N_7333,N_1859,N_2825);
and U7334 (N_7334,N_4066,N_3410);
xnor U7335 (N_7335,N_212,N_1594);
and U7336 (N_7336,N_2389,N_269);
nor U7337 (N_7337,N_4408,N_596);
xor U7338 (N_7338,N_2473,N_1688);
xnor U7339 (N_7339,N_40,N_2352);
or U7340 (N_7340,N_4202,N_3317);
and U7341 (N_7341,N_2621,N_1115);
or U7342 (N_7342,N_3768,N_3438);
xor U7343 (N_7343,N_2379,N_3389);
nor U7344 (N_7344,N_3604,N_2496);
xor U7345 (N_7345,N_4208,N_1038);
or U7346 (N_7346,N_4797,N_2648);
and U7347 (N_7347,N_2527,N_388);
and U7348 (N_7348,N_825,N_1739);
nor U7349 (N_7349,N_4443,N_3773);
and U7350 (N_7350,N_1669,N_833);
nand U7351 (N_7351,N_1069,N_3437);
and U7352 (N_7352,N_4774,N_3798);
nor U7353 (N_7353,N_4326,N_481);
nor U7354 (N_7354,N_1225,N_1351);
nand U7355 (N_7355,N_2438,N_2423);
nor U7356 (N_7356,N_1551,N_2011);
nand U7357 (N_7357,N_4262,N_1247);
nand U7358 (N_7358,N_3260,N_2184);
and U7359 (N_7359,N_2608,N_4799);
and U7360 (N_7360,N_2874,N_1421);
nor U7361 (N_7361,N_4521,N_2013);
or U7362 (N_7362,N_870,N_23);
and U7363 (N_7363,N_3860,N_3523);
xnor U7364 (N_7364,N_2465,N_3728);
xor U7365 (N_7365,N_4580,N_1604);
nor U7366 (N_7366,N_838,N_4655);
xnor U7367 (N_7367,N_1976,N_2576);
xor U7368 (N_7368,N_3398,N_3877);
nand U7369 (N_7369,N_2939,N_1509);
nor U7370 (N_7370,N_3429,N_4936);
nor U7371 (N_7371,N_3934,N_742);
or U7372 (N_7372,N_4816,N_3539);
nand U7373 (N_7373,N_2801,N_164);
or U7374 (N_7374,N_1129,N_1093);
and U7375 (N_7375,N_1191,N_1474);
and U7376 (N_7376,N_2906,N_1778);
xnor U7377 (N_7377,N_2599,N_4051);
or U7378 (N_7378,N_1015,N_3767);
xnor U7379 (N_7379,N_3213,N_53);
nand U7380 (N_7380,N_1018,N_1827);
or U7381 (N_7381,N_2653,N_3498);
nand U7382 (N_7382,N_3737,N_227);
or U7383 (N_7383,N_2194,N_1981);
nand U7384 (N_7384,N_2053,N_414);
or U7385 (N_7385,N_2783,N_922);
xor U7386 (N_7386,N_2944,N_939);
and U7387 (N_7387,N_2431,N_1699);
xor U7388 (N_7388,N_600,N_1180);
xnor U7389 (N_7389,N_2727,N_4305);
nand U7390 (N_7390,N_4297,N_3208);
and U7391 (N_7391,N_2091,N_2395);
and U7392 (N_7392,N_2092,N_3516);
and U7393 (N_7393,N_4099,N_805);
and U7394 (N_7394,N_134,N_436);
nor U7395 (N_7395,N_2503,N_27);
xor U7396 (N_7396,N_2947,N_1059);
and U7397 (N_7397,N_310,N_2966);
nand U7398 (N_7398,N_348,N_1938);
nor U7399 (N_7399,N_863,N_2084);
nand U7400 (N_7400,N_2129,N_721);
and U7401 (N_7401,N_2821,N_1727);
and U7402 (N_7402,N_4275,N_766);
nor U7403 (N_7403,N_4233,N_2935);
xor U7404 (N_7404,N_4743,N_3871);
nor U7405 (N_7405,N_4718,N_683);
nor U7406 (N_7406,N_2962,N_1352);
nor U7407 (N_7407,N_4394,N_1880);
xor U7408 (N_7408,N_4704,N_2327);
or U7409 (N_7409,N_4119,N_4966);
nand U7410 (N_7410,N_1559,N_2943);
xnor U7411 (N_7411,N_4632,N_864);
or U7412 (N_7412,N_2307,N_3400);
nand U7413 (N_7413,N_4700,N_4438);
nor U7414 (N_7414,N_16,N_1915);
nor U7415 (N_7415,N_3291,N_887);
or U7416 (N_7416,N_1000,N_1568);
nor U7417 (N_7417,N_2349,N_1241);
and U7418 (N_7418,N_1523,N_754);
xnor U7419 (N_7419,N_137,N_2195);
or U7420 (N_7420,N_895,N_2919);
and U7421 (N_7421,N_2059,N_704);
nand U7422 (N_7422,N_2297,N_4736);
nand U7423 (N_7423,N_1168,N_228);
nor U7424 (N_7424,N_3329,N_757);
nand U7425 (N_7425,N_3179,N_762);
nand U7426 (N_7426,N_2815,N_1852);
nor U7427 (N_7427,N_4047,N_1986);
and U7428 (N_7428,N_1636,N_205);
xnor U7429 (N_7429,N_3951,N_1165);
or U7430 (N_7430,N_885,N_3263);
nand U7431 (N_7431,N_1917,N_4195);
nor U7432 (N_7432,N_2600,N_2949);
or U7433 (N_7433,N_2208,N_3063);
or U7434 (N_7434,N_2003,N_1143);
and U7435 (N_7435,N_1397,N_4916);
xor U7436 (N_7436,N_806,N_13);
or U7437 (N_7437,N_397,N_1091);
nor U7438 (N_7438,N_4030,N_3577);
nand U7439 (N_7439,N_3542,N_169);
or U7440 (N_7440,N_3130,N_4173);
nand U7441 (N_7441,N_877,N_3186);
or U7442 (N_7442,N_8,N_54);
and U7443 (N_7443,N_3093,N_3340);
nand U7444 (N_7444,N_2601,N_4720);
nand U7445 (N_7445,N_3541,N_286);
nor U7446 (N_7446,N_2981,N_167);
nand U7447 (N_7447,N_324,N_3068);
xnor U7448 (N_7448,N_2739,N_2586);
or U7449 (N_7449,N_4269,N_1765);
nand U7450 (N_7450,N_2953,N_4420);
nand U7451 (N_7451,N_3444,N_4965);
nand U7452 (N_7452,N_2057,N_3167);
nand U7453 (N_7453,N_964,N_4418);
nor U7454 (N_7454,N_2310,N_849);
nor U7455 (N_7455,N_1005,N_461);
nor U7456 (N_7456,N_534,N_4090);
xor U7457 (N_7457,N_1173,N_1207);
nand U7458 (N_7458,N_4591,N_1682);
xnor U7459 (N_7459,N_1329,N_3056);
or U7460 (N_7460,N_2818,N_4827);
nor U7461 (N_7461,N_829,N_3701);
xor U7462 (N_7462,N_1357,N_2646);
and U7463 (N_7463,N_4426,N_1392);
or U7464 (N_7464,N_3360,N_732);
nand U7465 (N_7465,N_1176,N_4519);
and U7466 (N_7466,N_4678,N_548);
nand U7467 (N_7467,N_1864,N_1125);
or U7468 (N_7468,N_2574,N_4534);
or U7469 (N_7469,N_1473,N_1531);
nand U7470 (N_7470,N_1330,N_1899);
nand U7471 (N_7471,N_2592,N_3);
nor U7472 (N_7472,N_225,N_506);
xor U7473 (N_7473,N_1605,N_2558);
nand U7474 (N_7474,N_3614,N_997);
and U7475 (N_7475,N_3503,N_3760);
or U7476 (N_7476,N_2959,N_2293);
xor U7477 (N_7477,N_3723,N_70);
xor U7478 (N_7478,N_1348,N_532);
nand U7479 (N_7479,N_4573,N_2497);
xor U7480 (N_7480,N_2135,N_3490);
or U7481 (N_7481,N_4870,N_1666);
nand U7482 (N_7482,N_4328,N_3559);
nand U7483 (N_7483,N_3259,N_2596);
xnor U7484 (N_7484,N_3455,N_677);
nand U7485 (N_7485,N_4234,N_3343);
nor U7486 (N_7486,N_3365,N_3573);
nor U7487 (N_7487,N_1570,N_3623);
and U7488 (N_7488,N_2976,N_4371);
and U7489 (N_7489,N_4499,N_3669);
nand U7490 (N_7490,N_803,N_2778);
or U7491 (N_7491,N_4862,N_1719);
nand U7492 (N_7492,N_693,N_2475);
xor U7493 (N_7493,N_1628,N_1931);
nand U7494 (N_7494,N_2123,N_28);
xor U7495 (N_7495,N_3675,N_585);
or U7496 (N_7496,N_3851,N_4590);
and U7497 (N_7497,N_425,N_4241);
nor U7498 (N_7498,N_731,N_4809);
and U7499 (N_7499,N_3973,N_1373);
nand U7500 (N_7500,N_3747,N_338);
or U7501 (N_7501,N_1994,N_2542);
nor U7502 (N_7502,N_1013,N_1612);
and U7503 (N_7503,N_4462,N_3199);
xnor U7504 (N_7504,N_2440,N_3314);
and U7505 (N_7505,N_348,N_2263);
and U7506 (N_7506,N_1858,N_4607);
and U7507 (N_7507,N_889,N_3245);
and U7508 (N_7508,N_2899,N_3856);
xnor U7509 (N_7509,N_2514,N_826);
nand U7510 (N_7510,N_4855,N_4930);
or U7511 (N_7511,N_1110,N_4445);
or U7512 (N_7512,N_1538,N_4809);
and U7513 (N_7513,N_3083,N_2875);
xor U7514 (N_7514,N_2940,N_3348);
nand U7515 (N_7515,N_1206,N_4154);
xnor U7516 (N_7516,N_3535,N_4619);
or U7517 (N_7517,N_2993,N_182);
and U7518 (N_7518,N_4523,N_3185);
xnor U7519 (N_7519,N_1101,N_3251);
xor U7520 (N_7520,N_2025,N_3414);
xor U7521 (N_7521,N_1068,N_4948);
xor U7522 (N_7522,N_2309,N_1184);
xnor U7523 (N_7523,N_3543,N_3999);
or U7524 (N_7524,N_4537,N_1891);
nor U7525 (N_7525,N_948,N_4732);
xor U7526 (N_7526,N_3370,N_3857);
nand U7527 (N_7527,N_2579,N_4193);
xor U7528 (N_7528,N_1433,N_1944);
xor U7529 (N_7529,N_1021,N_1627);
nor U7530 (N_7530,N_796,N_3200);
or U7531 (N_7531,N_3317,N_4220);
and U7532 (N_7532,N_2722,N_1331);
nor U7533 (N_7533,N_3273,N_306);
and U7534 (N_7534,N_2757,N_4817);
and U7535 (N_7535,N_1911,N_3418);
nand U7536 (N_7536,N_1622,N_2898);
or U7537 (N_7537,N_577,N_4439);
xnor U7538 (N_7538,N_1185,N_1361);
or U7539 (N_7539,N_3889,N_140);
nor U7540 (N_7540,N_2675,N_3578);
and U7541 (N_7541,N_1931,N_68);
xnor U7542 (N_7542,N_4232,N_521);
or U7543 (N_7543,N_3896,N_817);
or U7544 (N_7544,N_1110,N_636);
nor U7545 (N_7545,N_2222,N_759);
nor U7546 (N_7546,N_3432,N_37);
and U7547 (N_7547,N_21,N_392);
nor U7548 (N_7548,N_3459,N_421);
and U7549 (N_7549,N_4167,N_1133);
and U7550 (N_7550,N_278,N_4899);
and U7551 (N_7551,N_2495,N_2173);
and U7552 (N_7552,N_3204,N_3164);
or U7553 (N_7553,N_1210,N_1128);
nor U7554 (N_7554,N_4388,N_3602);
nor U7555 (N_7555,N_1784,N_4611);
and U7556 (N_7556,N_1225,N_3356);
xnor U7557 (N_7557,N_3992,N_2047);
nor U7558 (N_7558,N_3987,N_2221);
or U7559 (N_7559,N_3504,N_1231);
and U7560 (N_7560,N_4609,N_4479);
nand U7561 (N_7561,N_2746,N_2976);
nor U7562 (N_7562,N_2416,N_682);
xor U7563 (N_7563,N_2832,N_3420);
or U7564 (N_7564,N_3967,N_4225);
and U7565 (N_7565,N_3129,N_2735);
and U7566 (N_7566,N_3499,N_3762);
and U7567 (N_7567,N_2615,N_2395);
and U7568 (N_7568,N_616,N_2656);
xor U7569 (N_7569,N_1215,N_3659);
or U7570 (N_7570,N_2866,N_1130);
nand U7571 (N_7571,N_2554,N_4565);
and U7572 (N_7572,N_4023,N_922);
nor U7573 (N_7573,N_436,N_4656);
or U7574 (N_7574,N_3818,N_2531);
nand U7575 (N_7575,N_154,N_4674);
nand U7576 (N_7576,N_3686,N_3524);
nor U7577 (N_7577,N_3378,N_2773);
nand U7578 (N_7578,N_1037,N_794);
or U7579 (N_7579,N_2595,N_2439);
xor U7580 (N_7580,N_2913,N_1814);
or U7581 (N_7581,N_86,N_1524);
xnor U7582 (N_7582,N_3202,N_2472);
nand U7583 (N_7583,N_615,N_4361);
or U7584 (N_7584,N_4675,N_2562);
and U7585 (N_7585,N_4577,N_2085);
or U7586 (N_7586,N_3965,N_30);
nor U7587 (N_7587,N_426,N_2595);
xor U7588 (N_7588,N_2220,N_1145);
or U7589 (N_7589,N_2805,N_3442);
xnor U7590 (N_7590,N_3747,N_2543);
nor U7591 (N_7591,N_109,N_2681);
and U7592 (N_7592,N_3996,N_3362);
or U7593 (N_7593,N_2401,N_3);
or U7594 (N_7594,N_3606,N_3905);
or U7595 (N_7595,N_1283,N_3499);
nor U7596 (N_7596,N_1408,N_3840);
or U7597 (N_7597,N_2332,N_1469);
or U7598 (N_7598,N_3444,N_4551);
nand U7599 (N_7599,N_180,N_629);
xor U7600 (N_7600,N_1690,N_2425);
nand U7601 (N_7601,N_3924,N_3742);
or U7602 (N_7602,N_3469,N_484);
or U7603 (N_7603,N_354,N_2679);
nor U7604 (N_7604,N_2311,N_2214);
or U7605 (N_7605,N_2915,N_3503);
or U7606 (N_7606,N_3250,N_1682);
or U7607 (N_7607,N_3593,N_1799);
nand U7608 (N_7608,N_3827,N_2882);
nor U7609 (N_7609,N_4191,N_1543);
xor U7610 (N_7610,N_3181,N_2715);
nand U7611 (N_7611,N_2734,N_4884);
and U7612 (N_7612,N_3403,N_4566);
or U7613 (N_7613,N_1311,N_2282);
nor U7614 (N_7614,N_2963,N_4591);
and U7615 (N_7615,N_2148,N_233);
nand U7616 (N_7616,N_4007,N_1503);
or U7617 (N_7617,N_2785,N_1419);
nor U7618 (N_7618,N_594,N_3822);
and U7619 (N_7619,N_47,N_2247);
or U7620 (N_7620,N_326,N_3871);
and U7621 (N_7621,N_2914,N_442);
and U7622 (N_7622,N_3430,N_4907);
xnor U7623 (N_7623,N_3177,N_4753);
and U7624 (N_7624,N_1688,N_4021);
or U7625 (N_7625,N_2598,N_2868);
xnor U7626 (N_7626,N_2716,N_3779);
nor U7627 (N_7627,N_1739,N_3293);
or U7628 (N_7628,N_3121,N_3607);
and U7629 (N_7629,N_4640,N_4075);
or U7630 (N_7630,N_2031,N_4461);
nand U7631 (N_7631,N_3693,N_4904);
nor U7632 (N_7632,N_2567,N_4921);
nand U7633 (N_7633,N_3721,N_203);
nand U7634 (N_7634,N_4358,N_4379);
or U7635 (N_7635,N_4813,N_3064);
and U7636 (N_7636,N_2664,N_1286);
nor U7637 (N_7637,N_1141,N_1789);
nor U7638 (N_7638,N_4022,N_4668);
and U7639 (N_7639,N_3854,N_2940);
or U7640 (N_7640,N_2961,N_2297);
and U7641 (N_7641,N_4645,N_3919);
and U7642 (N_7642,N_2920,N_2234);
or U7643 (N_7643,N_426,N_1029);
and U7644 (N_7644,N_542,N_4322);
or U7645 (N_7645,N_3059,N_2692);
nor U7646 (N_7646,N_4720,N_3324);
or U7647 (N_7647,N_2202,N_590);
xor U7648 (N_7648,N_2667,N_822);
nand U7649 (N_7649,N_3756,N_682);
or U7650 (N_7650,N_3425,N_4038);
nand U7651 (N_7651,N_934,N_203);
nand U7652 (N_7652,N_2455,N_4633);
xnor U7653 (N_7653,N_4489,N_2439);
and U7654 (N_7654,N_3441,N_319);
or U7655 (N_7655,N_3938,N_1342);
nor U7656 (N_7656,N_2539,N_3501);
xor U7657 (N_7657,N_2572,N_322);
and U7658 (N_7658,N_44,N_117);
and U7659 (N_7659,N_1545,N_133);
or U7660 (N_7660,N_4933,N_326);
nand U7661 (N_7661,N_2267,N_3488);
and U7662 (N_7662,N_4040,N_3952);
nor U7663 (N_7663,N_2701,N_3563);
or U7664 (N_7664,N_2439,N_1238);
or U7665 (N_7665,N_2874,N_1464);
nand U7666 (N_7666,N_461,N_639);
and U7667 (N_7667,N_1112,N_3732);
or U7668 (N_7668,N_2994,N_1131);
and U7669 (N_7669,N_3772,N_267);
and U7670 (N_7670,N_3864,N_3234);
nand U7671 (N_7671,N_2858,N_4282);
nand U7672 (N_7672,N_3717,N_3555);
or U7673 (N_7673,N_2579,N_2778);
nor U7674 (N_7674,N_3622,N_3238);
and U7675 (N_7675,N_1428,N_3971);
or U7676 (N_7676,N_2891,N_4686);
nand U7677 (N_7677,N_4895,N_4533);
nor U7678 (N_7678,N_867,N_2152);
and U7679 (N_7679,N_4694,N_4145);
nand U7680 (N_7680,N_1418,N_508);
or U7681 (N_7681,N_2225,N_1420);
or U7682 (N_7682,N_2476,N_3785);
xnor U7683 (N_7683,N_1329,N_3216);
or U7684 (N_7684,N_2083,N_686);
and U7685 (N_7685,N_2156,N_1349);
nor U7686 (N_7686,N_866,N_2312);
nand U7687 (N_7687,N_2426,N_2810);
nor U7688 (N_7688,N_1987,N_3912);
xnor U7689 (N_7689,N_4405,N_207);
or U7690 (N_7690,N_531,N_1077);
nor U7691 (N_7691,N_1109,N_324);
nor U7692 (N_7692,N_3212,N_1908);
nand U7693 (N_7693,N_4574,N_1081);
nor U7694 (N_7694,N_1639,N_4433);
or U7695 (N_7695,N_4288,N_1694);
nor U7696 (N_7696,N_2425,N_2499);
and U7697 (N_7697,N_90,N_1929);
xor U7698 (N_7698,N_2193,N_1790);
nand U7699 (N_7699,N_113,N_4113);
nor U7700 (N_7700,N_4343,N_3043);
and U7701 (N_7701,N_189,N_3416);
nor U7702 (N_7702,N_3171,N_1507);
nor U7703 (N_7703,N_699,N_3504);
nor U7704 (N_7704,N_3062,N_4352);
nand U7705 (N_7705,N_4590,N_2179);
and U7706 (N_7706,N_2879,N_3467);
nor U7707 (N_7707,N_1751,N_413);
xor U7708 (N_7708,N_2445,N_113);
nor U7709 (N_7709,N_511,N_1306);
and U7710 (N_7710,N_1843,N_4857);
nand U7711 (N_7711,N_145,N_2123);
and U7712 (N_7712,N_1595,N_2705);
or U7713 (N_7713,N_3324,N_3833);
and U7714 (N_7714,N_962,N_4503);
or U7715 (N_7715,N_200,N_3832);
or U7716 (N_7716,N_1987,N_3772);
nand U7717 (N_7717,N_1124,N_744);
nor U7718 (N_7718,N_2905,N_2336);
nor U7719 (N_7719,N_1642,N_490);
and U7720 (N_7720,N_341,N_3506);
nand U7721 (N_7721,N_2573,N_3659);
and U7722 (N_7722,N_4240,N_4481);
nor U7723 (N_7723,N_2488,N_4578);
nor U7724 (N_7724,N_2901,N_2487);
nor U7725 (N_7725,N_852,N_3500);
nor U7726 (N_7726,N_4160,N_4829);
xor U7727 (N_7727,N_3161,N_3235);
nand U7728 (N_7728,N_122,N_699);
nand U7729 (N_7729,N_3348,N_18);
nor U7730 (N_7730,N_4626,N_665);
or U7731 (N_7731,N_2326,N_708);
or U7732 (N_7732,N_425,N_1906);
and U7733 (N_7733,N_2643,N_4481);
nand U7734 (N_7734,N_2086,N_912);
xor U7735 (N_7735,N_3223,N_255);
nor U7736 (N_7736,N_4514,N_961);
xor U7737 (N_7737,N_3699,N_1083);
or U7738 (N_7738,N_3347,N_922);
nand U7739 (N_7739,N_3089,N_2255);
or U7740 (N_7740,N_1871,N_476);
nor U7741 (N_7741,N_4350,N_3151);
nand U7742 (N_7742,N_3532,N_3682);
nand U7743 (N_7743,N_4121,N_498);
xor U7744 (N_7744,N_2753,N_4915);
and U7745 (N_7745,N_4811,N_2287);
nand U7746 (N_7746,N_4913,N_3041);
or U7747 (N_7747,N_3409,N_3105);
nand U7748 (N_7748,N_3938,N_4892);
nor U7749 (N_7749,N_1197,N_984);
nor U7750 (N_7750,N_2451,N_4724);
nand U7751 (N_7751,N_4253,N_1206);
nand U7752 (N_7752,N_3069,N_4942);
or U7753 (N_7753,N_2596,N_657);
xor U7754 (N_7754,N_2017,N_1275);
xor U7755 (N_7755,N_3246,N_2252);
xnor U7756 (N_7756,N_2406,N_2683);
xnor U7757 (N_7757,N_3675,N_252);
or U7758 (N_7758,N_4336,N_3161);
nand U7759 (N_7759,N_1759,N_3841);
and U7760 (N_7760,N_3440,N_4898);
nor U7761 (N_7761,N_4406,N_1489);
xnor U7762 (N_7762,N_3727,N_1604);
or U7763 (N_7763,N_408,N_877);
nor U7764 (N_7764,N_1072,N_4414);
or U7765 (N_7765,N_3109,N_265);
xor U7766 (N_7766,N_3878,N_2668);
xnor U7767 (N_7767,N_3014,N_3910);
and U7768 (N_7768,N_2829,N_4185);
nand U7769 (N_7769,N_2877,N_3721);
or U7770 (N_7770,N_4449,N_1643);
or U7771 (N_7771,N_305,N_2895);
xor U7772 (N_7772,N_3074,N_3706);
and U7773 (N_7773,N_332,N_2160);
nand U7774 (N_7774,N_4822,N_3651);
nor U7775 (N_7775,N_26,N_2439);
nor U7776 (N_7776,N_277,N_4355);
nand U7777 (N_7777,N_2593,N_2253);
and U7778 (N_7778,N_1989,N_229);
nand U7779 (N_7779,N_81,N_3006);
xnor U7780 (N_7780,N_1485,N_4540);
xnor U7781 (N_7781,N_517,N_1751);
nand U7782 (N_7782,N_1027,N_2204);
nor U7783 (N_7783,N_326,N_4722);
nand U7784 (N_7784,N_581,N_1191);
and U7785 (N_7785,N_3328,N_4197);
xnor U7786 (N_7786,N_514,N_1367);
nand U7787 (N_7787,N_4651,N_4267);
nand U7788 (N_7788,N_110,N_2283);
or U7789 (N_7789,N_4187,N_2446);
nor U7790 (N_7790,N_3603,N_1436);
nand U7791 (N_7791,N_957,N_2156);
nor U7792 (N_7792,N_3863,N_2159);
and U7793 (N_7793,N_2913,N_2808);
or U7794 (N_7794,N_4089,N_4656);
or U7795 (N_7795,N_2211,N_4321);
and U7796 (N_7796,N_2554,N_1268);
nor U7797 (N_7797,N_1805,N_3326);
or U7798 (N_7798,N_3169,N_2521);
nand U7799 (N_7799,N_3503,N_4114);
nand U7800 (N_7800,N_2514,N_4404);
nor U7801 (N_7801,N_4578,N_2284);
nand U7802 (N_7802,N_1580,N_854);
nor U7803 (N_7803,N_2692,N_3631);
and U7804 (N_7804,N_1993,N_4223);
or U7805 (N_7805,N_2499,N_3540);
xor U7806 (N_7806,N_661,N_4688);
nand U7807 (N_7807,N_4059,N_4260);
xor U7808 (N_7808,N_1043,N_157);
xor U7809 (N_7809,N_1911,N_3595);
or U7810 (N_7810,N_1892,N_1699);
xor U7811 (N_7811,N_3061,N_101);
nand U7812 (N_7812,N_3285,N_1267);
and U7813 (N_7813,N_4738,N_4787);
nor U7814 (N_7814,N_3997,N_3527);
xnor U7815 (N_7815,N_4171,N_4486);
and U7816 (N_7816,N_3402,N_3072);
or U7817 (N_7817,N_702,N_3196);
or U7818 (N_7818,N_1059,N_2578);
nand U7819 (N_7819,N_4534,N_2186);
xnor U7820 (N_7820,N_3991,N_4807);
nand U7821 (N_7821,N_1719,N_4268);
and U7822 (N_7822,N_1929,N_2236);
nor U7823 (N_7823,N_4543,N_4203);
and U7824 (N_7824,N_867,N_4492);
nand U7825 (N_7825,N_3691,N_3098);
and U7826 (N_7826,N_1578,N_800);
nand U7827 (N_7827,N_842,N_501);
xnor U7828 (N_7828,N_3575,N_3448);
nor U7829 (N_7829,N_2773,N_74);
or U7830 (N_7830,N_1288,N_2633);
and U7831 (N_7831,N_2403,N_1068);
and U7832 (N_7832,N_3691,N_3892);
nand U7833 (N_7833,N_1877,N_4189);
xor U7834 (N_7834,N_3721,N_4818);
or U7835 (N_7835,N_960,N_95);
and U7836 (N_7836,N_2374,N_2479);
or U7837 (N_7837,N_846,N_50);
xor U7838 (N_7838,N_3279,N_2599);
nor U7839 (N_7839,N_1419,N_3443);
nor U7840 (N_7840,N_4181,N_299);
or U7841 (N_7841,N_3179,N_417);
and U7842 (N_7842,N_3433,N_1339);
and U7843 (N_7843,N_1855,N_2550);
nand U7844 (N_7844,N_1620,N_3183);
nor U7845 (N_7845,N_2863,N_2868);
nand U7846 (N_7846,N_1152,N_561);
xor U7847 (N_7847,N_2721,N_2309);
and U7848 (N_7848,N_2983,N_4894);
and U7849 (N_7849,N_418,N_2252);
nand U7850 (N_7850,N_1080,N_4300);
nand U7851 (N_7851,N_901,N_2630);
nand U7852 (N_7852,N_4740,N_2283);
nand U7853 (N_7853,N_2233,N_2170);
and U7854 (N_7854,N_2274,N_2462);
nor U7855 (N_7855,N_1417,N_2371);
xor U7856 (N_7856,N_4244,N_3902);
nand U7857 (N_7857,N_3545,N_1986);
nor U7858 (N_7858,N_3174,N_584);
nor U7859 (N_7859,N_3960,N_3084);
and U7860 (N_7860,N_4692,N_979);
nand U7861 (N_7861,N_722,N_2483);
nor U7862 (N_7862,N_3856,N_2248);
nand U7863 (N_7863,N_2285,N_312);
nor U7864 (N_7864,N_663,N_3191);
or U7865 (N_7865,N_924,N_2600);
or U7866 (N_7866,N_3973,N_1001);
xnor U7867 (N_7867,N_1632,N_2623);
nor U7868 (N_7868,N_1865,N_903);
and U7869 (N_7869,N_1135,N_2074);
nand U7870 (N_7870,N_3686,N_3443);
xnor U7871 (N_7871,N_3203,N_3924);
xor U7872 (N_7872,N_3762,N_2830);
xor U7873 (N_7873,N_2518,N_4893);
nor U7874 (N_7874,N_4885,N_409);
nor U7875 (N_7875,N_1401,N_2491);
xnor U7876 (N_7876,N_1549,N_135);
nand U7877 (N_7877,N_3146,N_3063);
and U7878 (N_7878,N_3511,N_4855);
or U7879 (N_7879,N_4685,N_3921);
nor U7880 (N_7880,N_1565,N_343);
or U7881 (N_7881,N_4767,N_686);
nor U7882 (N_7882,N_4849,N_371);
or U7883 (N_7883,N_4458,N_2315);
nor U7884 (N_7884,N_4343,N_663);
nand U7885 (N_7885,N_4263,N_176);
nand U7886 (N_7886,N_4823,N_4758);
xor U7887 (N_7887,N_1417,N_2206);
nor U7888 (N_7888,N_178,N_1544);
and U7889 (N_7889,N_763,N_631);
nor U7890 (N_7890,N_4381,N_1346);
nand U7891 (N_7891,N_4647,N_89);
and U7892 (N_7892,N_4976,N_2640);
or U7893 (N_7893,N_2214,N_4642);
and U7894 (N_7894,N_847,N_3486);
or U7895 (N_7895,N_1416,N_4984);
nor U7896 (N_7896,N_3929,N_4628);
and U7897 (N_7897,N_596,N_390);
nand U7898 (N_7898,N_1182,N_2896);
or U7899 (N_7899,N_2820,N_4903);
and U7900 (N_7900,N_2189,N_2582);
xor U7901 (N_7901,N_1088,N_3471);
nor U7902 (N_7902,N_1258,N_284);
nand U7903 (N_7903,N_3902,N_2556);
and U7904 (N_7904,N_3307,N_3401);
nand U7905 (N_7905,N_4836,N_3814);
xnor U7906 (N_7906,N_1406,N_1170);
nand U7907 (N_7907,N_2389,N_4263);
nand U7908 (N_7908,N_3480,N_4510);
or U7909 (N_7909,N_4878,N_700);
or U7910 (N_7910,N_4042,N_4773);
nor U7911 (N_7911,N_4908,N_3598);
nand U7912 (N_7912,N_1730,N_348);
or U7913 (N_7913,N_1092,N_1638);
xor U7914 (N_7914,N_4901,N_1473);
nor U7915 (N_7915,N_3771,N_4300);
xnor U7916 (N_7916,N_1617,N_1874);
nor U7917 (N_7917,N_4625,N_4156);
and U7918 (N_7918,N_4238,N_4595);
nor U7919 (N_7919,N_4960,N_3670);
and U7920 (N_7920,N_4827,N_1079);
nor U7921 (N_7921,N_4355,N_3579);
or U7922 (N_7922,N_2357,N_1066);
xnor U7923 (N_7923,N_3812,N_899);
xnor U7924 (N_7924,N_3797,N_99);
or U7925 (N_7925,N_3186,N_2299);
nor U7926 (N_7926,N_2272,N_4467);
and U7927 (N_7927,N_1210,N_743);
and U7928 (N_7928,N_1352,N_4810);
nand U7929 (N_7929,N_601,N_3567);
or U7930 (N_7930,N_3795,N_4408);
xnor U7931 (N_7931,N_397,N_114);
xnor U7932 (N_7932,N_1815,N_2902);
nand U7933 (N_7933,N_3760,N_1821);
nor U7934 (N_7934,N_3420,N_2256);
or U7935 (N_7935,N_3498,N_3398);
nand U7936 (N_7936,N_2684,N_780);
nand U7937 (N_7937,N_3433,N_4605);
and U7938 (N_7938,N_4088,N_2384);
nor U7939 (N_7939,N_4242,N_4926);
xor U7940 (N_7940,N_134,N_3315);
or U7941 (N_7941,N_1868,N_4924);
xnor U7942 (N_7942,N_1635,N_3799);
or U7943 (N_7943,N_1014,N_2208);
nand U7944 (N_7944,N_3395,N_1315);
xnor U7945 (N_7945,N_1375,N_1270);
nand U7946 (N_7946,N_1593,N_4567);
nor U7947 (N_7947,N_4933,N_2287);
or U7948 (N_7948,N_3246,N_2702);
or U7949 (N_7949,N_4851,N_4626);
nor U7950 (N_7950,N_567,N_3865);
and U7951 (N_7951,N_4585,N_1036);
nor U7952 (N_7952,N_3957,N_3043);
xor U7953 (N_7953,N_2285,N_738);
nor U7954 (N_7954,N_4760,N_1874);
nor U7955 (N_7955,N_2549,N_1976);
or U7956 (N_7956,N_1014,N_4276);
nor U7957 (N_7957,N_862,N_4394);
nor U7958 (N_7958,N_3155,N_2171);
nand U7959 (N_7959,N_480,N_3983);
or U7960 (N_7960,N_1799,N_3511);
nand U7961 (N_7961,N_535,N_4076);
xor U7962 (N_7962,N_1415,N_3035);
and U7963 (N_7963,N_4439,N_4182);
and U7964 (N_7964,N_1307,N_2923);
nor U7965 (N_7965,N_4400,N_524);
and U7966 (N_7966,N_2539,N_2827);
xnor U7967 (N_7967,N_1143,N_2676);
or U7968 (N_7968,N_2242,N_2755);
and U7969 (N_7969,N_2582,N_4436);
or U7970 (N_7970,N_978,N_383);
or U7971 (N_7971,N_1456,N_3212);
or U7972 (N_7972,N_4401,N_2660);
nor U7973 (N_7973,N_2256,N_4589);
and U7974 (N_7974,N_3373,N_3733);
nor U7975 (N_7975,N_1274,N_3767);
nand U7976 (N_7976,N_2982,N_1111);
or U7977 (N_7977,N_931,N_3640);
xnor U7978 (N_7978,N_4076,N_1096);
or U7979 (N_7979,N_3441,N_701);
nor U7980 (N_7980,N_3606,N_4670);
nor U7981 (N_7981,N_4461,N_2968);
or U7982 (N_7982,N_2282,N_10);
nand U7983 (N_7983,N_4521,N_4010);
or U7984 (N_7984,N_2744,N_802);
nor U7985 (N_7985,N_4390,N_4260);
xnor U7986 (N_7986,N_1695,N_521);
nand U7987 (N_7987,N_4558,N_4767);
xor U7988 (N_7988,N_410,N_1334);
nand U7989 (N_7989,N_3170,N_2400);
nand U7990 (N_7990,N_3412,N_1444);
nor U7991 (N_7991,N_1788,N_2113);
or U7992 (N_7992,N_1887,N_2035);
and U7993 (N_7993,N_1676,N_4924);
and U7994 (N_7994,N_798,N_4236);
or U7995 (N_7995,N_2264,N_2237);
and U7996 (N_7996,N_4116,N_2043);
nand U7997 (N_7997,N_3939,N_3272);
nor U7998 (N_7998,N_3858,N_4049);
nand U7999 (N_7999,N_2924,N_2613);
nor U8000 (N_8000,N_1854,N_269);
and U8001 (N_8001,N_1792,N_1245);
and U8002 (N_8002,N_4879,N_3235);
or U8003 (N_8003,N_4031,N_1606);
and U8004 (N_8004,N_4532,N_4995);
xnor U8005 (N_8005,N_3438,N_1891);
or U8006 (N_8006,N_4003,N_3199);
nor U8007 (N_8007,N_2382,N_2612);
xnor U8008 (N_8008,N_4228,N_4095);
and U8009 (N_8009,N_1384,N_2550);
or U8010 (N_8010,N_2612,N_3756);
nor U8011 (N_8011,N_1748,N_4506);
nor U8012 (N_8012,N_1064,N_2070);
nand U8013 (N_8013,N_3803,N_3220);
nor U8014 (N_8014,N_185,N_4772);
nor U8015 (N_8015,N_2450,N_2268);
nand U8016 (N_8016,N_377,N_53);
nand U8017 (N_8017,N_3027,N_3981);
xor U8018 (N_8018,N_3388,N_961);
or U8019 (N_8019,N_1814,N_3090);
or U8020 (N_8020,N_3811,N_4989);
nor U8021 (N_8021,N_1921,N_2351);
nor U8022 (N_8022,N_928,N_3308);
and U8023 (N_8023,N_2744,N_4679);
xor U8024 (N_8024,N_3567,N_2123);
nand U8025 (N_8025,N_2523,N_4718);
and U8026 (N_8026,N_137,N_2386);
nor U8027 (N_8027,N_996,N_1724);
xor U8028 (N_8028,N_208,N_364);
or U8029 (N_8029,N_494,N_543);
and U8030 (N_8030,N_1024,N_363);
nand U8031 (N_8031,N_4139,N_2589);
and U8032 (N_8032,N_3130,N_2767);
or U8033 (N_8033,N_229,N_1008);
nand U8034 (N_8034,N_4594,N_4712);
nand U8035 (N_8035,N_2718,N_3026);
or U8036 (N_8036,N_595,N_669);
and U8037 (N_8037,N_4719,N_777);
or U8038 (N_8038,N_2686,N_1705);
xnor U8039 (N_8039,N_1284,N_724);
or U8040 (N_8040,N_4886,N_326);
or U8041 (N_8041,N_2168,N_4174);
nand U8042 (N_8042,N_2338,N_4906);
nand U8043 (N_8043,N_130,N_1831);
and U8044 (N_8044,N_3410,N_2148);
or U8045 (N_8045,N_1306,N_4314);
and U8046 (N_8046,N_1115,N_4456);
or U8047 (N_8047,N_2122,N_4458);
nand U8048 (N_8048,N_3480,N_3793);
nor U8049 (N_8049,N_2565,N_3377);
or U8050 (N_8050,N_2820,N_3207);
nand U8051 (N_8051,N_2654,N_2554);
nor U8052 (N_8052,N_217,N_1759);
xnor U8053 (N_8053,N_419,N_2093);
xor U8054 (N_8054,N_4569,N_4484);
xnor U8055 (N_8055,N_1868,N_1522);
nor U8056 (N_8056,N_2914,N_4939);
nand U8057 (N_8057,N_4584,N_2231);
and U8058 (N_8058,N_4134,N_2063);
and U8059 (N_8059,N_1508,N_2289);
nand U8060 (N_8060,N_2993,N_107);
nand U8061 (N_8061,N_992,N_4185);
and U8062 (N_8062,N_858,N_709);
and U8063 (N_8063,N_2844,N_1492);
nor U8064 (N_8064,N_4110,N_1702);
xor U8065 (N_8065,N_486,N_1014);
xnor U8066 (N_8066,N_1941,N_1543);
xor U8067 (N_8067,N_4809,N_1230);
or U8068 (N_8068,N_570,N_714);
nor U8069 (N_8069,N_1619,N_935);
xor U8070 (N_8070,N_249,N_1613);
nor U8071 (N_8071,N_2632,N_715);
or U8072 (N_8072,N_1690,N_583);
nor U8073 (N_8073,N_1490,N_4439);
nand U8074 (N_8074,N_3515,N_1674);
nor U8075 (N_8075,N_1750,N_1104);
xnor U8076 (N_8076,N_1988,N_3591);
xnor U8077 (N_8077,N_2760,N_1520);
nand U8078 (N_8078,N_4495,N_1988);
nand U8079 (N_8079,N_3930,N_1604);
and U8080 (N_8080,N_2431,N_3088);
nor U8081 (N_8081,N_172,N_4814);
nand U8082 (N_8082,N_1294,N_1063);
or U8083 (N_8083,N_4296,N_409);
or U8084 (N_8084,N_738,N_1689);
nor U8085 (N_8085,N_3363,N_3540);
and U8086 (N_8086,N_1661,N_202);
nor U8087 (N_8087,N_3916,N_4574);
nor U8088 (N_8088,N_253,N_2079);
nor U8089 (N_8089,N_4723,N_3058);
or U8090 (N_8090,N_4612,N_1527);
or U8091 (N_8091,N_1994,N_1176);
nand U8092 (N_8092,N_1299,N_2127);
and U8093 (N_8093,N_2606,N_1680);
nor U8094 (N_8094,N_4877,N_4774);
and U8095 (N_8095,N_3407,N_3179);
xnor U8096 (N_8096,N_3227,N_2439);
xor U8097 (N_8097,N_3119,N_818);
nand U8098 (N_8098,N_2190,N_4299);
and U8099 (N_8099,N_1503,N_1947);
nand U8100 (N_8100,N_956,N_3391);
nor U8101 (N_8101,N_132,N_1853);
nand U8102 (N_8102,N_3317,N_3724);
and U8103 (N_8103,N_1562,N_4924);
nand U8104 (N_8104,N_3470,N_910);
and U8105 (N_8105,N_693,N_3686);
or U8106 (N_8106,N_2130,N_4788);
and U8107 (N_8107,N_1411,N_1932);
nor U8108 (N_8108,N_507,N_697);
xor U8109 (N_8109,N_581,N_3646);
and U8110 (N_8110,N_933,N_4324);
and U8111 (N_8111,N_4737,N_2446);
nor U8112 (N_8112,N_2989,N_1038);
and U8113 (N_8113,N_928,N_2896);
xnor U8114 (N_8114,N_3893,N_3965);
nor U8115 (N_8115,N_207,N_548);
xor U8116 (N_8116,N_3070,N_2179);
xnor U8117 (N_8117,N_1388,N_3235);
nand U8118 (N_8118,N_4618,N_3196);
and U8119 (N_8119,N_1076,N_266);
xnor U8120 (N_8120,N_382,N_2262);
nor U8121 (N_8121,N_1513,N_989);
and U8122 (N_8122,N_4145,N_4120);
and U8123 (N_8123,N_2822,N_2921);
or U8124 (N_8124,N_468,N_2915);
or U8125 (N_8125,N_4509,N_3778);
nand U8126 (N_8126,N_1842,N_4308);
and U8127 (N_8127,N_4045,N_3915);
nand U8128 (N_8128,N_4977,N_4208);
and U8129 (N_8129,N_3451,N_4653);
and U8130 (N_8130,N_463,N_1467);
and U8131 (N_8131,N_4489,N_4658);
xnor U8132 (N_8132,N_211,N_4341);
nor U8133 (N_8133,N_3343,N_2351);
xor U8134 (N_8134,N_2175,N_2);
xor U8135 (N_8135,N_2215,N_423);
and U8136 (N_8136,N_890,N_3229);
nor U8137 (N_8137,N_4684,N_938);
xor U8138 (N_8138,N_2043,N_3802);
xnor U8139 (N_8139,N_2028,N_1344);
nand U8140 (N_8140,N_2037,N_2055);
or U8141 (N_8141,N_3585,N_448);
and U8142 (N_8142,N_2381,N_4256);
xnor U8143 (N_8143,N_2284,N_2944);
and U8144 (N_8144,N_4224,N_3574);
or U8145 (N_8145,N_2651,N_2209);
and U8146 (N_8146,N_3863,N_2215);
and U8147 (N_8147,N_2933,N_1055);
nor U8148 (N_8148,N_119,N_4232);
nand U8149 (N_8149,N_2200,N_421);
nand U8150 (N_8150,N_1176,N_2167);
or U8151 (N_8151,N_2564,N_3707);
xnor U8152 (N_8152,N_225,N_2603);
nand U8153 (N_8153,N_1566,N_701);
nor U8154 (N_8154,N_1901,N_3490);
nand U8155 (N_8155,N_1132,N_3531);
nor U8156 (N_8156,N_3726,N_4797);
nor U8157 (N_8157,N_3829,N_2949);
and U8158 (N_8158,N_918,N_2317);
and U8159 (N_8159,N_1869,N_3075);
nand U8160 (N_8160,N_202,N_4206);
xor U8161 (N_8161,N_605,N_250);
xnor U8162 (N_8162,N_4715,N_2617);
or U8163 (N_8163,N_2216,N_645);
nand U8164 (N_8164,N_2418,N_4060);
nor U8165 (N_8165,N_1423,N_4189);
and U8166 (N_8166,N_4505,N_4363);
nor U8167 (N_8167,N_764,N_2780);
nor U8168 (N_8168,N_47,N_3675);
nor U8169 (N_8169,N_1037,N_179);
nand U8170 (N_8170,N_3386,N_3351);
or U8171 (N_8171,N_2247,N_197);
nand U8172 (N_8172,N_1125,N_1842);
or U8173 (N_8173,N_340,N_1721);
nand U8174 (N_8174,N_3676,N_1345);
nor U8175 (N_8175,N_997,N_3414);
or U8176 (N_8176,N_4251,N_3276);
or U8177 (N_8177,N_522,N_3091);
nand U8178 (N_8178,N_3498,N_38);
nor U8179 (N_8179,N_4445,N_560);
xor U8180 (N_8180,N_27,N_901);
nor U8181 (N_8181,N_3446,N_3920);
and U8182 (N_8182,N_1705,N_487);
nand U8183 (N_8183,N_1810,N_980);
nor U8184 (N_8184,N_627,N_4845);
and U8185 (N_8185,N_661,N_1727);
xnor U8186 (N_8186,N_2288,N_3349);
nand U8187 (N_8187,N_227,N_3109);
or U8188 (N_8188,N_4877,N_3669);
or U8189 (N_8189,N_2316,N_2872);
xnor U8190 (N_8190,N_4688,N_3989);
and U8191 (N_8191,N_2251,N_34);
nor U8192 (N_8192,N_2305,N_4885);
xor U8193 (N_8193,N_4179,N_807);
nand U8194 (N_8194,N_2164,N_2897);
and U8195 (N_8195,N_4963,N_4347);
xnor U8196 (N_8196,N_962,N_4662);
nand U8197 (N_8197,N_4086,N_1624);
nor U8198 (N_8198,N_4584,N_2548);
and U8199 (N_8199,N_2153,N_831);
nor U8200 (N_8200,N_4758,N_4087);
nor U8201 (N_8201,N_1242,N_4825);
xnor U8202 (N_8202,N_2854,N_3589);
and U8203 (N_8203,N_1355,N_3737);
xor U8204 (N_8204,N_4589,N_1033);
nor U8205 (N_8205,N_3208,N_901);
nor U8206 (N_8206,N_3036,N_162);
and U8207 (N_8207,N_1142,N_967);
nand U8208 (N_8208,N_679,N_2922);
nor U8209 (N_8209,N_4960,N_4778);
nor U8210 (N_8210,N_823,N_2758);
or U8211 (N_8211,N_2426,N_4546);
or U8212 (N_8212,N_3539,N_4721);
and U8213 (N_8213,N_2934,N_1392);
nor U8214 (N_8214,N_3163,N_3115);
or U8215 (N_8215,N_468,N_3074);
xor U8216 (N_8216,N_2282,N_111);
and U8217 (N_8217,N_4364,N_326);
and U8218 (N_8218,N_575,N_3832);
and U8219 (N_8219,N_3848,N_943);
and U8220 (N_8220,N_574,N_1287);
nor U8221 (N_8221,N_1338,N_3631);
or U8222 (N_8222,N_1384,N_584);
or U8223 (N_8223,N_1610,N_3593);
and U8224 (N_8224,N_3360,N_1753);
nor U8225 (N_8225,N_2975,N_1815);
nor U8226 (N_8226,N_2330,N_1216);
and U8227 (N_8227,N_4392,N_2049);
xor U8228 (N_8228,N_4105,N_2739);
nor U8229 (N_8229,N_4702,N_4121);
and U8230 (N_8230,N_2402,N_2546);
nor U8231 (N_8231,N_1179,N_763);
and U8232 (N_8232,N_4937,N_3289);
nor U8233 (N_8233,N_597,N_4394);
or U8234 (N_8234,N_2282,N_1683);
or U8235 (N_8235,N_3982,N_3258);
and U8236 (N_8236,N_749,N_3719);
or U8237 (N_8237,N_2859,N_3455);
and U8238 (N_8238,N_4576,N_4416);
xnor U8239 (N_8239,N_691,N_2589);
nor U8240 (N_8240,N_1288,N_1930);
nor U8241 (N_8241,N_1733,N_2680);
or U8242 (N_8242,N_4323,N_833);
xor U8243 (N_8243,N_295,N_2848);
nand U8244 (N_8244,N_740,N_1482);
and U8245 (N_8245,N_2371,N_134);
nor U8246 (N_8246,N_4918,N_2789);
or U8247 (N_8247,N_4577,N_3471);
or U8248 (N_8248,N_4832,N_2667);
or U8249 (N_8249,N_353,N_3240);
or U8250 (N_8250,N_2484,N_1575);
or U8251 (N_8251,N_1329,N_2732);
or U8252 (N_8252,N_1260,N_4813);
or U8253 (N_8253,N_1219,N_1678);
nand U8254 (N_8254,N_2930,N_10);
nor U8255 (N_8255,N_805,N_264);
nand U8256 (N_8256,N_3906,N_3745);
nor U8257 (N_8257,N_2520,N_4527);
nand U8258 (N_8258,N_312,N_3457);
nand U8259 (N_8259,N_3833,N_1173);
nand U8260 (N_8260,N_1618,N_329);
and U8261 (N_8261,N_4189,N_3347);
nor U8262 (N_8262,N_34,N_3940);
nor U8263 (N_8263,N_1701,N_4897);
xor U8264 (N_8264,N_4345,N_3441);
nand U8265 (N_8265,N_2931,N_730);
xnor U8266 (N_8266,N_4916,N_1150);
or U8267 (N_8267,N_4636,N_3282);
nor U8268 (N_8268,N_566,N_3549);
and U8269 (N_8269,N_2179,N_2399);
xnor U8270 (N_8270,N_2617,N_1310);
xor U8271 (N_8271,N_4861,N_4248);
or U8272 (N_8272,N_1843,N_2802);
or U8273 (N_8273,N_1188,N_8);
nor U8274 (N_8274,N_3194,N_3951);
nand U8275 (N_8275,N_3585,N_188);
nand U8276 (N_8276,N_1004,N_2829);
or U8277 (N_8277,N_831,N_2980);
or U8278 (N_8278,N_2061,N_1730);
xor U8279 (N_8279,N_4544,N_3034);
xor U8280 (N_8280,N_933,N_3039);
nor U8281 (N_8281,N_1378,N_3870);
nor U8282 (N_8282,N_2902,N_2323);
and U8283 (N_8283,N_1674,N_287);
nand U8284 (N_8284,N_1035,N_1791);
or U8285 (N_8285,N_3753,N_1945);
or U8286 (N_8286,N_4730,N_4082);
nor U8287 (N_8287,N_4544,N_2910);
nand U8288 (N_8288,N_761,N_2092);
nor U8289 (N_8289,N_1030,N_844);
and U8290 (N_8290,N_2769,N_472);
or U8291 (N_8291,N_2341,N_2686);
xor U8292 (N_8292,N_4321,N_584);
xnor U8293 (N_8293,N_2524,N_4105);
nor U8294 (N_8294,N_2659,N_3564);
or U8295 (N_8295,N_3966,N_3919);
nor U8296 (N_8296,N_4811,N_4267);
or U8297 (N_8297,N_3958,N_4917);
xor U8298 (N_8298,N_1919,N_3227);
nand U8299 (N_8299,N_1924,N_1999);
nand U8300 (N_8300,N_2877,N_2980);
and U8301 (N_8301,N_1906,N_4475);
xor U8302 (N_8302,N_4287,N_286);
nor U8303 (N_8303,N_1442,N_2691);
or U8304 (N_8304,N_2883,N_2733);
and U8305 (N_8305,N_4474,N_2773);
nand U8306 (N_8306,N_2744,N_886);
or U8307 (N_8307,N_3599,N_884);
or U8308 (N_8308,N_1107,N_19);
nor U8309 (N_8309,N_1209,N_880);
and U8310 (N_8310,N_4586,N_355);
or U8311 (N_8311,N_556,N_1230);
nand U8312 (N_8312,N_2624,N_910);
xor U8313 (N_8313,N_2787,N_2287);
and U8314 (N_8314,N_1883,N_1962);
xnor U8315 (N_8315,N_4082,N_3161);
nand U8316 (N_8316,N_4990,N_2685);
and U8317 (N_8317,N_2410,N_4731);
xnor U8318 (N_8318,N_2417,N_2611);
nor U8319 (N_8319,N_1339,N_2761);
nor U8320 (N_8320,N_3063,N_4558);
xor U8321 (N_8321,N_4119,N_132);
or U8322 (N_8322,N_1551,N_3652);
and U8323 (N_8323,N_1511,N_4812);
xnor U8324 (N_8324,N_1816,N_2172);
nand U8325 (N_8325,N_1732,N_3171);
nor U8326 (N_8326,N_601,N_4506);
nand U8327 (N_8327,N_2258,N_3698);
xnor U8328 (N_8328,N_3607,N_2046);
or U8329 (N_8329,N_715,N_4313);
nor U8330 (N_8330,N_606,N_2047);
and U8331 (N_8331,N_1085,N_2205);
and U8332 (N_8332,N_3447,N_3168);
xnor U8333 (N_8333,N_4275,N_1397);
nand U8334 (N_8334,N_3972,N_4315);
xor U8335 (N_8335,N_4594,N_3250);
and U8336 (N_8336,N_3168,N_1035);
or U8337 (N_8337,N_4470,N_3963);
and U8338 (N_8338,N_3220,N_2976);
xnor U8339 (N_8339,N_432,N_4520);
nor U8340 (N_8340,N_656,N_4632);
or U8341 (N_8341,N_4427,N_902);
nor U8342 (N_8342,N_2213,N_374);
nand U8343 (N_8343,N_3161,N_490);
nor U8344 (N_8344,N_3414,N_441);
or U8345 (N_8345,N_989,N_3078);
or U8346 (N_8346,N_3484,N_4807);
xnor U8347 (N_8347,N_2590,N_306);
nand U8348 (N_8348,N_4269,N_2239);
xor U8349 (N_8349,N_3208,N_534);
xnor U8350 (N_8350,N_4111,N_2898);
or U8351 (N_8351,N_1552,N_2450);
or U8352 (N_8352,N_3642,N_3790);
and U8353 (N_8353,N_135,N_2581);
and U8354 (N_8354,N_3637,N_429);
nor U8355 (N_8355,N_1626,N_3571);
nor U8356 (N_8356,N_218,N_1319);
xnor U8357 (N_8357,N_1738,N_3463);
nor U8358 (N_8358,N_198,N_2621);
or U8359 (N_8359,N_4815,N_3131);
xnor U8360 (N_8360,N_3469,N_2258);
xnor U8361 (N_8361,N_3511,N_2054);
nand U8362 (N_8362,N_3512,N_3746);
xnor U8363 (N_8363,N_4298,N_2912);
nand U8364 (N_8364,N_799,N_4083);
xnor U8365 (N_8365,N_4360,N_3153);
nand U8366 (N_8366,N_952,N_1539);
nand U8367 (N_8367,N_2237,N_2696);
and U8368 (N_8368,N_1220,N_3100);
nand U8369 (N_8369,N_1346,N_2095);
or U8370 (N_8370,N_4374,N_690);
and U8371 (N_8371,N_4018,N_4921);
nand U8372 (N_8372,N_1678,N_821);
nor U8373 (N_8373,N_880,N_2236);
nand U8374 (N_8374,N_3309,N_3970);
and U8375 (N_8375,N_582,N_635);
nand U8376 (N_8376,N_526,N_3875);
and U8377 (N_8377,N_1366,N_4546);
nand U8378 (N_8378,N_3740,N_1102);
nor U8379 (N_8379,N_2488,N_3111);
xnor U8380 (N_8380,N_3033,N_4045);
nand U8381 (N_8381,N_371,N_4460);
and U8382 (N_8382,N_4370,N_1323);
xnor U8383 (N_8383,N_4538,N_3522);
and U8384 (N_8384,N_632,N_3121);
nor U8385 (N_8385,N_1420,N_974);
nand U8386 (N_8386,N_1527,N_2820);
and U8387 (N_8387,N_2041,N_1081);
or U8388 (N_8388,N_173,N_4252);
nand U8389 (N_8389,N_2904,N_220);
nor U8390 (N_8390,N_1504,N_2356);
or U8391 (N_8391,N_4867,N_3097);
nor U8392 (N_8392,N_4657,N_1305);
and U8393 (N_8393,N_1606,N_2340);
nor U8394 (N_8394,N_1876,N_183);
and U8395 (N_8395,N_4175,N_2308);
nor U8396 (N_8396,N_2611,N_4601);
xnor U8397 (N_8397,N_2356,N_4625);
xor U8398 (N_8398,N_3671,N_689);
and U8399 (N_8399,N_1360,N_465);
nor U8400 (N_8400,N_4503,N_1386);
xor U8401 (N_8401,N_1701,N_2431);
or U8402 (N_8402,N_3150,N_3633);
and U8403 (N_8403,N_2400,N_564);
xnor U8404 (N_8404,N_4381,N_2813);
or U8405 (N_8405,N_3382,N_1945);
nand U8406 (N_8406,N_3872,N_2528);
xnor U8407 (N_8407,N_1922,N_4453);
nor U8408 (N_8408,N_244,N_1534);
and U8409 (N_8409,N_1334,N_1532);
or U8410 (N_8410,N_1621,N_283);
nand U8411 (N_8411,N_1690,N_862);
nor U8412 (N_8412,N_1933,N_3127);
and U8413 (N_8413,N_2203,N_2536);
and U8414 (N_8414,N_3296,N_707);
or U8415 (N_8415,N_4549,N_4785);
nand U8416 (N_8416,N_4596,N_833);
nand U8417 (N_8417,N_509,N_2974);
and U8418 (N_8418,N_2664,N_4607);
and U8419 (N_8419,N_325,N_2795);
nand U8420 (N_8420,N_2388,N_775);
or U8421 (N_8421,N_2524,N_4677);
and U8422 (N_8422,N_3427,N_2966);
and U8423 (N_8423,N_2088,N_4458);
nor U8424 (N_8424,N_4245,N_2994);
and U8425 (N_8425,N_3653,N_2349);
nor U8426 (N_8426,N_4073,N_4720);
and U8427 (N_8427,N_1101,N_3480);
nand U8428 (N_8428,N_1091,N_504);
nand U8429 (N_8429,N_4188,N_4094);
nor U8430 (N_8430,N_2014,N_3218);
nor U8431 (N_8431,N_197,N_3883);
nand U8432 (N_8432,N_1469,N_1426);
nand U8433 (N_8433,N_3955,N_2753);
xor U8434 (N_8434,N_1504,N_870);
xor U8435 (N_8435,N_3710,N_4446);
nor U8436 (N_8436,N_778,N_1163);
nor U8437 (N_8437,N_2280,N_4455);
nor U8438 (N_8438,N_388,N_757);
xor U8439 (N_8439,N_3921,N_740);
xor U8440 (N_8440,N_1884,N_1819);
nor U8441 (N_8441,N_4416,N_170);
or U8442 (N_8442,N_1027,N_1232);
nand U8443 (N_8443,N_1923,N_1193);
or U8444 (N_8444,N_4235,N_3039);
and U8445 (N_8445,N_2430,N_107);
nand U8446 (N_8446,N_4806,N_3526);
and U8447 (N_8447,N_4581,N_2091);
nor U8448 (N_8448,N_1266,N_2659);
nor U8449 (N_8449,N_516,N_703);
xnor U8450 (N_8450,N_1485,N_3648);
nand U8451 (N_8451,N_1118,N_978);
nand U8452 (N_8452,N_386,N_1359);
nand U8453 (N_8453,N_4369,N_754);
and U8454 (N_8454,N_4308,N_3966);
nand U8455 (N_8455,N_3316,N_2907);
and U8456 (N_8456,N_1245,N_2687);
nor U8457 (N_8457,N_409,N_2002);
nand U8458 (N_8458,N_4739,N_10);
or U8459 (N_8459,N_2366,N_2037);
or U8460 (N_8460,N_204,N_778);
xnor U8461 (N_8461,N_4509,N_302);
nor U8462 (N_8462,N_1877,N_3125);
nor U8463 (N_8463,N_2652,N_1003);
or U8464 (N_8464,N_1425,N_3296);
nor U8465 (N_8465,N_4283,N_2740);
nor U8466 (N_8466,N_1249,N_1665);
nor U8467 (N_8467,N_70,N_4733);
or U8468 (N_8468,N_3429,N_1348);
xnor U8469 (N_8469,N_2814,N_835);
nand U8470 (N_8470,N_2780,N_3654);
and U8471 (N_8471,N_3238,N_2423);
nand U8472 (N_8472,N_1209,N_4986);
nor U8473 (N_8473,N_2493,N_4189);
nor U8474 (N_8474,N_2711,N_729);
nand U8475 (N_8475,N_844,N_4406);
or U8476 (N_8476,N_1010,N_3929);
nand U8477 (N_8477,N_1862,N_3382);
xor U8478 (N_8478,N_2570,N_3520);
and U8479 (N_8479,N_2277,N_339);
and U8480 (N_8480,N_1809,N_4762);
and U8481 (N_8481,N_1764,N_4284);
and U8482 (N_8482,N_2854,N_3839);
nand U8483 (N_8483,N_4513,N_2274);
nand U8484 (N_8484,N_2692,N_2850);
nor U8485 (N_8485,N_3068,N_1855);
and U8486 (N_8486,N_3463,N_4318);
and U8487 (N_8487,N_993,N_1857);
and U8488 (N_8488,N_122,N_4661);
nand U8489 (N_8489,N_3021,N_1735);
xnor U8490 (N_8490,N_1180,N_1527);
xnor U8491 (N_8491,N_3593,N_496);
nand U8492 (N_8492,N_828,N_1552);
xor U8493 (N_8493,N_4039,N_2370);
nor U8494 (N_8494,N_3726,N_1916);
nand U8495 (N_8495,N_2118,N_1466);
nor U8496 (N_8496,N_1846,N_1254);
nor U8497 (N_8497,N_582,N_4289);
or U8498 (N_8498,N_4264,N_897);
and U8499 (N_8499,N_4581,N_4753);
nand U8500 (N_8500,N_474,N_1343);
xnor U8501 (N_8501,N_1689,N_4596);
nor U8502 (N_8502,N_1902,N_2442);
or U8503 (N_8503,N_4661,N_597);
nand U8504 (N_8504,N_2539,N_1333);
xnor U8505 (N_8505,N_62,N_4632);
or U8506 (N_8506,N_4634,N_3787);
and U8507 (N_8507,N_1182,N_1665);
xnor U8508 (N_8508,N_1963,N_100);
nand U8509 (N_8509,N_853,N_2827);
nor U8510 (N_8510,N_4122,N_216);
xor U8511 (N_8511,N_4863,N_2272);
nand U8512 (N_8512,N_607,N_23);
xor U8513 (N_8513,N_3875,N_4336);
and U8514 (N_8514,N_4704,N_1081);
xor U8515 (N_8515,N_4286,N_4524);
nor U8516 (N_8516,N_1345,N_3404);
nand U8517 (N_8517,N_4254,N_3606);
or U8518 (N_8518,N_3448,N_420);
nor U8519 (N_8519,N_3579,N_2259);
nor U8520 (N_8520,N_4651,N_3148);
nand U8521 (N_8521,N_4896,N_3116);
and U8522 (N_8522,N_2422,N_844);
and U8523 (N_8523,N_4457,N_4091);
xnor U8524 (N_8524,N_3477,N_2110);
or U8525 (N_8525,N_559,N_1599);
and U8526 (N_8526,N_2381,N_2768);
or U8527 (N_8527,N_3556,N_3359);
and U8528 (N_8528,N_2957,N_3766);
nand U8529 (N_8529,N_2364,N_3216);
nor U8530 (N_8530,N_2073,N_943);
nand U8531 (N_8531,N_1006,N_1888);
or U8532 (N_8532,N_1782,N_4872);
and U8533 (N_8533,N_650,N_2776);
nor U8534 (N_8534,N_3999,N_3058);
nor U8535 (N_8535,N_1925,N_854);
nand U8536 (N_8536,N_4842,N_3805);
or U8537 (N_8537,N_1168,N_1811);
or U8538 (N_8538,N_2610,N_1090);
or U8539 (N_8539,N_4983,N_1617);
nand U8540 (N_8540,N_1287,N_2091);
or U8541 (N_8541,N_1524,N_1560);
nor U8542 (N_8542,N_3547,N_564);
xnor U8543 (N_8543,N_2405,N_3231);
xnor U8544 (N_8544,N_2696,N_4267);
xor U8545 (N_8545,N_4230,N_1440);
or U8546 (N_8546,N_3575,N_1308);
nand U8547 (N_8547,N_2676,N_905);
or U8548 (N_8548,N_2204,N_170);
nand U8549 (N_8549,N_2921,N_4416);
xnor U8550 (N_8550,N_1388,N_2609);
nor U8551 (N_8551,N_3881,N_4837);
xnor U8552 (N_8552,N_1870,N_768);
nor U8553 (N_8553,N_477,N_4942);
nor U8554 (N_8554,N_2248,N_4116);
or U8555 (N_8555,N_1629,N_3333);
or U8556 (N_8556,N_647,N_4832);
and U8557 (N_8557,N_2125,N_894);
or U8558 (N_8558,N_2425,N_2687);
nor U8559 (N_8559,N_1712,N_1714);
nand U8560 (N_8560,N_4645,N_1102);
and U8561 (N_8561,N_2451,N_4102);
xnor U8562 (N_8562,N_3168,N_2738);
nor U8563 (N_8563,N_3262,N_2148);
xor U8564 (N_8564,N_1755,N_924);
nor U8565 (N_8565,N_1739,N_4313);
xnor U8566 (N_8566,N_1398,N_3331);
nor U8567 (N_8567,N_2876,N_4023);
and U8568 (N_8568,N_546,N_3198);
nor U8569 (N_8569,N_2178,N_1586);
xor U8570 (N_8570,N_4721,N_3765);
nor U8571 (N_8571,N_119,N_1098);
and U8572 (N_8572,N_4314,N_2440);
nand U8573 (N_8573,N_2417,N_2718);
nand U8574 (N_8574,N_18,N_3449);
and U8575 (N_8575,N_1782,N_2670);
nor U8576 (N_8576,N_4423,N_1358);
nand U8577 (N_8577,N_4770,N_3629);
nor U8578 (N_8578,N_2953,N_3915);
or U8579 (N_8579,N_4523,N_1953);
and U8580 (N_8580,N_4586,N_1510);
xnor U8581 (N_8581,N_2299,N_3385);
or U8582 (N_8582,N_1969,N_2812);
xor U8583 (N_8583,N_533,N_3105);
or U8584 (N_8584,N_3649,N_1229);
or U8585 (N_8585,N_4230,N_2392);
nor U8586 (N_8586,N_1820,N_1359);
nor U8587 (N_8587,N_3016,N_3115);
or U8588 (N_8588,N_3899,N_4199);
or U8589 (N_8589,N_3402,N_252);
or U8590 (N_8590,N_3725,N_2021);
or U8591 (N_8591,N_874,N_663);
or U8592 (N_8592,N_701,N_192);
nor U8593 (N_8593,N_435,N_1458);
xnor U8594 (N_8594,N_1171,N_2343);
xor U8595 (N_8595,N_3759,N_2333);
and U8596 (N_8596,N_3860,N_3611);
and U8597 (N_8597,N_4011,N_4568);
nand U8598 (N_8598,N_3713,N_3436);
nor U8599 (N_8599,N_2748,N_4817);
xnor U8600 (N_8600,N_1856,N_114);
nor U8601 (N_8601,N_4670,N_3449);
nor U8602 (N_8602,N_2954,N_1270);
nand U8603 (N_8603,N_3159,N_1937);
and U8604 (N_8604,N_1085,N_4476);
nor U8605 (N_8605,N_1056,N_4395);
xor U8606 (N_8606,N_1658,N_3499);
or U8607 (N_8607,N_4120,N_4812);
nor U8608 (N_8608,N_2326,N_422);
and U8609 (N_8609,N_3376,N_2830);
xnor U8610 (N_8610,N_4705,N_3413);
nor U8611 (N_8611,N_3762,N_2916);
or U8612 (N_8612,N_4972,N_4346);
xor U8613 (N_8613,N_3385,N_7);
nor U8614 (N_8614,N_3307,N_3398);
xnor U8615 (N_8615,N_952,N_2780);
xnor U8616 (N_8616,N_1591,N_4237);
xnor U8617 (N_8617,N_904,N_4603);
nand U8618 (N_8618,N_1714,N_4999);
nand U8619 (N_8619,N_3787,N_3211);
xor U8620 (N_8620,N_4277,N_486);
and U8621 (N_8621,N_4945,N_857);
nand U8622 (N_8622,N_3991,N_2);
nor U8623 (N_8623,N_1888,N_2122);
nand U8624 (N_8624,N_2625,N_3172);
or U8625 (N_8625,N_19,N_2724);
nand U8626 (N_8626,N_1491,N_2898);
and U8627 (N_8627,N_2685,N_1373);
nor U8628 (N_8628,N_623,N_2311);
or U8629 (N_8629,N_1222,N_290);
xnor U8630 (N_8630,N_440,N_4232);
nand U8631 (N_8631,N_4147,N_3310);
nand U8632 (N_8632,N_1646,N_3907);
or U8633 (N_8633,N_4931,N_1529);
or U8634 (N_8634,N_2885,N_731);
xor U8635 (N_8635,N_2075,N_1805);
xor U8636 (N_8636,N_2741,N_3840);
and U8637 (N_8637,N_1878,N_1839);
and U8638 (N_8638,N_3040,N_3224);
nor U8639 (N_8639,N_2172,N_3851);
or U8640 (N_8640,N_3162,N_3549);
nor U8641 (N_8641,N_4032,N_4897);
or U8642 (N_8642,N_107,N_3276);
or U8643 (N_8643,N_4260,N_565);
nand U8644 (N_8644,N_1396,N_626);
or U8645 (N_8645,N_1805,N_2280);
nor U8646 (N_8646,N_609,N_1592);
or U8647 (N_8647,N_4464,N_1668);
and U8648 (N_8648,N_4529,N_416);
and U8649 (N_8649,N_4858,N_2682);
xnor U8650 (N_8650,N_4173,N_3219);
nor U8651 (N_8651,N_2675,N_1847);
xnor U8652 (N_8652,N_4875,N_233);
or U8653 (N_8653,N_2167,N_4062);
nor U8654 (N_8654,N_4370,N_1974);
or U8655 (N_8655,N_2824,N_4724);
and U8656 (N_8656,N_3042,N_4303);
xnor U8657 (N_8657,N_3645,N_2970);
nand U8658 (N_8658,N_4471,N_838);
xor U8659 (N_8659,N_4393,N_1495);
and U8660 (N_8660,N_29,N_2016);
nor U8661 (N_8661,N_233,N_4930);
and U8662 (N_8662,N_3722,N_4815);
or U8663 (N_8663,N_4868,N_4489);
nand U8664 (N_8664,N_4201,N_3036);
or U8665 (N_8665,N_3514,N_1498);
or U8666 (N_8666,N_4899,N_3707);
nand U8667 (N_8667,N_3206,N_96);
or U8668 (N_8668,N_2471,N_4403);
or U8669 (N_8669,N_2125,N_4251);
nand U8670 (N_8670,N_3159,N_481);
nand U8671 (N_8671,N_2983,N_2819);
nand U8672 (N_8672,N_1723,N_112);
xnor U8673 (N_8673,N_1920,N_3534);
xor U8674 (N_8674,N_2928,N_4223);
xnor U8675 (N_8675,N_135,N_4574);
and U8676 (N_8676,N_4068,N_4931);
nand U8677 (N_8677,N_4402,N_4436);
or U8678 (N_8678,N_875,N_2336);
or U8679 (N_8679,N_2461,N_955);
nand U8680 (N_8680,N_2111,N_1477);
or U8681 (N_8681,N_1819,N_2145);
nor U8682 (N_8682,N_3959,N_3224);
or U8683 (N_8683,N_2566,N_4472);
xor U8684 (N_8684,N_4234,N_2630);
or U8685 (N_8685,N_4983,N_1998);
nand U8686 (N_8686,N_4765,N_3815);
xnor U8687 (N_8687,N_1207,N_2257);
xor U8688 (N_8688,N_3725,N_367);
or U8689 (N_8689,N_1409,N_1109);
nand U8690 (N_8690,N_3592,N_1408);
nand U8691 (N_8691,N_2685,N_336);
nor U8692 (N_8692,N_4691,N_406);
and U8693 (N_8693,N_1202,N_3495);
or U8694 (N_8694,N_4064,N_4566);
or U8695 (N_8695,N_3532,N_1935);
nand U8696 (N_8696,N_481,N_3000);
nor U8697 (N_8697,N_3307,N_4974);
nor U8698 (N_8698,N_4578,N_139);
nand U8699 (N_8699,N_344,N_394);
and U8700 (N_8700,N_951,N_3810);
and U8701 (N_8701,N_4502,N_4430);
and U8702 (N_8702,N_4449,N_3896);
and U8703 (N_8703,N_1615,N_3703);
nor U8704 (N_8704,N_3299,N_2170);
nand U8705 (N_8705,N_2978,N_1016);
and U8706 (N_8706,N_3314,N_1689);
nand U8707 (N_8707,N_4454,N_813);
nor U8708 (N_8708,N_2822,N_563);
xnor U8709 (N_8709,N_4124,N_1050);
xor U8710 (N_8710,N_2468,N_1088);
nor U8711 (N_8711,N_2405,N_3668);
nand U8712 (N_8712,N_3265,N_2604);
nand U8713 (N_8713,N_4777,N_3210);
or U8714 (N_8714,N_3969,N_2108);
and U8715 (N_8715,N_2720,N_2771);
xnor U8716 (N_8716,N_3608,N_566);
nand U8717 (N_8717,N_794,N_1299);
nor U8718 (N_8718,N_1390,N_746);
or U8719 (N_8719,N_4308,N_27);
or U8720 (N_8720,N_246,N_2373);
xnor U8721 (N_8721,N_2795,N_4840);
xnor U8722 (N_8722,N_3888,N_4087);
or U8723 (N_8723,N_689,N_1222);
nand U8724 (N_8724,N_340,N_4229);
nand U8725 (N_8725,N_3356,N_1950);
nand U8726 (N_8726,N_2799,N_462);
nor U8727 (N_8727,N_811,N_4140);
nand U8728 (N_8728,N_2507,N_2796);
and U8729 (N_8729,N_2235,N_4571);
and U8730 (N_8730,N_3617,N_2667);
xnor U8731 (N_8731,N_4993,N_3993);
and U8732 (N_8732,N_1497,N_2969);
xor U8733 (N_8733,N_3338,N_4734);
or U8734 (N_8734,N_3742,N_3297);
or U8735 (N_8735,N_4394,N_4942);
or U8736 (N_8736,N_2132,N_4333);
and U8737 (N_8737,N_4630,N_3326);
xor U8738 (N_8738,N_2342,N_3120);
or U8739 (N_8739,N_1432,N_4644);
and U8740 (N_8740,N_3939,N_1511);
nand U8741 (N_8741,N_2728,N_479);
or U8742 (N_8742,N_4496,N_1988);
nand U8743 (N_8743,N_2077,N_1177);
and U8744 (N_8744,N_4504,N_1179);
nand U8745 (N_8745,N_215,N_772);
nand U8746 (N_8746,N_3952,N_1061);
xnor U8747 (N_8747,N_1631,N_2535);
nand U8748 (N_8748,N_1852,N_4998);
and U8749 (N_8749,N_2193,N_1619);
nor U8750 (N_8750,N_2795,N_3919);
xor U8751 (N_8751,N_408,N_2967);
xnor U8752 (N_8752,N_380,N_126);
and U8753 (N_8753,N_324,N_1540);
and U8754 (N_8754,N_1885,N_793);
nor U8755 (N_8755,N_4058,N_144);
xor U8756 (N_8756,N_4153,N_4214);
nor U8757 (N_8757,N_1843,N_4790);
xor U8758 (N_8758,N_4509,N_2197);
nor U8759 (N_8759,N_4055,N_1483);
nor U8760 (N_8760,N_806,N_3190);
and U8761 (N_8761,N_497,N_1492);
xor U8762 (N_8762,N_3400,N_1110);
nor U8763 (N_8763,N_4802,N_3041);
nor U8764 (N_8764,N_3292,N_1425);
nand U8765 (N_8765,N_4317,N_2693);
nor U8766 (N_8766,N_97,N_4222);
nor U8767 (N_8767,N_2607,N_1468);
nor U8768 (N_8768,N_2040,N_4192);
and U8769 (N_8769,N_2502,N_1008);
and U8770 (N_8770,N_2621,N_2211);
xor U8771 (N_8771,N_1685,N_2762);
xnor U8772 (N_8772,N_765,N_3202);
nor U8773 (N_8773,N_3597,N_4845);
or U8774 (N_8774,N_3915,N_1281);
nand U8775 (N_8775,N_2121,N_863);
nor U8776 (N_8776,N_3533,N_1961);
xor U8777 (N_8777,N_2623,N_3184);
or U8778 (N_8778,N_1322,N_2708);
nand U8779 (N_8779,N_2687,N_1126);
nor U8780 (N_8780,N_1281,N_1250);
xor U8781 (N_8781,N_1276,N_628);
nor U8782 (N_8782,N_3289,N_848);
nor U8783 (N_8783,N_3421,N_119);
nor U8784 (N_8784,N_3064,N_4816);
or U8785 (N_8785,N_3235,N_2651);
nand U8786 (N_8786,N_1080,N_3278);
xor U8787 (N_8787,N_3997,N_24);
nand U8788 (N_8788,N_4728,N_853);
nand U8789 (N_8789,N_3702,N_2589);
xnor U8790 (N_8790,N_4213,N_3213);
and U8791 (N_8791,N_706,N_4409);
nor U8792 (N_8792,N_3932,N_1824);
xor U8793 (N_8793,N_3690,N_2139);
nand U8794 (N_8794,N_4131,N_1259);
nand U8795 (N_8795,N_777,N_3843);
nand U8796 (N_8796,N_1688,N_3158);
xnor U8797 (N_8797,N_2118,N_2590);
nor U8798 (N_8798,N_1111,N_748);
nand U8799 (N_8799,N_4187,N_963);
xor U8800 (N_8800,N_1989,N_2023);
nand U8801 (N_8801,N_2502,N_1448);
xor U8802 (N_8802,N_285,N_3089);
and U8803 (N_8803,N_3557,N_2005);
or U8804 (N_8804,N_666,N_2628);
nand U8805 (N_8805,N_4487,N_1077);
and U8806 (N_8806,N_2776,N_3769);
nor U8807 (N_8807,N_3798,N_1993);
and U8808 (N_8808,N_988,N_2237);
xor U8809 (N_8809,N_2979,N_236);
or U8810 (N_8810,N_979,N_1215);
nand U8811 (N_8811,N_734,N_2831);
nor U8812 (N_8812,N_2349,N_4001);
nor U8813 (N_8813,N_117,N_2009);
nor U8814 (N_8814,N_1932,N_944);
nor U8815 (N_8815,N_1850,N_3899);
or U8816 (N_8816,N_4279,N_873);
nand U8817 (N_8817,N_1231,N_1065);
or U8818 (N_8818,N_3817,N_366);
or U8819 (N_8819,N_4562,N_2025);
and U8820 (N_8820,N_241,N_4757);
nor U8821 (N_8821,N_4348,N_1766);
or U8822 (N_8822,N_4747,N_255);
and U8823 (N_8823,N_1600,N_4651);
or U8824 (N_8824,N_727,N_4073);
nand U8825 (N_8825,N_1153,N_2504);
and U8826 (N_8826,N_2482,N_778);
nand U8827 (N_8827,N_1884,N_3816);
nand U8828 (N_8828,N_2257,N_130);
or U8829 (N_8829,N_4486,N_265);
nor U8830 (N_8830,N_417,N_3116);
or U8831 (N_8831,N_353,N_1303);
nor U8832 (N_8832,N_816,N_1078);
and U8833 (N_8833,N_1582,N_4900);
nor U8834 (N_8834,N_1681,N_4331);
or U8835 (N_8835,N_1684,N_2385);
xor U8836 (N_8836,N_718,N_2218);
nor U8837 (N_8837,N_2374,N_2204);
nor U8838 (N_8838,N_2714,N_3865);
nor U8839 (N_8839,N_1160,N_4260);
xor U8840 (N_8840,N_650,N_1934);
xnor U8841 (N_8841,N_4284,N_4050);
xor U8842 (N_8842,N_1398,N_4149);
or U8843 (N_8843,N_1531,N_2363);
xnor U8844 (N_8844,N_3048,N_830);
nand U8845 (N_8845,N_2721,N_130);
and U8846 (N_8846,N_4672,N_308);
or U8847 (N_8847,N_76,N_2723);
nor U8848 (N_8848,N_3376,N_126);
and U8849 (N_8849,N_4483,N_4421);
nor U8850 (N_8850,N_416,N_607);
and U8851 (N_8851,N_4366,N_1793);
nor U8852 (N_8852,N_2877,N_4457);
nand U8853 (N_8853,N_3511,N_1413);
or U8854 (N_8854,N_2857,N_3080);
or U8855 (N_8855,N_1556,N_712);
nor U8856 (N_8856,N_216,N_4270);
and U8857 (N_8857,N_4733,N_3282);
or U8858 (N_8858,N_7,N_4793);
or U8859 (N_8859,N_1957,N_3404);
nand U8860 (N_8860,N_2010,N_3762);
and U8861 (N_8861,N_2446,N_2942);
and U8862 (N_8862,N_3629,N_1965);
xnor U8863 (N_8863,N_2114,N_3497);
nand U8864 (N_8864,N_4057,N_643);
or U8865 (N_8865,N_4097,N_3106);
and U8866 (N_8866,N_3587,N_2736);
nand U8867 (N_8867,N_4251,N_3738);
nand U8868 (N_8868,N_1075,N_3024);
nand U8869 (N_8869,N_4092,N_1574);
and U8870 (N_8870,N_37,N_696);
or U8871 (N_8871,N_326,N_2761);
nor U8872 (N_8872,N_3488,N_1601);
or U8873 (N_8873,N_2906,N_3176);
or U8874 (N_8874,N_3775,N_3702);
nor U8875 (N_8875,N_4914,N_330);
and U8876 (N_8876,N_4909,N_4688);
or U8877 (N_8877,N_685,N_112);
nand U8878 (N_8878,N_2071,N_1031);
and U8879 (N_8879,N_253,N_2623);
xnor U8880 (N_8880,N_1676,N_4471);
or U8881 (N_8881,N_4338,N_2356);
nor U8882 (N_8882,N_1631,N_1404);
xnor U8883 (N_8883,N_2356,N_3628);
and U8884 (N_8884,N_3640,N_4308);
or U8885 (N_8885,N_1391,N_2993);
and U8886 (N_8886,N_2475,N_4646);
xnor U8887 (N_8887,N_2210,N_1886);
nand U8888 (N_8888,N_4616,N_2607);
or U8889 (N_8889,N_741,N_3312);
nor U8890 (N_8890,N_1075,N_2222);
nor U8891 (N_8891,N_2674,N_3543);
nor U8892 (N_8892,N_2440,N_638);
xnor U8893 (N_8893,N_1332,N_2477);
nand U8894 (N_8894,N_783,N_4760);
xor U8895 (N_8895,N_3664,N_2460);
and U8896 (N_8896,N_236,N_3196);
and U8897 (N_8897,N_4272,N_484);
xor U8898 (N_8898,N_739,N_624);
and U8899 (N_8899,N_1885,N_4072);
nand U8900 (N_8900,N_3653,N_4635);
nor U8901 (N_8901,N_2790,N_3673);
nor U8902 (N_8902,N_463,N_1734);
nor U8903 (N_8903,N_527,N_3469);
and U8904 (N_8904,N_4603,N_1332);
nor U8905 (N_8905,N_2350,N_3430);
nand U8906 (N_8906,N_3140,N_4986);
and U8907 (N_8907,N_4379,N_241);
nor U8908 (N_8908,N_3038,N_2111);
xnor U8909 (N_8909,N_3684,N_531);
and U8910 (N_8910,N_2317,N_3193);
nand U8911 (N_8911,N_4840,N_1216);
or U8912 (N_8912,N_2163,N_3549);
and U8913 (N_8913,N_3256,N_4568);
xnor U8914 (N_8914,N_2936,N_3153);
xor U8915 (N_8915,N_444,N_445);
and U8916 (N_8916,N_1706,N_3508);
or U8917 (N_8917,N_2812,N_1327);
and U8918 (N_8918,N_1554,N_4918);
and U8919 (N_8919,N_4193,N_270);
nand U8920 (N_8920,N_3299,N_1563);
nor U8921 (N_8921,N_1508,N_1158);
nor U8922 (N_8922,N_3909,N_20);
and U8923 (N_8923,N_4674,N_4134);
nor U8924 (N_8924,N_4089,N_4940);
nand U8925 (N_8925,N_1815,N_115);
and U8926 (N_8926,N_3739,N_1657);
nor U8927 (N_8927,N_3614,N_1225);
or U8928 (N_8928,N_2381,N_2103);
nor U8929 (N_8929,N_4861,N_993);
nand U8930 (N_8930,N_1865,N_670);
nand U8931 (N_8931,N_1137,N_1828);
or U8932 (N_8932,N_2362,N_4036);
nand U8933 (N_8933,N_3021,N_2002);
xnor U8934 (N_8934,N_4073,N_1697);
or U8935 (N_8935,N_3930,N_3120);
nor U8936 (N_8936,N_1918,N_1103);
or U8937 (N_8937,N_1536,N_3175);
or U8938 (N_8938,N_1539,N_3765);
nor U8939 (N_8939,N_4096,N_2243);
or U8940 (N_8940,N_4407,N_2605);
or U8941 (N_8941,N_4138,N_1829);
xor U8942 (N_8942,N_2024,N_3172);
nand U8943 (N_8943,N_4450,N_4730);
and U8944 (N_8944,N_482,N_2494);
nand U8945 (N_8945,N_2061,N_4784);
or U8946 (N_8946,N_3457,N_4562);
and U8947 (N_8947,N_2803,N_3529);
and U8948 (N_8948,N_3416,N_4701);
and U8949 (N_8949,N_436,N_900);
nor U8950 (N_8950,N_788,N_203);
nor U8951 (N_8951,N_3943,N_3066);
nand U8952 (N_8952,N_394,N_2042);
nand U8953 (N_8953,N_411,N_3087);
and U8954 (N_8954,N_2265,N_220);
xor U8955 (N_8955,N_4394,N_3096);
nor U8956 (N_8956,N_266,N_3030);
nand U8957 (N_8957,N_1690,N_4254);
xnor U8958 (N_8958,N_2216,N_87);
or U8959 (N_8959,N_1043,N_4794);
nor U8960 (N_8960,N_4381,N_4355);
nor U8961 (N_8961,N_4501,N_1488);
and U8962 (N_8962,N_3612,N_1121);
and U8963 (N_8963,N_57,N_1062);
nor U8964 (N_8964,N_1372,N_412);
and U8965 (N_8965,N_3316,N_308);
or U8966 (N_8966,N_3429,N_2845);
nand U8967 (N_8967,N_4889,N_2755);
and U8968 (N_8968,N_3947,N_1875);
nand U8969 (N_8969,N_2971,N_2577);
or U8970 (N_8970,N_1953,N_797);
nor U8971 (N_8971,N_2874,N_3143);
nor U8972 (N_8972,N_1495,N_518);
or U8973 (N_8973,N_1908,N_1339);
xor U8974 (N_8974,N_4625,N_566);
and U8975 (N_8975,N_1965,N_4904);
and U8976 (N_8976,N_487,N_4419);
nor U8977 (N_8977,N_711,N_3833);
and U8978 (N_8978,N_207,N_2769);
and U8979 (N_8979,N_1020,N_2981);
or U8980 (N_8980,N_613,N_4649);
and U8981 (N_8981,N_1402,N_3196);
nor U8982 (N_8982,N_3680,N_115);
and U8983 (N_8983,N_936,N_837);
nor U8984 (N_8984,N_1296,N_4982);
and U8985 (N_8985,N_3498,N_1795);
xnor U8986 (N_8986,N_2672,N_2372);
or U8987 (N_8987,N_2042,N_1249);
nor U8988 (N_8988,N_3879,N_94);
and U8989 (N_8989,N_2664,N_3535);
xor U8990 (N_8990,N_3166,N_3892);
or U8991 (N_8991,N_3042,N_500);
xnor U8992 (N_8992,N_4992,N_1375);
nor U8993 (N_8993,N_1476,N_4617);
nor U8994 (N_8994,N_1442,N_471);
and U8995 (N_8995,N_614,N_367);
or U8996 (N_8996,N_144,N_2957);
nor U8997 (N_8997,N_2468,N_4641);
or U8998 (N_8998,N_1692,N_2563);
and U8999 (N_8999,N_638,N_3406);
or U9000 (N_9000,N_3928,N_4040);
and U9001 (N_9001,N_2404,N_3764);
xor U9002 (N_9002,N_4536,N_2979);
nor U9003 (N_9003,N_1255,N_966);
xor U9004 (N_9004,N_4049,N_2617);
nor U9005 (N_9005,N_1908,N_626);
nor U9006 (N_9006,N_3427,N_432);
nor U9007 (N_9007,N_887,N_4920);
xor U9008 (N_9008,N_3653,N_3675);
and U9009 (N_9009,N_2141,N_1281);
or U9010 (N_9010,N_779,N_1845);
nor U9011 (N_9011,N_175,N_2142);
nand U9012 (N_9012,N_4359,N_4870);
nand U9013 (N_9013,N_2651,N_4459);
nor U9014 (N_9014,N_2420,N_4502);
and U9015 (N_9015,N_283,N_1389);
and U9016 (N_9016,N_3008,N_1362);
nand U9017 (N_9017,N_2400,N_3713);
and U9018 (N_9018,N_2790,N_939);
nand U9019 (N_9019,N_824,N_1183);
nor U9020 (N_9020,N_1590,N_1429);
and U9021 (N_9021,N_2972,N_4185);
nor U9022 (N_9022,N_1701,N_1115);
nand U9023 (N_9023,N_4425,N_448);
or U9024 (N_9024,N_967,N_2065);
and U9025 (N_9025,N_4025,N_3383);
nor U9026 (N_9026,N_3717,N_4080);
nor U9027 (N_9027,N_4009,N_2150);
xnor U9028 (N_9028,N_4174,N_1817);
nor U9029 (N_9029,N_2691,N_4703);
and U9030 (N_9030,N_650,N_2038);
xor U9031 (N_9031,N_3453,N_3235);
nand U9032 (N_9032,N_1499,N_4031);
nand U9033 (N_9033,N_2364,N_1609);
xor U9034 (N_9034,N_3929,N_4613);
or U9035 (N_9035,N_107,N_2953);
xnor U9036 (N_9036,N_694,N_4878);
and U9037 (N_9037,N_2283,N_4916);
nand U9038 (N_9038,N_2285,N_413);
nand U9039 (N_9039,N_599,N_2539);
and U9040 (N_9040,N_1113,N_4803);
xnor U9041 (N_9041,N_3710,N_4644);
or U9042 (N_9042,N_4792,N_2207);
and U9043 (N_9043,N_3250,N_2397);
and U9044 (N_9044,N_577,N_172);
and U9045 (N_9045,N_4990,N_1259);
or U9046 (N_9046,N_4077,N_2993);
or U9047 (N_9047,N_4457,N_1709);
or U9048 (N_9048,N_931,N_77);
xor U9049 (N_9049,N_570,N_289);
nor U9050 (N_9050,N_522,N_444);
nand U9051 (N_9051,N_3414,N_102);
nand U9052 (N_9052,N_1358,N_2065);
nand U9053 (N_9053,N_4145,N_2993);
or U9054 (N_9054,N_353,N_3134);
nand U9055 (N_9055,N_2951,N_2698);
xor U9056 (N_9056,N_2278,N_1482);
or U9057 (N_9057,N_3390,N_1369);
and U9058 (N_9058,N_3934,N_2218);
nand U9059 (N_9059,N_1508,N_747);
and U9060 (N_9060,N_4452,N_2755);
or U9061 (N_9061,N_4213,N_1261);
xor U9062 (N_9062,N_4301,N_4772);
xor U9063 (N_9063,N_2181,N_1720);
and U9064 (N_9064,N_4401,N_2139);
nand U9065 (N_9065,N_4064,N_4763);
nor U9066 (N_9066,N_3100,N_2327);
nand U9067 (N_9067,N_2514,N_2963);
xnor U9068 (N_9068,N_3985,N_440);
xnor U9069 (N_9069,N_4759,N_2196);
nor U9070 (N_9070,N_139,N_3201);
nor U9071 (N_9071,N_4946,N_1086);
and U9072 (N_9072,N_2773,N_3237);
xor U9073 (N_9073,N_780,N_558);
nor U9074 (N_9074,N_2324,N_406);
xor U9075 (N_9075,N_1644,N_448);
or U9076 (N_9076,N_4997,N_1031);
xnor U9077 (N_9077,N_1612,N_3636);
nor U9078 (N_9078,N_601,N_854);
nor U9079 (N_9079,N_1735,N_1135);
nand U9080 (N_9080,N_2350,N_3124);
nor U9081 (N_9081,N_2550,N_4301);
xnor U9082 (N_9082,N_4998,N_1339);
nor U9083 (N_9083,N_476,N_252);
nand U9084 (N_9084,N_4902,N_313);
nand U9085 (N_9085,N_3748,N_1428);
nor U9086 (N_9086,N_3529,N_779);
and U9087 (N_9087,N_1469,N_3033);
nand U9088 (N_9088,N_4657,N_2613);
xnor U9089 (N_9089,N_2025,N_623);
or U9090 (N_9090,N_1850,N_3768);
nor U9091 (N_9091,N_195,N_4717);
and U9092 (N_9092,N_2442,N_3573);
or U9093 (N_9093,N_3497,N_2148);
and U9094 (N_9094,N_3695,N_4172);
xor U9095 (N_9095,N_986,N_2959);
and U9096 (N_9096,N_581,N_3200);
xor U9097 (N_9097,N_2940,N_99);
nand U9098 (N_9098,N_823,N_4992);
xnor U9099 (N_9099,N_2336,N_754);
xor U9100 (N_9100,N_62,N_4868);
nand U9101 (N_9101,N_1973,N_4554);
and U9102 (N_9102,N_120,N_4734);
nor U9103 (N_9103,N_1480,N_2459);
or U9104 (N_9104,N_2246,N_679);
nor U9105 (N_9105,N_277,N_1183);
nor U9106 (N_9106,N_3940,N_511);
xnor U9107 (N_9107,N_3090,N_1754);
or U9108 (N_9108,N_1121,N_4907);
nor U9109 (N_9109,N_93,N_2041);
nand U9110 (N_9110,N_3273,N_3540);
or U9111 (N_9111,N_3946,N_3728);
and U9112 (N_9112,N_2540,N_2773);
or U9113 (N_9113,N_1689,N_4804);
xnor U9114 (N_9114,N_3816,N_3110);
xnor U9115 (N_9115,N_1874,N_4269);
or U9116 (N_9116,N_1957,N_3069);
nor U9117 (N_9117,N_3591,N_2275);
nor U9118 (N_9118,N_1181,N_1421);
nor U9119 (N_9119,N_4251,N_4188);
or U9120 (N_9120,N_3448,N_407);
or U9121 (N_9121,N_4800,N_3142);
xnor U9122 (N_9122,N_3763,N_2391);
or U9123 (N_9123,N_1433,N_1080);
nand U9124 (N_9124,N_4751,N_4688);
nand U9125 (N_9125,N_4978,N_1109);
and U9126 (N_9126,N_3998,N_860);
and U9127 (N_9127,N_1428,N_4752);
and U9128 (N_9128,N_4873,N_4232);
nand U9129 (N_9129,N_1991,N_1329);
nor U9130 (N_9130,N_3858,N_2888);
or U9131 (N_9131,N_454,N_2693);
and U9132 (N_9132,N_1210,N_2699);
nor U9133 (N_9133,N_3157,N_1253);
or U9134 (N_9134,N_463,N_842);
or U9135 (N_9135,N_3223,N_4141);
nand U9136 (N_9136,N_1401,N_892);
nor U9137 (N_9137,N_288,N_3568);
or U9138 (N_9138,N_699,N_4388);
nand U9139 (N_9139,N_40,N_3536);
xor U9140 (N_9140,N_3718,N_311);
and U9141 (N_9141,N_2982,N_803);
and U9142 (N_9142,N_4541,N_3807);
or U9143 (N_9143,N_4381,N_4181);
or U9144 (N_9144,N_2311,N_4435);
and U9145 (N_9145,N_3931,N_3249);
and U9146 (N_9146,N_3280,N_1123);
nand U9147 (N_9147,N_543,N_1367);
xor U9148 (N_9148,N_1913,N_1808);
and U9149 (N_9149,N_4898,N_2391);
or U9150 (N_9150,N_1036,N_1259);
nand U9151 (N_9151,N_3819,N_954);
xor U9152 (N_9152,N_2528,N_2869);
xnor U9153 (N_9153,N_1244,N_4145);
and U9154 (N_9154,N_2490,N_1519);
nand U9155 (N_9155,N_548,N_4999);
xnor U9156 (N_9156,N_734,N_422);
nor U9157 (N_9157,N_1088,N_2718);
or U9158 (N_9158,N_1033,N_2402);
nor U9159 (N_9159,N_4733,N_2066);
nor U9160 (N_9160,N_3478,N_3582);
and U9161 (N_9161,N_65,N_127);
nand U9162 (N_9162,N_4400,N_424);
xor U9163 (N_9163,N_3884,N_3459);
nand U9164 (N_9164,N_2010,N_2258);
or U9165 (N_9165,N_2110,N_487);
and U9166 (N_9166,N_697,N_3920);
nand U9167 (N_9167,N_2369,N_1053);
nand U9168 (N_9168,N_1736,N_3456);
xor U9169 (N_9169,N_4662,N_2579);
or U9170 (N_9170,N_1502,N_1535);
nand U9171 (N_9171,N_2788,N_4114);
nor U9172 (N_9172,N_4632,N_3140);
nor U9173 (N_9173,N_3309,N_3351);
nor U9174 (N_9174,N_538,N_1560);
or U9175 (N_9175,N_4148,N_1807);
xnor U9176 (N_9176,N_2962,N_1931);
xnor U9177 (N_9177,N_3270,N_2042);
or U9178 (N_9178,N_1177,N_1119);
nor U9179 (N_9179,N_3084,N_3313);
nand U9180 (N_9180,N_4837,N_2866);
xor U9181 (N_9181,N_2361,N_2752);
nand U9182 (N_9182,N_2032,N_3204);
or U9183 (N_9183,N_1240,N_3318);
nand U9184 (N_9184,N_4416,N_4388);
nand U9185 (N_9185,N_3613,N_1176);
and U9186 (N_9186,N_1814,N_755);
xor U9187 (N_9187,N_2697,N_3834);
xnor U9188 (N_9188,N_859,N_1581);
and U9189 (N_9189,N_1027,N_1425);
nor U9190 (N_9190,N_4796,N_1065);
nor U9191 (N_9191,N_2086,N_4120);
nor U9192 (N_9192,N_2328,N_1172);
or U9193 (N_9193,N_4715,N_3116);
nand U9194 (N_9194,N_2184,N_1842);
and U9195 (N_9195,N_515,N_1764);
nor U9196 (N_9196,N_4777,N_566);
or U9197 (N_9197,N_2374,N_902);
nor U9198 (N_9198,N_538,N_1387);
and U9199 (N_9199,N_2349,N_1444);
nand U9200 (N_9200,N_2463,N_360);
nand U9201 (N_9201,N_3363,N_4956);
nor U9202 (N_9202,N_3974,N_2998);
xor U9203 (N_9203,N_4737,N_843);
nor U9204 (N_9204,N_1611,N_3455);
nor U9205 (N_9205,N_3055,N_1989);
nand U9206 (N_9206,N_3211,N_617);
nor U9207 (N_9207,N_995,N_4291);
or U9208 (N_9208,N_896,N_3518);
nor U9209 (N_9209,N_2229,N_3615);
nand U9210 (N_9210,N_215,N_973);
xnor U9211 (N_9211,N_1800,N_1609);
nor U9212 (N_9212,N_496,N_42);
and U9213 (N_9213,N_3479,N_4245);
or U9214 (N_9214,N_4414,N_628);
nand U9215 (N_9215,N_1515,N_1831);
nor U9216 (N_9216,N_594,N_4010);
and U9217 (N_9217,N_366,N_1947);
and U9218 (N_9218,N_857,N_3527);
and U9219 (N_9219,N_1926,N_4674);
nand U9220 (N_9220,N_3110,N_4108);
or U9221 (N_9221,N_1936,N_461);
nand U9222 (N_9222,N_4165,N_153);
xor U9223 (N_9223,N_3487,N_2997);
or U9224 (N_9224,N_593,N_3093);
nand U9225 (N_9225,N_2332,N_2716);
and U9226 (N_9226,N_1049,N_1719);
or U9227 (N_9227,N_4503,N_1716);
and U9228 (N_9228,N_767,N_1284);
nor U9229 (N_9229,N_42,N_3187);
nand U9230 (N_9230,N_4090,N_3073);
nand U9231 (N_9231,N_1272,N_4720);
and U9232 (N_9232,N_4632,N_3985);
xnor U9233 (N_9233,N_2290,N_3623);
or U9234 (N_9234,N_3342,N_3714);
nand U9235 (N_9235,N_2596,N_1149);
and U9236 (N_9236,N_307,N_3291);
nor U9237 (N_9237,N_3035,N_2034);
and U9238 (N_9238,N_3439,N_3949);
or U9239 (N_9239,N_4677,N_96);
nand U9240 (N_9240,N_1125,N_2236);
xor U9241 (N_9241,N_2185,N_1760);
and U9242 (N_9242,N_4713,N_2699);
or U9243 (N_9243,N_280,N_2783);
nor U9244 (N_9244,N_3402,N_394);
xnor U9245 (N_9245,N_3924,N_1609);
nand U9246 (N_9246,N_3390,N_3018);
xnor U9247 (N_9247,N_2882,N_3254);
xnor U9248 (N_9248,N_219,N_3806);
or U9249 (N_9249,N_3699,N_4515);
and U9250 (N_9250,N_4736,N_3306);
nor U9251 (N_9251,N_1963,N_122);
and U9252 (N_9252,N_1566,N_4881);
or U9253 (N_9253,N_1715,N_3962);
xnor U9254 (N_9254,N_1181,N_1548);
xor U9255 (N_9255,N_514,N_3842);
and U9256 (N_9256,N_1525,N_3167);
and U9257 (N_9257,N_4662,N_64);
nand U9258 (N_9258,N_2862,N_3854);
nor U9259 (N_9259,N_819,N_1415);
and U9260 (N_9260,N_1717,N_3818);
and U9261 (N_9261,N_2283,N_3683);
nand U9262 (N_9262,N_4960,N_1289);
and U9263 (N_9263,N_3700,N_2986);
nor U9264 (N_9264,N_3424,N_1822);
nand U9265 (N_9265,N_4515,N_649);
or U9266 (N_9266,N_642,N_4055);
and U9267 (N_9267,N_1255,N_1560);
and U9268 (N_9268,N_3116,N_2745);
nand U9269 (N_9269,N_3285,N_4502);
and U9270 (N_9270,N_2210,N_3298);
and U9271 (N_9271,N_3355,N_2934);
nand U9272 (N_9272,N_1307,N_3555);
or U9273 (N_9273,N_3880,N_4529);
xnor U9274 (N_9274,N_2706,N_2798);
or U9275 (N_9275,N_1113,N_3209);
and U9276 (N_9276,N_942,N_4041);
xnor U9277 (N_9277,N_18,N_4575);
nand U9278 (N_9278,N_886,N_4208);
nand U9279 (N_9279,N_1459,N_117);
or U9280 (N_9280,N_2379,N_412);
xnor U9281 (N_9281,N_4406,N_502);
or U9282 (N_9282,N_1737,N_4357);
or U9283 (N_9283,N_2819,N_805);
or U9284 (N_9284,N_2481,N_2120);
nand U9285 (N_9285,N_4289,N_829);
or U9286 (N_9286,N_2956,N_764);
xor U9287 (N_9287,N_1055,N_301);
nand U9288 (N_9288,N_1436,N_3444);
nand U9289 (N_9289,N_3714,N_2202);
xnor U9290 (N_9290,N_2445,N_4779);
nand U9291 (N_9291,N_1722,N_3696);
and U9292 (N_9292,N_2450,N_2366);
nand U9293 (N_9293,N_228,N_2446);
and U9294 (N_9294,N_713,N_3427);
nand U9295 (N_9295,N_3954,N_2314);
xnor U9296 (N_9296,N_2378,N_3044);
xnor U9297 (N_9297,N_768,N_1609);
or U9298 (N_9298,N_2255,N_861);
xnor U9299 (N_9299,N_1671,N_1431);
xnor U9300 (N_9300,N_4758,N_22);
or U9301 (N_9301,N_4173,N_1439);
nand U9302 (N_9302,N_1317,N_3118);
or U9303 (N_9303,N_3245,N_2273);
xnor U9304 (N_9304,N_1146,N_4340);
nand U9305 (N_9305,N_4864,N_3391);
and U9306 (N_9306,N_156,N_2561);
or U9307 (N_9307,N_1252,N_2682);
nor U9308 (N_9308,N_604,N_3104);
nor U9309 (N_9309,N_1216,N_3214);
and U9310 (N_9310,N_173,N_4380);
nand U9311 (N_9311,N_2613,N_4179);
or U9312 (N_9312,N_3292,N_418);
nor U9313 (N_9313,N_3544,N_82);
or U9314 (N_9314,N_1101,N_2141);
nor U9315 (N_9315,N_224,N_4841);
nand U9316 (N_9316,N_4373,N_3853);
or U9317 (N_9317,N_8,N_2223);
or U9318 (N_9318,N_2641,N_3586);
xor U9319 (N_9319,N_178,N_4558);
and U9320 (N_9320,N_1532,N_2995);
xnor U9321 (N_9321,N_2617,N_2859);
nor U9322 (N_9322,N_982,N_3326);
or U9323 (N_9323,N_659,N_1310);
and U9324 (N_9324,N_4052,N_346);
nand U9325 (N_9325,N_3859,N_2707);
or U9326 (N_9326,N_1933,N_3707);
nand U9327 (N_9327,N_4464,N_733);
and U9328 (N_9328,N_792,N_4096);
xnor U9329 (N_9329,N_558,N_950);
xnor U9330 (N_9330,N_4585,N_3869);
or U9331 (N_9331,N_4317,N_2756);
nor U9332 (N_9332,N_471,N_590);
and U9333 (N_9333,N_2165,N_2852);
or U9334 (N_9334,N_3894,N_1703);
xor U9335 (N_9335,N_4090,N_4053);
xnor U9336 (N_9336,N_189,N_1440);
or U9337 (N_9337,N_3027,N_1168);
xnor U9338 (N_9338,N_3376,N_2763);
nand U9339 (N_9339,N_1143,N_1258);
nand U9340 (N_9340,N_1406,N_609);
and U9341 (N_9341,N_2702,N_4764);
nor U9342 (N_9342,N_3965,N_1230);
nand U9343 (N_9343,N_1518,N_2479);
nand U9344 (N_9344,N_4288,N_3106);
or U9345 (N_9345,N_1664,N_1622);
nand U9346 (N_9346,N_3135,N_119);
xnor U9347 (N_9347,N_1785,N_3968);
and U9348 (N_9348,N_2760,N_4360);
or U9349 (N_9349,N_739,N_3618);
and U9350 (N_9350,N_3468,N_4299);
nor U9351 (N_9351,N_392,N_3137);
xnor U9352 (N_9352,N_2656,N_4675);
and U9353 (N_9353,N_3514,N_4346);
nor U9354 (N_9354,N_1681,N_4114);
and U9355 (N_9355,N_1321,N_1770);
nand U9356 (N_9356,N_1818,N_2733);
or U9357 (N_9357,N_4405,N_645);
nand U9358 (N_9358,N_1217,N_2712);
nand U9359 (N_9359,N_1712,N_4802);
nand U9360 (N_9360,N_2111,N_2235);
xnor U9361 (N_9361,N_2246,N_1483);
nand U9362 (N_9362,N_2901,N_432);
and U9363 (N_9363,N_1759,N_2290);
or U9364 (N_9364,N_3191,N_3589);
nor U9365 (N_9365,N_3070,N_1723);
nand U9366 (N_9366,N_4562,N_1098);
nand U9367 (N_9367,N_2166,N_4247);
or U9368 (N_9368,N_1047,N_3906);
or U9369 (N_9369,N_3581,N_1550);
nor U9370 (N_9370,N_4413,N_4278);
nor U9371 (N_9371,N_271,N_2274);
xnor U9372 (N_9372,N_2883,N_3613);
nor U9373 (N_9373,N_4039,N_524);
nor U9374 (N_9374,N_4739,N_321);
xor U9375 (N_9375,N_4225,N_4789);
or U9376 (N_9376,N_89,N_4059);
nand U9377 (N_9377,N_3932,N_4622);
nor U9378 (N_9378,N_411,N_2358);
xnor U9379 (N_9379,N_1144,N_1558);
nand U9380 (N_9380,N_291,N_2705);
nand U9381 (N_9381,N_2396,N_580);
nor U9382 (N_9382,N_116,N_1470);
and U9383 (N_9383,N_2476,N_3036);
nand U9384 (N_9384,N_2906,N_1429);
nor U9385 (N_9385,N_1602,N_2888);
or U9386 (N_9386,N_4773,N_588);
nor U9387 (N_9387,N_3292,N_3199);
xnor U9388 (N_9388,N_3125,N_57);
xor U9389 (N_9389,N_3768,N_4591);
and U9390 (N_9390,N_1219,N_4046);
nor U9391 (N_9391,N_4722,N_339);
nand U9392 (N_9392,N_3635,N_2982);
nor U9393 (N_9393,N_2041,N_1954);
xor U9394 (N_9394,N_2113,N_3548);
or U9395 (N_9395,N_1355,N_3955);
and U9396 (N_9396,N_4371,N_4967);
nor U9397 (N_9397,N_4990,N_865);
nand U9398 (N_9398,N_2323,N_1578);
nand U9399 (N_9399,N_169,N_4150);
and U9400 (N_9400,N_783,N_4523);
nor U9401 (N_9401,N_4312,N_1393);
nor U9402 (N_9402,N_622,N_2453);
or U9403 (N_9403,N_2390,N_1314);
xor U9404 (N_9404,N_4982,N_494);
xnor U9405 (N_9405,N_2692,N_4294);
nor U9406 (N_9406,N_2783,N_4917);
nand U9407 (N_9407,N_1873,N_807);
nand U9408 (N_9408,N_3212,N_1798);
and U9409 (N_9409,N_943,N_432);
or U9410 (N_9410,N_1879,N_977);
nor U9411 (N_9411,N_769,N_2727);
or U9412 (N_9412,N_2286,N_548);
or U9413 (N_9413,N_3447,N_1236);
or U9414 (N_9414,N_333,N_3848);
xnor U9415 (N_9415,N_1228,N_505);
and U9416 (N_9416,N_92,N_3887);
or U9417 (N_9417,N_623,N_561);
and U9418 (N_9418,N_2755,N_2578);
xor U9419 (N_9419,N_2427,N_309);
nand U9420 (N_9420,N_69,N_2532);
xor U9421 (N_9421,N_3677,N_527);
or U9422 (N_9422,N_864,N_1435);
nand U9423 (N_9423,N_3066,N_3869);
nor U9424 (N_9424,N_4535,N_4036);
nand U9425 (N_9425,N_1288,N_2406);
nor U9426 (N_9426,N_1795,N_2952);
or U9427 (N_9427,N_680,N_2877);
nor U9428 (N_9428,N_1184,N_4026);
nor U9429 (N_9429,N_4132,N_701);
nor U9430 (N_9430,N_3942,N_4109);
nor U9431 (N_9431,N_3936,N_4616);
nor U9432 (N_9432,N_4862,N_3904);
xor U9433 (N_9433,N_3482,N_732);
and U9434 (N_9434,N_4116,N_3233);
nor U9435 (N_9435,N_2260,N_2729);
and U9436 (N_9436,N_1027,N_2406);
or U9437 (N_9437,N_3505,N_2508);
nor U9438 (N_9438,N_105,N_2417);
nand U9439 (N_9439,N_2457,N_2795);
or U9440 (N_9440,N_1707,N_2530);
and U9441 (N_9441,N_4514,N_3877);
nor U9442 (N_9442,N_3792,N_1345);
nand U9443 (N_9443,N_4829,N_2896);
nand U9444 (N_9444,N_3909,N_1416);
nor U9445 (N_9445,N_3343,N_1327);
xnor U9446 (N_9446,N_768,N_2343);
and U9447 (N_9447,N_3196,N_1506);
nor U9448 (N_9448,N_2881,N_4823);
or U9449 (N_9449,N_708,N_1281);
nand U9450 (N_9450,N_4685,N_2659);
nor U9451 (N_9451,N_1386,N_3752);
nand U9452 (N_9452,N_2590,N_801);
or U9453 (N_9453,N_4569,N_3582);
nand U9454 (N_9454,N_3234,N_4940);
or U9455 (N_9455,N_252,N_2123);
xor U9456 (N_9456,N_3799,N_100);
or U9457 (N_9457,N_68,N_1017);
nor U9458 (N_9458,N_2282,N_4484);
and U9459 (N_9459,N_751,N_2299);
nand U9460 (N_9460,N_3058,N_158);
xor U9461 (N_9461,N_3156,N_2129);
nor U9462 (N_9462,N_1301,N_577);
nand U9463 (N_9463,N_2715,N_4432);
nand U9464 (N_9464,N_3495,N_3700);
nor U9465 (N_9465,N_3625,N_1563);
xor U9466 (N_9466,N_2284,N_3327);
or U9467 (N_9467,N_88,N_3586);
nand U9468 (N_9468,N_2369,N_877);
nor U9469 (N_9469,N_1787,N_3716);
xor U9470 (N_9470,N_2780,N_4380);
and U9471 (N_9471,N_1950,N_1201);
xnor U9472 (N_9472,N_31,N_654);
xor U9473 (N_9473,N_1654,N_4273);
nand U9474 (N_9474,N_2904,N_1764);
nor U9475 (N_9475,N_2612,N_3798);
and U9476 (N_9476,N_1405,N_4759);
nor U9477 (N_9477,N_2487,N_1634);
xor U9478 (N_9478,N_3171,N_692);
or U9479 (N_9479,N_1624,N_2052);
or U9480 (N_9480,N_998,N_1047);
nor U9481 (N_9481,N_524,N_3825);
xnor U9482 (N_9482,N_2594,N_3930);
or U9483 (N_9483,N_1011,N_2639);
nand U9484 (N_9484,N_1945,N_1575);
nor U9485 (N_9485,N_2937,N_982);
xor U9486 (N_9486,N_2184,N_197);
xnor U9487 (N_9487,N_3974,N_947);
xnor U9488 (N_9488,N_4724,N_1753);
nand U9489 (N_9489,N_3470,N_2588);
xor U9490 (N_9490,N_3689,N_4306);
nand U9491 (N_9491,N_2196,N_1960);
xnor U9492 (N_9492,N_2435,N_768);
and U9493 (N_9493,N_187,N_4635);
and U9494 (N_9494,N_4444,N_3394);
nand U9495 (N_9495,N_3012,N_1188);
and U9496 (N_9496,N_189,N_829);
nand U9497 (N_9497,N_1236,N_4472);
and U9498 (N_9498,N_3216,N_613);
or U9499 (N_9499,N_413,N_1916);
nand U9500 (N_9500,N_953,N_2102);
xnor U9501 (N_9501,N_3075,N_135);
nand U9502 (N_9502,N_1762,N_4516);
or U9503 (N_9503,N_263,N_103);
or U9504 (N_9504,N_1761,N_1118);
or U9505 (N_9505,N_4741,N_4950);
nand U9506 (N_9506,N_623,N_3682);
nand U9507 (N_9507,N_197,N_122);
xnor U9508 (N_9508,N_3657,N_1121);
nand U9509 (N_9509,N_2895,N_4037);
nand U9510 (N_9510,N_4798,N_663);
and U9511 (N_9511,N_4885,N_2967);
nor U9512 (N_9512,N_4976,N_1494);
and U9513 (N_9513,N_2990,N_4071);
nor U9514 (N_9514,N_4746,N_2849);
nand U9515 (N_9515,N_1695,N_2213);
nand U9516 (N_9516,N_744,N_2272);
nor U9517 (N_9517,N_651,N_4323);
and U9518 (N_9518,N_4603,N_2616);
or U9519 (N_9519,N_1619,N_170);
and U9520 (N_9520,N_2938,N_4030);
or U9521 (N_9521,N_2180,N_835);
or U9522 (N_9522,N_3604,N_4211);
xnor U9523 (N_9523,N_306,N_2646);
and U9524 (N_9524,N_2035,N_4964);
and U9525 (N_9525,N_3365,N_723);
and U9526 (N_9526,N_2999,N_2842);
nand U9527 (N_9527,N_4065,N_1916);
nor U9528 (N_9528,N_1554,N_1080);
nand U9529 (N_9529,N_4527,N_2449);
nand U9530 (N_9530,N_2988,N_1274);
or U9531 (N_9531,N_3258,N_1685);
xor U9532 (N_9532,N_3065,N_1801);
or U9533 (N_9533,N_1286,N_490);
and U9534 (N_9534,N_1340,N_1185);
or U9535 (N_9535,N_2326,N_772);
xnor U9536 (N_9536,N_1375,N_2582);
or U9537 (N_9537,N_2623,N_4412);
nand U9538 (N_9538,N_3820,N_3559);
or U9539 (N_9539,N_2266,N_1137);
nor U9540 (N_9540,N_3393,N_542);
and U9541 (N_9541,N_2604,N_2267);
and U9542 (N_9542,N_458,N_3746);
and U9543 (N_9543,N_3590,N_3067);
nor U9544 (N_9544,N_4182,N_3724);
nor U9545 (N_9545,N_4915,N_193);
nand U9546 (N_9546,N_460,N_1311);
nor U9547 (N_9547,N_397,N_4408);
nor U9548 (N_9548,N_4870,N_3951);
or U9549 (N_9549,N_3971,N_3535);
xor U9550 (N_9550,N_4257,N_1729);
xor U9551 (N_9551,N_4446,N_3455);
and U9552 (N_9552,N_582,N_4748);
or U9553 (N_9553,N_1217,N_1283);
and U9554 (N_9554,N_1985,N_403);
nand U9555 (N_9555,N_2694,N_221);
nand U9556 (N_9556,N_630,N_674);
nor U9557 (N_9557,N_4382,N_4628);
nand U9558 (N_9558,N_2304,N_2591);
nor U9559 (N_9559,N_1702,N_4937);
or U9560 (N_9560,N_494,N_2971);
nor U9561 (N_9561,N_3293,N_3306);
nor U9562 (N_9562,N_2016,N_1412);
and U9563 (N_9563,N_4379,N_2671);
or U9564 (N_9564,N_1340,N_4727);
nor U9565 (N_9565,N_1360,N_4105);
xnor U9566 (N_9566,N_1216,N_938);
nand U9567 (N_9567,N_68,N_3275);
nand U9568 (N_9568,N_2597,N_3949);
or U9569 (N_9569,N_2430,N_1912);
and U9570 (N_9570,N_2174,N_30);
xor U9571 (N_9571,N_3108,N_4337);
nand U9572 (N_9572,N_3425,N_15);
xor U9573 (N_9573,N_684,N_1805);
nand U9574 (N_9574,N_3576,N_4864);
xnor U9575 (N_9575,N_4239,N_1809);
xnor U9576 (N_9576,N_2129,N_2184);
nand U9577 (N_9577,N_4250,N_885);
or U9578 (N_9578,N_3221,N_1067);
or U9579 (N_9579,N_2731,N_197);
and U9580 (N_9580,N_2617,N_1990);
nand U9581 (N_9581,N_1056,N_2788);
nand U9582 (N_9582,N_543,N_4606);
nor U9583 (N_9583,N_658,N_2092);
and U9584 (N_9584,N_3972,N_913);
nand U9585 (N_9585,N_4690,N_2253);
and U9586 (N_9586,N_2959,N_954);
nand U9587 (N_9587,N_3267,N_3671);
xnor U9588 (N_9588,N_2610,N_3374);
xnor U9589 (N_9589,N_3790,N_3012);
nor U9590 (N_9590,N_247,N_555);
and U9591 (N_9591,N_491,N_4878);
nand U9592 (N_9592,N_3813,N_4607);
or U9593 (N_9593,N_4512,N_2491);
xor U9594 (N_9594,N_3910,N_650);
xnor U9595 (N_9595,N_1343,N_45);
nor U9596 (N_9596,N_953,N_4446);
and U9597 (N_9597,N_1143,N_3810);
nand U9598 (N_9598,N_4838,N_298);
nor U9599 (N_9599,N_4961,N_3846);
nor U9600 (N_9600,N_396,N_763);
xnor U9601 (N_9601,N_3861,N_1558);
and U9602 (N_9602,N_4975,N_3413);
nand U9603 (N_9603,N_4002,N_1035);
and U9604 (N_9604,N_471,N_2228);
nor U9605 (N_9605,N_4978,N_1619);
and U9606 (N_9606,N_560,N_1124);
xnor U9607 (N_9607,N_4234,N_3598);
nand U9608 (N_9608,N_4610,N_1601);
nor U9609 (N_9609,N_505,N_2872);
xor U9610 (N_9610,N_3118,N_759);
xnor U9611 (N_9611,N_4191,N_3004);
and U9612 (N_9612,N_663,N_1330);
and U9613 (N_9613,N_2671,N_4753);
or U9614 (N_9614,N_2597,N_9);
and U9615 (N_9615,N_3717,N_3045);
xnor U9616 (N_9616,N_2633,N_1728);
and U9617 (N_9617,N_1519,N_109);
xnor U9618 (N_9618,N_4716,N_4400);
and U9619 (N_9619,N_1692,N_4817);
or U9620 (N_9620,N_1514,N_3975);
nor U9621 (N_9621,N_735,N_1571);
xnor U9622 (N_9622,N_396,N_2467);
and U9623 (N_9623,N_4056,N_4646);
nand U9624 (N_9624,N_186,N_1150);
nand U9625 (N_9625,N_2835,N_4706);
nor U9626 (N_9626,N_1457,N_1259);
xnor U9627 (N_9627,N_4366,N_3747);
nor U9628 (N_9628,N_3809,N_2040);
xnor U9629 (N_9629,N_1895,N_1097);
nand U9630 (N_9630,N_480,N_3004);
and U9631 (N_9631,N_3762,N_3586);
xor U9632 (N_9632,N_4935,N_4809);
xnor U9633 (N_9633,N_3023,N_4339);
nand U9634 (N_9634,N_468,N_3990);
nor U9635 (N_9635,N_4588,N_3936);
and U9636 (N_9636,N_1115,N_2287);
nand U9637 (N_9637,N_2548,N_4840);
or U9638 (N_9638,N_4428,N_22);
or U9639 (N_9639,N_3490,N_1347);
or U9640 (N_9640,N_2537,N_4926);
xnor U9641 (N_9641,N_3188,N_4782);
and U9642 (N_9642,N_1335,N_1346);
nor U9643 (N_9643,N_4439,N_1458);
or U9644 (N_9644,N_2566,N_3092);
nor U9645 (N_9645,N_4960,N_3995);
xor U9646 (N_9646,N_3887,N_4051);
nor U9647 (N_9647,N_729,N_1086);
xnor U9648 (N_9648,N_4144,N_4794);
xor U9649 (N_9649,N_3569,N_4415);
nor U9650 (N_9650,N_4826,N_4837);
or U9651 (N_9651,N_4864,N_3933);
and U9652 (N_9652,N_2376,N_2773);
or U9653 (N_9653,N_4995,N_5);
or U9654 (N_9654,N_834,N_3367);
nor U9655 (N_9655,N_3421,N_3539);
nand U9656 (N_9656,N_4081,N_1104);
nand U9657 (N_9657,N_2880,N_1254);
xnor U9658 (N_9658,N_4962,N_1349);
xor U9659 (N_9659,N_50,N_3704);
xnor U9660 (N_9660,N_987,N_2709);
or U9661 (N_9661,N_2736,N_2336);
and U9662 (N_9662,N_2080,N_998);
nor U9663 (N_9663,N_440,N_3424);
nand U9664 (N_9664,N_318,N_1125);
and U9665 (N_9665,N_1890,N_347);
nor U9666 (N_9666,N_306,N_1217);
nand U9667 (N_9667,N_515,N_3877);
xor U9668 (N_9668,N_1567,N_1371);
xnor U9669 (N_9669,N_2633,N_2447);
nor U9670 (N_9670,N_3553,N_1047);
or U9671 (N_9671,N_576,N_1350);
and U9672 (N_9672,N_334,N_1911);
nand U9673 (N_9673,N_4539,N_3126);
or U9674 (N_9674,N_3507,N_1635);
xnor U9675 (N_9675,N_860,N_75);
or U9676 (N_9676,N_1842,N_3153);
and U9677 (N_9677,N_4002,N_1179);
or U9678 (N_9678,N_2752,N_561);
or U9679 (N_9679,N_14,N_2745);
xnor U9680 (N_9680,N_1902,N_1846);
xnor U9681 (N_9681,N_1148,N_3542);
xnor U9682 (N_9682,N_1365,N_3870);
xor U9683 (N_9683,N_1369,N_3924);
nor U9684 (N_9684,N_508,N_43);
nand U9685 (N_9685,N_3218,N_656);
or U9686 (N_9686,N_1575,N_4010);
and U9687 (N_9687,N_2644,N_1882);
nor U9688 (N_9688,N_2200,N_2759);
xnor U9689 (N_9689,N_4208,N_2609);
xor U9690 (N_9690,N_1795,N_1482);
nand U9691 (N_9691,N_556,N_1396);
or U9692 (N_9692,N_3272,N_2142);
nand U9693 (N_9693,N_1293,N_3031);
and U9694 (N_9694,N_3762,N_2120);
and U9695 (N_9695,N_3820,N_1304);
nor U9696 (N_9696,N_3285,N_3217);
and U9697 (N_9697,N_1346,N_1937);
nand U9698 (N_9698,N_229,N_4765);
nand U9699 (N_9699,N_1823,N_2023);
nor U9700 (N_9700,N_2573,N_4738);
nand U9701 (N_9701,N_2338,N_1090);
nand U9702 (N_9702,N_191,N_3615);
or U9703 (N_9703,N_2731,N_2048);
and U9704 (N_9704,N_3644,N_1352);
nor U9705 (N_9705,N_4022,N_1701);
nor U9706 (N_9706,N_2036,N_3513);
nor U9707 (N_9707,N_834,N_2785);
or U9708 (N_9708,N_4851,N_1268);
and U9709 (N_9709,N_3941,N_3707);
and U9710 (N_9710,N_4044,N_2528);
nand U9711 (N_9711,N_867,N_925);
xor U9712 (N_9712,N_283,N_862);
and U9713 (N_9713,N_3678,N_1356);
and U9714 (N_9714,N_4160,N_3017);
or U9715 (N_9715,N_2688,N_1046);
nand U9716 (N_9716,N_1880,N_36);
nand U9717 (N_9717,N_4707,N_782);
xnor U9718 (N_9718,N_570,N_3404);
nand U9719 (N_9719,N_4290,N_2347);
nand U9720 (N_9720,N_4611,N_1944);
nor U9721 (N_9721,N_3522,N_334);
or U9722 (N_9722,N_2963,N_596);
nand U9723 (N_9723,N_970,N_892);
nand U9724 (N_9724,N_3064,N_1020);
or U9725 (N_9725,N_2841,N_2110);
nor U9726 (N_9726,N_2121,N_652);
nor U9727 (N_9727,N_3238,N_4851);
nand U9728 (N_9728,N_2364,N_473);
or U9729 (N_9729,N_1330,N_2653);
nand U9730 (N_9730,N_1560,N_513);
nand U9731 (N_9731,N_3067,N_4733);
or U9732 (N_9732,N_1214,N_1640);
nor U9733 (N_9733,N_3855,N_970);
nor U9734 (N_9734,N_4171,N_2045);
or U9735 (N_9735,N_1701,N_1240);
nand U9736 (N_9736,N_942,N_629);
nand U9737 (N_9737,N_4591,N_4130);
xor U9738 (N_9738,N_1180,N_394);
nor U9739 (N_9739,N_4301,N_2481);
xor U9740 (N_9740,N_4693,N_611);
or U9741 (N_9741,N_2163,N_2721);
or U9742 (N_9742,N_2145,N_3914);
xnor U9743 (N_9743,N_3059,N_504);
nand U9744 (N_9744,N_1263,N_321);
and U9745 (N_9745,N_3707,N_1489);
xnor U9746 (N_9746,N_2620,N_1460);
xnor U9747 (N_9747,N_1970,N_1143);
and U9748 (N_9748,N_4651,N_3482);
nand U9749 (N_9749,N_3367,N_4601);
nand U9750 (N_9750,N_1918,N_4771);
xnor U9751 (N_9751,N_1431,N_358);
or U9752 (N_9752,N_2100,N_3794);
and U9753 (N_9753,N_345,N_2850);
nor U9754 (N_9754,N_1156,N_719);
nor U9755 (N_9755,N_2541,N_3837);
xnor U9756 (N_9756,N_3067,N_4659);
or U9757 (N_9757,N_1468,N_3950);
nor U9758 (N_9758,N_3221,N_1566);
and U9759 (N_9759,N_1427,N_3247);
nand U9760 (N_9760,N_3335,N_2966);
xor U9761 (N_9761,N_54,N_3640);
nand U9762 (N_9762,N_3888,N_4192);
and U9763 (N_9763,N_3577,N_1976);
nand U9764 (N_9764,N_4798,N_1244);
and U9765 (N_9765,N_549,N_3280);
nor U9766 (N_9766,N_1170,N_4316);
xnor U9767 (N_9767,N_3691,N_863);
xnor U9768 (N_9768,N_1284,N_4591);
and U9769 (N_9769,N_4077,N_3090);
and U9770 (N_9770,N_17,N_2169);
xor U9771 (N_9771,N_563,N_1282);
nor U9772 (N_9772,N_1700,N_1303);
nor U9773 (N_9773,N_4684,N_1072);
or U9774 (N_9774,N_1687,N_701);
or U9775 (N_9775,N_854,N_1481);
or U9776 (N_9776,N_283,N_207);
and U9777 (N_9777,N_3017,N_276);
and U9778 (N_9778,N_543,N_508);
and U9779 (N_9779,N_2746,N_2911);
nand U9780 (N_9780,N_453,N_4570);
xnor U9781 (N_9781,N_4112,N_3395);
nor U9782 (N_9782,N_1869,N_2165);
nor U9783 (N_9783,N_3361,N_4182);
or U9784 (N_9784,N_4110,N_2600);
and U9785 (N_9785,N_2004,N_1114);
xor U9786 (N_9786,N_2768,N_1942);
xor U9787 (N_9787,N_3052,N_264);
and U9788 (N_9788,N_1910,N_2705);
nand U9789 (N_9789,N_4051,N_456);
nand U9790 (N_9790,N_4216,N_898);
nand U9791 (N_9791,N_1296,N_2745);
xnor U9792 (N_9792,N_4864,N_4631);
nor U9793 (N_9793,N_4832,N_2091);
and U9794 (N_9794,N_3342,N_3722);
and U9795 (N_9795,N_4087,N_4455);
and U9796 (N_9796,N_876,N_2008);
and U9797 (N_9797,N_3493,N_2975);
xnor U9798 (N_9798,N_16,N_1621);
nand U9799 (N_9799,N_3886,N_1927);
nand U9800 (N_9800,N_3533,N_1288);
nand U9801 (N_9801,N_3039,N_1271);
xor U9802 (N_9802,N_2897,N_1558);
and U9803 (N_9803,N_112,N_1621);
nor U9804 (N_9804,N_4968,N_4880);
nor U9805 (N_9805,N_1556,N_753);
nand U9806 (N_9806,N_4984,N_1029);
nand U9807 (N_9807,N_2055,N_3963);
nand U9808 (N_9808,N_1408,N_1752);
nor U9809 (N_9809,N_308,N_1893);
xnor U9810 (N_9810,N_424,N_3805);
nand U9811 (N_9811,N_55,N_2042);
and U9812 (N_9812,N_2819,N_1921);
and U9813 (N_9813,N_4438,N_4690);
nor U9814 (N_9814,N_1756,N_2723);
xnor U9815 (N_9815,N_58,N_3494);
and U9816 (N_9816,N_3922,N_3569);
or U9817 (N_9817,N_1192,N_127);
xor U9818 (N_9818,N_1581,N_1089);
or U9819 (N_9819,N_2349,N_4178);
and U9820 (N_9820,N_1518,N_2140);
xnor U9821 (N_9821,N_300,N_4997);
or U9822 (N_9822,N_2377,N_2598);
and U9823 (N_9823,N_3815,N_2873);
and U9824 (N_9824,N_1026,N_2119);
and U9825 (N_9825,N_4458,N_4692);
nor U9826 (N_9826,N_4673,N_4722);
nand U9827 (N_9827,N_2470,N_444);
xnor U9828 (N_9828,N_750,N_3213);
and U9829 (N_9829,N_3005,N_751);
or U9830 (N_9830,N_469,N_445);
nand U9831 (N_9831,N_4409,N_4774);
nand U9832 (N_9832,N_4561,N_1025);
nand U9833 (N_9833,N_1002,N_1455);
and U9834 (N_9834,N_1262,N_586);
or U9835 (N_9835,N_3678,N_2699);
nor U9836 (N_9836,N_1089,N_4308);
or U9837 (N_9837,N_815,N_207);
and U9838 (N_9838,N_4726,N_4856);
and U9839 (N_9839,N_4032,N_2566);
xor U9840 (N_9840,N_3867,N_546);
and U9841 (N_9841,N_3395,N_2948);
or U9842 (N_9842,N_497,N_2905);
xor U9843 (N_9843,N_2604,N_2589);
or U9844 (N_9844,N_89,N_4056);
or U9845 (N_9845,N_2235,N_3876);
xor U9846 (N_9846,N_4051,N_163);
nor U9847 (N_9847,N_3842,N_3234);
xnor U9848 (N_9848,N_450,N_3037);
xor U9849 (N_9849,N_4936,N_4439);
and U9850 (N_9850,N_782,N_4251);
and U9851 (N_9851,N_2935,N_2692);
xnor U9852 (N_9852,N_4821,N_4568);
nor U9853 (N_9853,N_88,N_1454);
nand U9854 (N_9854,N_4600,N_184);
xor U9855 (N_9855,N_1430,N_3874);
nor U9856 (N_9856,N_365,N_4882);
xor U9857 (N_9857,N_1701,N_4687);
or U9858 (N_9858,N_3965,N_241);
and U9859 (N_9859,N_4463,N_4913);
or U9860 (N_9860,N_1085,N_4806);
nor U9861 (N_9861,N_654,N_206);
and U9862 (N_9862,N_2773,N_3494);
and U9863 (N_9863,N_1475,N_1241);
or U9864 (N_9864,N_31,N_4502);
nor U9865 (N_9865,N_1182,N_2746);
and U9866 (N_9866,N_4172,N_1728);
or U9867 (N_9867,N_4458,N_14);
or U9868 (N_9868,N_919,N_1203);
nor U9869 (N_9869,N_4627,N_3770);
or U9870 (N_9870,N_3203,N_1053);
or U9871 (N_9871,N_2578,N_3162);
nand U9872 (N_9872,N_1834,N_717);
nand U9873 (N_9873,N_3350,N_464);
nand U9874 (N_9874,N_4087,N_2242);
nand U9875 (N_9875,N_4558,N_2308);
or U9876 (N_9876,N_850,N_1478);
and U9877 (N_9877,N_4869,N_4763);
xnor U9878 (N_9878,N_2388,N_1059);
nand U9879 (N_9879,N_556,N_4076);
nand U9880 (N_9880,N_678,N_1380);
nand U9881 (N_9881,N_363,N_3359);
and U9882 (N_9882,N_4972,N_4516);
xnor U9883 (N_9883,N_2339,N_321);
and U9884 (N_9884,N_1338,N_3820);
and U9885 (N_9885,N_3528,N_3230);
xor U9886 (N_9886,N_3611,N_1890);
or U9887 (N_9887,N_605,N_2998);
nand U9888 (N_9888,N_1258,N_3558);
xor U9889 (N_9889,N_4236,N_46);
or U9890 (N_9890,N_3689,N_2474);
nand U9891 (N_9891,N_742,N_1265);
or U9892 (N_9892,N_3560,N_2784);
nand U9893 (N_9893,N_276,N_2144);
xnor U9894 (N_9894,N_280,N_4156);
nand U9895 (N_9895,N_2758,N_3884);
xnor U9896 (N_9896,N_4258,N_2417);
nor U9897 (N_9897,N_4074,N_3599);
nand U9898 (N_9898,N_2055,N_4934);
nor U9899 (N_9899,N_3126,N_1964);
nand U9900 (N_9900,N_1362,N_4469);
xor U9901 (N_9901,N_1652,N_1237);
nand U9902 (N_9902,N_2245,N_1196);
xor U9903 (N_9903,N_2816,N_4814);
nand U9904 (N_9904,N_3174,N_1447);
and U9905 (N_9905,N_4114,N_4044);
xor U9906 (N_9906,N_2701,N_1432);
and U9907 (N_9907,N_1227,N_4061);
or U9908 (N_9908,N_2335,N_4159);
or U9909 (N_9909,N_1423,N_3289);
nor U9910 (N_9910,N_3413,N_987);
nand U9911 (N_9911,N_980,N_3426);
or U9912 (N_9912,N_4455,N_4740);
or U9913 (N_9913,N_4166,N_2419);
nor U9914 (N_9914,N_2475,N_1645);
nor U9915 (N_9915,N_47,N_1829);
and U9916 (N_9916,N_2250,N_2646);
xor U9917 (N_9917,N_3731,N_3425);
xor U9918 (N_9918,N_195,N_3758);
xor U9919 (N_9919,N_637,N_1187);
nand U9920 (N_9920,N_2953,N_164);
xnor U9921 (N_9921,N_2316,N_3222);
nand U9922 (N_9922,N_453,N_240);
nand U9923 (N_9923,N_4723,N_2278);
nor U9924 (N_9924,N_2296,N_4924);
nand U9925 (N_9925,N_319,N_320);
and U9926 (N_9926,N_3522,N_2997);
or U9927 (N_9927,N_3696,N_3144);
nor U9928 (N_9928,N_2668,N_2856);
nand U9929 (N_9929,N_2651,N_1081);
nand U9930 (N_9930,N_1938,N_4506);
nor U9931 (N_9931,N_3776,N_1627);
nor U9932 (N_9932,N_4514,N_4138);
and U9933 (N_9933,N_3011,N_2700);
xor U9934 (N_9934,N_1839,N_2712);
and U9935 (N_9935,N_3224,N_1423);
nor U9936 (N_9936,N_2515,N_1681);
and U9937 (N_9937,N_1402,N_253);
xor U9938 (N_9938,N_875,N_4043);
nor U9939 (N_9939,N_1795,N_3950);
nand U9940 (N_9940,N_3361,N_2664);
nor U9941 (N_9941,N_1222,N_2826);
nor U9942 (N_9942,N_3545,N_4894);
and U9943 (N_9943,N_2060,N_2759);
or U9944 (N_9944,N_4909,N_4053);
nand U9945 (N_9945,N_3983,N_3604);
and U9946 (N_9946,N_771,N_1203);
xnor U9947 (N_9947,N_4786,N_4404);
nor U9948 (N_9948,N_2255,N_1664);
nand U9949 (N_9949,N_3247,N_555);
and U9950 (N_9950,N_3266,N_4569);
or U9951 (N_9951,N_3009,N_1733);
nand U9952 (N_9952,N_4371,N_609);
and U9953 (N_9953,N_3210,N_3081);
or U9954 (N_9954,N_1166,N_2524);
xnor U9955 (N_9955,N_2998,N_1617);
xor U9956 (N_9956,N_247,N_952);
or U9957 (N_9957,N_535,N_3157);
nand U9958 (N_9958,N_4692,N_1131);
xor U9959 (N_9959,N_1975,N_2960);
and U9960 (N_9960,N_3591,N_3280);
and U9961 (N_9961,N_4480,N_2895);
nor U9962 (N_9962,N_1625,N_495);
nand U9963 (N_9963,N_1234,N_935);
and U9964 (N_9964,N_2075,N_67);
nor U9965 (N_9965,N_3268,N_4317);
and U9966 (N_9966,N_3901,N_1250);
nand U9967 (N_9967,N_565,N_1336);
and U9968 (N_9968,N_3776,N_3114);
nor U9969 (N_9969,N_2718,N_4049);
xor U9970 (N_9970,N_2813,N_4044);
or U9971 (N_9971,N_3886,N_3844);
nand U9972 (N_9972,N_2293,N_3515);
and U9973 (N_9973,N_296,N_4049);
nor U9974 (N_9974,N_235,N_4224);
nor U9975 (N_9975,N_688,N_1352);
xor U9976 (N_9976,N_298,N_323);
and U9977 (N_9977,N_4766,N_2726);
nor U9978 (N_9978,N_0,N_375);
xor U9979 (N_9979,N_2628,N_2135);
xor U9980 (N_9980,N_1362,N_1144);
nand U9981 (N_9981,N_3279,N_3405);
xor U9982 (N_9982,N_3946,N_4725);
nor U9983 (N_9983,N_4526,N_1834);
or U9984 (N_9984,N_3443,N_3233);
nor U9985 (N_9985,N_1114,N_915);
or U9986 (N_9986,N_1784,N_4503);
xnor U9987 (N_9987,N_2777,N_1273);
or U9988 (N_9988,N_195,N_1493);
and U9989 (N_9989,N_3973,N_3083);
or U9990 (N_9990,N_3046,N_2296);
nor U9991 (N_9991,N_163,N_1548);
nand U9992 (N_9992,N_2792,N_1880);
nand U9993 (N_9993,N_1151,N_3311);
or U9994 (N_9994,N_4274,N_2403);
xor U9995 (N_9995,N_1901,N_4855);
nor U9996 (N_9996,N_707,N_4194);
nor U9997 (N_9997,N_3751,N_1489);
or U9998 (N_9998,N_2503,N_680);
nor U9999 (N_9999,N_2536,N_3369);
and U10000 (N_10000,N_6612,N_7455);
nand U10001 (N_10001,N_7708,N_7937);
xor U10002 (N_10002,N_6787,N_7269);
and U10003 (N_10003,N_9302,N_6890);
or U10004 (N_10004,N_8315,N_5189);
nor U10005 (N_10005,N_8799,N_7390);
and U10006 (N_10006,N_9341,N_5835);
nor U10007 (N_10007,N_6798,N_6386);
or U10008 (N_10008,N_8027,N_8192);
or U10009 (N_10009,N_8493,N_9046);
or U10010 (N_10010,N_7252,N_9343);
or U10011 (N_10011,N_8890,N_9154);
and U10012 (N_10012,N_7572,N_5433);
and U10013 (N_10013,N_8109,N_6791);
or U10014 (N_10014,N_8767,N_5174);
and U10015 (N_10015,N_5507,N_5371);
or U10016 (N_10016,N_5150,N_5532);
nand U10017 (N_10017,N_7313,N_8569);
and U10018 (N_10018,N_5916,N_7817);
and U10019 (N_10019,N_6194,N_9015);
or U10020 (N_10020,N_6807,N_5207);
or U10021 (N_10021,N_9811,N_7635);
or U10022 (N_10022,N_8586,N_8445);
nor U10023 (N_10023,N_6792,N_5938);
nand U10024 (N_10024,N_7767,N_5977);
or U10025 (N_10025,N_7992,N_7470);
xor U10026 (N_10026,N_9573,N_7758);
nor U10027 (N_10027,N_8984,N_8936);
xor U10028 (N_10028,N_6972,N_8159);
and U10029 (N_10029,N_7122,N_7051);
nand U10030 (N_10030,N_9394,N_9178);
or U10031 (N_10031,N_8145,N_9685);
and U10032 (N_10032,N_5588,N_9859);
or U10033 (N_10033,N_5432,N_9952);
nand U10034 (N_10034,N_9171,N_7245);
nand U10035 (N_10035,N_9540,N_6647);
and U10036 (N_10036,N_6493,N_8536);
and U10037 (N_10037,N_8419,N_9554);
xnor U10038 (N_10038,N_5165,N_9894);
or U10039 (N_10039,N_7955,N_8979);
or U10040 (N_10040,N_8089,N_8047);
or U10041 (N_10041,N_9215,N_9626);
nor U10042 (N_10042,N_5267,N_5701);
xor U10043 (N_10043,N_8637,N_5519);
xnor U10044 (N_10044,N_7536,N_5358);
xnor U10045 (N_10045,N_9909,N_7238);
xor U10046 (N_10046,N_9580,N_6070);
nand U10047 (N_10047,N_5461,N_9333);
or U10048 (N_10048,N_9442,N_7739);
or U10049 (N_10049,N_8189,N_5661);
nand U10050 (N_10050,N_8584,N_7186);
nor U10051 (N_10051,N_7532,N_7451);
nand U10052 (N_10052,N_5338,N_7383);
xnor U10053 (N_10053,N_7369,N_5065);
xor U10054 (N_10054,N_7466,N_6433);
or U10055 (N_10055,N_6492,N_8059);
xnor U10056 (N_10056,N_9972,N_5126);
or U10057 (N_10057,N_9831,N_9793);
or U10058 (N_10058,N_5648,N_6764);
or U10059 (N_10059,N_5868,N_8300);
nor U10060 (N_10060,N_7454,N_9471);
nor U10061 (N_10061,N_7449,N_9487);
and U10062 (N_10062,N_8770,N_5955);
or U10063 (N_10063,N_9574,N_7934);
and U10064 (N_10064,N_5687,N_7240);
nand U10065 (N_10065,N_5000,N_5720);
nor U10066 (N_10066,N_7611,N_7738);
xor U10067 (N_10067,N_7358,N_5344);
nand U10068 (N_10068,N_5986,N_8093);
and U10069 (N_10069,N_7113,N_6131);
nor U10070 (N_10070,N_8039,N_8313);
and U10071 (N_10071,N_7669,N_8910);
xnor U10072 (N_10072,N_7634,N_9469);
xor U10073 (N_10073,N_6412,N_6626);
nor U10074 (N_10074,N_6494,N_7178);
nand U10075 (N_10075,N_7018,N_5926);
nor U10076 (N_10076,N_8169,N_6738);
nand U10077 (N_10077,N_6533,N_8121);
or U10078 (N_10078,N_5812,N_8128);
nand U10079 (N_10079,N_8641,N_6047);
or U10080 (N_10080,N_9322,N_7056);
nor U10081 (N_10081,N_8748,N_8015);
or U10082 (N_10082,N_6835,N_7980);
xnor U10083 (N_10083,N_8807,N_7082);
and U10084 (N_10084,N_7216,N_9695);
and U10085 (N_10085,N_9130,N_9364);
nand U10086 (N_10086,N_9990,N_5998);
nor U10087 (N_10087,N_9851,N_7865);
and U10088 (N_10088,N_5345,N_7479);
xnor U10089 (N_10089,N_6713,N_7893);
xor U10090 (N_10090,N_5272,N_8593);
nor U10091 (N_10091,N_7165,N_5269);
and U10092 (N_10092,N_7914,N_7655);
xnor U10093 (N_10093,N_5503,N_9681);
or U10094 (N_10094,N_9604,N_9133);
and U10095 (N_10095,N_9558,N_6260);
nand U10096 (N_10096,N_9782,N_5427);
xor U10097 (N_10097,N_5993,N_5699);
nand U10098 (N_10098,N_7671,N_8787);
xnor U10099 (N_10099,N_8363,N_5036);
and U10100 (N_10100,N_9423,N_5747);
xor U10101 (N_10101,N_9643,N_6368);
and U10102 (N_10102,N_5458,N_6023);
nand U10103 (N_10103,N_8268,N_8706);
nand U10104 (N_10104,N_6853,N_5192);
xnor U10105 (N_10105,N_8395,N_9294);
xnor U10106 (N_10106,N_9629,N_9867);
nor U10107 (N_10107,N_7291,N_9662);
xnor U10108 (N_10108,N_8620,N_8307);
or U10109 (N_10109,N_7920,N_6134);
xnor U10110 (N_10110,N_8398,N_7345);
xor U10111 (N_10111,N_6629,N_5195);
and U10112 (N_10112,N_5513,N_5003);
xor U10113 (N_10113,N_6042,N_8446);
nand U10114 (N_10114,N_7840,N_8610);
and U10115 (N_10115,N_6037,N_6689);
nand U10116 (N_10116,N_5653,N_8800);
nor U10117 (N_10117,N_6693,N_8777);
and U10118 (N_10118,N_8980,N_9837);
or U10119 (N_10119,N_5869,N_5575);
or U10120 (N_10120,N_5329,N_5078);
or U10121 (N_10121,N_6151,N_8238);
nand U10122 (N_10122,N_9823,N_5956);
nand U10123 (N_10123,N_5657,N_7828);
and U10124 (N_10124,N_7166,N_7521);
nor U10125 (N_10125,N_7347,N_8476);
xnor U10126 (N_10126,N_5792,N_5999);
nand U10127 (N_10127,N_8505,N_6739);
and U10128 (N_10128,N_6348,N_6053);
or U10129 (N_10129,N_8467,N_6487);
xnor U10130 (N_10130,N_5819,N_7206);
nand U10131 (N_10131,N_7901,N_9435);
nand U10132 (N_10132,N_8306,N_5350);
nor U10133 (N_10133,N_6586,N_9739);
and U10134 (N_10134,N_8549,N_6676);
and U10135 (N_10135,N_8104,N_9158);
and U10136 (N_10136,N_9609,N_7499);
xor U10137 (N_10137,N_6050,N_9798);
nor U10138 (N_10138,N_8064,N_9977);
nor U10139 (N_10139,N_9592,N_8209);
nand U10140 (N_10140,N_6414,N_8905);
xor U10141 (N_10141,N_7031,N_8289);
nand U10142 (N_10142,N_6589,N_5054);
and U10143 (N_10143,N_9856,N_6341);
nor U10144 (N_10144,N_6927,N_5316);
xor U10145 (N_10145,N_9680,N_8858);
xor U10146 (N_10146,N_9637,N_8625);
and U10147 (N_10147,N_6902,N_9671);
xor U10148 (N_10148,N_9264,N_6240);
nand U10149 (N_10149,N_9624,N_9450);
and U10150 (N_10150,N_8718,N_8599);
nand U10151 (N_10151,N_8119,N_7411);
and U10152 (N_10152,N_9970,N_6737);
nand U10153 (N_10153,N_8551,N_6674);
xnor U10154 (N_10154,N_9594,N_5216);
nand U10155 (N_10155,N_9188,N_7385);
xnor U10156 (N_10156,N_6219,N_6865);
or U10157 (N_10157,N_5063,N_8733);
and U10158 (N_10158,N_8875,N_7157);
and U10159 (N_10159,N_6954,N_7613);
and U10160 (N_10160,N_6376,N_6499);
nor U10161 (N_10161,N_5965,N_6292);
and U10162 (N_10162,N_9813,N_9221);
nand U10163 (N_10163,N_7748,N_9845);
or U10164 (N_10164,N_7373,N_7300);
nand U10165 (N_10165,N_7881,N_5487);
or U10166 (N_10166,N_7853,N_7978);
and U10167 (N_10167,N_9848,N_6572);
or U10168 (N_10168,N_7052,N_9721);
xor U10169 (N_10169,N_6277,N_7426);
and U10170 (N_10170,N_5277,N_7107);
or U10171 (N_10171,N_7101,N_7441);
nand U10172 (N_10172,N_8686,N_6296);
nand U10173 (N_10173,N_9863,N_6583);
and U10174 (N_10174,N_6382,N_6684);
or U10175 (N_10175,N_9974,N_6011);
or U10176 (N_10176,N_6671,N_5688);
nor U10177 (N_10177,N_6052,N_8992);
nand U10178 (N_10178,N_8491,N_5136);
or U10179 (N_10179,N_5061,N_6261);
nor U10180 (N_10180,N_7714,N_9765);
nand U10181 (N_10181,N_5450,N_6093);
or U10182 (N_10182,N_5582,N_7020);
or U10183 (N_10183,N_7394,N_8006);
xor U10184 (N_10184,N_8811,N_5927);
nor U10185 (N_10185,N_7519,N_7477);
nor U10186 (N_10186,N_6478,N_8785);
nand U10187 (N_10187,N_9076,N_6518);
xor U10188 (N_10188,N_9193,N_5408);
nor U10189 (N_10189,N_7340,N_8069);
and U10190 (N_10190,N_7808,N_6621);
nand U10191 (N_10191,N_6112,N_8283);
and U10192 (N_10192,N_7179,N_6138);
xnor U10193 (N_10193,N_9224,N_5900);
nand U10194 (N_10194,N_7006,N_8911);
or U10195 (N_10195,N_5012,N_9225);
nand U10196 (N_10196,N_6966,N_5611);
xor U10197 (N_10197,N_8801,N_6654);
and U10198 (N_10198,N_8776,N_8458);
nor U10199 (N_10199,N_7067,N_7354);
nand U10200 (N_10200,N_5415,N_5028);
and U10201 (N_10201,N_9049,N_5883);
and U10202 (N_10202,N_9960,N_9752);
or U10203 (N_10203,N_5183,N_6646);
xor U10204 (N_10204,N_9289,N_7585);
xnor U10205 (N_10205,N_7303,N_7977);
nor U10206 (N_10206,N_6982,N_6658);
and U10207 (N_10207,N_6127,N_8893);
xnor U10208 (N_10208,N_8110,N_8346);
and U10209 (N_10209,N_9281,N_6440);
nand U10210 (N_10210,N_6722,N_8316);
nor U10211 (N_10211,N_7173,N_5631);
or U10212 (N_10212,N_8070,N_5206);
xor U10213 (N_10213,N_5780,N_8614);
nand U10214 (N_10214,N_9879,N_7400);
xnor U10215 (N_10215,N_6400,N_7017);
or U10216 (N_10216,N_5009,N_8929);
nand U10217 (N_10217,N_9925,N_6020);
nand U10218 (N_10218,N_5590,N_8634);
xnor U10219 (N_10219,N_8161,N_9598);
and U10220 (N_10220,N_5475,N_8691);
nand U10221 (N_10221,N_9611,N_5262);
xor U10222 (N_10222,N_6229,N_6098);
or U10223 (N_10223,N_7744,N_6455);
or U10224 (N_10224,N_9452,N_5055);
and U10225 (N_10225,N_5242,N_5710);
or U10226 (N_10226,N_8966,N_7794);
xor U10227 (N_10227,N_5765,N_9503);
nand U10228 (N_10228,N_9597,N_8367);
or U10229 (N_10229,N_6078,N_6209);
and U10230 (N_10230,N_6895,N_6504);
and U10231 (N_10231,N_7849,N_5423);
nand U10232 (N_10232,N_8741,N_7311);
nand U10233 (N_10233,N_7594,N_6636);
or U10234 (N_10234,N_7612,N_5705);
xnor U10235 (N_10235,N_6265,N_5325);
nor U10236 (N_10236,N_8232,N_5299);
or U10237 (N_10237,N_6177,N_5011);
nand U10238 (N_10238,N_5978,N_5296);
or U10239 (N_10239,N_9987,N_8642);
xor U10240 (N_10240,N_9185,N_5846);
or U10241 (N_10241,N_5894,N_6210);
xor U10242 (N_10242,N_5839,N_5075);
or U10243 (N_10243,N_9141,N_7185);
nor U10244 (N_10244,N_8378,N_8387);
or U10245 (N_10245,N_6014,N_5084);
nor U10246 (N_10246,N_7388,N_6863);
nand U10247 (N_10247,N_8612,N_6809);
xor U10248 (N_10248,N_6017,N_5693);
xor U10249 (N_10249,N_8023,N_9267);
or U10250 (N_10250,N_9904,N_8223);
xnor U10251 (N_10251,N_7484,N_6514);
xor U10252 (N_10252,N_6378,N_9169);
or U10253 (N_10253,N_7312,N_5604);
nor U10254 (N_10254,N_8727,N_6900);
nand U10255 (N_10255,N_5505,N_9490);
or U10256 (N_10256,N_8298,N_9696);
nand U10257 (N_10257,N_8848,N_9905);
nor U10258 (N_10258,N_8564,N_6875);
or U10259 (N_10259,N_8738,N_9128);
xor U10260 (N_10260,N_7771,N_8225);
or U10261 (N_10261,N_5334,N_9432);
or U10262 (N_10262,N_8680,N_9989);
or U10263 (N_10263,N_8894,N_9144);
nand U10264 (N_10264,N_7352,N_8348);
xor U10265 (N_10265,N_7030,N_5392);
and U10266 (N_10266,N_6384,N_9004);
xor U10267 (N_10267,N_6105,N_8291);
nor U10268 (N_10268,N_7827,N_6590);
or U10269 (N_10269,N_8388,N_8420);
or U10270 (N_10270,N_7951,N_9196);
xor U10271 (N_10271,N_5319,N_9483);
nor U10272 (N_10272,N_7599,N_7085);
xor U10273 (N_10273,N_6527,N_9565);
and U10274 (N_10274,N_8186,N_9843);
or U10275 (N_10275,N_9235,N_8560);
or U10276 (N_10276,N_5630,N_5733);
xor U10277 (N_10277,N_7831,N_9918);
xor U10278 (N_10278,N_6959,N_9967);
xnor U10279 (N_10279,N_5464,N_6565);
and U10280 (N_10280,N_5741,N_9043);
and U10281 (N_10281,N_5952,N_9242);
or U10282 (N_10282,N_5179,N_8945);
nor U10283 (N_10283,N_9395,N_6948);
nor U10284 (N_10284,N_7142,N_8917);
or U10285 (N_10285,N_5259,N_7545);
or U10286 (N_10286,N_6641,N_8390);
nand U10287 (N_10287,N_8834,N_9104);
and U10288 (N_10288,N_9650,N_5173);
and U10289 (N_10289,N_9167,N_8502);
and U10290 (N_10290,N_7452,N_6842);
and U10291 (N_10291,N_9430,N_6735);
xnor U10292 (N_10292,N_9468,N_6611);
and U10293 (N_10293,N_5468,N_8961);
xor U10294 (N_10294,N_6907,N_6197);
and U10295 (N_10295,N_9148,N_5832);
nand U10296 (N_10296,N_7284,N_9189);
nor U10297 (N_10297,N_9922,N_9186);
xor U10298 (N_10298,N_6387,N_8026);
xor U10299 (N_10299,N_8521,N_7327);
or U10300 (N_10300,N_5945,N_7762);
and U10301 (N_10301,N_5558,N_8604);
and U10302 (N_10302,N_8255,N_9805);
xor U10303 (N_10303,N_5915,N_9942);
and U10304 (N_10304,N_9214,N_5625);
and U10305 (N_10305,N_6221,N_7250);
xor U10306 (N_10306,N_5095,N_8662);
xnor U10307 (N_10307,N_5904,N_7190);
nor U10308 (N_10308,N_6161,N_7026);
or U10309 (N_10309,N_5947,N_5390);
and U10310 (N_10310,N_9438,N_9481);
and U10311 (N_10311,N_5535,N_9460);
and U10312 (N_10312,N_8566,N_5434);
or U10313 (N_10313,N_7633,N_5542);
or U10314 (N_10314,N_9033,N_9710);
or U10315 (N_10315,N_5237,N_6508);
xor U10316 (N_10316,N_5265,N_8772);
xnor U10317 (N_10317,N_7834,N_5837);
nor U10318 (N_10318,N_5606,N_9220);
xor U10319 (N_10319,N_7604,N_9852);
or U10320 (N_10320,N_5762,N_9377);
nand U10321 (N_10321,N_8364,N_5031);
nor U10322 (N_10322,N_8784,N_6095);
xor U10323 (N_10323,N_9243,N_7077);
and U10324 (N_10324,N_7387,N_5902);
nor U10325 (N_10325,N_6822,N_5293);
nor U10326 (N_10326,N_8631,N_9497);
or U10327 (N_10327,N_5896,N_5218);
nor U10328 (N_10328,N_5895,N_9374);
nor U10329 (N_10329,N_8728,N_6289);
xnor U10330 (N_10330,N_9314,N_6019);
xnor U10331 (N_10331,N_5933,N_6018);
or U10332 (N_10332,N_5983,N_9495);
xor U10333 (N_10333,N_6769,N_7010);
and U10334 (N_10334,N_5671,N_5781);
nor U10335 (N_10335,N_9253,N_8783);
nand U10336 (N_10336,N_7653,N_9090);
and U10337 (N_10337,N_5928,N_9795);
xor U10338 (N_10338,N_5320,N_7458);
nand U10339 (N_10339,N_8941,N_6402);
xnor U10340 (N_10340,N_6274,N_8515);
xnor U10341 (N_10341,N_6709,N_7571);
or U10342 (N_10342,N_5827,N_9032);
and U10343 (N_10343,N_6136,N_9953);
and U10344 (N_10344,N_6354,N_8163);
or U10345 (N_10345,N_5892,N_7508);
and U10346 (N_10346,N_8361,N_5806);
nor U10347 (N_10347,N_5641,N_8466);
nand U10348 (N_10348,N_6649,N_9808);
nand U10349 (N_10349,N_9719,N_6215);
or U10350 (N_10350,N_6771,N_9262);
xnor U10351 (N_10351,N_9628,N_9962);
and U10352 (N_10352,N_9916,N_7880);
and U10353 (N_10353,N_6252,N_5992);
nand U10354 (N_10354,N_7086,N_9998);
nor U10355 (N_10355,N_6068,N_9037);
xnor U10356 (N_10356,N_5644,N_6313);
nor U10357 (N_10357,N_5351,N_8946);
and U10358 (N_10358,N_8274,N_6846);
and U10359 (N_10359,N_5520,N_6638);
nor U10360 (N_10360,N_9008,N_9238);
or U10361 (N_10361,N_9071,N_8176);
nand U10362 (N_10362,N_9286,N_7861);
xor U10363 (N_10363,N_7877,N_7209);
or U10364 (N_10364,N_7450,N_7089);
or U10365 (N_10365,N_5348,N_7679);
nor U10366 (N_10366,N_6377,N_7218);
xnor U10367 (N_10367,N_6760,N_7770);
xor U10368 (N_10368,N_7236,N_5950);
nand U10369 (N_10369,N_7862,N_6468);
nand U10370 (N_10370,N_7887,N_9526);
xnor U10371 (N_10371,N_5960,N_6743);
nand U10372 (N_10372,N_9191,N_9511);
nand U10373 (N_10373,N_5953,N_6434);
xor U10374 (N_10374,N_5457,N_7732);
or U10375 (N_10375,N_8165,N_5431);
and U10376 (N_10376,N_9280,N_6423);
nand U10377 (N_10377,N_6765,N_9480);
nor U10378 (N_10378,N_5473,N_8889);
xnor U10379 (N_10379,N_6775,N_7562);
xnor U10380 (N_10380,N_8253,N_6507);
xnor U10381 (N_10381,N_9445,N_6845);
nor U10382 (N_10382,N_6168,N_9521);
xor U10383 (N_10383,N_5280,N_8791);
and U10384 (N_10384,N_8724,N_5514);
and U10385 (N_10385,N_6861,N_7971);
nor U10386 (N_10386,N_7414,N_9891);
xor U10387 (N_10387,N_6135,N_5559);
xor U10388 (N_10388,N_9986,N_7445);
or U10389 (N_10389,N_5860,N_6146);
or U10390 (N_10390,N_7988,N_7210);
or U10391 (N_10391,N_6352,N_6406);
nand U10392 (N_10392,N_8843,N_8948);
xnor U10393 (N_10393,N_6594,N_8456);
nand U10394 (N_10394,N_5180,N_8734);
xor U10395 (N_10395,N_6970,N_9202);
nand U10396 (N_10396,N_5776,N_9530);
nor U10397 (N_10397,N_8494,N_6027);
xor U10398 (N_10398,N_9176,N_7592);
xnor U10399 (N_10399,N_8661,N_6981);
or U10400 (N_10400,N_9951,N_7682);
and U10401 (N_10401,N_6272,N_5290);
or U10402 (N_10402,N_5186,N_7034);
nand U10403 (N_10403,N_9621,N_7343);
nand U10404 (N_10404,N_7167,N_7005);
and U10405 (N_10405,N_9386,N_6830);
xor U10406 (N_10406,N_8341,N_5638);
nand U10407 (N_10407,N_9051,N_6322);
nand U10408 (N_10408,N_6685,N_7697);
nor U10409 (N_10409,N_8603,N_8831);
nand U10410 (N_10410,N_8107,N_9689);
nor U10411 (N_10411,N_8191,N_5021);
nand U10412 (N_10412,N_6998,N_9372);
nor U10413 (N_10413,N_9486,N_5110);
or U10414 (N_10414,N_6388,N_7324);
or U10415 (N_10415,N_6033,N_9534);
and U10416 (N_10416,N_9712,N_7700);
or U10417 (N_10417,N_9682,N_9042);
xor U10418 (N_10418,N_7069,N_6064);
nand U10419 (N_10419,N_9964,N_5069);
and U10420 (N_10420,N_5633,N_9160);
xor U10421 (N_10421,N_8439,N_7513);
xnor U10422 (N_10422,N_7919,N_6497);
or U10423 (N_10423,N_8938,N_7693);
or U10424 (N_10424,N_8160,N_9647);
xor U10425 (N_10425,N_6208,N_9906);
or U10426 (N_10426,N_6779,N_8447);
and U10427 (N_10427,N_8927,N_6453);
and U10428 (N_10428,N_8489,N_9840);
nand U10429 (N_10429,N_6385,N_5106);
nor U10430 (N_10430,N_7106,N_7362);
xor U10431 (N_10431,N_7743,N_5330);
xor U10432 (N_10432,N_9866,N_7856);
nor U10433 (N_10433,N_5147,N_9587);
nand U10434 (N_10434,N_7836,N_5988);
nor U10435 (N_10435,N_8973,N_9885);
and U10436 (N_10436,N_7678,N_5990);
xnor U10437 (N_10437,N_9640,N_5964);
nor U10438 (N_10438,N_9874,N_8652);
or U10439 (N_10439,N_6852,N_7436);
xor U10440 (N_10440,N_5997,N_5362);
or U10441 (N_10441,N_5292,N_6872);
or U10442 (N_10442,N_7683,N_5703);
nor U10443 (N_10443,N_6443,N_9287);
xor U10444 (N_10444,N_7108,N_5248);
nor U10445 (N_10445,N_6338,N_9389);
and U10446 (N_10446,N_8233,N_9600);
or U10447 (N_10447,N_6543,N_8276);
nand U10448 (N_10448,N_7263,N_9896);
nor U10449 (N_10449,N_6608,N_9822);
nand U10450 (N_10450,N_8953,N_8919);
and U10451 (N_10451,N_9608,N_9409);
nand U10452 (N_10452,N_7422,N_6333);
and U10453 (N_10453,N_6949,N_5629);
and U10454 (N_10454,N_8437,N_7197);
and U10455 (N_10455,N_6169,N_8162);
nand U10456 (N_10456,N_9993,N_5496);
and U10457 (N_10457,N_9672,N_9550);
or U10458 (N_10458,N_5056,N_5568);
xor U10459 (N_10459,N_6263,N_5082);
or U10460 (N_10460,N_7591,N_7336);
or U10461 (N_10461,N_7493,N_9402);
or U10462 (N_10462,N_6202,N_9946);
nand U10463 (N_10463,N_6396,N_7995);
and U10464 (N_10464,N_6206,N_6575);
nand U10465 (N_10465,N_8256,N_7412);
xor U10466 (N_10466,N_6314,N_7550);
and U10467 (N_10467,N_7879,N_9125);
and U10468 (N_10468,N_9161,N_5281);
nand U10469 (N_10469,N_5306,N_5470);
nor U10470 (N_10470,N_5111,N_6938);
xor U10471 (N_10471,N_8018,N_5359);
nor U10472 (N_10472,N_9783,N_9317);
nand U10473 (N_10473,N_9115,N_5261);
or U10474 (N_10474,N_6650,N_6803);
and U10475 (N_10475,N_9746,N_8669);
or U10476 (N_10476,N_9664,N_9010);
and U10477 (N_10477,N_7651,N_7801);
xnor U10478 (N_10478,N_9111,N_9505);
xnor U10479 (N_10479,N_8750,N_8281);
and U10480 (N_10480,N_7766,N_9387);
nand U10481 (N_10481,N_7009,N_6726);
nor U10482 (N_10482,N_6489,N_8898);
nand U10483 (N_10483,N_8947,N_5282);
xnor U10484 (N_10484,N_8383,N_9216);
or U10485 (N_10485,N_5845,N_9126);
nand U10486 (N_10486,N_6164,N_5074);
xnor U10487 (N_10487,N_9052,N_6606);
and U10488 (N_10488,N_9023,N_8579);
and U10489 (N_10489,N_8832,N_6288);
or U10490 (N_10490,N_6355,N_9239);
or U10491 (N_10491,N_8019,N_8257);
xor U10492 (N_10492,N_7259,N_6308);
or U10493 (N_10493,N_6906,N_7755);
or U10494 (N_10494,N_9212,N_7268);
or U10495 (N_10495,N_8701,N_9441);
or U10496 (N_10496,N_6082,N_6061);
or U10497 (N_10497,N_9641,N_9602);
or U10498 (N_10498,N_9902,N_6069);
or U10499 (N_10499,N_7799,N_8155);
and U10500 (N_10500,N_6926,N_6117);
nor U10501 (N_10501,N_8366,N_9496);
or U10502 (N_10502,N_7650,N_6717);
nand U10503 (N_10503,N_7658,N_8958);
or U10504 (N_10504,N_9062,N_9258);
nand U10505 (N_10505,N_6516,N_7731);
xor U10506 (N_10506,N_6266,N_5726);
and U10507 (N_10507,N_6451,N_9864);
nand U10508 (N_10508,N_8968,N_8380);
xor U10509 (N_10509,N_9996,N_8406);
nor U10510 (N_10510,N_6987,N_5969);
or U10511 (N_10511,N_9649,N_6075);
or U10512 (N_10512,N_7746,N_6413);
xnor U10513 (N_10513,N_6975,N_8804);
and U10514 (N_10514,N_8099,N_5763);
or U10515 (N_10515,N_7180,N_7673);
nor U10516 (N_10516,N_6235,N_7695);
and U10517 (N_10517,N_8697,N_6609);
nor U10518 (N_10518,N_7320,N_9344);
xnor U10519 (N_10519,N_7686,N_7636);
and U10520 (N_10520,N_5044,N_8060);
and U10521 (N_10521,N_8971,N_9777);
or U10522 (N_10522,N_9701,N_9679);
nand U10523 (N_10523,N_6564,N_5833);
or U10524 (N_10524,N_8972,N_7644);
nand U10525 (N_10525,N_6299,N_8550);
nand U10526 (N_10526,N_9311,N_5096);
nand U10527 (N_10527,N_9581,N_7765);
nor U10528 (N_10528,N_6567,N_5053);
xor U10529 (N_10529,N_5424,N_7567);
xnor U10530 (N_10530,N_6298,N_8700);
nand U10531 (N_10531,N_5029,N_9447);
nand U10532 (N_10532,N_8759,N_5683);
nor U10533 (N_10533,N_8114,N_5783);
or U10534 (N_10534,N_6311,N_9862);
xor U10535 (N_10535,N_5639,N_5305);
nor U10536 (N_10536,N_8106,N_9532);
nand U10537 (N_10537,N_8517,N_7864);
or U10538 (N_10538,N_8371,N_8925);
and U10539 (N_10539,N_9226,N_9200);
nor U10540 (N_10540,N_9814,N_5903);
nor U10541 (N_10541,N_6997,N_8818);
xor U10542 (N_10542,N_8934,N_6408);
xnor U10543 (N_10543,N_9217,N_6502);
and U10544 (N_10544,N_5241,N_8085);
and U10545 (N_10545,N_6063,N_7293);
and U10546 (N_10546,N_9801,N_8224);
xor U10547 (N_10547,N_7022,N_5740);
xnor U10548 (N_10548,N_9375,N_6869);
nand U10549 (N_10549,N_9120,N_7846);
nand U10550 (N_10550,N_9729,N_7566);
nand U10551 (N_10551,N_6476,N_5899);
nand U10552 (N_10552,N_6896,N_9523);
or U10553 (N_10553,N_7378,N_8506);
nor U10554 (N_10554,N_9557,N_8824);
or U10555 (N_10555,N_5596,N_7384);
or U10556 (N_10556,N_5877,N_7858);
xnor U10557 (N_10557,N_7734,N_6932);
and U10558 (N_10558,N_7013,N_5574);
and U10559 (N_10559,N_5419,N_5660);
and U10560 (N_10560,N_6864,N_9228);
and U10561 (N_10561,N_8646,N_8487);
or U10562 (N_10562,N_7570,N_9183);
nor U10563 (N_10563,N_6255,N_9948);
xor U10564 (N_10564,N_8563,N_5249);
nor U10565 (N_10565,N_6871,N_6983);
or U10566 (N_10566,N_7672,N_6617);
xnor U10567 (N_10567,N_8763,N_9779);
nand U10568 (N_10568,N_5737,N_5337);
nor U10569 (N_10569,N_8613,N_5561);
xor U10570 (N_10570,N_7249,N_5219);
and U10571 (N_10571,N_8782,N_5579);
nor U10572 (N_10572,N_7265,N_6933);
nor U10573 (N_10573,N_7943,N_6025);
and U10574 (N_10574,N_6544,N_6915);
and U10575 (N_10575,N_6262,N_9254);
nor U10576 (N_10576,N_9316,N_9418);
nand U10577 (N_10577,N_5815,N_5250);
and U10578 (N_10578,N_8384,N_6513);
nor U10579 (N_10579,N_9378,N_9923);
or U10580 (N_10580,N_9473,N_9871);
xor U10581 (N_10581,N_6046,N_7397);
and U10582 (N_10582,N_7274,N_7956);
xor U10583 (N_10583,N_5948,N_5210);
nor U10584 (N_10584,N_9061,N_8974);
nand U10585 (N_10585,N_6913,N_5906);
nand U10586 (N_10586,N_9045,N_6154);
or U10587 (N_10587,N_7898,N_6256);
nand U10588 (N_10588,N_9002,N_6885);
or U10589 (N_10589,N_6305,N_5805);
nor U10590 (N_10590,N_6422,N_7927);
xor U10591 (N_10591,N_6304,N_6245);
and U10592 (N_10592,N_5322,N_6883);
nand U10593 (N_10593,N_5205,N_5848);
nor U10594 (N_10594,N_7174,N_5546);
nor U10595 (N_10595,N_8338,N_8053);
and U10596 (N_10596,N_9198,N_5238);
nor U10597 (N_10597,N_6373,N_7684);
xor U10598 (N_10598,N_7928,N_5402);
nor U10599 (N_10599,N_8617,N_9583);
xnor U10600 (N_10600,N_6142,N_5794);
nor U10601 (N_10601,N_9553,N_5381);
and U10602 (N_10602,N_9307,N_6062);
xnor U10603 (N_10603,N_7407,N_8479);
nor U10604 (N_10604,N_8731,N_5672);
or U10605 (N_10605,N_5771,N_5156);
or U10606 (N_10606,N_9152,N_9544);
and U10607 (N_10607,N_8351,N_7478);
xor U10608 (N_10608,N_7033,N_7440);
nand U10609 (N_10609,N_6699,N_8722);
or U10610 (N_10610,N_9119,N_7504);
nand U10611 (N_10611,N_6397,N_5972);
or U10612 (N_10612,N_6519,N_9778);
nand U10613 (N_10613,N_9610,N_7626);
nand U10614 (N_10614,N_5247,N_8547);
xnor U10615 (N_10615,N_6889,N_5668);
xnor U10616 (N_10616,N_5254,N_6401);
and U10617 (N_10617,N_7952,N_8305);
nor U10618 (N_10618,N_9363,N_5033);
nand U10619 (N_10619,N_8758,N_5941);
nand U10620 (N_10620,N_5049,N_9142);
xnor U10621 (N_10621,N_5439,N_5550);
and U10622 (N_10622,N_6613,N_7229);
or U10623 (N_10623,N_8535,N_6149);
xor U10624 (N_10624,N_5816,N_5062);
or U10625 (N_10625,N_8336,N_7147);
or U10626 (N_10626,N_5343,N_7102);
and U10627 (N_10627,N_6480,N_8385);
nor U10628 (N_10628,N_7172,N_9282);
xnor U10629 (N_10629,N_5711,N_9293);
nor U10630 (N_10630,N_9563,N_8666);
nor U10631 (N_10631,N_7524,N_6772);
xor U10632 (N_10632,N_9757,N_6556);
or U10633 (N_10633,N_9113,N_8649);
nor U10634 (N_10634,N_5526,N_7989);
xnor U10635 (N_10635,N_5996,N_8086);
nand U10636 (N_10636,N_8624,N_6270);
xor U10637 (N_10637,N_9535,N_8326);
and U10638 (N_10638,N_8344,N_9937);
or U10639 (N_10639,N_9659,N_8484);
nand U10640 (N_10640,N_5152,N_8193);
nor U10641 (N_10641,N_8863,N_9295);
nand U10642 (N_10642,N_5212,N_6343);
nand U10643 (N_10643,N_8149,N_9846);
or U10644 (N_10644,N_7170,N_6976);
xnor U10645 (N_10645,N_9485,N_6774);
or U10646 (N_10646,N_8538,N_5889);
nor U10647 (N_10647,N_9181,N_5321);
xor U10648 (N_10648,N_6327,N_6411);
nor U10649 (N_10649,N_5962,N_9950);
and U10650 (N_10650,N_9519,N_8869);
nand U10651 (N_10651,N_7616,N_6424);
or U10652 (N_10652,N_5522,N_8333);
and U10653 (N_10653,N_6351,N_5852);
nor U10654 (N_10654,N_9278,N_7539);
nand U10655 (N_10655,N_7593,N_5438);
or U10656 (N_10656,N_7181,N_5730);
nand U10657 (N_10657,N_9371,N_7699);
or U10658 (N_10658,N_7912,N_7510);
and U10659 (N_10659,N_6701,N_5623);
and U10660 (N_10660,N_8805,N_5445);
xor U10661 (N_10661,N_5336,N_9321);
nand U10662 (N_10662,N_6877,N_9617);
and U10663 (N_10663,N_7812,N_6766);
and U10664 (N_10664,N_6941,N_5052);
xor U10665 (N_10665,N_5166,N_9978);
and U10666 (N_10666,N_7711,N_8391);
xor U10667 (N_10667,N_6284,N_7561);
nor U10668 (N_10668,N_9698,N_5235);
nor U10669 (N_10669,N_5311,N_8857);
nand U10670 (N_10670,N_5626,N_9069);
or U10671 (N_10671,N_9678,N_7317);
and U10672 (N_10672,N_9531,N_9050);
nor U10673 (N_10673,N_6374,N_8623);
nor U10674 (N_10674,N_5379,N_9651);
nand U10675 (N_10675,N_8977,N_9329);
or U10676 (N_10676,N_7742,N_5667);
nor U10677 (N_10677,N_7903,N_8609);
nand U10678 (N_10678,N_5501,N_8229);
nor U10679 (N_10679,N_6920,N_8001);
nand U10680 (N_10680,N_7296,N_5239);
and U10681 (N_10681,N_9320,N_5732);
and U10682 (N_10682,N_6418,N_5177);
nor U10683 (N_10683,N_8498,N_7137);
and U10684 (N_10684,N_6318,N_9203);
or U10685 (N_10685,N_9585,N_5171);
nand U10686 (N_10686,N_6267,N_6681);
or U10687 (N_10687,N_6416,N_7845);
xnor U10688 (N_10688,N_9123,N_9005);
xnor U10689 (N_10689,N_9296,N_5383);
nor U10690 (N_10690,N_9421,N_6486);
and U10691 (N_10691,N_5856,N_5234);
xor U10692 (N_10692,N_7344,N_7404);
xor U10693 (N_10693,N_6107,N_5070);
xor U10694 (N_10694,N_5447,N_6568);
or U10695 (N_10695,N_6868,N_7444);
and U10696 (N_10696,N_7489,N_8567);
and U10697 (N_10697,N_9803,N_6084);
nand U10698 (N_10698,N_7747,N_7638);
and U10699 (N_10699,N_7625,N_5340);
or U10700 (N_10700,N_8810,N_6751);
nand U10701 (N_10701,N_7224,N_9654);
nand U10702 (N_10702,N_7749,N_5676);
nor U10703 (N_10703,N_8931,N_5738);
and U10704 (N_10704,N_9872,N_9959);
or U10705 (N_10705,N_7628,N_7709);
nor U10706 (N_10706,N_6035,N_9173);
and U10707 (N_10707,N_6100,N_9728);
xnor U10708 (N_10708,N_9634,N_5942);
and U10709 (N_10709,N_6758,N_5497);
xnor U10710 (N_10710,N_7917,N_6279);
xor U10711 (N_10711,N_7544,N_7701);
and U10712 (N_10712,N_5728,N_7806);
nand U10713 (N_10713,N_8115,N_8856);
and U10714 (N_10714,N_7223,N_6977);
nand U10715 (N_10715,N_6928,N_9121);
nand U10716 (N_10716,N_8773,N_8066);
xor U10717 (N_10717,N_8354,N_9449);
nor U10718 (N_10718,N_6698,N_7605);
nand U10719 (N_10719,N_8267,N_8113);
and U10720 (N_10720,N_8308,N_9068);
xnor U10721 (N_10721,N_5577,N_9562);
xor U10722 (N_10722,N_9131,N_7289);
and U10723 (N_10723,N_9638,N_9539);
or U10724 (N_10724,N_9163,N_8200);
or U10725 (N_10725,N_7514,N_5678);
and U10726 (N_10726,N_7933,N_7795);
nor U10727 (N_10727,N_5213,N_5570);
xor U10728 (N_10728,N_7964,N_9089);
and U10729 (N_10729,N_9601,N_5744);
or U10730 (N_10730,N_5367,N_7648);
or U10731 (N_10731,N_6032,N_7044);
or U10732 (N_10732,N_5236,N_9330);
or U10733 (N_10733,N_5418,N_9100);
nand U10734 (N_10734,N_6733,N_7787);
xnor U10735 (N_10735,N_8073,N_8814);
or U10736 (N_10736,N_9065,N_6950);
nor U10737 (N_10737,N_5842,N_9802);
xnor U10738 (N_10738,N_8352,N_7065);
nand U10739 (N_10739,N_9096,N_9413);
and U10740 (N_10740,N_7970,N_7437);
nand U10741 (N_10741,N_7431,N_5863);
or U10742 (N_10742,N_9661,N_6767);
and U10743 (N_10743,N_6113,N_5170);
or U10744 (N_10744,N_5328,N_7637);
and U10745 (N_10745,N_7200,N_8347);
xor U10746 (N_10746,N_5163,N_7011);
nor U10747 (N_10747,N_9359,N_9029);
nor U10748 (N_10748,N_8138,N_9136);
nand U10749 (N_10749,N_6239,N_8650);
nor U10750 (N_10750,N_9194,N_7945);
nor U10751 (N_10751,N_8368,N_9011);
nor U10752 (N_10752,N_8534,N_6389);
or U10753 (N_10753,N_9475,N_7012);
nand U10754 (N_10754,N_8990,N_8527);
xnor U10755 (N_10755,N_8516,N_9263);
xor U10756 (N_10756,N_7016,N_9332);
nand U10757 (N_10757,N_7475,N_6850);
xnor U10758 (N_10758,N_5656,N_7822);
xnor U10759 (N_10759,N_5790,N_7242);
or U10760 (N_10760,N_7557,N_5168);
and U10761 (N_10761,N_7133,N_5911);
nor U10762 (N_10762,N_6559,N_8962);
or U10763 (N_10763,N_9512,N_5605);
xor U10764 (N_10764,N_5884,N_7883);
nor U10765 (N_10765,N_7019,N_5417);
and U10766 (N_10766,N_8522,N_7588);
xor U10767 (N_10767,N_7213,N_6483);
xnor U10768 (N_10768,N_6789,N_7506);
or U10769 (N_10769,N_8781,N_6784);
and U10770 (N_10770,N_8852,N_8143);
or U10771 (N_10771,N_7351,N_8845);
xor U10772 (N_10772,N_7888,N_8975);
and U10773 (N_10773,N_6419,N_8993);
nand U10774 (N_10774,N_7380,N_7253);
and U10775 (N_10775,N_8241,N_8587);
and U10776 (N_10776,N_5452,N_9079);
and U10777 (N_10777,N_9092,N_8259);
nor U10778 (N_10778,N_7835,N_8822);
and U10779 (N_10779,N_5025,N_8837);
or U10780 (N_10780,N_7088,N_5893);
nor U10781 (N_10781,N_9352,N_6728);
nor U10782 (N_10782,N_8172,N_8815);
xnor U10783 (N_10783,N_6935,N_5713);
nor U10784 (N_10784,N_5981,N_9809);
nand U10785 (N_10785,N_6282,N_9012);
nand U10786 (N_10786,N_9911,N_7460);
and U10787 (N_10787,N_7642,N_6837);
and U10788 (N_10788,N_5580,N_6663);
nor U10789 (N_10789,N_6734,N_8041);
or U10790 (N_10790,N_6326,N_6417);
nor U10791 (N_10791,N_8696,N_6325);
and U10792 (N_10792,N_8978,N_9179);
or U10793 (N_10793,N_7365,N_9187);
nor U10794 (N_10794,N_9758,N_8250);
nand U10795 (N_10795,N_6329,N_7457);
nand U10796 (N_10796,N_6918,N_6749);
nor U10797 (N_10797,N_9351,N_6457);
and U10798 (N_10798,N_5108,N_9855);
and U10799 (N_10799,N_5677,N_7913);
or U10800 (N_10800,N_6554,N_9819);
nor U10801 (N_10801,N_7090,N_9013);
and U10802 (N_10802,N_9059,N_6704);
or U10803 (N_10803,N_9064,N_9501);
nor U10804 (N_10804,N_5482,N_7528);
or U10805 (N_10805,N_7002,N_7192);
nor U10806 (N_10806,N_7963,N_5498);
nand U10807 (N_10807,N_6021,N_8392);
or U10808 (N_10808,N_6962,N_8422);
nor U10809 (N_10809,N_9889,N_9981);
nand U10810 (N_10810,N_7665,N_9091);
and U10811 (N_10811,N_5050,N_8244);
and U10812 (N_10812,N_7761,N_8749);
nand U10813 (N_10813,N_9472,N_6407);
nand U10814 (N_10814,N_5613,N_8955);
and U10815 (N_10815,N_6573,N_8471);
and U10816 (N_10816,N_5393,N_5256);
nor U10817 (N_10817,N_7676,N_6506);
nand U10818 (N_10818,N_9841,N_6752);
and U10819 (N_10819,N_5557,N_9829);
nand U10820 (N_10820,N_6226,N_8404);
or U10821 (N_10821,N_5339,N_6436);
or U10822 (N_10822,N_7129,N_7471);
or U10823 (N_10823,N_6725,N_7021);
xor U10824 (N_10824,N_8071,N_8098);
or U10825 (N_10825,N_6691,N_7111);
or U10826 (N_10826,N_7418,N_5356);
xnor U10827 (N_10827,N_8939,N_6184);
xor U10828 (N_10828,N_5910,N_7869);
or U10829 (N_10829,N_6952,N_6220);
xor U10830 (N_10830,N_9255,N_9958);
nor U10831 (N_10831,N_8320,N_9861);
nor U10832 (N_10832,N_9555,N_7099);
nor U10833 (N_10833,N_7121,N_5167);
xor U10834 (N_10834,N_6570,N_5485);
nor U10835 (N_10835,N_7750,N_8332);
and U10836 (N_10836,N_9733,N_8709);
nand U10837 (N_10837,N_8578,N_9957);
and U10838 (N_10838,N_6781,N_9516);
and U10839 (N_10839,N_8675,N_5211);
nand U10840 (N_10840,N_6297,N_6546);
or U10841 (N_10841,N_6620,N_8747);
xor U10842 (N_10842,N_8685,N_7270);
and U10843 (N_10843,N_8851,N_5222);
and U10844 (N_10844,N_5886,N_5836);
nor U10845 (N_10845,N_6446,N_9569);
xor U10846 (N_10846,N_9645,N_8216);
or U10847 (N_10847,N_5430,N_5536);
and U10848 (N_10848,N_9510,N_8648);
xnor U10849 (N_10849,N_7979,N_5722);
or U10850 (N_10850,N_8827,N_8139);
xor U10851 (N_10851,N_9939,N_6473);
nor U10852 (N_10852,N_6218,N_7807);
xnor U10853 (N_10853,N_8230,N_8956);
and U10854 (N_10854,N_7821,N_8218);
nand U10855 (N_10855,N_8277,N_5714);
nand U10856 (N_10856,N_5227,N_8896);
nand U10857 (N_10857,N_7389,N_6122);
and U10858 (N_10858,N_5537,N_7729);
nor U10859 (N_10859,N_7892,N_8127);
and U10860 (N_10860,N_7941,N_9443);
xnor U10861 (N_10861,N_5386,N_8739);
nor U10862 (N_10862,N_7215,N_5357);
nand U10863 (N_10863,N_8125,N_6174);
nor U10864 (N_10864,N_8874,N_7386);
or U10865 (N_10865,N_7960,N_5959);
and U10866 (N_10866,N_6395,N_7930);
nor U10867 (N_10867,N_9973,N_8544);
nor U10868 (N_10868,N_6688,N_5490);
nor U10869 (N_10869,N_6827,N_6466);
nor U10870 (N_10870,N_5365,N_5594);
nand U10871 (N_10871,N_8205,N_7670);
and U10872 (N_10872,N_6205,N_7641);
and U10873 (N_10873,N_5276,N_9806);
nand U10874 (N_10874,N_6409,N_9035);
or U10875 (N_10875,N_7294,N_7225);
xor U10876 (N_10876,N_5544,N_9506);
and U10877 (N_10877,N_9482,N_5788);
nor U10878 (N_10878,N_6866,N_8078);
or U10879 (N_10879,N_9812,N_7007);
xor U10880 (N_10880,N_8626,N_9219);
nor U10881 (N_10881,N_6330,N_8438);
xnor U10882 (N_10882,N_5403,N_7302);
or U10883 (N_10883,N_7851,N_8414);
nor U10884 (N_10884,N_8234,N_8682);
or U10885 (N_10885,N_7710,N_5083);
or U10886 (N_10886,N_6182,N_9164);
nor U10887 (N_10887,N_6799,N_6331);
and U10888 (N_10888,N_8142,N_6587);
or U10889 (N_10889,N_8813,N_5861);
or U10890 (N_10890,N_8768,N_5102);
nand U10891 (N_10891,N_6110,N_8401);
xnor U10892 (N_10892,N_8462,N_5370);
nor U10893 (N_10893,N_8683,N_8714);
and U10894 (N_10894,N_6186,N_7949);
nor U10895 (N_10895,N_5042,N_9056);
and U10896 (N_10896,N_8674,N_5731);
nor U10897 (N_10897,N_7353,N_6615);
or U10898 (N_10898,N_5342,N_9529);
or U10899 (N_10899,N_9590,N_8627);
xnor U10900 (N_10900,N_7382,N_5857);
or U10901 (N_10901,N_7290,N_6225);
or U10902 (N_10902,N_9677,N_7523);
nor U10903 (N_10903,N_9034,N_6099);
or U10904 (N_10904,N_6365,N_7171);
nand U10905 (N_10905,N_8657,N_9357);
nor U10906 (N_10906,N_9797,N_9336);
nand U10907 (N_10907,N_9552,N_8058);
xor U10908 (N_10908,N_8492,N_9353);
xor U10909 (N_10909,N_7076,N_9319);
xor U10910 (N_10910,N_9982,N_9842);
xnor U10911 (N_10911,N_7578,N_5968);
or U10912 (N_10912,N_6452,N_8094);
and U10913 (N_10913,N_6085,N_5129);
or U10914 (N_10914,N_9675,N_8157);
nor U10915 (N_10915,N_9030,N_8702);
and U10916 (N_10916,N_5907,N_6757);
or U10917 (N_10917,N_9824,N_8179);
nor U10918 (N_10918,N_7376,N_5184);
nand U10919 (N_10919,N_5966,N_7624);
and U10920 (N_10920,N_6337,N_6783);
xor U10921 (N_10921,N_8989,N_8999);
xnor U10922 (N_10922,N_8158,N_5037);
or U10923 (N_10923,N_7659,N_8786);
and U10924 (N_10924,N_8872,N_5279);
nand U10925 (N_10925,N_5634,N_7779);
xor U10926 (N_10926,N_8033,N_5414);
or U10927 (N_10927,N_9047,N_6076);
and U10928 (N_10928,N_7116,N_8762);
nor U10929 (N_10929,N_7733,N_9299);
nand U10930 (N_10930,N_9399,N_8821);
and U10931 (N_10931,N_8878,N_5724);
or U10932 (N_10932,N_7516,N_7043);
xnor U10933 (N_10933,N_8790,N_7622);
or U10934 (N_10934,N_6958,N_7907);
xnor U10935 (N_10935,N_6815,N_8735);
nor U10936 (N_10936,N_6028,N_8672);
xnor U10937 (N_10937,N_9018,N_6702);
or U10938 (N_10938,N_5405,N_8509);
xnor U10939 (N_10939,N_6285,N_9247);
or U10940 (N_10940,N_7433,N_7333);
and U10941 (N_10941,N_7756,N_5940);
or U10942 (N_10942,N_9467,N_8651);
and U10943 (N_10943,N_9204,N_5020);
and U10944 (N_10944,N_9538,N_8285);
nand U10945 (N_10945,N_9899,N_9887);
nand U10946 (N_10946,N_7975,N_9588);
nand U10947 (N_10947,N_5291,N_7691);
and U10948 (N_10948,N_6364,N_7976);
or U10949 (N_10949,N_5891,N_7527);
and U10950 (N_10950,N_6802,N_7652);
nand U10951 (N_10951,N_7254,N_7310);
and U10952 (N_10952,N_5100,N_8168);
nor U10953 (N_10953,N_5823,N_9599);
and U10954 (N_10954,N_9994,N_7632);
nand U10955 (N_10955,N_7654,N_9576);
nor U10956 (N_10956,N_8140,N_9274);
or U10957 (N_10957,N_9773,N_7824);
and U10958 (N_10958,N_9014,N_5609);
xnor U10959 (N_10959,N_8987,N_7486);
or U10960 (N_10960,N_9384,N_7318);
nor U10961 (N_10961,N_5761,N_7212);
nand U10962 (N_10962,N_8319,N_6931);
nor U10963 (N_10963,N_5937,N_5500);
nand U10964 (N_10964,N_8753,N_5436);
or U10965 (N_10965,N_6716,N_7161);
and U10966 (N_10966,N_6244,N_6339);
nand U10967 (N_10967,N_9249,N_7331);
xor U10968 (N_10968,N_8688,N_5670);
or U10969 (N_10969,N_5851,N_9633);
and U10970 (N_10970,N_7680,N_9424);
nand U10971 (N_10971,N_9205,N_9077);
and U10972 (N_10972,N_9210,N_5455);
xor U10973 (N_10973,N_7275,N_8573);
and U10974 (N_10974,N_7403,N_9072);
nand U10975 (N_10975,N_7110,N_9498);
and U10976 (N_10976,N_9355,N_8022);
nor U10977 (N_10977,N_7375,N_6960);
or U10978 (N_10978,N_6712,N_8671);
xnor U10979 (N_10979,N_8920,N_8942);
xor U10980 (N_10980,N_6662,N_5681);
or U10981 (N_10981,N_6665,N_9098);
or U10982 (N_10982,N_5864,N_5268);
nor U10983 (N_10983,N_6232,N_5302);
and U10984 (N_10984,N_8325,N_5113);
and U10985 (N_10985,N_6163,N_5598);
nand U10986 (N_10986,N_6855,N_7921);
or U10987 (N_10987,N_9038,N_9109);
or U10988 (N_10988,N_5038,N_8949);
nor U10989 (N_10989,N_9301,N_9127);
or U10990 (N_10990,N_8097,N_9172);
or U10991 (N_10991,N_6074,N_9414);
nand U10992 (N_10992,N_5140,N_9858);
nand U10993 (N_10993,N_7829,N_8005);
nand U10994 (N_10994,N_9514,N_9082);
nor U10995 (N_10995,N_5509,N_6625);
xor U10996 (N_10996,N_8409,N_7055);
nor U10997 (N_10997,N_9315,N_6503);
or U10998 (N_10998,N_8301,N_6477);
xnor U10999 (N_10999,N_6008,N_6657);
nor U11000 (N_11000,N_5217,N_6470);
xor U11001 (N_11001,N_6475,N_6635);
nor U11002 (N_11002,N_9979,N_9405);
or U11003 (N_11003,N_8816,N_5451);
and U11004 (N_11004,N_5098,N_9944);
xnor U11005 (N_11005,N_8435,N_7675);
nor U11006 (N_11006,N_6579,N_9406);
xor U11007 (N_11007,N_6198,N_5862);
nand U11008 (N_11008,N_9306,N_7003);
nand U11009 (N_11009,N_8170,N_5865);
and U11010 (N_11010,N_7615,N_9658);
nor U11011 (N_11011,N_5872,N_5828);
or U11012 (N_11012,N_9398,N_5531);
xnor U11013 (N_11013,N_6814,N_9108);
xnor U11014 (N_11014,N_8237,N_8825);
nor U11015 (N_11015,N_7704,N_7037);
or U11016 (N_11016,N_7297,N_7103);
xor U11017 (N_11017,N_5273,N_8247);
or U11018 (N_11018,N_5647,N_5153);
xor U11019 (N_11019,N_6888,N_9149);
and U11020 (N_11020,N_9910,N_8061);
xnor U11021 (N_11021,N_5719,N_8198);
or U11022 (N_11022,N_5749,N_9373);
or U11023 (N_11023,N_6576,N_7432);
or U11024 (N_11024,N_7707,N_7283);
xor U11025 (N_11025,N_9368,N_8242);
and U11026 (N_11026,N_9727,N_8895);
xor U11027 (N_11027,N_8201,N_7876);
nand U11028 (N_11028,N_9568,N_5584);
or U11029 (N_11029,N_7759,N_6930);
nand U11030 (N_11030,N_5109,N_7647);
or U11031 (N_11031,N_7745,N_8251);
nand U11032 (N_11032,N_5802,N_9078);
xnor U11033 (N_11033,N_9792,N_9095);
and U11034 (N_11034,N_6133,N_5918);
nor U11035 (N_11035,N_5796,N_5176);
nor U11036 (N_11036,N_9623,N_8180);
xnor U11037 (N_11037,N_7125,N_6026);
xor U11038 (N_11038,N_5619,N_5782);
and U11039 (N_11039,N_6777,N_8432);
or U11040 (N_11040,N_9401,N_6723);
nor U11041 (N_11041,N_7145,N_5394);
nor U11042 (N_11042,N_8933,N_8133);
nand U11043 (N_11043,N_6652,N_6222);
and U11044 (N_11044,N_5298,N_9709);
nor U11045 (N_11045,N_9749,N_8362);
xnor U11046 (N_11046,N_7498,N_9300);
nand U11047 (N_11047,N_6898,N_9124);
nand U11048 (N_11048,N_9880,N_5914);
or U11049 (N_11049,N_5303,N_5352);
and U11050 (N_11050,N_9961,N_7443);
nand U11051 (N_11051,N_8797,N_9595);
or U11052 (N_11052,N_6072,N_6320);
nand U11053 (N_11053,N_8072,N_5406);
nor U11054 (N_11054,N_5045,N_8830);
nor U11055 (N_11055,N_7549,N_6087);
or U11056 (N_11056,N_7260,N_9877);
xnor U11057 (N_11057,N_7462,N_8658);
xnor U11058 (N_11058,N_7419,N_9828);
and U11059 (N_11059,N_8293,N_9466);
or U11060 (N_11060,N_8273,N_9245);
nand U11061 (N_11061,N_9536,N_8693);
nand U11062 (N_11062,N_9244,N_7526);
nand U11063 (N_11063,N_5809,N_7825);
nand U11064 (N_11064,N_9687,N_8046);
nor U11065 (N_11065,N_8111,N_5521);
and U11066 (N_11066,N_6268,N_8141);
xnor U11067 (N_11067,N_6909,N_7890);
and U11068 (N_11068,N_7889,N_5442);
or U11069 (N_11069,N_7024,N_6963);
nor U11070 (N_11070,N_8334,N_8105);
nand U11071 (N_11071,N_6132,N_9735);
or U11072 (N_11072,N_8323,N_9457);
or U11073 (N_11073,N_7886,N_9434);
or U11074 (N_11074,N_8986,N_6192);
nand U11075 (N_11075,N_7015,N_6180);
nor U11076 (N_11076,N_5324,N_5759);
or U11077 (N_11077,N_7332,N_9788);
and U11078 (N_11078,N_8860,N_6886);
nand U11079 (N_11079,N_5510,N_6391);
xor U11080 (N_11080,N_8374,N_8765);
nor U11081 (N_11081,N_7645,N_7130);
xor U11082 (N_11082,N_7916,N_7639);
nand U11083 (N_11083,N_7428,N_6969);
nor U11084 (N_11084,N_6618,N_7127);
nor U11085 (N_11085,N_5257,N_9927);
nand U11086 (N_11086,N_5849,N_8423);
and U11087 (N_11087,N_8365,N_8377);
and U11088 (N_11088,N_9578,N_8855);
xor U11089 (N_11089,N_5460,N_8357);
nor U11090 (N_11090,N_5215,N_7773);
and U11091 (N_11091,N_7399,N_5576);
nand U11092 (N_11092,N_5784,N_8376);
nor U11093 (N_11093,N_7468,N_9044);
or U11094 (N_11094,N_5006,N_9075);
nand U11095 (N_11095,N_9620,N_6661);
nor U11096 (N_11096,N_7435,N_5375);
or U11097 (N_11097,N_9589,N_8525);
nor U11098 (N_11098,N_8867,N_6051);
or U11099 (N_11099,N_9618,N_9850);
or U11100 (N_11100,N_7194,N_7996);
xnor U11101 (N_11101,N_9800,N_5597);
nor U11102 (N_11102,N_7227,N_9708);
and U11103 (N_11103,N_7398,N_7461);
nor U11104 (N_11104,N_8882,N_9213);
nand U11105 (N_11105,N_6291,N_5015);
nor U11106 (N_11106,N_7124,N_9114);
xnor U11107 (N_11107,N_5534,N_8327);
xnor U11108 (N_11108,N_7146,N_7520);
or U11109 (N_11109,N_7776,N_7367);
xor U11110 (N_11110,N_7287,N_5831);
nor U11111 (N_11111,N_8429,N_7543);
nor U11112 (N_11112,N_9584,N_8202);
xor U11113 (N_11113,N_9285,N_6447);
nand U11114 (N_11114,N_6227,N_8932);
nand U11115 (N_11115,N_6172,N_9184);
and U11116 (N_11116,N_9237,N_9268);
or U11117 (N_11117,N_8865,N_5214);
xnor U11118 (N_11118,N_9422,N_7602);
nand U11119 (N_11119,N_6089,N_7609);
nand U11120 (N_11120,N_6910,N_6849);
xnor U11121 (N_11121,N_9081,N_7292);
and U11122 (N_11122,N_8495,N_6129);
nor U11123 (N_11123,N_8243,N_6642);
and U11124 (N_11124,N_6740,N_8288);
or U11125 (N_11125,N_9669,N_9479);
or U11126 (N_11126,N_7546,N_5587);
or U11127 (N_11127,N_6088,N_8744);
and U11128 (N_11128,N_9094,N_7783);
xor U11129 (N_11129,N_9878,N_5275);
xor U11130 (N_11130,N_6217,N_8190);
or U11131 (N_11131,N_8270,N_6651);
nor U11132 (N_11132,N_5421,N_5817);
or U11133 (N_11133,N_9162,N_6157);
nor U11134 (N_11134,N_9298,N_6705);
nor U11135 (N_11135,N_8812,N_6214);
nor U11136 (N_11136,N_8519,N_6847);
xor U11137 (N_11137,N_7091,N_7726);
xor U11138 (N_11138,N_6332,N_6399);
or U11139 (N_11139,N_9857,N_8803);
nor U11140 (N_11140,N_6614,N_6363);
nand U11141 (N_11141,N_8206,N_8000);
or U11142 (N_11142,N_6048,N_5175);
nand U11143 (N_11143,N_5989,N_8055);
and U11144 (N_11144,N_6130,N_5444);
or U11145 (N_11145,N_8965,N_5014);
and U11146 (N_11146,N_7760,N_6114);
nand U11147 (N_11147,N_7328,N_6526);
or U11148 (N_11148,N_9360,N_9388);
and U11149 (N_11149,N_5448,N_9917);
nand U11150 (N_11150,N_7900,N_5363);
nor U11151 (N_11151,N_9361,N_5967);
and U11152 (N_11152,N_5834,N_6893);
nand U11153 (N_11153,N_8269,N_8036);
nor U11154 (N_11154,N_6360,N_6346);
nand U11155 (N_11155,N_8017,N_6286);
nor U11156 (N_11156,N_7820,N_8611);
and U11157 (N_11157,N_6302,N_6585);
nand U11158 (N_11158,N_7631,N_7062);
nor U11159 (N_11159,N_5270,N_9836);
or U11160 (N_11160,N_8204,N_8771);
xor U11161 (N_11161,N_7464,N_8726);
and U11162 (N_11162,N_7560,N_9502);
and U11163 (N_11163,N_7685,N_6840);
xnor U11164 (N_11164,N_8619,N_7045);
and U11165 (N_11165,N_8151,N_9966);
or U11166 (N_11166,N_8908,N_7793);
nand U11167 (N_11167,N_9713,N_9754);
nor U11168 (N_11168,N_9560,N_9507);
and U11169 (N_11169,N_5854,N_9380);
and U11170 (N_11170,N_9383,N_6444);
or U11171 (N_11171,N_5079,N_8004);
and U11172 (N_11172,N_6523,N_7195);
nor U11173 (N_11173,N_9591,N_5811);
nor U11174 (N_11174,N_6191,N_5361);
nand U11175 (N_11175,N_8226,N_7349);
nand U11176 (N_11176,N_6204,N_6371);
nand U11177 (N_11177,N_8148,N_7608);
or U11178 (N_11178,N_9810,N_7994);
or U11179 (N_11179,N_6426,N_6678);
xor U11180 (N_11180,N_5354,N_9084);
nand U11181 (N_11181,N_7243,N_5991);
nor U11182 (N_11182,N_9429,N_7603);
xnor U11183 (N_11183,N_6211,N_6643);
or U11184 (N_11184,N_5346,N_6510);
and U11185 (N_11185,N_5919,N_6578);
nand U11186 (N_11186,N_8740,N_9093);
and U11187 (N_11187,N_5128,N_6666);
or U11188 (N_11188,N_8034,N_5440);
nor U11189 (N_11189,N_7072,N_7535);
xor U11190 (N_11190,N_9145,N_7371);
and U11191 (N_11191,N_8330,N_9572);
nand U11192 (N_11192,N_6090,N_9517);
or U11193 (N_11193,N_5949,N_9275);
nor U11194 (N_11194,N_6778,N_9711);
nor U11195 (N_11195,N_8117,N_8130);
nand U11196 (N_11196,N_7789,N_8588);
nor U11197 (N_11197,N_5840,N_5300);
nand U11198 (N_11198,N_7804,N_9020);
and U11199 (N_11199,N_9582,N_5850);
or U11200 (N_11200,N_5157,N_5103);
and U11201 (N_11201,N_8295,N_9656);
or U11202 (N_11202,N_7070,N_6213);
nor U11203 (N_11203,N_8144,N_6022);
and U11204 (N_11204,N_6181,N_7097);
and U11205 (N_11205,N_7854,N_6054);
or U11206 (N_11206,N_6276,N_6145);
or U11207 (N_11207,N_7692,N_7078);
nand U11208 (N_11208,N_6449,N_9915);
nor U11209 (N_11209,N_6175,N_6525);
nand U11210 (N_11210,N_7132,N_8118);
nor U11211 (N_11211,N_9938,N_9197);
and U11212 (N_11212,N_9349,N_8636);
nor U11213 (N_11213,N_5441,N_5870);
nor U11214 (N_11214,N_9327,N_7342);
nand U11215 (N_11215,N_6934,N_9053);
nor U11216 (N_11216,N_9988,N_5718);
and U11217 (N_11217,N_9236,N_8695);
and U11218 (N_11218,N_6957,N_9983);
xor U11219 (N_11219,N_5355,N_8329);
or U11220 (N_11220,N_7456,N_8252);
or U11221 (N_11221,N_9784,N_7694);
and U11222 (N_11222,N_5628,N_9453);
nor U11223 (N_11223,N_6430,N_6591);
xor U11224 (N_11224,N_8853,N_5284);
or U11225 (N_11225,N_7541,N_7500);
or U11226 (N_11226,N_8451,N_7703);
xor U11227 (N_11227,N_9834,N_8694);
or U11228 (N_11228,N_5097,N_6369);
and U11229 (N_11229,N_7792,N_9117);
xor U11230 (N_11230,N_7790,N_8944);
xnor U11231 (N_11231,N_5048,N_5288);
and U11232 (N_11232,N_8548,N_8029);
and U11233 (N_11233,N_9985,N_6839);
or U11234 (N_11234,N_8507,N_7429);
nand U11235 (N_11235,N_6040,N_9211);
xor U11236 (N_11236,N_5881,N_5245);
or U11237 (N_11237,N_7618,N_8703);
and U11238 (N_11238,N_5246,N_5925);
nand U11239 (N_11239,N_6328,N_7392);
nand U11240 (N_11240,N_5204,N_9022);
nand U11241 (N_11241,N_7120,N_8880);
nor U11242 (N_11242,N_5484,N_7774);
xnor U11243 (N_11243,N_6825,N_7833);
nand U11244 (N_11244,N_6993,N_8297);
and U11245 (N_11245,N_5260,N_8065);
nand U11246 (N_11246,N_6832,N_9688);
nand U11247 (N_11247,N_6710,N_9310);
and U11248 (N_11248,N_7982,N_5391);
nand U11249 (N_11249,N_5085,N_9513);
nand U11250 (N_11250,N_7569,N_6660);
nand U11251 (N_11251,N_5308,N_5518);
nor U11252 (N_11252,N_5770,N_6605);
and U11253 (N_11253,N_9548,N_5567);
and U11254 (N_11254,N_6746,N_9543);
and U11255 (N_11255,N_9478,N_5528);
xnor U11256 (N_11256,N_9787,N_9791);
and U11257 (N_11257,N_9775,N_7334);
nor U11258 (N_11258,N_9949,N_8847);
nand U11259 (N_11259,N_9407,N_9815);
and U11260 (N_11260,N_8841,N_8840);
xnor U11261 (N_11261,N_6603,N_6880);
nand U11262 (N_11262,N_6770,N_7533);
nand U11263 (N_11263,N_8988,N_8452);
xnor U11264 (N_11264,N_6882,N_6183);
or U11265 (N_11265,N_7233,N_7540);
and U11266 (N_11266,N_7809,N_6335);
and U11267 (N_11267,N_7073,N_7459);
or U11268 (N_11268,N_9704,N_7839);
or U11269 (N_11269,N_6009,N_9748);
and U11270 (N_11270,N_6903,N_7442);
xnor U11271 (N_11271,N_9954,N_7075);
and U11272 (N_11272,N_7885,N_6708);
and U11273 (N_11273,N_5181,N_5224);
nor U11274 (N_11274,N_7039,N_7702);
xnor U11275 (N_11275,N_5758,N_7939);
nor U11276 (N_11276,N_8074,N_5480);
nand U11277 (N_11277,N_6193,N_5088);
nor U11278 (N_11278,N_5323,N_6106);
nor U11279 (N_11279,N_6207,N_7957);
xnor U11280 (N_11280,N_6231,N_5529);
xnor U11281 (N_11281,N_5756,N_9080);
and U11282 (N_11282,N_9420,N_9724);
and U11283 (N_11283,N_7534,N_8687);
and U11284 (N_11284,N_5453,N_6101);
xor U11285 (N_11285,N_5266,N_6248);
or U11286 (N_11286,N_8052,N_6600);
nor U11287 (N_11287,N_7617,N_9190);
and U11288 (N_11288,N_6000,N_9139);
and U11289 (N_11289,N_7424,N_9309);
or U11290 (N_11290,N_7784,N_5120);
or U11291 (N_11291,N_7241,N_9463);
xor U11292 (N_11292,N_7689,N_7512);
and U11293 (N_11293,N_9914,N_5124);
xor U11294 (N_11294,N_7158,N_8417);
or U11295 (N_11295,N_5081,N_8545);
nor U11296 (N_11296,N_7232,N_5255);
or U11297 (N_11297,N_7059,N_6805);
or U11298 (N_11298,N_5149,N_6761);
or U11299 (N_11299,N_9703,N_6002);
nand U11300 (N_11300,N_9630,N_6454);
nor U11301 (N_11301,N_9461,N_9847);
nand U11302 (N_11302,N_7623,N_9520);
or U11303 (N_11303,N_8846,N_5810);
nor U11304 (N_11304,N_8030,N_8195);
nor U11305 (N_11305,N_8601,N_8091);
nor U11306 (N_11306,N_5208,N_6992);
or U11307 (N_11307,N_9567,N_5307);
and U11308 (N_11308,N_9366,N_6912);
nor U11309 (N_11309,N_8829,N_9718);
or U11310 (N_11310,N_8885,N_7972);
and U11311 (N_11311,N_9385,N_7138);
nand U11312 (N_11312,N_9347,N_9639);
nand U11313 (N_11313,N_7286,N_8937);
nand U11314 (N_11314,N_8485,N_6562);
xor U11315 (N_11315,N_5368,N_6030);
or U11316 (N_11316,N_5491,N_5285);
nor U11317 (N_11317,N_5858,N_9006);
nand U11318 (N_11318,N_8643,N_5690);
and U11319 (N_11319,N_5395,N_7586);
or U11320 (N_11320,N_7630,N_6472);
nand U11321 (N_11321,N_9345,N_8453);
nand U11322 (N_11322,N_5739,N_9743);
xnor U11323 (N_11323,N_9575,N_8178);
nor U11324 (N_11324,N_5495,N_7769);
and U11325 (N_11325,N_7406,N_7754);
or U11326 (N_11326,N_5578,N_8512);
or U11327 (N_11327,N_7258,N_9339);
nand U11328 (N_11328,N_5409,N_9796);
nor U11329 (N_11329,N_8318,N_7381);
xnor U11330 (N_11330,N_7222,N_6541);
and U11331 (N_11331,N_8581,N_6152);
xor U11332 (N_11332,N_9175,N_8723);
nor U11333 (N_11333,N_9367,N_5539);
xor U11334 (N_11334,N_5764,N_5373);
nor U11335 (N_11335,N_6012,N_6015);
and U11336 (N_11336,N_8716,N_8084);
nor U11337 (N_11337,N_7751,N_8561);
xnor U11338 (N_11338,N_7721,N_5664);
nand U11339 (N_11339,N_6247,N_9528);
and U11340 (N_11340,N_7160,N_7496);
xor U11341 (N_11341,N_7843,N_8272);
and U11342 (N_11342,N_9105,N_7954);
xor U11343 (N_11343,N_6501,N_7511);
xnor U11344 (N_11344,N_7068,N_8559);
or U11345 (N_11345,N_9835,N_5137);
nand U11346 (N_11346,N_8037,N_8501);
nand U11347 (N_11347,N_9631,N_5198);
xor U11348 (N_11348,N_6808,N_7279);
nor U11349 (N_11349,N_9028,N_6465);
nand U11350 (N_11350,N_6083,N_9947);
or U11351 (N_11351,N_6659,N_7211);
xnor U11352 (N_11352,N_6905,N_7619);
and U11353 (N_11353,N_8079,N_6881);
and U11354 (N_11354,N_8844,N_8056);
nor U11355 (N_11355,N_9912,N_8842);
xor U11356 (N_11356,N_6857,N_7646);
xor U11357 (N_11357,N_8664,N_6978);
or U11358 (N_11358,N_9066,N_6664);
xor U11359 (N_11359,N_8063,N_8183);
nor U11360 (N_11360,N_5013,N_9277);
nor U11361 (N_11361,N_6742,N_9248);
or U11362 (N_11362,N_5793,N_8231);
xnor U11363 (N_11363,N_6309,N_7505);
nand U11364 (N_11364,N_7063,N_7029);
and U11365 (N_11365,N_7948,N_8324);
or U11366 (N_11366,N_6081,N_5244);
nor U11367 (N_11367,N_8565,N_8442);
or U11368 (N_11368,N_5093,N_5511);
xnor U11369 (N_11369,N_7152,N_6038);
nor U11370 (N_11370,N_8632,N_9419);
or U11371 (N_11371,N_7897,N_6160);
or U11372 (N_11372,N_6563,N_6860);
nand U11373 (N_11373,N_5615,N_9883);
xnor U11374 (N_11374,N_5209,N_7531);
xor U11375 (N_11375,N_7842,N_8951);
nor U11376 (N_11376,N_6137,N_5471);
xnor U11377 (N_11377,N_7558,N_8203);
xnor U11378 (N_11378,N_6250,N_8426);
xor U11379 (N_11379,N_8184,N_6460);
nand U11380 (N_11380,N_7736,N_8991);
xor U11381 (N_11381,N_5066,N_5695);
and U11382 (N_11382,N_7408,N_6086);
or U11383 (N_11383,N_8752,N_8260);
and U11384 (N_11384,N_8254,N_6582);
and U11385 (N_11385,N_9627,N_6680);
nor U11386 (N_11386,N_5547,N_5389);
xor U11387 (N_11387,N_7522,N_9533);
xor U11388 (N_11388,N_7781,N_6124);
xnor U11389 (N_11389,N_5873,N_8571);
and U11390 (N_11390,N_8883,N_8031);
and U11391 (N_11391,N_5995,N_5252);
xnor U11392 (N_11392,N_5133,N_5387);
or U11393 (N_11393,N_6428,N_5768);
nor U11394 (N_11394,N_6599,N_7950);
or U11395 (N_11395,N_8468,N_6551);
and U11396 (N_11396,N_8957,N_5380);
xnor U11397 (N_11397,N_6862,N_5508);
or U11398 (N_11398,N_9875,N_6607);
nor U11399 (N_11399,N_5274,N_5404);
or U11400 (N_11400,N_9903,N_9288);
nand U11401 (N_11401,N_9995,N_6697);
nand U11402 (N_11402,N_9963,N_7144);
nor U11403 (N_11403,N_9577,N_6471);
xor U11404 (N_11404,N_6307,N_6150);
xor U11405 (N_11405,N_7722,N_7922);
nand U11406 (N_11406,N_5378,N_6524);
xor U11407 (N_11407,N_5040,N_8443);
xor U11408 (N_11408,N_7105,N_8286);
nor U11409 (N_11409,N_8418,N_9138);
or U11410 (N_11410,N_5130,N_6321);
nor U11411 (N_11411,N_7330,N_9926);
nor U11412 (N_11412,N_8322,N_6720);
nand U11413 (N_11413,N_9652,N_8135);
nand U11414 (N_11414,N_7472,N_5801);
nand U11415 (N_11415,N_6474,N_8048);
and U11416 (N_11416,N_9635,N_8590);
xnor U11417 (N_11417,N_7355,N_8959);
and U11418 (N_11418,N_5976,N_9892);
and U11419 (N_11419,N_6817,N_9340);
and U11420 (N_11420,N_8510,N_7041);
or U11421 (N_11421,N_8808,N_8556);
nor U11422 (N_11422,N_6096,N_9755);
or U11423 (N_11423,N_7234,N_7182);
xnor U11424 (N_11424,N_8210,N_7187);
nor U11425 (N_11425,N_7696,N_8788);
nand U11426 (N_11426,N_9283,N_5178);
or U11427 (N_11427,N_8340,N_6748);
nor U11428 (N_11428,N_5622,N_7517);
nand U11429 (N_11429,N_8950,N_9898);
nor U11430 (N_11430,N_9272,N_5435);
xnor U11431 (N_11431,N_8864,N_8524);
and U11432 (N_11432,N_8076,N_8258);
nand U11433 (N_11433,N_9556,N_8659);
nor U11434 (N_11434,N_7668,N_8859);
and U11435 (N_11435,N_5164,N_7494);
and U11436 (N_11436,N_9860,N_6677);
and U11437 (N_11437,N_6943,N_9593);
nor U11438 (N_11438,N_6223,N_9515);
and U11439 (N_11439,N_6711,N_6679);
xnor U11440 (N_11440,N_8655,N_5243);
or U11441 (N_11441,N_8436,N_5866);
xnor U11442 (N_11442,N_8399,N_7911);
nand U11443 (N_11443,N_5086,N_7084);
nand U11444 (N_11444,N_8914,N_7797);
or U11445 (N_11445,N_8836,N_9870);
and U11446 (N_11446,N_7942,N_5099);
and U11447 (N_11447,N_6166,N_6750);
and U11448 (N_11448,N_7306,N_9632);
nor U11449 (N_11449,N_5715,N_5125);
or U11450 (N_11450,N_9934,N_5685);
nor U11451 (N_11451,N_5360,N_7143);
and U11452 (N_11452,N_9527,N_6557);
or U11453 (N_11453,N_7868,N_9048);
xnor U11454 (N_11454,N_7559,N_6584);
nand U11455 (N_11455,N_7891,N_9971);
and U11456 (N_11456,N_8431,N_5101);
nor U11457 (N_11457,N_9919,N_5220);
and U11458 (N_11458,N_6831,N_5610);
or U11459 (N_11459,N_6281,N_5985);
and U11460 (N_11460,N_8504,N_5614);
and U11461 (N_11461,N_9097,N_7199);
nand U11462 (N_11462,N_7131,N_6951);
and U11463 (N_11463,N_9041,N_5476);
and U11464 (N_11464,N_6271,N_5472);
xor U11465 (N_11465,N_9025,N_6672);
nand U11466 (N_11466,N_9665,N_6324);
nor U11467 (N_11467,N_5493,N_9009);
nor U11468 (N_11468,N_5278,N_5202);
and U11469 (N_11469,N_8838,N_9830);
nor U11470 (N_11470,N_6203,N_5068);
nand U11471 (N_11471,N_5595,N_8433);
and U11472 (N_11472,N_9465,N_6230);
and U11473 (N_11473,N_7035,N_5880);
or U11474 (N_11474,N_6123,N_5090);
nor U11475 (N_11475,N_8725,N_6092);
or U11476 (N_11476,N_9907,N_7649);
or U11477 (N_11477,N_8457,N_8464);
nand U11478 (N_11478,N_6058,N_7162);
or U11479 (N_11479,N_9541,N_8042);
xnor U11480 (N_11480,N_8358,N_7818);
or U11481 (N_11481,N_8480,N_8088);
and U11482 (N_11482,N_7932,N_6065);
nor U11483 (N_11483,N_5963,N_8769);
and U11484 (N_11484,N_6560,N_8103);
and U11485 (N_11485,N_6055,N_7713);
nor U11486 (N_11486,N_5867,N_9931);
and U11487 (N_11487,N_7830,N_7001);
and U11488 (N_11488,N_5112,N_7752);
and U11489 (N_11489,N_8689,N_6616);
and U11490 (N_11490,N_8116,N_8793);
or U11491 (N_11491,N_7782,N_8412);
nand U11492 (N_11492,N_5680,N_5116);
xor U11493 (N_11493,N_5621,N_6438);
and U11494 (N_11494,N_7081,N_7346);
xnor U11495 (N_11495,N_5565,N_8670);
nor U11496 (N_11496,N_5727,N_5481);
nand U11497 (N_11497,N_9223,N_8353);
or U11498 (N_11498,N_5841,N_6813);
and U11499 (N_11499,N_6729,N_8057);
xor U11500 (N_11500,N_7850,N_9693);
xnor U11501 (N_11501,N_5104,N_9807);
or U11502 (N_11502,N_7987,N_8849);
or U11503 (N_11503,N_8120,N_8309);
and U11504 (N_11504,N_9106,N_6294);
and U11505 (N_11505,N_8490,N_8175);
nor U11506 (N_11506,N_8370,N_8886);
and U11507 (N_11507,N_9655,N_5822);
or U11508 (N_11508,N_9653,N_6873);
nor U11509 (N_11509,N_7576,N_8043);
nand U11510 (N_11510,N_7597,N_6558);
or U11511 (N_11511,N_9284,N_5022);
and U11512 (N_11512,N_6381,N_7203);
nor U11513 (N_11513,N_5637,N_8552);
nor U11514 (N_11514,N_5349,N_8647);
and U11515 (N_11515,N_5376,N_5197);
or U11516 (N_11516,N_9716,N_5777);
nor U11517 (N_11517,N_6879,N_8397);
xor U11518 (N_11518,N_7938,N_8528);
xor U11519 (N_11519,N_5200,N_6280);
xnor U11520 (N_11520,N_6067,N_9768);
xnor U11521 (N_11521,N_7529,N_5226);
nor U11522 (N_11522,N_9292,N_7814);
xnor U11523 (N_11523,N_7093,N_7737);
xnor U11524 (N_11524,N_6639,N_7530);
and U11525 (N_11525,N_5107,N_5658);
or U11526 (N_11526,N_5874,N_5697);
and U11527 (N_11527,N_8690,N_9425);
and U11528 (N_11528,N_6694,N_6974);
nor U11529 (N_11529,N_6901,N_6724);
xnor U11530 (N_11530,N_6592,N_5627);
or U11531 (N_11531,N_5694,N_5301);
nand U11532 (N_11532,N_7725,N_8766);
nand U11533 (N_11533,N_5310,N_6405);
nor U11534 (N_11534,N_8798,N_7319);
or U11535 (N_11535,N_5608,N_7791);
or U11536 (N_11536,N_5545,N_6201);
and U11537 (N_11537,N_9766,N_5077);
or U11538 (N_11538,N_9250,N_9684);
xnor U11539 (N_11539,N_8639,N_9741);
xor U11540 (N_11540,N_7469,N_8496);
nand U11541 (N_11541,N_9088,N_8077);
and U11542 (N_11542,N_8751,N_7847);
xor U11543 (N_11543,N_9699,N_7405);
nor U11544 (N_11544,N_6383,N_8087);
nand U11545 (N_11545,N_8321,N_9417);
or U11546 (N_11546,N_6059,N_5043);
nand U11547 (N_11547,N_5117,N_9232);
nand U11548 (N_11548,N_9491,N_5135);
xor U11549 (N_11549,N_6509,N_7607);
and U11550 (N_11550,N_8854,N_9816);
and U11551 (N_11551,N_7811,N_9799);
nor U11552 (N_11552,N_5830,N_8013);
or U11553 (N_11553,N_7004,N_9024);
or U11554 (N_11554,N_7997,N_9622);
xnor U11555 (N_11555,N_7046,N_6878);
nor U11556 (N_11556,N_5541,N_8736);
nor U11557 (N_11557,N_9579,N_6102);
and U11558 (N_11558,N_7163,N_9208);
xnor U11559 (N_11559,N_5795,N_8994);
nand U11560 (N_11560,N_5060,N_9431);
and U11561 (N_11561,N_5426,N_6776);
nand U11562 (N_11562,N_6287,N_6317);
nand U11563 (N_11563,N_5030,N_8425);
or U11564 (N_11564,N_7264,N_6491);
nor U11565 (N_11565,N_7338,N_9731);
nor U11566 (N_11566,N_6390,N_8475);
and U11567 (N_11567,N_9259,N_9039);
nor U11568 (N_11568,N_5913,N_6985);
and U11569 (N_11569,N_6682,N_6892);
or U11570 (N_11570,N_9545,N_8328);
xor U11571 (N_11571,N_7025,N_5898);
nand U11572 (N_11572,N_7304,N_8024);
nor U11573 (N_11573,N_9433,N_7474);
nand U11574 (N_11574,N_6548,N_9397);
nor U11575 (N_11575,N_9794,N_6366);
xnor U11576 (N_11576,N_6334,N_7156);
or U11577 (N_11577,N_6462,N_6566);
xnor U11578 (N_11578,N_5416,N_9415);
xnor U11579 (N_11579,N_5201,N_8606);
nand U11580 (N_11580,N_9518,N_8926);
nor U11581 (N_11581,N_9180,N_5709);
xor U11582 (N_11582,N_8794,N_9040);
xor U11583 (N_11583,N_7094,N_5755);
and U11584 (N_11584,N_7815,N_5980);
or U11585 (N_11585,N_5400,N_5139);
or U11586 (N_11586,N_5767,N_8823);
nor U11587 (N_11587,N_8589,N_9606);
or U11588 (N_11588,N_7590,N_8576);
or U11589 (N_11589,N_8884,N_6796);
xor U11590 (N_11590,N_8789,N_5313);
xor U11591 (N_11591,N_8477,N_8903);
and U11592 (N_11592,N_6700,N_8952);
nand U11593 (N_11593,N_5640,N_9839);
nand U11594 (N_11594,N_6212,N_8554);
nand U11595 (N_11595,N_9222,N_5707);
and U11596 (N_11596,N_7272,N_9747);
and U11597 (N_11597,N_8428,N_5571);
nor U11598 (N_11598,N_7175,N_7053);
nand U11599 (N_11599,N_5616,N_9750);
nand U11600 (N_11600,N_6675,N_9350);
nand U11601 (N_11601,N_8444,N_9706);
nand U11602 (N_11602,N_9054,N_6995);
nand U11603 (N_11603,N_6640,N_7128);
nor U11604 (N_11604,N_7796,N_8520);
or U11605 (N_11605,N_9881,N_5523);
or U11606 (N_11606,N_8985,N_8775);
or U11607 (N_11607,N_6899,N_7434);
nor U11608 (N_11608,N_7537,N_6041);
and U11609 (N_11609,N_5855,N_9229);
xor U11610 (N_11610,N_6630,N_6623);
or U11611 (N_11611,N_7785,N_5059);
nand U11612 (N_11612,N_6921,N_5654);
xor U11613 (N_11613,N_8129,N_5871);
nor U11614 (N_11614,N_9086,N_8185);
or U11615 (N_11615,N_8302,N_7918);
xnor U11616 (N_11616,N_9767,N_5073);
or U11617 (N_11617,N_5662,N_5632);
and U11618 (N_11618,N_5592,N_9734);
nor U11619 (N_11619,N_9821,N_9276);
or U11620 (N_11620,N_9737,N_5987);
nand U11621 (N_11621,N_8873,N_9644);
or U11622 (N_11622,N_9192,N_5875);
nand U11623 (N_11623,N_8054,N_9642);
xor U11624 (N_11624,N_6763,N_6464);
and U11625 (N_11625,N_6645,N_8294);
nor U11626 (N_11626,N_8503,N_8002);
nand U11627 (N_11627,N_7395,N_7401);
xor U11628 (N_11628,N_9393,N_9230);
nor U11629 (N_11629,N_9817,N_7183);
or U11630 (N_11630,N_7148,N_6823);
xnor U11631 (N_11631,N_6549,N_7981);
nor U11632 (N_11632,N_6259,N_5132);
xnor U11633 (N_11633,N_9021,N_8916);
nor U11634 (N_11634,N_9241,N_7990);
or U11635 (N_11635,N_5775,N_9427);
and U11636 (N_11636,N_6812,N_5882);
nand U11637 (N_11637,N_7164,N_5071);
nand U11638 (N_11638,N_6834,N_8474);
xor U11639 (N_11639,N_7986,N_9943);
and U11640 (N_11640,N_7660,N_8954);
and U11641 (N_11641,N_5253,N_5650);
xnor U11642 (N_11642,N_6867,N_6937);
xor U11643 (N_11643,N_8470,N_8174);
and U11644 (N_11644,N_5746,N_8930);
or U11645 (N_11645,N_5779,N_6908);
nor U11646 (N_11646,N_9786,N_5752);
nand U11647 (N_11647,N_7798,N_8839);
xor U11648 (N_11648,N_7280,N_7228);
xnor U11649 (N_11649,N_5826,N_9935);
nor U11650 (N_11650,N_6420,N_8481);
xnor U11651 (N_11651,N_6790,N_5145);
or U11652 (N_11652,N_6574,N_9826);
or U11653 (N_11653,N_8488,N_7476);
nand U11654 (N_11654,N_8995,N_7047);
or U11655 (N_11655,N_8508,N_6273);
or U11656 (N_11656,N_6111,N_9873);
nand U11657 (N_11657,N_7255,N_7251);
nor U11658 (N_11658,N_9458,N_8235);
nor U11659 (N_11659,N_5643,N_5076);
xnor U11660 (N_11660,N_7363,N_8411);
xor U11661 (N_11661,N_6851,N_9334);
xor U11662 (N_11662,N_8562,N_5878);
and U11663 (N_11663,N_9854,N_7261);
nor U11664 (N_11664,N_5193,N_7763);
and U11665 (N_11665,N_5589,N_7772);
nor U11666 (N_11666,N_5459,N_5753);
or U11667 (N_11667,N_8638,N_8598);
and U11668 (N_11668,N_6290,N_6344);
and U11669 (N_11669,N_8558,N_8580);
xnor U11670 (N_11670,N_6010,N_8173);
and U11671 (N_11671,N_6668,N_6631);
and U11672 (N_11672,N_9207,N_8595);
nand U11673 (N_11673,N_7028,N_9663);
nor U11674 (N_11674,N_6176,N_9818);
xnor U11675 (N_11675,N_8996,N_9168);
and U11676 (N_11676,N_7281,N_8876);
and U11677 (N_11677,N_8375,N_6843);
nand U11678 (N_11678,N_5901,N_8645);
nor U11679 (N_11679,N_7141,N_7657);
xor U11680 (N_11680,N_6550,N_7816);
and U11681 (N_11681,N_8913,N_6001);
xor U11682 (N_11682,N_5563,N_9692);
or U11683 (N_11683,N_7074,N_6005);
and U11684 (N_11684,N_7627,N_6398);
nand U11685 (N_11685,N_9720,N_8912);
or U11686 (N_11686,N_7940,N_9759);
or U11687 (N_11687,N_7202,N_6295);
and U11688 (N_11688,N_8715,N_7730);
nand U11689 (N_11689,N_6596,N_8862);
and U11690 (N_11690,N_5735,N_9260);
and U11691 (N_11691,N_7961,N_8756);
nor U11692 (N_11692,N_8100,N_6165);
nor U11693 (N_11693,N_7247,N_6522);
nor U11694 (N_11694,N_6786,N_9551);
and U11695 (N_11695,N_8940,N_6686);
nor U11696 (N_11696,N_6345,N_8040);
xnor U11697 (N_11697,N_5922,N_9412);
nor U11698 (N_11698,N_7515,N_8236);
nor U11699 (N_11699,N_5562,N_8795);
and U11700 (N_11700,N_5934,N_8122);
nand U11701 (N_11701,N_5787,N_9666);
xnor U11702 (N_11702,N_9888,N_8826);
nand U11703 (N_11703,N_7584,N_5931);
nand U11704 (N_11704,N_6894,N_7273);
nand U11705 (N_11705,N_9690,N_8679);
and U11706 (N_11706,N_7844,N_9354);
xnor U11707 (N_11707,N_5560,N_5384);
or U11708 (N_11708,N_7305,N_9780);
and U11709 (N_11709,N_5859,N_8879);
and U11710 (N_11710,N_5353,N_9101);
and U11711 (N_11711,N_7552,N_6079);
nand U11712 (N_11712,N_6990,N_6942);
or U11713 (N_11713,N_5723,N_8819);
nand U11714 (N_11714,N_8051,N_6246);
or U11715 (N_11715,N_9252,N_8699);
nor U11716 (N_11716,N_7967,N_7246);
and U11717 (N_11717,N_8265,N_7357);
and U11718 (N_11718,N_5698,N_7301);
nor U11719 (N_11719,N_6118,N_5002);
xnor U11720 (N_11720,N_8263,N_9147);
nor U11721 (N_11721,N_5682,N_7565);
nand U11722 (N_11722,N_5552,N_5160);
nor U11723 (N_11723,N_6644,N_6056);
nand U11724 (N_11724,N_6538,N_7803);
nand U11725 (N_11725,N_5251,N_8400);
nand U11726 (N_11726,N_7402,N_8045);
nor U11727 (N_11727,N_5751,N_7497);
xnor U11728 (N_11728,N_6870,N_5151);
and U11729 (N_11729,N_7595,N_8473);
and U11730 (N_11730,N_5769,N_8511);
and U11731 (N_11731,N_5663,N_7092);
and U11732 (N_11732,N_5704,N_9936);
and U11733 (N_11733,N_7878,N_7427);
nand U11734 (N_11734,N_8901,N_9561);
or U11735 (N_11735,N_7563,N_8707);
and U11736 (N_11736,N_9365,N_9625);
nand U11737 (N_11737,N_7079,N_6884);
or U11738 (N_11738,N_9137,N_8472);
nand U11739 (N_11739,N_8459,N_6569);
and U11740 (N_11740,N_6060,N_9269);
or U11741 (N_11741,N_5564,N_5228);
nand U11742 (N_11742,N_8704,N_8712);
xor U11743 (N_11743,N_5712,N_6370);
xnor U11744 (N_11744,N_5754,N_8542);
or U11745 (N_11745,N_6610,N_9566);
xnor U11746 (N_11746,N_7780,N_5454);
nor U11747 (N_11747,N_7555,N_7348);
nor U11748 (N_11748,N_6848,N_8983);
nor U11749 (N_11749,N_8553,N_7149);
xnor U11750 (N_11750,N_8284,N_8570);
xor U11751 (N_11751,N_5169,N_7134);
nor U11752 (N_11752,N_5847,N_8080);
and U11753 (N_11753,N_5743,N_5885);
xor U11754 (N_11754,N_6669,N_6531);
nand U11755 (N_11755,N_8454,N_7495);
and U11756 (N_11756,N_6251,N_8271);
and U11757 (N_11757,N_5469,N_6530);
nor U11758 (N_11758,N_8083,N_6189);
nand U11759 (N_11759,N_7307,N_5182);
or U11760 (N_11760,N_5936,N_7606);
xnor U11761 (N_11761,N_7741,N_7438);
nand U11762 (N_11762,N_8555,N_6485);
and U11763 (N_11763,N_9151,N_8032);
nand U11764 (N_11764,N_6824,N_9019);
xnor U11765 (N_11765,N_8541,N_6788);
nand U11766 (N_11766,N_7080,N_6441);
and U11767 (N_11767,N_5543,N_5921);
and U11768 (N_11768,N_7189,N_6891);
or U11769 (N_11769,N_8605,N_5347);
and U11770 (N_11770,N_5920,N_7083);
nand U11771 (N_11771,N_5645,N_8261);
or U11772 (N_11772,N_9660,N_9439);
nor U11773 (N_11773,N_7848,N_5824);
and U11774 (N_11774,N_8067,N_9279);
nand U11775 (N_11775,N_8539,N_7071);
nand U11776 (N_11776,N_8137,N_6461);
nor U11777 (N_11777,N_9007,N_9789);
nor U11778 (N_11778,N_9636,N_7220);
nand U11779 (N_11779,N_6656,N_7036);
xnor U11780 (N_11780,N_8386,N_9901);
xnor U11781 (N_11781,N_6045,N_9965);
nand U11782 (N_11782,N_9455,N_5443);
and U11783 (N_11783,N_5929,N_7267);
nand U11784 (N_11784,N_7374,N_5642);
and U11785 (N_11785,N_6810,N_7104);
xnor U11786 (N_11786,N_8602,N_7573);
nand U11787 (N_11787,N_6692,N_6782);
and U11788 (N_11788,N_6833,N_5412);
and U11789 (N_11789,N_7060,N_8523);
or U11790 (N_11790,N_8219,N_6224);
nand U11791 (N_11791,N_5617,N_9975);
xor U11792 (N_11792,N_6706,N_6601);
and U11793 (N_11793,N_6392,N_9318);
nor U11794 (N_11794,N_8396,N_8150);
nor U11795 (N_11795,N_8463,N_9382);
or U11796 (N_11796,N_5467,N_9605);
nand U11797 (N_11797,N_6753,N_7802);
or U11798 (N_11798,N_5717,N_7038);
xnor U11799 (N_11799,N_9326,N_5548);
xor U11800 (N_11800,N_7139,N_6604);
and U11801 (N_11801,N_9908,N_9099);
nor U11802 (N_11802,N_6632,N_7909);
nor U11803 (N_11803,N_5533,N_6057);
or U11804 (N_11804,N_7285,N_8997);
xor U11805 (N_11805,N_8698,N_7321);
nand U11806 (N_11806,N_6598,N_5315);
and U11807 (N_11807,N_7140,N_6278);
nor U11808 (N_11808,N_7706,N_9723);
and U11809 (N_11809,N_8282,N_9240);
nand U11810 (N_11810,N_6463,N_6911);
nor U11811 (N_11811,N_7184,N_8349);
or U11812 (N_11812,N_8214,N_5674);
nor U11813 (N_11813,N_9135,N_6306);
or U11814 (N_11814,N_7777,N_6561);
nor U11815 (N_11815,N_6984,N_5141);
xnor U11816 (N_11816,N_5669,N_8663);
nand U11817 (N_11817,N_7556,N_9676);
or U11818 (N_11818,N_7574,N_8684);
or U11819 (N_11819,N_7221,N_8616);
xnor U11820 (N_11820,N_9504,N_6141);
nand U11821 (N_11821,N_6233,N_9444);
or U11822 (N_11822,N_9900,N_7492);
nor U11823 (N_11823,N_8540,N_9271);
xor U11824 (N_11824,N_9261,N_7724);
nor U11825 (N_11825,N_8720,N_5388);
and U11826 (N_11826,N_9890,N_7587);
and U11827 (N_11827,N_6953,N_6380);
and U11828 (N_11828,N_7965,N_9410);
and U11829 (N_11829,N_9700,N_9744);
nor U11830 (N_11830,N_5162,N_6236);
and U11831 (N_11831,N_6747,N_5410);
nor U11832 (N_11832,N_7117,N_5905);
nand U11833 (N_11833,N_8629,N_9924);
xor U11834 (N_11834,N_6571,N_6097);
nand U11835 (N_11835,N_7553,N_8147);
nand U11836 (N_11836,N_9155,N_7991);
and U11837 (N_11837,N_9895,N_6153);
or U11838 (N_11838,N_6741,N_6968);
or U11839 (N_11839,N_5258,N_8608);
xnor U11840 (N_11840,N_6459,N_6488);
xor U11841 (N_11841,N_7361,N_8543);
xnor U11842 (N_11842,N_6257,N_9612);
nor U11843 (N_11843,N_5374,N_7600);
or U11844 (N_11844,N_6973,N_9762);
xor U11845 (N_11845,N_9945,N_6826);
xor U11846 (N_11846,N_9524,N_5072);
nor U11847 (N_11847,N_7482,N_5398);
or U11848 (N_11848,N_6732,N_8705);
or U11849 (N_11849,N_9897,N_7467);
and U11850 (N_11850,N_5019,N_5196);
or U11851 (N_11851,N_6336,N_7944);
and U11852 (N_11852,N_8461,N_7453);
or U11853 (N_11853,N_9146,N_6916);
and U11854 (N_11854,N_7904,N_8618);
nor U11855 (N_11855,N_8711,N_5486);
and U11856 (N_11856,N_6013,N_8806);
or U11857 (N_11857,N_5686,N_9893);
and U11858 (N_11858,N_7100,N_7042);
and U11859 (N_11859,N_7735,N_9619);
xor U11860 (N_11860,N_6156,N_7538);
xor U11861 (N_11861,N_7391,N_6500);
and U11862 (N_11862,N_9227,N_6253);
or U11863 (N_11863,N_7151,N_6806);
nor U11864 (N_11864,N_6820,N_6731);
nor U11865 (N_11865,N_5774,N_7542);
and U11866 (N_11866,N_5556,N_7656);
nand U11867 (N_11867,N_5158,N_9492);
nand U11868 (N_11868,N_7596,N_9003);
xor U11869 (N_11869,N_5844,N_7360);
nor U11870 (N_11870,N_6811,N_9199);
and U11871 (N_11871,N_5332,N_8167);
nand U11872 (N_11872,N_7805,N_9060);
xnor U11873 (N_11873,N_9657,N_7681);
or U11874 (N_11874,N_5700,N_8654);
and U11875 (N_11875,N_6736,N_5377);
nand U11876 (N_11876,N_8828,N_5890);
and U11877 (N_11877,N_6999,N_8582);
nand U11878 (N_11878,N_8035,N_5593);
or U11879 (N_11879,N_6588,N_7480);
xnor U11880 (N_11880,N_5569,N_7993);
xnor U11881 (N_11881,N_5524,N_7064);
nor U11882 (N_11882,N_7598,N_9760);
nand U11883 (N_11883,N_8778,N_6904);
nor U11884 (N_11884,N_9484,N_9324);
nor U11885 (N_11885,N_6171,N_7936);
nor U11886 (N_11886,N_6185,N_5420);
xor U11887 (N_11887,N_9984,N_9648);
and U11888 (N_11888,N_7926,N_5057);
nor U11889 (N_11889,N_7935,N_8621);
xor U11890 (N_11890,N_6116,N_8518);
and U11891 (N_11891,N_8416,N_5119);
nand U11892 (N_11892,N_9305,N_9233);
and U11893 (N_11893,N_6293,N_8025);
or U11894 (N_11894,N_9929,N_5786);
xnor U11895 (N_11895,N_7159,N_7838);
nand U11896 (N_11896,N_8833,N_9694);
and U11897 (N_11897,N_5144,N_7219);
nand U11898 (N_11898,N_6349,N_9913);
nor U11899 (N_11899,N_8644,N_7910);
xnor U11900 (N_11900,N_5429,N_6241);
or U11901 (N_11901,N_6448,N_8742);
or U11902 (N_11902,N_7448,N_5618);
and U11903 (N_11903,N_5799,N_8924);
xor U11904 (N_11904,N_6721,N_9110);
and U11905 (N_11905,N_5757,N_8403);
xnor U11906 (N_11906,N_6624,N_6456);
nand U11907 (N_11907,N_6897,N_6719);
or U11908 (N_11908,N_6794,N_7205);
nor U11909 (N_11909,N_5803,N_5620);
nand U11910 (N_11910,N_7368,N_5230);
and U11911 (N_11911,N_5326,N_8591);
and U11912 (N_11912,N_8208,N_5295);
xor U11913 (N_11913,N_9992,N_7323);
xnor U11914 (N_11914,N_6310,N_8653);
or U11915 (N_11915,N_9707,N_7837);
and U11916 (N_11916,N_5603,N_7589);
nor U11917 (N_11917,N_6190,N_6744);
xnor U11918 (N_11918,N_9265,N_8708);
xnor U11919 (N_11919,N_9691,N_8187);
and U11920 (N_11920,N_6144,N_6357);
nor U11921 (N_11921,N_9774,N_8382);
and U11922 (N_11922,N_5566,N_7379);
nand U11923 (N_11923,N_5428,N_8410);
xor U11924 (N_11924,N_5973,N_7554);
nand U11925 (N_11925,N_6581,N_8044);
nand U11926 (N_11926,N_7277,N_6024);
xor U11927 (N_11927,N_9683,N_9338);
xnor U11928 (N_11928,N_9055,N_6439);
xor U11929 (N_11929,N_7214,N_6801);
nor U11930 (N_11930,N_5736,N_5555);
xor U11931 (N_11931,N_8532,N_9087);
xnor U11932 (N_11932,N_5399,N_7322);
and U11933 (N_11933,N_5958,N_7372);
and U11934 (N_11934,N_9085,N_7423);
nand U11935 (N_11935,N_5372,N_6353);
or U11936 (N_11936,N_7416,N_5046);
or U11937 (N_11937,N_8574,N_7896);
or U11938 (N_11938,N_5264,N_8969);
nor U11939 (N_11939,N_8102,N_7359);
nand U11940 (N_11940,N_6695,N_6979);
nor U11941 (N_11941,N_8633,N_9454);
nor U11942 (N_11942,N_9356,N_7257);
nand U11943 (N_11943,N_8194,N_8667);
xnor U11944 (N_11944,N_6819,N_9697);
xnor U11945 (N_11945,N_9218,N_5199);
nand U11946 (N_11946,N_5327,N_5146);
and U11947 (N_11947,N_5286,N_9297);
or U11948 (N_11948,N_9369,N_6986);
nand U11949 (N_11949,N_9348,N_7114);
nand U11950 (N_11950,N_9362,N_7953);
or U11951 (N_11951,N_5530,N_9358);
nor U11952 (N_11952,N_8719,N_7723);
or U11953 (N_11953,N_9616,N_6029);
and U11954 (N_11954,N_7819,N_7946);
xnor U11955 (N_11955,N_7705,N_7813);
xnor U11956 (N_11956,N_7370,N_9853);
nand U11957 (N_11957,N_9785,N_9928);
nor U11958 (N_11958,N_8871,N_6829);
nor U11959 (N_11959,N_5804,N_9820);
or U11960 (N_11960,N_9346,N_5517);
nor U11961 (N_11961,N_5975,N_6996);
and U11962 (N_11962,N_6773,N_8673);
nor U11963 (N_11963,N_6170,N_9166);
nand U11964 (N_11964,N_8188,N_9074);
xor U11965 (N_11965,N_5271,N_8287);
nor U11966 (N_11966,N_8101,N_8049);
nand U11967 (N_11967,N_8817,N_8407);
or U11968 (N_11968,N_5492,N_8892);
or U11969 (N_11969,N_5591,N_7985);
and U11970 (N_11970,N_5051,N_9291);
or U11971 (N_11971,N_5479,N_5161);
xnor U11972 (N_11972,N_9067,N_8415);
and U11973 (N_11973,N_9886,N_9546);
nor U11974 (N_11974,N_5785,N_9763);
and U11975 (N_11975,N_5789,N_7329);
nand U11976 (N_11976,N_9790,N_6955);
nor U11977 (N_11977,N_8394,N_5696);
nand U11978 (N_11978,N_8640,N_6162);
nand U11979 (N_11979,N_5979,N_6804);
and U11980 (N_11980,N_8681,N_7712);
nor U11981 (N_11981,N_7580,N_7974);
xor U11982 (N_11982,N_5818,N_6505);
xor U11983 (N_11983,N_5341,N_7719);
nor U11984 (N_11984,N_9266,N_6887);
nor U11985 (N_11985,N_5778,N_9376);
xnor U11986 (N_11986,N_9868,N_9270);
nor U11987 (N_11987,N_5233,N_9940);
nor U11988 (N_11988,N_5143,N_6515);
nor U11989 (N_11989,N_6039,N_6356);
and U11990 (N_11990,N_7201,N_8373);
and U11991 (N_11991,N_5385,N_6435);
or U11992 (N_11992,N_8597,N_7800);
xor U11993 (N_11993,N_9603,N_5016);
and U11994 (N_11994,N_7061,N_7871);
xor U11995 (N_11995,N_8943,N_5813);
and U11996 (N_11996,N_6498,N_9770);
nor U11997 (N_11997,N_6316,N_6425);
and U11998 (N_11998,N_6361,N_8530);
and U11999 (N_11999,N_5474,N_6925);
nand U12000 (N_12000,N_6340,N_8500);
xor U12001 (N_12001,N_5115,N_6147);
nand U12002 (N_12002,N_8557,N_9159);
or U12003 (N_12003,N_6707,N_5601);
nand U12004 (N_12004,N_5666,N_7764);
or U12005 (N_12005,N_8381,N_5909);
and U12006 (N_12006,N_7894,N_7507);
nor U12007 (N_12007,N_5191,N_8220);
nand U12008 (N_12008,N_9073,N_5024);
xnor U12009 (N_12009,N_7564,N_9476);
nor U12010 (N_12010,N_7112,N_8717);
and U12011 (N_12011,N_8909,N_8350);
or U12012 (N_12012,N_8245,N_6856);
and U12013 (N_12013,N_7155,N_8906);
and U12014 (N_12014,N_7579,N_6467);
nor U12015 (N_12015,N_8011,N_6539);
nand U12016 (N_12016,N_7674,N_7620);
xnor U12017 (N_12017,N_7176,N_7867);
and U12018 (N_12018,N_8729,N_8881);
xnor U12019 (N_12019,N_5716,N_5923);
xor U12020 (N_12020,N_8356,N_6655);
nand U12021 (N_12021,N_6429,N_5791);
xor U12022 (N_12022,N_9083,N_5797);
xor U12023 (N_12023,N_7908,N_7959);
xnor U12024 (N_12024,N_5114,N_9570);
nor U12025 (N_12025,N_9165,N_9607);
or U12026 (N_12026,N_7040,N_5499);
nand U12027 (N_12027,N_6945,N_6043);
or U12028 (N_12028,N_7098,N_5734);
or U12029 (N_12029,N_5772,N_7577);
and U12030 (N_12030,N_6517,N_7188);
nor U12031 (N_12031,N_5970,N_6036);
and U12032 (N_12032,N_9379,N_7778);
or U12033 (N_12033,N_8455,N_5425);
and U12034 (N_12034,N_7298,N_6481);
xor U12035 (N_12035,N_7687,N_7485);
and U12036 (N_12036,N_7239,N_6923);
xor U12037 (N_12037,N_7207,N_9738);
nor U12038 (N_12038,N_6445,N_9396);
and U12039 (N_12039,N_6917,N_5312);
or U12040 (N_12040,N_8096,N_8331);
and U12041 (N_12041,N_7491,N_7698);
xor U12042 (N_12042,N_6403,N_7237);
or U12043 (N_12043,N_7473,N_8575);
nor U12044 (N_12044,N_8676,N_5318);
and U12045 (N_12045,N_5607,N_7621);
and U12046 (N_12046,N_9328,N_5506);
or U12047 (N_12047,N_8465,N_5957);
nand U12048 (N_12048,N_6980,N_7581);
xnor U12049 (N_12049,N_5745,N_9761);
xnor U12050 (N_12050,N_6520,N_5488);
nand U12051 (N_12051,N_6944,N_8075);
or U12052 (N_12052,N_5602,N_7718);
and U12053 (N_12053,N_7667,N_7335);
nor U12054 (N_12054,N_9063,N_6537);
nor U12055 (N_12055,N_5825,N_8514);
or U12056 (N_12056,N_5080,N_7895);
or U12057 (N_12057,N_5369,N_8249);
nand U12058 (N_12058,N_7866,N_7196);
nor U12059 (N_12059,N_5635,N_8572);
nand U12060 (N_12060,N_7666,N_8108);
xor U12061 (N_12061,N_6994,N_7050);
xnor U12062 (N_12062,N_6696,N_9933);
nor U12063 (N_12063,N_8003,N_8181);
or U12064 (N_12064,N_9549,N_6836);
xnor U12065 (N_12065,N_5954,N_5984);
nand U12066 (N_12066,N_8583,N_6552);
nor U12067 (N_12067,N_9156,N_8628);
or U12068 (N_12068,N_6238,N_5961);
or U12069 (N_12069,N_5142,N_8339);
nor U12070 (N_12070,N_6633,N_6479);
nand U12071 (N_12071,N_5304,N_8482);
xor U12072 (N_12072,N_6421,N_7525);
or U12073 (N_12073,N_6511,N_7208);
or U12074 (N_12074,N_9331,N_7509);
or U12075 (N_12075,N_7663,N_6529);
and U12076 (N_12076,N_7924,N_8568);
and U12077 (N_12077,N_8483,N_9736);
and U12078 (N_12078,N_8710,N_9509);
nor U12079 (N_12079,N_9586,N_8215);
and U12080 (N_12080,N_9844,N_5766);
and U12081 (N_12081,N_7115,N_7119);
or U12082 (N_12082,N_9776,N_8967);
nand U12083 (N_12083,N_6431,N_5229);
and U12084 (N_12084,N_5924,N_8850);
xor U12085 (N_12085,N_8393,N_5939);
xor U12086 (N_12086,N_9827,N_6971);
and U12087 (N_12087,N_5240,N_9930);
xnor U12088 (N_12088,N_6315,N_8007);
nand U12089 (N_12089,N_8577,N_6482);
nor U12090 (N_12090,N_7899,N_9969);
or U12091 (N_12091,N_8887,N_9470);
and U12092 (N_12092,N_9070,N_7518);
or U12093 (N_12093,N_7308,N_8737);
nor U12094 (N_12094,N_6347,N_8050);
or U12095 (N_12095,N_9001,N_6196);
nand U12096 (N_12096,N_7662,N_6155);
nand U12097 (N_12097,N_7872,N_5001);
and U12098 (N_12098,N_7425,N_7410);
nand U12099 (N_12099,N_6269,N_7925);
xor U12100 (N_12100,N_9547,N_9804);
xnor U12101 (N_12101,N_5437,N_5148);
and U12102 (N_12102,N_5651,N_8660);
nor U12103 (N_12103,N_8303,N_7463);
and U12104 (N_12104,N_8335,N_8212);
nor U12105 (N_12105,N_5586,N_5702);
or U12106 (N_12106,N_7873,N_8126);
and U12107 (N_12107,N_8497,N_5008);
xor U12108 (N_12108,N_7008,N_7852);
xnor U12109 (N_12109,N_9884,N_7057);
nand U12110 (N_12110,N_5185,N_9000);
nand U12111 (N_12111,N_6956,N_6703);
nor U12112 (N_12112,N_6795,N_8152);
xnor U12113 (N_12113,N_7629,N_9955);
or U12114 (N_12114,N_7929,N_5814);
and U12115 (N_12115,N_9116,N_9717);
or U12116 (N_12116,N_5225,N_8678);
nor U12117 (N_12117,N_8630,N_8337);
or U12118 (N_12118,N_8092,N_7350);
nor U12119 (N_12119,N_5943,N_6922);
and U12120 (N_12120,N_8136,N_5773);
nand U12121 (N_12121,N_7316,N_8982);
xnor U12122 (N_12122,N_6301,N_6200);
xnor U12123 (N_12123,N_5032,N_6119);
and U12124 (N_12124,N_8413,N_7884);
nand U12125 (N_12125,N_8868,N_5121);
nand U12126 (N_12126,N_8764,N_9726);
nand U12127 (N_12127,N_8928,N_9150);
or U12128 (N_12128,N_6415,N_9571);
or U12129 (N_12129,N_6967,N_7266);
and U12130 (N_12130,N_8721,N_6577);
and U12131 (N_12131,N_9742,N_7568);
xnor U12132 (N_12132,N_5456,N_8792);
xor U12133 (N_12133,N_8677,N_5411);
nand U12134 (N_12134,N_8780,N_7193);
and U12135 (N_12135,N_9170,N_5982);
xor U12136 (N_12136,N_7998,N_7309);
and U12137 (N_12137,N_8730,N_9865);
xor U12138 (N_12138,N_8460,N_8095);
xor U12139 (N_12139,N_6249,N_6874);
nand U12140 (N_12140,N_8424,N_5289);
nand U12141 (N_12141,N_5335,N_6077);
and U12142 (N_12142,N_7377,N_6929);
and U12143 (N_12143,N_6555,N_7547);
or U12144 (N_12144,N_5887,N_9488);
and U12145 (N_12145,N_9781,N_7096);
or U12146 (N_12146,N_5820,N_6965);
and U12147 (N_12147,N_8008,N_6187);
or U12148 (N_12148,N_6553,N_8132);
or U12149 (N_12149,N_7439,N_9325);
xor U12150 (N_12150,N_7715,N_6358);
xor U12151 (N_12151,N_5665,N_7717);
or U12152 (N_12152,N_8211,N_5122);
and U12153 (N_12153,N_5725,N_8264);
or U12154 (N_12154,N_7915,N_8112);
nand U12155 (N_12155,N_5525,N_6673);
nor U12156 (N_12156,N_9304,N_9876);
or U12157 (N_12157,N_7027,N_8310);
and U12158 (N_12158,N_6828,N_8622);
and U12159 (N_12159,N_6115,N_8434);
or U12160 (N_12160,N_6964,N_5005);
and U12161 (N_12161,N_8870,N_7420);
xor U12162 (N_12162,N_7490,N_7583);
and U12163 (N_12163,N_6379,N_8010);
or U12164 (N_12164,N_8146,N_6006);
nor U12165 (N_12165,N_6188,N_9725);
and U12166 (N_12166,N_6637,N_5659);
nor U12167 (N_12167,N_7727,N_9251);
and U12168 (N_12168,N_6991,N_7049);
or U12169 (N_12169,N_8314,N_5413);
and U12170 (N_12170,N_7855,N_7874);
nor U12171 (N_12171,N_9390,N_9751);
or U12172 (N_12172,N_9670,N_9440);
or U12173 (N_12173,N_8355,N_6094);
nand U12174 (N_12174,N_9500,N_8526);
or U12175 (N_12175,N_6108,N_7154);
xor U12176 (N_12176,N_9140,N_9416);
and U12177 (N_12177,N_6195,N_5935);
xnor U12178 (N_12178,N_8369,N_9102);
nor U12179 (N_12179,N_6139,N_8897);
or U12180 (N_12180,N_6427,N_9668);
xor U12181 (N_12181,N_6158,N_8585);
nand U12182 (N_12182,N_8153,N_8131);
xnor U12183 (N_12183,N_6542,N_5515);
nor U12184 (N_12184,N_8754,N_6540);
nor U12185 (N_12185,N_9976,N_9057);
nand U12186 (N_12186,N_7337,N_5287);
or U12187 (N_12187,N_8171,N_7487);
xor U12188 (N_12188,N_9323,N_8499);
or U12189 (N_12189,N_7198,N_5760);
and U12190 (N_12190,N_6947,N_9968);
xnor U12191 (N_12191,N_5689,N_6469);
xor U12192 (N_12192,N_7875,N_5058);
nand U12193 (N_12193,N_6004,N_9182);
and U12194 (N_12194,N_5951,N_6216);
xnor U12195 (N_12195,N_6109,N_9153);
nand U12196 (N_12196,N_7168,N_8430);
xnor U12197 (N_12197,N_8877,N_8342);
or U12198 (N_12198,N_6179,N_8533);
nor U12199 (N_12199,N_8196,N_6648);
and U12200 (N_12200,N_5194,N_9508);
nor U12201 (N_12201,N_8891,N_9493);
xnor U12202 (N_12202,N_6838,N_6375);
and U12203 (N_12203,N_5187,N_9564);
nor U12204 (N_12204,N_6323,N_6450);
nand U12205 (N_12205,N_7364,N_8665);
or U12206 (N_12206,N_5573,N_6173);
nor U12207 (N_12207,N_9174,N_9313);
nor U12208 (N_12208,N_7788,N_6350);
xnor U12209 (N_12209,N_9112,N_5554);
nand U12210 (N_12210,N_9381,N_5599);
or U12211 (N_12211,N_7860,N_5572);
and U12212 (N_12212,N_9134,N_6545);
nand U12213 (N_12213,N_6372,N_9921);
or U12214 (N_12214,N_5087,N_5551);
xor U12215 (N_12215,N_9201,N_7465);
or U12216 (N_12216,N_8014,N_9715);
xor U12217 (N_12217,N_7823,N_9730);
or U12218 (N_12218,N_9991,N_7832);
xor U12219 (N_12219,N_5540,N_6044);
or U12220 (N_12220,N_5123,N_7643);
or U12221 (N_12221,N_9542,N_5489);
nand U12222 (N_12222,N_5231,N_5463);
nor U12223 (N_12223,N_9209,N_8299);
and U12224 (N_12224,N_6125,N_6858);
nand U12225 (N_12225,N_8123,N_5750);
and U12226 (N_12226,N_6714,N_7356);
and U12227 (N_12227,N_7341,N_7775);
nand U12228 (N_12228,N_5188,N_6627);
or U12229 (N_12229,N_6140,N_9596);
nand U12230 (N_12230,N_5221,N_6821);
nand U12231 (N_12231,N_7610,N_6595);
nor U12232 (N_12232,N_6727,N_5748);
nand U12233 (N_12233,N_9428,N_5912);
nand U12234 (N_12234,N_7226,N_5821);
xnor U12235 (N_12235,N_8405,N_7923);
or U12236 (N_12236,N_6319,N_5466);
nor U12237 (N_12237,N_5172,N_6283);
and U12238 (N_12238,N_6924,N_9290);
nor U12239 (N_12239,N_5908,N_8028);
or U12240 (N_12240,N_5708,N_6091);
xor U12241 (N_12241,N_9342,N_7153);
and U12242 (N_12242,N_6961,N_5018);
or U12243 (N_12243,N_6754,N_6653);
and U12244 (N_12244,N_6936,N_9031);
nand U12245 (N_12245,N_5742,N_9206);
nor U12246 (N_12246,N_6066,N_9732);
nor U12247 (N_12247,N_7271,N_9494);
xor U12248 (N_12248,N_7863,N_9408);
nor U12249 (N_12249,N_8820,N_8907);
nor U12250 (N_12250,N_5154,N_9446);
nor U12251 (N_12251,N_6919,N_5624);
and U12252 (N_12252,N_8529,N_8904);
and U12253 (N_12253,N_9838,N_7366);
nand U12254 (N_12254,N_5396,N_5721);
and U12255 (N_12255,N_6228,N_8246);
or U12256 (N_12256,N_9273,N_7931);
or U12257 (N_12257,N_7841,N_5449);
xnor U12258 (N_12258,N_6103,N_8372);
nor U12259 (N_12259,N_7135,N_6593);
or U12260 (N_12260,N_8760,N_8478);
xor U12261 (N_12261,N_8227,N_8312);
nor U12262 (N_12262,N_6534,N_5004);
xnor U12263 (N_12263,N_8317,N_5138);
xor U12264 (N_12264,N_9231,N_6003);
and U12265 (N_12265,N_6797,N_8922);
nand U12266 (N_12266,N_8902,N_7768);
nand U12267 (N_12267,N_8266,N_8668);
nor U12268 (N_12268,N_6940,N_7720);
xor U12269 (N_12269,N_5407,N_8239);
nand U12270 (N_12270,N_6619,N_8207);
nor U12271 (N_12271,N_8915,N_8359);
or U12272 (N_12272,N_8020,N_7601);
nor U12273 (N_12273,N_9980,N_6946);
xor U12274 (N_12274,N_7664,N_8379);
nor U12275 (N_12275,N_6016,N_5729);
nor U12276 (N_12276,N_5585,N_5512);
or U12277 (N_12277,N_9404,N_8600);
nor U12278 (N_12278,N_9195,N_8960);
or U12279 (N_12279,N_5843,N_6242);
nor U12280 (N_12280,N_9997,N_7054);
nor U12281 (N_12281,N_8779,N_9456);
nand U12282 (N_12282,N_8761,N_6762);
nor U12283 (N_12283,N_8692,N_5798);
and U12284 (N_12284,N_7278,N_6484);
nand U12285 (N_12285,N_7688,N_6404);
xor U12286 (N_12286,N_8596,N_6300);
and U12287 (N_12287,N_5673,N_7299);
and U12288 (N_12288,N_9403,N_7282);
or U12289 (N_12289,N_5829,N_9303);
and U12290 (N_12290,N_7947,N_9132);
xor U12291 (N_12291,N_5317,N_8635);
nand U12292 (N_12292,N_9337,N_7640);
and U12293 (N_12293,N_7421,N_7150);
xnor U12294 (N_12294,N_7177,N_6458);
and U12295 (N_12295,N_5223,N_8449);
and U12296 (N_12296,N_9753,N_7882);
xnor U12297 (N_12297,N_6521,N_5091);
or U12298 (N_12298,N_6121,N_6532);
nand U12299 (N_12299,N_9143,N_7446);
or U12300 (N_12300,N_7048,N_7126);
nand U12301 (N_12301,N_9833,N_7314);
xnor U12302 (N_12302,N_5853,N_8240);
nor U12303 (N_12303,N_7905,N_9537);
nand U12304 (N_12304,N_8156,N_9016);
xor U12305 (N_12305,N_7136,N_7095);
nor U12306 (N_12306,N_8866,N_9234);
or U12307 (N_12307,N_5366,N_9474);
nor U12308 (N_12308,N_7109,N_6234);
nor U12309 (N_12309,N_5876,N_9391);
or U12310 (N_12310,N_7032,N_8304);
xor U12311 (N_12311,N_8082,N_6683);
nand U12312 (N_12312,N_5026,N_5314);
and U12313 (N_12313,N_8062,N_9436);
nand U12314 (N_12314,N_9499,N_5422);
and U12315 (N_12315,N_6690,N_8746);
nand U12316 (N_12316,N_8280,N_9832);
or U12317 (N_12317,N_8796,N_5483);
and U12318 (N_12318,N_7969,N_8835);
nand U12319 (N_12319,N_6844,N_9335);
or U12320 (N_12320,N_5808,N_7415);
nor U12321 (N_12321,N_8164,N_7413);
or U12322 (N_12322,N_7966,N_8009);
or U12323 (N_12323,N_9027,N_7058);
or U12324 (N_12324,N_7575,N_7256);
and U12325 (N_12325,N_5679,N_8166);
and U12326 (N_12326,N_5035,N_8513);
and U12327 (N_12327,N_7315,N_8213);
nor U12328 (N_12328,N_7661,N_5684);
nand U12329 (N_12329,N_7123,N_6362);
nand U12330 (N_12330,N_7204,N_8421);
xnor U12331 (N_12331,N_5897,N_9772);
nand U12332 (N_12332,N_5397,N_7614);
nor U12333 (N_12333,N_9613,N_9256);
or U12334 (N_12334,N_9103,N_8275);
nor U12335 (N_12335,N_8012,N_7810);
or U12336 (N_12336,N_8615,N_5502);
nand U12337 (N_12337,N_8592,N_6490);
or U12338 (N_12338,N_8440,N_8221);
nand U12339 (N_12339,N_9714,N_8888);
nor U12340 (N_12340,N_8546,N_9489);
and U12341 (N_12341,N_8935,N_5382);
xnor U12342 (N_12342,N_6178,N_9932);
or U12343 (N_12343,N_6535,N_5692);
nor U12344 (N_12344,N_8016,N_8745);
nand U12345 (N_12345,N_9559,N_5027);
nor U12346 (N_12346,N_9118,N_6432);
nor U12347 (N_12347,N_7396,N_8389);
or U12348 (N_12348,N_6718,N_8755);
xnor U12349 (N_12349,N_6367,N_7118);
nor U12350 (N_12350,N_7325,N_6495);
nor U12351 (N_12351,N_8861,N_5494);
xor U12352 (N_12352,N_6687,N_7217);
or U12353 (N_12353,N_8311,N_8222);
or U12354 (N_12354,N_5612,N_7276);
xor U12355 (N_12355,N_6547,N_6602);
xnor U12356 (N_12356,N_8918,N_5134);
xnor U12357 (N_12357,N_6167,N_6394);
and U12358 (N_12358,N_9036,N_5446);
nor U12359 (N_12359,N_8802,N_6104);
or U12360 (N_12360,N_7326,N_6243);
xnor U12361 (N_12361,N_9451,N_6536);
nor U12362 (N_12362,N_7983,N_6989);
and U12363 (N_12363,N_6988,N_6785);
nand U12364 (N_12364,N_5465,N_7973);
nand U12365 (N_12365,N_7740,N_8402);
and U12366 (N_12366,N_8757,N_9722);
or U12367 (N_12367,N_9058,N_8923);
nand U12368 (N_12368,N_6264,N_9686);
xor U12369 (N_12369,N_5462,N_8081);
or U12370 (N_12370,N_9920,N_5331);
nor U12371 (N_12371,N_6670,N_7430);
nand U12372 (N_12372,N_9956,N_6254);
xnor U12373 (N_12373,N_5581,N_6800);
and U12374 (N_12374,N_8290,N_7288);
nor U12375 (N_12375,N_8441,N_6148);
xor U12376 (N_12376,N_8408,N_9667);
and U12377 (N_12377,N_9614,N_7728);
xnor U12378 (N_12378,N_7906,N_7968);
and U12379 (N_12379,N_6080,N_5675);
nand U12380 (N_12380,N_9825,N_8296);
nor U12381 (N_12381,N_5888,N_9459);
nor U12382 (N_12382,N_7677,N_7501);
xor U12383 (N_12383,N_5041,N_9017);
or U12384 (N_12384,N_8450,N_5706);
or U12385 (N_12385,N_7393,N_6159);
nand U12386 (N_12386,N_9392,N_8998);
and U12387 (N_12387,N_8963,N_5646);
and U12388 (N_12388,N_9705,N_5971);
and U12389 (N_12389,N_5946,N_5294);
or U12390 (N_12390,N_9882,N_6597);
nor U12391 (N_12391,N_8607,N_6914);
nor U12392 (N_12392,N_5039,N_5538);
xnor U12393 (N_12393,N_7551,N_6780);
nor U12394 (N_12394,N_7248,N_7962);
nand U12395 (N_12395,N_7488,N_9756);
or U12396 (N_12396,N_6303,N_8921);
and U12397 (N_12397,N_6031,N_9107);
and U12398 (N_12398,N_5649,N_5504);
nand U12399 (N_12399,N_7984,N_6755);
and U12400 (N_12400,N_6143,N_9522);
or U12401 (N_12401,N_6628,N_6071);
nand U12402 (N_12402,N_9448,N_5232);
nor U12403 (N_12403,N_5527,N_9129);
nor U12404 (N_12404,N_8068,N_7244);
xnor U12405 (N_12405,N_9771,N_6634);
or U12406 (N_12406,N_7066,N_5838);
xor U12407 (N_12407,N_6275,N_7826);
xor U12408 (N_12408,N_8197,N_8278);
nand U12409 (N_12409,N_7000,N_5064);
nand U12410 (N_12410,N_7191,N_5159);
nand U12411 (N_12411,N_6622,N_7786);
nor U12412 (N_12412,N_8486,N_9257);
and U12413 (N_12413,N_7023,N_9740);
and U12414 (N_12414,N_5067,N_8531);
nand U12415 (N_12415,N_9400,N_6128);
and U12416 (N_12416,N_8124,N_5600);
or U12417 (N_12417,N_5364,N_6410);
and U12418 (N_12418,N_7231,N_8469);
or U12419 (N_12419,N_9769,N_5263);
nor U12420 (N_12420,N_5092,N_6359);
nand U12421 (N_12421,N_7502,N_9411);
and U12422 (N_12422,N_7014,N_9941);
nand U12423 (N_12423,N_8899,N_6793);
or U12424 (N_12424,N_5478,N_6120);
nand U12425 (N_12425,N_6667,N_5655);
or U12426 (N_12426,N_7262,N_5309);
nor U12427 (N_12427,N_6496,N_5017);
nor U12428 (N_12428,N_9674,N_8713);
and U12429 (N_12429,N_8427,N_6007);
nand U12430 (N_12430,N_7690,N_5691);
and U12431 (N_12431,N_7503,N_7417);
nand U12432 (N_12432,N_9312,N_9764);
xnor U12433 (N_12433,N_6859,N_9869);
nand U12434 (N_12434,N_9525,N_5118);
nand U12435 (N_12435,N_9370,N_5131);
or U12436 (N_12436,N_8343,N_9177);
nand U12437 (N_12437,N_6258,N_6816);
nor U12438 (N_12438,N_6580,N_8976);
and U12439 (N_12439,N_6393,N_6759);
nand U12440 (N_12440,N_5636,N_8537);
nand U12441 (N_12441,N_6745,N_6442);
and U12442 (N_12442,N_8199,N_5549);
or U12443 (N_12443,N_6312,N_8248);
and U12444 (N_12444,N_6715,N_8217);
and U12445 (N_12445,N_6528,N_5930);
nor U12446 (N_12446,N_8809,N_9702);
or U12447 (N_12447,N_7481,N_9615);
nand U12448 (N_12448,N_8448,N_7716);
nand U12449 (N_12449,N_8345,N_5283);
nand U12450 (N_12450,N_8656,N_5023);
xnor U12451 (N_12451,N_7902,N_7999);
nand U12452 (N_12452,N_5879,N_8292);
and U12453 (N_12453,N_5583,N_6237);
nor U12454 (N_12454,N_7548,N_9745);
nand U12455 (N_12455,N_8743,N_9246);
or U12456 (N_12456,N_5190,N_6034);
nand U12457 (N_12457,N_7859,N_8154);
or U12458 (N_12458,N_9464,N_7757);
nand U12459 (N_12459,N_5994,N_5516);
xor U12460 (N_12460,N_5007,N_7230);
or U12461 (N_12461,N_8021,N_9477);
and U12462 (N_12462,N_8900,N_6073);
nand U12463 (N_12463,N_8177,N_8182);
nand U12464 (N_12464,N_8732,N_8090);
xnor U12465 (N_12465,N_6939,N_8970);
nand U12466 (N_12466,N_5297,N_6126);
xor U12467 (N_12467,N_7087,N_8594);
or U12468 (N_12468,N_6342,N_8774);
or U12469 (N_12469,N_5477,N_5155);
xor U12470 (N_12470,N_7582,N_8279);
nand U12471 (N_12471,N_9462,N_7753);
nor U12472 (N_12472,N_8038,N_8262);
xor U12473 (N_12473,N_5047,N_7958);
xor U12474 (N_12474,N_5932,N_9026);
xnor U12475 (N_12475,N_5203,N_6841);
xnor U12476 (N_12476,N_8964,N_6854);
or U12477 (N_12477,N_9157,N_5034);
xnor U12478 (N_12478,N_5094,N_5807);
nand U12479 (N_12479,N_6756,N_5333);
and U12480 (N_12480,N_5089,N_9673);
xor U12481 (N_12481,N_5800,N_6768);
xor U12482 (N_12482,N_5105,N_7235);
or U12483 (N_12483,N_9122,N_9426);
xnor U12484 (N_12484,N_7870,N_5401);
or U12485 (N_12485,N_6876,N_9437);
nor U12486 (N_12486,N_8981,N_5944);
nand U12487 (N_12487,N_5127,N_5652);
or U12488 (N_12488,N_9308,N_8134);
xnor U12489 (N_12489,N_7857,N_6512);
and U12490 (N_12490,N_7295,N_7409);
nand U12491 (N_12491,N_7339,N_5010);
xor U12492 (N_12492,N_6049,N_6730);
xnor U12493 (N_12493,N_6199,N_9999);
xor U12494 (N_12494,N_5917,N_7483);
nand U12495 (N_12495,N_6818,N_8360);
or U12496 (N_12496,N_7169,N_9646);
or U12497 (N_12497,N_8228,N_7447);
or U12498 (N_12498,N_5553,N_5974);
nor U12499 (N_12499,N_9849,N_6437);
nand U12500 (N_12500,N_5535,N_9914);
and U12501 (N_12501,N_9339,N_5456);
and U12502 (N_12502,N_6653,N_6726);
or U12503 (N_12503,N_9968,N_8850);
and U12504 (N_12504,N_5547,N_7704);
and U12505 (N_12505,N_8058,N_8708);
nand U12506 (N_12506,N_8486,N_9880);
nand U12507 (N_12507,N_8694,N_9729);
nand U12508 (N_12508,N_6790,N_8712);
and U12509 (N_12509,N_6587,N_7689);
or U12510 (N_12510,N_5356,N_5309);
nor U12511 (N_12511,N_9691,N_7928);
nand U12512 (N_12512,N_7973,N_5273);
and U12513 (N_12513,N_9104,N_5838);
nand U12514 (N_12514,N_9155,N_7458);
and U12515 (N_12515,N_5236,N_6840);
and U12516 (N_12516,N_7433,N_8393);
nand U12517 (N_12517,N_6711,N_9539);
or U12518 (N_12518,N_9463,N_9955);
nand U12519 (N_12519,N_5464,N_6239);
and U12520 (N_12520,N_9088,N_8292);
or U12521 (N_12521,N_8922,N_8566);
nor U12522 (N_12522,N_6302,N_6419);
nor U12523 (N_12523,N_9997,N_8045);
nor U12524 (N_12524,N_7224,N_6490);
nand U12525 (N_12525,N_9933,N_9839);
and U12526 (N_12526,N_7354,N_7268);
and U12527 (N_12527,N_5179,N_6034);
nand U12528 (N_12528,N_9079,N_8519);
xor U12529 (N_12529,N_8877,N_7920);
nand U12530 (N_12530,N_6229,N_6717);
xnor U12531 (N_12531,N_9245,N_9335);
xor U12532 (N_12532,N_8599,N_9320);
or U12533 (N_12533,N_5279,N_9114);
and U12534 (N_12534,N_6284,N_6350);
or U12535 (N_12535,N_9767,N_7578);
nand U12536 (N_12536,N_6524,N_9116);
and U12537 (N_12537,N_9756,N_5438);
or U12538 (N_12538,N_9145,N_5921);
nand U12539 (N_12539,N_8103,N_6253);
nand U12540 (N_12540,N_5910,N_7287);
or U12541 (N_12541,N_9345,N_8455);
and U12542 (N_12542,N_8700,N_6647);
xor U12543 (N_12543,N_7187,N_5776);
and U12544 (N_12544,N_6425,N_9145);
xnor U12545 (N_12545,N_8391,N_8328);
nor U12546 (N_12546,N_7544,N_6668);
or U12547 (N_12547,N_6626,N_7703);
or U12548 (N_12548,N_6266,N_9720);
nor U12549 (N_12549,N_5487,N_9376);
xnor U12550 (N_12550,N_5439,N_7392);
nand U12551 (N_12551,N_8434,N_9574);
xnor U12552 (N_12552,N_7199,N_8808);
nand U12553 (N_12553,N_6164,N_6439);
nand U12554 (N_12554,N_9266,N_8490);
xor U12555 (N_12555,N_9369,N_8258);
or U12556 (N_12556,N_8029,N_8882);
nor U12557 (N_12557,N_7726,N_9145);
nor U12558 (N_12558,N_7444,N_7752);
nand U12559 (N_12559,N_5587,N_9914);
and U12560 (N_12560,N_9451,N_9815);
or U12561 (N_12561,N_7756,N_5023);
nor U12562 (N_12562,N_9022,N_7593);
and U12563 (N_12563,N_9727,N_6260);
nor U12564 (N_12564,N_6877,N_6043);
xor U12565 (N_12565,N_8747,N_8650);
nand U12566 (N_12566,N_6843,N_6073);
xor U12567 (N_12567,N_8309,N_5225);
or U12568 (N_12568,N_7759,N_6554);
or U12569 (N_12569,N_6615,N_6741);
or U12570 (N_12570,N_9426,N_9363);
and U12571 (N_12571,N_7598,N_5949);
nand U12572 (N_12572,N_6234,N_5798);
xnor U12573 (N_12573,N_9575,N_9381);
and U12574 (N_12574,N_8298,N_7541);
nor U12575 (N_12575,N_7138,N_6552);
or U12576 (N_12576,N_5758,N_6442);
nand U12577 (N_12577,N_8805,N_8207);
nand U12578 (N_12578,N_7742,N_8454);
or U12579 (N_12579,N_7046,N_5616);
xor U12580 (N_12580,N_6658,N_9914);
nand U12581 (N_12581,N_9253,N_9315);
and U12582 (N_12582,N_6070,N_9315);
nand U12583 (N_12583,N_7193,N_9346);
and U12584 (N_12584,N_7312,N_5426);
nor U12585 (N_12585,N_9844,N_6150);
or U12586 (N_12586,N_9625,N_5511);
and U12587 (N_12587,N_7438,N_6674);
nand U12588 (N_12588,N_6524,N_9589);
and U12589 (N_12589,N_5664,N_5337);
or U12590 (N_12590,N_7649,N_8455);
nand U12591 (N_12591,N_7537,N_7613);
or U12592 (N_12592,N_6615,N_9158);
or U12593 (N_12593,N_9647,N_8708);
xnor U12594 (N_12594,N_6753,N_6138);
or U12595 (N_12595,N_7449,N_7133);
xnor U12596 (N_12596,N_7911,N_8244);
nor U12597 (N_12597,N_8308,N_7897);
or U12598 (N_12598,N_7368,N_9907);
or U12599 (N_12599,N_8707,N_6838);
or U12600 (N_12600,N_6687,N_6116);
nand U12601 (N_12601,N_8748,N_6501);
nor U12602 (N_12602,N_6956,N_7974);
and U12603 (N_12603,N_8706,N_7277);
xnor U12604 (N_12604,N_9222,N_7115);
or U12605 (N_12605,N_8221,N_5540);
nor U12606 (N_12606,N_8746,N_8796);
and U12607 (N_12607,N_7731,N_6000);
and U12608 (N_12608,N_5830,N_9573);
xor U12609 (N_12609,N_7822,N_6297);
xor U12610 (N_12610,N_5601,N_8070);
nand U12611 (N_12611,N_8763,N_6108);
or U12612 (N_12612,N_5847,N_6064);
nand U12613 (N_12613,N_9457,N_6153);
nand U12614 (N_12614,N_7172,N_8113);
nor U12615 (N_12615,N_9189,N_5675);
or U12616 (N_12616,N_6758,N_5172);
xnor U12617 (N_12617,N_5628,N_5676);
nand U12618 (N_12618,N_5613,N_9906);
xnor U12619 (N_12619,N_5876,N_6735);
and U12620 (N_12620,N_9642,N_9740);
and U12621 (N_12621,N_9154,N_8236);
or U12622 (N_12622,N_5615,N_9814);
xnor U12623 (N_12623,N_8271,N_9333);
xor U12624 (N_12624,N_7450,N_5783);
nor U12625 (N_12625,N_8553,N_9647);
or U12626 (N_12626,N_8224,N_8739);
and U12627 (N_12627,N_9741,N_5306);
xor U12628 (N_12628,N_7018,N_6382);
nand U12629 (N_12629,N_9654,N_8651);
nor U12630 (N_12630,N_9830,N_7345);
xor U12631 (N_12631,N_6791,N_5350);
nand U12632 (N_12632,N_8222,N_6245);
and U12633 (N_12633,N_7730,N_5583);
nand U12634 (N_12634,N_8435,N_9984);
or U12635 (N_12635,N_6269,N_9876);
nor U12636 (N_12636,N_8408,N_9310);
xor U12637 (N_12637,N_8189,N_5025);
or U12638 (N_12638,N_6984,N_9348);
nand U12639 (N_12639,N_7023,N_7356);
or U12640 (N_12640,N_7529,N_8969);
nand U12641 (N_12641,N_5822,N_9867);
or U12642 (N_12642,N_9033,N_9055);
or U12643 (N_12643,N_5682,N_6395);
xnor U12644 (N_12644,N_8224,N_9174);
or U12645 (N_12645,N_8378,N_6643);
and U12646 (N_12646,N_9420,N_5814);
xnor U12647 (N_12647,N_9481,N_9306);
nor U12648 (N_12648,N_9089,N_6818);
nor U12649 (N_12649,N_6638,N_8235);
and U12650 (N_12650,N_5946,N_6557);
and U12651 (N_12651,N_5306,N_7982);
or U12652 (N_12652,N_6356,N_6545);
nand U12653 (N_12653,N_9884,N_9862);
nand U12654 (N_12654,N_9819,N_6107);
nand U12655 (N_12655,N_7660,N_8736);
and U12656 (N_12656,N_5887,N_7932);
or U12657 (N_12657,N_5386,N_7073);
xnor U12658 (N_12658,N_6442,N_6830);
and U12659 (N_12659,N_9159,N_6110);
or U12660 (N_12660,N_5480,N_8832);
or U12661 (N_12661,N_5144,N_7991);
nand U12662 (N_12662,N_6044,N_5955);
or U12663 (N_12663,N_6191,N_5064);
xnor U12664 (N_12664,N_7546,N_5731);
nor U12665 (N_12665,N_5266,N_9758);
nand U12666 (N_12666,N_5399,N_8473);
or U12667 (N_12667,N_5859,N_7626);
nor U12668 (N_12668,N_5969,N_8527);
nand U12669 (N_12669,N_8975,N_8815);
nor U12670 (N_12670,N_9007,N_8033);
xnor U12671 (N_12671,N_5370,N_8052);
or U12672 (N_12672,N_8975,N_8009);
or U12673 (N_12673,N_7379,N_9170);
or U12674 (N_12674,N_8478,N_9213);
nor U12675 (N_12675,N_7223,N_8016);
xor U12676 (N_12676,N_8023,N_7350);
nor U12677 (N_12677,N_9200,N_9652);
nand U12678 (N_12678,N_9817,N_9696);
nor U12679 (N_12679,N_5310,N_7647);
nor U12680 (N_12680,N_8507,N_5980);
xnor U12681 (N_12681,N_9775,N_8648);
xnor U12682 (N_12682,N_7029,N_9464);
or U12683 (N_12683,N_9371,N_7067);
xor U12684 (N_12684,N_8450,N_8134);
and U12685 (N_12685,N_5129,N_6841);
and U12686 (N_12686,N_9569,N_6409);
nand U12687 (N_12687,N_5304,N_6677);
nand U12688 (N_12688,N_9296,N_6240);
nand U12689 (N_12689,N_8745,N_5150);
and U12690 (N_12690,N_8117,N_8074);
nand U12691 (N_12691,N_5334,N_6534);
nor U12692 (N_12692,N_5679,N_5920);
xor U12693 (N_12693,N_9836,N_9800);
nand U12694 (N_12694,N_5056,N_6670);
nand U12695 (N_12695,N_5182,N_9645);
nand U12696 (N_12696,N_5672,N_7170);
or U12697 (N_12697,N_8569,N_5857);
nor U12698 (N_12698,N_9453,N_8449);
nand U12699 (N_12699,N_5211,N_7469);
nor U12700 (N_12700,N_6857,N_5273);
nand U12701 (N_12701,N_6486,N_7082);
and U12702 (N_12702,N_6808,N_6124);
xor U12703 (N_12703,N_9429,N_9880);
xor U12704 (N_12704,N_8990,N_6023);
xor U12705 (N_12705,N_6310,N_7891);
xnor U12706 (N_12706,N_9264,N_5632);
xor U12707 (N_12707,N_6164,N_5360);
xor U12708 (N_12708,N_6285,N_5194);
or U12709 (N_12709,N_6090,N_6777);
and U12710 (N_12710,N_7099,N_6329);
nand U12711 (N_12711,N_7891,N_9279);
and U12712 (N_12712,N_9057,N_9469);
nor U12713 (N_12713,N_8743,N_6980);
nand U12714 (N_12714,N_6005,N_6258);
nand U12715 (N_12715,N_8636,N_6986);
nor U12716 (N_12716,N_9456,N_9868);
or U12717 (N_12717,N_8470,N_6807);
or U12718 (N_12718,N_6963,N_6763);
or U12719 (N_12719,N_5893,N_9639);
nand U12720 (N_12720,N_9824,N_5846);
nand U12721 (N_12721,N_5017,N_8749);
or U12722 (N_12722,N_9142,N_7457);
xor U12723 (N_12723,N_6980,N_5649);
nor U12724 (N_12724,N_8792,N_5655);
or U12725 (N_12725,N_7594,N_9074);
nand U12726 (N_12726,N_5786,N_9435);
xor U12727 (N_12727,N_5847,N_8058);
or U12728 (N_12728,N_6294,N_5655);
or U12729 (N_12729,N_5842,N_9556);
nor U12730 (N_12730,N_7984,N_8839);
nand U12731 (N_12731,N_7860,N_8793);
xnor U12732 (N_12732,N_6138,N_5080);
and U12733 (N_12733,N_7302,N_7872);
nand U12734 (N_12734,N_9046,N_5756);
nand U12735 (N_12735,N_5351,N_8796);
xnor U12736 (N_12736,N_9025,N_6881);
or U12737 (N_12737,N_5177,N_6551);
xnor U12738 (N_12738,N_8763,N_8685);
and U12739 (N_12739,N_7033,N_9755);
and U12740 (N_12740,N_7306,N_9362);
nand U12741 (N_12741,N_9990,N_9641);
xor U12742 (N_12742,N_9520,N_9850);
nand U12743 (N_12743,N_6199,N_5664);
nor U12744 (N_12744,N_6941,N_8985);
or U12745 (N_12745,N_7207,N_9892);
nand U12746 (N_12746,N_5129,N_7053);
and U12747 (N_12747,N_7509,N_9030);
or U12748 (N_12748,N_6798,N_7263);
xor U12749 (N_12749,N_9114,N_5606);
nand U12750 (N_12750,N_6835,N_5871);
nand U12751 (N_12751,N_9603,N_9858);
and U12752 (N_12752,N_5332,N_8914);
xor U12753 (N_12753,N_8039,N_8694);
and U12754 (N_12754,N_5966,N_7073);
nor U12755 (N_12755,N_7179,N_7593);
and U12756 (N_12756,N_8274,N_9542);
and U12757 (N_12757,N_6567,N_6666);
xnor U12758 (N_12758,N_7573,N_8110);
or U12759 (N_12759,N_7395,N_5868);
or U12760 (N_12760,N_6579,N_8777);
nand U12761 (N_12761,N_6581,N_5953);
nor U12762 (N_12762,N_9220,N_9483);
nand U12763 (N_12763,N_6922,N_9724);
and U12764 (N_12764,N_9582,N_9950);
nand U12765 (N_12765,N_8487,N_8681);
nor U12766 (N_12766,N_5404,N_8601);
and U12767 (N_12767,N_8887,N_6845);
and U12768 (N_12768,N_7235,N_5756);
xnor U12769 (N_12769,N_7408,N_8089);
nor U12770 (N_12770,N_9782,N_7983);
xor U12771 (N_12771,N_8607,N_6629);
xor U12772 (N_12772,N_8942,N_5621);
or U12773 (N_12773,N_5468,N_8550);
or U12774 (N_12774,N_9973,N_8595);
and U12775 (N_12775,N_6405,N_8738);
or U12776 (N_12776,N_5999,N_5129);
nand U12777 (N_12777,N_5772,N_5415);
xnor U12778 (N_12778,N_7585,N_6782);
xnor U12779 (N_12779,N_5583,N_5473);
or U12780 (N_12780,N_9487,N_8953);
and U12781 (N_12781,N_6817,N_6709);
nor U12782 (N_12782,N_6623,N_5315);
xor U12783 (N_12783,N_8059,N_6110);
or U12784 (N_12784,N_8625,N_5669);
xnor U12785 (N_12785,N_9744,N_9566);
and U12786 (N_12786,N_6880,N_5528);
xor U12787 (N_12787,N_8483,N_5880);
or U12788 (N_12788,N_5666,N_9975);
nand U12789 (N_12789,N_7485,N_5341);
nand U12790 (N_12790,N_9776,N_9544);
xnor U12791 (N_12791,N_7920,N_7576);
nor U12792 (N_12792,N_6746,N_5435);
or U12793 (N_12793,N_8808,N_9574);
or U12794 (N_12794,N_5095,N_6373);
nand U12795 (N_12795,N_5572,N_5422);
xnor U12796 (N_12796,N_6621,N_7739);
nor U12797 (N_12797,N_6135,N_9929);
and U12798 (N_12798,N_9789,N_9340);
nand U12799 (N_12799,N_8625,N_5813);
and U12800 (N_12800,N_9507,N_8899);
xor U12801 (N_12801,N_8893,N_9723);
and U12802 (N_12802,N_7751,N_9738);
nand U12803 (N_12803,N_5627,N_7795);
xnor U12804 (N_12804,N_9468,N_9966);
or U12805 (N_12805,N_5899,N_6697);
or U12806 (N_12806,N_7080,N_5437);
nor U12807 (N_12807,N_5572,N_5403);
nor U12808 (N_12808,N_5885,N_6592);
and U12809 (N_12809,N_9884,N_8201);
or U12810 (N_12810,N_5266,N_5878);
nand U12811 (N_12811,N_5477,N_7280);
and U12812 (N_12812,N_6860,N_9400);
nor U12813 (N_12813,N_7408,N_6074);
xor U12814 (N_12814,N_8001,N_9096);
xor U12815 (N_12815,N_8369,N_8979);
and U12816 (N_12816,N_6903,N_5739);
and U12817 (N_12817,N_9329,N_6207);
xor U12818 (N_12818,N_8406,N_7591);
nor U12819 (N_12819,N_6624,N_5475);
and U12820 (N_12820,N_7441,N_6946);
nor U12821 (N_12821,N_5608,N_6340);
xnor U12822 (N_12822,N_8823,N_7660);
xor U12823 (N_12823,N_8044,N_7293);
nor U12824 (N_12824,N_5111,N_5737);
nand U12825 (N_12825,N_8085,N_8349);
nand U12826 (N_12826,N_7111,N_7880);
nor U12827 (N_12827,N_7738,N_8220);
xnor U12828 (N_12828,N_7906,N_5830);
nand U12829 (N_12829,N_7002,N_6787);
nand U12830 (N_12830,N_7358,N_8211);
nand U12831 (N_12831,N_9382,N_9487);
nand U12832 (N_12832,N_7709,N_5204);
and U12833 (N_12833,N_8431,N_5514);
nor U12834 (N_12834,N_7024,N_7407);
nor U12835 (N_12835,N_5412,N_5660);
or U12836 (N_12836,N_9791,N_5944);
or U12837 (N_12837,N_8210,N_5308);
nor U12838 (N_12838,N_9311,N_9228);
nor U12839 (N_12839,N_5485,N_5433);
or U12840 (N_12840,N_9921,N_9993);
xnor U12841 (N_12841,N_9631,N_9183);
xor U12842 (N_12842,N_9803,N_7662);
nand U12843 (N_12843,N_8583,N_7404);
xor U12844 (N_12844,N_7020,N_9949);
nand U12845 (N_12845,N_9016,N_5518);
or U12846 (N_12846,N_6347,N_9230);
and U12847 (N_12847,N_6852,N_7518);
nand U12848 (N_12848,N_7369,N_6197);
and U12849 (N_12849,N_6681,N_6171);
or U12850 (N_12850,N_7088,N_7529);
or U12851 (N_12851,N_6218,N_7597);
xnor U12852 (N_12852,N_6831,N_5941);
nand U12853 (N_12853,N_6043,N_8233);
or U12854 (N_12854,N_8330,N_8596);
and U12855 (N_12855,N_8473,N_8999);
and U12856 (N_12856,N_7842,N_7633);
and U12857 (N_12857,N_5162,N_7302);
nor U12858 (N_12858,N_8015,N_5165);
xor U12859 (N_12859,N_5156,N_9147);
nand U12860 (N_12860,N_8609,N_8906);
or U12861 (N_12861,N_5488,N_5246);
or U12862 (N_12862,N_9300,N_5358);
or U12863 (N_12863,N_6461,N_7447);
or U12864 (N_12864,N_7190,N_5835);
nor U12865 (N_12865,N_8652,N_5323);
nand U12866 (N_12866,N_8014,N_6337);
nand U12867 (N_12867,N_5136,N_5716);
or U12868 (N_12868,N_6654,N_5301);
xor U12869 (N_12869,N_7002,N_6524);
xor U12870 (N_12870,N_5516,N_8624);
and U12871 (N_12871,N_5555,N_7685);
xnor U12872 (N_12872,N_8606,N_9550);
or U12873 (N_12873,N_6025,N_7786);
or U12874 (N_12874,N_5151,N_5849);
and U12875 (N_12875,N_8060,N_5041);
or U12876 (N_12876,N_5026,N_8778);
nor U12877 (N_12877,N_9023,N_6672);
xnor U12878 (N_12878,N_8116,N_7005);
and U12879 (N_12879,N_8516,N_6659);
and U12880 (N_12880,N_6256,N_8397);
xnor U12881 (N_12881,N_6586,N_8622);
or U12882 (N_12882,N_8335,N_5513);
xnor U12883 (N_12883,N_7486,N_5705);
xnor U12884 (N_12884,N_8139,N_9541);
and U12885 (N_12885,N_8389,N_8460);
nand U12886 (N_12886,N_6100,N_9661);
nor U12887 (N_12887,N_6006,N_5534);
or U12888 (N_12888,N_5020,N_7058);
and U12889 (N_12889,N_9579,N_5567);
or U12890 (N_12890,N_8823,N_5063);
or U12891 (N_12891,N_7202,N_8920);
or U12892 (N_12892,N_7700,N_7770);
nand U12893 (N_12893,N_7038,N_5828);
and U12894 (N_12894,N_6870,N_7467);
xnor U12895 (N_12895,N_8732,N_9786);
xnor U12896 (N_12896,N_7563,N_8295);
or U12897 (N_12897,N_8592,N_6695);
nor U12898 (N_12898,N_7462,N_5060);
xor U12899 (N_12899,N_7392,N_7345);
or U12900 (N_12900,N_8226,N_7072);
nand U12901 (N_12901,N_8856,N_5701);
xor U12902 (N_12902,N_7900,N_7258);
nand U12903 (N_12903,N_9888,N_9492);
or U12904 (N_12904,N_6502,N_6433);
xor U12905 (N_12905,N_5642,N_7660);
nand U12906 (N_12906,N_7977,N_6810);
or U12907 (N_12907,N_6564,N_7549);
xor U12908 (N_12908,N_7362,N_7507);
nor U12909 (N_12909,N_8758,N_8825);
nand U12910 (N_12910,N_6021,N_6604);
xnor U12911 (N_12911,N_6231,N_7495);
xnor U12912 (N_12912,N_9202,N_8552);
xnor U12913 (N_12913,N_6286,N_7194);
xor U12914 (N_12914,N_8845,N_8523);
nor U12915 (N_12915,N_7143,N_6143);
nand U12916 (N_12916,N_6269,N_9916);
or U12917 (N_12917,N_7441,N_8773);
nand U12918 (N_12918,N_7692,N_7820);
and U12919 (N_12919,N_9619,N_5664);
nand U12920 (N_12920,N_6588,N_8385);
nor U12921 (N_12921,N_5165,N_5538);
nor U12922 (N_12922,N_8286,N_7060);
xnor U12923 (N_12923,N_9343,N_7499);
xnor U12924 (N_12924,N_5572,N_5002);
or U12925 (N_12925,N_9518,N_7138);
nor U12926 (N_12926,N_6444,N_7607);
xnor U12927 (N_12927,N_6201,N_6675);
nand U12928 (N_12928,N_7609,N_8388);
nand U12929 (N_12929,N_5549,N_5301);
or U12930 (N_12930,N_6749,N_5283);
and U12931 (N_12931,N_7007,N_8302);
and U12932 (N_12932,N_7310,N_7063);
nand U12933 (N_12933,N_5179,N_8272);
nand U12934 (N_12934,N_7363,N_6210);
xor U12935 (N_12935,N_7187,N_9789);
and U12936 (N_12936,N_9360,N_6940);
nor U12937 (N_12937,N_5500,N_5788);
nand U12938 (N_12938,N_8304,N_8394);
or U12939 (N_12939,N_8312,N_8721);
xnor U12940 (N_12940,N_8979,N_6774);
xor U12941 (N_12941,N_6795,N_9531);
nand U12942 (N_12942,N_8964,N_7087);
nor U12943 (N_12943,N_5581,N_5222);
and U12944 (N_12944,N_5070,N_8294);
and U12945 (N_12945,N_6119,N_8694);
xnor U12946 (N_12946,N_8861,N_9162);
nor U12947 (N_12947,N_7087,N_6809);
xnor U12948 (N_12948,N_9691,N_8577);
nor U12949 (N_12949,N_5833,N_7830);
nor U12950 (N_12950,N_6855,N_6367);
or U12951 (N_12951,N_6459,N_7296);
xnor U12952 (N_12952,N_6256,N_6123);
xor U12953 (N_12953,N_7672,N_9805);
or U12954 (N_12954,N_6468,N_7112);
xnor U12955 (N_12955,N_5946,N_9250);
xnor U12956 (N_12956,N_6519,N_9008);
or U12957 (N_12957,N_8639,N_6673);
or U12958 (N_12958,N_9599,N_5745);
and U12959 (N_12959,N_8468,N_9154);
nand U12960 (N_12960,N_9472,N_5405);
xnor U12961 (N_12961,N_9705,N_8724);
xor U12962 (N_12962,N_7681,N_9122);
nand U12963 (N_12963,N_7123,N_8439);
xor U12964 (N_12964,N_9065,N_5381);
nor U12965 (N_12965,N_9775,N_9943);
nor U12966 (N_12966,N_5014,N_8923);
or U12967 (N_12967,N_5021,N_9866);
nor U12968 (N_12968,N_7056,N_7267);
and U12969 (N_12969,N_6375,N_9987);
nor U12970 (N_12970,N_9001,N_6504);
nor U12971 (N_12971,N_8876,N_8330);
or U12972 (N_12972,N_7942,N_8212);
nor U12973 (N_12973,N_7653,N_8701);
xor U12974 (N_12974,N_7569,N_6924);
nand U12975 (N_12975,N_8719,N_5015);
nor U12976 (N_12976,N_9087,N_7512);
nand U12977 (N_12977,N_9864,N_9598);
and U12978 (N_12978,N_5779,N_9084);
xnor U12979 (N_12979,N_8107,N_9624);
nor U12980 (N_12980,N_6967,N_6791);
xnor U12981 (N_12981,N_7429,N_6235);
nor U12982 (N_12982,N_7704,N_5863);
or U12983 (N_12983,N_5932,N_8083);
nor U12984 (N_12984,N_6434,N_7843);
nand U12985 (N_12985,N_7771,N_5863);
nand U12986 (N_12986,N_8718,N_7628);
or U12987 (N_12987,N_6573,N_9999);
nand U12988 (N_12988,N_5048,N_5562);
xnor U12989 (N_12989,N_6609,N_8178);
and U12990 (N_12990,N_7941,N_9810);
and U12991 (N_12991,N_6347,N_8292);
or U12992 (N_12992,N_8382,N_5409);
or U12993 (N_12993,N_9300,N_9042);
nand U12994 (N_12994,N_5995,N_5543);
xnor U12995 (N_12995,N_6768,N_9886);
xor U12996 (N_12996,N_6498,N_8767);
xnor U12997 (N_12997,N_5827,N_7475);
and U12998 (N_12998,N_7834,N_8251);
xor U12999 (N_12999,N_6721,N_5474);
and U13000 (N_13000,N_5077,N_7181);
nand U13001 (N_13001,N_6998,N_6704);
or U13002 (N_13002,N_7581,N_5660);
nand U13003 (N_13003,N_8812,N_6145);
xnor U13004 (N_13004,N_5717,N_9145);
and U13005 (N_13005,N_5864,N_8367);
nand U13006 (N_13006,N_5887,N_8815);
xnor U13007 (N_13007,N_6009,N_6757);
xnor U13008 (N_13008,N_8101,N_8578);
or U13009 (N_13009,N_8799,N_8421);
nor U13010 (N_13010,N_6726,N_8903);
and U13011 (N_13011,N_6797,N_7832);
or U13012 (N_13012,N_8451,N_5298);
or U13013 (N_13013,N_6660,N_9993);
xnor U13014 (N_13014,N_8054,N_9646);
nor U13015 (N_13015,N_9496,N_8888);
or U13016 (N_13016,N_7888,N_6042);
xor U13017 (N_13017,N_9596,N_7028);
xor U13018 (N_13018,N_6720,N_6555);
nor U13019 (N_13019,N_7192,N_9631);
nor U13020 (N_13020,N_6700,N_6389);
and U13021 (N_13021,N_5117,N_6318);
xor U13022 (N_13022,N_9466,N_6171);
or U13023 (N_13023,N_5080,N_6352);
nand U13024 (N_13024,N_8742,N_6461);
nand U13025 (N_13025,N_5152,N_6805);
or U13026 (N_13026,N_9612,N_7374);
or U13027 (N_13027,N_8545,N_6189);
xor U13028 (N_13028,N_9590,N_6625);
xor U13029 (N_13029,N_7956,N_9903);
and U13030 (N_13030,N_9774,N_7110);
xnor U13031 (N_13031,N_9235,N_5275);
nor U13032 (N_13032,N_9649,N_6901);
nand U13033 (N_13033,N_9213,N_5857);
nand U13034 (N_13034,N_9796,N_9610);
xnor U13035 (N_13035,N_6174,N_5711);
nand U13036 (N_13036,N_5360,N_5384);
nor U13037 (N_13037,N_6402,N_9817);
and U13038 (N_13038,N_5841,N_8762);
nor U13039 (N_13039,N_7133,N_6828);
nand U13040 (N_13040,N_8332,N_6722);
nor U13041 (N_13041,N_5161,N_8720);
xnor U13042 (N_13042,N_8612,N_7645);
or U13043 (N_13043,N_6994,N_7573);
nand U13044 (N_13044,N_9944,N_8416);
and U13045 (N_13045,N_8978,N_9554);
and U13046 (N_13046,N_9362,N_6269);
nor U13047 (N_13047,N_9140,N_9163);
or U13048 (N_13048,N_7211,N_5313);
and U13049 (N_13049,N_6662,N_5116);
xnor U13050 (N_13050,N_6712,N_6562);
or U13051 (N_13051,N_5207,N_6677);
or U13052 (N_13052,N_7596,N_7579);
and U13053 (N_13053,N_7903,N_9502);
and U13054 (N_13054,N_8627,N_5672);
nor U13055 (N_13055,N_7059,N_8694);
xnor U13056 (N_13056,N_6590,N_6905);
xnor U13057 (N_13057,N_9921,N_5772);
nand U13058 (N_13058,N_9129,N_6772);
and U13059 (N_13059,N_9609,N_8384);
and U13060 (N_13060,N_5215,N_7385);
nand U13061 (N_13061,N_8433,N_9754);
or U13062 (N_13062,N_7271,N_6563);
or U13063 (N_13063,N_6724,N_6238);
or U13064 (N_13064,N_8713,N_9063);
nor U13065 (N_13065,N_6784,N_9542);
xor U13066 (N_13066,N_6592,N_8138);
xor U13067 (N_13067,N_6356,N_5652);
nor U13068 (N_13068,N_5592,N_5616);
xor U13069 (N_13069,N_9189,N_7916);
and U13070 (N_13070,N_7157,N_5345);
nor U13071 (N_13071,N_9571,N_5711);
xnor U13072 (N_13072,N_6557,N_5535);
or U13073 (N_13073,N_8836,N_7711);
xor U13074 (N_13074,N_5670,N_9314);
and U13075 (N_13075,N_6046,N_9256);
nor U13076 (N_13076,N_5386,N_6024);
nand U13077 (N_13077,N_8119,N_7132);
or U13078 (N_13078,N_8308,N_7276);
and U13079 (N_13079,N_6178,N_5490);
xnor U13080 (N_13080,N_8832,N_7474);
and U13081 (N_13081,N_8461,N_8124);
xor U13082 (N_13082,N_5436,N_8751);
nor U13083 (N_13083,N_8644,N_7222);
nor U13084 (N_13084,N_9083,N_7916);
nor U13085 (N_13085,N_7551,N_5116);
nand U13086 (N_13086,N_5579,N_7801);
and U13087 (N_13087,N_8856,N_7946);
nand U13088 (N_13088,N_6882,N_8633);
xnor U13089 (N_13089,N_8356,N_5349);
xnor U13090 (N_13090,N_7150,N_7660);
nand U13091 (N_13091,N_9540,N_7702);
nor U13092 (N_13092,N_5433,N_6076);
and U13093 (N_13093,N_9275,N_7433);
nand U13094 (N_13094,N_6025,N_9962);
xor U13095 (N_13095,N_9704,N_8202);
nor U13096 (N_13096,N_7124,N_7231);
nand U13097 (N_13097,N_5225,N_8408);
and U13098 (N_13098,N_6128,N_6466);
and U13099 (N_13099,N_8044,N_7035);
xor U13100 (N_13100,N_8740,N_5170);
nand U13101 (N_13101,N_7374,N_9548);
and U13102 (N_13102,N_6266,N_8320);
xnor U13103 (N_13103,N_9566,N_5196);
xor U13104 (N_13104,N_8275,N_6504);
and U13105 (N_13105,N_6185,N_5915);
and U13106 (N_13106,N_6337,N_9894);
or U13107 (N_13107,N_5182,N_8458);
and U13108 (N_13108,N_8052,N_6169);
nor U13109 (N_13109,N_7340,N_7720);
nor U13110 (N_13110,N_7259,N_9279);
nand U13111 (N_13111,N_8191,N_9084);
nor U13112 (N_13112,N_7599,N_7160);
or U13113 (N_13113,N_7053,N_7963);
nand U13114 (N_13114,N_9950,N_7185);
and U13115 (N_13115,N_8450,N_6840);
or U13116 (N_13116,N_7995,N_6970);
and U13117 (N_13117,N_7591,N_6648);
nor U13118 (N_13118,N_9861,N_6298);
and U13119 (N_13119,N_6849,N_8161);
nand U13120 (N_13120,N_9747,N_5646);
or U13121 (N_13121,N_5765,N_8635);
xor U13122 (N_13122,N_7210,N_6749);
and U13123 (N_13123,N_8915,N_6887);
or U13124 (N_13124,N_7961,N_7239);
nor U13125 (N_13125,N_9435,N_6645);
nor U13126 (N_13126,N_7330,N_7902);
nor U13127 (N_13127,N_9851,N_6031);
nand U13128 (N_13128,N_5957,N_5288);
nor U13129 (N_13129,N_8073,N_8347);
nor U13130 (N_13130,N_9981,N_9427);
or U13131 (N_13131,N_8275,N_6703);
xor U13132 (N_13132,N_7925,N_9914);
nor U13133 (N_13133,N_5212,N_9426);
nor U13134 (N_13134,N_6545,N_8186);
nor U13135 (N_13135,N_5936,N_5589);
xor U13136 (N_13136,N_5033,N_8032);
or U13137 (N_13137,N_9573,N_5861);
nor U13138 (N_13138,N_7862,N_7327);
nand U13139 (N_13139,N_9320,N_9854);
or U13140 (N_13140,N_9267,N_7402);
xnor U13141 (N_13141,N_6761,N_7964);
xnor U13142 (N_13142,N_5332,N_5880);
or U13143 (N_13143,N_6060,N_9223);
or U13144 (N_13144,N_5594,N_8537);
and U13145 (N_13145,N_6570,N_7573);
or U13146 (N_13146,N_9625,N_9992);
nand U13147 (N_13147,N_5878,N_5420);
or U13148 (N_13148,N_8122,N_9960);
nand U13149 (N_13149,N_5071,N_8924);
nor U13150 (N_13150,N_8281,N_5384);
nor U13151 (N_13151,N_6109,N_8137);
and U13152 (N_13152,N_6288,N_6076);
and U13153 (N_13153,N_9956,N_7451);
and U13154 (N_13154,N_6599,N_5029);
xor U13155 (N_13155,N_8314,N_5690);
or U13156 (N_13156,N_8882,N_8219);
xor U13157 (N_13157,N_9244,N_7892);
and U13158 (N_13158,N_7153,N_5830);
nand U13159 (N_13159,N_8931,N_6693);
nand U13160 (N_13160,N_5625,N_8185);
and U13161 (N_13161,N_5816,N_8429);
nand U13162 (N_13162,N_8212,N_7256);
nand U13163 (N_13163,N_9897,N_6641);
xor U13164 (N_13164,N_7094,N_9918);
nor U13165 (N_13165,N_7981,N_9350);
xnor U13166 (N_13166,N_6552,N_5314);
and U13167 (N_13167,N_7760,N_7047);
or U13168 (N_13168,N_9512,N_7021);
nand U13169 (N_13169,N_9267,N_6554);
nor U13170 (N_13170,N_8705,N_7079);
nand U13171 (N_13171,N_9743,N_6602);
or U13172 (N_13172,N_8620,N_5573);
or U13173 (N_13173,N_9046,N_6504);
or U13174 (N_13174,N_7371,N_8163);
or U13175 (N_13175,N_8036,N_9052);
nand U13176 (N_13176,N_8523,N_7094);
xnor U13177 (N_13177,N_8105,N_7200);
nand U13178 (N_13178,N_9332,N_7026);
and U13179 (N_13179,N_6130,N_8571);
and U13180 (N_13180,N_7533,N_9439);
and U13181 (N_13181,N_8582,N_7195);
nor U13182 (N_13182,N_7532,N_5954);
and U13183 (N_13183,N_9563,N_7702);
or U13184 (N_13184,N_8165,N_5275);
nand U13185 (N_13185,N_5445,N_5263);
nand U13186 (N_13186,N_6495,N_9006);
nand U13187 (N_13187,N_5475,N_6819);
xnor U13188 (N_13188,N_7146,N_5733);
nand U13189 (N_13189,N_7202,N_8727);
and U13190 (N_13190,N_5575,N_9656);
and U13191 (N_13191,N_9645,N_8360);
or U13192 (N_13192,N_8361,N_6805);
and U13193 (N_13193,N_7781,N_7659);
nand U13194 (N_13194,N_7042,N_8645);
xor U13195 (N_13195,N_9829,N_8402);
and U13196 (N_13196,N_8801,N_9806);
and U13197 (N_13197,N_6763,N_9572);
and U13198 (N_13198,N_5054,N_7693);
and U13199 (N_13199,N_5751,N_7561);
and U13200 (N_13200,N_9879,N_6180);
nor U13201 (N_13201,N_8037,N_7784);
or U13202 (N_13202,N_6564,N_7027);
xor U13203 (N_13203,N_9703,N_8264);
or U13204 (N_13204,N_7895,N_9590);
nand U13205 (N_13205,N_9633,N_9223);
or U13206 (N_13206,N_7882,N_6249);
nor U13207 (N_13207,N_8859,N_7982);
or U13208 (N_13208,N_5584,N_8217);
or U13209 (N_13209,N_5796,N_5151);
and U13210 (N_13210,N_5885,N_8919);
xnor U13211 (N_13211,N_5318,N_5703);
and U13212 (N_13212,N_7715,N_8106);
nand U13213 (N_13213,N_8214,N_8560);
or U13214 (N_13214,N_9653,N_9091);
or U13215 (N_13215,N_5765,N_5898);
or U13216 (N_13216,N_7564,N_7396);
nor U13217 (N_13217,N_5999,N_8916);
nand U13218 (N_13218,N_7910,N_7621);
xor U13219 (N_13219,N_7277,N_9589);
or U13220 (N_13220,N_6839,N_6584);
nor U13221 (N_13221,N_5751,N_8230);
nand U13222 (N_13222,N_6665,N_9704);
nand U13223 (N_13223,N_9587,N_7842);
and U13224 (N_13224,N_5884,N_7411);
nor U13225 (N_13225,N_6844,N_5058);
and U13226 (N_13226,N_5836,N_6594);
nor U13227 (N_13227,N_5209,N_8431);
and U13228 (N_13228,N_5666,N_5557);
or U13229 (N_13229,N_5561,N_7161);
or U13230 (N_13230,N_7672,N_6634);
nor U13231 (N_13231,N_6787,N_5018);
xor U13232 (N_13232,N_9619,N_5773);
and U13233 (N_13233,N_7878,N_9996);
and U13234 (N_13234,N_8882,N_9971);
or U13235 (N_13235,N_8758,N_7755);
nor U13236 (N_13236,N_9245,N_9874);
and U13237 (N_13237,N_6805,N_7888);
nand U13238 (N_13238,N_5657,N_9456);
or U13239 (N_13239,N_9563,N_9265);
nor U13240 (N_13240,N_7243,N_8663);
nor U13241 (N_13241,N_5657,N_6360);
and U13242 (N_13242,N_9811,N_9496);
xnor U13243 (N_13243,N_6971,N_8070);
nor U13244 (N_13244,N_8709,N_5998);
nand U13245 (N_13245,N_5941,N_6674);
xnor U13246 (N_13246,N_8861,N_9708);
and U13247 (N_13247,N_7284,N_7212);
nor U13248 (N_13248,N_5011,N_7372);
xor U13249 (N_13249,N_6315,N_5565);
nand U13250 (N_13250,N_6720,N_8734);
xor U13251 (N_13251,N_8323,N_7765);
or U13252 (N_13252,N_8833,N_8135);
xor U13253 (N_13253,N_8377,N_6957);
xnor U13254 (N_13254,N_5590,N_6504);
xnor U13255 (N_13255,N_7038,N_5899);
nor U13256 (N_13256,N_8746,N_9975);
or U13257 (N_13257,N_5038,N_9519);
nor U13258 (N_13258,N_5462,N_8369);
and U13259 (N_13259,N_9722,N_9177);
xnor U13260 (N_13260,N_7256,N_7117);
and U13261 (N_13261,N_7807,N_9065);
and U13262 (N_13262,N_6590,N_5651);
nor U13263 (N_13263,N_5026,N_6591);
nor U13264 (N_13264,N_9481,N_5624);
and U13265 (N_13265,N_8544,N_7216);
or U13266 (N_13266,N_6124,N_5863);
xnor U13267 (N_13267,N_9427,N_8908);
nor U13268 (N_13268,N_8107,N_6581);
nand U13269 (N_13269,N_5603,N_7609);
or U13270 (N_13270,N_7642,N_6924);
nand U13271 (N_13271,N_8446,N_5969);
xor U13272 (N_13272,N_6442,N_6737);
or U13273 (N_13273,N_9951,N_5757);
and U13274 (N_13274,N_7218,N_8207);
nor U13275 (N_13275,N_6467,N_7421);
xor U13276 (N_13276,N_8151,N_9272);
and U13277 (N_13277,N_5383,N_9807);
or U13278 (N_13278,N_8659,N_6637);
nor U13279 (N_13279,N_9600,N_8731);
nand U13280 (N_13280,N_7775,N_9813);
and U13281 (N_13281,N_8355,N_9891);
nor U13282 (N_13282,N_6265,N_9817);
nor U13283 (N_13283,N_7684,N_9411);
xnor U13284 (N_13284,N_5293,N_5894);
nor U13285 (N_13285,N_6693,N_9463);
xnor U13286 (N_13286,N_7233,N_9936);
nand U13287 (N_13287,N_5557,N_9273);
nor U13288 (N_13288,N_6405,N_8609);
nand U13289 (N_13289,N_6208,N_7015);
xnor U13290 (N_13290,N_8486,N_8819);
xnor U13291 (N_13291,N_7242,N_8069);
and U13292 (N_13292,N_6874,N_5578);
and U13293 (N_13293,N_7348,N_5694);
or U13294 (N_13294,N_6424,N_6967);
nand U13295 (N_13295,N_9082,N_8762);
xor U13296 (N_13296,N_5652,N_5943);
nand U13297 (N_13297,N_5395,N_9528);
nand U13298 (N_13298,N_8949,N_5679);
xor U13299 (N_13299,N_5568,N_9948);
or U13300 (N_13300,N_9792,N_6759);
nor U13301 (N_13301,N_6107,N_6883);
nand U13302 (N_13302,N_5599,N_9018);
nor U13303 (N_13303,N_7139,N_6073);
and U13304 (N_13304,N_6863,N_9466);
xnor U13305 (N_13305,N_9108,N_9480);
and U13306 (N_13306,N_7327,N_9607);
nand U13307 (N_13307,N_9726,N_5834);
or U13308 (N_13308,N_9979,N_5339);
nand U13309 (N_13309,N_8987,N_7375);
xor U13310 (N_13310,N_9345,N_5513);
xor U13311 (N_13311,N_6467,N_7973);
and U13312 (N_13312,N_8206,N_6537);
and U13313 (N_13313,N_7745,N_7320);
xor U13314 (N_13314,N_7696,N_6312);
xor U13315 (N_13315,N_6068,N_8482);
and U13316 (N_13316,N_5999,N_7648);
or U13317 (N_13317,N_7354,N_7342);
nand U13318 (N_13318,N_8374,N_5591);
xor U13319 (N_13319,N_6000,N_6664);
nor U13320 (N_13320,N_5259,N_9467);
or U13321 (N_13321,N_5169,N_7456);
xor U13322 (N_13322,N_8406,N_7803);
or U13323 (N_13323,N_6941,N_7810);
and U13324 (N_13324,N_6857,N_7822);
nand U13325 (N_13325,N_5773,N_9231);
xnor U13326 (N_13326,N_6648,N_5742);
nand U13327 (N_13327,N_5970,N_5358);
nand U13328 (N_13328,N_7654,N_6208);
and U13329 (N_13329,N_7227,N_8584);
and U13330 (N_13330,N_8397,N_7417);
xnor U13331 (N_13331,N_8366,N_5082);
nand U13332 (N_13332,N_5712,N_7851);
nand U13333 (N_13333,N_5187,N_8426);
and U13334 (N_13334,N_5082,N_5303);
and U13335 (N_13335,N_8806,N_8642);
and U13336 (N_13336,N_8484,N_8639);
or U13337 (N_13337,N_9569,N_6635);
nor U13338 (N_13338,N_9420,N_5521);
or U13339 (N_13339,N_7629,N_9560);
xnor U13340 (N_13340,N_8440,N_6793);
and U13341 (N_13341,N_9299,N_9978);
xnor U13342 (N_13342,N_7184,N_7917);
and U13343 (N_13343,N_6989,N_9351);
and U13344 (N_13344,N_9951,N_5037);
or U13345 (N_13345,N_9095,N_7785);
xnor U13346 (N_13346,N_8052,N_9982);
xor U13347 (N_13347,N_8958,N_7962);
and U13348 (N_13348,N_8321,N_6636);
or U13349 (N_13349,N_6898,N_6273);
and U13350 (N_13350,N_8472,N_6363);
and U13351 (N_13351,N_7658,N_7550);
xor U13352 (N_13352,N_9242,N_8473);
nor U13353 (N_13353,N_8858,N_5445);
and U13354 (N_13354,N_6506,N_9960);
xnor U13355 (N_13355,N_9220,N_9061);
nor U13356 (N_13356,N_5444,N_7086);
and U13357 (N_13357,N_8074,N_6759);
or U13358 (N_13358,N_8055,N_8184);
nor U13359 (N_13359,N_9896,N_5217);
and U13360 (N_13360,N_9389,N_6509);
nor U13361 (N_13361,N_7553,N_9496);
nor U13362 (N_13362,N_6284,N_8386);
or U13363 (N_13363,N_9472,N_8647);
nand U13364 (N_13364,N_7159,N_5908);
nor U13365 (N_13365,N_9770,N_7429);
xnor U13366 (N_13366,N_7557,N_6996);
nand U13367 (N_13367,N_6869,N_7515);
or U13368 (N_13368,N_7753,N_9764);
nor U13369 (N_13369,N_7738,N_7129);
or U13370 (N_13370,N_6443,N_8080);
and U13371 (N_13371,N_9694,N_8507);
and U13372 (N_13372,N_6132,N_9454);
and U13373 (N_13373,N_5437,N_9863);
nor U13374 (N_13374,N_5033,N_5058);
nand U13375 (N_13375,N_7633,N_9176);
or U13376 (N_13376,N_8385,N_8075);
nand U13377 (N_13377,N_8775,N_5557);
or U13378 (N_13378,N_9341,N_9120);
xor U13379 (N_13379,N_8195,N_8200);
xor U13380 (N_13380,N_7367,N_9730);
nand U13381 (N_13381,N_8821,N_5968);
and U13382 (N_13382,N_7858,N_8772);
nor U13383 (N_13383,N_9293,N_6102);
and U13384 (N_13384,N_6050,N_7216);
xor U13385 (N_13385,N_5344,N_7185);
and U13386 (N_13386,N_8283,N_9217);
and U13387 (N_13387,N_8671,N_5758);
and U13388 (N_13388,N_7532,N_8929);
nor U13389 (N_13389,N_6681,N_6083);
or U13390 (N_13390,N_6556,N_6326);
and U13391 (N_13391,N_9958,N_8892);
xnor U13392 (N_13392,N_8221,N_5631);
or U13393 (N_13393,N_5584,N_6212);
xnor U13394 (N_13394,N_7842,N_8017);
nand U13395 (N_13395,N_7092,N_6549);
nor U13396 (N_13396,N_8422,N_5387);
and U13397 (N_13397,N_9206,N_9995);
xnor U13398 (N_13398,N_6738,N_7757);
or U13399 (N_13399,N_8499,N_8498);
or U13400 (N_13400,N_6490,N_8683);
and U13401 (N_13401,N_5799,N_6563);
or U13402 (N_13402,N_5138,N_5067);
or U13403 (N_13403,N_5956,N_7767);
nand U13404 (N_13404,N_9829,N_8456);
nand U13405 (N_13405,N_7254,N_5193);
nand U13406 (N_13406,N_9351,N_6554);
nor U13407 (N_13407,N_5341,N_8650);
and U13408 (N_13408,N_5863,N_8085);
and U13409 (N_13409,N_5796,N_5008);
or U13410 (N_13410,N_7436,N_7684);
and U13411 (N_13411,N_6122,N_9801);
nand U13412 (N_13412,N_9975,N_6092);
xor U13413 (N_13413,N_5116,N_9369);
nand U13414 (N_13414,N_7030,N_8109);
and U13415 (N_13415,N_8880,N_6855);
xor U13416 (N_13416,N_9165,N_6379);
nand U13417 (N_13417,N_7913,N_7044);
and U13418 (N_13418,N_5307,N_5690);
xnor U13419 (N_13419,N_5695,N_8887);
nor U13420 (N_13420,N_8853,N_8129);
nor U13421 (N_13421,N_6087,N_7097);
and U13422 (N_13422,N_5981,N_6345);
nand U13423 (N_13423,N_8637,N_8111);
xor U13424 (N_13424,N_7544,N_8206);
nor U13425 (N_13425,N_5757,N_6291);
nand U13426 (N_13426,N_9196,N_9151);
and U13427 (N_13427,N_7283,N_8063);
nor U13428 (N_13428,N_7150,N_8272);
nand U13429 (N_13429,N_6242,N_5276);
or U13430 (N_13430,N_7951,N_7524);
nor U13431 (N_13431,N_7684,N_7946);
and U13432 (N_13432,N_6617,N_5119);
nor U13433 (N_13433,N_8760,N_8019);
or U13434 (N_13434,N_5016,N_8263);
and U13435 (N_13435,N_5262,N_5479);
xor U13436 (N_13436,N_9189,N_5908);
xnor U13437 (N_13437,N_9368,N_5148);
nor U13438 (N_13438,N_8321,N_8474);
or U13439 (N_13439,N_5802,N_6787);
nand U13440 (N_13440,N_9173,N_8092);
xor U13441 (N_13441,N_9376,N_6283);
nor U13442 (N_13442,N_9704,N_5847);
xnor U13443 (N_13443,N_7942,N_5189);
xor U13444 (N_13444,N_8157,N_6796);
xor U13445 (N_13445,N_8806,N_8965);
and U13446 (N_13446,N_8666,N_7049);
xor U13447 (N_13447,N_5222,N_6068);
nand U13448 (N_13448,N_9008,N_9878);
or U13449 (N_13449,N_7817,N_8457);
nand U13450 (N_13450,N_9866,N_8550);
and U13451 (N_13451,N_7361,N_5741);
nand U13452 (N_13452,N_9976,N_5349);
or U13453 (N_13453,N_5576,N_8356);
and U13454 (N_13454,N_8701,N_9967);
xor U13455 (N_13455,N_9486,N_9957);
xnor U13456 (N_13456,N_6381,N_5604);
nor U13457 (N_13457,N_7156,N_7554);
nor U13458 (N_13458,N_5922,N_7686);
nor U13459 (N_13459,N_5490,N_6221);
and U13460 (N_13460,N_6633,N_9096);
nor U13461 (N_13461,N_6050,N_6072);
or U13462 (N_13462,N_6882,N_6180);
nor U13463 (N_13463,N_6638,N_9721);
and U13464 (N_13464,N_8016,N_8941);
nand U13465 (N_13465,N_7287,N_5701);
or U13466 (N_13466,N_9691,N_7380);
xnor U13467 (N_13467,N_9016,N_8027);
or U13468 (N_13468,N_5190,N_5044);
xor U13469 (N_13469,N_5306,N_8423);
nand U13470 (N_13470,N_8982,N_8133);
xnor U13471 (N_13471,N_7453,N_9404);
xnor U13472 (N_13472,N_5478,N_6725);
xnor U13473 (N_13473,N_7041,N_7550);
nand U13474 (N_13474,N_8434,N_8200);
nor U13475 (N_13475,N_7998,N_8847);
xor U13476 (N_13476,N_6369,N_9751);
or U13477 (N_13477,N_6467,N_5311);
and U13478 (N_13478,N_6823,N_9171);
or U13479 (N_13479,N_6510,N_7152);
and U13480 (N_13480,N_8373,N_9582);
and U13481 (N_13481,N_9325,N_8463);
xor U13482 (N_13482,N_9322,N_9684);
or U13483 (N_13483,N_8808,N_8634);
and U13484 (N_13484,N_7265,N_6298);
nand U13485 (N_13485,N_6903,N_6484);
or U13486 (N_13486,N_8924,N_7114);
nand U13487 (N_13487,N_5906,N_5897);
or U13488 (N_13488,N_7245,N_8529);
nor U13489 (N_13489,N_6914,N_9136);
nor U13490 (N_13490,N_6654,N_7063);
or U13491 (N_13491,N_7021,N_5818);
and U13492 (N_13492,N_7815,N_8486);
nand U13493 (N_13493,N_6805,N_5565);
and U13494 (N_13494,N_9289,N_6606);
nor U13495 (N_13495,N_8023,N_5607);
nor U13496 (N_13496,N_9979,N_6394);
and U13497 (N_13497,N_6018,N_7021);
or U13498 (N_13498,N_8266,N_5027);
xor U13499 (N_13499,N_8105,N_6910);
nand U13500 (N_13500,N_7951,N_5193);
and U13501 (N_13501,N_8518,N_5972);
nor U13502 (N_13502,N_8928,N_5466);
nor U13503 (N_13503,N_9262,N_7429);
nand U13504 (N_13504,N_6783,N_5777);
or U13505 (N_13505,N_5386,N_5252);
nor U13506 (N_13506,N_8489,N_9608);
xnor U13507 (N_13507,N_5014,N_9254);
nand U13508 (N_13508,N_5722,N_6772);
and U13509 (N_13509,N_8743,N_7912);
nand U13510 (N_13510,N_9590,N_8289);
xnor U13511 (N_13511,N_6694,N_9834);
nor U13512 (N_13512,N_9754,N_8147);
and U13513 (N_13513,N_7994,N_6438);
nor U13514 (N_13514,N_6296,N_9303);
xor U13515 (N_13515,N_9355,N_6081);
nor U13516 (N_13516,N_8874,N_8882);
nand U13517 (N_13517,N_6549,N_8681);
nand U13518 (N_13518,N_5265,N_5916);
or U13519 (N_13519,N_5468,N_5825);
and U13520 (N_13520,N_9806,N_6710);
and U13521 (N_13521,N_7085,N_9154);
or U13522 (N_13522,N_7721,N_5373);
and U13523 (N_13523,N_8813,N_6497);
xor U13524 (N_13524,N_5776,N_7763);
or U13525 (N_13525,N_5344,N_8091);
xor U13526 (N_13526,N_8094,N_5556);
nor U13527 (N_13527,N_7221,N_5773);
and U13528 (N_13528,N_7273,N_8455);
nand U13529 (N_13529,N_7201,N_6754);
or U13530 (N_13530,N_7232,N_5409);
nor U13531 (N_13531,N_7005,N_5707);
nand U13532 (N_13532,N_9964,N_9916);
nand U13533 (N_13533,N_7560,N_5430);
and U13534 (N_13534,N_5196,N_9762);
nor U13535 (N_13535,N_8563,N_5126);
or U13536 (N_13536,N_6628,N_8540);
nand U13537 (N_13537,N_7059,N_8156);
and U13538 (N_13538,N_5729,N_5960);
nor U13539 (N_13539,N_5792,N_5834);
nand U13540 (N_13540,N_5813,N_9095);
and U13541 (N_13541,N_9858,N_6205);
nand U13542 (N_13542,N_5060,N_6970);
and U13543 (N_13543,N_8936,N_6049);
or U13544 (N_13544,N_9387,N_5812);
and U13545 (N_13545,N_5235,N_5671);
nand U13546 (N_13546,N_9174,N_9805);
xor U13547 (N_13547,N_5039,N_7857);
or U13548 (N_13548,N_7997,N_9163);
nand U13549 (N_13549,N_9440,N_7284);
and U13550 (N_13550,N_9520,N_6734);
and U13551 (N_13551,N_9816,N_9701);
nand U13552 (N_13552,N_6063,N_5511);
nor U13553 (N_13553,N_7439,N_8253);
or U13554 (N_13554,N_6042,N_8153);
nor U13555 (N_13555,N_5949,N_6021);
or U13556 (N_13556,N_6845,N_8769);
nand U13557 (N_13557,N_6944,N_7185);
or U13558 (N_13558,N_6219,N_6076);
nand U13559 (N_13559,N_5056,N_9829);
nor U13560 (N_13560,N_9889,N_6625);
or U13561 (N_13561,N_9828,N_9656);
nor U13562 (N_13562,N_8792,N_8948);
and U13563 (N_13563,N_5437,N_7046);
nand U13564 (N_13564,N_5186,N_5351);
nand U13565 (N_13565,N_9102,N_6066);
nor U13566 (N_13566,N_9654,N_7556);
xnor U13567 (N_13567,N_9644,N_7241);
and U13568 (N_13568,N_9431,N_6378);
xnor U13569 (N_13569,N_6039,N_9465);
or U13570 (N_13570,N_5233,N_5662);
or U13571 (N_13571,N_7075,N_9418);
or U13572 (N_13572,N_7130,N_9847);
xnor U13573 (N_13573,N_6076,N_6750);
nand U13574 (N_13574,N_8657,N_5221);
nand U13575 (N_13575,N_6636,N_5743);
nor U13576 (N_13576,N_5868,N_8008);
or U13577 (N_13577,N_6346,N_6039);
nor U13578 (N_13578,N_5362,N_9019);
nand U13579 (N_13579,N_8632,N_7674);
or U13580 (N_13580,N_6731,N_6696);
nand U13581 (N_13581,N_6703,N_7202);
xnor U13582 (N_13582,N_9848,N_9394);
xnor U13583 (N_13583,N_7249,N_7153);
nand U13584 (N_13584,N_6194,N_8351);
nand U13585 (N_13585,N_6755,N_8045);
and U13586 (N_13586,N_6383,N_5152);
nor U13587 (N_13587,N_5900,N_7361);
xor U13588 (N_13588,N_7395,N_5349);
nor U13589 (N_13589,N_6464,N_8532);
nand U13590 (N_13590,N_8750,N_5582);
and U13591 (N_13591,N_7551,N_7555);
or U13592 (N_13592,N_9119,N_8485);
and U13593 (N_13593,N_5455,N_6912);
nand U13594 (N_13594,N_6197,N_5422);
nand U13595 (N_13595,N_9244,N_6483);
or U13596 (N_13596,N_9678,N_5894);
or U13597 (N_13597,N_8958,N_5152);
or U13598 (N_13598,N_8823,N_6162);
nand U13599 (N_13599,N_8539,N_6672);
or U13600 (N_13600,N_8461,N_9494);
nor U13601 (N_13601,N_6787,N_8530);
nor U13602 (N_13602,N_9018,N_9661);
nand U13603 (N_13603,N_9730,N_7518);
nor U13604 (N_13604,N_8139,N_5094);
or U13605 (N_13605,N_8450,N_5679);
nand U13606 (N_13606,N_6258,N_6266);
nand U13607 (N_13607,N_6946,N_9217);
or U13608 (N_13608,N_5730,N_8185);
nor U13609 (N_13609,N_9863,N_5890);
and U13610 (N_13610,N_9477,N_6481);
or U13611 (N_13611,N_5872,N_8635);
or U13612 (N_13612,N_6854,N_7127);
xor U13613 (N_13613,N_6117,N_7300);
xnor U13614 (N_13614,N_9531,N_6218);
and U13615 (N_13615,N_9787,N_6218);
or U13616 (N_13616,N_9426,N_5093);
nor U13617 (N_13617,N_9430,N_5707);
xor U13618 (N_13618,N_6971,N_9091);
nor U13619 (N_13619,N_5036,N_8542);
nor U13620 (N_13620,N_9485,N_5534);
or U13621 (N_13621,N_7550,N_9095);
xnor U13622 (N_13622,N_9750,N_6053);
xnor U13623 (N_13623,N_8825,N_9156);
or U13624 (N_13624,N_9074,N_5392);
xor U13625 (N_13625,N_9891,N_8765);
xnor U13626 (N_13626,N_8837,N_7177);
nor U13627 (N_13627,N_7192,N_5546);
xnor U13628 (N_13628,N_7406,N_6862);
and U13629 (N_13629,N_6520,N_5572);
nand U13630 (N_13630,N_9864,N_6477);
nand U13631 (N_13631,N_7743,N_9663);
xor U13632 (N_13632,N_5141,N_6368);
or U13633 (N_13633,N_7830,N_5373);
and U13634 (N_13634,N_9543,N_7326);
and U13635 (N_13635,N_8909,N_5042);
xnor U13636 (N_13636,N_9949,N_9144);
or U13637 (N_13637,N_5748,N_8422);
nor U13638 (N_13638,N_9921,N_8819);
nor U13639 (N_13639,N_9820,N_5223);
nand U13640 (N_13640,N_8698,N_6156);
and U13641 (N_13641,N_9819,N_8338);
or U13642 (N_13642,N_8399,N_5639);
nand U13643 (N_13643,N_6701,N_8839);
nand U13644 (N_13644,N_9479,N_7554);
nor U13645 (N_13645,N_6872,N_7953);
xnor U13646 (N_13646,N_6367,N_6523);
nor U13647 (N_13647,N_5781,N_6759);
and U13648 (N_13648,N_7142,N_9015);
xor U13649 (N_13649,N_6911,N_7539);
and U13650 (N_13650,N_6675,N_8860);
and U13651 (N_13651,N_8619,N_5262);
nor U13652 (N_13652,N_9814,N_7990);
nor U13653 (N_13653,N_8776,N_6377);
xor U13654 (N_13654,N_9999,N_7314);
nor U13655 (N_13655,N_7409,N_9216);
and U13656 (N_13656,N_8385,N_8733);
and U13657 (N_13657,N_8901,N_7040);
nand U13658 (N_13658,N_7021,N_5594);
nand U13659 (N_13659,N_8342,N_5464);
nor U13660 (N_13660,N_8005,N_6073);
xnor U13661 (N_13661,N_7643,N_9137);
xor U13662 (N_13662,N_7755,N_8763);
and U13663 (N_13663,N_5476,N_8949);
nor U13664 (N_13664,N_8691,N_9925);
xnor U13665 (N_13665,N_8278,N_9927);
nor U13666 (N_13666,N_9914,N_9143);
xor U13667 (N_13667,N_9527,N_6174);
and U13668 (N_13668,N_6757,N_8512);
xnor U13669 (N_13669,N_9537,N_5010);
nand U13670 (N_13670,N_7575,N_8228);
and U13671 (N_13671,N_8920,N_8339);
nand U13672 (N_13672,N_9157,N_9768);
nor U13673 (N_13673,N_9694,N_6515);
nand U13674 (N_13674,N_7809,N_9860);
nor U13675 (N_13675,N_9303,N_7104);
or U13676 (N_13676,N_7622,N_5001);
and U13677 (N_13677,N_6384,N_9924);
or U13678 (N_13678,N_8159,N_6825);
nand U13679 (N_13679,N_7798,N_9389);
xnor U13680 (N_13680,N_8696,N_5955);
nand U13681 (N_13681,N_6969,N_7149);
and U13682 (N_13682,N_7791,N_9422);
and U13683 (N_13683,N_6210,N_6123);
nor U13684 (N_13684,N_7586,N_5000);
and U13685 (N_13685,N_7505,N_7542);
nand U13686 (N_13686,N_5615,N_6487);
nor U13687 (N_13687,N_8555,N_5734);
nand U13688 (N_13688,N_6081,N_7329);
and U13689 (N_13689,N_6961,N_5929);
or U13690 (N_13690,N_8583,N_5397);
nand U13691 (N_13691,N_8624,N_7299);
nand U13692 (N_13692,N_7547,N_5809);
xor U13693 (N_13693,N_8050,N_8121);
or U13694 (N_13694,N_7359,N_5032);
or U13695 (N_13695,N_5904,N_6205);
nand U13696 (N_13696,N_7999,N_8706);
and U13697 (N_13697,N_6655,N_5044);
nand U13698 (N_13698,N_8436,N_6619);
or U13699 (N_13699,N_5626,N_8765);
xnor U13700 (N_13700,N_9473,N_8703);
nand U13701 (N_13701,N_8075,N_9356);
and U13702 (N_13702,N_9064,N_7690);
nor U13703 (N_13703,N_5357,N_9708);
or U13704 (N_13704,N_7777,N_6189);
or U13705 (N_13705,N_5309,N_6407);
nor U13706 (N_13706,N_5751,N_8496);
or U13707 (N_13707,N_7927,N_8786);
xor U13708 (N_13708,N_7733,N_5216);
xor U13709 (N_13709,N_6433,N_5995);
and U13710 (N_13710,N_8938,N_8653);
xnor U13711 (N_13711,N_8797,N_5244);
or U13712 (N_13712,N_9502,N_5977);
nor U13713 (N_13713,N_6833,N_6868);
and U13714 (N_13714,N_7556,N_9606);
nand U13715 (N_13715,N_5844,N_7492);
xnor U13716 (N_13716,N_7670,N_7661);
nand U13717 (N_13717,N_7046,N_5404);
nand U13718 (N_13718,N_7771,N_8528);
and U13719 (N_13719,N_9694,N_8611);
and U13720 (N_13720,N_8264,N_5286);
xnor U13721 (N_13721,N_5084,N_8003);
and U13722 (N_13722,N_8958,N_9616);
nand U13723 (N_13723,N_9538,N_7236);
nand U13724 (N_13724,N_8903,N_8466);
nor U13725 (N_13725,N_5790,N_7799);
and U13726 (N_13726,N_7136,N_7963);
or U13727 (N_13727,N_9000,N_8980);
nor U13728 (N_13728,N_8291,N_9135);
and U13729 (N_13729,N_8641,N_5874);
nor U13730 (N_13730,N_8778,N_5110);
or U13731 (N_13731,N_8444,N_6065);
xor U13732 (N_13732,N_5739,N_7073);
and U13733 (N_13733,N_8889,N_9159);
or U13734 (N_13734,N_8871,N_9220);
and U13735 (N_13735,N_8913,N_6042);
nand U13736 (N_13736,N_6004,N_9243);
nor U13737 (N_13737,N_5245,N_9708);
nand U13738 (N_13738,N_5278,N_7579);
nand U13739 (N_13739,N_6425,N_9609);
and U13740 (N_13740,N_9017,N_5567);
nor U13741 (N_13741,N_5907,N_5529);
xnor U13742 (N_13742,N_8541,N_8632);
and U13743 (N_13743,N_7676,N_7179);
xor U13744 (N_13744,N_7275,N_6330);
or U13745 (N_13745,N_9347,N_7749);
nor U13746 (N_13746,N_5516,N_6503);
nand U13747 (N_13747,N_9702,N_8711);
xnor U13748 (N_13748,N_7697,N_9297);
and U13749 (N_13749,N_8831,N_5588);
nor U13750 (N_13750,N_6840,N_9710);
xnor U13751 (N_13751,N_6346,N_5999);
or U13752 (N_13752,N_8226,N_5783);
nor U13753 (N_13753,N_5228,N_8140);
and U13754 (N_13754,N_7575,N_8209);
or U13755 (N_13755,N_5261,N_5320);
or U13756 (N_13756,N_7372,N_9051);
and U13757 (N_13757,N_5413,N_8867);
xor U13758 (N_13758,N_6191,N_8882);
nand U13759 (N_13759,N_8408,N_9940);
nor U13760 (N_13760,N_5934,N_9043);
nand U13761 (N_13761,N_8788,N_8524);
nand U13762 (N_13762,N_9113,N_6904);
nand U13763 (N_13763,N_6773,N_8387);
xor U13764 (N_13764,N_7492,N_8956);
nand U13765 (N_13765,N_9488,N_5097);
and U13766 (N_13766,N_8733,N_8363);
and U13767 (N_13767,N_9979,N_5311);
and U13768 (N_13768,N_8472,N_8025);
nor U13769 (N_13769,N_8983,N_8984);
nand U13770 (N_13770,N_7279,N_6229);
nor U13771 (N_13771,N_7232,N_5564);
or U13772 (N_13772,N_5773,N_7415);
nor U13773 (N_13773,N_5786,N_7764);
xor U13774 (N_13774,N_7733,N_8673);
nand U13775 (N_13775,N_8284,N_7813);
and U13776 (N_13776,N_6836,N_6079);
xor U13777 (N_13777,N_7980,N_5251);
xor U13778 (N_13778,N_6400,N_7766);
xnor U13779 (N_13779,N_7361,N_9207);
or U13780 (N_13780,N_8700,N_6725);
nor U13781 (N_13781,N_8137,N_7446);
nor U13782 (N_13782,N_6654,N_7140);
nand U13783 (N_13783,N_9546,N_8609);
nor U13784 (N_13784,N_8889,N_8508);
nand U13785 (N_13785,N_6436,N_6807);
or U13786 (N_13786,N_8553,N_8088);
and U13787 (N_13787,N_6639,N_8826);
nand U13788 (N_13788,N_8003,N_9295);
nor U13789 (N_13789,N_8221,N_8683);
xor U13790 (N_13790,N_9405,N_6646);
nand U13791 (N_13791,N_5899,N_5353);
xnor U13792 (N_13792,N_6261,N_5101);
nor U13793 (N_13793,N_7001,N_5131);
xor U13794 (N_13794,N_5518,N_6645);
xor U13795 (N_13795,N_9845,N_5450);
or U13796 (N_13796,N_8541,N_7146);
and U13797 (N_13797,N_8766,N_5193);
nand U13798 (N_13798,N_6751,N_9693);
or U13799 (N_13799,N_8904,N_9347);
and U13800 (N_13800,N_5714,N_9776);
nand U13801 (N_13801,N_9814,N_7886);
or U13802 (N_13802,N_8781,N_5155);
or U13803 (N_13803,N_8809,N_5936);
nand U13804 (N_13804,N_7618,N_8524);
nand U13805 (N_13805,N_9459,N_7157);
nor U13806 (N_13806,N_7189,N_8465);
nand U13807 (N_13807,N_6514,N_5330);
nor U13808 (N_13808,N_6165,N_6295);
nand U13809 (N_13809,N_5411,N_8944);
and U13810 (N_13810,N_9205,N_6301);
nand U13811 (N_13811,N_9850,N_8952);
nand U13812 (N_13812,N_9059,N_5593);
xor U13813 (N_13813,N_7465,N_6629);
or U13814 (N_13814,N_9279,N_8364);
or U13815 (N_13815,N_7319,N_5675);
or U13816 (N_13816,N_5175,N_9300);
nor U13817 (N_13817,N_7476,N_7767);
nor U13818 (N_13818,N_6839,N_5856);
or U13819 (N_13819,N_9940,N_7110);
and U13820 (N_13820,N_8077,N_5001);
nand U13821 (N_13821,N_6472,N_5928);
and U13822 (N_13822,N_8816,N_8164);
xor U13823 (N_13823,N_9314,N_9390);
and U13824 (N_13824,N_8457,N_7837);
xnor U13825 (N_13825,N_9250,N_6323);
xnor U13826 (N_13826,N_7682,N_8509);
xnor U13827 (N_13827,N_9618,N_7667);
nor U13828 (N_13828,N_8633,N_6786);
xor U13829 (N_13829,N_5341,N_8803);
xnor U13830 (N_13830,N_8634,N_7183);
nor U13831 (N_13831,N_9807,N_6367);
and U13832 (N_13832,N_9345,N_8057);
xor U13833 (N_13833,N_5481,N_7323);
xor U13834 (N_13834,N_8096,N_5686);
nand U13835 (N_13835,N_5226,N_8163);
nor U13836 (N_13836,N_9970,N_5673);
nand U13837 (N_13837,N_9472,N_6502);
or U13838 (N_13838,N_6131,N_6991);
xor U13839 (N_13839,N_8793,N_9361);
xor U13840 (N_13840,N_5520,N_7187);
or U13841 (N_13841,N_7771,N_9133);
and U13842 (N_13842,N_5214,N_6062);
or U13843 (N_13843,N_7821,N_8401);
or U13844 (N_13844,N_6923,N_6329);
nor U13845 (N_13845,N_5405,N_8626);
nand U13846 (N_13846,N_7020,N_5577);
or U13847 (N_13847,N_6986,N_9930);
and U13848 (N_13848,N_8941,N_5743);
and U13849 (N_13849,N_8669,N_5323);
xor U13850 (N_13850,N_7187,N_5322);
nand U13851 (N_13851,N_8661,N_5845);
or U13852 (N_13852,N_9686,N_5770);
nor U13853 (N_13853,N_7125,N_6651);
and U13854 (N_13854,N_9748,N_5239);
nor U13855 (N_13855,N_8886,N_8188);
and U13856 (N_13856,N_8960,N_6598);
nor U13857 (N_13857,N_7705,N_9380);
nand U13858 (N_13858,N_6128,N_5464);
nand U13859 (N_13859,N_7508,N_6690);
xnor U13860 (N_13860,N_9385,N_8991);
or U13861 (N_13861,N_5314,N_8039);
and U13862 (N_13862,N_5377,N_5018);
nand U13863 (N_13863,N_9170,N_6426);
or U13864 (N_13864,N_8178,N_5241);
and U13865 (N_13865,N_8919,N_8154);
nand U13866 (N_13866,N_6123,N_5290);
nand U13867 (N_13867,N_6025,N_9261);
nor U13868 (N_13868,N_6691,N_8404);
xor U13869 (N_13869,N_6915,N_9408);
and U13870 (N_13870,N_7470,N_5848);
and U13871 (N_13871,N_8472,N_6581);
or U13872 (N_13872,N_9908,N_9458);
nand U13873 (N_13873,N_9798,N_7046);
xor U13874 (N_13874,N_7842,N_7020);
and U13875 (N_13875,N_8627,N_7378);
nand U13876 (N_13876,N_8245,N_5663);
nand U13877 (N_13877,N_5977,N_6643);
or U13878 (N_13878,N_6037,N_8191);
and U13879 (N_13879,N_7526,N_8021);
xnor U13880 (N_13880,N_9881,N_7785);
or U13881 (N_13881,N_8249,N_7501);
nand U13882 (N_13882,N_6840,N_6769);
nand U13883 (N_13883,N_5909,N_6415);
nor U13884 (N_13884,N_7497,N_6892);
or U13885 (N_13885,N_9166,N_6787);
nand U13886 (N_13886,N_5352,N_6201);
xnor U13887 (N_13887,N_9162,N_8592);
xnor U13888 (N_13888,N_8456,N_9476);
and U13889 (N_13889,N_6222,N_8472);
nand U13890 (N_13890,N_8162,N_7804);
xor U13891 (N_13891,N_9068,N_7080);
xnor U13892 (N_13892,N_8288,N_5829);
nor U13893 (N_13893,N_5851,N_6322);
nor U13894 (N_13894,N_5658,N_8628);
and U13895 (N_13895,N_7387,N_6845);
and U13896 (N_13896,N_8060,N_6999);
and U13897 (N_13897,N_9381,N_6131);
nor U13898 (N_13898,N_7661,N_7509);
xor U13899 (N_13899,N_6490,N_8799);
and U13900 (N_13900,N_9779,N_6428);
nor U13901 (N_13901,N_8177,N_5642);
or U13902 (N_13902,N_5459,N_7082);
and U13903 (N_13903,N_8468,N_8617);
and U13904 (N_13904,N_9770,N_5495);
xor U13905 (N_13905,N_7480,N_6876);
or U13906 (N_13906,N_8502,N_5666);
and U13907 (N_13907,N_5623,N_7600);
and U13908 (N_13908,N_7125,N_9790);
xor U13909 (N_13909,N_5834,N_7858);
or U13910 (N_13910,N_5641,N_8020);
xnor U13911 (N_13911,N_7409,N_8660);
or U13912 (N_13912,N_7655,N_7475);
or U13913 (N_13913,N_9508,N_8501);
and U13914 (N_13914,N_5444,N_8688);
nand U13915 (N_13915,N_6854,N_9288);
nand U13916 (N_13916,N_8870,N_5044);
or U13917 (N_13917,N_5086,N_9574);
and U13918 (N_13918,N_8703,N_9358);
and U13919 (N_13919,N_6509,N_8033);
nor U13920 (N_13920,N_8086,N_9235);
xnor U13921 (N_13921,N_8235,N_9498);
and U13922 (N_13922,N_5518,N_7944);
nor U13923 (N_13923,N_7501,N_7859);
and U13924 (N_13924,N_6815,N_5041);
xnor U13925 (N_13925,N_7048,N_5268);
xnor U13926 (N_13926,N_7396,N_5353);
or U13927 (N_13927,N_8075,N_5506);
nand U13928 (N_13928,N_5587,N_7156);
nand U13929 (N_13929,N_5689,N_7148);
and U13930 (N_13930,N_8617,N_5946);
xnor U13931 (N_13931,N_7507,N_6471);
or U13932 (N_13932,N_9243,N_9408);
xor U13933 (N_13933,N_8504,N_6244);
xnor U13934 (N_13934,N_5365,N_7286);
xor U13935 (N_13935,N_9745,N_8030);
nor U13936 (N_13936,N_8929,N_5466);
nand U13937 (N_13937,N_6199,N_8461);
xor U13938 (N_13938,N_5112,N_5928);
or U13939 (N_13939,N_6343,N_6394);
nor U13940 (N_13940,N_6629,N_6746);
and U13941 (N_13941,N_7722,N_6905);
and U13942 (N_13942,N_6424,N_6195);
nand U13943 (N_13943,N_7446,N_6164);
nor U13944 (N_13944,N_7452,N_6179);
and U13945 (N_13945,N_9846,N_9301);
nor U13946 (N_13946,N_7133,N_7964);
nor U13947 (N_13947,N_6993,N_8380);
xnor U13948 (N_13948,N_5028,N_8960);
xnor U13949 (N_13949,N_6464,N_6633);
nor U13950 (N_13950,N_5603,N_8252);
or U13951 (N_13951,N_8331,N_9379);
nand U13952 (N_13952,N_7144,N_6983);
nor U13953 (N_13953,N_5684,N_5633);
nand U13954 (N_13954,N_9869,N_6978);
nor U13955 (N_13955,N_5531,N_9623);
or U13956 (N_13956,N_9522,N_8298);
nor U13957 (N_13957,N_5224,N_5040);
nand U13958 (N_13958,N_5959,N_7534);
or U13959 (N_13959,N_6578,N_8887);
xnor U13960 (N_13960,N_7241,N_9193);
nor U13961 (N_13961,N_7910,N_9372);
nand U13962 (N_13962,N_6595,N_7185);
or U13963 (N_13963,N_6895,N_6525);
xor U13964 (N_13964,N_7261,N_6923);
and U13965 (N_13965,N_5703,N_9314);
nand U13966 (N_13966,N_5074,N_7618);
and U13967 (N_13967,N_8449,N_8015);
xnor U13968 (N_13968,N_9940,N_8252);
nor U13969 (N_13969,N_5818,N_7891);
and U13970 (N_13970,N_5311,N_8663);
nand U13971 (N_13971,N_6664,N_6553);
nand U13972 (N_13972,N_9535,N_5887);
or U13973 (N_13973,N_8189,N_5865);
or U13974 (N_13974,N_7747,N_6978);
nand U13975 (N_13975,N_8792,N_7613);
and U13976 (N_13976,N_9720,N_8596);
and U13977 (N_13977,N_9367,N_5432);
nor U13978 (N_13978,N_7653,N_8112);
xor U13979 (N_13979,N_7409,N_8875);
xor U13980 (N_13980,N_5589,N_6812);
xor U13981 (N_13981,N_7819,N_6693);
and U13982 (N_13982,N_5529,N_5544);
and U13983 (N_13983,N_9397,N_8460);
xor U13984 (N_13984,N_8421,N_5819);
and U13985 (N_13985,N_6176,N_8995);
nor U13986 (N_13986,N_5857,N_7890);
and U13987 (N_13987,N_5441,N_6427);
or U13988 (N_13988,N_5952,N_9014);
or U13989 (N_13989,N_7473,N_6501);
or U13990 (N_13990,N_6222,N_7265);
or U13991 (N_13991,N_8690,N_5026);
nand U13992 (N_13992,N_6856,N_6343);
or U13993 (N_13993,N_7358,N_6946);
nor U13994 (N_13994,N_8712,N_9859);
nor U13995 (N_13995,N_5748,N_7917);
xor U13996 (N_13996,N_7300,N_8505);
nand U13997 (N_13997,N_8189,N_5698);
nand U13998 (N_13998,N_9300,N_8255);
nor U13999 (N_13999,N_7396,N_5793);
or U14000 (N_14000,N_5774,N_8508);
nor U14001 (N_14001,N_8927,N_6483);
xor U14002 (N_14002,N_6880,N_5934);
and U14003 (N_14003,N_5493,N_8927);
and U14004 (N_14004,N_7350,N_8621);
and U14005 (N_14005,N_7333,N_5519);
and U14006 (N_14006,N_7701,N_5514);
xor U14007 (N_14007,N_7329,N_5517);
xor U14008 (N_14008,N_6866,N_8524);
or U14009 (N_14009,N_6428,N_7410);
nand U14010 (N_14010,N_8556,N_7467);
nand U14011 (N_14011,N_5850,N_6904);
and U14012 (N_14012,N_9163,N_9551);
and U14013 (N_14013,N_9414,N_8519);
and U14014 (N_14014,N_9570,N_8240);
or U14015 (N_14015,N_5507,N_9134);
nor U14016 (N_14016,N_8441,N_8920);
or U14017 (N_14017,N_8308,N_8592);
xnor U14018 (N_14018,N_8941,N_9358);
xnor U14019 (N_14019,N_6073,N_7189);
and U14020 (N_14020,N_5199,N_6259);
or U14021 (N_14021,N_5259,N_7172);
or U14022 (N_14022,N_7571,N_7791);
or U14023 (N_14023,N_9765,N_7646);
and U14024 (N_14024,N_9550,N_9194);
nor U14025 (N_14025,N_9545,N_7116);
and U14026 (N_14026,N_7656,N_6618);
xnor U14027 (N_14027,N_6035,N_6664);
and U14028 (N_14028,N_5851,N_8024);
xnor U14029 (N_14029,N_5748,N_6713);
and U14030 (N_14030,N_5333,N_5956);
nor U14031 (N_14031,N_6934,N_7491);
and U14032 (N_14032,N_5925,N_5094);
xor U14033 (N_14033,N_9551,N_5180);
xnor U14034 (N_14034,N_7311,N_7034);
nand U14035 (N_14035,N_9553,N_6693);
nor U14036 (N_14036,N_5482,N_6205);
nand U14037 (N_14037,N_6079,N_6952);
and U14038 (N_14038,N_5786,N_7072);
and U14039 (N_14039,N_9100,N_5281);
nor U14040 (N_14040,N_7739,N_5337);
and U14041 (N_14041,N_8352,N_5001);
nand U14042 (N_14042,N_5567,N_6205);
nor U14043 (N_14043,N_7777,N_5878);
and U14044 (N_14044,N_9594,N_5187);
and U14045 (N_14045,N_8582,N_8366);
and U14046 (N_14046,N_6134,N_6288);
or U14047 (N_14047,N_5556,N_5343);
nor U14048 (N_14048,N_9574,N_7215);
xor U14049 (N_14049,N_9816,N_7392);
nand U14050 (N_14050,N_7510,N_6903);
xnor U14051 (N_14051,N_9004,N_9025);
nand U14052 (N_14052,N_5687,N_7119);
nand U14053 (N_14053,N_9614,N_9603);
and U14054 (N_14054,N_6536,N_9408);
and U14055 (N_14055,N_8234,N_6603);
or U14056 (N_14056,N_5565,N_6708);
or U14057 (N_14057,N_7012,N_5604);
and U14058 (N_14058,N_7697,N_5770);
nor U14059 (N_14059,N_5626,N_5499);
xnor U14060 (N_14060,N_8462,N_8597);
xnor U14061 (N_14061,N_9324,N_6553);
xnor U14062 (N_14062,N_8598,N_8210);
nor U14063 (N_14063,N_9475,N_8054);
and U14064 (N_14064,N_5791,N_6050);
or U14065 (N_14065,N_8172,N_6447);
xnor U14066 (N_14066,N_7363,N_8660);
xor U14067 (N_14067,N_9504,N_8884);
xnor U14068 (N_14068,N_9431,N_7540);
xnor U14069 (N_14069,N_6685,N_6094);
or U14070 (N_14070,N_9201,N_6995);
xor U14071 (N_14071,N_8468,N_6384);
nand U14072 (N_14072,N_9105,N_8674);
and U14073 (N_14073,N_8118,N_5763);
nand U14074 (N_14074,N_7084,N_8284);
or U14075 (N_14075,N_6738,N_8697);
or U14076 (N_14076,N_5567,N_9836);
and U14077 (N_14077,N_9234,N_9341);
or U14078 (N_14078,N_5348,N_9732);
and U14079 (N_14079,N_7243,N_6447);
xor U14080 (N_14080,N_6439,N_5988);
nand U14081 (N_14081,N_9582,N_7870);
and U14082 (N_14082,N_9163,N_9311);
xor U14083 (N_14083,N_7856,N_6321);
nand U14084 (N_14084,N_7929,N_8288);
and U14085 (N_14085,N_9392,N_9734);
and U14086 (N_14086,N_8052,N_7685);
and U14087 (N_14087,N_5982,N_9783);
nor U14088 (N_14088,N_6398,N_9791);
xnor U14089 (N_14089,N_8927,N_5027);
nor U14090 (N_14090,N_6280,N_8104);
xor U14091 (N_14091,N_8920,N_6586);
xor U14092 (N_14092,N_9711,N_9566);
nor U14093 (N_14093,N_8379,N_7674);
nor U14094 (N_14094,N_7972,N_9247);
or U14095 (N_14095,N_6346,N_8127);
nand U14096 (N_14096,N_5526,N_5098);
or U14097 (N_14097,N_8269,N_8113);
nor U14098 (N_14098,N_6363,N_5001);
nor U14099 (N_14099,N_8204,N_8469);
or U14100 (N_14100,N_7407,N_5994);
and U14101 (N_14101,N_9284,N_8802);
or U14102 (N_14102,N_6405,N_6449);
xor U14103 (N_14103,N_6675,N_6854);
nor U14104 (N_14104,N_9179,N_6352);
xor U14105 (N_14105,N_8475,N_8123);
nor U14106 (N_14106,N_8813,N_7847);
or U14107 (N_14107,N_8274,N_7208);
nor U14108 (N_14108,N_6093,N_8701);
xnor U14109 (N_14109,N_8235,N_5170);
and U14110 (N_14110,N_9056,N_5795);
or U14111 (N_14111,N_7755,N_8513);
or U14112 (N_14112,N_8919,N_5899);
nand U14113 (N_14113,N_8510,N_9960);
xnor U14114 (N_14114,N_7022,N_6503);
nor U14115 (N_14115,N_9868,N_6419);
xor U14116 (N_14116,N_8903,N_9432);
and U14117 (N_14117,N_8223,N_9851);
xnor U14118 (N_14118,N_6610,N_6167);
nand U14119 (N_14119,N_9235,N_6542);
nor U14120 (N_14120,N_5007,N_5439);
xor U14121 (N_14121,N_6765,N_9629);
or U14122 (N_14122,N_5831,N_6877);
or U14123 (N_14123,N_7114,N_6273);
nand U14124 (N_14124,N_6752,N_8470);
nand U14125 (N_14125,N_5926,N_8316);
and U14126 (N_14126,N_6069,N_6448);
or U14127 (N_14127,N_7019,N_6785);
nand U14128 (N_14128,N_6212,N_8233);
nand U14129 (N_14129,N_6728,N_9604);
and U14130 (N_14130,N_7152,N_6778);
nand U14131 (N_14131,N_9940,N_6549);
nand U14132 (N_14132,N_7986,N_5370);
nand U14133 (N_14133,N_5733,N_5510);
and U14134 (N_14134,N_5646,N_8086);
or U14135 (N_14135,N_6878,N_8895);
nand U14136 (N_14136,N_6495,N_7320);
nor U14137 (N_14137,N_7347,N_6053);
and U14138 (N_14138,N_8238,N_6988);
or U14139 (N_14139,N_8979,N_6326);
xor U14140 (N_14140,N_7042,N_7790);
xnor U14141 (N_14141,N_9675,N_5941);
or U14142 (N_14142,N_5644,N_9899);
and U14143 (N_14143,N_9177,N_9107);
and U14144 (N_14144,N_7713,N_9404);
or U14145 (N_14145,N_7495,N_9310);
nand U14146 (N_14146,N_6917,N_5507);
xnor U14147 (N_14147,N_5618,N_7480);
nand U14148 (N_14148,N_6256,N_8353);
and U14149 (N_14149,N_8529,N_8340);
nor U14150 (N_14150,N_6792,N_9572);
nand U14151 (N_14151,N_6479,N_5756);
nor U14152 (N_14152,N_7323,N_7817);
nand U14153 (N_14153,N_8657,N_9802);
or U14154 (N_14154,N_9762,N_8758);
xnor U14155 (N_14155,N_9356,N_5448);
nand U14156 (N_14156,N_8887,N_7474);
and U14157 (N_14157,N_7732,N_7224);
or U14158 (N_14158,N_7687,N_9525);
or U14159 (N_14159,N_9840,N_5245);
and U14160 (N_14160,N_6492,N_8803);
nor U14161 (N_14161,N_9006,N_7181);
or U14162 (N_14162,N_5158,N_9080);
or U14163 (N_14163,N_5576,N_9478);
or U14164 (N_14164,N_8735,N_5735);
nand U14165 (N_14165,N_9100,N_6557);
nand U14166 (N_14166,N_6662,N_9602);
xor U14167 (N_14167,N_9469,N_8097);
or U14168 (N_14168,N_9113,N_6013);
nor U14169 (N_14169,N_5934,N_6977);
nor U14170 (N_14170,N_9976,N_5937);
nor U14171 (N_14171,N_8316,N_7934);
and U14172 (N_14172,N_5864,N_7899);
xor U14173 (N_14173,N_6119,N_8928);
and U14174 (N_14174,N_7558,N_6778);
nor U14175 (N_14175,N_8805,N_6984);
or U14176 (N_14176,N_8734,N_7716);
and U14177 (N_14177,N_5529,N_9209);
nor U14178 (N_14178,N_5442,N_7231);
nand U14179 (N_14179,N_5223,N_8848);
nand U14180 (N_14180,N_9938,N_6047);
or U14181 (N_14181,N_7146,N_6085);
nor U14182 (N_14182,N_7056,N_6989);
nor U14183 (N_14183,N_7008,N_7488);
xor U14184 (N_14184,N_9522,N_7934);
nand U14185 (N_14185,N_8578,N_9979);
nor U14186 (N_14186,N_7780,N_7074);
or U14187 (N_14187,N_8867,N_9420);
or U14188 (N_14188,N_7125,N_9121);
and U14189 (N_14189,N_7565,N_6507);
nor U14190 (N_14190,N_5131,N_5552);
nand U14191 (N_14191,N_9327,N_6170);
or U14192 (N_14192,N_8393,N_6287);
nand U14193 (N_14193,N_6970,N_8728);
nand U14194 (N_14194,N_8193,N_9409);
or U14195 (N_14195,N_8984,N_5715);
or U14196 (N_14196,N_7604,N_7875);
and U14197 (N_14197,N_9601,N_9314);
xor U14198 (N_14198,N_8640,N_7685);
xnor U14199 (N_14199,N_7388,N_5531);
xor U14200 (N_14200,N_8771,N_9292);
or U14201 (N_14201,N_9910,N_8012);
and U14202 (N_14202,N_6569,N_5912);
xor U14203 (N_14203,N_8508,N_5494);
or U14204 (N_14204,N_6519,N_5502);
nor U14205 (N_14205,N_6728,N_5757);
nor U14206 (N_14206,N_5289,N_9499);
xor U14207 (N_14207,N_9694,N_6443);
nor U14208 (N_14208,N_8752,N_8866);
nor U14209 (N_14209,N_8108,N_7652);
nand U14210 (N_14210,N_5223,N_9367);
nand U14211 (N_14211,N_5503,N_8679);
xnor U14212 (N_14212,N_7879,N_7451);
or U14213 (N_14213,N_7569,N_6248);
xnor U14214 (N_14214,N_7013,N_5655);
or U14215 (N_14215,N_8956,N_9163);
xor U14216 (N_14216,N_5523,N_9544);
or U14217 (N_14217,N_8624,N_9340);
or U14218 (N_14218,N_7485,N_5065);
or U14219 (N_14219,N_8696,N_8127);
and U14220 (N_14220,N_9698,N_9531);
or U14221 (N_14221,N_6720,N_5882);
xor U14222 (N_14222,N_7449,N_9021);
and U14223 (N_14223,N_7490,N_5720);
xor U14224 (N_14224,N_8602,N_5805);
and U14225 (N_14225,N_6465,N_9668);
xor U14226 (N_14226,N_9443,N_9851);
or U14227 (N_14227,N_7647,N_6323);
and U14228 (N_14228,N_7145,N_9493);
and U14229 (N_14229,N_7841,N_9649);
or U14230 (N_14230,N_6820,N_8963);
and U14231 (N_14231,N_7223,N_6119);
and U14232 (N_14232,N_8337,N_9725);
and U14233 (N_14233,N_9821,N_8796);
and U14234 (N_14234,N_8099,N_5019);
nand U14235 (N_14235,N_5215,N_7631);
or U14236 (N_14236,N_5609,N_9182);
and U14237 (N_14237,N_9327,N_9069);
or U14238 (N_14238,N_5018,N_5124);
or U14239 (N_14239,N_5110,N_9480);
or U14240 (N_14240,N_5558,N_8475);
and U14241 (N_14241,N_9363,N_5727);
xnor U14242 (N_14242,N_9984,N_5334);
nor U14243 (N_14243,N_6831,N_7037);
xnor U14244 (N_14244,N_5753,N_9861);
and U14245 (N_14245,N_8670,N_8493);
and U14246 (N_14246,N_6600,N_8010);
and U14247 (N_14247,N_6285,N_6398);
xnor U14248 (N_14248,N_7653,N_8427);
nor U14249 (N_14249,N_6335,N_6829);
and U14250 (N_14250,N_8523,N_5152);
and U14251 (N_14251,N_7779,N_9373);
or U14252 (N_14252,N_6558,N_7165);
nor U14253 (N_14253,N_7508,N_9048);
and U14254 (N_14254,N_5052,N_9404);
xnor U14255 (N_14255,N_5553,N_8526);
or U14256 (N_14256,N_7088,N_5091);
xor U14257 (N_14257,N_7960,N_5645);
nor U14258 (N_14258,N_9133,N_6995);
or U14259 (N_14259,N_5979,N_5844);
and U14260 (N_14260,N_7473,N_8734);
and U14261 (N_14261,N_5209,N_9186);
nor U14262 (N_14262,N_9844,N_9144);
xor U14263 (N_14263,N_7125,N_6183);
or U14264 (N_14264,N_5172,N_6614);
nand U14265 (N_14265,N_6367,N_8206);
nand U14266 (N_14266,N_8976,N_8947);
and U14267 (N_14267,N_6942,N_8305);
nor U14268 (N_14268,N_5059,N_7358);
and U14269 (N_14269,N_5128,N_8116);
xor U14270 (N_14270,N_8415,N_9888);
nor U14271 (N_14271,N_8201,N_8664);
xor U14272 (N_14272,N_7771,N_5351);
xnor U14273 (N_14273,N_7451,N_7142);
nor U14274 (N_14274,N_9042,N_8828);
and U14275 (N_14275,N_9089,N_8739);
or U14276 (N_14276,N_9801,N_7825);
and U14277 (N_14277,N_8669,N_8404);
or U14278 (N_14278,N_5630,N_8087);
xor U14279 (N_14279,N_7253,N_7706);
and U14280 (N_14280,N_9826,N_8188);
nand U14281 (N_14281,N_6345,N_8038);
and U14282 (N_14282,N_9994,N_7386);
xnor U14283 (N_14283,N_9495,N_6355);
nand U14284 (N_14284,N_7271,N_6723);
and U14285 (N_14285,N_5543,N_6436);
nand U14286 (N_14286,N_9493,N_6629);
nor U14287 (N_14287,N_6380,N_6907);
or U14288 (N_14288,N_7527,N_8122);
nand U14289 (N_14289,N_6243,N_9940);
or U14290 (N_14290,N_8361,N_6895);
and U14291 (N_14291,N_5196,N_8915);
nand U14292 (N_14292,N_6901,N_6326);
xor U14293 (N_14293,N_7470,N_8111);
or U14294 (N_14294,N_5233,N_9243);
or U14295 (N_14295,N_9116,N_5458);
and U14296 (N_14296,N_6929,N_6193);
nand U14297 (N_14297,N_5611,N_8431);
nor U14298 (N_14298,N_8612,N_6676);
and U14299 (N_14299,N_8040,N_6094);
nand U14300 (N_14300,N_9163,N_7756);
and U14301 (N_14301,N_7102,N_5123);
nand U14302 (N_14302,N_9858,N_6393);
nor U14303 (N_14303,N_7108,N_6787);
or U14304 (N_14304,N_7095,N_6187);
and U14305 (N_14305,N_8359,N_9030);
and U14306 (N_14306,N_6974,N_5860);
nand U14307 (N_14307,N_7653,N_9486);
nor U14308 (N_14308,N_5585,N_9538);
or U14309 (N_14309,N_9839,N_5338);
nand U14310 (N_14310,N_8321,N_6479);
xnor U14311 (N_14311,N_7355,N_6653);
or U14312 (N_14312,N_7099,N_6033);
xnor U14313 (N_14313,N_5691,N_8908);
nand U14314 (N_14314,N_7505,N_5751);
or U14315 (N_14315,N_9800,N_6017);
xor U14316 (N_14316,N_9173,N_7857);
nand U14317 (N_14317,N_6678,N_5278);
xnor U14318 (N_14318,N_6211,N_8198);
xor U14319 (N_14319,N_6412,N_9768);
or U14320 (N_14320,N_6878,N_5498);
or U14321 (N_14321,N_5725,N_8782);
or U14322 (N_14322,N_6486,N_8671);
or U14323 (N_14323,N_9781,N_8147);
nor U14324 (N_14324,N_7727,N_6122);
nand U14325 (N_14325,N_6597,N_8132);
nor U14326 (N_14326,N_8948,N_5882);
and U14327 (N_14327,N_9112,N_7276);
and U14328 (N_14328,N_6661,N_8706);
nand U14329 (N_14329,N_8493,N_6820);
or U14330 (N_14330,N_5904,N_8700);
and U14331 (N_14331,N_5612,N_9135);
or U14332 (N_14332,N_6248,N_8537);
nand U14333 (N_14333,N_9979,N_7299);
xnor U14334 (N_14334,N_9616,N_5474);
or U14335 (N_14335,N_7433,N_7043);
nand U14336 (N_14336,N_6416,N_5265);
xnor U14337 (N_14337,N_6659,N_5259);
or U14338 (N_14338,N_7519,N_5057);
nand U14339 (N_14339,N_7737,N_8573);
nand U14340 (N_14340,N_9743,N_6715);
and U14341 (N_14341,N_8326,N_9160);
or U14342 (N_14342,N_6035,N_6725);
and U14343 (N_14343,N_8745,N_8609);
xor U14344 (N_14344,N_9959,N_6692);
or U14345 (N_14345,N_8953,N_9870);
nand U14346 (N_14346,N_6586,N_5809);
nand U14347 (N_14347,N_8053,N_7687);
nand U14348 (N_14348,N_6358,N_8874);
and U14349 (N_14349,N_9908,N_8685);
xnor U14350 (N_14350,N_5559,N_5975);
and U14351 (N_14351,N_6164,N_8653);
and U14352 (N_14352,N_6352,N_5273);
xnor U14353 (N_14353,N_7657,N_6291);
or U14354 (N_14354,N_8106,N_5424);
and U14355 (N_14355,N_5497,N_5474);
nand U14356 (N_14356,N_7372,N_9259);
xnor U14357 (N_14357,N_7120,N_5064);
nor U14358 (N_14358,N_5894,N_9525);
xor U14359 (N_14359,N_6839,N_7555);
xnor U14360 (N_14360,N_6434,N_6216);
xor U14361 (N_14361,N_8449,N_6256);
xnor U14362 (N_14362,N_9466,N_8060);
xnor U14363 (N_14363,N_5775,N_7875);
nand U14364 (N_14364,N_9397,N_6775);
or U14365 (N_14365,N_9116,N_8859);
or U14366 (N_14366,N_8073,N_6975);
xnor U14367 (N_14367,N_9012,N_5244);
xnor U14368 (N_14368,N_6410,N_6612);
nor U14369 (N_14369,N_8995,N_7088);
nor U14370 (N_14370,N_6070,N_8998);
nand U14371 (N_14371,N_7059,N_9659);
nor U14372 (N_14372,N_9830,N_6786);
nand U14373 (N_14373,N_8939,N_7035);
or U14374 (N_14374,N_9431,N_6266);
or U14375 (N_14375,N_8686,N_7125);
nand U14376 (N_14376,N_8083,N_6809);
nand U14377 (N_14377,N_5945,N_5415);
xor U14378 (N_14378,N_8219,N_8027);
xor U14379 (N_14379,N_9985,N_9553);
or U14380 (N_14380,N_7648,N_6574);
nand U14381 (N_14381,N_9801,N_6845);
xor U14382 (N_14382,N_8912,N_7064);
xnor U14383 (N_14383,N_7609,N_8826);
or U14384 (N_14384,N_5759,N_5289);
nor U14385 (N_14385,N_7150,N_5841);
xor U14386 (N_14386,N_8255,N_8078);
nand U14387 (N_14387,N_5343,N_5866);
and U14388 (N_14388,N_5084,N_9355);
or U14389 (N_14389,N_9889,N_7226);
xor U14390 (N_14390,N_5317,N_9232);
nor U14391 (N_14391,N_8022,N_6302);
or U14392 (N_14392,N_5590,N_6341);
nor U14393 (N_14393,N_6149,N_7280);
xor U14394 (N_14394,N_6166,N_9367);
or U14395 (N_14395,N_5939,N_9959);
nand U14396 (N_14396,N_8556,N_9141);
xnor U14397 (N_14397,N_5626,N_5072);
or U14398 (N_14398,N_6953,N_6767);
nand U14399 (N_14399,N_5774,N_9242);
or U14400 (N_14400,N_5088,N_9117);
or U14401 (N_14401,N_6739,N_8440);
nor U14402 (N_14402,N_7638,N_6218);
and U14403 (N_14403,N_8695,N_8143);
nand U14404 (N_14404,N_5976,N_6547);
or U14405 (N_14405,N_9898,N_9195);
or U14406 (N_14406,N_8242,N_9097);
and U14407 (N_14407,N_7560,N_9422);
and U14408 (N_14408,N_8036,N_8071);
or U14409 (N_14409,N_6667,N_9744);
xnor U14410 (N_14410,N_9977,N_8443);
or U14411 (N_14411,N_5006,N_9927);
and U14412 (N_14412,N_7987,N_9220);
xor U14413 (N_14413,N_6485,N_5592);
nor U14414 (N_14414,N_9819,N_8776);
nand U14415 (N_14415,N_5768,N_8926);
nor U14416 (N_14416,N_7578,N_8248);
nand U14417 (N_14417,N_8847,N_9521);
nand U14418 (N_14418,N_7975,N_7057);
nor U14419 (N_14419,N_5786,N_6415);
and U14420 (N_14420,N_7563,N_6939);
xor U14421 (N_14421,N_8598,N_5068);
xor U14422 (N_14422,N_6480,N_7028);
and U14423 (N_14423,N_8112,N_7951);
or U14424 (N_14424,N_5170,N_6085);
or U14425 (N_14425,N_5351,N_6427);
and U14426 (N_14426,N_8977,N_5608);
nor U14427 (N_14427,N_7932,N_8986);
nor U14428 (N_14428,N_9160,N_7884);
xor U14429 (N_14429,N_8188,N_6932);
and U14430 (N_14430,N_9698,N_5379);
nor U14431 (N_14431,N_8183,N_8333);
nor U14432 (N_14432,N_7293,N_6943);
or U14433 (N_14433,N_5210,N_8509);
and U14434 (N_14434,N_7682,N_9565);
or U14435 (N_14435,N_8348,N_5902);
nand U14436 (N_14436,N_6996,N_5612);
or U14437 (N_14437,N_7363,N_9112);
and U14438 (N_14438,N_7581,N_6220);
or U14439 (N_14439,N_7771,N_8969);
or U14440 (N_14440,N_6733,N_8443);
nor U14441 (N_14441,N_9193,N_7851);
xor U14442 (N_14442,N_8485,N_9500);
xor U14443 (N_14443,N_6677,N_9985);
nor U14444 (N_14444,N_8019,N_9042);
nor U14445 (N_14445,N_7870,N_8891);
xor U14446 (N_14446,N_9827,N_9506);
and U14447 (N_14447,N_5685,N_7540);
xor U14448 (N_14448,N_7012,N_6550);
and U14449 (N_14449,N_8900,N_9756);
nor U14450 (N_14450,N_7071,N_8105);
and U14451 (N_14451,N_8822,N_5894);
and U14452 (N_14452,N_6217,N_7975);
and U14453 (N_14453,N_7353,N_7480);
and U14454 (N_14454,N_5294,N_8952);
nor U14455 (N_14455,N_6660,N_7566);
nor U14456 (N_14456,N_5794,N_8068);
and U14457 (N_14457,N_5586,N_6747);
nand U14458 (N_14458,N_9345,N_8713);
xor U14459 (N_14459,N_6032,N_7489);
nand U14460 (N_14460,N_6966,N_5702);
nand U14461 (N_14461,N_9757,N_9527);
xor U14462 (N_14462,N_9975,N_7300);
and U14463 (N_14463,N_5212,N_9529);
xor U14464 (N_14464,N_5360,N_8836);
nor U14465 (N_14465,N_7453,N_8039);
nor U14466 (N_14466,N_9009,N_5940);
nor U14467 (N_14467,N_8974,N_5800);
nor U14468 (N_14468,N_7665,N_9392);
and U14469 (N_14469,N_7125,N_7221);
and U14470 (N_14470,N_8234,N_6686);
and U14471 (N_14471,N_9118,N_7464);
or U14472 (N_14472,N_5397,N_6637);
nand U14473 (N_14473,N_9436,N_6060);
nand U14474 (N_14474,N_9537,N_8565);
or U14475 (N_14475,N_9426,N_6319);
nand U14476 (N_14476,N_7877,N_6278);
nand U14477 (N_14477,N_9450,N_8154);
nor U14478 (N_14478,N_5243,N_9689);
nor U14479 (N_14479,N_6800,N_9951);
xor U14480 (N_14480,N_6718,N_7954);
or U14481 (N_14481,N_7450,N_5872);
xor U14482 (N_14482,N_6262,N_7640);
or U14483 (N_14483,N_6296,N_5197);
nor U14484 (N_14484,N_6410,N_9034);
nand U14485 (N_14485,N_8244,N_5181);
nor U14486 (N_14486,N_9577,N_8574);
and U14487 (N_14487,N_6202,N_9275);
or U14488 (N_14488,N_7161,N_7941);
or U14489 (N_14489,N_9564,N_8500);
or U14490 (N_14490,N_6798,N_8927);
nand U14491 (N_14491,N_9647,N_8264);
xor U14492 (N_14492,N_6134,N_6344);
and U14493 (N_14493,N_8028,N_6481);
or U14494 (N_14494,N_9817,N_9407);
nand U14495 (N_14495,N_8057,N_7140);
or U14496 (N_14496,N_8621,N_6577);
nor U14497 (N_14497,N_8386,N_5660);
xor U14498 (N_14498,N_5751,N_7935);
or U14499 (N_14499,N_5784,N_7509);
or U14500 (N_14500,N_5810,N_9759);
nor U14501 (N_14501,N_6733,N_8873);
xor U14502 (N_14502,N_6603,N_9049);
xnor U14503 (N_14503,N_8152,N_7365);
nand U14504 (N_14504,N_7391,N_8352);
nor U14505 (N_14505,N_7705,N_6309);
xor U14506 (N_14506,N_9201,N_6695);
xor U14507 (N_14507,N_6972,N_6429);
and U14508 (N_14508,N_8221,N_5626);
nand U14509 (N_14509,N_7757,N_6434);
nor U14510 (N_14510,N_9099,N_6719);
or U14511 (N_14511,N_9240,N_6801);
xor U14512 (N_14512,N_6642,N_7073);
nor U14513 (N_14513,N_9220,N_7608);
or U14514 (N_14514,N_5046,N_6213);
xor U14515 (N_14515,N_9557,N_5258);
xnor U14516 (N_14516,N_5969,N_9412);
nor U14517 (N_14517,N_9522,N_7728);
and U14518 (N_14518,N_5482,N_7885);
or U14519 (N_14519,N_9534,N_9635);
xnor U14520 (N_14520,N_9252,N_7892);
or U14521 (N_14521,N_8813,N_6838);
and U14522 (N_14522,N_9622,N_6922);
or U14523 (N_14523,N_8566,N_9465);
nor U14524 (N_14524,N_6157,N_6831);
nor U14525 (N_14525,N_9902,N_7146);
or U14526 (N_14526,N_7880,N_8556);
nor U14527 (N_14527,N_6072,N_9002);
and U14528 (N_14528,N_7130,N_8393);
and U14529 (N_14529,N_7105,N_8148);
nand U14530 (N_14530,N_9966,N_7281);
nand U14531 (N_14531,N_8036,N_6273);
or U14532 (N_14532,N_6276,N_6992);
nand U14533 (N_14533,N_7274,N_6316);
and U14534 (N_14534,N_8701,N_5817);
xor U14535 (N_14535,N_9922,N_8789);
nor U14536 (N_14536,N_5862,N_5902);
nand U14537 (N_14537,N_5305,N_5140);
nor U14538 (N_14538,N_9749,N_8183);
and U14539 (N_14539,N_6139,N_5720);
or U14540 (N_14540,N_7064,N_9109);
and U14541 (N_14541,N_8812,N_8274);
or U14542 (N_14542,N_7282,N_5532);
and U14543 (N_14543,N_8448,N_6151);
nor U14544 (N_14544,N_6327,N_5543);
or U14545 (N_14545,N_6324,N_7235);
and U14546 (N_14546,N_5195,N_7228);
nor U14547 (N_14547,N_9695,N_7291);
nand U14548 (N_14548,N_7717,N_8750);
xor U14549 (N_14549,N_8051,N_6412);
and U14550 (N_14550,N_8958,N_5146);
nor U14551 (N_14551,N_8406,N_9540);
xnor U14552 (N_14552,N_9221,N_9832);
or U14553 (N_14553,N_8711,N_8927);
nand U14554 (N_14554,N_6167,N_9530);
xnor U14555 (N_14555,N_9584,N_7192);
nor U14556 (N_14556,N_7671,N_6500);
nand U14557 (N_14557,N_5718,N_8436);
nand U14558 (N_14558,N_5632,N_8311);
and U14559 (N_14559,N_8859,N_7688);
nor U14560 (N_14560,N_7445,N_8081);
xor U14561 (N_14561,N_5019,N_8672);
or U14562 (N_14562,N_6199,N_6755);
nand U14563 (N_14563,N_9916,N_6238);
nor U14564 (N_14564,N_9170,N_5956);
nand U14565 (N_14565,N_7702,N_9576);
and U14566 (N_14566,N_8871,N_7186);
xnor U14567 (N_14567,N_9858,N_5428);
nor U14568 (N_14568,N_5164,N_9129);
or U14569 (N_14569,N_8086,N_5584);
or U14570 (N_14570,N_8025,N_9952);
nand U14571 (N_14571,N_5414,N_5547);
nand U14572 (N_14572,N_6987,N_5446);
and U14573 (N_14573,N_8937,N_6801);
or U14574 (N_14574,N_9568,N_6274);
xor U14575 (N_14575,N_9980,N_8596);
xnor U14576 (N_14576,N_9092,N_6063);
or U14577 (N_14577,N_9449,N_6586);
nand U14578 (N_14578,N_9938,N_7912);
or U14579 (N_14579,N_5564,N_6426);
or U14580 (N_14580,N_9589,N_6131);
xnor U14581 (N_14581,N_9185,N_9321);
or U14582 (N_14582,N_8774,N_9939);
nand U14583 (N_14583,N_8281,N_6143);
nor U14584 (N_14584,N_9876,N_8408);
nor U14585 (N_14585,N_5445,N_6940);
and U14586 (N_14586,N_5070,N_8445);
and U14587 (N_14587,N_7614,N_8351);
xor U14588 (N_14588,N_8584,N_5120);
and U14589 (N_14589,N_8399,N_7665);
and U14590 (N_14590,N_9565,N_5356);
nor U14591 (N_14591,N_7404,N_5443);
nor U14592 (N_14592,N_6224,N_5583);
nand U14593 (N_14593,N_6136,N_8040);
nor U14594 (N_14594,N_5416,N_9396);
or U14595 (N_14595,N_9890,N_6649);
nor U14596 (N_14596,N_7715,N_7989);
nand U14597 (N_14597,N_5199,N_8641);
or U14598 (N_14598,N_6961,N_9115);
xnor U14599 (N_14599,N_9909,N_9357);
and U14600 (N_14600,N_8143,N_5910);
and U14601 (N_14601,N_8292,N_8293);
nor U14602 (N_14602,N_5007,N_9051);
and U14603 (N_14603,N_8658,N_6043);
and U14604 (N_14604,N_6931,N_9607);
or U14605 (N_14605,N_8329,N_9407);
nand U14606 (N_14606,N_6664,N_6602);
and U14607 (N_14607,N_5492,N_8895);
nor U14608 (N_14608,N_9825,N_8413);
nor U14609 (N_14609,N_8108,N_5252);
xor U14610 (N_14610,N_7300,N_9258);
and U14611 (N_14611,N_5424,N_6005);
and U14612 (N_14612,N_5063,N_7712);
or U14613 (N_14613,N_7050,N_8246);
xnor U14614 (N_14614,N_8696,N_5954);
nand U14615 (N_14615,N_8753,N_6517);
or U14616 (N_14616,N_6056,N_7144);
nor U14617 (N_14617,N_7708,N_6744);
nor U14618 (N_14618,N_7782,N_6920);
and U14619 (N_14619,N_5600,N_7893);
nor U14620 (N_14620,N_9892,N_7071);
or U14621 (N_14621,N_9257,N_7582);
xor U14622 (N_14622,N_6212,N_8359);
and U14623 (N_14623,N_5797,N_5498);
nor U14624 (N_14624,N_6017,N_6577);
nor U14625 (N_14625,N_8205,N_5053);
xor U14626 (N_14626,N_9687,N_7171);
and U14627 (N_14627,N_7963,N_6758);
and U14628 (N_14628,N_9237,N_5570);
and U14629 (N_14629,N_9912,N_6069);
xor U14630 (N_14630,N_9481,N_6658);
and U14631 (N_14631,N_6489,N_8854);
xnor U14632 (N_14632,N_5019,N_6466);
or U14633 (N_14633,N_6447,N_7525);
nor U14634 (N_14634,N_5834,N_9431);
xor U14635 (N_14635,N_8156,N_6794);
and U14636 (N_14636,N_8799,N_5930);
and U14637 (N_14637,N_8588,N_9053);
nor U14638 (N_14638,N_9848,N_8417);
or U14639 (N_14639,N_8607,N_5871);
or U14640 (N_14640,N_6778,N_6214);
or U14641 (N_14641,N_8783,N_6713);
and U14642 (N_14642,N_8153,N_5798);
nand U14643 (N_14643,N_7014,N_7259);
xor U14644 (N_14644,N_7310,N_6881);
xnor U14645 (N_14645,N_9160,N_6186);
nor U14646 (N_14646,N_9098,N_8562);
and U14647 (N_14647,N_9760,N_5883);
xnor U14648 (N_14648,N_5604,N_5366);
nor U14649 (N_14649,N_7162,N_6966);
nor U14650 (N_14650,N_9877,N_6945);
nor U14651 (N_14651,N_5339,N_5784);
nand U14652 (N_14652,N_5058,N_5706);
nand U14653 (N_14653,N_8736,N_7565);
nand U14654 (N_14654,N_8002,N_8760);
or U14655 (N_14655,N_9995,N_8749);
and U14656 (N_14656,N_9672,N_5191);
nand U14657 (N_14657,N_7308,N_9305);
xnor U14658 (N_14658,N_7051,N_7562);
nand U14659 (N_14659,N_8903,N_8213);
nor U14660 (N_14660,N_6911,N_5096);
or U14661 (N_14661,N_5533,N_5045);
nor U14662 (N_14662,N_5935,N_5712);
and U14663 (N_14663,N_9867,N_6757);
and U14664 (N_14664,N_7385,N_5968);
xor U14665 (N_14665,N_9284,N_7861);
and U14666 (N_14666,N_8856,N_6453);
nor U14667 (N_14667,N_6892,N_5252);
nor U14668 (N_14668,N_5746,N_7965);
nand U14669 (N_14669,N_5235,N_6510);
xor U14670 (N_14670,N_5032,N_9182);
nor U14671 (N_14671,N_8022,N_7558);
xnor U14672 (N_14672,N_5731,N_5992);
xnor U14673 (N_14673,N_7333,N_5161);
and U14674 (N_14674,N_7168,N_6193);
or U14675 (N_14675,N_7533,N_7367);
nand U14676 (N_14676,N_7948,N_9692);
nor U14677 (N_14677,N_6160,N_7494);
nor U14678 (N_14678,N_9106,N_9858);
nand U14679 (N_14679,N_8222,N_8081);
nand U14680 (N_14680,N_5478,N_5148);
and U14681 (N_14681,N_6747,N_6487);
or U14682 (N_14682,N_9783,N_8048);
or U14683 (N_14683,N_9266,N_5420);
xor U14684 (N_14684,N_8659,N_6363);
xor U14685 (N_14685,N_9409,N_8970);
xor U14686 (N_14686,N_5610,N_5305);
nor U14687 (N_14687,N_6780,N_6799);
nand U14688 (N_14688,N_7922,N_8579);
and U14689 (N_14689,N_6233,N_8835);
xnor U14690 (N_14690,N_8290,N_7632);
nor U14691 (N_14691,N_9766,N_9819);
nor U14692 (N_14692,N_8805,N_6855);
nor U14693 (N_14693,N_6061,N_6743);
or U14694 (N_14694,N_9280,N_8780);
xor U14695 (N_14695,N_5121,N_8872);
nand U14696 (N_14696,N_7863,N_8115);
nor U14697 (N_14697,N_8002,N_9404);
nand U14698 (N_14698,N_9566,N_6355);
nand U14699 (N_14699,N_6684,N_9326);
nor U14700 (N_14700,N_5315,N_6699);
and U14701 (N_14701,N_9344,N_6950);
or U14702 (N_14702,N_6010,N_6233);
or U14703 (N_14703,N_6042,N_8229);
nor U14704 (N_14704,N_9426,N_5557);
and U14705 (N_14705,N_6540,N_6477);
nor U14706 (N_14706,N_9464,N_7222);
or U14707 (N_14707,N_5727,N_9562);
xor U14708 (N_14708,N_6436,N_5795);
or U14709 (N_14709,N_6999,N_6348);
or U14710 (N_14710,N_8206,N_7690);
nor U14711 (N_14711,N_5416,N_7495);
or U14712 (N_14712,N_7461,N_9950);
xor U14713 (N_14713,N_5916,N_9881);
or U14714 (N_14714,N_6733,N_5697);
and U14715 (N_14715,N_5203,N_5988);
xnor U14716 (N_14716,N_9160,N_5083);
nand U14717 (N_14717,N_7676,N_8239);
nand U14718 (N_14718,N_9302,N_7149);
nand U14719 (N_14719,N_9338,N_8441);
xnor U14720 (N_14720,N_9354,N_7212);
or U14721 (N_14721,N_8467,N_8410);
and U14722 (N_14722,N_9824,N_5458);
or U14723 (N_14723,N_5597,N_8087);
nor U14724 (N_14724,N_6408,N_7601);
or U14725 (N_14725,N_7276,N_6594);
nor U14726 (N_14726,N_6697,N_7360);
xnor U14727 (N_14727,N_7838,N_9448);
or U14728 (N_14728,N_7105,N_5378);
nor U14729 (N_14729,N_9043,N_5484);
nand U14730 (N_14730,N_8356,N_6002);
or U14731 (N_14731,N_8975,N_9933);
and U14732 (N_14732,N_6869,N_6258);
xor U14733 (N_14733,N_7612,N_5944);
xor U14734 (N_14734,N_9658,N_8668);
nor U14735 (N_14735,N_8084,N_6025);
nor U14736 (N_14736,N_7970,N_6943);
nor U14737 (N_14737,N_6967,N_9595);
or U14738 (N_14738,N_6185,N_9979);
nand U14739 (N_14739,N_8254,N_6919);
or U14740 (N_14740,N_9939,N_8749);
nand U14741 (N_14741,N_9439,N_9378);
xnor U14742 (N_14742,N_9581,N_5163);
nand U14743 (N_14743,N_9951,N_6564);
xnor U14744 (N_14744,N_7247,N_6126);
or U14745 (N_14745,N_5374,N_8660);
nor U14746 (N_14746,N_9538,N_5729);
nand U14747 (N_14747,N_6135,N_8323);
xor U14748 (N_14748,N_8641,N_7142);
nand U14749 (N_14749,N_9016,N_9991);
nor U14750 (N_14750,N_5715,N_6856);
or U14751 (N_14751,N_9285,N_9293);
or U14752 (N_14752,N_5586,N_5042);
nor U14753 (N_14753,N_7972,N_9914);
xor U14754 (N_14754,N_6648,N_9363);
nor U14755 (N_14755,N_9407,N_8234);
or U14756 (N_14756,N_5589,N_8577);
nor U14757 (N_14757,N_9923,N_8666);
or U14758 (N_14758,N_8265,N_9295);
nor U14759 (N_14759,N_8855,N_7019);
xnor U14760 (N_14760,N_9734,N_6824);
or U14761 (N_14761,N_8072,N_6251);
nor U14762 (N_14762,N_9127,N_7654);
or U14763 (N_14763,N_9332,N_8856);
or U14764 (N_14764,N_9659,N_5589);
nor U14765 (N_14765,N_7917,N_8819);
nand U14766 (N_14766,N_5840,N_8452);
nor U14767 (N_14767,N_7998,N_8345);
xnor U14768 (N_14768,N_7927,N_8500);
xor U14769 (N_14769,N_6515,N_7338);
nor U14770 (N_14770,N_8956,N_9783);
and U14771 (N_14771,N_7907,N_7659);
and U14772 (N_14772,N_9167,N_9020);
xor U14773 (N_14773,N_6054,N_7266);
xnor U14774 (N_14774,N_8012,N_8827);
nand U14775 (N_14775,N_9035,N_5317);
nor U14776 (N_14776,N_6452,N_8798);
and U14777 (N_14777,N_6651,N_7291);
and U14778 (N_14778,N_5929,N_8317);
nor U14779 (N_14779,N_8046,N_9789);
or U14780 (N_14780,N_8707,N_8624);
nand U14781 (N_14781,N_9898,N_5947);
xnor U14782 (N_14782,N_7678,N_5858);
and U14783 (N_14783,N_5748,N_7140);
and U14784 (N_14784,N_5715,N_7752);
nand U14785 (N_14785,N_6160,N_7905);
nor U14786 (N_14786,N_5492,N_5757);
nor U14787 (N_14787,N_6150,N_8212);
nand U14788 (N_14788,N_8968,N_5571);
nand U14789 (N_14789,N_8057,N_7030);
and U14790 (N_14790,N_5605,N_5213);
and U14791 (N_14791,N_7013,N_6007);
nand U14792 (N_14792,N_7024,N_6890);
nand U14793 (N_14793,N_9500,N_9393);
and U14794 (N_14794,N_9411,N_7587);
xor U14795 (N_14795,N_8788,N_9875);
xnor U14796 (N_14796,N_5318,N_9946);
nand U14797 (N_14797,N_9250,N_7109);
nor U14798 (N_14798,N_7845,N_5399);
or U14799 (N_14799,N_8443,N_7509);
nor U14800 (N_14800,N_5174,N_9721);
xor U14801 (N_14801,N_5221,N_7181);
xor U14802 (N_14802,N_9151,N_5231);
xnor U14803 (N_14803,N_7101,N_9258);
and U14804 (N_14804,N_6682,N_7118);
and U14805 (N_14805,N_7913,N_8431);
nor U14806 (N_14806,N_8037,N_9856);
nand U14807 (N_14807,N_6697,N_5996);
and U14808 (N_14808,N_9901,N_9485);
and U14809 (N_14809,N_6423,N_5103);
and U14810 (N_14810,N_6585,N_6603);
or U14811 (N_14811,N_8305,N_8501);
nor U14812 (N_14812,N_8399,N_6685);
and U14813 (N_14813,N_7449,N_6338);
or U14814 (N_14814,N_5662,N_7878);
xor U14815 (N_14815,N_6703,N_9135);
and U14816 (N_14816,N_9529,N_7927);
nand U14817 (N_14817,N_9152,N_8814);
nand U14818 (N_14818,N_9408,N_9078);
or U14819 (N_14819,N_9110,N_8796);
nor U14820 (N_14820,N_5214,N_8401);
and U14821 (N_14821,N_8128,N_7861);
and U14822 (N_14822,N_9933,N_9188);
or U14823 (N_14823,N_6240,N_8829);
nand U14824 (N_14824,N_6488,N_9226);
or U14825 (N_14825,N_6784,N_8718);
xor U14826 (N_14826,N_8909,N_9569);
nand U14827 (N_14827,N_8269,N_6724);
nor U14828 (N_14828,N_6735,N_5000);
nor U14829 (N_14829,N_5264,N_9529);
or U14830 (N_14830,N_5292,N_5785);
nand U14831 (N_14831,N_9146,N_7454);
xor U14832 (N_14832,N_7635,N_6516);
or U14833 (N_14833,N_6153,N_6623);
and U14834 (N_14834,N_7577,N_9491);
nor U14835 (N_14835,N_8972,N_5749);
and U14836 (N_14836,N_7160,N_9280);
and U14837 (N_14837,N_6551,N_7461);
or U14838 (N_14838,N_8228,N_7975);
xnor U14839 (N_14839,N_9976,N_6708);
or U14840 (N_14840,N_8590,N_7961);
and U14841 (N_14841,N_9172,N_7988);
and U14842 (N_14842,N_6360,N_9025);
and U14843 (N_14843,N_5150,N_7777);
nand U14844 (N_14844,N_9364,N_5583);
nor U14845 (N_14845,N_5012,N_8335);
or U14846 (N_14846,N_5843,N_7335);
and U14847 (N_14847,N_9346,N_8912);
xor U14848 (N_14848,N_9088,N_7628);
and U14849 (N_14849,N_8830,N_9094);
or U14850 (N_14850,N_6901,N_7200);
xnor U14851 (N_14851,N_7052,N_8321);
or U14852 (N_14852,N_6126,N_7023);
or U14853 (N_14853,N_6593,N_5174);
nand U14854 (N_14854,N_5843,N_6140);
nand U14855 (N_14855,N_7328,N_8506);
xnor U14856 (N_14856,N_5332,N_7892);
nand U14857 (N_14857,N_5820,N_7260);
and U14858 (N_14858,N_8424,N_5230);
nand U14859 (N_14859,N_9463,N_6175);
and U14860 (N_14860,N_8345,N_9942);
nor U14861 (N_14861,N_8289,N_6971);
nor U14862 (N_14862,N_8169,N_9548);
or U14863 (N_14863,N_5860,N_7878);
and U14864 (N_14864,N_5510,N_5730);
nand U14865 (N_14865,N_7149,N_7837);
nand U14866 (N_14866,N_5276,N_8363);
nor U14867 (N_14867,N_5996,N_9892);
xnor U14868 (N_14868,N_5373,N_7143);
and U14869 (N_14869,N_5410,N_6480);
nor U14870 (N_14870,N_5884,N_8203);
nand U14871 (N_14871,N_8665,N_6729);
xnor U14872 (N_14872,N_9226,N_8603);
and U14873 (N_14873,N_8306,N_8940);
nor U14874 (N_14874,N_9483,N_8410);
nor U14875 (N_14875,N_5575,N_5882);
nor U14876 (N_14876,N_8426,N_5861);
nor U14877 (N_14877,N_8190,N_8972);
and U14878 (N_14878,N_6478,N_6264);
and U14879 (N_14879,N_6198,N_6269);
or U14880 (N_14880,N_7984,N_9673);
nor U14881 (N_14881,N_6710,N_7345);
nor U14882 (N_14882,N_5211,N_7331);
xor U14883 (N_14883,N_8203,N_8892);
xor U14884 (N_14884,N_6050,N_5895);
xor U14885 (N_14885,N_9146,N_6170);
and U14886 (N_14886,N_6152,N_9776);
xnor U14887 (N_14887,N_7912,N_9338);
nor U14888 (N_14888,N_6175,N_6452);
or U14889 (N_14889,N_8538,N_9283);
or U14890 (N_14890,N_7318,N_5381);
nor U14891 (N_14891,N_7856,N_9323);
xnor U14892 (N_14892,N_5983,N_5313);
and U14893 (N_14893,N_5975,N_8432);
and U14894 (N_14894,N_7547,N_5986);
xor U14895 (N_14895,N_8133,N_7081);
nand U14896 (N_14896,N_5813,N_8172);
or U14897 (N_14897,N_7409,N_8798);
and U14898 (N_14898,N_8744,N_9271);
nand U14899 (N_14899,N_6181,N_7088);
or U14900 (N_14900,N_7406,N_5692);
and U14901 (N_14901,N_5321,N_9849);
xnor U14902 (N_14902,N_6542,N_8470);
nand U14903 (N_14903,N_7415,N_8639);
nor U14904 (N_14904,N_7054,N_5257);
xnor U14905 (N_14905,N_5277,N_9340);
nor U14906 (N_14906,N_5577,N_7333);
nor U14907 (N_14907,N_8823,N_6657);
and U14908 (N_14908,N_7021,N_8740);
or U14909 (N_14909,N_7306,N_6777);
nand U14910 (N_14910,N_8343,N_8623);
xor U14911 (N_14911,N_7423,N_5222);
and U14912 (N_14912,N_5437,N_6951);
nor U14913 (N_14913,N_6770,N_8104);
or U14914 (N_14914,N_8746,N_7998);
nand U14915 (N_14915,N_9171,N_6589);
xnor U14916 (N_14916,N_9183,N_7221);
and U14917 (N_14917,N_8779,N_8777);
nor U14918 (N_14918,N_6579,N_7512);
or U14919 (N_14919,N_6537,N_9325);
nand U14920 (N_14920,N_7551,N_5824);
nand U14921 (N_14921,N_7927,N_6956);
and U14922 (N_14922,N_8196,N_8148);
or U14923 (N_14923,N_9284,N_7162);
nand U14924 (N_14924,N_7393,N_5136);
nand U14925 (N_14925,N_7988,N_9591);
nand U14926 (N_14926,N_9949,N_6814);
nand U14927 (N_14927,N_8462,N_6016);
or U14928 (N_14928,N_7614,N_5758);
and U14929 (N_14929,N_9313,N_7334);
xnor U14930 (N_14930,N_7075,N_9107);
and U14931 (N_14931,N_8727,N_9214);
and U14932 (N_14932,N_6956,N_8205);
or U14933 (N_14933,N_5161,N_7524);
nor U14934 (N_14934,N_9643,N_7712);
xnor U14935 (N_14935,N_9968,N_9865);
nand U14936 (N_14936,N_8086,N_9908);
and U14937 (N_14937,N_9164,N_9198);
nor U14938 (N_14938,N_8215,N_8359);
and U14939 (N_14939,N_5230,N_8616);
nand U14940 (N_14940,N_5376,N_5768);
nor U14941 (N_14941,N_8974,N_5584);
or U14942 (N_14942,N_6316,N_7083);
and U14943 (N_14943,N_9334,N_6468);
and U14944 (N_14944,N_7724,N_6568);
and U14945 (N_14945,N_8801,N_6826);
nor U14946 (N_14946,N_5322,N_9419);
and U14947 (N_14947,N_9064,N_8243);
nor U14948 (N_14948,N_8400,N_8579);
or U14949 (N_14949,N_6182,N_9393);
or U14950 (N_14950,N_9737,N_7460);
and U14951 (N_14951,N_5597,N_6452);
nor U14952 (N_14952,N_5145,N_6256);
nand U14953 (N_14953,N_9110,N_9130);
or U14954 (N_14954,N_7326,N_5852);
and U14955 (N_14955,N_6970,N_8756);
nand U14956 (N_14956,N_9163,N_6445);
or U14957 (N_14957,N_5569,N_7579);
nor U14958 (N_14958,N_7875,N_6339);
xnor U14959 (N_14959,N_6377,N_7516);
xor U14960 (N_14960,N_5319,N_9070);
and U14961 (N_14961,N_6079,N_8705);
xor U14962 (N_14962,N_7123,N_6956);
or U14963 (N_14963,N_7345,N_7215);
nor U14964 (N_14964,N_7846,N_9513);
nand U14965 (N_14965,N_5658,N_9608);
and U14966 (N_14966,N_5264,N_8222);
nand U14967 (N_14967,N_8544,N_8418);
and U14968 (N_14968,N_9115,N_6205);
nor U14969 (N_14969,N_9461,N_9871);
nor U14970 (N_14970,N_6553,N_7471);
xnor U14971 (N_14971,N_7181,N_7110);
nand U14972 (N_14972,N_7638,N_9782);
nor U14973 (N_14973,N_7122,N_7404);
nor U14974 (N_14974,N_5583,N_6019);
nor U14975 (N_14975,N_8640,N_6833);
and U14976 (N_14976,N_6802,N_6094);
nand U14977 (N_14977,N_5309,N_7019);
or U14978 (N_14978,N_5538,N_6691);
nor U14979 (N_14979,N_9434,N_5964);
and U14980 (N_14980,N_9552,N_7812);
nand U14981 (N_14981,N_7341,N_8188);
nand U14982 (N_14982,N_7695,N_5999);
nor U14983 (N_14983,N_8232,N_5798);
xor U14984 (N_14984,N_8183,N_9450);
nor U14985 (N_14985,N_9981,N_7827);
nor U14986 (N_14986,N_8076,N_9309);
nand U14987 (N_14987,N_5625,N_7754);
and U14988 (N_14988,N_6775,N_6230);
nor U14989 (N_14989,N_9722,N_7250);
nor U14990 (N_14990,N_6479,N_7352);
or U14991 (N_14991,N_5124,N_5105);
and U14992 (N_14992,N_5813,N_5293);
nand U14993 (N_14993,N_7518,N_5380);
nand U14994 (N_14994,N_7333,N_7495);
or U14995 (N_14995,N_6040,N_8313);
nor U14996 (N_14996,N_7891,N_8130);
nand U14997 (N_14997,N_5814,N_5257);
xnor U14998 (N_14998,N_7202,N_6496);
and U14999 (N_14999,N_9224,N_7510);
xnor UO_0 (O_0,N_12539,N_10425);
xnor UO_1 (O_1,N_13254,N_13912);
xnor UO_2 (O_2,N_12010,N_13512);
xor UO_3 (O_3,N_10415,N_14262);
xnor UO_4 (O_4,N_13853,N_14582);
nor UO_5 (O_5,N_11196,N_14638);
and UO_6 (O_6,N_13202,N_12354);
or UO_7 (O_7,N_12293,N_12860);
nor UO_8 (O_8,N_11963,N_12516);
xnor UO_9 (O_9,N_11943,N_10770);
nor UO_10 (O_10,N_14669,N_13720);
and UO_11 (O_11,N_14910,N_14257);
nor UO_12 (O_12,N_12885,N_13669);
xnor UO_13 (O_13,N_10785,N_14415);
xor UO_14 (O_14,N_13023,N_10499);
and UO_15 (O_15,N_11348,N_12740);
nor UO_16 (O_16,N_12490,N_11947);
xnor UO_17 (O_17,N_10374,N_12323);
xnor UO_18 (O_18,N_10059,N_13580);
or UO_19 (O_19,N_12224,N_14572);
nor UO_20 (O_20,N_12245,N_13192);
xnor UO_21 (O_21,N_11991,N_13726);
or UO_22 (O_22,N_14732,N_11909);
nor UO_23 (O_23,N_10687,N_14026);
nand UO_24 (O_24,N_12544,N_12814);
and UO_25 (O_25,N_12597,N_11336);
nand UO_26 (O_26,N_10962,N_13919);
or UO_27 (O_27,N_14537,N_14567);
nor UO_28 (O_28,N_13969,N_10203);
nor UO_29 (O_29,N_14474,N_13977);
nor UO_30 (O_30,N_10658,N_12165);
nand UO_31 (O_31,N_11685,N_10718);
nand UO_32 (O_32,N_11143,N_13155);
or UO_33 (O_33,N_12441,N_14431);
xnor UO_34 (O_34,N_12664,N_13947);
nand UO_35 (O_35,N_14557,N_13431);
nand UO_36 (O_36,N_13397,N_12784);
nand UO_37 (O_37,N_13160,N_13523);
xor UO_38 (O_38,N_12731,N_12134);
xnor UO_39 (O_39,N_14115,N_10406);
nand UO_40 (O_40,N_13129,N_12983);
or UO_41 (O_41,N_12098,N_13648);
nand UO_42 (O_42,N_10812,N_13266);
xnor UO_43 (O_43,N_14300,N_11037);
xor UO_44 (O_44,N_11571,N_10971);
and UO_45 (O_45,N_13649,N_13894);
nand UO_46 (O_46,N_11334,N_13865);
xor UO_47 (O_47,N_13722,N_14937);
and UO_48 (O_48,N_12581,N_11278);
and UO_49 (O_49,N_10528,N_14734);
nand UO_50 (O_50,N_10503,N_10582);
nor UO_51 (O_51,N_13561,N_10175);
or UO_52 (O_52,N_13609,N_11326);
nor UO_53 (O_53,N_13142,N_14286);
nor UO_54 (O_54,N_12919,N_12495);
and UO_55 (O_55,N_14811,N_11830);
nand UO_56 (O_56,N_13480,N_13634);
or UO_57 (O_57,N_10001,N_11263);
and UO_58 (O_58,N_11740,N_14364);
xor UO_59 (O_59,N_11727,N_14491);
xor UO_60 (O_60,N_10826,N_13372);
or UO_61 (O_61,N_12262,N_14902);
and UO_62 (O_62,N_14563,N_11033);
xor UO_63 (O_63,N_11429,N_13723);
nand UO_64 (O_64,N_13540,N_10608);
and UO_65 (O_65,N_13509,N_13717);
nor UO_66 (O_66,N_10646,N_14195);
or UO_67 (O_67,N_14691,N_10701);
nand UO_68 (O_68,N_14890,N_13219);
nand UO_69 (O_69,N_13315,N_13406);
nor UO_70 (O_70,N_11098,N_10989);
nor UO_71 (O_71,N_10678,N_10730);
xor UO_72 (O_72,N_11205,N_13823);
or UO_73 (O_73,N_14751,N_13873);
nand UO_74 (O_74,N_12431,N_14067);
or UO_75 (O_75,N_14113,N_13670);
nand UO_76 (O_76,N_10549,N_14879);
nand UO_77 (O_77,N_12219,N_11668);
and UO_78 (O_78,N_12788,N_10560);
nor UO_79 (O_79,N_10155,N_14701);
and UO_80 (O_80,N_12990,N_11243);
and UO_81 (O_81,N_13757,N_10916);
nand UO_82 (O_82,N_12179,N_13225);
and UO_83 (O_83,N_13495,N_13205);
nor UO_84 (O_84,N_10859,N_12632);
xnor UO_85 (O_85,N_14769,N_10974);
nand UO_86 (O_86,N_10093,N_13439);
or UO_87 (O_87,N_12153,N_13345);
nand UO_88 (O_88,N_10768,N_11951);
or UO_89 (O_89,N_11523,N_14590);
or UO_90 (O_90,N_11390,N_14965);
nor UO_91 (O_91,N_10869,N_13761);
nand UO_92 (O_92,N_13471,N_10047);
nor UO_93 (O_93,N_12133,N_10171);
or UO_94 (O_94,N_10286,N_12463);
or UO_95 (O_95,N_14361,N_12921);
nor UO_96 (O_96,N_13195,N_11745);
nand UO_97 (O_97,N_11979,N_12160);
or UO_98 (O_98,N_11564,N_10934);
xnor UO_99 (O_99,N_10665,N_12511);
nand UO_100 (O_100,N_13917,N_10275);
xor UO_101 (O_101,N_10553,N_11107);
xnor UO_102 (O_102,N_12774,N_10355);
nor UO_103 (O_103,N_12585,N_14839);
or UO_104 (O_104,N_13404,N_12605);
xor UO_105 (O_105,N_12720,N_11242);
nor UO_106 (O_106,N_13991,N_14551);
or UO_107 (O_107,N_12980,N_11531);
nand UO_108 (O_108,N_12791,N_13945);
xnor UO_109 (O_109,N_14331,N_13908);
nand UO_110 (O_110,N_10961,N_13223);
nand UO_111 (O_111,N_13456,N_11455);
xnor UO_112 (O_112,N_11756,N_13555);
nor UO_113 (O_113,N_13455,N_11366);
nor UO_114 (O_114,N_11709,N_13138);
nand UO_115 (O_115,N_13140,N_14127);
and UO_116 (O_116,N_13828,N_14840);
or UO_117 (O_117,N_10903,N_11015);
and UO_118 (O_118,N_12209,N_10131);
nor UO_119 (O_119,N_11050,N_13855);
nor UO_120 (O_120,N_13748,N_11082);
or UO_121 (O_121,N_14201,N_13256);
and UO_122 (O_122,N_13876,N_12369);
and UO_123 (O_123,N_14939,N_12538);
xor UO_124 (O_124,N_12743,N_13167);
and UO_125 (O_125,N_12096,N_11984);
and UO_126 (O_126,N_12662,N_11898);
or UO_127 (O_127,N_12566,N_13758);
nor UO_128 (O_128,N_13369,N_14072);
xnor UO_129 (O_129,N_13144,N_10757);
and UO_130 (O_130,N_11043,N_13238);
nor UO_131 (O_131,N_11539,N_10284);
and UO_132 (O_132,N_12491,N_13549);
or UO_133 (O_133,N_10241,N_12373);
and UO_134 (O_134,N_13323,N_10583);
nand UO_135 (O_135,N_11781,N_14588);
and UO_136 (O_136,N_12531,N_12271);
nor UO_137 (O_137,N_13856,N_13029);
nor UO_138 (O_138,N_12828,N_14176);
and UO_139 (O_139,N_13714,N_11762);
or UO_140 (O_140,N_10140,N_13652);
nor UO_141 (O_141,N_10009,N_12008);
or UO_142 (O_142,N_10194,N_13162);
nand UO_143 (O_143,N_14509,N_10992);
or UO_144 (O_144,N_13527,N_13172);
xnor UO_145 (O_145,N_12150,N_11081);
or UO_146 (O_146,N_11852,N_12036);
nor UO_147 (O_147,N_12750,N_11777);
nand UO_148 (O_148,N_12830,N_11871);
nand UO_149 (O_149,N_14712,N_13545);
and UO_150 (O_150,N_12767,N_13858);
or UO_151 (O_151,N_13579,N_11642);
or UO_152 (O_152,N_13055,N_13412);
and UO_153 (O_153,N_13115,N_14544);
xnor UO_154 (O_154,N_11617,N_11450);
or UO_155 (O_155,N_13211,N_12813);
nor UO_156 (O_156,N_12418,N_12877);
and UO_157 (O_157,N_10966,N_12685);
nand UO_158 (O_158,N_12532,N_13067);
nand UO_159 (O_159,N_14493,N_14335);
nor UO_160 (O_160,N_13452,N_13534);
or UO_161 (O_161,N_11467,N_14150);
xnor UO_162 (O_162,N_10359,N_11809);
nor UO_163 (O_163,N_10045,N_14314);
xnor UO_164 (O_164,N_14158,N_13065);
nor UO_165 (O_165,N_14741,N_10016);
or UO_166 (O_166,N_10294,N_14786);
nor UO_167 (O_167,N_14155,N_14889);
nand UO_168 (O_168,N_14011,N_13241);
nor UO_169 (O_169,N_12971,N_12005);
and UO_170 (O_170,N_12059,N_12678);
nor UO_171 (O_171,N_10523,N_12782);
xnor UO_172 (O_172,N_14145,N_13571);
xnor UO_173 (O_173,N_14467,N_10682);
and UO_174 (O_174,N_14059,N_10710);
nor UO_175 (O_175,N_11346,N_14355);
xor UO_176 (O_176,N_10711,N_14713);
xor UO_177 (O_177,N_11784,N_14032);
and UO_178 (O_178,N_12831,N_10402);
nor UO_179 (O_179,N_12805,N_13169);
xor UO_180 (O_180,N_12999,N_14773);
nand UO_181 (O_181,N_10790,N_14081);
nor UO_182 (O_182,N_14216,N_11361);
nand UO_183 (O_183,N_10606,N_14546);
or UO_184 (O_184,N_10860,N_10664);
xor UO_185 (O_185,N_13793,N_14800);
xnor UO_186 (O_186,N_12568,N_11847);
and UO_187 (O_187,N_10955,N_12241);
nand UO_188 (O_188,N_13773,N_10732);
nor UO_189 (O_189,N_11799,N_13304);
or UO_190 (O_190,N_13967,N_13262);
xor UO_191 (O_191,N_13885,N_13791);
nor UO_192 (O_192,N_11882,N_13015);
or UO_193 (O_193,N_11733,N_12368);
nor UO_194 (O_194,N_11952,N_13230);
and UO_195 (O_195,N_14193,N_11464);
nor UO_196 (O_196,N_13850,N_10972);
or UO_197 (O_197,N_12304,N_14325);
xor UO_198 (O_198,N_10489,N_12004);
and UO_199 (O_199,N_14141,N_14627);
xnor UO_200 (O_200,N_12291,N_10361);
or UO_201 (O_201,N_12996,N_14337);
nand UO_202 (O_202,N_13951,N_12034);
nor UO_203 (O_203,N_13840,N_10917);
nor UO_204 (O_204,N_11344,N_14687);
and UO_205 (O_205,N_13104,N_14525);
nor UO_206 (O_206,N_11227,N_10628);
xor UO_207 (O_207,N_10685,N_10807);
xnor UO_208 (O_208,N_10931,N_10272);
and UO_209 (O_209,N_13366,N_11404);
nor UO_210 (O_210,N_14256,N_13292);
nand UO_211 (O_211,N_11028,N_10429);
nand UO_212 (O_212,N_10106,N_12487);
and UO_213 (O_213,N_14204,N_11048);
and UO_214 (O_214,N_10126,N_14104);
and UO_215 (O_215,N_11108,N_10833);
or UO_216 (O_216,N_14768,N_11920);
and UO_217 (O_217,N_11794,N_14297);
and UO_218 (O_218,N_13827,N_13498);
nand UO_219 (O_219,N_12902,N_12890);
xor UO_220 (O_220,N_14457,N_13197);
nand UO_221 (O_221,N_12019,N_10067);
and UO_222 (O_222,N_10127,N_10023);
and UO_223 (O_223,N_12534,N_14724);
xor UO_224 (O_224,N_12480,N_13656);
or UO_225 (O_225,N_10576,N_11662);
and UO_226 (O_226,N_11890,N_13039);
and UO_227 (O_227,N_10689,N_14774);
nand UO_228 (O_228,N_10465,N_11282);
nand UO_229 (O_229,N_13923,N_14404);
and UO_230 (O_230,N_11634,N_11510);
xnor UO_231 (O_231,N_12312,N_13389);
xnor UO_232 (O_232,N_13796,N_11965);
nand UO_233 (O_233,N_13764,N_13116);
and UO_234 (O_234,N_10511,N_13124);
nor UO_235 (O_235,N_10236,N_10543);
xor UO_236 (O_236,N_12269,N_10882);
or UO_237 (O_237,N_12922,N_10987);
and UO_238 (O_238,N_13459,N_13227);
xnor UO_239 (O_239,N_11322,N_13267);
and UO_240 (O_240,N_14877,N_13554);
nor UO_241 (O_241,N_13487,N_11454);
or UO_242 (O_242,N_13505,N_14156);
nand UO_243 (O_243,N_10021,N_12176);
nor UO_244 (O_244,N_11097,N_11428);
and UO_245 (O_245,N_13765,N_13121);
nand UO_246 (O_246,N_11257,N_10477);
nor UO_247 (O_247,N_13216,N_12540);
and UO_248 (O_248,N_13595,N_10360);
or UO_249 (O_249,N_11482,N_13000);
nand UO_250 (O_250,N_12763,N_11011);
nand UO_251 (O_251,N_11252,N_11106);
nor UO_252 (O_252,N_11583,N_13653);
nand UO_253 (O_253,N_13598,N_10736);
and UO_254 (O_254,N_13848,N_10592);
xor UO_255 (O_255,N_10868,N_13413);
nor UO_256 (O_256,N_12391,N_10124);
and UO_257 (O_257,N_13678,N_14927);
and UO_258 (O_258,N_14086,N_13302);
or UO_259 (O_259,N_14685,N_10037);
or UO_260 (O_260,N_14911,N_14565);
or UO_261 (O_261,N_10358,N_11000);
nand UO_262 (O_262,N_10423,N_11542);
and UO_263 (O_263,N_10846,N_12970);
or UO_264 (O_264,N_14548,N_11060);
nor UO_265 (O_265,N_12185,N_13259);
and UO_266 (O_266,N_13785,N_14153);
and UO_267 (O_267,N_10110,N_12000);
nor UO_268 (O_268,N_10516,N_14830);
or UO_269 (O_269,N_12332,N_11453);
xor UO_270 (O_270,N_10270,N_14266);
nor UO_271 (O_271,N_11451,N_12497);
nor UO_272 (O_272,N_10788,N_12546);
xor UO_273 (O_273,N_10453,N_10419);
or UO_274 (O_274,N_14705,N_12212);
nor UO_275 (O_275,N_12721,N_12189);
or UO_276 (O_276,N_13157,N_13043);
or UO_277 (O_277,N_11371,N_14182);
and UO_278 (O_278,N_14425,N_13616);
nand UO_279 (O_279,N_14370,N_12693);
xor UO_280 (O_280,N_14663,N_10836);
or UO_281 (O_281,N_13644,N_11174);
nor UO_282 (O_282,N_12178,N_10483);
nor UO_283 (O_283,N_11760,N_12633);
or UO_284 (O_284,N_14143,N_13994);
and UO_285 (O_285,N_14674,N_13910);
nor UO_286 (O_286,N_11981,N_11912);
xor UO_287 (O_287,N_13407,N_11360);
and UO_288 (O_288,N_10815,N_11658);
nor UO_289 (O_289,N_13575,N_13798);
or UO_290 (O_290,N_11591,N_12327);
xor UO_291 (O_291,N_10324,N_12865);
nand UO_292 (O_292,N_13953,N_14717);
xor UO_293 (O_293,N_11300,N_10211);
nand UO_294 (O_294,N_10558,N_13154);
and UO_295 (O_295,N_12954,N_14043);
nor UO_296 (O_296,N_11526,N_12726);
or UO_297 (O_297,N_13012,N_14432);
and UO_298 (O_298,N_14673,N_11166);
nand UO_299 (O_299,N_14186,N_14842);
and UO_300 (O_300,N_10493,N_14244);
xor UO_301 (O_301,N_14538,N_13935);
or UO_302 (O_302,N_12553,N_10574);
nor UO_303 (O_303,N_14715,N_11054);
nand UO_304 (O_304,N_14988,N_11163);
and UO_305 (O_305,N_10748,N_10417);
and UO_306 (O_306,N_14004,N_14387);
and UO_307 (O_307,N_12085,N_10052);
or UO_308 (O_308,N_11316,N_11665);
and UO_309 (O_309,N_12635,N_11609);
xor UO_310 (O_310,N_10262,N_10876);
and UO_311 (O_311,N_10670,N_10497);
or UO_312 (O_312,N_14392,N_10967);
xnor UO_313 (O_313,N_12582,N_10615);
nand UO_314 (O_314,N_12547,N_12968);
nand UO_315 (O_315,N_14992,N_11397);
xnor UO_316 (O_316,N_12131,N_11115);
xnor UO_317 (O_317,N_12058,N_10285);
nand UO_318 (O_318,N_11815,N_14154);
or UO_319 (O_319,N_14313,N_11647);
and UO_320 (O_320,N_14429,N_10180);
nand UO_321 (O_321,N_14063,N_12002);
and UO_322 (O_322,N_14307,N_12158);
nor UO_323 (O_323,N_10669,N_13287);
and UO_324 (O_324,N_14273,N_10264);
nand UO_325 (O_325,N_11832,N_12783);
nand UO_326 (O_326,N_10344,N_10901);
xor UO_327 (O_327,N_14731,N_12408);
nand UO_328 (O_328,N_13221,N_13989);
and UO_329 (O_329,N_12173,N_11051);
and UO_330 (O_330,N_12742,N_12929);
or UO_331 (O_331,N_10986,N_13332);
nand UO_332 (O_332,N_14486,N_14192);
or UO_333 (O_333,N_11804,N_10808);
and UO_334 (O_334,N_12233,N_10518);
and UO_335 (O_335,N_13863,N_13640);
nor UO_336 (O_336,N_10874,N_12437);
or UO_337 (O_337,N_12851,N_10572);
xor UO_338 (O_338,N_10829,N_13081);
nor UO_339 (O_339,N_14519,N_10793);
xnor UO_340 (O_340,N_11798,N_13544);
nor UO_341 (O_341,N_12659,N_10214);
and UO_342 (O_342,N_11931,N_14900);
xor UO_343 (O_343,N_14242,N_12677);
or UO_344 (O_344,N_13775,N_12526);
nor UO_345 (O_345,N_11442,N_14978);
and UO_346 (O_346,N_11905,N_12840);
and UO_347 (O_347,N_13447,N_14743);
nand UO_348 (O_348,N_12350,N_12389);
or UO_349 (O_349,N_11565,N_12223);
xor UO_350 (O_350,N_13478,N_14821);
nand UO_351 (O_351,N_12956,N_12683);
nand UO_352 (O_352,N_13474,N_10291);
nand UO_353 (O_353,N_12045,N_13668);
xor UO_354 (O_354,N_10357,N_13422);
or UO_355 (O_355,N_14570,N_10050);
or UO_356 (O_356,N_12658,N_12939);
and UO_357 (O_357,N_11739,N_13106);
nor UO_358 (O_358,N_13054,N_12386);
or UO_359 (O_359,N_11992,N_12292);
and UO_360 (O_360,N_10196,N_11114);
nand UO_361 (O_361,N_13747,N_12679);
xor UO_362 (O_362,N_14865,N_10157);
nor UO_363 (O_363,N_12355,N_14826);
nand UO_364 (O_364,N_11047,N_12681);
nor UO_365 (O_365,N_10899,N_10176);
and UO_366 (O_366,N_12289,N_13318);
nor UO_367 (O_367,N_13751,N_11836);
xor UO_368 (O_368,N_10708,N_10662);
nor UO_369 (O_369,N_10648,N_11006);
xnor UO_370 (O_370,N_10130,N_13606);
or UO_371 (O_371,N_10227,N_10030);
or UO_372 (O_372,N_10134,N_12103);
and UO_373 (O_373,N_12232,N_14250);
or UO_374 (O_374,N_13260,N_11228);
and UO_375 (O_375,N_12716,N_13263);
nor UO_376 (O_376,N_14147,N_12148);
and UO_377 (O_377,N_11825,N_14569);
or UO_378 (O_378,N_13299,N_10950);
nand UO_379 (O_379,N_12994,N_12957);
nor UO_380 (O_380,N_11751,N_12594);
xor UO_381 (O_381,N_11528,N_12878);
nor UO_382 (O_382,N_11408,N_11874);
xor UO_383 (O_383,N_12772,N_12626);
or UO_384 (O_384,N_11562,N_12348);
and UO_385 (O_385,N_14989,N_14146);
xnor UO_386 (O_386,N_14936,N_11008);
nand UO_387 (O_387,N_11925,N_12573);
and UO_388 (O_388,N_14012,N_11295);
nor UO_389 (O_389,N_14274,N_14872);
or UO_390 (O_390,N_12338,N_11239);
nand UO_391 (O_391,N_13641,N_14219);
or UO_392 (O_392,N_12567,N_12443);
and UO_393 (O_393,N_13188,N_13822);
nand UO_394 (O_394,N_12069,N_13377);
and UO_395 (O_395,N_11650,N_10132);
and UO_396 (O_396,N_13305,N_10635);
or UO_397 (O_397,N_10340,N_11970);
nor UO_398 (O_398,N_10173,N_12607);
nand UO_399 (O_399,N_12151,N_10542);
nand UO_400 (O_400,N_14948,N_13792);
nand UO_401 (O_401,N_11085,N_10006);
and UO_402 (O_402,N_13661,N_13731);
nand UO_403 (O_403,N_10936,N_13343);
or UO_404 (O_404,N_14915,N_10526);
nor UO_405 (O_405,N_14048,N_10496);
and UO_406 (O_406,N_13118,N_12610);
xor UO_407 (O_407,N_11119,N_10000);
and UO_408 (O_408,N_14535,N_13985);
xor UO_409 (O_409,N_12834,N_14133);
xor UO_410 (O_410,N_13165,N_12230);
or UO_411 (O_411,N_13420,N_11413);
xor UO_412 (O_412,N_10775,N_12125);
nor UO_413 (O_413,N_11285,N_13907);
or UO_414 (O_414,N_14479,N_10512);
nor UO_415 (O_415,N_11962,N_10424);
and UO_416 (O_416,N_11645,N_14152);
xnor UO_417 (O_417,N_11335,N_10276);
or UO_418 (O_418,N_14844,N_14088);
xor UO_419 (O_419,N_12116,N_11613);
or UO_420 (O_420,N_11619,N_11863);
or UO_421 (O_421,N_12712,N_11864);
nand UO_422 (O_422,N_14946,N_11463);
xor UO_423 (O_423,N_11381,N_13161);
and UO_424 (O_424,N_11140,N_14407);
and UO_425 (O_425,N_10305,N_12548);
or UO_426 (O_426,N_11374,N_12175);
and UO_427 (O_427,N_13100,N_13125);
xnor UO_428 (O_428,N_11367,N_14453);
or UO_429 (O_429,N_12274,N_13373);
and UO_430 (O_430,N_11469,N_14738);
nor UO_431 (O_431,N_10347,N_11975);
nor UO_432 (O_432,N_10842,N_13166);
nor UO_433 (O_433,N_14103,N_14390);
xor UO_434 (O_434,N_13470,N_13303);
and UO_435 (O_435,N_12517,N_11724);
nor UO_436 (O_436,N_13780,N_11059);
and UO_437 (O_437,N_13603,N_10022);
and UO_438 (O_438,N_13484,N_13007);
xor UO_439 (O_439,N_12222,N_10098);
or UO_440 (O_440,N_14697,N_12231);
or UO_441 (O_441,N_12667,N_14166);
or UO_442 (O_442,N_11176,N_10018);
nor UO_443 (O_443,N_12401,N_10265);
nor UO_444 (O_444,N_13079,N_14629);
or UO_445 (O_445,N_12663,N_13918);
and UO_446 (O_446,N_13813,N_14973);
xnor UO_447 (O_447,N_10521,N_12628);
or UO_448 (O_448,N_13326,N_13082);
nand UO_449 (O_449,N_12471,N_13849);
and UO_450 (O_450,N_14688,N_10271);
xor UO_451 (O_451,N_10554,N_11556);
or UO_452 (O_452,N_10591,N_14498);
or UO_453 (O_453,N_10088,N_13027);
or UO_454 (O_454,N_10816,N_14510);
xor UO_455 (O_455,N_10259,N_11330);
xnor UO_456 (O_456,N_12780,N_12916);
nand UO_457 (O_457,N_10181,N_12604);
and UO_458 (O_458,N_13298,N_12188);
xnor UO_459 (O_459,N_10599,N_12102);
nand UO_460 (O_460,N_13390,N_14600);
xor UO_461 (O_461,N_13837,N_10680);
and UO_462 (O_462,N_11741,N_12670);
nand UO_463 (O_463,N_10529,N_13537);
or UO_464 (O_464,N_13683,N_14210);
nand UO_465 (O_465,N_14601,N_13997);
nand UO_466 (O_466,N_14234,N_10224);
nand UO_467 (O_467,N_13701,N_13122);
nand UO_468 (O_468,N_11587,N_11862);
nor UO_469 (O_469,N_10172,N_11950);
and UO_470 (O_470,N_13570,N_14980);
nand UO_471 (O_471,N_12768,N_14477);
or UO_472 (O_472,N_12328,N_11160);
nor UO_473 (O_473,N_10300,N_11811);
or UO_474 (O_474,N_12887,N_14740);
nand UO_475 (O_475,N_11299,N_13525);
nand UO_476 (O_476,N_10811,N_11405);
nor UO_477 (O_477,N_10197,N_11250);
nor UO_478 (O_478,N_14709,N_13199);
and UO_479 (O_479,N_14982,N_13429);
or UO_480 (O_480,N_14670,N_13972);
or UO_481 (O_481,N_12524,N_11091);
nor UO_482 (O_482,N_13386,N_12859);
or UO_483 (O_483,N_10908,N_10650);
nor UO_484 (O_484,N_12697,N_10527);
nor UO_485 (O_485,N_14446,N_12962);
nor UO_486 (O_486,N_14276,N_13882);
or UO_487 (O_487,N_14620,N_11262);
xor UO_488 (O_488,N_13690,N_12550);
and UO_489 (O_489,N_10354,N_11456);
and UO_490 (O_490,N_14135,N_12060);
xor UO_491 (O_491,N_11823,N_14753);
nor UO_492 (O_492,N_11235,N_12079);
xnor UO_493 (O_493,N_12329,N_13767);
nand UO_494 (O_494,N_12948,N_13803);
nor UO_495 (O_495,N_13463,N_10484);
or UO_496 (O_496,N_13024,N_11310);
or UO_497 (O_497,N_10422,N_14173);
or UO_498 (O_498,N_14287,N_10947);
and UO_499 (O_499,N_14892,N_11080);
nor UO_500 (O_500,N_14861,N_14016);
or UO_501 (O_501,N_14635,N_11099);
xor UO_502 (O_502,N_13589,N_10267);
nand UO_503 (O_503,N_10647,N_14875);
nand UO_504 (O_504,N_14211,N_11723);
nor UO_505 (O_505,N_12115,N_11324);
or UO_506 (O_506,N_12884,N_14969);
nand UO_507 (O_507,N_13280,N_13719);
or UO_508 (O_508,N_14666,N_10613);
xor UO_509 (O_509,N_12218,N_13890);
nand UO_510 (O_510,N_13153,N_11796);
xnor UO_511 (O_511,N_10299,N_13394);
and UO_512 (O_512,N_14924,N_12300);
nand UO_513 (O_513,N_11072,N_10996);
xor UO_514 (O_514,N_14267,N_14652);
or UO_515 (O_515,N_12513,N_10912);
or UO_516 (O_516,N_10228,N_13272);
nand UO_517 (O_517,N_11768,N_11093);
or UO_518 (O_518,N_13031,N_10724);
and UO_519 (O_519,N_12871,N_14227);
or UO_520 (O_520,N_14799,N_13902);
nor UO_521 (O_521,N_10199,N_10438);
nand UO_522 (O_522,N_10261,N_11261);
or UO_523 (O_523,N_13312,N_13421);
xor UO_524 (O_524,N_11158,N_14531);
nor UO_525 (O_525,N_14472,N_11786);
nand UO_526 (O_526,N_11365,N_12704);
and UO_527 (O_527,N_10924,N_13307);
or UO_528 (O_528,N_12904,N_13679);
xnor UO_529 (O_529,N_14634,N_13092);
nor UO_530 (O_530,N_11031,N_14802);
nor UO_531 (O_531,N_11449,N_12623);
nand UO_532 (O_532,N_13949,N_11661);
nand UO_533 (O_533,N_14792,N_12326);
xor UO_534 (O_534,N_10301,N_13869);
and UO_535 (O_535,N_12192,N_14918);
and UO_536 (O_536,N_14541,N_10304);
and UO_537 (O_537,N_11287,N_10941);
nor UO_538 (O_538,N_12282,N_14630);
xor UO_539 (O_539,N_10169,N_10195);
xor UO_540 (O_540,N_13826,N_11507);
or UO_541 (O_541,N_13419,N_13105);
nor UO_542 (O_542,N_11924,N_10764);
or UO_543 (O_543,N_12808,N_12883);
or UO_544 (O_544,N_12769,N_12062);
or UO_545 (O_545,N_12512,N_12022);
and UO_546 (O_546,N_13879,N_14396);
or UO_547 (O_547,N_14109,N_11218);
or UO_548 (O_548,N_14232,N_12816);
and UO_549 (O_549,N_14851,N_11121);
and UO_550 (O_550,N_10885,N_10010);
xnor UO_551 (O_551,N_10803,N_11308);
or UO_552 (O_552,N_11671,N_11581);
and UO_553 (O_553,N_11315,N_10626);
or UO_554 (O_554,N_12199,N_13513);
or UO_555 (O_555,N_13235,N_13996);
nand UO_556 (O_556,N_14850,N_14695);
nand UO_557 (O_557,N_13770,N_10209);
xnor UO_558 (O_558,N_13786,N_13592);
nand UO_559 (O_559,N_14694,N_11364);
nor UO_560 (O_560,N_11648,N_10937);
and UO_561 (O_561,N_11549,N_10392);
or UO_562 (O_562,N_12770,N_10729);
nor UO_563 (O_563,N_11069,N_13095);
and UO_564 (O_564,N_13415,N_11204);
nand UO_565 (O_565,N_13176,N_14766);
nor UO_566 (O_566,N_13638,N_13884);
or UO_567 (O_567,N_13026,N_12457);
xnor UO_568 (O_568,N_11104,N_14021);
nand UO_569 (O_569,N_12063,N_14029);
xnor UO_570 (O_570,N_12964,N_10125);
or UO_571 (O_571,N_14595,N_14386);
or UO_572 (O_572,N_11624,N_11268);
xor UO_573 (O_573,N_12592,N_13712);
nand UO_574 (O_574,N_14755,N_12759);
and UO_575 (O_575,N_13437,N_11949);
and UO_576 (O_576,N_11168,N_14101);
or UO_577 (O_577,N_11370,N_11424);
nor UO_578 (O_578,N_13428,N_14343);
nor UO_579 (O_579,N_11873,N_11625);
nor UO_580 (O_580,N_11976,N_13763);
xor UO_581 (O_581,N_11164,N_13276);
and UO_582 (O_582,N_13839,N_13915);
nand UO_583 (O_583,N_11638,N_14416);
and UO_584 (O_584,N_10540,N_11972);
xor UO_585 (O_585,N_12213,N_13030);
nor UO_586 (O_586,N_12593,N_11563);
and UO_587 (O_587,N_11802,N_10587);
xor UO_588 (O_588,N_14761,N_10544);
xor UO_589 (O_589,N_14061,N_10025);
or UO_590 (O_590,N_14323,N_12779);
xor UO_591 (O_591,N_14255,N_11078);
xor UO_592 (O_592,N_13357,N_14986);
nor UO_593 (O_593,N_14448,N_10982);
xor UO_594 (O_594,N_12114,N_11032);
and UO_595 (O_595,N_10019,N_12198);
and UO_596 (O_596,N_11731,N_12479);
or UO_597 (O_597,N_11684,N_12372);
and UO_598 (O_598,N_11659,N_13499);
xnor UO_599 (O_599,N_14348,N_14105);
nor UO_600 (O_600,N_14882,N_10975);
nand UO_601 (O_601,N_12376,N_14735);
nand UO_602 (O_602,N_13599,N_11846);
nand UO_603 (O_603,N_13133,N_10500);
nand UO_604 (O_604,N_13718,N_11214);
nor UO_605 (O_605,N_14793,N_12317);
or UO_606 (O_606,N_13231,N_13939);
xor UO_607 (O_607,N_14347,N_10935);
and UO_608 (O_608,N_13604,N_12162);
or UO_609 (O_609,N_14598,N_10221);
or UO_610 (O_610,N_14483,N_11894);
nor UO_611 (O_611,N_13355,N_12451);
xor UO_612 (O_612,N_10129,N_11736);
nor UO_613 (O_613,N_12319,N_13435);
nand UO_614 (O_614,N_14249,N_13245);
xor UO_615 (O_615,N_14475,N_13284);
nand UO_616 (O_616,N_10238,N_14552);
nor UO_617 (O_617,N_11036,N_13306);
and UO_618 (O_618,N_12618,N_12107);
nand UO_619 (O_619,N_14490,N_11907);
and UO_620 (O_620,N_11394,N_12747);
or UO_621 (O_621,N_13132,N_13063);
nor UO_622 (O_622,N_12986,N_10420);
nand UO_623 (O_623,N_14804,N_14955);
xnor UO_624 (O_624,N_13817,N_14665);
and UO_625 (O_625,N_12021,N_14095);
xnor UO_626 (O_626,N_11900,N_11915);
or UO_627 (O_627,N_11485,N_10747);
xnor UO_628 (O_628,N_13721,N_11154);
nand UO_629 (O_629,N_11416,N_14898);
xnor UO_630 (O_630,N_11459,N_14116);
nor UO_631 (O_631,N_11987,N_13959);
nor UO_632 (O_632,N_13033,N_12024);
xor UO_633 (O_633,N_11660,N_14828);
nor UO_634 (O_634,N_13584,N_10721);
or UO_635 (O_635,N_12313,N_12577);
and UO_636 (O_636,N_13164,N_10752);
and UO_637 (O_637,N_14338,N_12033);
nand UO_638 (O_638,N_12729,N_12384);
or UO_639 (O_639,N_13253,N_12172);
nand UO_640 (O_640,N_14863,N_14742);
or UO_641 (O_641,N_14923,N_14046);
and UO_642 (O_642,N_13964,N_14646);
xnor UO_643 (O_643,N_12932,N_11329);
nor UO_644 (O_644,N_12208,N_12803);
nand UO_645 (O_645,N_13834,N_11116);
xnor UO_646 (O_646,N_13654,N_10517);
and UO_647 (O_647,N_13271,N_12843);
and UO_648 (O_648,N_14106,N_14438);
nand UO_649 (O_649,N_11603,N_11669);
and UO_650 (O_650,N_11708,N_10765);
nand UO_651 (O_651,N_10893,N_13096);
or UO_652 (O_652,N_12735,N_10642);
and UO_653 (O_653,N_10911,N_13136);
nand UO_654 (O_654,N_13466,N_14958);
or UO_655 (O_655,N_12489,N_14178);
nor UO_656 (O_656,N_10843,N_10866);
or UO_657 (O_657,N_14699,N_10979);
xor UO_658 (O_658,N_11246,N_10008);
or UO_659 (O_659,N_11680,N_12616);
nor UO_660 (O_660,N_10923,N_11133);
nand UO_661 (O_661,N_13152,N_10679);
nor UO_662 (O_662,N_13725,N_14311);
nor UO_663 (O_663,N_12421,N_10352);
xnor UO_664 (O_664,N_14995,N_11180);
nand UO_665 (O_665,N_14422,N_11994);
nor UO_666 (O_666,N_10806,N_13094);
xnor UO_667 (O_667,N_12417,N_11582);
xnor UO_668 (O_668,N_12995,N_13944);
nand UO_669 (O_669,N_11961,N_13832);
and UO_670 (O_670,N_13028,N_11753);
xnor UO_671 (O_671,N_13625,N_14456);
or UO_672 (O_672,N_10005,N_10498);
xor UO_673 (O_673,N_10174,N_11935);
and UO_674 (O_674,N_14703,N_13035);
and UO_675 (O_675,N_11586,N_10993);
and UO_676 (O_676,N_14945,N_11129);
nor UO_677 (O_677,N_13517,N_12882);
nand UO_678 (O_678,N_13936,N_13900);
and UO_679 (O_679,N_11123,N_11229);
nor UO_680 (O_680,N_10588,N_10178);
xnor UO_681 (O_681,N_12100,N_10248);
or UO_682 (O_682,N_10190,N_13017);
and UO_683 (O_683,N_14677,N_14661);
xnor UO_684 (O_684,N_10389,N_11593);
and UO_685 (O_685,N_10160,N_11363);
nor UO_686 (O_686,N_14881,N_11899);
nor UO_687 (O_687,N_10492,N_13085);
nor UO_688 (O_688,N_12599,N_12456);
nand UO_689 (O_689,N_12675,N_11435);
nor UO_690 (O_690,N_14217,N_10753);
and UO_691 (O_691,N_13203,N_14702);
nand UO_692 (O_692,N_10257,N_14928);
or UO_693 (O_693,N_14938,N_12316);
and UO_694 (O_694,N_13821,N_12752);
and UO_695 (O_695,N_12164,N_10437);
and UO_696 (O_696,N_13034,N_11842);
and UO_697 (O_697,N_13460,N_13859);
and UO_698 (O_698,N_14649,N_12089);
nand UO_699 (O_699,N_12765,N_13815);
nand UO_700 (O_700,N_13185,N_13388);
and UO_701 (O_701,N_10504,N_11530);
and UO_702 (O_702,N_12627,N_13131);
xor UO_703 (O_703,N_13209,N_10886);
nand UO_704 (O_704,N_14042,N_11199);
nor UO_705 (O_705,N_11157,N_13117);
and UO_706 (O_706,N_10036,N_14324);
nand UO_707 (O_707,N_10601,N_14962);
nand UO_708 (O_708,N_13285,N_14129);
and UO_709 (O_709,N_14207,N_11610);
xor UO_710 (O_710,N_10434,N_12093);
nor UO_711 (O_711,N_13633,N_14991);
and UO_712 (O_712,N_12400,N_10015);
or UO_713 (O_713,N_13728,N_10137);
nor UO_714 (O_714,N_13800,N_10692);
and UO_715 (O_715,N_10457,N_11957);
and UO_716 (O_716,N_11495,N_12006);
xnor UO_717 (O_717,N_14527,N_10920);
and UO_718 (O_718,N_10433,N_14420);
and UO_719 (O_719,N_14489,N_12026);
nand UO_720 (O_720,N_10328,N_11734);
or UO_721 (O_721,N_11923,N_10334);
xor UO_722 (O_722,N_10915,N_12787);
and UO_723 (O_723,N_14071,N_14612);
and UO_724 (O_724,N_14533,N_10713);
or UO_725 (O_725,N_14841,N_11850);
xnor UO_726 (O_726,N_13593,N_14760);
and UO_727 (O_727,N_12724,N_12436);
and UO_728 (O_728,N_10318,N_10474);
or UO_729 (O_729,N_13926,N_10439);
and UO_730 (O_730,N_11457,N_13619);
xnor UO_731 (O_731,N_10990,N_12419);
nor UO_732 (O_732,N_12477,N_10268);
xor UO_733 (O_733,N_13675,N_13296);
nor UO_734 (O_734,N_11990,N_13261);
nor UO_735 (O_735,N_10659,N_12937);
and UO_736 (O_736,N_11525,N_14611);
or UO_737 (O_737,N_14970,N_10607);
nor UO_738 (O_738,N_14024,N_13494);
nor UO_739 (O_739,N_14259,N_14499);
and UO_740 (O_740,N_12433,N_14684);
nand UO_741 (O_741,N_12702,N_14680);
and UO_742 (O_742,N_14414,N_11679);
nor UO_743 (O_743,N_11128,N_11267);
xor UO_744 (O_744,N_11234,N_13635);
xnor UO_745 (O_745,N_14066,N_14121);
nand UO_746 (O_746,N_13680,N_13819);
or UO_747 (O_747,N_11226,N_12672);
or UO_748 (O_748,N_11146,N_13752);
and UO_749 (O_749,N_13073,N_12833);
nor UO_750 (O_750,N_12118,N_12701);
or UO_751 (O_751,N_10720,N_12365);
xor UO_752 (O_752,N_11732,N_10705);
or UO_753 (O_753,N_11656,N_10258);
and UO_754 (O_754,N_13289,N_14080);
nor UO_755 (O_755,N_13614,N_11458);
xnor UO_756 (O_756,N_12446,N_10951);
nor UO_757 (O_757,N_12362,N_11189);
nand UO_758 (O_758,N_12298,N_11182);
nand UO_759 (O_759,N_12556,N_11269);
nor UO_760 (O_760,N_10017,N_13732);
and UO_761 (O_761,N_13783,N_13349);
and UO_762 (O_762,N_13204,N_12737);
or UO_763 (O_763,N_12204,N_14780);
xnor UO_764 (O_764,N_11718,N_10421);
or UO_765 (O_765,N_13196,N_12306);
and UO_766 (O_766,N_12154,N_10085);
nand UO_767 (O_767,N_10569,N_14727);
xor UO_768 (O_768,N_13414,N_10397);
nor UO_769 (O_769,N_14511,N_11946);
or UO_770 (O_770,N_13006,N_14465);
nor UO_771 (O_771,N_12650,N_14302);
xor UO_772 (O_772,N_10311,N_14532);
xor UO_773 (O_773,N_12819,N_14679);
nor UO_774 (O_774,N_14454,N_12571);
or UO_775 (O_775,N_13341,N_12719);
and UO_776 (O_776,N_13110,N_14831);
xnor UO_777 (O_777,N_10123,N_12357);
or UO_778 (O_778,N_11693,N_12829);
nand UO_779 (O_779,N_14704,N_10156);
nor UO_780 (O_780,N_13802,N_13961);
nor UO_781 (O_781,N_13448,N_13149);
nor UO_782 (O_782,N_12307,N_10135);
xnor UO_783 (O_783,N_11838,N_10063);
or UO_784 (O_784,N_11996,N_12434);
xor UO_785 (O_785,N_11328,N_10725);
xnor UO_786 (O_786,N_12958,N_11159);
and UO_787 (O_787,N_11673,N_10168);
or UO_788 (O_788,N_11908,N_11219);
nor UO_789 (O_789,N_11145,N_14808);
and UO_790 (O_790,N_10351,N_12947);
nor UO_791 (O_791,N_12799,N_12159);
and UO_792 (O_792,N_12170,N_12047);
or UO_793 (O_793,N_13548,N_11238);
xnor UO_794 (O_794,N_10675,N_12612);
xor UO_795 (O_795,N_14340,N_12560);
xor UO_796 (O_796,N_13632,N_12206);
or UO_797 (O_797,N_14540,N_10373);
and UO_798 (O_798,N_12268,N_11698);
nor UO_799 (O_799,N_11780,N_13268);
nand UO_800 (O_800,N_12344,N_13806);
nor UO_801 (O_801,N_13171,N_10827);
nand UO_802 (O_802,N_10887,N_14874);
nand UO_803 (O_803,N_12920,N_10703);
xor UO_804 (O_804,N_12341,N_13992);
or UO_805 (O_805,N_10296,N_14746);
and UO_806 (O_806,N_13941,N_12267);
and UO_807 (O_807,N_12643,N_14480);
nand UO_808 (O_808,N_14450,N_12478);
and UO_809 (O_809,N_14399,N_10714);
nor UO_810 (O_810,N_10003,N_10479);
nor UO_811 (O_811,N_12126,N_14794);
xnor UO_812 (O_812,N_12012,N_10309);
nand UO_813 (O_813,N_11695,N_11643);
and UO_814 (O_814,N_10462,N_11806);
or UO_815 (O_815,N_14035,N_11904);
or UO_816 (O_816,N_10159,N_10077);
nand UO_817 (O_817,N_13955,N_13739);
xor UO_818 (O_818,N_11694,N_14658);
xor UO_819 (O_819,N_12309,N_13344);
nand UO_820 (O_820,N_14609,N_12445);
and UO_821 (O_821,N_11019,N_14140);
or UO_822 (O_822,N_10191,N_11061);
nor UO_823 (O_823,N_11604,N_14442);
and UO_824 (O_824,N_12924,N_14094);
and UO_825 (O_825,N_14864,N_11848);
nand UO_826 (O_826,N_11588,N_12998);
and UO_827 (O_827,N_14577,N_10871);
nand UO_828 (O_828,N_10146,N_11029);
and UO_829 (O_829,N_13514,N_14838);
and UO_830 (O_830,N_11480,N_10573);
and UO_831 (O_831,N_11602,N_14607);
nor UO_832 (O_832,N_14228,N_10201);
nand UO_833 (O_833,N_12129,N_11743);
and UO_834 (O_834,N_11052,N_12917);
or UO_835 (O_835,N_13655,N_11274);
nand UO_836 (O_836,N_13846,N_12074);
and UO_837 (O_837,N_12333,N_14006);
nand UO_838 (O_838,N_10820,N_11558);
xor UO_839 (O_839,N_12070,N_10095);
nor UO_840 (O_840,N_14064,N_13328);
nand UO_841 (O_841,N_12943,N_10288);
xor UO_842 (O_842,N_10364,N_12798);
nor UO_843 (O_843,N_14051,N_13867);
or UO_844 (O_844,N_10107,N_13948);
or UO_845 (O_845,N_13218,N_12554);
xnor UO_846 (O_846,N_11297,N_12242);
and UO_847 (O_847,N_11005,N_13531);
and UO_848 (O_848,N_13968,N_10282);
nor UO_849 (O_849,N_13727,N_13168);
or UO_850 (O_850,N_11776,N_13922);
nor UO_851 (O_851,N_12235,N_14099);
and UO_852 (O_852,N_10447,N_11758);
nor UO_853 (O_853,N_12700,N_13522);
nor UO_854 (O_854,N_13768,N_11677);
xnor UO_855 (O_855,N_10167,N_12310);
nor UO_856 (O_856,N_10323,N_10452);
nor UO_857 (O_857,N_14504,N_11441);
or UO_858 (O_858,N_13288,N_10672);
nand UO_859 (O_859,N_14585,N_14587);
xor UO_860 (O_860,N_11313,N_11200);
and UO_861 (O_861,N_13182,N_14357);
xor UO_862 (O_862,N_14798,N_12536);
nor UO_863 (O_863,N_10823,N_12285);
or UO_864 (O_864,N_12197,N_13249);
and UO_865 (O_865,N_11291,N_14065);
or UO_866 (O_866,N_10368,N_13493);
nor UO_867 (O_867,N_12161,N_12264);
nand UO_868 (O_868,N_13685,N_10550);
nor UO_869 (O_869,N_11529,N_12493);
and UO_870 (O_870,N_14640,N_10247);
nand UO_871 (O_871,N_11771,N_13676);
xor UO_872 (O_872,N_10577,N_12521);
nand UO_873 (O_873,N_14443,N_13542);
or UO_874 (O_874,N_10464,N_11775);
and UO_875 (O_875,N_11594,N_12911);
or UO_876 (O_876,N_14860,N_10004);
and UO_877 (O_877,N_10217,N_13984);
and UO_878 (O_878,N_14516,N_14956);
or UO_879 (O_879,N_12790,N_12515);
xnor UO_880 (O_880,N_12710,N_11255);
and UO_881 (O_881,N_12589,N_11521);
nor UO_882 (O_882,N_10799,N_12869);
nand UO_883 (O_883,N_10777,N_14764);
and UO_884 (O_884,N_10824,N_11432);
nand UO_885 (O_885,N_12541,N_13931);
and UO_886 (O_886,N_13405,N_10609);
and UO_887 (O_887,N_10163,N_14225);
xnor UO_888 (O_888,N_13921,N_12163);
or UO_889 (O_889,N_14981,N_11552);
xor UO_890 (O_890,N_13340,N_13481);
xor UO_891 (O_891,N_12686,N_11244);
xnor UO_892 (O_892,N_11465,N_12504);
and UO_893 (O_893,N_14941,N_12127);
or UO_894 (O_894,N_10400,N_12844);
and UO_895 (O_895,N_14824,N_10548);
or UO_896 (O_896,N_14326,N_10330);
and UO_897 (O_897,N_14790,N_11020);
nor UO_898 (O_898,N_14885,N_12506);
nand UO_899 (O_899,N_14384,N_10013);
or UO_900 (O_900,N_11822,N_10772);
nand UO_901 (O_901,N_10973,N_14076);
xor UO_902 (O_902,N_12817,N_13611);
nor UO_903 (O_903,N_14151,N_12243);
xor UO_904 (O_904,N_10256,N_12343);
xnor UO_905 (O_905,N_14628,N_12751);
nand UO_906 (O_906,N_11839,N_14819);
nor UO_907 (O_907,N_10333,N_13060);
or UO_908 (O_908,N_14632,N_12933);
nor UO_909 (O_909,N_12621,N_13352);
nor UO_910 (O_910,N_10918,N_14082);
and UO_911 (O_911,N_14690,N_14169);
nand UO_912 (O_912,N_11017,N_13938);
nor UO_913 (O_913,N_11755,N_10319);
or UO_914 (O_914,N_10865,N_14395);
nor UO_915 (O_915,N_12037,N_13430);
xnor UO_916 (O_916,N_14179,N_12804);
nor UO_917 (O_917,N_11837,N_10476);
or UO_918 (O_918,N_13620,N_11075);
xor UO_919 (O_919,N_14818,N_10653);
nor UO_920 (O_920,N_11653,N_13971);
nor UO_921 (O_921,N_10712,N_14079);
nand UO_922 (O_922,N_10964,N_14678);
nor UO_923 (O_923,N_11113,N_13385);
and UO_924 (O_924,N_10501,N_12614);
xor UO_925 (O_925,N_10058,N_12396);
or UO_926 (O_926,N_10939,N_14767);
and UO_927 (O_927,N_11151,N_11260);
nor UO_928 (O_928,N_13558,N_14241);
and UO_929 (O_929,N_11845,N_10317);
and UO_930 (O_930,N_10467,N_13191);
nand UO_931 (O_931,N_13594,N_11461);
or UO_932 (O_932,N_10468,N_12866);
or UO_933 (O_933,N_13424,N_12657);
nor UO_934 (O_934,N_13313,N_12174);
xor UO_935 (O_935,N_10789,N_13179);
nand UO_936 (O_936,N_10922,N_10778);
and UO_937 (O_937,N_10605,N_12893);
nand UO_938 (O_938,N_12823,N_14683);
and UO_939 (O_939,N_13483,N_11859);
and UO_940 (O_940,N_12518,N_13189);
and UO_941 (O_941,N_11702,N_10877);
and UO_942 (O_942,N_12907,N_10206);
and UO_943 (O_943,N_12936,N_11476);
and UO_944 (O_944,N_12991,N_12388);
or UO_945 (O_945,N_12056,N_11787);
nor UO_946 (O_946,N_10810,N_12600);
or UO_947 (O_947,N_12979,N_14409);
or UO_948 (O_948,N_14001,N_11162);
nor UO_949 (O_949,N_14410,N_11167);
and UO_950 (O_950,N_12989,N_11635);
nand UO_951 (O_951,N_11341,N_13078);
or UO_952 (O_952,N_12023,N_13091);
or UO_953 (O_953,N_12183,N_11191);
xor UO_954 (O_954,N_11002,N_12299);
or UO_955 (O_955,N_12263,N_14377);
nor UO_956 (O_956,N_14251,N_11007);
nand UO_957 (O_957,N_14625,N_13569);
xor UO_958 (O_958,N_13273,N_13874);
nand UO_959 (O_959,N_13551,N_12692);
and UO_960 (O_960,N_13119,N_14312);
or UO_961 (O_961,N_10404,N_14583);
and UO_962 (O_962,N_12360,N_10148);
or UO_963 (O_963,N_11560,N_13314);
nand UO_964 (O_964,N_11259,N_11312);
xnor UO_965 (O_965,N_12624,N_12455);
nand UO_966 (O_966,N_14614,N_11922);
and UO_967 (O_967,N_11323,N_10120);
and UO_968 (O_968,N_13743,N_13844);
nor UO_969 (O_969,N_10630,N_11627);
nor UO_970 (O_970,N_11620,N_12486);
and UO_971 (O_971,N_12459,N_11395);
xnor UO_972 (O_972,N_10381,N_12345);
and UO_973 (O_973,N_13325,N_11754);
or UO_974 (O_974,N_12064,N_10716);
xnor UO_975 (O_975,N_12193,N_10584);
and UO_976 (O_976,N_12013,N_14891);
or UO_977 (O_977,N_13801,N_14296);
nor UO_978 (O_978,N_14383,N_13898);
xor UO_979 (O_979,N_10762,N_11986);
nor UO_980 (O_980,N_11233,N_12195);
or UO_981 (O_981,N_11217,N_14380);
and UO_982 (O_982,N_12366,N_11867);
or UO_983 (O_983,N_13364,N_11980);
xnor UO_984 (O_984,N_12625,N_11487);
xnor UO_985 (O_985,N_14268,N_12305);
nand UO_986 (O_986,N_10435,N_12052);
xnor UO_987 (O_987,N_14943,N_11418);
or UO_988 (O_988,N_13294,N_10339);
nand UO_989 (O_989,N_10115,N_12836);
xnor UO_990 (O_990,N_14492,N_10322);
nand UO_991 (O_991,N_12755,N_12565);
or UO_992 (O_992,N_10862,N_14556);
nor UO_993 (O_993,N_10640,N_13048);
xnor UO_994 (O_994,N_12598,N_13693);
or UO_995 (O_995,N_10983,N_14139);
nor UO_996 (O_996,N_13101,N_14445);
and UO_997 (O_997,N_11995,N_14057);
xor UO_998 (O_998,N_10520,N_11388);
nor UO_999 (O_999,N_10902,N_11928);
nand UO_1000 (O_1000,N_10633,N_10938);
nor UO_1001 (O_1001,N_14168,N_14814);
xnor UO_1002 (O_1002,N_13426,N_11666);
nor UO_1003 (O_1003,N_10041,N_10755);
and UO_1004 (O_1004,N_13290,N_11201);
nand UO_1005 (O_1005,N_14284,N_10617);
nand UO_1006 (O_1006,N_10696,N_14759);
and UO_1007 (O_1007,N_13730,N_14175);
xor UO_1008 (O_1008,N_10798,N_13083);
nand UO_1009 (O_1009,N_10969,N_14553);
xnor UO_1010 (O_1010,N_13762,N_11865);
nand UO_1011 (O_1011,N_10905,N_12112);
or UO_1012 (O_1012,N_13795,N_14812);
or UO_1013 (O_1013,N_10965,N_13864);
xor UO_1014 (O_1014,N_10551,N_11125);
nand UO_1015 (O_1015,N_13716,N_10377);
and UO_1016 (O_1016,N_14157,N_14358);
or UO_1017 (O_1017,N_11590,N_10342);
and UO_1018 (O_1018,N_10835,N_12132);
nand UO_1019 (O_1019,N_12584,N_10403);
nor UO_1020 (O_1020,N_11670,N_14295);
xnor UO_1021 (O_1021,N_14613,N_12068);
nor UO_1022 (O_1022,N_11944,N_11883);
and UO_1023 (O_1023,N_12825,N_14762);
and UO_1024 (O_1024,N_10449,N_12636);
nand UO_1025 (O_1025,N_12054,N_12613);
nor UO_1026 (O_1026,N_12214,N_10481);
xnor UO_1027 (O_1027,N_13539,N_14056);
nand UO_1028 (O_1028,N_10759,N_12284);
nor UO_1029 (O_1029,N_14372,N_11735);
nor UO_1030 (O_1030,N_13339,N_11955);
nand UO_1031 (O_1031,N_11503,N_13954);
and UO_1032 (O_1032,N_11437,N_14716);
xor UO_1033 (O_1033,N_14654,N_10888);
xor UO_1034 (O_1034,N_10567,N_11089);
nor UO_1035 (O_1035,N_10097,N_12321);
nand UO_1036 (O_1036,N_12088,N_11929);
or UO_1037 (O_1037,N_14305,N_12325);
or UO_1038 (O_1038,N_13666,N_11038);
or UO_1039 (O_1039,N_14895,N_11152);
nor UO_1040 (O_1040,N_13507,N_11831);
or UO_1041 (O_1041,N_14487,N_12181);
nor UO_1042 (O_1042,N_12027,N_10891);
nand UO_1043 (O_1043,N_11314,N_12275);
nor UO_1044 (O_1044,N_12982,N_10557);
xnor UO_1045 (O_1045,N_10307,N_12167);
xnor UO_1046 (O_1046,N_13269,N_14481);
and UO_1047 (O_1047,N_10719,N_10913);
or UO_1048 (O_1048,N_11618,N_10235);
xnor UO_1049 (O_1049,N_13145,N_12756);
or UO_1050 (O_1050,N_10055,N_13560);
nor UO_1051 (O_1051,N_10470,N_13139);
nor UO_1052 (O_1052,N_11493,N_10952);
and UO_1053 (O_1053,N_13872,N_11141);
nor UO_1054 (O_1054,N_12458,N_10274);
xnor UO_1055 (O_1055,N_10445,N_11541);
nor UO_1056 (O_1056,N_13870,N_10208);
nand UO_1057 (O_1057,N_14184,N_10149);
nand UO_1058 (O_1058,N_10144,N_11202);
or UO_1059 (O_1059,N_14639,N_14571);
or UO_1060 (O_1060,N_13980,N_13543);
nand UO_1061 (O_1061,N_11649,N_11077);
nor UO_1062 (O_1062,N_14177,N_13605);
nand UO_1063 (O_1063,N_14341,N_14096);
and UO_1064 (O_1064,N_14003,N_13825);
and UO_1065 (O_1065,N_11589,N_12622);
and UO_1066 (O_1066,N_11362,N_14170);
nor UO_1067 (O_1067,N_10651,N_10099);
or UO_1068 (O_1068,N_10290,N_10145);
nor UO_1069 (O_1069,N_14275,N_12016);
xor UO_1070 (O_1070,N_12558,N_12032);
xor UO_1071 (O_1071,N_10405,N_11767);
or UO_1072 (O_1072,N_13686,N_11707);
and UO_1073 (O_1073,N_11948,N_12469);
xor UO_1074 (O_1074,N_13782,N_10281);
nand UO_1075 (O_1075,N_10391,N_10188);
nand UO_1076 (O_1076,N_10313,N_14122);
xnor UO_1077 (O_1077,N_10263,N_13695);
and UO_1078 (O_1078,N_10552,N_12946);
nor UO_1079 (O_1079,N_14222,N_10580);
or UO_1080 (O_1080,N_14508,N_11289);
xor UO_1081 (O_1081,N_14903,N_14944);
xnor UO_1082 (O_1082,N_11927,N_13465);
nor UO_1083 (O_1083,N_10394,N_10255);
or UO_1084 (O_1084,N_11782,N_14788);
and UO_1085 (O_1085,N_10761,N_14801);
xor UO_1086 (O_1086,N_11254,N_10076);
and UO_1087 (O_1087,N_10165,N_13847);
nor UO_1088 (O_1088,N_13597,N_10490);
or UO_1089 (O_1089,N_10695,N_13983);
or UO_1090 (O_1090,N_11056,N_14869);
xor UO_1091 (O_1091,N_10997,N_11414);
nor UO_1092 (O_1092,N_10741,N_14897);
nand UO_1093 (O_1093,N_10800,N_10801);
xnor UO_1094 (O_1094,N_14471,N_10745);
nand UO_1095 (O_1095,N_10727,N_14530);
nand UO_1096 (O_1096,N_12897,N_12961);
nor UO_1097 (O_1097,N_11039,N_14000);
nor UO_1098 (O_1098,N_12393,N_13878);
nand UO_1099 (O_1099,N_11761,N_11801);
or UO_1100 (O_1100,N_12862,N_10150);
or UO_1101 (O_1101,N_13363,N_10702);
or UO_1102 (O_1102,N_14451,N_14351);
nor UO_1103 (O_1103,N_13358,N_13163);
xnor UO_1104 (O_1104,N_13103,N_14904);
nand UO_1105 (O_1105,N_14772,N_14459);
nand UO_1106 (O_1106,N_12501,N_14108);
xor UO_1107 (O_1107,N_12910,N_12143);
or UO_1108 (O_1108,N_10297,N_11538);
xnor UO_1109 (O_1109,N_11357,N_13496);
or UO_1110 (O_1110,N_12853,N_12331);
or UO_1111 (O_1111,N_12453,N_12426);
xnor UO_1112 (O_1112,N_10945,N_14596);
nor UO_1113 (O_1113,N_11496,N_12377);
nand UO_1114 (O_1114,N_14005,N_12634);
and UO_1115 (O_1115,N_14290,N_11916);
xnor UO_1116 (O_1116,N_11283,N_14171);
xor UO_1117 (O_1117,N_11532,N_10805);
xnor UO_1118 (O_1118,N_11511,N_11392);
nand UO_1119 (O_1119,N_13857,N_11715);
or UO_1120 (O_1120,N_13960,N_13321);
xnor UO_1121 (O_1121,N_13845,N_11575);
and UO_1122 (O_1122,N_10524,N_12247);
xnor UO_1123 (O_1123,N_13128,N_13098);
or UO_1124 (O_1124,N_14853,N_11359);
nor UO_1125 (O_1125,N_14894,N_11058);
nor UO_1126 (O_1126,N_10040,N_12992);
nor UO_1127 (O_1127,N_11829,N_14580);
and UO_1128 (O_1128,N_12171,N_14180);
nand UO_1129 (O_1129,N_12379,N_11041);
nor UO_1130 (O_1130,N_13032,N_12276);
and UO_1131 (O_1131,N_14292,N_14845);
or UO_1132 (O_1132,N_12244,N_10942);
or UO_1133 (O_1133,N_12049,N_10927);
or UO_1134 (O_1134,N_10631,N_14272);
nor UO_1135 (O_1135,N_12609,N_11778);
or UO_1136 (O_1136,N_12324,N_10114);
nand UO_1137 (O_1137,N_13794,N_11035);
or UO_1138 (O_1138,N_13041,N_12053);
xnor UO_1139 (O_1139,N_13127,N_14084);
xor UO_1140 (O_1140,N_13143,N_14528);
xnor UO_1141 (O_1141,N_11595,N_14359);
nor UO_1142 (O_1142,N_11475,N_10079);
nand UO_1143 (O_1143,N_12071,N_14352);
nor UO_1144 (O_1144,N_13443,N_10495);
and UO_1145 (O_1145,N_11042,N_11795);
nor UO_1146 (O_1146,N_14825,N_12352);
and UO_1147 (O_1147,N_14905,N_11579);
nand UO_1148 (O_1148,N_12086,N_14455);
and UO_1149 (O_1149,N_13976,N_12718);
and UO_1150 (O_1150,N_12467,N_14469);
nand UO_1151 (O_1151,N_10598,N_13596);
and UO_1152 (O_1152,N_10151,N_14664);
nand UO_1153 (O_1153,N_12984,N_11265);
xnor UO_1154 (O_1154,N_10456,N_13778);
xor UO_1155 (O_1155,N_11222,N_11999);
nand UO_1156 (O_1156,N_10958,N_11884);
xor UO_1157 (O_1157,N_13637,N_14126);
nand UO_1158 (O_1158,N_11132,N_10395);
nand UO_1159 (O_1159,N_14435,N_11105);
nor UO_1160 (O_1160,N_14784,N_11722);
or UO_1161 (O_1161,N_12429,N_12858);
xor UO_1162 (O_1162,N_11471,N_14651);
xor UO_1163 (O_1163,N_13087,N_12978);
or UO_1164 (O_1164,N_13657,N_11960);
and UO_1165 (O_1165,N_14183,N_10892);
or UO_1166 (O_1166,N_11841,N_10440);
xnor UO_1167 (O_1167,N_14976,N_12028);
or UO_1168 (O_1168,N_12789,N_14373);
xnor UO_1169 (O_1169,N_14440,N_10735);
nor UO_1170 (O_1170,N_10416,N_12207);
or UO_1171 (O_1171,N_14100,N_12416);
xnor UO_1172 (O_1172,N_10610,N_12399);
xor UO_1173 (O_1173,N_11964,N_14226);
and UO_1174 (O_1174,N_11053,N_11446);
nor UO_1175 (O_1175,N_13479,N_12492);
and UO_1176 (O_1176,N_12318,N_14748);
or UO_1177 (O_1177,N_13995,N_14700);
nand UO_1178 (O_1178,N_12595,N_11553);
nand UO_1179 (O_1179,N_14110,N_10329);
and UO_1180 (O_1180,N_14243,N_13247);
nor UO_1181 (O_1181,N_13458,N_12908);
nand UO_1182 (O_1182,N_11913,N_10325);
and UO_1183 (O_1183,N_14536,N_11137);
or UO_1184 (O_1184,N_10207,N_10002);
nand UO_1185 (O_1185,N_13608,N_13601);
xnor UO_1186 (O_1186,N_13277,N_12655);
and UO_1187 (O_1187,N_11142,N_13838);
xor UO_1188 (O_1188,N_13787,N_12146);
nor UO_1189 (O_1189,N_10568,N_14926);
and UO_1190 (O_1190,N_14417,N_14999);
nand UO_1191 (O_1191,N_12236,N_13681);
nor UO_1192 (O_1192,N_11296,N_11389);
xor UO_1193 (O_1193,N_13662,N_11869);
nand UO_1194 (O_1194,N_11934,N_13308);
or UO_1195 (O_1195,N_10363,N_10062);
nor UO_1196 (O_1196,N_12691,N_12981);
and UO_1197 (O_1197,N_11853,N_10818);
or UO_1198 (O_1198,N_11623,N_13816);
nor UO_1199 (O_1199,N_10454,N_12349);
xnor UO_1200 (O_1200,N_10043,N_10231);
nor UO_1201 (O_1201,N_12177,N_12498);
and UO_1202 (O_1202,N_12639,N_12413);
or UO_1203 (O_1203,N_13320,N_13586);
nor UO_1204 (O_1204,N_10897,N_12082);
and UO_1205 (O_1205,N_11083,N_14097);
nand UO_1206 (O_1206,N_11270,N_12676);
xnor UO_1207 (O_1207,N_12654,N_12094);
nor UO_1208 (O_1208,N_11433,N_10020);
nand UO_1209 (O_1209,N_14566,N_11067);
or UO_1210 (O_1210,N_14912,N_13049);
or UO_1211 (O_1211,N_14354,N_11444);
or UO_1212 (O_1212,N_13956,N_10819);
and UO_1213 (O_1213,N_12669,N_12533);
nand UO_1214 (O_1214,N_11277,N_13330);
or UO_1215 (O_1215,N_14040,N_11769);
nand UO_1216 (O_1216,N_11062,N_13896);
or UO_1217 (O_1217,N_12835,N_10432);
and UO_1218 (O_1218,N_13979,N_10278);
xor UO_1219 (O_1219,N_14901,N_12473);
nand UO_1220 (O_1220,N_14855,N_12966);
or UO_1221 (O_1221,N_10293,N_13410);
xor UO_1222 (O_1222,N_14236,N_11683);
nand UO_1223 (O_1223,N_11065,N_14518);
nor UO_1224 (O_1224,N_14681,N_10698);
nor UO_1225 (O_1225,N_10316,N_11208);
xnor UO_1226 (O_1226,N_13014,N_10999);
nor UO_1227 (O_1227,N_14985,N_11712);
and UO_1228 (O_1228,N_12084,N_10726);
xnor UO_1229 (O_1229,N_14854,N_11403);
or UO_1230 (O_1230,N_14579,N_12629);
nor UO_1231 (O_1231,N_10995,N_10365);
xor UO_1232 (O_1232,N_11023,N_14870);
or UO_1233 (O_1233,N_13705,N_10378);
and UO_1234 (O_1234,N_14722,N_12846);
and UO_1235 (O_1235,N_12296,N_14837);
xnor UO_1236 (O_1236,N_10185,N_14181);
nor UO_1237 (O_1237,N_14960,N_11567);
and UO_1238 (O_1238,N_11317,N_12900);
or UO_1239 (O_1239,N_10656,N_11858);
nor UO_1240 (O_1240,N_14963,N_14747);
nand UO_1241 (O_1241,N_10645,N_11349);
or UO_1242 (O_1242,N_13433,N_12259);
nor UO_1243 (O_1243,N_13559,N_10625);
xnor UO_1244 (O_1244,N_11989,N_11055);
and UO_1245 (O_1245,N_11288,N_10471);
nor UO_1246 (O_1246,N_13036,N_10370);
nor UO_1247 (O_1247,N_11293,N_13533);
xnor UO_1248 (O_1248,N_13141,N_12545);
and UO_1249 (O_1249,N_12905,N_10219);
and UO_1250 (O_1250,N_10091,N_13510);
xnor UO_1251 (O_1251,N_14190,N_11318);
xnor UO_1252 (O_1252,N_14977,N_13518);
and UO_1253 (O_1253,N_10218,N_13811);
xnor UO_1254 (O_1254,N_11231,N_12728);
xnor UO_1255 (O_1255,N_11585,N_11118);
nor UO_1256 (O_1256,N_13526,N_14010);
xor UO_1257 (O_1257,N_12221,N_14711);
nand UO_1258 (O_1258,N_14198,N_14636);
and UO_1259 (O_1259,N_11003,N_12342);
or UO_1260 (O_1260,N_12749,N_12543);
nor UO_1261 (O_1261,N_10910,N_13123);
nor UO_1262 (O_1262,N_11350,N_10007);
and UO_1263 (O_1263,N_13588,N_11198);
xnor UO_1264 (O_1264,N_14261,N_11203);
and UO_1265 (O_1265,N_12569,N_10514);
nor UO_1266 (O_1266,N_10220,N_12330);
xor UO_1267 (O_1267,N_12375,N_10898);
and UO_1268 (O_1268,N_14240,N_11892);
xnor UO_1269 (O_1269,N_14494,N_11534);
nor UO_1270 (O_1270,N_13206,N_11179);
xor UO_1271 (O_1271,N_10065,N_11537);
xnor UO_1272 (O_1272,N_12044,N_10957);
xnor UO_1273 (O_1273,N_12409,N_10644);
and UO_1274 (O_1274,N_10754,N_10202);
or UO_1275 (O_1275,N_13159,N_10838);
nor UO_1276 (O_1276,N_11686,N_11614);
or UO_1277 (O_1277,N_12727,N_11888);
xor UO_1278 (O_1278,N_11632,N_14389);
xor UO_1279 (O_1279,N_11307,N_12590);
or UO_1280 (O_1280,N_10946,N_14782);
nor UO_1281 (O_1281,N_10448,N_13282);
and UO_1282 (O_1282,N_14200,N_13490);
nand UO_1283 (O_1283,N_12220,N_14829);
or UO_1284 (O_1284,N_14027,N_14327);
and UO_1285 (O_1285,N_13692,N_12246);
and UO_1286 (O_1286,N_10787,N_13740);
xor UO_1287 (O_1287,N_14339,N_14345);
xor UO_1288 (O_1288,N_11122,N_10627);
nor UO_1289 (O_1289,N_12928,N_13999);
nor UO_1290 (O_1290,N_13854,N_10742);
and UO_1291 (O_1291,N_10676,N_11877);
xor UO_1292 (O_1292,N_10384,N_12705);
or UO_1293 (O_1293,N_12739,N_13981);
or UO_1294 (O_1294,N_12687,N_10353);
nand UO_1295 (O_1295,N_10154,N_11933);
and UO_1296 (O_1296,N_12940,N_13888);
and UO_1297 (O_1297,N_13387,N_11343);
nand UO_1298 (O_1298,N_13382,N_11462);
nand UO_1299 (O_1299,N_10611,N_11325);
nor UO_1300 (O_1300,N_14039,N_12909);
nor UO_1301 (O_1301,N_14062,N_13170);
and UO_1302 (O_1302,N_14162,N_14014);
xnor UO_1303 (O_1303,N_12753,N_10244);
or UO_1304 (O_1304,N_14655,N_10306);
and UO_1305 (O_1305,N_11126,N_10034);
or UO_1306 (O_1306,N_10407,N_10212);
xor UO_1307 (O_1307,N_13425,N_10948);
nor UO_1308 (O_1308,N_12525,N_11153);
and UO_1309 (O_1309,N_11247,N_14401);
nand UO_1310 (O_1310,N_10412,N_10533);
and UO_1311 (O_1311,N_13934,N_12868);
or UO_1312 (O_1312,N_10575,N_14843);
or UO_1313 (O_1313,N_11546,N_13234);
or UO_1314 (O_1314,N_10878,N_12601);
or UO_1315 (O_1315,N_11165,N_13904);
or UO_1316 (O_1316,N_13892,N_11747);
and UO_1317 (O_1317,N_14672,N_13651);
nor UO_1318 (O_1318,N_10637,N_14304);
nand UO_1319 (O_1319,N_10506,N_14575);
and UO_1320 (O_1320,N_11236,N_14797);
and UO_1321 (O_1321,N_11347,N_14090);
xor UO_1322 (O_1322,N_10250,N_11173);
nor UO_1323 (O_1323,N_11211,N_10634);
xnor UO_1324 (O_1324,N_10251,N_14739);
nand UO_1325 (O_1325,N_13058,N_11704);
nor UO_1326 (O_1326,N_13445,N_13489);
xor UO_1327 (O_1327,N_10229,N_13630);
xor UO_1328 (O_1328,N_11713,N_12551);
xnor UO_1329 (O_1329,N_10715,N_12363);
nand UO_1330 (O_1330,N_13310,N_11178);
xnor UO_1331 (O_1331,N_12194,N_12725);
nor UO_1332 (O_1332,N_13930,N_14093);
nand UO_1333 (O_1333,N_10919,N_10802);
and UO_1334 (O_1334,N_12405,N_14375);
nor UO_1335 (O_1335,N_13066,N_10709);
nor UO_1336 (O_1336,N_10593,N_12785);
or UO_1337 (O_1337,N_11084,N_13360);
xnor UO_1338 (O_1338,N_10057,N_12578);
nor UO_1339 (O_1339,N_10101,N_10401);
or UO_1340 (O_1340,N_11120,N_13475);
and UO_1341 (O_1341,N_14730,N_11967);
nor UO_1342 (O_1342,N_14561,N_11969);
nor UO_1343 (O_1343,N_12680,N_11584);
xnor UO_1344 (O_1344,N_14427,N_14464);
xor UO_1345 (O_1345,N_12225,N_11398);
xnor UO_1346 (O_1346,N_11439,N_14328);
and UO_1347 (O_1347,N_12520,N_10458);
nand UO_1348 (O_1348,N_14402,N_10738);
and UO_1349 (O_1349,N_13932,N_10906);
and UO_1350 (O_1350,N_12527,N_12564);
or UO_1351 (O_1351,N_13520,N_14131);
or UO_1352 (O_1352,N_14591,N_10026);
nor UO_1353 (O_1353,N_14344,N_13400);
xor UO_1354 (O_1354,N_12237,N_12987);
and UO_1355 (O_1355,N_10455,N_13957);
nor UO_1356 (O_1356,N_13476,N_10108);
and UO_1357 (O_1357,N_14823,N_13114);
nand UO_1358 (O_1358,N_11544,N_11640);
nand UO_1359 (O_1359,N_11438,N_14506);
nand UO_1360 (O_1360,N_12280,N_13353);
or UO_1361 (O_1361,N_10451,N_14114);
xnor UO_1362 (O_1362,N_10414,N_13137);
and UO_1363 (O_1363,N_12290,N_13511);
or UO_1364 (O_1364,N_12076,N_10666);
nor UO_1365 (O_1365,N_12881,N_10472);
nand UO_1366 (O_1366,N_14301,N_10051);
or UO_1367 (O_1367,N_13647,N_11494);
nor UO_1368 (O_1368,N_10840,N_13381);
or UO_1369 (O_1369,N_12414,N_11988);
or UO_1370 (O_1370,N_14507,N_11566);
or UO_1371 (O_1371,N_11550,N_14847);
nor UO_1372 (O_1372,N_11977,N_11303);
or UO_1373 (O_1373,N_10277,N_11383);
nor UO_1374 (O_1374,N_12017,N_14185);
and UO_1375 (O_1375,N_12353,N_10332);
nor UO_1376 (O_1376,N_14917,N_11193);
or UO_1377 (O_1377,N_13622,N_11423);
and UO_1378 (O_1378,N_10746,N_13694);
and UO_1379 (O_1379,N_11866,N_11517);
and UO_1380 (O_1380,N_12707,N_12239);
or UO_1381 (O_1381,N_14618,N_14447);
and UO_1382 (O_1382,N_10853,N_11535);
xnor UO_1383 (O_1383,N_10187,N_12248);
nand UO_1384 (O_1384,N_14138,N_12254);
or UO_1385 (O_1385,N_11856,N_13215);
and UO_1386 (O_1386,N_12121,N_13877);
nand UO_1387 (O_1387,N_12781,N_11514);
nand UO_1388 (O_1388,N_12119,N_13736);
and UO_1389 (O_1389,N_12468,N_10809);
nor UO_1390 (O_1390,N_11071,N_10907);
nand UO_1391 (O_1391,N_12673,N_11628);
nor UO_1392 (O_1392,N_11719,N_10739);
nand UO_1393 (O_1393,N_11966,N_13564);
nand UO_1394 (O_1394,N_13528,N_13226);
nand UO_1395 (O_1395,N_14054,N_14294);
and UO_1396 (O_1396,N_13438,N_10603);
or UO_1397 (O_1397,N_12810,N_13198);
nor UO_1398 (O_1398,N_11386,N_13080);
nor UO_1399 (O_1399,N_11710,N_14968);
and UO_1400 (O_1400,N_12850,N_12711);
nor UO_1401 (O_1401,N_14074,N_14578);
nand UO_1402 (O_1402,N_12339,N_12382);
nor UO_1403 (O_1403,N_12483,N_12935);
xor UO_1404 (O_1404,N_13975,N_10042);
or UO_1405 (O_1405,N_11749,N_13379);
nand UO_1406 (O_1406,N_11147,N_13607);
nor UO_1407 (O_1407,N_11631,N_10970);
xnor UO_1408 (O_1408,N_10475,N_11827);
nand UO_1409 (O_1409,N_10035,N_14208);
nor UO_1410 (O_1410,N_14779,N_12430);
or UO_1411 (O_1411,N_13691,N_12320);
or UO_1412 (O_1412,N_10864,N_13587);
and UO_1413 (O_1413,N_12732,N_13724);
nor UO_1414 (O_1414,N_12653,N_13760);
nand UO_1415 (O_1415,N_11355,N_14371);
or UO_1416 (O_1416,N_10222,N_11169);
xor UO_1417 (O_1417,N_13986,N_10776);
xnor UO_1418 (O_1418,N_12849,N_11942);
and UO_1419 (O_1419,N_12949,N_11486);
and UO_1420 (O_1420,N_13350,N_13432);
nor UO_1421 (O_1421,N_12951,N_10443);
or UO_1422 (O_1422,N_14631,N_12464);
nor UO_1423 (O_1423,N_10847,N_14983);
nand UO_1424 (O_1424,N_11835,N_11730);
and UO_1425 (O_1425,N_13799,N_11737);
xor UO_1426 (O_1426,N_13916,N_14049);
and UO_1427 (O_1427,N_11861,N_14497);
and UO_1428 (O_1428,N_13010,N_14188);
nand UO_1429 (O_1429,N_13391,N_11181);
nor UO_1430 (O_1430,N_11849,N_11512);
nor UO_1431 (O_1431,N_14568,N_11022);
nor UO_1432 (O_1432,N_12602,N_13665);
xor UO_1433 (O_1433,N_13658,N_13278);
nand UO_1434 (O_1434,N_13933,N_10087);
xnor UO_1435 (O_1435,N_10884,N_11554);
xnor UO_1436 (O_1436,N_12631,N_11652);
nor UO_1437 (O_1437,N_11044,N_11024);
nand UO_1438 (O_1438,N_11468,N_14009);
nor UO_1439 (O_1439,N_12435,N_14846);
xor UO_1440 (O_1440,N_14656,N_11854);
nand UO_1441 (O_1441,N_12113,N_14979);
nor UO_1442 (O_1442,N_14356,N_12557);
nand UO_1443 (O_1443,N_13347,N_14549);
or UO_1444 (O_1444,N_11721,N_10740);
nand UO_1445 (O_1445,N_10849,N_10260);
xnor UO_1446 (O_1446,N_11138,N_11779);
xor UO_1447 (O_1447,N_10771,N_11073);
and UO_1448 (O_1448,N_11417,N_13759);
xor UO_1449 (O_1449,N_13126,N_14723);
nor UO_1450 (O_1450,N_11256,N_10832);
xor UO_1451 (O_1451,N_12510,N_10118);
and UO_1452 (O_1452,N_10683,N_10786);
xnor UO_1453 (O_1453,N_12014,N_12690);
xnor UO_1454 (O_1454,N_12462,N_11688);
and UO_1455 (O_1455,N_10782,N_12460);
nand UO_1456 (O_1456,N_10932,N_12741);
xor UO_1457 (O_1457,N_12228,N_12499);
nand UO_1458 (O_1458,N_13741,N_10379);
xor UO_1459 (O_1459,N_14199,N_11111);
and UO_1460 (O_1460,N_13913,N_14610);
and UO_1461 (O_1461,N_12334,N_14330);
xor UO_1462 (O_1462,N_13744,N_10519);
xnor UO_1463 (O_1463,N_10390,N_11833);
and UO_1464 (O_1464,N_13376,N_11814);
nor UO_1465 (O_1465,N_12668,N_13659);
xnor UO_1466 (O_1466,N_11014,N_11876);
xor UO_1467 (O_1467,N_11748,N_11095);
nand UO_1468 (O_1468,N_10534,N_10032);
nor UO_1469 (O_1469,N_13297,N_10968);
nor UO_1470 (O_1470,N_12758,N_14933);
and UO_1471 (O_1471,N_14288,N_14452);
xnor UO_1472 (O_1472,N_11376,N_12449);
nand UO_1473 (O_1473,N_10657,N_14316);
and UO_1474 (O_1474,N_14245,N_11816);
or UO_1475 (O_1475,N_14648,N_13663);
or UO_1476 (O_1476,N_14031,N_14187);
nor UO_1477 (O_1477,N_10226,N_13461);
or UO_1478 (O_1478,N_11224,N_12186);
and UO_1479 (O_1479,N_13368,N_12135);
or UO_1480 (O_1480,N_10837,N_10758);
xor UO_1481 (O_1481,N_10133,N_11207);
and UO_1482 (O_1482,N_14164,N_10070);
xor UO_1483 (O_1483,N_10371,N_12953);
and UO_1484 (O_1484,N_14008,N_14346);
nor UO_1485 (O_1485,N_10170,N_12485);
nand UO_1486 (O_1486,N_14698,N_12730);
nor UO_1487 (O_1487,N_14935,N_13502);
nand UO_1488 (O_1488,N_13236,N_11577);
or UO_1489 (O_1489,N_13181,N_11744);
nand UO_1490 (O_1490,N_12278,N_13911);
nor UO_1491 (O_1491,N_11763,N_14218);
xor UO_1492 (O_1492,N_12370,N_11881);
xnor UO_1493 (O_1493,N_11803,N_10784);
and UO_1494 (O_1494,N_12802,N_10223);
nor UO_1495 (O_1495,N_13102,N_10056);
nor UO_1496 (O_1496,N_13075,N_11629);
nor UO_1497 (O_1497,N_11016,N_10348);
or UO_1498 (O_1498,N_10717,N_10844);
nor UO_1499 (O_1499,N_14221,N_13401);
and UO_1500 (O_1500,N_11012,N_14174);
and UO_1501 (O_1501,N_12715,N_10510);
xnor UO_1502 (O_1502,N_13237,N_11337);
nor UO_1503 (O_1503,N_13998,N_10804);
or UO_1504 (O_1504,N_11372,N_13351);
xor UO_1505 (O_1505,N_13148,N_13184);
nand UO_1506 (O_1506,N_10690,N_12040);
xor UO_1507 (O_1507,N_10205,N_14247);
nand UO_1508 (O_1508,N_14871,N_14277);
and UO_1509 (O_1509,N_14117,N_13699);
xnor UO_1510 (O_1510,N_12035,N_14378);
or UO_1511 (O_1511,N_14033,N_14322);
xor UO_1512 (O_1512,N_13367,N_12931);
xor UO_1513 (O_1513,N_11253,N_11321);
and UO_1514 (O_1514,N_13213,N_11774);
or UO_1515 (O_1515,N_14034,N_10478);
nor UO_1516 (O_1516,N_12311,N_14726);
nand UO_1517 (O_1517,N_11880,N_13503);
xnor UO_1518 (O_1518,N_13464,N_13756);
xnor UO_1519 (O_1519,N_13210,N_13504);
nand UO_1520 (O_1520,N_13403,N_13242);
or UO_1521 (O_1521,N_13581,N_14013);
or UO_1522 (O_1522,N_13281,N_13887);
and UO_1523 (O_1523,N_10949,N_10502);
nor UO_1524 (O_1524,N_13045,N_14547);
xor UO_1525 (O_1525,N_12766,N_11049);
or UO_1526 (O_1526,N_14908,N_10488);
xor UO_1527 (O_1527,N_10856,N_10734);
nor UO_1528 (O_1528,N_12403,N_11279);
xnor UO_1529 (O_1529,N_11101,N_10078);
xor UO_1530 (O_1530,N_14934,N_13536);
nor UO_1531 (O_1531,N_13488,N_11759);
xnor UO_1532 (O_1532,N_12385,N_11637);
nor UO_1533 (O_1533,N_11353,N_14966);
nand UO_1534 (O_1534,N_11911,N_12277);
xor UO_1535 (O_1535,N_11543,N_12128);
and UO_1536 (O_1536,N_10469,N_11286);
xnor UO_1537 (O_1537,N_12252,N_10411);
nand UO_1538 (O_1538,N_12535,N_10872);
or UO_1539 (O_1539,N_14605,N_10100);
nand UO_1540 (O_1540,N_10960,N_12661);
nand UO_1541 (O_1541,N_14309,N_11699);
nor UO_1542 (O_1542,N_10086,N_11606);
xor UO_1543 (O_1543,N_11574,N_12960);
nand UO_1544 (O_1544,N_14112,N_11973);
nand UO_1545 (O_1545,N_11021,N_14603);
and UO_1546 (O_1546,N_10691,N_11633);
xor UO_1547 (O_1547,N_11171,N_10797);
nand UO_1548 (O_1548,N_14642,N_11930);
nand UO_1549 (O_1549,N_10850,N_13927);
or UO_1550 (O_1550,N_11885,N_13454);
or UO_1551 (O_1551,N_14018,N_13901);
and UO_1552 (O_1552,N_10117,N_14264);
xnor UO_1553 (O_1553,N_14706,N_14771);
or UO_1554 (O_1554,N_13396,N_10825);
xnor UO_1555 (O_1555,N_12744,N_14682);
or UO_1556 (O_1556,N_10555,N_11369);
nand UO_1557 (O_1557,N_12514,N_10090);
nor UO_1558 (O_1558,N_13808,N_10166);
nand UO_1559 (O_1559,N_10763,N_13190);
nor UO_1560 (O_1560,N_12139,N_11788);
nor UO_1561 (O_1561,N_13446,N_10694);
or UO_1562 (O_1562,N_11248,N_14512);
nand UO_1563 (O_1563,N_14085,N_14714);
xor UO_1564 (O_1564,N_13111,N_12090);
nand UO_1565 (O_1565,N_12447,N_13194);
nor UO_1566 (O_1566,N_14584,N_10396);
nor UO_1567 (O_1567,N_12689,N_11411);
nor UO_1568 (O_1568,N_14087,N_10998);
nand UO_1569 (O_1569,N_14473,N_13711);
and UO_1570 (O_1570,N_14848,N_10925);
or UO_1571 (O_1571,N_11910,N_12771);
xor UO_1572 (O_1572,N_14597,N_10216);
and UO_1573 (O_1573,N_10038,N_14931);
xnor UO_1574 (O_1574,N_11155,N_12500);
and UO_1575 (O_1575,N_11982,N_11504);
nor UO_1576 (O_1576,N_12202,N_13709);
and UO_1577 (O_1577,N_10122,N_13354);
xor UO_1578 (O_1578,N_11611,N_14258);
and UO_1579 (O_1579,N_13978,N_10813);
nor UO_1580 (O_1580,N_13881,N_13812);
xnor UO_1581 (O_1581,N_11672,N_13582);
or UO_1582 (O_1582,N_14368,N_14391);
or UO_1583 (O_1583,N_10783,N_12975);
xor UO_1584 (O_1584,N_14235,N_12745);
xor UO_1585 (O_1585,N_14564,N_10388);
xnor UO_1586 (O_1586,N_11110,N_14733);
xnor UO_1587 (O_1587,N_12039,N_12642);
or UO_1588 (O_1588,N_14576,N_14671);
or UO_1589 (O_1589,N_12315,N_13449);
nor UO_1590 (O_1590,N_13418,N_12003);
xor UO_1591 (O_1591,N_12930,N_11939);
or UO_1592 (O_1592,N_11703,N_12322);
nor UO_1593 (O_1593,N_14736,N_10459);
nor UO_1594 (O_1594,N_12481,N_13899);
nand UO_1595 (O_1595,N_14594,N_13090);
xor UO_1596 (O_1596,N_12927,N_10012);
and UO_1597 (O_1597,N_10444,N_14832);
or UO_1598 (O_1598,N_13875,N_12559);
nand UO_1599 (O_1599,N_10830,N_13883);
xor UO_1600 (O_1600,N_10287,N_12842);
xor UO_1601 (O_1601,N_13346,N_12537);
nor UO_1602 (O_1602,N_11896,N_10186);
and UO_1603 (O_1603,N_13784,N_11621);
xnor UO_1604 (O_1604,N_11692,N_13384);
or UO_1605 (O_1605,N_11170,N_10663);
or UO_1606 (O_1606,N_14606,N_14770);
nor UO_1607 (O_1607,N_13645,N_11206);
and UO_1608 (O_1608,N_14206,N_12260);
and UO_1609 (O_1609,N_10024,N_13704);
xor UO_1610 (O_1610,N_14444,N_11921);
and UO_1611 (O_1611,N_10337,N_14816);
or UO_1612 (O_1612,N_14360,N_13279);
or UO_1613 (O_1613,N_13334,N_12988);
and UO_1614 (O_1614,N_10362,N_11932);
and UO_1615 (O_1615,N_14676,N_10338);
and UO_1616 (O_1616,N_12596,N_14167);
xor UO_1617 (O_1617,N_12872,N_12580);
nand UO_1618 (O_1618,N_11515,N_11596);
nor UO_1619 (O_1619,N_14215,N_13567);
nor UO_1620 (O_1620,N_10654,N_14615);
xor UO_1621 (O_1621,N_14045,N_13380);
xnor UO_1622 (O_1622,N_13258,N_14942);
nor UO_1623 (O_1623,N_12892,N_14381);
or UO_1624 (O_1624,N_13178,N_13013);
nand UO_1625 (O_1625,N_10240,N_10183);
xnor UO_1626 (O_1626,N_11378,N_12200);
nor UO_1627 (O_1627,N_13664,N_12251);
xnor UO_1628 (O_1628,N_11127,N_10245);
xnor UO_1629 (O_1629,N_12562,N_10480);
or UO_1630 (O_1630,N_10426,N_11320);
nand UO_1631 (O_1631,N_13019,N_14203);
nor UO_1632 (O_1632,N_10845,N_11440);
or UO_1633 (O_1633,N_11102,N_11917);
and UO_1634 (O_1634,N_13070,N_14342);
nand UO_1635 (O_1635,N_13193,N_11936);
nand UO_1636 (O_1636,N_13486,N_13831);
nand UO_1637 (O_1637,N_14306,N_13316);
nor UO_1638 (O_1638,N_10189,N_12106);
nand UO_1639 (O_1639,N_12818,N_10896);
or UO_1640 (O_1640,N_10064,N_10641);
nor UO_1641 (O_1641,N_12684,N_11001);
and UO_1642 (O_1642,N_11879,N_13820);
or UO_1643 (O_1643,N_12415,N_11473);
nor UO_1644 (O_1644,N_13317,N_12861);
or UO_1645 (O_1645,N_13295,N_11045);
or UO_1646 (O_1646,N_14070,N_11599);
or UO_1647 (O_1647,N_11245,N_11379);
xor UO_1648 (O_1648,N_11792,N_11561);
and UO_1649 (O_1649,N_13889,N_10372);
nand UO_1650 (O_1650,N_12007,N_11063);
or UO_1651 (O_1651,N_13809,N_12748);
and UO_1652 (O_1652,N_11139,N_11998);
xor UO_1653 (O_1653,N_14675,N_14002);
and UO_1654 (O_1654,N_10530,N_13472);
and UO_1655 (O_1655,N_14282,N_11290);
nor UO_1656 (O_1656,N_13687,N_11430);
or UO_1657 (O_1657,N_11810,N_11559);
and UO_1658 (O_1658,N_11891,N_12821);
nor UO_1659 (O_1659,N_13365,N_14279);
nand UO_1660 (O_1660,N_12101,N_13469);
nand UO_1661 (O_1661,N_11292,N_12879);
and UO_1662 (O_1662,N_14836,N_13963);
and UO_1663 (O_1663,N_14278,N_11284);
and UO_1664 (O_1664,N_13436,N_12838);
nor UO_1665 (O_1665,N_11555,N_10273);
xnor UO_1666 (O_1666,N_10177,N_13093);
nand UO_1667 (O_1667,N_11622,N_13468);
and UO_1668 (O_1668,N_13650,N_12061);
xor UO_1669 (O_1669,N_11834,N_12714);
xor UO_1670 (O_1670,N_12432,N_12392);
or UO_1671 (O_1671,N_14686,N_10565);
or UO_1672 (O_1672,N_11445,N_14906);
nand UO_1673 (O_1673,N_11194,N_10320);
nand UO_1674 (O_1674,N_13557,N_11800);
and UO_1675 (O_1675,N_12250,N_13244);
xor UO_1676 (O_1676,N_14388,N_14856);
and UO_1677 (O_1677,N_10930,N_13617);
nand UO_1678 (O_1678,N_12286,N_11393);
nand UO_1679 (O_1679,N_12157,N_14718);
nand UO_1680 (O_1680,N_10581,N_14815);
and UO_1681 (O_1681,N_10723,N_12180);
xor UO_1682 (O_1682,N_14805,N_13891);
and UO_1683 (O_1683,N_14896,N_10704);
and UO_1684 (O_1684,N_11551,N_12147);
and UO_1685 (O_1685,N_10089,N_14047);
nand UO_1686 (O_1686,N_13749,N_10857);
or UO_1687 (O_1687,N_11826,N_10578);
xor UO_1688 (O_1688,N_11519,N_11509);
xnor UO_1689 (O_1689,N_13500,N_13893);
xor UO_1690 (O_1690,N_10619,N_11940);
nor UO_1691 (O_1691,N_12945,N_14852);
and UO_1692 (O_1692,N_12955,N_14280);
nand UO_1693 (O_1693,N_14990,N_10851);
nor UO_1694 (O_1694,N_13576,N_11066);
or UO_1695 (O_1695,N_12097,N_13929);
xnor UO_1696 (O_1696,N_14940,N_10418);
and UO_1697 (O_1697,N_13275,N_11860);
or UO_1698 (O_1698,N_11477,N_13228);
and UO_1699 (O_1699,N_11249,N_10349);
xor UO_1700 (O_1700,N_12795,N_12792);
xor UO_1701 (O_1701,N_13924,N_14265);
nor UO_1702 (O_1702,N_12356,N_13300);
and UO_1703 (O_1703,N_12072,N_11422);
xnor UO_1704 (O_1704,N_12722,N_12694);
and UO_1705 (O_1705,N_13251,N_11197);
or UO_1706 (O_1706,N_11889,N_14974);
nand UO_1707 (O_1707,N_11954,N_11641);
nand UO_1708 (O_1708,N_11086,N_12130);
xnor UO_1709 (O_1709,N_13311,N_10242);
xnor UO_1710 (O_1710,N_12105,N_12648);
nor UO_1711 (O_1711,N_12227,N_14925);
xnor UO_1712 (O_1712,N_14501,N_12976);
nand UO_1713 (O_1713,N_12015,N_10743);
or UO_1714 (O_1714,N_14754,N_14291);
nor UO_1715 (O_1715,N_12301,N_12394);
and UO_1716 (O_1716,N_10116,N_13291);
or UO_1717 (O_1717,N_14559,N_13451);
nand UO_1718 (O_1718,N_14189,N_11906);
nand UO_1719 (O_1719,N_10636,N_14514);
or UO_1720 (O_1720,N_10629,N_11306);
or UO_1721 (O_1721,N_12826,N_12347);
and UO_1722 (O_1722,N_10926,N_12297);
or UO_1723 (O_1723,N_13336,N_12359);
xnor UO_1724 (O_1724,N_14920,N_13453);
nand UO_1725 (O_1725,N_10612,N_13022);
nand UO_1726 (O_1726,N_14543,N_13563);
or UO_1727 (O_1727,N_14608,N_10505);
nor UO_1728 (O_1728,N_11547,N_14362);
xnor UO_1729 (O_1729,N_10138,N_11616);
or UO_1730 (O_1730,N_13220,N_14405);
and UO_1731 (O_1731,N_14333,N_14111);
xnor UO_1732 (O_1732,N_13940,N_11447);
or UO_1733 (O_1733,N_11785,N_12083);
nand UO_1734 (O_1734,N_10668,N_10431);
or UO_1735 (O_1735,N_13623,N_14412);
and UO_1736 (O_1736,N_11524,N_11094);
xnor UO_1737 (O_1737,N_11557,N_14367);
and UO_1738 (O_1738,N_14796,N_14505);
or UO_1739 (O_1739,N_14880,N_11926);
or UO_1740 (O_1740,N_12764,N_11434);
xor UO_1741 (O_1741,N_12901,N_11333);
and UO_1742 (O_1742,N_14132,N_13395);
xnor UO_1743 (O_1743,N_13550,N_11070);
xnor UO_1744 (O_1744,N_10509,N_10105);
nand UO_1745 (O_1745,N_14083,N_10310);
and UO_1746 (O_1746,N_14349,N_12660);
nor UO_1747 (O_1747,N_13207,N_14775);
nor UO_1748 (O_1748,N_12786,N_10828);
nand UO_1749 (O_1749,N_14785,N_13038);
nand UO_1750 (O_1750,N_11420,N_12723);
xor UO_1751 (O_1751,N_13777,N_11750);
and UO_1752 (O_1752,N_13672,N_11729);
nor UO_1753 (O_1753,N_10376,N_13130);
or UO_1754 (O_1754,N_14400,N_10302);
or UO_1755 (O_1755,N_12314,N_12380);
nand UO_1756 (O_1756,N_10442,N_14868);
nor UO_1757 (O_1757,N_11639,N_13252);
or UO_1758 (O_1758,N_12057,N_13217);
xor UO_1759 (O_1759,N_14077,N_11410);
xor UO_1760 (O_1760,N_14728,N_10446);
nand UO_1761 (O_1761,N_10817,N_14873);
nand UO_1762 (O_1762,N_10895,N_13107);
nor UO_1763 (O_1763,N_11663,N_10494);
nand UO_1764 (O_1764,N_12454,N_13335);
nand UO_1765 (O_1765,N_12257,N_13535);
nor UO_1766 (O_1766,N_10450,N_12120);
nand UO_1767 (O_1767,N_13408,N_14376);
or UO_1768 (O_1768,N_14602,N_14075);
xor UO_1769 (O_1769,N_12555,N_13708);
nand UO_1770 (O_1770,N_13524,N_14136);
nor UO_1771 (O_1771,N_11088,N_10046);
nand UO_1772 (O_1772,N_12906,N_12378);
and UO_1773 (O_1773,N_13552,N_12549);
or UO_1774 (O_1774,N_13040,N_14886);
nor UO_1775 (O_1775,N_10210,N_12422);
and UO_1776 (O_1776,N_13393,N_14998);
or UO_1777 (O_1777,N_11578,N_12412);
or UO_1778 (O_1778,N_11266,N_13392);
and UO_1779 (O_1779,N_10112,N_14130);
xor UO_1780 (O_1780,N_12030,N_13843);
and UO_1781 (O_1781,N_13056,N_11319);
xnor UO_1782 (O_1782,N_14091,N_12424);
or UO_1783 (O_1783,N_11682,N_14092);
nand UO_1784 (O_1784,N_14161,N_11828);
and UO_1785 (O_1785,N_14281,N_12666);
or UO_1786 (O_1786,N_10535,N_10681);
nor UO_1787 (O_1787,N_11415,N_14233);
nor UO_1788 (O_1788,N_14363,N_14725);
and UO_1789 (O_1789,N_12529,N_12734);
xnor UO_1790 (O_1790,N_14426,N_12811);
or UO_1791 (O_1791,N_13943,N_11264);
nand UO_1792 (O_1792,N_11026,N_14513);
and UO_1793 (O_1793,N_14205,N_10991);
nand UO_1794 (O_1794,N_14460,N_11764);
xor UO_1795 (O_1795,N_14124,N_11241);
xnor UO_1796 (O_1796,N_13158,N_14485);
and UO_1797 (O_1797,N_13319,N_14554);
nor UO_1798 (O_1798,N_12210,N_14317);
or UO_1799 (O_1799,N_14293,N_10546);
nor UO_1800 (O_1800,N_14949,N_11646);
and UO_1801 (O_1801,N_14238,N_11983);
and UO_1802 (O_1802,N_12926,N_12294);
xor UO_1803 (O_1803,N_10054,N_11280);
xor UO_1804 (O_1804,N_10706,N_12099);
xor UO_1805 (O_1805,N_13804,N_11351);
xor UO_1806 (O_1806,N_14827,N_12591);
nor UO_1807 (O_1807,N_10900,N_13696);
or UO_1808 (O_1808,N_12461,N_14015);
nand UO_1809 (O_1809,N_14822,N_13214);
xor UO_1810 (O_1810,N_14972,N_12450);
xnor UO_1811 (O_1811,N_13553,N_12145);
nor UO_1812 (O_1812,N_10083,N_11213);
nand UO_1813 (O_1813,N_11691,N_12997);
xor UO_1814 (O_1814,N_13416,N_13240);
and UO_1815 (O_1815,N_11527,N_12465);
nor UO_1816 (O_1816,N_11373,N_12383);
nor UO_1817 (O_1817,N_13928,N_14030);
and UO_1818 (O_1818,N_13573,N_14260);
xor UO_1819 (O_1819,N_10769,N_13150);
nor UO_1820 (O_1820,N_14332,N_14971);
xnor UO_1821 (O_1821,N_13274,N_13624);
or UO_1822 (O_1822,N_13337,N_13327);
or UO_1823 (O_1823,N_10779,N_10249);
nor UO_1824 (O_1824,N_11870,N_12046);
nor UO_1825 (O_1825,N_12570,N_14120);
nor UO_1826 (O_1826,N_13970,N_11978);
nor UO_1827 (O_1827,N_13750,N_12706);
nand UO_1828 (O_1828,N_14379,N_11878);
xnor UO_1829 (O_1829,N_11220,N_10614);
nand UO_1830 (O_1830,N_12201,N_12109);
or UO_1831 (O_1831,N_13021,N_10944);
xor UO_1832 (O_1832,N_10984,N_12149);
or UO_1833 (O_1833,N_13146,N_10326);
or UO_1834 (O_1834,N_13772,N_10940);
xor UO_1835 (O_1835,N_13338,N_12136);
nor UO_1836 (O_1836,N_11427,N_14657);
and UO_1837 (O_1837,N_14545,N_10298);
or UO_1838 (O_1838,N_14993,N_10066);
nand UO_1839 (O_1839,N_12530,N_11791);
nor UO_1840 (O_1840,N_14213,N_10620);
and UO_1841 (O_1841,N_14523,N_14419);
nand UO_1842 (O_1842,N_11997,N_14807);
and UO_1843 (O_1843,N_10624,N_14022);
xor UO_1844 (O_1844,N_14789,N_10889);
nor UO_1845 (O_1845,N_11230,N_10589);
nor UO_1846 (O_1846,N_10369,N_14470);
or UO_1847 (O_1847,N_12974,N_13950);
xor UO_1848 (O_1848,N_13613,N_11484);
xor UO_1849 (O_1849,N_14708,N_14624);
or UO_1850 (O_1850,N_13842,N_10538);
nor UO_1851 (O_1851,N_11674,N_13684);
nor UO_1852 (O_1852,N_13962,N_11605);
nor UO_1853 (O_1853,N_12561,N_11407);
nand UO_1854 (O_1854,N_12482,N_14252);
and UO_1855 (O_1855,N_11506,N_14539);
xor UO_1856 (O_1856,N_10119,N_10536);
and UO_1857 (O_1857,N_10408,N_13988);
nand UO_1858 (O_1858,N_13071,N_14719);
and UO_1859 (O_1859,N_10563,N_14626);
nor UO_1860 (O_1860,N_12952,N_14997);
nor UO_1861 (O_1861,N_11993,N_13713);
or UO_1862 (O_1862,N_10858,N_10594);
xnor UO_1863 (O_1863,N_14795,N_14866);
and UO_1864 (O_1864,N_13062,N_12918);
nor UO_1865 (O_1865,N_11068,N_12652);
nor UO_1866 (O_1866,N_14321,N_11790);
and UO_1867 (O_1867,N_12649,N_11338);
and UO_1868 (O_1868,N_11752,N_12308);
xnor UO_1869 (O_1869,N_11820,N_13374);
or UO_1870 (O_1870,N_10639,N_11772);
or UO_1871 (O_1871,N_13615,N_12439);
and UO_1872 (O_1872,N_13897,N_12031);
xor UO_1873 (O_1873,N_14922,N_13836);
nor UO_1874 (O_1874,N_10269,N_14165);
nand UO_1875 (O_1875,N_13342,N_14403);
or UO_1876 (O_1876,N_13627,N_13906);
nor UO_1877 (O_1877,N_14089,N_12651);
nand UO_1878 (O_1878,N_11738,N_13246);
and UO_1879 (O_1879,N_12216,N_14604);
or UO_1880 (O_1880,N_14776,N_10655);
and UO_1881 (O_1881,N_13776,N_11273);
or UO_1882 (O_1882,N_13020,N_13689);
or UO_1883 (O_1883,N_11412,N_12807);
xnor UO_1884 (O_1884,N_10848,N_11657);
nand UO_1885 (O_1885,N_14038,N_10981);
and UO_1886 (O_1886,N_13841,N_12266);
nor UO_1887 (O_1887,N_12406,N_12470);
nand UO_1888 (O_1888,N_12395,N_11655);
xnor UO_1889 (O_1889,N_10356,N_10904);
and UO_1890 (O_1890,N_12588,N_14142);
nand UO_1891 (O_1891,N_11872,N_10954);
or UO_1892 (O_1892,N_14336,N_11466);
nand UO_1893 (O_1893,N_10674,N_12258);
nor UO_1894 (O_1894,N_12340,N_12708);
xnor UO_1895 (O_1895,N_13450,N_14589);
xnor UO_1896 (O_1896,N_12969,N_11302);
nand UO_1897 (O_1897,N_11251,N_10111);
xnor UO_1898 (O_1898,N_10643,N_13626);
or UO_1899 (O_1899,N_14817,N_12215);
xnor UO_1900 (O_1900,N_12182,N_12283);
xnor UO_1901 (O_1901,N_14996,N_14413);
xnor UO_1902 (O_1902,N_10867,N_12620);
xnor UO_1903 (O_1903,N_12066,N_12346);
or UO_1904 (O_1904,N_13880,N_13286);
nor UO_1905 (O_1905,N_14424,N_12358);
xor UO_1906 (O_1906,N_10508,N_10980);
nand UO_1907 (O_1907,N_14382,N_12381);
nor UO_1908 (O_1908,N_11327,N_10230);
or UO_1909 (O_1909,N_10541,N_10234);
nor UO_1910 (O_1910,N_10515,N_11117);
xnor UO_1911 (O_1911,N_10547,N_11391);
nor UO_1912 (O_1912,N_13612,N_14393);
xnor UO_1913 (O_1913,N_11714,N_10661);
nor UO_1914 (O_1914,N_13061,N_10831);
and UO_1915 (O_1915,N_11608,N_13774);
nand UO_1916 (O_1916,N_14123,N_11027);
nand UO_1917 (O_1917,N_14191,N_13629);
and UO_1918 (O_1918,N_10031,N_13628);
nand UO_1919 (O_1919,N_12476,N_12091);
xnor UO_1920 (O_1920,N_10943,N_14833);
nor UO_1921 (O_1921,N_12205,N_10744);
xor UO_1922 (O_1922,N_11607,N_11479);
nand UO_1923 (O_1923,N_10102,N_12190);
or UO_1924 (O_1924,N_14721,N_14884);
and UO_1925 (O_1925,N_13621,N_10841);
xor UO_1926 (O_1926,N_12168,N_12647);
nor UO_1927 (O_1927,N_12144,N_13243);
nand UO_1928 (O_1928,N_13715,N_12423);
and UO_1929 (O_1929,N_12166,N_10184);
nand UO_1930 (O_1930,N_13255,N_11813);
or UO_1931 (O_1931,N_14643,N_14028);
and UO_1932 (O_1932,N_11136,N_13671);
or UO_1933 (O_1933,N_11013,N_13909);
xnor UO_1934 (O_1934,N_13097,N_10596);
or UO_1935 (O_1935,N_10345,N_14520);
nand UO_1936 (O_1936,N_11696,N_12367);
and UO_1937 (O_1937,N_11844,N_12029);
nor UO_1938 (O_1938,N_10564,N_14558);
or UO_1939 (O_1939,N_13781,N_12420);
nor UO_1940 (O_1940,N_13508,N_14653);
nand UO_1941 (O_1941,N_14500,N_12466);
or UO_1942 (O_1942,N_10161,N_12985);
nand UO_1943 (O_1943,N_12777,N_12542);
and UO_1944 (O_1944,N_13485,N_10049);
xnor UO_1945 (O_1945,N_10652,N_12579);
xnor UO_1946 (O_1946,N_13521,N_12899);
and UO_1947 (O_1947,N_12281,N_10225);
or UO_1948 (O_1948,N_11382,N_12824);
and UO_1949 (O_1949,N_11190,N_12502);
and UO_1950 (O_1950,N_14060,N_10084);
or UO_1951 (O_1951,N_10213,N_11701);
or UO_1952 (O_1952,N_12812,N_10855);
xnor UO_1953 (O_1953,N_14478,N_11436);
and UO_1954 (O_1954,N_14020,N_14209);
or UO_1955 (O_1955,N_14720,N_14482);
and UO_1956 (O_1956,N_11716,N_10193);
nor UO_1957 (O_1957,N_13677,N_14619);
or UO_1958 (O_1958,N_11773,N_13618);
and UO_1959 (O_1959,N_12963,N_14555);
or UO_1960 (O_1960,N_14160,N_13135);
nor UO_1961 (O_1961,N_14550,N_14418);
and UO_1962 (O_1962,N_14659,N_12203);
nand UO_1963 (O_1963,N_13270,N_11483);
or UO_1964 (O_1964,N_12407,N_12688);
or UO_1965 (O_1965,N_13108,N_10618);
or UO_1966 (O_1966,N_11223,N_11215);
xor UO_1967 (O_1967,N_12575,N_11187);
or UO_1968 (O_1968,N_12073,N_12587);
xor UO_1969 (O_1969,N_12519,N_13547);
and UO_1970 (O_1970,N_12110,N_11124);
or UO_1971 (O_1971,N_10623,N_13324);
or UO_1972 (O_1972,N_12965,N_10861);
or UO_1973 (O_1973,N_14433,N_11971);
nand UO_1974 (O_1974,N_11664,N_13501);
nand UO_1975 (O_1975,N_12137,N_11276);
and UO_1976 (O_1976,N_12191,N_14783);
xnor UO_1977 (O_1977,N_10486,N_11765);
nand UO_1978 (O_1978,N_13745,N_10756);
xor UO_1979 (O_1979,N_13361,N_14149);
and UO_1980 (O_1980,N_14562,N_12302);
xor UO_1981 (O_1981,N_12874,N_12913);
xnor UO_1982 (O_1982,N_12253,N_14248);
nor UO_1983 (O_1983,N_13375,N_10410);
nand UO_1984 (O_1984,N_11793,N_11209);
or UO_1985 (O_1985,N_12867,N_11812);
xnor UO_1986 (O_1986,N_12075,N_13411);
nand UO_1987 (O_1987,N_13283,N_14778);
and UO_1988 (O_1988,N_12508,N_10466);
nand UO_1989 (O_1989,N_11135,N_13497);
and UO_1990 (O_1990,N_11057,N_13333);
nor UO_1991 (O_1991,N_11580,N_14303);
nor UO_1992 (O_1992,N_12941,N_11272);
or UO_1993 (O_1993,N_10693,N_13871);
or UO_1994 (O_1994,N_11309,N_10441);
xnor UO_1995 (O_1995,N_12993,N_14929);
and UO_1996 (O_1996,N_11004,N_13639);
nand UO_1997 (O_1997,N_11576,N_12041);
and UO_1998 (O_1998,N_14230,N_10914);
nor UO_1999 (O_1999,N_11717,N_10873);
endmodule