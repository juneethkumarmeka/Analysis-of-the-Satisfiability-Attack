module basic_2500_25000_3000_25_levels_10xor_4(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999;
or U0 (N_0,In_741,In_2362);
nor U1 (N_1,In_332,In_2009);
nand U2 (N_2,In_1846,In_2264);
xnor U3 (N_3,In_574,In_1399);
nor U4 (N_4,In_1038,In_1835);
nor U5 (N_5,In_837,In_2066);
xnor U6 (N_6,In_15,In_471);
nand U7 (N_7,In_218,In_1071);
and U8 (N_8,In_2171,In_275);
nor U9 (N_9,In_853,In_844);
xor U10 (N_10,In_1438,In_337);
nor U11 (N_11,In_2206,In_2368);
xor U12 (N_12,In_801,In_1173);
nor U13 (N_13,In_599,In_2297);
xnor U14 (N_14,In_344,In_2234);
xor U15 (N_15,In_1431,In_1903);
and U16 (N_16,In_1840,In_1356);
or U17 (N_17,In_1333,In_1497);
nand U18 (N_18,In_526,In_1755);
nand U19 (N_19,In_1691,In_988);
nand U20 (N_20,In_1437,In_1077);
nand U21 (N_21,In_1853,In_433);
nor U22 (N_22,In_809,In_1666);
and U23 (N_23,In_1486,In_380);
nor U24 (N_24,In_2486,In_958);
or U25 (N_25,In_2281,In_2011);
and U26 (N_26,In_1396,In_871);
nor U27 (N_27,In_1563,In_1007);
nor U28 (N_28,In_1641,In_1810);
xor U29 (N_29,In_1440,In_1093);
nand U30 (N_30,In_2284,In_2496);
nand U31 (N_31,In_1229,In_2378);
and U32 (N_32,In_750,In_919);
nand U33 (N_33,In_1752,In_695);
and U34 (N_34,In_2044,In_894);
nand U35 (N_35,In_927,In_989);
nor U36 (N_36,In_2217,In_852);
and U37 (N_37,In_1867,In_2299);
xnor U38 (N_38,In_30,In_1490);
or U39 (N_39,In_1579,In_999);
and U40 (N_40,In_502,In_1717);
and U41 (N_41,In_805,In_167);
and U42 (N_42,In_1900,In_444);
xnor U43 (N_43,In_1032,In_1513);
or U44 (N_44,In_354,In_628);
and U45 (N_45,In_702,In_1605);
and U46 (N_46,In_1714,In_2448);
or U47 (N_47,In_2177,In_81);
nand U48 (N_48,In_87,In_1545);
and U49 (N_49,In_469,In_1599);
nor U50 (N_50,In_688,In_1448);
nor U51 (N_51,In_1028,In_651);
or U52 (N_52,In_464,In_1557);
nand U53 (N_53,In_1912,In_1943);
xnor U54 (N_54,In_2466,In_1530);
nand U55 (N_55,In_1811,In_2157);
nor U56 (N_56,In_1451,In_1461);
and U57 (N_57,In_1842,In_1978);
xor U58 (N_58,In_296,In_1672);
or U59 (N_59,In_864,In_933);
and U60 (N_60,In_2000,In_279);
nand U61 (N_61,In_2189,In_2006);
nand U62 (N_62,In_1073,In_1331);
xnor U63 (N_63,In_292,In_585);
nand U64 (N_64,In_1577,In_727);
xor U65 (N_65,In_730,In_2382);
nor U66 (N_66,In_2344,In_1705);
nand U67 (N_67,In_1583,In_2393);
or U68 (N_68,In_1155,In_869);
nor U69 (N_69,In_257,In_495);
or U70 (N_70,In_2335,In_1242);
nor U71 (N_71,In_2012,In_2019);
and U72 (N_72,In_940,In_1823);
nor U73 (N_73,In_2439,In_1962);
nand U74 (N_74,In_973,In_2174);
nor U75 (N_75,In_1467,In_390);
or U76 (N_76,In_2455,In_1056);
xnor U77 (N_77,In_1013,In_69);
nand U78 (N_78,In_1041,In_2256);
nand U79 (N_79,In_1266,In_1020);
xnor U80 (N_80,In_726,In_1296);
or U81 (N_81,In_2470,In_2111);
and U82 (N_82,In_1571,In_2016);
xnor U83 (N_83,In_2031,In_2034);
nand U84 (N_84,In_1997,In_2330);
nor U85 (N_85,In_2384,In_169);
nor U86 (N_86,In_1015,In_24);
and U87 (N_87,In_439,In_348);
xor U88 (N_88,In_482,In_385);
xor U89 (N_89,In_393,In_2262);
and U90 (N_90,In_422,In_1427);
nand U91 (N_91,In_1170,In_731);
or U92 (N_92,In_1342,In_445);
and U93 (N_93,In_357,In_58);
or U94 (N_94,In_2039,In_2208);
nand U95 (N_95,In_56,In_1094);
or U96 (N_96,In_37,In_429);
nor U97 (N_97,In_216,In_589);
or U98 (N_98,In_2027,In_1243);
nor U99 (N_99,In_1021,In_1446);
xor U100 (N_100,In_388,In_879);
or U101 (N_101,In_2225,In_2422);
xor U102 (N_102,In_545,In_1830);
nor U103 (N_103,In_1036,In_2246);
and U104 (N_104,In_639,In_2205);
and U105 (N_105,In_607,In_114);
nor U106 (N_106,In_2360,In_2464);
xor U107 (N_107,In_995,In_787);
or U108 (N_108,In_1559,In_2190);
or U109 (N_109,In_909,In_1471);
or U110 (N_110,In_515,In_165);
xor U111 (N_111,In_1286,In_492);
nor U112 (N_112,In_1368,In_1487);
or U113 (N_113,In_478,In_1673);
xor U114 (N_114,In_276,In_499);
nor U115 (N_115,In_1759,In_341);
xnor U116 (N_116,In_711,In_1152);
or U117 (N_117,In_67,In_1227);
and U118 (N_118,In_249,In_66);
nor U119 (N_119,In_2210,In_2159);
nor U120 (N_120,In_1350,In_16);
and U121 (N_121,In_398,In_360);
nor U122 (N_122,In_2449,In_2168);
and U123 (N_123,In_2351,In_1532);
xnor U124 (N_124,In_387,In_1147);
and U125 (N_125,In_534,In_2417);
or U126 (N_126,In_1580,In_2101);
and U127 (N_127,In_1249,In_1768);
or U128 (N_128,In_412,In_2093);
nor U129 (N_129,In_1332,In_925);
and U130 (N_130,In_1313,In_774);
and U131 (N_131,In_850,In_2338);
xnor U132 (N_132,In_1125,In_1265);
xor U133 (N_133,In_1773,In_1955);
nand U134 (N_134,In_1709,In_729);
and U135 (N_135,In_855,In_1153);
nor U136 (N_136,In_548,In_2004);
nand U137 (N_137,In_238,In_1697);
or U138 (N_138,In_1345,In_1087);
and U139 (N_139,In_2383,In_818);
nor U140 (N_140,In_1099,In_704);
and U141 (N_141,In_2107,In_1283);
nor U142 (N_142,In_1185,In_2228);
nor U143 (N_143,In_1841,In_912);
or U144 (N_144,In_1126,In_1880);
or U145 (N_145,In_551,In_2235);
nor U146 (N_146,In_1181,In_1863);
or U147 (N_147,In_2251,In_1062);
xor U148 (N_148,In_1831,In_366);
xnor U149 (N_149,In_1587,In_2002);
nor U150 (N_150,In_1561,In_2421);
nor U151 (N_151,In_578,In_1683);
nand U152 (N_152,In_703,In_1740);
or U153 (N_153,In_1798,In_1988);
or U154 (N_154,In_2279,In_1570);
nor U155 (N_155,In_2267,In_1963);
xor U156 (N_156,In_991,In_2261);
nor U157 (N_157,In_1377,In_2114);
and U158 (N_158,In_2186,In_1800);
or U159 (N_159,In_778,In_2347);
and U160 (N_160,In_142,In_2325);
and U161 (N_161,In_816,In_1460);
and U162 (N_162,In_1116,In_1108);
and U163 (N_163,In_435,In_1732);
and U164 (N_164,In_880,In_486);
and U165 (N_165,In_448,In_566);
or U166 (N_166,In_27,In_459);
nand U167 (N_167,In_2062,In_2143);
and U168 (N_168,In_1820,In_2275);
and U169 (N_169,In_840,In_1419);
or U170 (N_170,In_1716,In_1980);
or U171 (N_171,In_1945,In_2124);
xor U172 (N_172,In_61,In_1888);
nand U173 (N_173,In_440,In_769);
nand U174 (N_174,In_671,In_2373);
nand U175 (N_175,In_94,In_1837);
and U176 (N_176,In_1707,In_996);
nand U177 (N_177,In_1290,In_60);
xor U178 (N_178,In_594,In_1151);
nor U179 (N_179,In_1104,In_99);
or U180 (N_180,In_1874,In_1075);
xnor U181 (N_181,In_792,In_2078);
nor U182 (N_182,In_2428,In_1877);
nor U183 (N_183,In_2434,In_568);
xnor U184 (N_184,In_1310,In_267);
xnor U185 (N_185,In_590,In_969);
nand U186 (N_186,In_1107,In_23);
or U187 (N_187,In_2154,In_1336);
and U188 (N_188,In_2165,In_320);
or U189 (N_189,In_569,In_1211);
xnor U190 (N_190,In_1002,In_1293);
and U191 (N_191,In_1416,In_1726);
and U192 (N_192,In_1277,In_728);
and U193 (N_193,In_2028,In_1967);
or U194 (N_194,In_725,In_2241);
xnor U195 (N_195,In_1989,In_2468);
nor U196 (N_196,In_1034,In_2088);
nand U197 (N_197,In_1189,In_1479);
nor U198 (N_198,In_1162,In_1654);
xnor U199 (N_199,In_665,In_2444);
nor U200 (N_200,In_1700,In_1141);
xnor U201 (N_201,In_524,In_1534);
xnor U202 (N_202,In_1627,In_1982);
nand U203 (N_203,In_713,In_2071);
nand U204 (N_204,In_2243,In_705);
or U205 (N_205,In_1857,In_1710);
nand U206 (N_206,In_100,In_13);
and U207 (N_207,In_1085,In_214);
nand U208 (N_208,In_2460,In_2491);
nand U209 (N_209,In_2179,In_2112);
xnor U210 (N_210,In_1589,In_442);
or U211 (N_211,In_2084,In_309);
nand U212 (N_212,In_795,In_1337);
and U213 (N_213,In_1839,In_1897);
and U214 (N_214,In_1334,In_1936);
or U215 (N_215,In_633,In_137);
nor U216 (N_216,In_552,In_2119);
and U217 (N_217,In_1423,In_1402);
nor U218 (N_218,In_1262,In_2318);
xor U219 (N_219,In_179,In_2076);
nor U220 (N_220,In_1044,In_586);
xnor U221 (N_221,In_473,In_978);
nor U222 (N_222,In_1953,In_1893);
xnor U223 (N_223,In_1971,In_694);
xnor U224 (N_224,In_1426,In_1119);
and U225 (N_225,In_1158,In_1680);
xnor U226 (N_226,In_954,In_1414);
and U227 (N_227,In_289,In_2479);
and U228 (N_228,In_981,In_1715);
nor U229 (N_229,In_1782,In_1433);
nor U230 (N_230,In_431,In_274);
or U231 (N_231,In_1976,In_1515);
nand U232 (N_232,In_1896,In_2254);
and U233 (N_233,In_897,In_685);
or U234 (N_234,In_2472,In_1655);
and U235 (N_235,In_755,In_781);
xor U236 (N_236,In_561,In_902);
and U237 (N_237,In_807,In_1592);
and U238 (N_238,In_191,In_1168);
nor U239 (N_239,In_162,In_1059);
or U240 (N_240,In_2103,In_734);
xor U241 (N_241,In_106,In_131);
xor U242 (N_242,In_2024,In_2369);
or U243 (N_243,In_1043,In_168);
and U244 (N_244,In_377,In_224);
xnor U245 (N_245,In_1081,In_197);
xor U246 (N_246,In_111,In_378);
xor U247 (N_247,In_1338,In_753);
nand U248 (N_248,In_468,In_2415);
xor U249 (N_249,In_1394,In_262);
nand U250 (N_250,In_1393,In_959);
xor U251 (N_251,In_2278,In_135);
or U252 (N_252,In_889,In_2113);
nand U253 (N_253,In_491,In_19);
and U254 (N_254,In_1648,In_1470);
nand U255 (N_255,In_686,In_406);
nor U256 (N_256,In_1001,In_2280);
xor U257 (N_257,In_88,In_183);
and U258 (N_258,In_1795,In_1991);
nand U259 (N_259,In_2086,In_895);
nor U260 (N_260,In_535,In_1324);
or U261 (N_261,In_2072,In_1380);
nand U262 (N_262,In_1979,In_992);
xor U263 (N_263,In_339,In_1581);
or U264 (N_264,In_1407,In_294);
or U265 (N_265,In_301,In_700);
nand U266 (N_266,In_1864,In_392);
nand U267 (N_267,In_353,In_1814);
nand U268 (N_268,In_775,In_434);
and U269 (N_269,In_122,In_536);
or U270 (N_270,In_1847,In_384);
or U271 (N_271,In_985,In_2258);
nand U272 (N_272,In_1502,In_2075);
nand U273 (N_273,In_884,In_1805);
or U274 (N_274,In_1088,In_1042);
and U275 (N_275,In_1016,In_0);
xor U276 (N_276,In_2129,In_1959);
and U277 (N_277,In_2437,In_963);
xnor U278 (N_278,In_1466,In_2425);
and U279 (N_279,In_2222,In_1022);
nand U280 (N_280,In_2381,In_1496);
nand U281 (N_281,In_635,In_219);
nor U282 (N_282,In_881,In_2277);
or U283 (N_283,In_1425,In_1983);
nor U284 (N_284,In_2478,In_557);
or U285 (N_285,In_558,In_605);
or U286 (N_286,In_474,In_2257);
or U287 (N_287,In_2252,In_1871);
or U288 (N_288,In_2495,In_1204);
or U289 (N_289,In_347,In_972);
nor U290 (N_290,In_29,In_1165);
and U291 (N_291,In_656,In_1111);
or U292 (N_292,In_441,In_1960);
or U293 (N_293,In_784,In_321);
nand U294 (N_294,In_145,In_2282);
nand U295 (N_295,In_1475,In_2357);
and U296 (N_296,In_1731,In_173);
nor U297 (N_297,In_1499,In_982);
xnor U298 (N_298,In_546,In_359);
xor U299 (N_299,In_1808,In_358);
and U300 (N_300,In_2355,In_1972);
and U301 (N_301,In_1052,In_653);
nand U302 (N_302,In_1698,In_1363);
xor U303 (N_303,In_2286,In_1913);
nand U304 (N_304,In_1272,In_1067);
nand U305 (N_305,In_1564,In_1112);
nand U306 (N_306,In_1634,In_654);
nor U307 (N_307,In_2010,In_643);
nand U308 (N_308,In_2013,In_663);
nor U309 (N_309,In_2183,In_556);
nand U310 (N_310,In_231,In_1027);
xnor U311 (N_311,In_1120,In_1230);
nor U312 (N_312,In_1878,In_693);
or U313 (N_313,In_230,In_1614);
nor U314 (N_314,In_1617,In_698);
and U315 (N_315,In_1183,In_225);
xor U316 (N_316,In_1033,In_2390);
xor U317 (N_317,In_1434,In_1636);
nor U318 (N_318,In_2120,In_1160);
nand U319 (N_319,In_1939,In_1196);
nor U320 (N_320,In_2008,In_119);
nor U321 (N_321,In_1488,In_1319);
or U322 (N_322,In_1215,In_1082);
or U323 (N_323,In_1794,In_1734);
or U324 (N_324,In_1205,In_2483);
xor U325 (N_325,In_2400,In_305);
nand U326 (N_326,In_1103,In_185);
xor U327 (N_327,In_767,In_1253);
nand U328 (N_328,In_1373,In_836);
nor U329 (N_329,In_1809,In_314);
or U330 (N_330,In_961,In_2118);
and U331 (N_331,In_1259,In_1615);
or U332 (N_332,In_2387,In_112);
or U333 (N_333,In_450,In_12);
xor U334 (N_334,In_865,In_2317);
nand U335 (N_335,In_773,In_1708);
and U336 (N_336,In_1750,In_1083);
and U337 (N_337,In_277,In_984);
xor U338 (N_338,In_993,In_1779);
and U339 (N_339,In_1439,In_608);
nand U340 (N_340,In_1722,In_637);
and U341 (N_341,In_1558,In_733);
or U342 (N_342,In_252,In_193);
and U343 (N_343,In_1626,In_38);
nor U344 (N_344,In_248,In_229);
or U345 (N_345,In_791,In_505);
nand U346 (N_346,In_48,In_1124);
xor U347 (N_347,In_1238,In_198);
nand U348 (N_348,In_126,In_1421);
nand U349 (N_349,In_1737,In_1480);
or U350 (N_350,In_1965,In_346);
and U351 (N_351,In_2414,In_1667);
or U352 (N_352,In_2323,In_140);
nand U353 (N_353,In_1994,In_655);
or U354 (N_354,In_1629,In_2110);
xor U355 (N_355,In_362,In_2049);
xor U356 (N_356,In_916,In_428);
nand U357 (N_357,In_1026,In_1870);
and U358 (N_358,In_2042,In_2269);
xor U359 (N_359,In_2176,In_1287);
nand U360 (N_360,In_1931,In_2097);
nor U361 (N_361,In_1449,In_1999);
nand U362 (N_362,In_680,In_2056);
and U363 (N_363,In_1413,In_1933);
xnor U364 (N_364,In_2404,In_1273);
nor U365 (N_365,In_2331,In_2022);
nor U366 (N_366,In_1092,In_2116);
xor U367 (N_367,In_1330,In_242);
xor U368 (N_368,In_141,In_188);
nor U369 (N_369,In_2123,In_929);
xnor U370 (N_370,In_1610,In_2339);
xnor U371 (N_371,In_300,In_649);
nor U372 (N_372,In_1096,In_1494);
nand U373 (N_373,In_2310,In_2445);
nand U374 (N_374,In_2302,In_1618);
or U375 (N_375,In_2366,In_564);
or U376 (N_376,In_2346,In_555);
xnor U377 (N_377,In_668,In_2054);
xor U378 (N_378,In_2380,In_1996);
and U379 (N_379,In_310,In_1248);
nor U380 (N_380,In_1105,In_1757);
xnor U381 (N_381,In_1646,In_1188);
and U382 (N_382,In_715,In_1905);
xnor U383 (N_383,In_1404,In_115);
nor U384 (N_384,In_1019,In_906);
and U385 (N_385,In_1157,In_793);
nor U386 (N_386,In_945,In_1541);
or U387 (N_387,In_1721,In_2487);
xor U388 (N_388,In_45,In_290);
nor U389 (N_389,In_1037,In_1279);
xor U390 (N_390,In_2301,In_977);
nand U391 (N_391,In_2152,In_2232);
or U392 (N_392,In_416,In_2342);
nor U393 (N_393,In_870,In_2140);
nor U394 (N_394,In_2020,In_1844);
nand U395 (N_395,In_2272,In_1251);
and U396 (N_396,In_1894,In_1929);
nor U397 (N_397,In_325,In_2391);
xnor U398 (N_398,In_2151,In_677);
or U399 (N_399,In_1053,In_511);
xor U400 (N_400,In_1348,In_676);
or U401 (N_401,In_1392,In_1584);
nand U402 (N_402,In_2480,In_470);
nand U403 (N_403,In_1241,In_1122);
xor U404 (N_404,In_1682,In_820);
nand U405 (N_405,In_1850,In_407);
and U406 (N_406,In_601,In_213);
and U407 (N_407,In_1372,In_1770);
xnor U408 (N_408,In_736,In_1314);
or U409 (N_409,In_547,In_1199);
nor U410 (N_410,In_1381,In_986);
nor U411 (N_411,In_1321,In_1628);
nand U412 (N_412,In_723,In_254);
nand U413 (N_413,In_2083,In_1379);
xor U414 (N_414,In_449,In_2372);
or U415 (N_415,In_1727,In_97);
nor U416 (N_416,In_176,In_610);
and U417 (N_417,In_1483,In_811);
or U418 (N_418,In_1703,In_1349);
and U419 (N_419,In_21,In_2195);
xor U420 (N_420,In_2287,In_2403);
or U421 (N_421,In_2055,In_2164);
xnor U422 (N_422,In_408,In_170);
or U423 (N_423,In_1482,In_1791);
nand U424 (N_424,In_1410,In_1526);
and U425 (N_425,In_2191,In_1200);
nor U426 (N_426,In_867,In_59);
and U427 (N_427,In_1383,In_2248);
xnor U428 (N_428,In_1764,In_132);
nand U429 (N_429,In_62,In_1254);
or U430 (N_430,In_1133,In_872);
nand U431 (N_431,In_2122,In_1031);
and U432 (N_432,In_2021,In_1213);
and U433 (N_433,In_226,In_1187);
nor U434 (N_434,In_883,In_1186);
xor U435 (N_435,In_57,In_1282);
nand U436 (N_436,In_2418,In_1370);
nand U437 (N_437,In_1555,In_1040);
nor U438 (N_438,In_2001,In_342);
nor U439 (N_439,In_2388,In_538);
nor U440 (N_440,In_1992,In_591);
nand U441 (N_441,In_2266,In_209);
or U442 (N_442,In_343,In_759);
and U443 (N_443,In_771,In_1068);
nand U444 (N_444,In_2050,In_2259);
nor U445 (N_445,In_1909,In_744);
xor U446 (N_446,In_1623,In_1358);
nand U447 (N_447,In_833,In_318);
or U448 (N_448,In_2386,In_1084);
xnor U449 (N_449,In_1514,In_638);
xor U450 (N_450,In_1920,In_463);
or U451 (N_451,In_1268,In_208);
xor U452 (N_452,In_523,In_1464);
or U453 (N_453,In_91,In_861);
nor U454 (N_454,In_1883,In_689);
nor U455 (N_455,In_2285,In_80);
xnor U456 (N_456,In_1866,In_265);
nand U457 (N_457,In_194,In_1987);
and U458 (N_458,In_550,In_297);
and U459 (N_459,In_121,In_1892);
and U460 (N_460,In_1728,In_2273);
or U461 (N_461,In_1885,In_1219);
nand U462 (N_462,In_1237,In_832);
nor U463 (N_463,In_1549,In_2401);
xnor U464 (N_464,In_1361,In_186);
or U465 (N_465,In_997,In_1619);
and U466 (N_466,In_2041,In_786);
xor U467 (N_467,In_1693,In_627);
xnor U468 (N_468,In_175,In_907);
and U469 (N_469,In_423,In_1301);
nand U470 (N_470,In_2461,In_609);
or U471 (N_471,In_109,In_2289);
nor U472 (N_472,In_2007,In_1591);
or U473 (N_473,In_1582,In_1825);
or U474 (N_474,In_2237,In_835);
xnor U475 (N_475,In_1024,In_1252);
xnor U476 (N_476,In_596,In_826);
nor U477 (N_477,In_2370,In_1391);
xnor U478 (N_478,In_1928,In_732);
nor U479 (N_479,In_1567,In_1403);
nand U480 (N_480,In_7,In_1832);
xnor U481 (N_481,In_2048,In_1910);
nor U482 (N_482,In_2136,In_2231);
nor U483 (N_483,In_2307,In_834);
and U484 (N_484,In_1220,In_1008);
or U485 (N_485,In_1005,In_2253);
xnor U486 (N_486,In_1940,In_1);
or U487 (N_487,In_2265,In_1239);
xor U488 (N_488,In_2288,In_857);
or U489 (N_489,In_2452,In_1207);
nand U490 (N_490,In_1528,In_661);
and U491 (N_491,In_1357,In_2218);
and U492 (N_492,In_2023,In_26);
nor U493 (N_493,In_1201,In_2399);
nor U494 (N_494,In_127,In_666);
or U495 (N_495,In_2202,In_159);
nor U496 (N_496,In_1142,In_2106);
nor U497 (N_497,In_1280,In_788);
and U498 (N_498,In_1453,In_1106);
and U499 (N_499,In_1762,In_207);
or U500 (N_500,In_764,In_32);
xor U501 (N_501,In_316,In_667);
nor U502 (N_502,In_1194,In_2484);
and U503 (N_503,In_2137,In_2115);
or U504 (N_504,In_1793,In_1339);
nor U505 (N_505,In_2402,In_1143);
nand U506 (N_506,In_2108,In_949);
nand U507 (N_507,In_1572,In_1596);
or U508 (N_508,In_1644,In_2316);
or U509 (N_509,In_941,In_848);
and U510 (N_510,In_63,In_2348);
or U511 (N_511,In_2300,In_2412);
nor U512 (N_512,In_2303,In_968);
xnor U513 (N_513,In_1374,In_1418);
nand U514 (N_514,In_2149,In_2395);
xnor U515 (N_515,In_1257,In_1649);
or U516 (N_516,In_664,In_1827);
and U517 (N_517,In_602,In_878);
or U518 (N_518,In_1518,In_1137);
and U519 (N_519,In_98,In_967);
and U520 (N_520,In_1539,In_1781);
and U521 (N_521,In_2385,In_772);
xnor U522 (N_522,In_891,In_1424);
and U523 (N_523,In_2204,In_1569);
nor U524 (N_524,In_866,In_150);
xnor U525 (N_525,In_708,In_1621);
xor U526 (N_526,In_1203,In_1602);
and U527 (N_527,In_125,In_699);
xnor U528 (N_528,In_785,In_133);
xor U529 (N_529,In_2291,In_636);
or U530 (N_530,In_1662,In_1302);
and U531 (N_531,In_2463,In_2296);
or U532 (N_532,In_1049,In_1246);
nor U533 (N_533,In_718,In_379);
xnor U534 (N_534,In_323,In_817);
or U535 (N_535,In_1304,In_1484);
and U536 (N_536,In_2471,In_859);
and U537 (N_537,In_2240,In_55);
nand U538 (N_538,In_1645,In_2431);
nor U539 (N_539,In_1723,In_2036);
xor U540 (N_540,In_1415,In_1510);
xnor U541 (N_541,In_2051,In_345);
xor U542 (N_542,In_350,In_2185);
nand U543 (N_543,In_1064,In_1552);
nand U544 (N_544,In_299,In_670);
and U545 (N_545,In_1788,In_420);
and U546 (N_546,In_1078,In_1291);
and U547 (N_547,In_288,In_1586);
and U548 (N_548,In_1647,In_1359);
and U549 (N_549,In_1694,In_1527);
xnor U550 (N_550,In_1669,In_2052);
nor U551 (N_551,In_1258,In_687);
xnor U552 (N_552,In_885,In_74);
xor U553 (N_553,In_1214,In_1921);
xnor U554 (N_554,In_485,In_979);
xor U555 (N_555,In_2311,In_1792);
xnor U556 (N_556,In_2450,In_255);
nor U557 (N_557,In_1384,In_1661);
nor U558 (N_558,In_1263,In_2005);
xnor U559 (N_559,In_1524,In_808);
xor U560 (N_560,In_2095,In_1886);
or U561 (N_561,In_223,In_2345);
or U562 (N_562,In_1197,In_1109);
nand U563 (N_563,In_854,In_1600);
nor U564 (N_564,In_1751,In_707);
xor U565 (N_565,In_110,In_272);
nand U566 (N_566,In_709,In_1365);
nor U567 (N_567,In_964,In_14);
nor U568 (N_568,In_1916,In_1450);
nor U569 (N_569,In_640,In_2242);
nor U570 (N_570,In_2215,In_951);
nor U571 (N_571,In_136,In_622);
nand U572 (N_572,In_2193,In_1590);
or U573 (N_573,In_2201,In_1689);
or U574 (N_574,In_512,In_539);
nand U575 (N_575,In_2436,In_1917);
and U576 (N_576,In_1961,In_935);
nor U577 (N_577,In_395,In_2292);
or U578 (N_578,In_2476,In_674);
nor U579 (N_579,In_934,In_1478);
xor U580 (N_580,In_178,In_1765);
nand U581 (N_581,In_372,In_1664);
or U582 (N_582,In_1098,In_2332);
nand U583 (N_583,In_679,In_2271);
nor U584 (N_584,In_1678,In_1889);
nor U585 (N_585,In_624,In_724);
or U586 (N_586,In_246,In_90);
or U587 (N_587,In_1505,In_892);
xor U588 (N_588,In_2309,In_266);
nand U589 (N_589,In_1430,In_2354);
nand U590 (N_590,In_239,In_490);
nand U591 (N_591,In_1472,In_1030);
xnor U592 (N_592,In_2126,In_371);
and U593 (N_593,In_335,In_483);
nor U594 (N_594,In_10,In_1535);
nand U595 (N_595,In_22,In_2238);
nand U596 (N_596,In_2410,In_2064);
or U597 (N_597,In_475,In_1547);
nand U598 (N_598,In_454,In_920);
nand U599 (N_599,In_748,In_1210);
xor U600 (N_600,In_749,In_1066);
xnor U601 (N_601,In_373,In_2407);
and U602 (N_602,In_232,In_648);
nand U603 (N_603,In_1401,In_684);
or U604 (N_604,In_1546,In_1743);
or U605 (N_605,In_1101,In_845);
xor U606 (N_606,In_1744,In_804);
and U607 (N_607,In_161,In_1074);
nand U608 (N_608,In_659,In_1307);
and U609 (N_609,In_1367,In_116);
or U610 (N_610,In_890,In_860);
and U611 (N_611,In_647,In_151);
nor U612 (N_612,In_1540,In_743);
nand U613 (N_613,In_757,In_1171);
nor U614 (N_614,In_199,In_567);
and U615 (N_615,In_394,In_2214);
nand U616 (N_616,In_641,In_1907);
xnor U617 (N_617,In_2188,In_1852);
or U618 (N_618,In_2375,In_697);
nor U619 (N_619,In_1090,In_1719);
xnor U620 (N_620,In_1512,In_1458);
nor U621 (N_621,In_1395,In_369);
and U622 (N_622,In_593,In_946);
or U623 (N_623,In_1914,In_754);
or U624 (N_624,In_815,In_701);
nand U625 (N_625,In_2182,In_196);
nand U626 (N_626,In_2192,In_2255);
nor U627 (N_627,In_1704,In_1630);
nor U628 (N_628,In_1686,In_768);
or U629 (N_629,In_899,In_1970);
or U630 (N_630,In_1784,In_2015);
nor U631 (N_631,In_1069,In_1981);
xor U632 (N_632,In_2321,In_1303);
nor U633 (N_633,In_1046,In_2090);
nand U634 (N_634,In_102,In_1355);
nor U635 (N_635,In_195,In_243);
and U636 (N_636,In_1576,In_1651);
nor U637 (N_637,In_1501,In_419);
xor U638 (N_638,In_631,In_2290);
nand U639 (N_639,In_1445,In_692);
and U640 (N_640,In_1816,In_1523);
nor U641 (N_641,In_806,In_2489);
nor U642 (N_642,In_2459,In_203);
and U643 (N_643,In_770,In_1761);
xor U644 (N_644,In_1315,In_1934);
or U645 (N_645,In_810,In_802);
nand U646 (N_646,In_1397,In_658);
or U647 (N_647,In_1977,In_2127);
and U648 (N_648,In_1276,In_404);
nand U649 (N_649,In_201,In_584);
nor U650 (N_650,In_738,In_107);
or U651 (N_651,In_2365,In_2058);
nor U652 (N_652,In_838,In_2219);
nand U653 (N_653,In_317,In_2227);
and U654 (N_654,In_740,In_1029);
nand U655 (N_655,In_2197,In_396);
nor U656 (N_656,In_2469,In_1701);
nor U657 (N_657,In_44,In_180);
xor U658 (N_658,In_931,In_190);
nand U659 (N_659,In_2067,In_1834);
and U660 (N_660,In_2465,In_451);
nor U661 (N_661,In_1441,In_2156);
nor U662 (N_662,In_1318,In_893);
or U663 (N_663,In_2038,In_1150);
xor U664 (N_664,In_2408,In_2364);
nand U665 (N_665,In_1944,In_776);
nor U666 (N_666,In_1221,In_1566);
or U667 (N_667,In_1544,In_579);
nand U668 (N_668,In_303,In_830);
nand U669 (N_669,In_1166,In_1670);
and U670 (N_670,In_874,In_619);
nor U671 (N_671,In_2037,In_2236);
xnor U672 (N_672,In_2270,In_625);
nand U673 (N_673,In_862,In_338);
nor U674 (N_674,In_2085,In_987);
nand U675 (N_675,In_913,In_1884);
or U676 (N_676,In_1256,In_825);
and U677 (N_677,In_1145,In_1625);
nor U678 (N_678,In_587,In_1269);
or U679 (N_679,In_1192,In_2035);
or U680 (N_680,In_2194,In_1134);
or U681 (N_681,In_1756,In_595);
or U682 (N_682,In_1659,In_1176);
xor U683 (N_683,In_1695,In_1696);
and U684 (N_684,In_2268,In_1216);
or U685 (N_685,In_1833,In_2184);
or U686 (N_686,In_957,In_1261);
xnor U687 (N_687,In_2153,In_2319);
or U688 (N_688,In_1890,In_2092);
nand U689 (N_689,In_476,In_39);
and U690 (N_690,In_1212,In_432);
and U691 (N_691,In_1278,In_1100);
or U692 (N_692,In_1521,In_51);
nor U693 (N_693,In_1456,In_1663);
nand U694 (N_694,In_1612,In_1730);
and U695 (N_695,In_1429,In_1298);
and U696 (N_696,In_1169,In_2198);
nand U697 (N_697,In_2481,In_2173);
nor U698 (N_698,In_2207,In_2030);
or U699 (N_699,In_286,In_559);
or U700 (N_700,In_1264,In_418);
nand U701 (N_701,In_1255,In_1240);
nor U702 (N_702,In_494,In_367);
xor U703 (N_703,In_1412,In_2249);
xor U704 (N_704,In_562,In_1938);
nor U705 (N_705,In_1735,In_2276);
nand U706 (N_706,In_1432,In_139);
and U707 (N_707,In_1560,In_1095);
xor U708 (N_708,In_1308,In_856);
xnor U709 (N_709,In_1585,In_1352);
nor U710 (N_710,In_876,In_2423);
or U711 (N_711,In_227,In_49);
and U712 (N_712,In_1573,In_2427);
nand U713 (N_713,In_1520,In_747);
nand U714 (N_714,In_2094,In_2263);
xnor U715 (N_715,In_1500,In_273);
or U716 (N_716,In_1006,In_308);
nor U717 (N_717,In_1766,In_1223);
xor U718 (N_718,In_898,In_217);
or U719 (N_719,In_1821,In_1946);
or U720 (N_720,In_537,In_1329);
nor U721 (N_721,In_1754,In_1778);
nor U722 (N_722,In_234,In_1725);
xor U723 (N_723,In_829,In_691);
and U724 (N_724,In_2130,In_2081);
and U725 (N_725,In_1542,In_158);
nor U726 (N_726,In_1749,In_2457);
nor U727 (N_727,In_293,In_1312);
or U728 (N_728,In_1144,In_1958);
xor U729 (N_729,In_282,In_1822);
and U730 (N_730,In_35,In_1986);
or U731 (N_731,In_364,In_2499);
xor U732 (N_732,In_1353,In_1736);
and U733 (N_733,In_1819,In_1217);
and U734 (N_734,In_256,In_370);
nor U735 (N_735,In_54,In_2025);
nor U736 (N_736,In_1091,In_355);
nand U737 (N_737,In_966,In_211);
nor U738 (N_738,In_1323,In_447);
nand U739 (N_739,In_1639,In_644);
xnor U740 (N_740,In_472,In_1974);
nor U741 (N_741,In_819,In_1010);
or U742 (N_742,In_2175,In_1371);
xor U743 (N_743,In_86,In_1447);
and U744 (N_744,In_1481,In_1012);
nand U745 (N_745,In_714,In_17);
nand U746 (N_746,In_1235,In_2061);
and U747 (N_747,In_120,In_2244);
and U748 (N_748,In_1469,In_2029);
xnor U749 (N_749,In_1760,In_2305);
and U750 (N_750,In_2134,In_376);
or U751 (N_751,In_40,In_2133);
nand U752 (N_752,In_6,In_1777);
or U753 (N_753,In_143,In_2091);
or U754 (N_754,In_1745,In_2145);
xor U755 (N_755,In_519,In_553);
nor U756 (N_756,In_85,In_34);
and U757 (N_757,In_549,In_1904);
and U758 (N_758,In_240,In_1003);
nor U759 (N_759,In_2441,In_2121);
nor U760 (N_760,In_1947,In_2053);
or U761 (N_761,In_1613,In_565);
nor U762 (N_762,In_827,In_1378);
nor U763 (N_763,In_96,In_541);
xor U764 (N_764,In_237,In_1369);
nand U765 (N_765,In_82,In_2328);
nor U766 (N_766,In_1604,In_2160);
or U767 (N_767,In_1132,In_1684);
nand U768 (N_768,In_89,In_1668);
nor U769 (N_769,In_1898,In_669);
nor U770 (N_770,In_1136,In_73);
or U771 (N_771,In_2014,In_315);
and U772 (N_772,In_1975,In_481);
nor U773 (N_773,In_1009,In_657);
or U774 (N_774,In_2314,In_250);
or U775 (N_775,In_1603,In_146);
and U776 (N_776,In_2040,In_1274);
or U777 (N_777,In_1164,In_436);
nor U778 (N_778,In_1851,In_259);
or U779 (N_779,In_1517,In_921);
and U780 (N_780,In_2245,In_349);
xor U781 (N_781,In_1004,In_660);
nand U782 (N_782,In_1608,In_313);
nor U783 (N_783,In_1924,In_911);
nor U784 (N_784,In_287,In_1070);
or U785 (N_785,In_84,In_1616);
nand U786 (N_786,In_603,In_937);
xor U787 (N_787,In_1452,In_626);
nand U788 (N_788,In_2315,In_970);
nand U789 (N_789,In_588,In_851);
nand U790 (N_790,In_1588,In_2324);
or U791 (N_791,In_908,In_334);
nand U792 (N_792,In_1285,In_93);
xor U793 (N_793,In_389,In_525);
and U794 (N_794,In_896,In_1802);
nor U795 (N_795,In_8,In_1812);
nand U796 (N_796,In_1813,In_1650);
nand U797 (N_797,In_1637,In_1182);
xor U798 (N_798,In_1899,In_1225);
nor U799 (N_799,In_2477,In_1632);
and U800 (N_800,In_1454,In_1681);
and U801 (N_801,In_1815,In_241);
nand U802 (N_802,In_147,In_1671);
nor U803 (N_803,In_1685,In_735);
nor U804 (N_804,In_2063,In_1861);
xnor U805 (N_805,In_746,In_1631);
nand U806 (N_806,In_544,In_458);
and U807 (N_807,In_2340,In_794);
xnor U808 (N_808,In_1014,In_813);
nor U809 (N_809,In_2313,In_877);
xnor U810 (N_810,In_783,In_888);
nand U811 (N_811,In_662,In_430);
nand U812 (N_812,In_1000,In_2070);
and U813 (N_813,In_465,In_1876);
xnor U814 (N_814,In_1317,In_1679);
xnor U815 (N_815,In_2247,In_577);
nor U816 (N_816,In_1462,In_1305);
nor U817 (N_817,In_1803,In_2349);
nand U818 (N_818,In_1758,In_1882);
xor U819 (N_819,In_905,In_1807);
or U820 (N_820,In_1018,In_1284);
or U821 (N_821,In_270,In_939);
xnor U822 (N_822,In_1504,In_261);
or U823 (N_823,In_763,In_1948);
nor U824 (N_824,In_582,In_33);
or U825 (N_825,In_2158,In_251);
nand U826 (N_826,In_189,In_737);
nand U827 (N_827,In_382,In_742);
nand U828 (N_828,In_336,In_975);
and U829 (N_829,In_1335,In_438);
xor U830 (N_830,In_1218,In_914);
or U831 (N_831,In_1748,In_134);
nor U832 (N_832,In_1039,In_2312);
or U833 (N_833,In_2333,In_822);
and U834 (N_834,In_117,In_618);
nor U835 (N_835,In_443,In_1829);
xor U836 (N_836,In_1923,In_1351);
and U837 (N_837,In_1875,In_1115);
xnor U838 (N_838,In_405,In_1017);
and U839 (N_839,In_2096,In_766);
nand U840 (N_840,In_2211,In_2420);
xor U841 (N_841,In_1161,In_1804);
nand U842 (N_842,In_1102,In_1492);
or U843 (N_843,In_720,In_2181);
nand U844 (N_844,In_144,In_2138);
xnor U845 (N_845,In_4,In_1674);
nand U846 (N_846,In_204,In_157);
nor U847 (N_847,In_1405,In_1473);
and U848 (N_848,In_1783,In_1733);
or U849 (N_849,In_983,In_72);
xor U850 (N_850,In_2079,In_2405);
or U851 (N_851,In_312,In_2146);
nor U852 (N_852,In_1611,In_2298);
xor U853 (N_853,In_2105,In_950);
or U854 (N_854,In_1950,In_2229);
xor U855 (N_855,In_247,In_563);
nand U856 (N_856,In_2167,In_123);
nor U857 (N_857,In_630,In_1343);
xor U858 (N_858,In_1344,In_1860);
nor U859 (N_859,In_148,In_2125);
or U860 (N_860,In_2170,In_2046);
nand U861 (N_861,In_2196,In_281);
or U862 (N_862,In_2367,In_930);
and U863 (N_863,In_612,In_1294);
and U864 (N_864,In_828,In_2396);
nor U865 (N_865,In_1593,In_796);
and U866 (N_866,In_1609,In_1417);
xnor U867 (N_867,In_1763,In_1956);
xor U868 (N_868,In_200,In_298);
nor U869 (N_869,In_1226,In_1859);
or U870 (N_870,In_952,In_790);
nand U871 (N_871,In_542,In_1951);
and U872 (N_872,In_1845,In_1468);
nand U873 (N_873,In_278,In_1643);
nand U874 (N_874,In_2162,In_1536);
nand U875 (N_875,In_683,In_598);
or U876 (N_876,In_375,In_260);
nor U877 (N_877,In_1620,In_322);
nand U878 (N_878,In_1154,In_1895);
xor U879 (N_879,In_1780,In_597);
xor U880 (N_880,In_1849,In_960);
xor U881 (N_881,In_2017,In_154);
or U882 (N_882,In_1129,In_1232);
xnor U883 (N_883,In_1271,In_1300);
nor U884 (N_884,In_1776,In_1117);
nand U885 (N_885,In_2074,In_311);
xnor U886 (N_886,In_2376,In_1949);
xor U887 (N_887,In_948,In_118);
and U888 (N_888,In_2494,In_926);
and U889 (N_889,In_222,In_938);
nand U890 (N_890,In_863,In_340);
nand U891 (N_891,In_1139,In_25);
xnor U892 (N_892,In_1657,In_1409);
xnor U893 (N_893,In_271,In_1364);
nor U894 (N_894,In_2406,In_466);
nor U895 (N_895,In_1288,In_1932);
and U896 (N_896,In_1131,In_690);
nor U897 (N_897,In_153,In_527);
and U898 (N_898,In_875,In_487);
nor U899 (N_899,In_2426,In_1489);
xor U900 (N_900,In_1177,In_283);
nand U901 (N_901,In_540,In_980);
nor U902 (N_902,In_1138,In_530);
nand U903 (N_903,In_1503,In_280);
or U904 (N_904,In_849,In_164);
nand U905 (N_905,In_2306,In_2322);
nor U906 (N_906,In_839,In_2398);
xnor U907 (N_907,In_104,In_1966);
nand U908 (N_908,In_488,In_1159);
or U909 (N_909,In_1688,In_2442);
nand U910 (N_910,In_1879,In_1818);
xnor U911 (N_911,In_446,In_1247);
nor U912 (N_912,In_83,In_696);
or U913 (N_913,In_1640,In_1562);
nand U914 (N_914,In_1598,In_592);
xnor U915 (N_915,In_616,In_2073);
and U916 (N_916,In_1548,In_2413);
nand U917 (N_917,In_1533,In_291);
nand U918 (N_918,In_1297,In_762);
nor U919 (N_919,In_399,In_1675);
nor U920 (N_920,In_138,In_571);
nand U921 (N_921,In_413,In_739);
nand U922 (N_922,In_1824,In_2068);
nand U923 (N_923,In_1702,In_1023);
or U924 (N_924,In_675,In_2147);
nand U925 (N_925,In_103,In_42);
xor U926 (N_926,In_215,In_758);
and U927 (N_927,In_2392,In_606);
or U928 (N_928,In_1642,In_615);
nor U929 (N_929,In_2432,In_2239);
nor U930 (N_930,In_1275,In_427);
and U931 (N_931,In_1769,In_2389);
nand U932 (N_932,In_717,In_1389);
and U933 (N_933,In_2150,In_497);
or U934 (N_934,In_583,In_1328);
xor U935 (N_935,In_841,In_1051);
or U936 (N_936,In_1790,In_64);
nor U937 (N_937,In_9,In_453);
nor U938 (N_938,In_2172,In_1236);
xnor U939 (N_939,In_391,In_678);
xnor U940 (N_940,In_1568,In_1076);
xor U941 (N_941,In_361,In_2482);
and U942 (N_942,In_531,In_1113);
and U943 (N_943,In_331,In_1060);
nor U944 (N_944,In_1382,In_800);
or U945 (N_945,In_1635,In_421);
nor U946 (N_946,In_1050,In_409);
nand U947 (N_947,In_1993,In_1508);
xnor U948 (N_948,In_1457,In_92);
or U949 (N_949,In_514,In_1712);
xor U950 (N_950,In_761,In_917);
and U951 (N_951,In_304,In_2274);
nand U952 (N_952,In_1724,In_152);
or U953 (N_953,In_2117,In_2069);
xnor U954 (N_954,In_1309,In_1706);
and U955 (N_955,In_1658,In_572);
and U956 (N_956,In_1806,In_1652);
nor U957 (N_957,In_947,In_1228);
xor U958 (N_958,In_1011,In_326);
nand U959 (N_959,In_1930,In_1123);
nand U960 (N_960,In_955,In_797);
or U961 (N_961,In_915,In_1887);
nor U962 (N_962,In_1935,In_2233);
nand U963 (N_963,In_1172,In_2098);
xor U964 (N_964,In_780,In_2341);
or U965 (N_965,In_1376,In_192);
or U966 (N_966,In_1127,In_1149);
xor U967 (N_967,In_1511,In_328);
nand U968 (N_968,In_1720,In_900);
nor U969 (N_969,In_1035,In_1167);
and U970 (N_970,In_1493,In_2166);
or U971 (N_971,In_1925,In_1198);
xnor U972 (N_972,In_1191,In_798);
xnor U973 (N_973,In_779,In_1498);
xor U974 (N_974,In_425,In_1195);
nor U975 (N_975,In_1128,In_2102);
nand U976 (N_976,In_1222,In_1848);
xnor U977 (N_977,In_1292,In_2352);
nor U978 (N_978,In_1915,In_1597);
and U979 (N_979,In_1406,In_18);
nand U980 (N_980,In_2326,In_2295);
and U981 (N_981,In_1455,In_1607);
nor U982 (N_982,In_2334,In_351);
nor U983 (N_983,In_53,In_2163);
or U984 (N_984,In_149,In_998);
or U985 (N_985,In_2203,In_923);
xor U986 (N_986,In_580,In_1525);
and U987 (N_987,In_1180,In_1320);
nand U988 (N_988,In_765,In_528);
or U989 (N_989,In_2047,In_1774);
and U990 (N_990,In_1836,In_1025);
and U991 (N_991,In_1927,In_1398);
nand U992 (N_992,In_1390,In_333);
or U993 (N_993,In_1436,In_1311);
nand U994 (N_994,In_1538,In_330);
nor U995 (N_995,In_263,In_130);
xnor U996 (N_996,In_2059,In_46);
nand U997 (N_997,In_2497,In_1911);
xnor U998 (N_998,In_1873,In_520);
or U999 (N_999,In_510,In_2356);
or U1000 (N_1000,In_1919,In_1729);
xnor U1001 (N_1001,N_680,In_1787);
or U1002 (N_1002,In_2308,N_870);
xor U1003 (N_1003,In_285,N_482);
xnor U1004 (N_1004,N_715,N_311);
nand U1005 (N_1005,In_1941,N_577);
or U1006 (N_1006,N_142,N_282);
and U1007 (N_1007,In_1156,N_404);
or U1008 (N_1008,N_745,In_2485);
nor U1009 (N_1009,N_818,In_936);
or U1010 (N_1010,In_2082,In_500);
nand U1011 (N_1011,In_1443,N_182);
nor U1012 (N_1012,In_623,In_2343);
nand U1013 (N_1013,N_733,N_171);
or U1014 (N_1014,N_533,In_1711);
nor U1015 (N_1015,In_1366,N_940);
nand U1016 (N_1016,N_55,N_502);
nand U1017 (N_1017,N_254,N_723);
or U1018 (N_1018,N_514,N_668);
and U1019 (N_1019,N_652,N_248);
and U1020 (N_1020,N_214,In_1687);
nor U1021 (N_1021,N_413,N_679);
nand U1022 (N_1022,N_930,In_1057);
or U1023 (N_1023,N_89,N_356);
nor U1024 (N_1024,N_335,N_503);
or U1025 (N_1025,N_250,N_63);
and U1026 (N_1026,N_763,N_830);
xor U1027 (N_1027,N_505,N_219);
nor U1028 (N_1028,N_168,In_1110);
xor U1029 (N_1029,In_789,In_620);
xnor U1030 (N_1030,N_93,N_865);
nand U1031 (N_1031,N_489,In_576);
or U1032 (N_1032,N_950,N_331);
nor U1033 (N_1033,N_327,N_972);
xor U1034 (N_1034,N_507,N_935);
nand U1035 (N_1035,In_2057,N_963);
nand U1036 (N_1036,N_806,In_1554);
or U1037 (N_1037,In_760,N_57);
and U1038 (N_1038,N_528,In_1753);
xnor U1039 (N_1039,N_585,N_881);
or U1040 (N_1040,N_895,N_589);
and U1041 (N_1041,N_307,In_356);
or U1042 (N_1042,N_395,N_56);
xnor U1043 (N_1043,In_2458,In_182);
or U1044 (N_1044,In_600,N_470);
nor U1045 (N_1045,N_41,In_461);
or U1046 (N_1046,N_179,N_522);
nor U1047 (N_1047,In_1485,N_884);
or U1048 (N_1048,In_1908,N_349);
nand U1049 (N_1049,N_394,N_675);
and U1050 (N_1050,In_2142,N_453);
and U1051 (N_1051,N_261,In_1231);
nand U1052 (N_1052,N_292,N_732);
or U1053 (N_1053,In_1519,N_218);
or U1054 (N_1054,N_31,In_1341);
and U1055 (N_1055,In_2379,In_1922);
xor U1056 (N_1056,In_1578,N_637);
xor U1057 (N_1057,N_405,In_20);
nor U1058 (N_1058,In_903,N_436);
nor U1059 (N_1059,N_88,In_2473);
and U1060 (N_1060,In_2419,N_925);
and U1061 (N_1061,N_676,In_108);
nand U1062 (N_1062,In_1507,In_1130);
or U1063 (N_1063,In_95,N_217);
nor U1064 (N_1064,N_53,N_360);
xor U1065 (N_1065,N_606,N_576);
and U1066 (N_1066,N_775,N_559);
or U1067 (N_1067,In_2453,N_280);
or U1068 (N_1068,In_1281,N_166);
nand U1069 (N_1069,N_875,N_600);
and U1070 (N_1070,In_1565,In_124);
or U1071 (N_1071,In_245,In_2224);
and U1072 (N_1072,In_508,In_268);
and U1073 (N_1073,N_648,N_802);
or U1074 (N_1074,In_1178,N_457);
or U1075 (N_1075,N_419,N_666);
or U1076 (N_1076,N_393,In_632);
or U1077 (N_1077,N_117,N_991);
xnor U1078 (N_1078,N_407,N_17);
nand U1079 (N_1079,In_821,N_302);
nor U1080 (N_1080,N_858,N_980);
nor U1081 (N_1081,N_324,N_534);
xor U1082 (N_1082,N_124,In_2109);
nand U1083 (N_1083,N_660,In_501);
and U1084 (N_1084,N_857,N_662);
or U1085 (N_1085,In_437,In_1299);
nand U1086 (N_1086,In_1148,In_1964);
xor U1087 (N_1087,In_1118,N_276);
xnor U1088 (N_1088,In_1746,N_328);
xor U1089 (N_1089,In_160,N_205);
nor U1090 (N_1090,N_177,In_484);
or U1091 (N_1091,N_60,N_764);
nand U1092 (N_1092,N_24,N_725);
xnor U1093 (N_1093,N_465,N_708);
or U1094 (N_1094,N_125,In_1543);
nand U1095 (N_1095,In_1340,N_661);
nor U1096 (N_1096,N_403,In_1624);
nand U1097 (N_1097,In_1556,N_456);
or U1098 (N_1098,In_363,N_201);
xnor U1099 (N_1099,In_962,N_455);
nand U1100 (N_1100,N_415,In_1387);
nand U1101 (N_1101,In_1747,N_582);
xnor U1102 (N_1102,In_2003,N_224);
and U1103 (N_1103,N_242,N_766);
nor U1104 (N_1104,N_796,N_878);
xnor U1105 (N_1105,N_614,N_946);
xnor U1106 (N_1106,N_230,In_426);
and U1107 (N_1107,In_368,N_401);
nand U1108 (N_1108,In_2178,N_584);
xnor U1109 (N_1109,N_665,In_942);
xnor U1110 (N_1110,N_834,N_195);
or U1111 (N_1111,N_397,In_1550);
nor U1112 (N_1112,N_686,In_621);
or U1113 (N_1113,N_770,N_959);
or U1114 (N_1114,N_718,N_653);
nor U1115 (N_1115,N_226,In_324);
or U1116 (N_1116,In_455,N_181);
nand U1117 (N_1117,N_841,In_1306);
nor U1118 (N_1118,N_549,N_104);
nor U1119 (N_1119,N_808,N_375);
xnor U1120 (N_1120,N_211,N_115);
nand U1121 (N_1121,In_2033,In_533);
xnor U1122 (N_1122,In_1926,N_43);
xnor U1123 (N_1123,N_674,N_444);
xnor U1124 (N_1124,N_535,N_304);
or U1125 (N_1125,N_640,N_377);
and U1126 (N_1126,N_787,N_500);
xor U1127 (N_1127,In_1234,In_2411);
or U1128 (N_1128,N_566,N_259);
nand U1129 (N_1129,N_898,N_267);
nand U1130 (N_1130,N_449,N_847);
nor U1131 (N_1131,In_814,N_748);
or U1132 (N_1132,In_284,N_418);
nor U1133 (N_1133,In_411,N_722);
or U1134 (N_1134,In_2135,In_479);
nor U1135 (N_1135,N_741,N_586);
nor U1136 (N_1136,In_2293,N_294);
and U1137 (N_1137,N_894,N_553);
nor U1138 (N_1138,N_683,N_663);
nor U1139 (N_1139,N_137,N_973);
xnor U1140 (N_1140,N_542,N_918);
xor U1141 (N_1141,N_762,N_938);
xnor U1142 (N_1142,N_23,In_1906);
and U1143 (N_1143,In_2498,N_622);
and U1144 (N_1144,N_59,In_381);
nor U1145 (N_1145,In_47,In_1797);
xor U1146 (N_1146,In_1738,In_489);
or U1147 (N_1147,In_1354,N_703);
nor U1148 (N_1148,In_1289,In_554);
nand U1149 (N_1149,N_684,In_575);
and U1150 (N_1150,N_493,N_420);
xnor U1151 (N_1151,N_599,N_146);
or U1152 (N_1152,N_915,N_739);
and U1153 (N_1153,N_61,In_2371);
or U1154 (N_1154,In_1055,N_701);
nand U1155 (N_1155,N_691,N_610);
nor U1156 (N_1156,N_461,N_620);
nor U1157 (N_1157,N_743,N_844);
or U1158 (N_1158,In_873,N_187);
and U1159 (N_1159,N_234,In_516);
and U1160 (N_1160,N_6,In_1522);
and U1161 (N_1161,N_742,N_220);
nor U1162 (N_1162,In_974,N_91);
nand U1163 (N_1163,N_207,N_162);
xor U1164 (N_1164,In_1653,N_501);
or U1165 (N_1165,In_532,N_800);
nor U1166 (N_1166,N_807,In_1206);
and U1167 (N_1167,In_1420,In_1690);
or U1168 (N_1168,N_283,N_447);
xnor U1169 (N_1169,N_408,N_598);
nand U1170 (N_1170,N_547,N_704);
xor U1171 (N_1171,N_885,N_497);
nand U1172 (N_1172,In_258,In_1868);
nor U1173 (N_1173,N_867,N_68);
nand U1174 (N_1174,N_76,N_445);
xor U1175 (N_1175,N_479,N_351);
xor U1176 (N_1176,N_659,In_1998);
and U1177 (N_1177,N_819,N_944);
nor U1178 (N_1178,In_269,N_651);
and U1179 (N_1179,In_1551,N_823);
and U1180 (N_1180,In_1739,N_848);
nor U1181 (N_1181,In_886,N_908);
xnor U1182 (N_1182,N_917,N_390);
nor U1183 (N_1183,In_521,In_756);
nand U1184 (N_1184,In_2409,In_1606);
nor U1185 (N_1185,N_968,N_82);
nand U1186 (N_1186,N_429,N_111);
nor U1187 (N_1187,N_695,In_573);
or U1188 (N_1188,N_545,N_243);
nand U1189 (N_1189,N_278,In_1843);
xnor U1190 (N_1190,N_359,N_340);
nand U1191 (N_1191,N_520,N_430);
nor U1192 (N_1192,N_962,N_145);
xor U1193 (N_1193,N_655,In_2212);
nor U1194 (N_1194,In_2493,In_943);
or U1195 (N_1195,In_509,N_936);
nand U1196 (N_1196,N_632,N_794);
nor U1197 (N_1197,N_941,In_2250);
xnor U1198 (N_1198,N_425,N_923);
nand U1199 (N_1199,N_212,N_28);
xnor U1200 (N_1200,N_761,N_105);
nor U1201 (N_1201,N_127,N_669);
and U1202 (N_1202,In_1375,N_860);
nor U1203 (N_1203,N_337,In_2424);
xor U1204 (N_1204,N_213,In_2128);
xnor U1205 (N_1205,N_295,N_564);
nor U1206 (N_1206,N_402,N_196);
and U1207 (N_1207,In_1089,In_2474);
or U1208 (N_1208,N_233,N_427);
and U1209 (N_1209,N_880,In_924);
and U1210 (N_1210,In_2353,N_869);
and U1211 (N_1211,N_828,N_624);
and U1212 (N_1212,N_175,N_816);
nand U1213 (N_1213,In_212,N_130);
and U1214 (N_1214,N_814,N_58);
xnor U1215 (N_1215,N_126,N_995);
nand U1216 (N_1216,In_75,N_805);
and U1217 (N_1217,N_116,N_474);
xnor U1218 (N_1218,N_906,N_631);
or U1219 (N_1219,N_799,N_438);
nor U1220 (N_1220,N_133,In_1801);
nand U1221 (N_1221,N_44,N_958);
and U1222 (N_1222,N_529,In_220);
nand U1223 (N_1223,N_713,In_205);
and U1224 (N_1224,N_312,In_1065);
xnor U1225 (N_1225,In_944,In_2087);
and U1226 (N_1226,N_308,N_391);
and U1227 (N_1227,In_990,N_37);
or U1228 (N_1228,N_439,In_1537);
and U1229 (N_1229,N_883,N_341);
nor U1230 (N_1230,N_478,N_149);
nor U1231 (N_1231,N_144,N_772);
nor U1232 (N_1232,In_1676,N_3);
nand U1233 (N_1233,N_778,In_1295);
nor U1234 (N_1234,N_738,In_513);
nor U1235 (N_1235,N_19,N_790);
nand U1236 (N_1236,N_728,N_971);
or U1237 (N_1237,N_231,N_483);
nor U1238 (N_1238,N_709,N_326);
nand U1239 (N_1239,In_1209,In_868);
nand U1240 (N_1240,In_462,N_147);
xnor U1241 (N_1241,In_751,In_1699);
or U1242 (N_1242,In_1121,N_0);
or U1243 (N_1243,N_705,N_605);
nand U1244 (N_1244,In_1250,In_1202);
nand U1245 (N_1245,N_992,N_939);
xnor U1246 (N_1246,N_210,In_163);
or U1247 (N_1247,N_71,N_203);
and U1248 (N_1248,In_1086,In_1509);
or U1249 (N_1249,In_128,N_410);
or U1250 (N_1250,N_275,N_325);
and U1251 (N_1251,N_833,N_50);
and U1252 (N_1252,N_384,N_638);
xor U1253 (N_1253,N_10,In_181);
and U1254 (N_1254,N_911,In_352);
nand U1255 (N_1255,In_1856,N_376);
or U1256 (N_1256,N_97,In_617);
xnor U1257 (N_1257,N_531,In_1942);
and U1258 (N_1258,N_942,N_480);
xor U1259 (N_1259,In_672,N_876);
nand U1260 (N_1260,N_897,In_1575);
or U1261 (N_1261,N_381,In_253);
nand U1262 (N_1262,N_993,In_645);
xor U1263 (N_1263,N_313,N_716);
xnor U1264 (N_1264,N_850,N_970);
nor U1265 (N_1265,N_774,N_400);
or U1266 (N_1266,In_156,N_256);
xnor U1267 (N_1267,In_710,In_36);
or U1268 (N_1268,N_488,N_277);
xnor U1269 (N_1269,N_21,N_52);
or U1270 (N_1270,N_154,N_252);
or U1271 (N_1271,In_1796,N_462);
nor U1272 (N_1272,N_815,N_654);
nand U1273 (N_1273,N_297,In_210);
xor U1274 (N_1274,In_1742,In_614);
nor U1275 (N_1275,In_1969,N_90);
xnor U1276 (N_1276,N_128,N_273);
nor U1277 (N_1277,N_927,N_39);
or U1278 (N_1278,N_639,In_1388);
nand U1279 (N_1279,N_172,In_1477);
and U1280 (N_1280,N_609,N_532);
nand U1281 (N_1281,N_15,N_481);
nor U1282 (N_1282,In_76,In_2199);
nor U1283 (N_1283,In_1322,N_650);
or U1284 (N_1284,N_689,N_26);
and U1285 (N_1285,In_1656,N_904);
nand U1286 (N_1286,N_229,N_697);
or U1287 (N_1287,N_47,N_69);
xnor U1288 (N_1288,N_344,N_386);
nor U1289 (N_1289,N_372,In_467);
or U1290 (N_1290,N_690,In_652);
nor U1291 (N_1291,In_417,In_1422);
and U1292 (N_1292,In_31,In_1408);
or U1293 (N_1293,N_682,N_392);
nor U1294 (N_1294,N_952,N_924);
nand U1295 (N_1295,N_781,In_184);
nand U1296 (N_1296,In_1045,N_804);
xnor U1297 (N_1297,N_72,In_1865);
nor U1298 (N_1298,N_471,In_1984);
or U1299 (N_1299,N_842,N_373);
nor U1300 (N_1300,N_817,In_1789);
and U1301 (N_1301,N_931,N_839);
and U1302 (N_1302,N_746,In_2327);
nor U1303 (N_1303,N_62,N_266);
nand U1304 (N_1304,In_236,In_2454);
or U1305 (N_1305,N_306,In_560);
nand U1306 (N_1306,In_831,N_621);
nand U1307 (N_1307,N_247,In_918);
and U1308 (N_1308,N_253,In_1633);
xnor U1309 (N_1309,In_673,In_1901);
nor U1310 (N_1310,In_2435,N_7);
nand U1311 (N_1311,N_657,N_587);
nor U1312 (N_1312,In_719,In_52);
nor U1313 (N_1313,N_720,In_1718);
xor U1314 (N_1314,In_2032,N_310);
nor U1315 (N_1315,N_274,N_121);
nor U1316 (N_1316,N_699,N_102);
nand U1317 (N_1317,N_710,N_527);
nand U1318 (N_1318,N_824,In_2104);
or U1319 (N_1319,N_996,N_131);
nand U1320 (N_1320,N_362,N_953);
nor U1321 (N_1321,N_518,In_295);
and U1322 (N_1322,N_74,N_204);
xor U1323 (N_1323,In_2397,N_871);
and U1324 (N_1324,N_106,In_1140);
or U1325 (N_1325,N_290,N_751);
nand U1326 (N_1326,In_78,N_590);
or U1327 (N_1327,N_571,In_2361);
nor U1328 (N_1328,N_949,In_994);
xnor U1329 (N_1329,In_2462,N_696);
and U1330 (N_1330,In_155,N_524);
xnor U1331 (N_1331,N_174,N_698);
nor U1332 (N_1332,N_836,In_976);
xor U1333 (N_1333,In_1660,In_2337);
and U1334 (N_1334,N_989,N_693);
nor U1335 (N_1335,In_1184,In_1347);
and U1336 (N_1336,N_148,In_901);
or U1337 (N_1337,N_13,N_86);
nor U1338 (N_1338,N_694,N_183);
nor U1339 (N_1339,In_2446,N_647);
xor U1340 (N_1340,N_985,N_873);
nand U1341 (N_1341,N_581,In_71);
and U1342 (N_1342,In_1063,N_951);
and U1343 (N_1343,N_442,N_160);
or U1344 (N_1344,N_299,In_1465);
nand U1345 (N_1345,In_2026,N_73);
and U1346 (N_1346,N_123,N_910);
or U1347 (N_1347,In_1079,N_730);
or U1348 (N_1348,N_150,In_2440);
xnor U1349 (N_1349,N_687,N_99);
nor U1350 (N_1350,N_494,N_626);
xnor U1351 (N_1351,N_630,N_492);
xnor U1352 (N_1352,N_998,N_336);
and U1353 (N_1353,N_246,N_664);
nor U1354 (N_1354,N_646,N_849);
nor U1355 (N_1355,In_2430,In_2077);
and U1356 (N_1356,N_486,N_792);
nand U1357 (N_1357,In_2443,In_965);
and U1358 (N_1358,N_672,In_629);
xor U1359 (N_1359,N_540,In_1516);
or U1360 (N_1360,N_932,N_974);
and U1361 (N_1361,N_530,N_42);
or U1362 (N_1362,In_1135,In_1444);
nor U1363 (N_1363,N_645,N_677);
or U1364 (N_1364,In_843,N_617);
nor U1365 (N_1365,N_263,N_9);
nand U1366 (N_1366,In_2488,N_338);
nor U1367 (N_1367,N_382,In_1190);
and U1368 (N_1368,N_426,N_827);
and U1369 (N_1369,In_2429,N_608);
or U1370 (N_1370,N_987,N_719);
nor U1371 (N_1371,In_971,In_2155);
nor U1372 (N_1372,N_550,In_2304);
nand U1373 (N_1373,N_788,N_907);
or U1374 (N_1374,In_174,In_1097);
nor U1375 (N_1375,In_2456,N_451);
nand U1376 (N_1376,N_346,In_11);
or U1377 (N_1377,In_50,N_364);
nor U1378 (N_1378,N_232,In_2490);
and U1379 (N_1379,N_159,N_70);
nor U1380 (N_1380,N_752,N_191);
xnor U1381 (N_1381,In_1476,In_402);
or U1382 (N_1382,N_832,In_302);
or U1383 (N_1383,In_101,N_431);
or U1384 (N_1384,In_1799,In_306);
nand U1385 (N_1385,N_291,N_943);
nand U1386 (N_1386,N_411,N_78);
nand U1387 (N_1387,N_756,N_811);
and U1388 (N_1388,N_113,N_563);
or U1389 (N_1389,N_579,N_475);
or U1390 (N_1390,N_846,N_433);
and U1391 (N_1391,N_285,N_38);
xnor U1392 (N_1392,In_799,N_797);
and U1393 (N_1393,In_2467,N_558);
or U1394 (N_1394,N_65,N_982);
nand U1395 (N_1395,N_750,N_122);
nor U1396 (N_1396,N_463,In_1713);
or U1397 (N_1397,N_443,N_414);
nor U1398 (N_1398,In_953,N_574);
xor U1399 (N_1399,N_84,N_859);
nand U1400 (N_1400,N_656,In_79);
and U1401 (N_1401,N_268,N_678);
xor U1402 (N_1402,N_198,N_416);
and U1403 (N_1403,In_1175,N_671);
or U1404 (N_1404,In_1325,N_618);
nand U1405 (N_1405,N_421,In_706);
nand U1406 (N_1406,In_777,N_813);
xnor U1407 (N_1407,N_25,N_706);
and U1408 (N_1408,N_966,N_322);
nand U1409 (N_1409,In_1400,N_464);
nand U1410 (N_1410,N_926,N_525);
or U1411 (N_1411,N_902,In_129);
or U1412 (N_1412,N_899,In_1386);
xor U1413 (N_1413,In_1459,In_2144);
xor U1414 (N_1414,N_851,In_503);
nor U1415 (N_1415,N_777,N_731);
nand U1416 (N_1416,N_649,In_2226);
and U1417 (N_1417,N_472,N_353);
nor U1418 (N_1418,N_20,In_2);
nand U1419 (N_1419,N_87,N_184);
nor U1420 (N_1420,In_1506,In_2320);
xnor U1421 (N_1421,In_1072,In_922);
xnor U1422 (N_1422,N_446,N_546);
nor U1423 (N_1423,In_1692,In_1772);
nor U1424 (N_1424,N_153,N_890);
xor U1425 (N_1425,N_644,N_235);
nand U1426 (N_1426,N_629,N_193);
nor U1427 (N_1427,N_485,N_216);
and U1428 (N_1428,In_904,In_1855);
xor U1429 (N_1429,N_837,N_983);
nor U1430 (N_1430,N_947,N_977);
or U1431 (N_1431,N_979,N_448);
nand U1432 (N_1432,In_2220,N_434);
xnor U1433 (N_1433,N_332,N_151);
or U1434 (N_1434,In_1316,N_602);
and U1435 (N_1435,In_452,In_2060);
nor U1436 (N_1436,In_68,N_134);
or U1437 (N_1437,N_901,N_109);
xor U1438 (N_1438,N_999,N_27);
and U1439 (N_1439,N_36,In_682);
xor U1440 (N_1440,In_1058,In_1260);
and U1441 (N_1441,In_1474,N_262);
nor U1442 (N_1442,N_754,N_826);
nor U1443 (N_1443,N_281,N_30);
and U1444 (N_1444,N_929,N_737);
nor U1445 (N_1445,N_424,N_496);
xnor U1446 (N_1446,In_2350,In_1838);
or U1447 (N_1447,In_1785,N_724);
and U1448 (N_1448,N_258,In_2141);
and U1449 (N_1449,In_2359,N_868);
nand U1450 (N_1450,In_858,N_484);
nor U1451 (N_1451,In_2169,N_192);
or U1452 (N_1452,N_810,N_592);
and U1453 (N_1453,N_173,In_1435);
nor U1454 (N_1454,N_539,N_239);
xor U1455 (N_1455,In_1826,In_2374);
nor U1456 (N_1456,In_932,N_785);
and U1457 (N_1457,In_517,N_238);
nand U1458 (N_1458,N_613,In_414);
nand U1459 (N_1459,N_368,N_757);
and U1460 (N_1460,N_357,In_2216);
nand U1461 (N_1461,N_206,N_358);
nand U1462 (N_1462,N_717,N_997);
nand U1463 (N_1463,N_903,N_760);
or U1464 (N_1464,N_627,N_625);
and U1465 (N_1465,N_264,In_43);
nand U1466 (N_1466,N_843,In_493);
xor U1467 (N_1467,In_2080,N_567);
nand U1468 (N_1468,In_1957,N_721);
xnor U1469 (N_1469,In_2475,N_396);
or U1470 (N_1470,In_177,In_910);
nor U1471 (N_1471,N_367,N_370);
nand U1472 (N_1472,N_565,N_948);
and U1473 (N_1473,N_5,N_912);
xor U1474 (N_1474,N_170,N_94);
xor U1475 (N_1475,In_457,In_1442);
nor U1476 (N_1476,N_2,N_132);
and U1477 (N_1477,N_852,In_1771);
nand U1478 (N_1478,N_92,N_383);
nand U1479 (N_1479,N_960,N_167);
or U1480 (N_1480,N_369,N_101);
and U1481 (N_1481,N_176,N_286);
nand U1482 (N_1482,N_284,N_225);
nor U1483 (N_1483,N_45,N_891);
or U1484 (N_1484,In_397,N_40);
and U1485 (N_1485,N_874,In_403);
nor U1486 (N_1486,N_783,In_1174);
nand U1487 (N_1487,N_33,N_18);
and U1488 (N_1488,N_459,N_378);
nor U1489 (N_1489,N_673,N_380);
xor U1490 (N_1490,N_921,In_752);
and U1491 (N_1491,In_2329,N_296);
nand U1492 (N_1492,N_506,N_441);
nand U1493 (N_1493,N_521,N_188);
and U1494 (N_1494,In_1224,In_206);
nand U1495 (N_1495,In_374,In_228);
nand U1496 (N_1496,N_569,In_681);
nor U1497 (N_1497,N_861,In_1267);
xor U1498 (N_1498,N_333,N_562);
or U1499 (N_1499,N_628,N_315);
or U1500 (N_1500,N_347,N_793);
and U1501 (N_1501,In_202,N_773);
and U1502 (N_1502,N_812,In_1918);
nand U1503 (N_1503,N_765,N_161);
and U1504 (N_1504,In_504,In_846);
nand U1505 (N_1505,N_305,N_854);
or U1506 (N_1506,N_825,In_1346);
and U1507 (N_1507,N_700,In_480);
nand U1508 (N_1508,N_244,N_707);
and U1509 (N_1509,N_301,N_555);
or U1510 (N_1510,In_650,N_964);
xor U1511 (N_1511,In_1954,N_11);
nand U1512 (N_1512,N_12,In_3);
nor U1513 (N_1513,N_409,N_279);
and U1514 (N_1514,In_2200,N_975);
nand U1515 (N_1515,N_893,N_821);
nor U1516 (N_1516,N_399,N_388);
nor U1517 (N_1517,N_537,N_499);
and U1518 (N_1518,In_2336,N_919);
nand U1519 (N_1519,N_711,N_965);
xor U1520 (N_1520,In_842,N_541);
and U1521 (N_1521,N_398,N_318);
xnor U1522 (N_1522,N_164,N_510);
or U1523 (N_1523,In_1061,In_1677);
xnor U1524 (N_1524,In_65,N_79);
nand U1525 (N_1525,In_2187,N_237);
or U1526 (N_1526,N_596,In_1817);
nand U1527 (N_1527,N_118,N_75);
nand U1528 (N_1528,In_887,N_136);
nor U1529 (N_1529,In_847,N_108);
and U1530 (N_1530,N_379,N_343);
or U1531 (N_1531,N_241,N_498);
xor U1532 (N_1532,N_512,N_432);
nor U1533 (N_1533,N_119,N_791);
or U1534 (N_1534,N_469,N_270);
and U1535 (N_1535,N_594,N_490);
nand U1536 (N_1536,In_604,In_716);
nand U1537 (N_1537,N_64,N_753);
nor U1538 (N_1538,In_1775,N_491);
xnor U1539 (N_1539,In_1741,N_120);
nand U1540 (N_1540,N_504,N_374);
or U1541 (N_1541,N_957,N_578);
nor U1542 (N_1542,N_920,N_667);
or U1543 (N_1543,In_2180,In_2416);
xnor U1544 (N_1544,N_889,N_352);
or U1545 (N_1545,N_34,In_264);
or U1546 (N_1546,N_990,N_112);
nand U1547 (N_1547,N_354,N_508);
xnor U1548 (N_1548,N_905,N_779);
or U1549 (N_1549,N_152,N_536);
xor U1550 (N_1550,N_615,N_984);
nand U1551 (N_1551,N_477,N_257);
and U1552 (N_1552,N_864,In_634);
and U1553 (N_1553,N_769,N_417);
and U1554 (N_1554,N_155,N_886);
or U1555 (N_1555,N_560,N_702);
or U1556 (N_1556,In_2283,In_2438);
and U1557 (N_1557,N_509,In_1463);
or U1558 (N_1558,N_887,N_994);
and U1559 (N_1559,In_1862,In_522);
nand U1560 (N_1560,In_1985,In_1327);
or U1561 (N_1561,N_937,In_1622);
xor U1562 (N_1562,N_557,In_2161);
or U1563 (N_1563,N_473,N_4);
and U1564 (N_1564,In_956,In_1360);
nor U1565 (N_1565,In_2148,N_298);
xnor U1566 (N_1566,N_517,N_129);
nor U1567 (N_1567,N_616,In_244);
xor U1568 (N_1568,In_2223,N_208);
and U1569 (N_1569,In_386,N_820);
or U1570 (N_1570,In_401,N_223);
xor U1571 (N_1571,N_289,N_892);
xnor U1572 (N_1572,N_759,N_423);
nor U1573 (N_1573,N_387,N_323);
xor U1574 (N_1574,N_789,N_978);
and U1575 (N_1575,In_2065,N_107);
nor U1576 (N_1576,N_85,In_1553);
and U1577 (N_1577,N_180,N_139);
nor U1578 (N_1578,N_366,N_872);
and U1579 (N_1579,In_2433,N_611);
nand U1580 (N_1580,N_169,In_928);
and U1581 (N_1581,N_245,N_227);
nor U1582 (N_1582,N_251,N_8);
and U1583 (N_1583,N_350,In_2447);
xor U1584 (N_1584,N_138,N_319);
nor U1585 (N_1585,N_476,N_185);
and U1586 (N_1586,In_722,N_228);
or U1587 (N_1587,N_636,In_1902);
xor U1588 (N_1588,In_2099,In_1952);
or U1589 (N_1589,N_782,N_1);
and U1590 (N_1590,N_685,N_729);
or U1591 (N_1591,In_2131,N_260);
nand U1592 (N_1592,In_1163,N_141);
nor U1593 (N_1593,N_986,N_389);
nand U1594 (N_1594,In_70,N_588);
and U1595 (N_1595,N_747,N_736);
nand U1596 (N_1596,N_726,N_240);
and U1597 (N_1597,N_543,N_856);
nand U1598 (N_1598,N_922,N_961);
or U1599 (N_1599,In_319,N_32);
or U1600 (N_1600,In_1208,N_516);
or U1601 (N_1601,N_361,In_1594);
nand U1602 (N_1602,In_1854,In_570);
nor U1603 (N_1603,In_460,N_422);
nand U1604 (N_1604,In_1114,N_916);
and U1605 (N_1605,In_235,N_976);
and U1606 (N_1606,N_450,In_1872);
and U1607 (N_1607,N_822,N_412);
and U1608 (N_1608,N_428,N_16);
nand U1609 (N_1609,N_293,In_2100);
nand U1610 (N_1610,N_303,N_339);
or U1611 (N_1611,N_801,In_5);
and U1612 (N_1612,N_853,In_1595);
nor U1613 (N_1613,N_272,In_1968);
nor U1614 (N_1614,In_882,In_105);
or U1615 (N_1615,N_454,N_48);
or U1616 (N_1616,In_2230,N_573);
nand U1617 (N_1617,In_712,N_321);
nor U1618 (N_1618,In_383,N_780);
and U1619 (N_1619,In_1891,N_271);
nor U1620 (N_1620,N_744,In_1245);
xnor U1621 (N_1621,In_506,In_307);
and U1622 (N_1622,N_755,N_934);
and U1623 (N_1623,N_269,In_518);
or U1624 (N_1624,N_334,In_1146);
xnor U1625 (N_1625,In_1767,N_515);
nand U1626 (N_1626,N_209,N_688);
nand U1627 (N_1627,N_163,In_1048);
and U1628 (N_1628,N_593,N_236);
or U1629 (N_1629,N_795,In_2221);
nor U1630 (N_1630,N_607,N_882);
nor U1631 (N_1631,In_1828,In_1411);
nand U1632 (N_1632,In_410,In_2260);
and U1633 (N_1633,N_371,N_329);
nand U1634 (N_1634,N_523,N_29);
nor U1635 (N_1635,N_727,N_194);
nand U1636 (N_1636,In_1080,In_2209);
nor U1637 (N_1637,N_642,N_288);
xor U1638 (N_1638,In_1233,N_855);
or U1639 (N_1639,N_956,N_435);
or U1640 (N_1640,In_400,N_158);
nand U1641 (N_1641,In_1869,N_135);
and U1642 (N_1642,N_95,N_554);
xor U1643 (N_1643,N_967,N_156);
and U1644 (N_1644,In_2394,In_171);
and U1645 (N_1645,In_1937,N_143);
or U1646 (N_1646,N_14,N_635);
xor U1647 (N_1647,N_348,N_487);
nor U1648 (N_1648,N_829,In_529);
or U1649 (N_1649,N_98,N_603);
xor U1650 (N_1650,N_49,N_863);
nor U1651 (N_1651,N_575,N_255);
nand U1652 (N_1652,N_561,N_749);
xor U1653 (N_1653,In_803,N_643);
xnor U1654 (N_1654,N_634,In_2132);
nand U1655 (N_1655,N_385,N_316);
nand U1656 (N_1656,In_642,In_507);
nand U1657 (N_1657,N_466,In_1193);
nor U1658 (N_1658,N_513,N_317);
and U1659 (N_1659,N_314,N_767);
nand U1660 (N_1660,N_96,N_467);
and U1661 (N_1661,In_1973,N_670);
and U1662 (N_1662,N_157,N_583);
nor U1663 (N_1663,N_189,N_345);
xnor U1664 (N_1664,N_202,N_437);
nand U1665 (N_1665,In_329,N_879);
nor U1666 (N_1666,N_758,In_1574);
or U1667 (N_1667,In_1428,N_110);
nor U1668 (N_1668,N_580,N_913);
and U1669 (N_1669,N_46,In_1665);
nand U1670 (N_1670,N_77,N_572);
nor U1671 (N_1671,N_838,N_845);
xor U1672 (N_1672,N_835,N_199);
xnor U1673 (N_1673,In_1385,N_734);
or U1674 (N_1674,N_249,N_771);
nand U1675 (N_1675,In_1270,In_415);
and U1676 (N_1676,N_570,N_365);
nor U1677 (N_1677,N_798,N_681);
nor U1678 (N_1678,N_165,In_41);
and U1679 (N_1679,N_735,N_103);
nor U1680 (N_1680,N_265,N_197);
or U1681 (N_1681,In_172,In_456);
and U1682 (N_1682,N_551,In_233);
nor U1683 (N_1683,N_215,N_330);
nor U1684 (N_1684,N_954,N_320);
or U1685 (N_1685,In_1858,N_190);
nor U1686 (N_1686,N_22,In_166);
nand U1687 (N_1687,N_309,N_928);
nor U1688 (N_1688,In_1495,In_1995);
xor U1689 (N_1689,N_300,In_2358);
xnor U1690 (N_1690,N_862,N_81);
xnor U1691 (N_1691,In_477,N_633);
or U1692 (N_1692,N_831,N_552);
nand U1693 (N_1693,In_2492,In_1638);
nor U1694 (N_1694,In_77,N_914);
nand U1695 (N_1695,In_2213,N_460);
xor U1696 (N_1696,N_612,N_988);
nand U1697 (N_1697,N_740,In_581);
nor U1698 (N_1698,N_595,In_812);
xor U1699 (N_1699,N_114,N_981);
nor U1700 (N_1700,N_548,N_619);
and U1701 (N_1701,N_80,N_786);
nor U1702 (N_1702,In_646,In_2089);
or U1703 (N_1703,N_955,In_721);
or U1704 (N_1704,N_363,N_840);
and U1705 (N_1705,In_498,In_1531);
or U1706 (N_1706,N_140,In_1491);
nor U1707 (N_1707,N_526,N_495);
nand U1708 (N_1708,N_287,N_784);
nor U1709 (N_1709,N_452,In_2451);
xor U1710 (N_1710,N_67,N_623);
nand U1711 (N_1711,N_66,N_100);
and U1712 (N_1712,In_327,N_809);
and U1713 (N_1713,N_714,N_342);
or U1714 (N_1714,N_468,In_1990);
xnor U1715 (N_1715,In_28,N_877);
xor U1716 (N_1716,In_2139,N_604);
and U1717 (N_1717,In_365,N_712);
nor U1718 (N_1718,In_1529,N_969);
nor U1719 (N_1719,In_1601,N_458);
nor U1720 (N_1720,N_597,In_824);
and U1721 (N_1721,In_1244,In_1362);
xnor U1722 (N_1722,N_83,In_1179);
nor U1723 (N_1723,In_2043,In_1047);
nand U1724 (N_1724,N_692,N_945);
or U1725 (N_1725,N_355,N_406);
xor U1726 (N_1726,N_35,N_568);
nand U1727 (N_1727,N_601,N_54);
xnor U1728 (N_1728,In_2363,N_888);
nand U1729 (N_1729,N_803,In_613);
or U1730 (N_1730,N_556,N_221);
or U1731 (N_1731,In_1054,In_1786);
xor U1732 (N_1732,N_591,N_909);
and U1733 (N_1733,N_519,In_543);
and U1734 (N_1734,In_1326,N_900);
nand U1735 (N_1735,N_538,N_641);
nor U1736 (N_1736,In_2294,In_187);
or U1737 (N_1737,N_933,In_113);
xnor U1738 (N_1738,N_200,N_896);
nand U1739 (N_1739,N_776,N_440);
nor U1740 (N_1740,In_782,In_496);
or U1741 (N_1741,N_511,In_2018);
or U1742 (N_1742,N_51,In_2045);
or U1743 (N_1743,In_221,N_186);
xnor U1744 (N_1744,N_178,In_823);
nor U1745 (N_1745,In_424,In_745);
and U1746 (N_1746,In_1881,N_544);
nor U1747 (N_1747,In_2377,In_611);
xnor U1748 (N_1748,N_658,N_768);
xor U1749 (N_1749,N_222,N_866);
nand U1750 (N_1750,In_352,N_378);
and U1751 (N_1751,N_477,In_513);
nand U1752 (N_1752,In_365,In_2416);
nand U1753 (N_1753,In_2492,N_854);
and U1754 (N_1754,N_537,N_543);
nand U1755 (N_1755,In_1174,In_681);
and U1756 (N_1756,In_212,N_552);
nor U1757 (N_1757,N_253,N_653);
nand U1758 (N_1758,N_320,N_609);
nand U1759 (N_1759,N_147,N_566);
nand U1760 (N_1760,N_834,In_814);
nand U1761 (N_1761,In_922,N_890);
and U1762 (N_1762,In_706,In_1140);
xor U1763 (N_1763,In_1718,N_125);
xor U1764 (N_1764,N_83,N_397);
or U1765 (N_1765,N_130,N_243);
or U1766 (N_1766,N_924,In_411);
or U1767 (N_1767,In_129,N_211);
nand U1768 (N_1768,In_71,In_823);
nand U1769 (N_1769,N_649,N_822);
nand U1770 (N_1770,In_503,N_62);
and U1771 (N_1771,In_302,In_2474);
nand U1772 (N_1772,In_506,N_685);
or U1773 (N_1773,N_300,N_228);
or U1774 (N_1774,In_1435,N_970);
nor U1775 (N_1775,N_806,In_417);
nand U1776 (N_1776,N_658,N_975);
xnor U1777 (N_1777,In_496,N_664);
xor U1778 (N_1778,N_394,N_923);
or U1779 (N_1779,In_533,N_243);
and U1780 (N_1780,N_224,N_927);
xor U1781 (N_1781,N_962,In_1692);
nor U1782 (N_1782,N_106,N_825);
nand U1783 (N_1783,N_706,In_1065);
nand U1784 (N_1784,N_445,N_350);
nor U1785 (N_1785,N_272,In_1420);
xnor U1786 (N_1786,N_49,N_624);
xnor U1787 (N_1787,N_493,N_12);
nor U1788 (N_1788,N_487,N_491);
and U1789 (N_1789,N_530,N_196);
nor U1790 (N_1790,N_377,In_1843);
nand U1791 (N_1791,In_1908,In_1208);
and U1792 (N_1792,In_799,N_678);
nand U1793 (N_1793,N_75,In_324);
and U1794 (N_1794,In_1638,N_335);
and U1795 (N_1795,In_2142,In_1148);
nand U1796 (N_1796,N_350,In_50);
xnor U1797 (N_1797,N_671,In_460);
nor U1798 (N_1798,N_957,N_272);
or U1799 (N_1799,N_205,N_374);
and U1800 (N_1800,N_880,N_361);
nor U1801 (N_1801,N_762,In_521);
or U1802 (N_1802,N_505,N_126);
nand U1803 (N_1803,N_205,N_579);
nand U1804 (N_1804,N_879,N_709);
and U1805 (N_1805,N_780,N_124);
and U1806 (N_1806,N_747,N_208);
and U1807 (N_1807,In_498,N_582);
or U1808 (N_1808,N_683,N_33);
nand U1809 (N_1809,N_675,N_10);
or U1810 (N_1810,In_1459,In_629);
or U1811 (N_1811,In_2350,In_484);
xor U1812 (N_1812,N_94,N_329);
and U1813 (N_1813,In_2082,N_0);
or U1814 (N_1814,N_300,In_264);
or U1815 (N_1815,N_769,N_345);
xor U1816 (N_1816,In_1985,N_189);
xor U1817 (N_1817,N_385,In_2180);
nand U1818 (N_1818,In_706,N_494);
or U1819 (N_1819,In_1594,N_948);
xor U1820 (N_1820,N_282,N_725);
and U1821 (N_1821,N_235,N_816);
nand U1822 (N_1822,N_741,In_1118);
or U1823 (N_1823,In_943,N_848);
and U1824 (N_1824,N_113,N_283);
xor U1825 (N_1825,N_74,N_348);
nor U1826 (N_1826,In_1190,N_838);
nor U1827 (N_1827,N_857,N_230);
nand U1828 (N_1828,N_171,N_802);
xnor U1829 (N_1829,In_1375,N_133);
and U1830 (N_1830,N_902,N_717);
and U1831 (N_1831,N_764,N_186);
xnor U1832 (N_1832,N_643,N_159);
nor U1833 (N_1833,N_515,In_2260);
and U1834 (N_1834,N_431,N_639);
and U1835 (N_1835,In_206,In_2294);
xor U1836 (N_1836,In_1476,N_404);
and U1837 (N_1837,N_961,N_465);
or U1838 (N_1838,In_2141,In_386);
or U1839 (N_1839,N_741,N_550);
nand U1840 (N_1840,N_668,In_1346);
nor U1841 (N_1841,In_212,N_134);
xor U1842 (N_1842,N_601,In_1676);
nor U1843 (N_1843,In_228,In_1746);
nor U1844 (N_1844,In_1202,N_431);
nand U1845 (N_1845,In_1786,N_726);
nand U1846 (N_1846,N_23,N_800);
nand U1847 (N_1847,N_59,In_2178);
or U1848 (N_1848,In_506,N_410);
nor U1849 (N_1849,N_829,N_186);
xor U1850 (N_1850,N_559,N_42);
xor U1851 (N_1851,N_964,N_322);
or U1852 (N_1852,In_1624,In_604);
xnor U1853 (N_1853,N_531,N_205);
nor U1854 (N_1854,In_1865,N_372);
nand U1855 (N_1855,N_49,N_741);
xor U1856 (N_1856,In_253,In_1529);
and U1857 (N_1857,N_6,In_521);
and U1858 (N_1858,N_361,N_802);
xor U1859 (N_1859,N_367,In_306);
and U1860 (N_1860,N_950,N_846);
nand U1861 (N_1861,N_325,In_634);
or U1862 (N_1862,N_152,In_1184);
xnor U1863 (N_1863,N_66,In_295);
or U1864 (N_1864,N_652,N_388);
xnor U1865 (N_1865,N_153,N_957);
or U1866 (N_1866,In_2336,In_171);
and U1867 (N_1867,N_726,N_860);
and U1868 (N_1868,N_303,N_47);
nand U1869 (N_1869,N_268,N_765);
and U1870 (N_1870,N_801,N_625);
xnor U1871 (N_1871,N_946,N_750);
or U1872 (N_1872,N_793,In_507);
or U1873 (N_1873,In_1665,N_943);
nor U1874 (N_1874,N_772,N_369);
and U1875 (N_1875,N_601,In_521);
and U1876 (N_1876,N_974,In_1656);
and U1877 (N_1877,N_369,In_1881);
nor U1878 (N_1878,N_236,N_122);
nor U1879 (N_1879,N_677,N_320);
nor U1880 (N_1880,N_959,N_908);
and U1881 (N_1881,N_760,N_990);
xnor U1882 (N_1882,N_808,In_11);
nor U1883 (N_1883,N_287,In_160);
and U1884 (N_1884,N_614,N_111);
nor U1885 (N_1885,In_1420,In_155);
xor U1886 (N_1886,N_72,N_905);
or U1887 (N_1887,N_51,In_1868);
xnor U1888 (N_1888,In_1465,In_1118);
xnor U1889 (N_1889,N_26,N_751);
and U1890 (N_1890,N_88,In_1858);
nand U1891 (N_1891,N_558,N_823);
xor U1892 (N_1892,In_1692,N_309);
and U1893 (N_1893,N_744,N_167);
nand U1894 (N_1894,N_770,In_2293);
xor U1895 (N_1895,N_425,N_741);
and U1896 (N_1896,N_840,N_197);
and U1897 (N_1897,In_235,N_6);
nand U1898 (N_1898,In_129,N_370);
xnor U1899 (N_1899,N_438,N_651);
nand U1900 (N_1900,N_804,N_858);
nor U1901 (N_1901,N_650,N_926);
nand U1902 (N_1902,N_353,N_751);
and U1903 (N_1903,N_5,In_352);
nor U1904 (N_1904,N_424,In_324);
or U1905 (N_1905,N_179,In_1250);
or U1906 (N_1906,N_86,In_751);
xor U1907 (N_1907,N_428,N_111);
xnor U1908 (N_1908,N_30,N_288);
and U1909 (N_1909,In_171,N_927);
nor U1910 (N_1910,N_125,N_924);
and U1911 (N_1911,N_510,N_464);
nor U1912 (N_1912,N_425,In_172);
or U1913 (N_1913,N_568,In_2283);
or U1914 (N_1914,In_1826,N_746);
nor U1915 (N_1915,N_522,N_394);
xnor U1916 (N_1916,N_93,In_1575);
xnor U1917 (N_1917,In_1785,N_63);
nor U1918 (N_1918,N_533,In_1385);
nor U1919 (N_1919,N_493,In_2379);
nor U1920 (N_1920,N_854,In_363);
xor U1921 (N_1921,In_2057,N_907);
or U1922 (N_1922,N_932,In_858);
and U1923 (N_1923,N_581,N_365);
nor U1924 (N_1924,In_2089,N_460);
xor U1925 (N_1925,N_719,N_30);
and U1926 (N_1926,N_990,In_2003);
and U1927 (N_1927,In_1465,N_125);
and U1928 (N_1928,N_217,In_1985);
or U1929 (N_1929,In_2490,In_2003);
nand U1930 (N_1930,N_164,N_159);
xnor U1931 (N_1931,N_453,N_76);
nand U1932 (N_1932,N_558,N_98);
or U1933 (N_1933,In_506,N_748);
nand U1934 (N_1934,N_336,N_486);
nor U1935 (N_1935,In_2308,N_509);
nor U1936 (N_1936,N_107,N_643);
or U1937 (N_1937,N_234,N_924);
nor U1938 (N_1938,N_225,N_164);
nor U1939 (N_1939,N_207,N_283);
and U1940 (N_1940,N_155,In_1595);
and U1941 (N_1941,N_639,N_930);
nor U1942 (N_1942,N_443,In_1114);
nand U1943 (N_1943,N_619,N_499);
or U1944 (N_1944,N_211,N_771);
nand U1945 (N_1945,N_199,N_450);
or U1946 (N_1946,N_677,N_817);
xor U1947 (N_1947,N_646,N_868);
and U1948 (N_1948,N_933,N_336);
xor U1949 (N_1949,N_77,N_445);
or U1950 (N_1950,N_871,N_81);
and U1951 (N_1951,N_169,In_2250);
nand U1952 (N_1952,N_203,N_143);
nand U1953 (N_1953,N_431,N_451);
xnor U1954 (N_1954,N_163,N_381);
or U1955 (N_1955,In_1193,N_565);
and U1956 (N_1956,In_503,In_1891);
nand U1957 (N_1957,N_499,N_236);
nor U1958 (N_1958,N_566,In_1388);
and U1959 (N_1959,N_456,N_744);
xnor U1960 (N_1960,N_30,N_967);
and U1961 (N_1961,N_522,N_177);
nor U1962 (N_1962,N_231,N_952);
or U1963 (N_1963,In_1741,N_847);
or U1964 (N_1964,N_471,N_518);
and U1965 (N_1965,N_894,In_1346);
nand U1966 (N_1966,In_1519,N_538);
nand U1967 (N_1967,In_1529,N_54);
or U1968 (N_1968,N_699,N_682);
xnor U1969 (N_1969,In_2187,N_441);
and U1970 (N_1970,N_942,N_216);
nand U1971 (N_1971,N_581,N_810);
nor U1972 (N_1972,N_790,N_733);
nand U1973 (N_1973,In_386,N_410);
nand U1974 (N_1974,N_543,In_645);
nor U1975 (N_1975,N_250,N_462);
and U1976 (N_1976,In_2456,N_695);
nor U1977 (N_1977,In_1202,N_801);
nor U1978 (N_1978,N_865,In_205);
and U1979 (N_1979,N_773,N_373);
and U1980 (N_1980,N_989,N_369);
and U1981 (N_1981,In_2060,N_277);
and U1982 (N_1982,N_836,N_113);
xor U1983 (N_1983,N_912,In_1606);
or U1984 (N_1984,In_479,N_362);
nor U1985 (N_1985,N_52,N_564);
or U1986 (N_1986,N_684,In_1387);
or U1987 (N_1987,N_644,N_856);
or U1988 (N_1988,In_324,N_633);
nand U1989 (N_1989,In_11,N_535);
xor U1990 (N_1990,N_600,N_661);
xor U1991 (N_1991,N_925,In_2336);
or U1992 (N_1992,In_1942,N_854);
nor U1993 (N_1993,N_47,In_1495);
or U1994 (N_1994,N_378,N_344);
xnor U1995 (N_1995,N_959,N_659);
and U1996 (N_1996,In_2220,N_328);
or U1997 (N_1997,N_693,N_888);
nor U1998 (N_1998,N_194,N_715);
and U1999 (N_1999,N_678,In_78);
nor U2000 (N_2000,N_1605,N_1873);
nand U2001 (N_2001,N_1661,N_1849);
or U2002 (N_2002,N_1125,N_1317);
and U2003 (N_2003,N_1530,N_1232);
nor U2004 (N_2004,N_1826,N_1914);
and U2005 (N_2005,N_1556,N_1336);
nor U2006 (N_2006,N_1299,N_1512);
or U2007 (N_2007,N_1811,N_1398);
and U2008 (N_2008,N_1380,N_1963);
nor U2009 (N_2009,N_1338,N_1272);
xor U2010 (N_2010,N_1074,N_1379);
or U2011 (N_2011,N_1886,N_1197);
or U2012 (N_2012,N_1840,N_1947);
or U2013 (N_2013,N_1083,N_1872);
nand U2014 (N_2014,N_1147,N_1846);
nand U2015 (N_2015,N_1607,N_1258);
nor U2016 (N_2016,N_1986,N_1511);
xnor U2017 (N_2017,N_1097,N_1725);
nand U2018 (N_2018,N_1807,N_1500);
and U2019 (N_2019,N_1797,N_1977);
nor U2020 (N_2020,N_1114,N_1227);
xnor U2021 (N_2021,N_1220,N_1773);
xnor U2022 (N_2022,N_1555,N_1766);
nand U2023 (N_2023,N_1681,N_1976);
nand U2024 (N_2024,N_1340,N_1505);
xnor U2025 (N_2025,N_1149,N_1396);
and U2026 (N_2026,N_1589,N_1824);
nor U2027 (N_2027,N_1858,N_1417);
nand U2028 (N_2028,N_1252,N_1208);
nand U2029 (N_2029,N_1603,N_1322);
and U2030 (N_2030,N_1009,N_1039);
xnor U2031 (N_2031,N_1950,N_1787);
or U2032 (N_2032,N_1597,N_1847);
and U2033 (N_2033,N_1779,N_1093);
xnor U2034 (N_2034,N_1163,N_1583);
or U2035 (N_2035,N_1890,N_1488);
nor U2036 (N_2036,N_1325,N_1566);
nand U2037 (N_2037,N_1819,N_1170);
nor U2038 (N_2038,N_1017,N_1407);
nor U2039 (N_2039,N_1011,N_1789);
or U2040 (N_2040,N_1301,N_1526);
and U2041 (N_2041,N_1572,N_1882);
and U2042 (N_2042,N_1187,N_1217);
nor U2043 (N_2043,N_1409,N_1831);
nand U2044 (N_2044,N_1007,N_1911);
or U2045 (N_2045,N_1860,N_1285);
and U2046 (N_2046,N_1867,N_1053);
and U2047 (N_2047,N_1710,N_1642);
xor U2048 (N_2048,N_1761,N_1075);
nand U2049 (N_2049,N_1198,N_1629);
nand U2050 (N_2050,N_1263,N_1884);
nor U2051 (N_2051,N_1416,N_1357);
or U2052 (N_2052,N_1988,N_1716);
xor U2053 (N_2053,N_1777,N_1763);
nor U2054 (N_2054,N_1062,N_1386);
nor U2055 (N_2055,N_1885,N_1660);
xor U2056 (N_2056,N_1800,N_1699);
xnor U2057 (N_2057,N_1016,N_1702);
or U2058 (N_2058,N_1203,N_1748);
and U2059 (N_2059,N_1120,N_1746);
xor U2060 (N_2060,N_1235,N_1997);
xnor U2061 (N_2061,N_1579,N_1656);
or U2062 (N_2062,N_1842,N_1767);
nand U2063 (N_2063,N_1598,N_1610);
or U2064 (N_2064,N_1506,N_1443);
and U2065 (N_2065,N_1538,N_1291);
and U2066 (N_2066,N_1672,N_1522);
xor U2067 (N_2067,N_1625,N_1048);
nand U2068 (N_2068,N_1080,N_1337);
and U2069 (N_2069,N_1814,N_1641);
nand U2070 (N_2070,N_1446,N_1085);
and U2071 (N_2071,N_1450,N_1617);
xor U2072 (N_2072,N_1843,N_1821);
xor U2073 (N_2073,N_1645,N_1167);
nand U2074 (N_2074,N_1164,N_1602);
nand U2075 (N_2075,N_1079,N_1411);
or U2076 (N_2076,N_1957,N_1816);
and U2077 (N_2077,N_1045,N_1102);
nand U2078 (N_2078,N_1376,N_1065);
nand U2079 (N_2079,N_1743,N_1833);
or U2080 (N_2080,N_1345,N_1528);
or U2081 (N_2081,N_1231,N_1736);
nor U2082 (N_2082,N_1124,N_1923);
xnor U2083 (N_2083,N_1503,N_1095);
or U2084 (N_2084,N_1837,N_1901);
nand U2085 (N_2085,N_1347,N_1920);
or U2086 (N_2086,N_1822,N_1434);
and U2087 (N_2087,N_1861,N_1611);
xor U2088 (N_2088,N_1334,N_1892);
xor U2089 (N_2089,N_1036,N_1713);
xnor U2090 (N_2090,N_1993,N_1276);
and U2091 (N_2091,N_1941,N_1119);
nor U2092 (N_2092,N_1883,N_1615);
xnor U2093 (N_2093,N_1937,N_1378);
nor U2094 (N_2094,N_1862,N_1518);
or U2095 (N_2095,N_1099,N_1513);
xnor U2096 (N_2096,N_1254,N_1212);
or U2097 (N_2097,N_1899,N_1444);
nand U2098 (N_2098,N_1658,N_1593);
nand U2099 (N_2099,N_1365,N_1367);
or U2100 (N_2100,N_1435,N_1620);
xor U2101 (N_2101,N_1823,N_1523);
nor U2102 (N_2102,N_1745,N_1280);
and U2103 (N_2103,N_1832,N_1253);
nand U2104 (N_2104,N_1240,N_1478);
or U2105 (N_2105,N_1935,N_1028);
xnor U2106 (N_2106,N_1349,N_1026);
xnor U2107 (N_2107,N_1490,N_1090);
nor U2108 (N_2108,N_1344,N_1876);
nor U2109 (N_2109,N_1155,N_1838);
and U2110 (N_2110,N_1968,N_1711);
xor U2111 (N_2111,N_1295,N_1096);
xnor U2112 (N_2112,N_1704,N_1659);
or U2113 (N_2113,N_1580,N_1408);
nand U2114 (N_2114,N_1183,N_1180);
nor U2115 (N_2115,N_1916,N_1738);
nand U2116 (N_2116,N_1390,N_1029);
nand U2117 (N_2117,N_1961,N_1161);
xnor U2118 (N_2118,N_1296,N_1186);
or U2119 (N_2119,N_1709,N_1448);
or U2120 (N_2120,N_1564,N_1588);
and U2121 (N_2121,N_1975,N_1030);
or U2122 (N_2122,N_1762,N_1479);
nor U2123 (N_2123,N_1524,N_1631);
or U2124 (N_2124,N_1493,N_1405);
or U2125 (N_2125,N_1126,N_1654);
and U2126 (N_2126,N_1496,N_1091);
xor U2127 (N_2127,N_1428,N_1744);
and U2128 (N_2128,N_1626,N_1735);
and U2129 (N_2129,N_1715,N_1550);
nor U2130 (N_2130,N_1893,N_1462);
nand U2131 (N_2131,N_1967,N_1801);
and U2132 (N_2132,N_1204,N_1297);
nor U2133 (N_2133,N_1201,N_1933);
nor U2134 (N_2134,N_1783,N_1023);
xor U2135 (N_2135,N_1207,N_1491);
or U2136 (N_2136,N_1078,N_1918);
nand U2137 (N_2137,N_1510,N_1841);
xor U2138 (N_2138,N_1592,N_1012);
xnor U2139 (N_2139,N_1540,N_1054);
xnor U2140 (N_2140,N_1969,N_1980);
and U2141 (N_2141,N_1752,N_1129);
nand U2142 (N_2142,N_1640,N_1088);
xnor U2143 (N_2143,N_1205,N_1393);
or U2144 (N_2144,N_1427,N_1382);
and U2145 (N_2145,N_1343,N_1655);
nand U2146 (N_2146,N_1723,N_1110);
xor U2147 (N_2147,N_1118,N_1989);
xnor U2148 (N_2148,N_1353,N_1994);
nor U2149 (N_2149,N_1117,N_1774);
or U2150 (N_2150,N_1902,N_1300);
nand U2151 (N_2151,N_1581,N_1547);
and U2152 (N_2152,N_1303,N_1150);
nand U2153 (N_2153,N_1314,N_1680);
or U2154 (N_2154,N_1638,N_1703);
nand U2155 (N_2155,N_1192,N_1596);
nand U2156 (N_2156,N_1894,N_1852);
nor U2157 (N_2157,N_1333,N_1475);
nor U2158 (N_2158,N_1246,N_1888);
nor U2159 (N_2159,N_1070,N_1829);
xor U2160 (N_2160,N_1895,N_1237);
and U2161 (N_2161,N_1728,N_1373);
xor U2162 (N_2162,N_1650,N_1594);
and U2163 (N_2163,N_1678,N_1109);
nor U2164 (N_2164,N_1696,N_1928);
xnor U2165 (N_2165,N_1193,N_1669);
xnor U2166 (N_2166,N_1487,N_1747);
nor U2167 (N_2167,N_1328,N_1987);
nor U2168 (N_2168,N_1828,N_1371);
nand U2169 (N_2169,N_1940,N_1845);
nand U2170 (N_2170,N_1750,N_1853);
nand U2171 (N_2171,N_1850,N_1754);
nand U2172 (N_2172,N_1174,N_1018);
and U2173 (N_2173,N_1414,N_1855);
or U2174 (N_2174,N_1794,N_1071);
and U2175 (N_2175,N_1684,N_1529);
xor U2176 (N_2176,N_1536,N_1308);
or U2177 (N_2177,N_1481,N_1908);
and U2178 (N_2178,N_1905,N_1804);
and U2179 (N_2179,N_1068,N_1226);
or U2180 (N_2180,N_1241,N_1058);
or U2181 (N_2181,N_1974,N_1881);
nor U2182 (N_2182,N_1310,N_1544);
nand U2183 (N_2183,N_1486,N_1552);
xnor U2184 (N_2184,N_1820,N_1509);
nand U2185 (N_2185,N_1447,N_1135);
or U2186 (N_2186,N_1910,N_1004);
and U2187 (N_2187,N_1959,N_1982);
xnor U2188 (N_2188,N_1692,N_1717);
nor U2189 (N_2189,N_1546,N_1087);
or U2190 (N_2190,N_1664,N_1483);
xnor U2191 (N_2191,N_1685,N_1250);
nor U2192 (N_2192,N_1104,N_1489);
nand U2193 (N_2193,N_1608,N_1422);
nand U2194 (N_2194,N_1366,N_1647);
nand U2195 (N_2195,N_1247,N_1595);
nor U2196 (N_2196,N_1306,N_1055);
nand U2197 (N_2197,N_1027,N_1288);
nand U2198 (N_2198,N_1775,N_1707);
xor U2199 (N_2199,N_1425,N_1484);
nand U2200 (N_2200,N_1168,N_1778);
and U2201 (N_2201,N_1000,N_1979);
nand U2202 (N_2202,N_1760,N_1674);
nor U2203 (N_2203,N_1047,N_1307);
and U2204 (N_2204,N_1809,N_1267);
nand U2205 (N_2205,N_1113,N_1724);
and U2206 (N_2206,N_1219,N_1929);
nor U2207 (N_2207,N_1255,N_1942);
nand U2208 (N_2208,N_1499,N_1041);
nand U2209 (N_2209,N_1172,N_1144);
or U2210 (N_2210,N_1477,N_1182);
xnor U2211 (N_2211,N_1952,N_1156);
and U2212 (N_2212,N_1412,N_1158);
or U2213 (N_2213,N_1131,N_1545);
xnor U2214 (N_2214,N_1903,N_1992);
nor U2215 (N_2215,N_1604,N_1930);
nand U2216 (N_2216,N_1962,N_1561);
or U2217 (N_2217,N_1244,N_1388);
and U2218 (N_2218,N_1067,N_1813);
or U2219 (N_2219,N_1209,N_1279);
nor U2220 (N_2220,N_1558,N_1983);
xnor U2221 (N_2221,N_1534,N_1358);
and U2222 (N_2222,N_1966,N_1264);
or U2223 (N_2223,N_1757,N_1931);
xor U2224 (N_2224,N_1420,N_1958);
nand U2225 (N_2225,N_1234,N_1739);
nand U2226 (N_2226,N_1426,N_1472);
xnor U2227 (N_2227,N_1939,N_1318);
nand U2228 (N_2228,N_1374,N_1363);
or U2229 (N_2229,N_1248,N_1557);
nor U2230 (N_2230,N_1415,N_1582);
and U2231 (N_2231,N_1854,N_1081);
and U2232 (N_2232,N_1651,N_1421);
and U2233 (N_2233,N_1865,N_1917);
or U2234 (N_2234,N_1494,N_1224);
and U2235 (N_2235,N_1525,N_1145);
and U2236 (N_2236,N_1900,N_1233);
xnor U2237 (N_2237,N_1229,N_1548);
nand U2238 (N_2238,N_1277,N_1706);
nand U2239 (N_2239,N_1348,N_1470);
xnor U2240 (N_2240,N_1984,N_1077);
or U2241 (N_2241,N_1430,N_1037);
and U2242 (N_2242,N_1159,N_1630);
nor U2243 (N_2243,N_1671,N_1830);
or U2244 (N_2244,N_1137,N_1298);
nand U2245 (N_2245,N_1906,N_1501);
nor U2246 (N_2246,N_1038,N_1619);
and U2247 (N_2247,N_1498,N_1316);
nor U2248 (N_2248,N_1364,N_1516);
or U2249 (N_2249,N_1342,N_1627);
and U2250 (N_2250,N_1200,N_1022);
xor U2251 (N_2251,N_1014,N_1476);
nand U2252 (N_2252,N_1520,N_1397);
and U2253 (N_2253,N_1568,N_1211);
nor U2254 (N_2254,N_1370,N_1278);
or U2255 (N_2255,N_1010,N_1798);
nor U2256 (N_2256,N_1266,N_1624);
nor U2257 (N_2257,N_1897,N_1944);
xor U2258 (N_2258,N_1817,N_1866);
nor U2259 (N_2259,N_1578,N_1889);
or U2260 (N_2260,N_1485,N_1864);
and U2261 (N_2261,N_1756,N_1575);
nand U2262 (N_2262,N_1835,N_1793);
nor U2263 (N_2263,N_1271,N_1469);
nor U2264 (N_2264,N_1262,N_1105);
nand U2265 (N_2265,N_1072,N_1352);
nand U2266 (N_2266,N_1265,N_1812);
nand U2267 (N_2267,N_1221,N_1999);
nand U2268 (N_2268,N_1537,N_1721);
or U2269 (N_2269,N_1152,N_1463);
nor U2270 (N_2270,N_1515,N_1805);
xnor U2271 (N_2271,N_1210,N_1391);
and U2272 (N_2272,N_1153,N_1392);
nor U2273 (N_2273,N_1178,N_1532);
xor U2274 (N_2274,N_1216,N_1290);
or U2275 (N_2275,N_1273,N_1176);
xnor U2276 (N_2276,N_1031,N_1926);
xnor U2277 (N_2277,N_1061,N_1875);
xnor U2278 (N_2278,N_1912,N_1433);
xnor U2279 (N_2279,N_1549,N_1006);
and U2280 (N_2280,N_1418,N_1973);
and U2281 (N_2281,N_1024,N_1245);
nand U2282 (N_2282,N_1141,N_1878);
or U2283 (N_2283,N_1718,N_1332);
xnor U2284 (N_2284,N_1693,N_1945);
or U2285 (N_2285,N_1107,N_1868);
nand U2286 (N_2286,N_1368,N_1051);
or U2287 (N_2287,N_1329,N_1199);
nor U2288 (N_2288,N_1586,N_1639);
nor U2289 (N_2289,N_1101,N_1169);
and U2290 (N_2290,N_1181,N_1175);
nand U2291 (N_2291,N_1554,N_1825);
xnor U2292 (N_2292,N_1034,N_1160);
xor U2293 (N_2293,N_1726,N_1733);
nand U2294 (N_2294,N_1740,N_1327);
nor U2295 (N_2295,N_1372,N_1331);
or U2296 (N_2296,N_1653,N_1003);
and U2297 (N_2297,N_1857,N_1880);
xnor U2298 (N_2298,N_1218,N_1727);
or U2299 (N_2299,N_1440,N_1050);
and U2300 (N_2300,N_1060,N_1064);
nand U2301 (N_2301,N_1441,N_1351);
xor U2302 (N_2302,N_1719,N_1682);
nand U2303 (N_2303,N_1714,N_1431);
or U2304 (N_2304,N_1970,N_1686);
and U2305 (N_2305,N_1749,N_1946);
and U2306 (N_2306,N_1304,N_1230);
or U2307 (N_2307,N_1891,N_1321);
or U2308 (N_2308,N_1335,N_1098);
or U2309 (N_2309,N_1646,N_1613);
and U2310 (N_2310,N_1844,N_1243);
nand U2311 (N_2311,N_1913,N_1657);
xnor U2312 (N_2312,N_1213,N_1785);
and U2313 (N_2313,N_1690,N_1020);
xor U2314 (N_2314,N_1151,N_1189);
or U2315 (N_2315,N_1251,N_1951);
and U2316 (N_2316,N_1543,N_1453);
nand U2317 (N_2317,N_1413,N_1765);
nand U2318 (N_2318,N_1565,N_1996);
nand U2319 (N_2319,N_1195,N_1236);
nor U2320 (N_2320,N_1179,N_1471);
nor U2321 (N_2321,N_1387,N_1551);
nand U2322 (N_2322,N_1571,N_1587);
nor U2323 (N_2323,N_1196,N_1438);
nor U2324 (N_2324,N_1577,N_1116);
and U2325 (N_2325,N_1429,N_1184);
or U2326 (N_2326,N_1312,N_1395);
and U2327 (N_2327,N_1720,N_1035);
and U2328 (N_2328,N_1652,N_1755);
xor U2329 (N_2329,N_1292,N_1375);
and U2330 (N_2330,N_1356,N_1998);
nand U2331 (N_2331,N_1519,N_1776);
or U2332 (N_2332,N_1863,N_1270);
nand U2333 (N_2333,N_1874,N_1008);
nand U2334 (N_2334,N_1410,N_1040);
or U2335 (N_2335,N_1698,N_1274);
or U2336 (N_2336,N_1089,N_1621);
nor U2337 (N_2337,N_1046,N_1015);
or U2338 (N_2338,N_1361,N_1005);
xor U2339 (N_2339,N_1456,N_1025);
nor U2340 (N_2340,N_1609,N_1792);
and U2341 (N_2341,N_1535,N_1474);
or U2342 (N_2342,N_1677,N_1103);
xor U2343 (N_2343,N_1032,N_1570);
xor U2344 (N_2344,N_1482,N_1442);
xor U2345 (N_2345,N_1339,N_1389);
nor U2346 (N_2346,N_1687,N_1130);
nand U2347 (N_2347,N_1585,N_1092);
nor U2348 (N_2348,N_1780,N_1601);
nor U2349 (N_2349,N_1286,N_1402);
xor U2350 (N_2350,N_1695,N_1445);
or U2351 (N_2351,N_1722,N_1697);
or U2352 (N_2352,N_1851,N_1249);
and U2353 (N_2353,N_1694,N_1454);
xnor U2354 (N_2354,N_1668,N_1013);
nand U2355 (N_2355,N_1121,N_1206);
nand U2356 (N_2356,N_1282,N_1399);
or U2357 (N_2357,N_1810,N_1790);
and U2358 (N_2358,N_1134,N_1173);
xnor U2359 (N_2359,N_1730,N_1675);
xor U2360 (N_2360,N_1260,N_1188);
or U2361 (N_2361,N_1781,N_1734);
xor U2362 (N_2362,N_1289,N_1533);
or U2363 (N_2363,N_1139,N_1964);
nand U2364 (N_2364,N_1791,N_1100);
nand U2365 (N_2365,N_1934,N_1667);
xnor U2366 (N_2366,N_1112,N_1369);
nor U2367 (N_2367,N_1887,N_1502);
nand U2368 (N_2368,N_1225,N_1590);
nand U2369 (N_2369,N_1185,N_1758);
nor U2370 (N_2370,N_1021,N_1737);
or U2371 (N_2371,N_1539,N_1381);
nor U2372 (N_2372,N_1936,N_1133);
and U2373 (N_2373,N_1788,N_1531);
nand U2374 (N_2374,N_1978,N_1729);
xor U2375 (N_2375,N_1806,N_1818);
nor U2376 (N_2376,N_1452,N_1559);
or U2377 (N_2377,N_1504,N_1799);
or U2378 (N_2378,N_1953,N_1042);
nor U2379 (N_2379,N_1157,N_1636);
xnor U2380 (N_2380,N_1848,N_1676);
nor U2381 (N_2381,N_1148,N_1839);
nor U2382 (N_2382,N_1691,N_1569);
or U2383 (N_2383,N_1394,N_1637);
nor U2384 (N_2384,N_1769,N_1073);
or U2385 (N_2385,N_1633,N_1877);
nand U2386 (N_2386,N_1359,N_1403);
xor U2387 (N_2387,N_1606,N_1741);
nor U2388 (N_2388,N_1283,N_1305);
or U2389 (N_2389,N_1424,N_1981);
and U2390 (N_2390,N_1122,N_1492);
or U2391 (N_2391,N_1127,N_1662);
nor U2392 (N_2392,N_1326,N_1069);
or U2393 (N_2393,N_1377,N_1449);
nand U2394 (N_2394,N_1753,N_1782);
nor U2395 (N_2395,N_1464,N_1287);
or U2396 (N_2396,N_1460,N_1495);
xnor U2397 (N_2397,N_1938,N_1896);
xnor U2398 (N_2398,N_1965,N_1665);
and U2399 (N_2399,N_1808,N_1261);
xor U2400 (N_2400,N_1439,N_1856);
or U2401 (N_2401,N_1106,N_1670);
nor U2402 (N_2402,N_1320,N_1632);
or U2403 (N_2403,N_1907,N_1527);
nor U2404 (N_2404,N_1898,N_1406);
xnor U2405 (N_2405,N_1731,N_1111);
xnor U2406 (N_2406,N_1057,N_1082);
or U2407 (N_2407,N_1772,N_1228);
or U2408 (N_2408,N_1870,N_1436);
nor U2409 (N_2409,N_1330,N_1385);
and U2410 (N_2410,N_1400,N_1927);
nor U2411 (N_2411,N_1796,N_1949);
or U2412 (N_2412,N_1214,N_1066);
nand U2413 (N_2413,N_1960,N_1284);
xor U2414 (N_2414,N_1458,N_1242);
and U2415 (N_2415,N_1128,N_1033);
xor U2416 (N_2416,N_1309,N_1784);
xor U2417 (N_2417,N_1751,N_1688);
or U2418 (N_2418,N_1084,N_1269);
xor U2419 (N_2419,N_1795,N_1076);
or U2420 (N_2420,N_1628,N_1256);
nand U2421 (N_2421,N_1311,N_1323);
or U2422 (N_2422,N_1764,N_1956);
nand U2423 (N_2423,N_1507,N_1275);
or U2424 (N_2424,N_1635,N_1985);
xor U2425 (N_2425,N_1455,N_1834);
nor U2426 (N_2426,N_1701,N_1384);
or U2427 (N_2427,N_1614,N_1770);
and U2428 (N_2428,N_1514,N_1467);
or U2429 (N_2429,N_1542,N_1324);
or U2430 (N_2430,N_1268,N_1712);
xor U2431 (N_2431,N_1612,N_1354);
nor U2432 (N_2432,N_1990,N_1742);
nor U2433 (N_2433,N_1803,N_1932);
or U2434 (N_2434,N_1052,N_1648);
or U2435 (N_2435,N_1281,N_1666);
and U2436 (N_2436,N_1644,N_1508);
and U2437 (N_2437,N_1223,N_1190);
nand U2438 (N_2438,N_1521,N_1705);
nand U2439 (N_2439,N_1465,N_1350);
or U2440 (N_2440,N_1643,N_1154);
xor U2441 (N_2441,N_1383,N_1759);
xnor U2442 (N_2442,N_1191,N_1497);
nand U2443 (N_2443,N_1708,N_1166);
and U2444 (N_2444,N_1215,N_1086);
or U2445 (N_2445,N_1001,N_1238);
nor U2446 (N_2446,N_1362,N_1859);
nor U2447 (N_2447,N_1584,N_1591);
nand U2448 (N_2448,N_1827,N_1553);
nand U2449 (N_2449,N_1401,N_1043);
nor U2450 (N_2450,N_1815,N_1562);
and U2451 (N_2451,N_1259,N_1871);
nor U2452 (N_2452,N_1404,N_1802);
or U2453 (N_2453,N_1315,N_1302);
or U2454 (N_2454,N_1056,N_1673);
nor U2455 (N_2455,N_1423,N_1732);
or U2456 (N_2456,N_1700,N_1239);
nand U2457 (N_2457,N_1517,N_1123);
xor U2458 (N_2458,N_1567,N_1616);
and U2459 (N_2459,N_1921,N_1634);
nand U2460 (N_2460,N_1257,N_1480);
nor U2461 (N_2461,N_1419,N_1915);
nor U2462 (N_2462,N_1768,N_1541);
nand U2463 (N_2463,N_1786,N_1771);
or U2464 (N_2464,N_1459,N_1649);
or U2465 (N_2465,N_1194,N_1955);
and U2466 (N_2466,N_1451,N_1222);
nor U2467 (N_2467,N_1143,N_1954);
xnor U2468 (N_2468,N_1360,N_1294);
nand U2469 (N_2469,N_1142,N_1943);
nor U2470 (N_2470,N_1171,N_1136);
and U2471 (N_2471,N_1576,N_1623);
or U2472 (N_2472,N_1044,N_1063);
nand U2473 (N_2473,N_1346,N_1108);
xor U2474 (N_2474,N_1457,N_1879);
xor U2475 (N_2475,N_1663,N_1341);
and U2476 (N_2476,N_1971,N_1293);
or U2477 (N_2477,N_1138,N_1991);
or U2478 (N_2478,N_1995,N_1002);
nor U2479 (N_2479,N_1600,N_1473);
xor U2480 (N_2480,N_1869,N_1622);
nor U2481 (N_2481,N_1165,N_1162);
and U2482 (N_2482,N_1049,N_1468);
and U2483 (N_2483,N_1599,N_1461);
and U2484 (N_2484,N_1972,N_1683);
nor U2485 (N_2485,N_1560,N_1948);
nor U2486 (N_2486,N_1319,N_1574);
and U2487 (N_2487,N_1924,N_1563);
nor U2488 (N_2488,N_1618,N_1059);
xor U2489 (N_2489,N_1679,N_1115);
xor U2490 (N_2490,N_1925,N_1909);
xnor U2491 (N_2491,N_1466,N_1132);
or U2492 (N_2492,N_1355,N_1922);
and U2493 (N_2493,N_1177,N_1836);
nand U2494 (N_2494,N_1146,N_1904);
or U2495 (N_2495,N_1437,N_1432);
and U2496 (N_2496,N_1919,N_1689);
xnor U2497 (N_2497,N_1140,N_1573);
nor U2498 (N_2498,N_1313,N_1202);
and U2499 (N_2499,N_1019,N_1094);
xor U2500 (N_2500,N_1318,N_1867);
nor U2501 (N_2501,N_1034,N_1009);
nor U2502 (N_2502,N_1492,N_1547);
xor U2503 (N_2503,N_1801,N_1110);
nor U2504 (N_2504,N_1377,N_1094);
nor U2505 (N_2505,N_1394,N_1910);
or U2506 (N_2506,N_1680,N_1641);
xnor U2507 (N_2507,N_1406,N_1226);
nor U2508 (N_2508,N_1433,N_1731);
nor U2509 (N_2509,N_1044,N_1118);
and U2510 (N_2510,N_1568,N_1561);
nor U2511 (N_2511,N_1062,N_1393);
or U2512 (N_2512,N_1108,N_1408);
xnor U2513 (N_2513,N_1183,N_1330);
nand U2514 (N_2514,N_1026,N_1533);
nand U2515 (N_2515,N_1909,N_1835);
nor U2516 (N_2516,N_1592,N_1947);
xnor U2517 (N_2517,N_1064,N_1509);
nor U2518 (N_2518,N_1069,N_1844);
nor U2519 (N_2519,N_1497,N_1918);
or U2520 (N_2520,N_1077,N_1157);
nand U2521 (N_2521,N_1547,N_1087);
xnor U2522 (N_2522,N_1541,N_1152);
or U2523 (N_2523,N_1090,N_1657);
nor U2524 (N_2524,N_1332,N_1605);
or U2525 (N_2525,N_1939,N_1773);
nor U2526 (N_2526,N_1911,N_1358);
xnor U2527 (N_2527,N_1881,N_1644);
nor U2528 (N_2528,N_1138,N_1598);
nor U2529 (N_2529,N_1817,N_1380);
or U2530 (N_2530,N_1770,N_1854);
nor U2531 (N_2531,N_1258,N_1208);
nor U2532 (N_2532,N_1079,N_1856);
xor U2533 (N_2533,N_1948,N_1138);
or U2534 (N_2534,N_1406,N_1077);
nor U2535 (N_2535,N_1407,N_1059);
nand U2536 (N_2536,N_1191,N_1553);
xor U2537 (N_2537,N_1222,N_1720);
or U2538 (N_2538,N_1227,N_1766);
nor U2539 (N_2539,N_1998,N_1116);
nand U2540 (N_2540,N_1812,N_1218);
xor U2541 (N_2541,N_1503,N_1472);
xor U2542 (N_2542,N_1399,N_1431);
nand U2543 (N_2543,N_1866,N_1118);
xnor U2544 (N_2544,N_1062,N_1225);
and U2545 (N_2545,N_1994,N_1896);
xnor U2546 (N_2546,N_1547,N_1089);
or U2547 (N_2547,N_1338,N_1312);
and U2548 (N_2548,N_1875,N_1111);
nand U2549 (N_2549,N_1878,N_1199);
xnor U2550 (N_2550,N_1232,N_1660);
nor U2551 (N_2551,N_1151,N_1027);
and U2552 (N_2552,N_1622,N_1744);
nand U2553 (N_2553,N_1960,N_1228);
or U2554 (N_2554,N_1800,N_1851);
nand U2555 (N_2555,N_1649,N_1564);
nand U2556 (N_2556,N_1488,N_1904);
nor U2557 (N_2557,N_1322,N_1938);
nand U2558 (N_2558,N_1296,N_1438);
nand U2559 (N_2559,N_1542,N_1742);
nand U2560 (N_2560,N_1076,N_1431);
xor U2561 (N_2561,N_1778,N_1415);
and U2562 (N_2562,N_1372,N_1054);
nand U2563 (N_2563,N_1913,N_1069);
and U2564 (N_2564,N_1551,N_1191);
xnor U2565 (N_2565,N_1605,N_1409);
or U2566 (N_2566,N_1789,N_1756);
nand U2567 (N_2567,N_1841,N_1044);
nand U2568 (N_2568,N_1481,N_1343);
nor U2569 (N_2569,N_1301,N_1944);
nand U2570 (N_2570,N_1086,N_1062);
nor U2571 (N_2571,N_1262,N_1754);
or U2572 (N_2572,N_1978,N_1752);
xor U2573 (N_2573,N_1966,N_1757);
and U2574 (N_2574,N_1680,N_1905);
or U2575 (N_2575,N_1474,N_1339);
xor U2576 (N_2576,N_1696,N_1608);
nor U2577 (N_2577,N_1737,N_1044);
xnor U2578 (N_2578,N_1193,N_1247);
and U2579 (N_2579,N_1600,N_1679);
or U2580 (N_2580,N_1752,N_1321);
nand U2581 (N_2581,N_1063,N_1452);
nand U2582 (N_2582,N_1750,N_1532);
nand U2583 (N_2583,N_1771,N_1873);
nor U2584 (N_2584,N_1576,N_1654);
or U2585 (N_2585,N_1352,N_1989);
and U2586 (N_2586,N_1725,N_1899);
nand U2587 (N_2587,N_1160,N_1682);
xor U2588 (N_2588,N_1140,N_1606);
nand U2589 (N_2589,N_1161,N_1515);
xnor U2590 (N_2590,N_1325,N_1352);
xnor U2591 (N_2591,N_1295,N_1146);
nand U2592 (N_2592,N_1586,N_1304);
or U2593 (N_2593,N_1759,N_1270);
or U2594 (N_2594,N_1083,N_1761);
or U2595 (N_2595,N_1570,N_1894);
or U2596 (N_2596,N_1366,N_1250);
and U2597 (N_2597,N_1961,N_1351);
xor U2598 (N_2598,N_1857,N_1004);
xor U2599 (N_2599,N_1856,N_1537);
xnor U2600 (N_2600,N_1330,N_1805);
and U2601 (N_2601,N_1697,N_1378);
nor U2602 (N_2602,N_1949,N_1671);
and U2603 (N_2603,N_1866,N_1147);
xor U2604 (N_2604,N_1585,N_1964);
xnor U2605 (N_2605,N_1851,N_1854);
and U2606 (N_2606,N_1576,N_1337);
or U2607 (N_2607,N_1977,N_1478);
nand U2608 (N_2608,N_1369,N_1795);
and U2609 (N_2609,N_1216,N_1908);
nand U2610 (N_2610,N_1478,N_1072);
and U2611 (N_2611,N_1116,N_1439);
nor U2612 (N_2612,N_1624,N_1344);
and U2613 (N_2613,N_1238,N_1661);
nor U2614 (N_2614,N_1636,N_1205);
nor U2615 (N_2615,N_1376,N_1777);
and U2616 (N_2616,N_1568,N_1841);
or U2617 (N_2617,N_1645,N_1870);
nand U2618 (N_2618,N_1308,N_1385);
xor U2619 (N_2619,N_1714,N_1638);
or U2620 (N_2620,N_1956,N_1794);
xnor U2621 (N_2621,N_1555,N_1183);
xor U2622 (N_2622,N_1556,N_1656);
xor U2623 (N_2623,N_1737,N_1905);
and U2624 (N_2624,N_1295,N_1521);
and U2625 (N_2625,N_1621,N_1680);
nand U2626 (N_2626,N_1354,N_1174);
xnor U2627 (N_2627,N_1996,N_1306);
xnor U2628 (N_2628,N_1848,N_1731);
nand U2629 (N_2629,N_1615,N_1981);
nand U2630 (N_2630,N_1279,N_1941);
and U2631 (N_2631,N_1964,N_1940);
and U2632 (N_2632,N_1149,N_1428);
nor U2633 (N_2633,N_1531,N_1757);
nor U2634 (N_2634,N_1141,N_1762);
nor U2635 (N_2635,N_1741,N_1431);
xnor U2636 (N_2636,N_1756,N_1967);
or U2637 (N_2637,N_1343,N_1510);
nor U2638 (N_2638,N_1578,N_1911);
and U2639 (N_2639,N_1555,N_1323);
nand U2640 (N_2640,N_1889,N_1204);
xnor U2641 (N_2641,N_1568,N_1483);
or U2642 (N_2642,N_1024,N_1763);
xor U2643 (N_2643,N_1657,N_1081);
nand U2644 (N_2644,N_1069,N_1609);
nor U2645 (N_2645,N_1733,N_1267);
nand U2646 (N_2646,N_1208,N_1193);
or U2647 (N_2647,N_1730,N_1063);
nand U2648 (N_2648,N_1053,N_1494);
xnor U2649 (N_2649,N_1459,N_1897);
or U2650 (N_2650,N_1107,N_1747);
nor U2651 (N_2651,N_1503,N_1983);
xnor U2652 (N_2652,N_1426,N_1505);
and U2653 (N_2653,N_1836,N_1209);
xnor U2654 (N_2654,N_1385,N_1674);
xnor U2655 (N_2655,N_1656,N_1085);
nor U2656 (N_2656,N_1267,N_1643);
and U2657 (N_2657,N_1573,N_1612);
and U2658 (N_2658,N_1020,N_1720);
nor U2659 (N_2659,N_1530,N_1442);
and U2660 (N_2660,N_1162,N_1114);
xnor U2661 (N_2661,N_1841,N_1634);
and U2662 (N_2662,N_1086,N_1690);
and U2663 (N_2663,N_1924,N_1504);
or U2664 (N_2664,N_1674,N_1094);
and U2665 (N_2665,N_1252,N_1212);
or U2666 (N_2666,N_1802,N_1178);
nand U2667 (N_2667,N_1527,N_1520);
xnor U2668 (N_2668,N_1793,N_1948);
and U2669 (N_2669,N_1352,N_1832);
nand U2670 (N_2670,N_1616,N_1593);
or U2671 (N_2671,N_1738,N_1829);
xnor U2672 (N_2672,N_1111,N_1866);
nand U2673 (N_2673,N_1498,N_1734);
nand U2674 (N_2674,N_1997,N_1369);
xnor U2675 (N_2675,N_1636,N_1206);
and U2676 (N_2676,N_1827,N_1457);
xnor U2677 (N_2677,N_1572,N_1831);
xor U2678 (N_2678,N_1828,N_1816);
nor U2679 (N_2679,N_1577,N_1119);
nor U2680 (N_2680,N_1283,N_1982);
and U2681 (N_2681,N_1532,N_1438);
nor U2682 (N_2682,N_1719,N_1764);
or U2683 (N_2683,N_1914,N_1706);
and U2684 (N_2684,N_1395,N_1360);
xnor U2685 (N_2685,N_1384,N_1432);
and U2686 (N_2686,N_1614,N_1667);
or U2687 (N_2687,N_1559,N_1060);
xnor U2688 (N_2688,N_1928,N_1612);
nand U2689 (N_2689,N_1408,N_1372);
xor U2690 (N_2690,N_1406,N_1901);
and U2691 (N_2691,N_1543,N_1456);
and U2692 (N_2692,N_1298,N_1421);
nand U2693 (N_2693,N_1301,N_1996);
xor U2694 (N_2694,N_1721,N_1084);
nor U2695 (N_2695,N_1500,N_1369);
nand U2696 (N_2696,N_1283,N_1233);
and U2697 (N_2697,N_1661,N_1270);
nand U2698 (N_2698,N_1638,N_1168);
nor U2699 (N_2699,N_1913,N_1373);
nand U2700 (N_2700,N_1540,N_1844);
and U2701 (N_2701,N_1381,N_1296);
xor U2702 (N_2702,N_1061,N_1975);
xnor U2703 (N_2703,N_1487,N_1192);
or U2704 (N_2704,N_1298,N_1509);
nor U2705 (N_2705,N_1281,N_1398);
nand U2706 (N_2706,N_1967,N_1185);
or U2707 (N_2707,N_1258,N_1157);
nand U2708 (N_2708,N_1025,N_1203);
nand U2709 (N_2709,N_1283,N_1094);
or U2710 (N_2710,N_1990,N_1435);
or U2711 (N_2711,N_1753,N_1431);
xor U2712 (N_2712,N_1067,N_1983);
nor U2713 (N_2713,N_1757,N_1615);
and U2714 (N_2714,N_1323,N_1993);
xor U2715 (N_2715,N_1820,N_1692);
nand U2716 (N_2716,N_1223,N_1755);
or U2717 (N_2717,N_1688,N_1670);
and U2718 (N_2718,N_1294,N_1933);
and U2719 (N_2719,N_1201,N_1903);
or U2720 (N_2720,N_1622,N_1683);
and U2721 (N_2721,N_1760,N_1136);
and U2722 (N_2722,N_1053,N_1457);
nand U2723 (N_2723,N_1781,N_1844);
nor U2724 (N_2724,N_1605,N_1169);
or U2725 (N_2725,N_1748,N_1409);
or U2726 (N_2726,N_1951,N_1556);
xnor U2727 (N_2727,N_1983,N_1732);
xnor U2728 (N_2728,N_1797,N_1945);
nor U2729 (N_2729,N_1082,N_1419);
nand U2730 (N_2730,N_1843,N_1972);
nor U2731 (N_2731,N_1431,N_1239);
and U2732 (N_2732,N_1134,N_1822);
nand U2733 (N_2733,N_1926,N_1548);
or U2734 (N_2734,N_1853,N_1344);
nor U2735 (N_2735,N_1201,N_1754);
xnor U2736 (N_2736,N_1279,N_1037);
or U2737 (N_2737,N_1188,N_1080);
nor U2738 (N_2738,N_1890,N_1356);
or U2739 (N_2739,N_1191,N_1316);
nand U2740 (N_2740,N_1385,N_1592);
xnor U2741 (N_2741,N_1379,N_1016);
xnor U2742 (N_2742,N_1311,N_1805);
and U2743 (N_2743,N_1262,N_1220);
or U2744 (N_2744,N_1908,N_1857);
nand U2745 (N_2745,N_1357,N_1030);
and U2746 (N_2746,N_1635,N_1044);
xnor U2747 (N_2747,N_1721,N_1027);
or U2748 (N_2748,N_1236,N_1276);
nor U2749 (N_2749,N_1745,N_1587);
and U2750 (N_2750,N_1005,N_1128);
or U2751 (N_2751,N_1764,N_1720);
nand U2752 (N_2752,N_1974,N_1441);
xor U2753 (N_2753,N_1310,N_1280);
or U2754 (N_2754,N_1355,N_1105);
nand U2755 (N_2755,N_1287,N_1937);
and U2756 (N_2756,N_1523,N_1186);
and U2757 (N_2757,N_1282,N_1393);
nor U2758 (N_2758,N_1933,N_1760);
nand U2759 (N_2759,N_1057,N_1929);
xor U2760 (N_2760,N_1603,N_1960);
xor U2761 (N_2761,N_1178,N_1546);
nor U2762 (N_2762,N_1419,N_1367);
and U2763 (N_2763,N_1679,N_1364);
nor U2764 (N_2764,N_1682,N_1535);
xnor U2765 (N_2765,N_1986,N_1688);
nand U2766 (N_2766,N_1620,N_1085);
or U2767 (N_2767,N_1097,N_1956);
and U2768 (N_2768,N_1403,N_1300);
xor U2769 (N_2769,N_1155,N_1262);
nand U2770 (N_2770,N_1670,N_1685);
xnor U2771 (N_2771,N_1368,N_1035);
and U2772 (N_2772,N_1045,N_1765);
nor U2773 (N_2773,N_1467,N_1989);
or U2774 (N_2774,N_1886,N_1881);
or U2775 (N_2775,N_1337,N_1689);
and U2776 (N_2776,N_1909,N_1376);
xnor U2777 (N_2777,N_1880,N_1136);
xor U2778 (N_2778,N_1829,N_1037);
nand U2779 (N_2779,N_1274,N_1800);
nand U2780 (N_2780,N_1142,N_1150);
nor U2781 (N_2781,N_1479,N_1032);
nor U2782 (N_2782,N_1077,N_1490);
nand U2783 (N_2783,N_1252,N_1479);
xnor U2784 (N_2784,N_1015,N_1257);
nand U2785 (N_2785,N_1612,N_1683);
nand U2786 (N_2786,N_1389,N_1634);
nand U2787 (N_2787,N_1621,N_1341);
nor U2788 (N_2788,N_1043,N_1169);
or U2789 (N_2789,N_1267,N_1732);
and U2790 (N_2790,N_1520,N_1485);
and U2791 (N_2791,N_1041,N_1175);
nor U2792 (N_2792,N_1024,N_1977);
or U2793 (N_2793,N_1900,N_1068);
and U2794 (N_2794,N_1937,N_1100);
and U2795 (N_2795,N_1943,N_1873);
and U2796 (N_2796,N_1863,N_1446);
xnor U2797 (N_2797,N_1335,N_1730);
and U2798 (N_2798,N_1230,N_1474);
or U2799 (N_2799,N_1991,N_1378);
nor U2800 (N_2800,N_1761,N_1791);
nand U2801 (N_2801,N_1236,N_1377);
nor U2802 (N_2802,N_1197,N_1202);
xnor U2803 (N_2803,N_1559,N_1221);
nor U2804 (N_2804,N_1101,N_1105);
nor U2805 (N_2805,N_1362,N_1694);
or U2806 (N_2806,N_1818,N_1496);
nand U2807 (N_2807,N_1367,N_1475);
xor U2808 (N_2808,N_1567,N_1220);
nand U2809 (N_2809,N_1635,N_1907);
or U2810 (N_2810,N_1067,N_1470);
nor U2811 (N_2811,N_1943,N_1756);
xor U2812 (N_2812,N_1261,N_1359);
nand U2813 (N_2813,N_1008,N_1388);
or U2814 (N_2814,N_1194,N_1606);
nand U2815 (N_2815,N_1891,N_1139);
xor U2816 (N_2816,N_1377,N_1916);
and U2817 (N_2817,N_1172,N_1402);
nand U2818 (N_2818,N_1862,N_1844);
or U2819 (N_2819,N_1251,N_1956);
nor U2820 (N_2820,N_1892,N_1168);
nor U2821 (N_2821,N_1174,N_1465);
and U2822 (N_2822,N_1018,N_1283);
and U2823 (N_2823,N_1546,N_1849);
and U2824 (N_2824,N_1201,N_1805);
and U2825 (N_2825,N_1952,N_1719);
xor U2826 (N_2826,N_1971,N_1737);
or U2827 (N_2827,N_1145,N_1893);
and U2828 (N_2828,N_1619,N_1360);
or U2829 (N_2829,N_1899,N_1329);
nand U2830 (N_2830,N_1977,N_1867);
or U2831 (N_2831,N_1660,N_1171);
xnor U2832 (N_2832,N_1894,N_1421);
xor U2833 (N_2833,N_1111,N_1499);
xnor U2834 (N_2834,N_1309,N_1520);
xor U2835 (N_2835,N_1047,N_1671);
nor U2836 (N_2836,N_1598,N_1373);
and U2837 (N_2837,N_1742,N_1827);
and U2838 (N_2838,N_1659,N_1380);
nor U2839 (N_2839,N_1518,N_1084);
xor U2840 (N_2840,N_1685,N_1424);
nor U2841 (N_2841,N_1863,N_1625);
and U2842 (N_2842,N_1555,N_1675);
and U2843 (N_2843,N_1822,N_1195);
nor U2844 (N_2844,N_1572,N_1151);
or U2845 (N_2845,N_1967,N_1527);
nand U2846 (N_2846,N_1692,N_1482);
and U2847 (N_2847,N_1902,N_1315);
xnor U2848 (N_2848,N_1926,N_1185);
nand U2849 (N_2849,N_1491,N_1412);
nor U2850 (N_2850,N_1182,N_1118);
nand U2851 (N_2851,N_1207,N_1650);
nor U2852 (N_2852,N_1909,N_1310);
nand U2853 (N_2853,N_1308,N_1427);
or U2854 (N_2854,N_1644,N_1509);
xnor U2855 (N_2855,N_1722,N_1195);
nor U2856 (N_2856,N_1418,N_1048);
nand U2857 (N_2857,N_1098,N_1037);
or U2858 (N_2858,N_1574,N_1790);
xor U2859 (N_2859,N_1071,N_1765);
xnor U2860 (N_2860,N_1070,N_1888);
nand U2861 (N_2861,N_1926,N_1938);
and U2862 (N_2862,N_1891,N_1901);
xor U2863 (N_2863,N_1564,N_1437);
nand U2864 (N_2864,N_1853,N_1984);
or U2865 (N_2865,N_1197,N_1068);
and U2866 (N_2866,N_1114,N_1158);
xor U2867 (N_2867,N_1317,N_1208);
nor U2868 (N_2868,N_1146,N_1867);
nor U2869 (N_2869,N_1850,N_1776);
nor U2870 (N_2870,N_1737,N_1489);
and U2871 (N_2871,N_1901,N_1360);
nor U2872 (N_2872,N_1328,N_1973);
xor U2873 (N_2873,N_1957,N_1628);
xnor U2874 (N_2874,N_1018,N_1113);
nand U2875 (N_2875,N_1522,N_1107);
nor U2876 (N_2876,N_1209,N_1340);
nand U2877 (N_2877,N_1915,N_1421);
xnor U2878 (N_2878,N_1440,N_1913);
or U2879 (N_2879,N_1234,N_1445);
xor U2880 (N_2880,N_1366,N_1134);
nand U2881 (N_2881,N_1234,N_1004);
nand U2882 (N_2882,N_1045,N_1183);
xnor U2883 (N_2883,N_1859,N_1928);
nor U2884 (N_2884,N_1572,N_1111);
nor U2885 (N_2885,N_1005,N_1351);
xnor U2886 (N_2886,N_1588,N_1744);
nor U2887 (N_2887,N_1384,N_1122);
nor U2888 (N_2888,N_1513,N_1439);
and U2889 (N_2889,N_1401,N_1570);
nand U2890 (N_2890,N_1149,N_1059);
or U2891 (N_2891,N_1930,N_1335);
xor U2892 (N_2892,N_1145,N_1386);
nor U2893 (N_2893,N_1888,N_1047);
xor U2894 (N_2894,N_1998,N_1565);
nand U2895 (N_2895,N_1894,N_1044);
xor U2896 (N_2896,N_1201,N_1867);
nand U2897 (N_2897,N_1472,N_1298);
and U2898 (N_2898,N_1868,N_1303);
or U2899 (N_2899,N_1540,N_1140);
or U2900 (N_2900,N_1244,N_1874);
nor U2901 (N_2901,N_1638,N_1002);
nor U2902 (N_2902,N_1590,N_1428);
or U2903 (N_2903,N_1458,N_1781);
and U2904 (N_2904,N_1233,N_1467);
nor U2905 (N_2905,N_1873,N_1918);
xnor U2906 (N_2906,N_1883,N_1619);
nand U2907 (N_2907,N_1192,N_1734);
and U2908 (N_2908,N_1119,N_1075);
nor U2909 (N_2909,N_1897,N_1003);
and U2910 (N_2910,N_1771,N_1995);
nand U2911 (N_2911,N_1397,N_1106);
xnor U2912 (N_2912,N_1913,N_1594);
xor U2913 (N_2913,N_1038,N_1969);
or U2914 (N_2914,N_1981,N_1218);
nor U2915 (N_2915,N_1484,N_1660);
xor U2916 (N_2916,N_1279,N_1027);
nand U2917 (N_2917,N_1288,N_1598);
nand U2918 (N_2918,N_1703,N_1565);
and U2919 (N_2919,N_1408,N_1144);
and U2920 (N_2920,N_1969,N_1856);
or U2921 (N_2921,N_1681,N_1423);
nand U2922 (N_2922,N_1362,N_1300);
and U2923 (N_2923,N_1190,N_1811);
nand U2924 (N_2924,N_1451,N_1672);
xnor U2925 (N_2925,N_1953,N_1876);
xnor U2926 (N_2926,N_1003,N_1604);
xor U2927 (N_2927,N_1219,N_1154);
or U2928 (N_2928,N_1042,N_1896);
nor U2929 (N_2929,N_1803,N_1540);
nand U2930 (N_2930,N_1161,N_1631);
and U2931 (N_2931,N_1827,N_1694);
nor U2932 (N_2932,N_1535,N_1835);
xor U2933 (N_2933,N_1685,N_1438);
and U2934 (N_2934,N_1639,N_1700);
or U2935 (N_2935,N_1425,N_1453);
nor U2936 (N_2936,N_1607,N_1474);
nor U2937 (N_2937,N_1007,N_1240);
or U2938 (N_2938,N_1313,N_1761);
and U2939 (N_2939,N_1923,N_1548);
or U2940 (N_2940,N_1516,N_1920);
or U2941 (N_2941,N_1873,N_1735);
or U2942 (N_2942,N_1509,N_1963);
nand U2943 (N_2943,N_1624,N_1572);
nand U2944 (N_2944,N_1661,N_1009);
nand U2945 (N_2945,N_1242,N_1771);
nor U2946 (N_2946,N_1221,N_1203);
nor U2947 (N_2947,N_1303,N_1862);
xnor U2948 (N_2948,N_1282,N_1694);
xor U2949 (N_2949,N_1325,N_1789);
and U2950 (N_2950,N_1909,N_1388);
and U2951 (N_2951,N_1801,N_1729);
and U2952 (N_2952,N_1173,N_1756);
and U2953 (N_2953,N_1354,N_1410);
nand U2954 (N_2954,N_1424,N_1634);
nand U2955 (N_2955,N_1780,N_1271);
nor U2956 (N_2956,N_1620,N_1194);
xnor U2957 (N_2957,N_1570,N_1286);
xnor U2958 (N_2958,N_1697,N_1905);
nor U2959 (N_2959,N_1396,N_1611);
nand U2960 (N_2960,N_1498,N_1156);
xor U2961 (N_2961,N_1723,N_1144);
xnor U2962 (N_2962,N_1099,N_1401);
xor U2963 (N_2963,N_1900,N_1645);
xor U2964 (N_2964,N_1957,N_1635);
nor U2965 (N_2965,N_1559,N_1763);
or U2966 (N_2966,N_1780,N_1732);
nand U2967 (N_2967,N_1520,N_1067);
nor U2968 (N_2968,N_1126,N_1272);
nor U2969 (N_2969,N_1285,N_1107);
xor U2970 (N_2970,N_1871,N_1644);
or U2971 (N_2971,N_1602,N_1547);
or U2972 (N_2972,N_1548,N_1886);
xnor U2973 (N_2973,N_1877,N_1923);
nand U2974 (N_2974,N_1479,N_1491);
and U2975 (N_2975,N_1830,N_1623);
and U2976 (N_2976,N_1754,N_1659);
nor U2977 (N_2977,N_1598,N_1835);
and U2978 (N_2978,N_1136,N_1368);
xnor U2979 (N_2979,N_1337,N_1250);
nand U2980 (N_2980,N_1707,N_1726);
nand U2981 (N_2981,N_1232,N_1670);
and U2982 (N_2982,N_1340,N_1021);
nor U2983 (N_2983,N_1729,N_1512);
xnor U2984 (N_2984,N_1315,N_1978);
or U2985 (N_2985,N_1063,N_1629);
xnor U2986 (N_2986,N_1499,N_1520);
nor U2987 (N_2987,N_1483,N_1002);
nor U2988 (N_2988,N_1367,N_1670);
nor U2989 (N_2989,N_1207,N_1765);
xnor U2990 (N_2990,N_1261,N_1477);
nand U2991 (N_2991,N_1831,N_1232);
or U2992 (N_2992,N_1480,N_1117);
xnor U2993 (N_2993,N_1731,N_1935);
and U2994 (N_2994,N_1381,N_1223);
and U2995 (N_2995,N_1964,N_1686);
nand U2996 (N_2996,N_1994,N_1481);
nand U2997 (N_2997,N_1772,N_1827);
or U2998 (N_2998,N_1417,N_1249);
xor U2999 (N_2999,N_1849,N_1093);
nor U3000 (N_3000,N_2458,N_2041);
nand U3001 (N_3001,N_2779,N_2300);
or U3002 (N_3002,N_2942,N_2734);
and U3003 (N_3003,N_2375,N_2024);
or U3004 (N_3004,N_2586,N_2612);
and U3005 (N_3005,N_2422,N_2156);
nand U3006 (N_3006,N_2327,N_2040);
and U3007 (N_3007,N_2240,N_2569);
nand U3008 (N_3008,N_2725,N_2190);
or U3009 (N_3009,N_2393,N_2672);
or U3010 (N_3010,N_2133,N_2906);
or U3011 (N_3011,N_2247,N_2466);
nand U3012 (N_3012,N_2033,N_2526);
or U3013 (N_3013,N_2799,N_2490);
and U3014 (N_3014,N_2936,N_2955);
or U3015 (N_3015,N_2086,N_2241);
or U3016 (N_3016,N_2217,N_2435);
nor U3017 (N_3017,N_2394,N_2005);
nor U3018 (N_3018,N_2379,N_2320);
and U3019 (N_3019,N_2027,N_2447);
nand U3020 (N_3020,N_2186,N_2968);
xor U3021 (N_3021,N_2022,N_2673);
or U3022 (N_3022,N_2355,N_2460);
nand U3023 (N_3023,N_2016,N_2860);
nor U3024 (N_3024,N_2110,N_2908);
or U3025 (N_3025,N_2287,N_2341);
or U3026 (N_3026,N_2228,N_2486);
and U3027 (N_3027,N_2351,N_2824);
xnor U3028 (N_3028,N_2315,N_2622);
or U3029 (N_3029,N_2214,N_2887);
xor U3030 (N_3030,N_2209,N_2210);
and U3031 (N_3031,N_2218,N_2260);
and U3032 (N_3032,N_2505,N_2912);
and U3033 (N_3033,N_2522,N_2161);
xnor U3034 (N_3034,N_2083,N_2122);
nand U3035 (N_3035,N_2120,N_2098);
nor U3036 (N_3036,N_2378,N_2426);
nand U3037 (N_3037,N_2476,N_2380);
and U3038 (N_3038,N_2028,N_2763);
and U3039 (N_3039,N_2001,N_2094);
and U3040 (N_3040,N_2674,N_2761);
xor U3041 (N_3041,N_2463,N_2227);
nand U3042 (N_3042,N_2025,N_2642);
or U3043 (N_3043,N_2268,N_2875);
and U3044 (N_3044,N_2578,N_2439);
nor U3045 (N_3045,N_2332,N_2191);
nor U3046 (N_3046,N_2482,N_2830);
and U3047 (N_3047,N_2599,N_2529);
nand U3048 (N_3048,N_2694,N_2539);
or U3049 (N_3049,N_2407,N_2931);
xnor U3050 (N_3050,N_2981,N_2733);
and U3051 (N_3051,N_2941,N_2534);
and U3052 (N_3052,N_2996,N_2135);
or U3053 (N_3053,N_2183,N_2974);
or U3054 (N_3054,N_2283,N_2629);
nand U3055 (N_3055,N_2454,N_2455);
or U3056 (N_3056,N_2969,N_2967);
xnor U3057 (N_3057,N_2462,N_2596);
nand U3058 (N_3058,N_2913,N_2959);
xnor U3059 (N_3059,N_2618,N_2078);
or U3060 (N_3060,N_2411,N_2232);
nand U3061 (N_3061,N_2049,N_2438);
nor U3062 (N_3062,N_2817,N_2286);
nor U3063 (N_3063,N_2990,N_2508);
xnor U3064 (N_3064,N_2499,N_2834);
nor U3065 (N_3065,N_2859,N_2924);
xnor U3066 (N_3066,N_2984,N_2684);
and U3067 (N_3067,N_2690,N_2117);
nor U3068 (N_3068,N_2160,N_2928);
or U3069 (N_3069,N_2155,N_2747);
nor U3070 (N_3070,N_2713,N_2487);
nand U3071 (N_3071,N_2903,N_2671);
and U3072 (N_3072,N_2639,N_2518);
nor U3073 (N_3073,N_2153,N_2964);
xnor U3074 (N_3074,N_2440,N_2960);
xor U3075 (N_3075,N_2445,N_2347);
or U3076 (N_3076,N_2146,N_2769);
and U3077 (N_3077,N_2802,N_2349);
or U3078 (N_3078,N_2800,N_2853);
nor U3079 (N_3079,N_2279,N_2409);
nand U3080 (N_3080,N_2090,N_2292);
and U3081 (N_3081,N_2669,N_2691);
and U3082 (N_3082,N_2130,N_2388);
nor U3083 (N_3083,N_2843,N_2814);
or U3084 (N_3084,N_2771,N_2009);
or U3085 (N_3085,N_2000,N_2148);
and U3086 (N_3086,N_2550,N_2405);
nand U3087 (N_3087,N_2889,N_2970);
nand U3088 (N_3088,N_2291,N_2961);
nand U3089 (N_3089,N_2204,N_2265);
xnor U3090 (N_3090,N_2354,N_2589);
nor U3091 (N_3091,N_2991,N_2625);
nand U3092 (N_3092,N_2591,N_2610);
and U3093 (N_3093,N_2696,N_2939);
and U3094 (N_3094,N_2087,N_2716);
nand U3095 (N_3095,N_2770,N_2328);
nand U3096 (N_3096,N_2031,N_2184);
nand U3097 (N_3097,N_2558,N_2004);
nand U3098 (N_3098,N_2012,N_2679);
nor U3099 (N_3099,N_2850,N_2051);
xnor U3100 (N_3100,N_2623,N_2630);
and U3101 (N_3101,N_2188,N_2751);
or U3102 (N_3102,N_2609,N_2333);
xnor U3103 (N_3103,N_2963,N_2838);
nor U3104 (N_3104,N_2119,N_2917);
or U3105 (N_3105,N_2192,N_2057);
and U3106 (N_3106,N_2434,N_2074);
and U3107 (N_3107,N_2791,N_2541);
or U3108 (N_3108,N_2911,N_2901);
xnor U3109 (N_3109,N_2938,N_2864);
nor U3110 (N_3110,N_2429,N_2731);
nand U3111 (N_3111,N_2549,N_2922);
or U3112 (N_3112,N_2421,N_2880);
nor U3113 (N_3113,N_2506,N_2840);
and U3114 (N_3114,N_2556,N_2430);
nor U3115 (N_3115,N_2801,N_2876);
xnor U3116 (N_3116,N_2567,N_2267);
nand U3117 (N_3117,N_2198,N_2857);
and U3118 (N_3118,N_2477,N_2396);
xor U3119 (N_3119,N_2348,N_2251);
nand U3120 (N_3120,N_2898,N_2593);
and U3121 (N_3121,N_2493,N_2091);
xnor U3122 (N_3122,N_2510,N_2965);
or U3123 (N_3123,N_2104,N_2785);
and U3124 (N_3124,N_2134,N_2836);
and U3125 (N_3125,N_2252,N_2322);
nand U3126 (N_3126,N_2065,N_2758);
nor U3127 (N_3127,N_2858,N_2688);
nand U3128 (N_3128,N_2902,N_2592);
or U3129 (N_3129,N_2196,N_2531);
or U3130 (N_3130,N_2743,N_2158);
nor U3131 (N_3131,N_2754,N_2281);
or U3132 (N_3132,N_2359,N_2194);
or U3133 (N_3133,N_2900,N_2606);
xnor U3134 (N_3134,N_2512,N_2331);
nand U3135 (N_3135,N_2737,N_2095);
nor U3136 (N_3136,N_2552,N_2709);
and U3137 (N_3137,N_2473,N_2695);
nand U3138 (N_3138,N_2835,N_2285);
and U3139 (N_3139,N_2132,N_2516);
or U3140 (N_3140,N_2631,N_2269);
nor U3141 (N_3141,N_2813,N_2804);
or U3142 (N_3142,N_2573,N_2329);
xor U3143 (N_3143,N_2114,N_2551);
or U3144 (N_3144,N_2729,N_2264);
or U3145 (N_3145,N_2073,N_2746);
nor U3146 (N_3146,N_2402,N_2271);
xor U3147 (N_3147,N_2920,N_2822);
or U3148 (N_3148,N_2019,N_2823);
or U3149 (N_3149,N_2878,N_2828);
nand U3150 (N_3150,N_2123,N_2256);
or U3151 (N_3151,N_2140,N_2220);
or U3152 (N_3152,N_2075,N_2389);
and U3153 (N_3153,N_2777,N_2284);
and U3154 (N_3154,N_2766,N_2614);
nor U3155 (N_3155,N_2459,N_2701);
nand U3156 (N_3156,N_2432,N_2185);
xnor U3157 (N_3157,N_2760,N_2142);
nand U3158 (N_3158,N_2635,N_2683);
xnor U3159 (N_3159,N_2894,N_2979);
nand U3160 (N_3160,N_2298,N_2837);
nor U3161 (N_3161,N_2374,N_2561);
or U3162 (N_3162,N_2598,N_2798);
xnor U3163 (N_3163,N_2293,N_2262);
nor U3164 (N_3164,N_2603,N_2316);
and U3165 (N_3165,N_2195,N_2170);
or U3166 (N_3166,N_2020,N_2239);
and U3167 (N_3167,N_2932,N_2301);
xor U3168 (N_3168,N_2403,N_2994);
nand U3169 (N_3169,N_2141,N_2047);
or U3170 (N_3170,N_2854,N_2096);
or U3171 (N_3171,N_2431,N_2414);
nand U3172 (N_3172,N_2011,N_2352);
nand U3173 (N_3173,N_2621,N_2719);
xnor U3174 (N_3174,N_2682,N_2494);
or U3175 (N_3175,N_2615,N_2034);
nand U3176 (N_3176,N_2590,N_2736);
and U3177 (N_3177,N_2226,N_2517);
xor U3178 (N_3178,N_2415,N_2562);
or U3179 (N_3179,N_2883,N_2907);
or U3180 (N_3180,N_2829,N_2233);
nand U3181 (N_3181,N_2579,N_2225);
and U3182 (N_3182,N_2200,N_2501);
xnor U3183 (N_3183,N_2498,N_2069);
and U3184 (N_3184,N_2923,N_2207);
and U3185 (N_3185,N_2786,N_2915);
xnor U3186 (N_3186,N_2594,N_2803);
xnor U3187 (N_3187,N_2360,N_2270);
or U3188 (N_3188,N_2735,N_2958);
nand U3189 (N_3189,N_2076,N_2787);
nor U3190 (N_3190,N_2987,N_2068);
nand U3191 (N_3191,N_2103,N_2066);
xor U3192 (N_3192,N_2503,N_2784);
nor U3193 (N_3193,N_2825,N_2914);
nor U3194 (N_3194,N_2282,N_2833);
nand U3195 (N_3195,N_2115,N_2436);
and U3196 (N_3196,N_2201,N_2324);
nand U3197 (N_3197,N_2753,N_2367);
xor U3198 (N_3198,N_2966,N_2852);
xor U3199 (N_3199,N_2179,N_2229);
xor U3200 (N_3200,N_2157,N_2916);
and U3201 (N_3201,N_2037,N_2111);
nor U3202 (N_3202,N_2613,N_2313);
nand U3203 (N_3203,N_2790,N_2178);
nand U3204 (N_3204,N_2846,N_2259);
xor U3205 (N_3205,N_2236,N_2385);
xor U3206 (N_3206,N_2481,N_2106);
xnor U3207 (N_3207,N_2988,N_2006);
xor U3208 (N_3208,N_2126,N_2205);
nor U3209 (N_3209,N_2774,N_2253);
nor U3210 (N_3210,N_2151,N_2152);
nand U3211 (N_3211,N_2577,N_2794);
and U3212 (N_3212,N_2404,N_2693);
xnor U3213 (N_3213,N_2278,N_2017);
nand U3214 (N_3214,N_2867,N_2149);
xnor U3215 (N_3215,N_2100,N_2206);
and U3216 (N_3216,N_2277,N_2419);
xor U3217 (N_3217,N_2811,N_2545);
and U3218 (N_3218,N_2084,N_2972);
nor U3219 (N_3219,N_2021,N_2125);
and U3220 (N_3220,N_2321,N_2056);
nor U3221 (N_3221,N_2273,N_2678);
nand U3222 (N_3222,N_2408,N_2399);
or U3223 (N_3223,N_2985,N_2871);
xnor U3224 (N_3224,N_2237,N_2035);
and U3225 (N_3225,N_2711,N_2309);
or U3226 (N_3226,N_2457,N_2652);
and U3227 (N_3227,N_2202,N_2842);
nand U3228 (N_3228,N_2870,N_2707);
xnor U3229 (N_3229,N_2536,N_2532);
xor U3230 (N_3230,N_2654,N_2274);
and U3231 (N_3231,N_2182,N_2509);
xnor U3232 (N_3232,N_2334,N_2128);
and U3233 (N_3233,N_2116,N_2013);
nor U3234 (N_3234,N_2139,N_2296);
and U3235 (N_3235,N_2492,N_2865);
and U3236 (N_3236,N_2423,N_2946);
or U3237 (N_3237,N_2193,N_2446);
nand U3238 (N_3238,N_2101,N_2497);
nand U3239 (N_3239,N_2645,N_2243);
and U3240 (N_3240,N_2588,N_2951);
nand U3241 (N_3241,N_2118,N_2620);
or U3242 (N_3242,N_2628,N_2370);
nor U3243 (N_3243,N_2189,N_2929);
or U3244 (N_3244,N_2372,N_2400);
or U3245 (N_3245,N_2741,N_2926);
nand U3246 (N_3246,N_2525,N_2995);
and U3247 (N_3247,N_2093,N_2676);
nor U3248 (N_3248,N_2659,N_2720);
nor U3249 (N_3249,N_2597,N_2235);
and U3250 (N_3250,N_2748,N_2732);
xnor U3251 (N_3251,N_2401,N_2983);
and U3252 (N_3252,N_2927,N_2892);
and U3253 (N_3253,N_2305,N_2410);
or U3254 (N_3254,N_2595,N_2956);
or U3255 (N_3255,N_2350,N_2658);
or U3256 (N_3256,N_2085,N_2780);
xor U3257 (N_3257,N_2167,N_2147);
or U3258 (N_3258,N_2042,N_2336);
nand U3259 (N_3259,N_2877,N_2976);
nor U3260 (N_3260,N_2893,N_2258);
nand U3261 (N_3261,N_2949,N_2993);
nor U3262 (N_3262,N_2986,N_2882);
or U3263 (N_3263,N_2699,N_2863);
nor U3264 (N_3264,N_2166,N_2089);
nor U3265 (N_3265,N_2063,N_2797);
nand U3266 (N_3266,N_2727,N_2039);
nor U3267 (N_3267,N_2570,N_2982);
xor U3268 (N_3268,N_2055,N_2181);
nand U3269 (N_3269,N_2003,N_2121);
nand U3270 (N_3270,N_2587,N_2318);
nand U3271 (N_3271,N_2472,N_2077);
nor U3272 (N_3272,N_2943,N_2685);
xor U3273 (N_3273,N_2353,N_2897);
nand U3274 (N_3274,N_2948,N_2624);
nor U3275 (N_3275,N_2715,N_2789);
and U3276 (N_3276,N_2323,N_2947);
xor U3277 (N_3277,N_2261,N_2124);
nor U3278 (N_3278,N_2187,N_2918);
and U3279 (N_3279,N_2879,N_2461);
or U3280 (N_3280,N_2317,N_2010);
and U3281 (N_3281,N_2046,N_2255);
and U3282 (N_3282,N_2881,N_2560);
xnor U3283 (N_3283,N_2962,N_2832);
nand U3284 (N_3284,N_2450,N_2627);
xor U3285 (N_3285,N_2776,N_2812);
nor U3286 (N_3286,N_2150,N_2504);
nand U3287 (N_3287,N_2029,N_2538);
xnor U3288 (N_3288,N_2957,N_2368);
xnor U3289 (N_3289,N_2997,N_2795);
nor U3290 (N_3290,N_2637,N_2809);
xnor U3291 (N_3291,N_2129,N_2174);
or U3292 (N_3292,N_2062,N_2444);
nand U3293 (N_3293,N_2921,N_2827);
nor U3294 (N_3294,N_2925,N_2088);
and U3295 (N_3295,N_2783,N_2714);
xnor U3296 (N_3296,N_2050,N_2663);
nand U3297 (N_3297,N_2548,N_2706);
and U3298 (N_3298,N_2513,N_2565);
nor U3299 (N_3299,N_2173,N_2632);
or U3300 (N_3300,N_2306,N_2805);
or U3301 (N_3301,N_2032,N_2165);
xor U3302 (N_3302,N_2940,N_2759);
or U3303 (N_3303,N_2666,N_2464);
or U3304 (N_3304,N_2199,N_2263);
and U3305 (N_3305,N_2775,N_2818);
nand U3306 (N_3306,N_2417,N_2527);
nand U3307 (N_3307,N_2427,N_2030);
or U3308 (N_3308,N_2819,N_2749);
and U3309 (N_3309,N_2081,N_2773);
or U3310 (N_3310,N_2471,N_2048);
or U3311 (N_3311,N_2668,N_2862);
and U3312 (N_3312,N_2568,N_2339);
nand U3313 (N_3313,N_2700,N_2977);
nand U3314 (N_3314,N_2395,N_2215);
nor U3315 (N_3315,N_2026,N_2249);
xnor U3316 (N_3316,N_2738,N_2954);
or U3317 (N_3317,N_2781,N_2250);
nand U3318 (N_3318,N_2045,N_2514);
xnor U3319 (N_3319,N_2014,N_2238);
and U3320 (N_3320,N_2782,N_2757);
xnor U3321 (N_3321,N_2392,N_2177);
or U3322 (N_3322,N_2154,N_2722);
nand U3323 (N_3323,N_2665,N_2145);
nand U3324 (N_3324,N_2762,N_2554);
or U3325 (N_3325,N_2869,N_2180);
nand U3326 (N_3326,N_2107,N_2888);
or U3327 (N_3327,N_2099,N_2686);
and U3328 (N_3328,N_2677,N_2386);
nor U3329 (N_3329,N_2953,N_2102);
and U3330 (N_3330,N_2484,N_2272);
and U3331 (N_3331,N_2650,N_2697);
nor U3332 (N_3332,N_2895,N_2788);
nand U3333 (N_3333,N_2608,N_2752);
or U3334 (N_3334,N_2266,N_2197);
nor U3335 (N_3335,N_2257,N_2750);
or U3336 (N_3336,N_2528,N_2377);
or U3337 (N_3337,N_2998,N_2079);
nand U3338 (N_3338,N_2520,N_2744);
nand U3339 (N_3339,N_2643,N_2335);
or U3340 (N_3340,N_2467,N_2885);
and U3341 (N_3341,N_2364,N_2043);
nand U3342 (N_3342,N_2213,N_2581);
nor U3343 (N_3343,N_2474,N_2952);
xor U3344 (N_3344,N_2601,N_2163);
nand U3345 (N_3345,N_2564,N_2764);
xnor U3346 (N_3346,N_2535,N_2136);
nor U3347 (N_3347,N_2537,N_2245);
xnor U3348 (N_3348,N_2905,N_2162);
xnor U3349 (N_3349,N_2168,N_2176);
nand U3350 (N_3350,N_2097,N_2469);
nand U3351 (N_3351,N_2058,N_2297);
xor U3352 (N_3352,N_2648,N_2244);
or U3353 (N_3353,N_2935,N_2007);
and U3354 (N_3354,N_2992,N_2294);
nand U3355 (N_3355,N_2708,N_2755);
and U3356 (N_3356,N_2383,N_2515);
or U3357 (N_3357,N_2018,N_2710);
xnor U3358 (N_3358,N_2675,N_2059);
nand U3359 (N_3359,N_2611,N_2127);
or U3360 (N_3360,N_2203,N_2616);
and U3361 (N_3361,N_2910,N_2826);
xor U3362 (N_3362,N_2299,N_2670);
xnor U3363 (N_3363,N_2646,N_2172);
or U3364 (N_3364,N_2574,N_2765);
nand U3365 (N_3365,N_2061,N_2680);
nor U3366 (N_3366,N_2023,N_2387);
and U3367 (N_3367,N_2989,N_2390);
nor U3368 (N_3368,N_2502,N_2999);
or U3369 (N_3369,N_2739,N_2756);
nor U3370 (N_3370,N_2718,N_2808);
and U3371 (N_3371,N_2656,N_2290);
nand U3372 (N_3372,N_2507,N_2767);
or U3373 (N_3373,N_2978,N_2662);
or U3374 (N_3374,N_2726,N_2617);
or U3375 (N_3375,N_2070,N_2868);
nand U3376 (N_3376,N_2137,N_2072);
or U3377 (N_3377,N_2071,N_2366);
and U3378 (N_3378,N_2816,N_2944);
nand U3379 (N_3379,N_2314,N_2636);
nor U3380 (N_3380,N_2357,N_2479);
xor U3381 (N_3381,N_2138,N_2358);
nand U3382 (N_3382,N_2443,N_2638);
nand U3383 (N_3383,N_2008,N_2442);
and U3384 (N_3384,N_2856,N_2778);
nor U3385 (N_3385,N_2742,N_2391);
nand U3386 (N_3386,N_2651,N_2343);
and U3387 (N_3387,N_2772,N_2304);
nor U3388 (N_3388,N_2376,N_2219);
xnor U3389 (N_3389,N_2950,N_2566);
nand U3390 (N_3390,N_2483,N_2563);
nand U3391 (N_3391,N_2530,N_2855);
xnor U3392 (N_3392,N_2441,N_2480);
nand U3393 (N_3393,N_2052,N_2821);
xor U3394 (N_3394,N_2433,N_2325);
or U3395 (N_3395,N_2082,N_2524);
and U3396 (N_3396,N_2839,N_2064);
nand U3397 (N_3397,N_2555,N_2092);
or U3398 (N_3398,N_2872,N_2724);
xor U3399 (N_3399,N_2848,N_2308);
and U3400 (N_3400,N_2345,N_2080);
and U3401 (N_3401,N_2382,N_2208);
nor U3402 (N_3402,N_2730,N_2649);
nor U3403 (N_3403,N_2425,N_2934);
nand U3404 (N_3404,N_2740,N_2640);
nand U3405 (N_3405,N_2311,N_2221);
and U3406 (N_3406,N_2807,N_2831);
xnor U3407 (N_3407,N_2216,N_2661);
nand U3408 (N_3408,N_2044,N_2413);
nand U3409 (N_3409,N_2511,N_2849);
nor U3410 (N_3410,N_2891,N_2820);
and U3411 (N_3411,N_2428,N_2346);
nor U3412 (N_3412,N_2144,N_2576);
nor U3413 (N_3413,N_2519,N_2384);
nor U3414 (N_3414,N_2692,N_2557);
and U3415 (N_3415,N_2488,N_2397);
nor U3416 (N_3416,N_2626,N_2131);
or U3417 (N_3417,N_2036,N_2164);
and U3418 (N_3418,N_2312,N_2448);
or U3419 (N_3419,N_2605,N_2424);
nor U3420 (N_3420,N_2641,N_2703);
and U3421 (N_3421,N_2365,N_2681);
and U3422 (N_3422,N_2234,N_2361);
xor U3423 (N_3423,N_2723,N_2851);
nor U3424 (N_3424,N_2452,N_2337);
or U3425 (N_3425,N_2288,N_2105);
or U3426 (N_3426,N_2371,N_2582);
and U3427 (N_3427,N_2246,N_2543);
nand U3428 (N_3428,N_2212,N_2108);
nor U3429 (N_3429,N_2810,N_2584);
and U3430 (N_3430,N_2705,N_2698);
or U3431 (N_3431,N_2873,N_2874);
nand U3432 (N_3432,N_2418,N_2398);
and U3433 (N_3433,N_2815,N_2175);
and U3434 (N_3434,N_2362,N_2721);
or U3435 (N_3435,N_2844,N_2495);
and U3436 (N_3436,N_2971,N_2619);
xnor U3437 (N_3437,N_2523,N_2053);
nor U3438 (N_3438,N_2465,N_2571);
nor U3439 (N_3439,N_2276,N_2067);
and U3440 (N_3440,N_2806,N_2542);
nand U3441 (N_3441,N_2224,N_2223);
xnor U3442 (N_3442,N_2230,N_2449);
and U3443 (N_3443,N_2406,N_2717);
nor U3444 (N_3444,N_2633,N_2704);
xor U3445 (N_3445,N_2338,N_2886);
xor U3446 (N_3446,N_2470,N_2687);
nand U3447 (N_3447,N_2899,N_2275);
nor U3448 (N_3448,N_2585,N_2973);
xor U3449 (N_3449,N_2496,N_2468);
nor U3450 (N_3450,N_2453,N_2657);
or U3451 (N_3451,N_2211,N_2344);
and U3452 (N_3452,N_2792,N_2572);
or U3453 (N_3453,N_2054,N_2745);
nor U3454 (N_3454,N_2500,N_2546);
nor U3455 (N_3455,N_2112,N_2109);
or U3456 (N_3456,N_2451,N_2478);
xor U3457 (N_3457,N_2363,N_2607);
nor U3458 (N_3458,N_2420,N_2667);
xnor U3459 (N_3459,N_2412,N_2060);
and U3460 (N_3460,N_2600,N_2544);
nand U3461 (N_3461,N_2583,N_2647);
nor U3462 (N_3462,N_2303,N_2289);
and U3463 (N_3463,N_2655,N_2793);
and U3464 (N_3464,N_2475,N_2373);
nor U3465 (N_3465,N_2307,N_2310);
or U3466 (N_3466,N_2861,N_2159);
or U3467 (N_3467,N_2171,N_2847);
xor U3468 (N_3468,N_2340,N_2521);
and U3469 (N_3469,N_2456,N_2896);
xor U3470 (N_3470,N_2330,N_2002);
xnor U3471 (N_3471,N_2437,N_2945);
xnor U3472 (N_3472,N_2845,N_2919);
nand U3473 (N_3473,N_2890,N_2559);
xor U3474 (N_3474,N_2866,N_2664);
xor U3475 (N_3475,N_2295,N_2602);
nand U3476 (N_3476,N_2796,N_2319);
and U3477 (N_3477,N_2689,N_2015);
nand U3478 (N_3478,N_2485,N_2937);
and U3479 (N_3479,N_2533,N_2381);
or U3480 (N_3480,N_2604,N_2768);
and U3481 (N_3481,N_2660,N_2547);
xnor U3482 (N_3482,N_2248,N_2143);
or U3483 (N_3483,N_2909,N_2231);
nor U3484 (N_3484,N_2113,N_2644);
nor U3485 (N_3485,N_2653,N_2728);
nor U3486 (N_3486,N_2342,N_2634);
xnor U3487 (N_3487,N_2326,N_2169);
nor U3488 (N_3488,N_2491,N_2930);
xor U3489 (N_3489,N_2933,N_2980);
nand U3490 (N_3490,N_2975,N_2369);
and U3491 (N_3491,N_2280,N_2302);
nand U3492 (N_3492,N_2553,N_2702);
xnor U3493 (N_3493,N_2222,N_2356);
nand U3494 (N_3494,N_2712,N_2841);
nor U3495 (N_3495,N_2904,N_2254);
nand U3496 (N_3496,N_2242,N_2575);
and U3497 (N_3497,N_2489,N_2416);
xor U3498 (N_3498,N_2540,N_2580);
and U3499 (N_3499,N_2038,N_2884);
or U3500 (N_3500,N_2319,N_2884);
nand U3501 (N_3501,N_2100,N_2735);
nand U3502 (N_3502,N_2014,N_2050);
or U3503 (N_3503,N_2425,N_2792);
or U3504 (N_3504,N_2710,N_2040);
and U3505 (N_3505,N_2208,N_2193);
nand U3506 (N_3506,N_2806,N_2225);
xnor U3507 (N_3507,N_2681,N_2363);
and U3508 (N_3508,N_2479,N_2035);
nand U3509 (N_3509,N_2257,N_2303);
or U3510 (N_3510,N_2008,N_2475);
nor U3511 (N_3511,N_2377,N_2077);
or U3512 (N_3512,N_2350,N_2748);
and U3513 (N_3513,N_2054,N_2004);
xnor U3514 (N_3514,N_2795,N_2497);
and U3515 (N_3515,N_2418,N_2900);
nand U3516 (N_3516,N_2600,N_2151);
or U3517 (N_3517,N_2975,N_2715);
or U3518 (N_3518,N_2028,N_2454);
xnor U3519 (N_3519,N_2433,N_2836);
and U3520 (N_3520,N_2127,N_2047);
xor U3521 (N_3521,N_2986,N_2052);
and U3522 (N_3522,N_2747,N_2044);
nand U3523 (N_3523,N_2965,N_2438);
nand U3524 (N_3524,N_2573,N_2775);
nor U3525 (N_3525,N_2856,N_2267);
nand U3526 (N_3526,N_2051,N_2011);
nand U3527 (N_3527,N_2831,N_2305);
or U3528 (N_3528,N_2705,N_2498);
and U3529 (N_3529,N_2685,N_2060);
and U3530 (N_3530,N_2032,N_2926);
nor U3531 (N_3531,N_2742,N_2901);
xor U3532 (N_3532,N_2019,N_2807);
nand U3533 (N_3533,N_2079,N_2083);
and U3534 (N_3534,N_2524,N_2722);
xor U3535 (N_3535,N_2921,N_2303);
nand U3536 (N_3536,N_2921,N_2876);
or U3537 (N_3537,N_2480,N_2979);
nor U3538 (N_3538,N_2374,N_2010);
nand U3539 (N_3539,N_2079,N_2885);
nor U3540 (N_3540,N_2712,N_2177);
or U3541 (N_3541,N_2026,N_2782);
and U3542 (N_3542,N_2739,N_2695);
nor U3543 (N_3543,N_2115,N_2823);
and U3544 (N_3544,N_2153,N_2960);
or U3545 (N_3545,N_2723,N_2557);
or U3546 (N_3546,N_2091,N_2753);
nor U3547 (N_3547,N_2090,N_2566);
xnor U3548 (N_3548,N_2060,N_2829);
or U3549 (N_3549,N_2100,N_2126);
nand U3550 (N_3550,N_2116,N_2917);
or U3551 (N_3551,N_2263,N_2031);
nor U3552 (N_3552,N_2951,N_2212);
or U3553 (N_3553,N_2021,N_2570);
nand U3554 (N_3554,N_2808,N_2198);
or U3555 (N_3555,N_2638,N_2028);
xnor U3556 (N_3556,N_2862,N_2926);
or U3557 (N_3557,N_2765,N_2037);
and U3558 (N_3558,N_2932,N_2953);
nor U3559 (N_3559,N_2283,N_2935);
and U3560 (N_3560,N_2100,N_2268);
nor U3561 (N_3561,N_2977,N_2567);
xor U3562 (N_3562,N_2079,N_2152);
or U3563 (N_3563,N_2960,N_2410);
nor U3564 (N_3564,N_2864,N_2647);
or U3565 (N_3565,N_2085,N_2824);
or U3566 (N_3566,N_2729,N_2420);
nor U3567 (N_3567,N_2615,N_2599);
nand U3568 (N_3568,N_2313,N_2621);
or U3569 (N_3569,N_2371,N_2181);
xor U3570 (N_3570,N_2518,N_2538);
nor U3571 (N_3571,N_2662,N_2532);
nand U3572 (N_3572,N_2022,N_2992);
and U3573 (N_3573,N_2639,N_2673);
nand U3574 (N_3574,N_2986,N_2519);
nor U3575 (N_3575,N_2726,N_2078);
xor U3576 (N_3576,N_2372,N_2426);
xor U3577 (N_3577,N_2518,N_2590);
and U3578 (N_3578,N_2996,N_2195);
or U3579 (N_3579,N_2205,N_2590);
nand U3580 (N_3580,N_2488,N_2454);
or U3581 (N_3581,N_2155,N_2692);
or U3582 (N_3582,N_2639,N_2495);
nor U3583 (N_3583,N_2450,N_2673);
and U3584 (N_3584,N_2144,N_2021);
and U3585 (N_3585,N_2306,N_2136);
or U3586 (N_3586,N_2202,N_2216);
xnor U3587 (N_3587,N_2045,N_2360);
nor U3588 (N_3588,N_2727,N_2624);
nor U3589 (N_3589,N_2979,N_2989);
nand U3590 (N_3590,N_2883,N_2839);
and U3591 (N_3591,N_2519,N_2615);
nand U3592 (N_3592,N_2665,N_2950);
nand U3593 (N_3593,N_2428,N_2797);
nand U3594 (N_3594,N_2497,N_2755);
xnor U3595 (N_3595,N_2212,N_2132);
or U3596 (N_3596,N_2660,N_2340);
or U3597 (N_3597,N_2196,N_2297);
or U3598 (N_3598,N_2028,N_2871);
or U3599 (N_3599,N_2643,N_2786);
and U3600 (N_3600,N_2197,N_2501);
nor U3601 (N_3601,N_2903,N_2407);
nor U3602 (N_3602,N_2085,N_2636);
nor U3603 (N_3603,N_2511,N_2049);
xnor U3604 (N_3604,N_2108,N_2664);
or U3605 (N_3605,N_2090,N_2841);
nand U3606 (N_3606,N_2145,N_2209);
nand U3607 (N_3607,N_2634,N_2983);
and U3608 (N_3608,N_2584,N_2436);
nor U3609 (N_3609,N_2924,N_2350);
nor U3610 (N_3610,N_2732,N_2323);
nor U3611 (N_3611,N_2496,N_2799);
or U3612 (N_3612,N_2402,N_2265);
nand U3613 (N_3613,N_2898,N_2156);
nor U3614 (N_3614,N_2392,N_2733);
nor U3615 (N_3615,N_2601,N_2593);
nor U3616 (N_3616,N_2230,N_2580);
nand U3617 (N_3617,N_2352,N_2320);
nor U3618 (N_3618,N_2369,N_2508);
nor U3619 (N_3619,N_2521,N_2199);
nor U3620 (N_3620,N_2852,N_2455);
nand U3621 (N_3621,N_2809,N_2562);
and U3622 (N_3622,N_2184,N_2740);
or U3623 (N_3623,N_2145,N_2586);
xnor U3624 (N_3624,N_2719,N_2740);
and U3625 (N_3625,N_2748,N_2286);
or U3626 (N_3626,N_2676,N_2495);
nor U3627 (N_3627,N_2443,N_2549);
nor U3628 (N_3628,N_2495,N_2059);
or U3629 (N_3629,N_2519,N_2817);
xor U3630 (N_3630,N_2749,N_2131);
xnor U3631 (N_3631,N_2209,N_2160);
xor U3632 (N_3632,N_2105,N_2586);
xnor U3633 (N_3633,N_2598,N_2444);
or U3634 (N_3634,N_2815,N_2919);
nor U3635 (N_3635,N_2479,N_2625);
nand U3636 (N_3636,N_2191,N_2171);
nor U3637 (N_3637,N_2704,N_2121);
and U3638 (N_3638,N_2195,N_2159);
nand U3639 (N_3639,N_2775,N_2597);
xnor U3640 (N_3640,N_2055,N_2182);
nand U3641 (N_3641,N_2613,N_2293);
xnor U3642 (N_3642,N_2693,N_2846);
xor U3643 (N_3643,N_2433,N_2813);
xnor U3644 (N_3644,N_2348,N_2057);
xnor U3645 (N_3645,N_2803,N_2232);
xor U3646 (N_3646,N_2648,N_2823);
xnor U3647 (N_3647,N_2648,N_2879);
or U3648 (N_3648,N_2636,N_2005);
or U3649 (N_3649,N_2051,N_2121);
xnor U3650 (N_3650,N_2229,N_2938);
nor U3651 (N_3651,N_2843,N_2211);
nor U3652 (N_3652,N_2128,N_2994);
and U3653 (N_3653,N_2454,N_2713);
or U3654 (N_3654,N_2694,N_2829);
nand U3655 (N_3655,N_2168,N_2601);
nand U3656 (N_3656,N_2516,N_2185);
or U3657 (N_3657,N_2281,N_2838);
xnor U3658 (N_3658,N_2464,N_2344);
and U3659 (N_3659,N_2642,N_2991);
nand U3660 (N_3660,N_2896,N_2638);
or U3661 (N_3661,N_2391,N_2822);
or U3662 (N_3662,N_2738,N_2167);
or U3663 (N_3663,N_2800,N_2869);
xnor U3664 (N_3664,N_2602,N_2866);
and U3665 (N_3665,N_2311,N_2501);
xor U3666 (N_3666,N_2999,N_2116);
or U3667 (N_3667,N_2478,N_2361);
xor U3668 (N_3668,N_2535,N_2489);
nand U3669 (N_3669,N_2150,N_2228);
or U3670 (N_3670,N_2741,N_2805);
or U3671 (N_3671,N_2711,N_2508);
nor U3672 (N_3672,N_2722,N_2327);
nand U3673 (N_3673,N_2894,N_2553);
nor U3674 (N_3674,N_2601,N_2913);
nor U3675 (N_3675,N_2010,N_2748);
xnor U3676 (N_3676,N_2240,N_2838);
and U3677 (N_3677,N_2642,N_2624);
nand U3678 (N_3678,N_2698,N_2067);
nand U3679 (N_3679,N_2495,N_2954);
or U3680 (N_3680,N_2848,N_2646);
nand U3681 (N_3681,N_2515,N_2027);
xnor U3682 (N_3682,N_2964,N_2727);
nand U3683 (N_3683,N_2036,N_2632);
nand U3684 (N_3684,N_2859,N_2976);
xnor U3685 (N_3685,N_2408,N_2313);
and U3686 (N_3686,N_2286,N_2755);
and U3687 (N_3687,N_2140,N_2295);
xor U3688 (N_3688,N_2383,N_2503);
and U3689 (N_3689,N_2663,N_2526);
nand U3690 (N_3690,N_2310,N_2583);
or U3691 (N_3691,N_2501,N_2791);
nor U3692 (N_3692,N_2725,N_2528);
and U3693 (N_3693,N_2907,N_2361);
xnor U3694 (N_3694,N_2737,N_2217);
or U3695 (N_3695,N_2467,N_2743);
nand U3696 (N_3696,N_2809,N_2752);
nand U3697 (N_3697,N_2094,N_2756);
or U3698 (N_3698,N_2697,N_2257);
nor U3699 (N_3699,N_2259,N_2643);
or U3700 (N_3700,N_2001,N_2718);
nor U3701 (N_3701,N_2889,N_2676);
or U3702 (N_3702,N_2337,N_2567);
and U3703 (N_3703,N_2324,N_2059);
nor U3704 (N_3704,N_2876,N_2234);
nand U3705 (N_3705,N_2331,N_2476);
xor U3706 (N_3706,N_2792,N_2290);
nor U3707 (N_3707,N_2852,N_2206);
nor U3708 (N_3708,N_2975,N_2461);
or U3709 (N_3709,N_2258,N_2789);
nand U3710 (N_3710,N_2905,N_2434);
xnor U3711 (N_3711,N_2199,N_2235);
nor U3712 (N_3712,N_2706,N_2253);
or U3713 (N_3713,N_2034,N_2172);
xor U3714 (N_3714,N_2731,N_2391);
nor U3715 (N_3715,N_2170,N_2234);
or U3716 (N_3716,N_2872,N_2292);
or U3717 (N_3717,N_2293,N_2920);
nand U3718 (N_3718,N_2824,N_2668);
or U3719 (N_3719,N_2340,N_2846);
xor U3720 (N_3720,N_2699,N_2199);
and U3721 (N_3721,N_2136,N_2130);
or U3722 (N_3722,N_2489,N_2760);
xor U3723 (N_3723,N_2455,N_2642);
and U3724 (N_3724,N_2375,N_2035);
or U3725 (N_3725,N_2431,N_2411);
nor U3726 (N_3726,N_2669,N_2630);
or U3727 (N_3727,N_2868,N_2799);
nand U3728 (N_3728,N_2382,N_2870);
nand U3729 (N_3729,N_2842,N_2213);
nand U3730 (N_3730,N_2698,N_2525);
nor U3731 (N_3731,N_2710,N_2412);
or U3732 (N_3732,N_2252,N_2133);
nor U3733 (N_3733,N_2372,N_2379);
and U3734 (N_3734,N_2917,N_2409);
nor U3735 (N_3735,N_2354,N_2298);
and U3736 (N_3736,N_2054,N_2935);
nand U3737 (N_3737,N_2539,N_2013);
nand U3738 (N_3738,N_2478,N_2679);
nand U3739 (N_3739,N_2151,N_2109);
nor U3740 (N_3740,N_2261,N_2868);
and U3741 (N_3741,N_2785,N_2363);
xor U3742 (N_3742,N_2492,N_2748);
nand U3743 (N_3743,N_2795,N_2821);
xnor U3744 (N_3744,N_2796,N_2417);
nor U3745 (N_3745,N_2684,N_2076);
nand U3746 (N_3746,N_2231,N_2069);
and U3747 (N_3747,N_2924,N_2194);
and U3748 (N_3748,N_2418,N_2343);
and U3749 (N_3749,N_2605,N_2833);
and U3750 (N_3750,N_2584,N_2126);
xor U3751 (N_3751,N_2400,N_2737);
xnor U3752 (N_3752,N_2838,N_2564);
and U3753 (N_3753,N_2316,N_2987);
nor U3754 (N_3754,N_2735,N_2647);
and U3755 (N_3755,N_2456,N_2505);
or U3756 (N_3756,N_2716,N_2586);
or U3757 (N_3757,N_2793,N_2958);
and U3758 (N_3758,N_2127,N_2146);
nand U3759 (N_3759,N_2253,N_2860);
nand U3760 (N_3760,N_2772,N_2986);
or U3761 (N_3761,N_2545,N_2842);
nand U3762 (N_3762,N_2244,N_2275);
and U3763 (N_3763,N_2394,N_2223);
nand U3764 (N_3764,N_2729,N_2274);
nor U3765 (N_3765,N_2470,N_2606);
nand U3766 (N_3766,N_2339,N_2445);
or U3767 (N_3767,N_2093,N_2817);
nand U3768 (N_3768,N_2288,N_2408);
xor U3769 (N_3769,N_2469,N_2031);
and U3770 (N_3770,N_2705,N_2016);
nor U3771 (N_3771,N_2706,N_2224);
nand U3772 (N_3772,N_2304,N_2317);
or U3773 (N_3773,N_2761,N_2582);
and U3774 (N_3774,N_2667,N_2064);
nor U3775 (N_3775,N_2000,N_2071);
nor U3776 (N_3776,N_2107,N_2892);
xor U3777 (N_3777,N_2160,N_2077);
nand U3778 (N_3778,N_2501,N_2677);
nand U3779 (N_3779,N_2131,N_2565);
and U3780 (N_3780,N_2871,N_2386);
or U3781 (N_3781,N_2225,N_2453);
and U3782 (N_3782,N_2177,N_2427);
and U3783 (N_3783,N_2949,N_2851);
nor U3784 (N_3784,N_2865,N_2206);
nor U3785 (N_3785,N_2393,N_2457);
nor U3786 (N_3786,N_2277,N_2513);
nand U3787 (N_3787,N_2744,N_2964);
nor U3788 (N_3788,N_2807,N_2502);
xnor U3789 (N_3789,N_2170,N_2063);
or U3790 (N_3790,N_2750,N_2216);
nand U3791 (N_3791,N_2557,N_2871);
nand U3792 (N_3792,N_2537,N_2449);
or U3793 (N_3793,N_2851,N_2989);
or U3794 (N_3794,N_2285,N_2806);
or U3795 (N_3795,N_2255,N_2386);
or U3796 (N_3796,N_2148,N_2583);
and U3797 (N_3797,N_2959,N_2576);
nor U3798 (N_3798,N_2488,N_2943);
or U3799 (N_3799,N_2828,N_2301);
nor U3800 (N_3800,N_2030,N_2508);
nor U3801 (N_3801,N_2916,N_2871);
and U3802 (N_3802,N_2701,N_2279);
nor U3803 (N_3803,N_2884,N_2957);
nor U3804 (N_3804,N_2862,N_2432);
and U3805 (N_3805,N_2102,N_2905);
xor U3806 (N_3806,N_2750,N_2343);
xnor U3807 (N_3807,N_2379,N_2065);
nand U3808 (N_3808,N_2431,N_2818);
or U3809 (N_3809,N_2144,N_2434);
or U3810 (N_3810,N_2659,N_2158);
xor U3811 (N_3811,N_2633,N_2199);
and U3812 (N_3812,N_2776,N_2303);
xnor U3813 (N_3813,N_2299,N_2225);
xor U3814 (N_3814,N_2270,N_2092);
nor U3815 (N_3815,N_2087,N_2074);
or U3816 (N_3816,N_2911,N_2569);
or U3817 (N_3817,N_2351,N_2924);
or U3818 (N_3818,N_2692,N_2384);
and U3819 (N_3819,N_2000,N_2646);
and U3820 (N_3820,N_2217,N_2059);
xor U3821 (N_3821,N_2151,N_2828);
and U3822 (N_3822,N_2829,N_2249);
or U3823 (N_3823,N_2528,N_2757);
or U3824 (N_3824,N_2342,N_2387);
nor U3825 (N_3825,N_2651,N_2729);
nand U3826 (N_3826,N_2070,N_2283);
xor U3827 (N_3827,N_2974,N_2119);
nor U3828 (N_3828,N_2795,N_2530);
xor U3829 (N_3829,N_2661,N_2985);
nor U3830 (N_3830,N_2514,N_2754);
or U3831 (N_3831,N_2242,N_2906);
and U3832 (N_3832,N_2185,N_2665);
xnor U3833 (N_3833,N_2389,N_2594);
nand U3834 (N_3834,N_2206,N_2257);
nand U3835 (N_3835,N_2309,N_2298);
nor U3836 (N_3836,N_2156,N_2457);
xnor U3837 (N_3837,N_2548,N_2038);
nor U3838 (N_3838,N_2832,N_2827);
nor U3839 (N_3839,N_2122,N_2675);
nand U3840 (N_3840,N_2622,N_2602);
nor U3841 (N_3841,N_2747,N_2241);
nor U3842 (N_3842,N_2526,N_2062);
nand U3843 (N_3843,N_2872,N_2814);
or U3844 (N_3844,N_2447,N_2888);
and U3845 (N_3845,N_2201,N_2024);
and U3846 (N_3846,N_2867,N_2426);
xor U3847 (N_3847,N_2532,N_2960);
xnor U3848 (N_3848,N_2493,N_2546);
and U3849 (N_3849,N_2099,N_2330);
nand U3850 (N_3850,N_2099,N_2635);
or U3851 (N_3851,N_2154,N_2457);
nand U3852 (N_3852,N_2137,N_2900);
nand U3853 (N_3853,N_2291,N_2292);
or U3854 (N_3854,N_2911,N_2724);
and U3855 (N_3855,N_2938,N_2231);
or U3856 (N_3856,N_2704,N_2209);
and U3857 (N_3857,N_2241,N_2598);
nor U3858 (N_3858,N_2353,N_2283);
or U3859 (N_3859,N_2851,N_2446);
nor U3860 (N_3860,N_2789,N_2858);
nor U3861 (N_3861,N_2323,N_2409);
nor U3862 (N_3862,N_2439,N_2856);
or U3863 (N_3863,N_2019,N_2955);
and U3864 (N_3864,N_2187,N_2153);
and U3865 (N_3865,N_2131,N_2476);
nand U3866 (N_3866,N_2419,N_2169);
or U3867 (N_3867,N_2184,N_2629);
or U3868 (N_3868,N_2733,N_2908);
nor U3869 (N_3869,N_2679,N_2429);
or U3870 (N_3870,N_2703,N_2083);
nand U3871 (N_3871,N_2197,N_2342);
or U3872 (N_3872,N_2405,N_2965);
or U3873 (N_3873,N_2830,N_2151);
and U3874 (N_3874,N_2087,N_2675);
nor U3875 (N_3875,N_2389,N_2127);
xor U3876 (N_3876,N_2067,N_2133);
or U3877 (N_3877,N_2774,N_2575);
nor U3878 (N_3878,N_2029,N_2727);
nor U3879 (N_3879,N_2787,N_2952);
or U3880 (N_3880,N_2290,N_2762);
nand U3881 (N_3881,N_2035,N_2993);
xor U3882 (N_3882,N_2984,N_2985);
or U3883 (N_3883,N_2801,N_2285);
nand U3884 (N_3884,N_2660,N_2591);
xnor U3885 (N_3885,N_2506,N_2173);
nand U3886 (N_3886,N_2659,N_2624);
and U3887 (N_3887,N_2865,N_2516);
xnor U3888 (N_3888,N_2653,N_2246);
xnor U3889 (N_3889,N_2252,N_2610);
nor U3890 (N_3890,N_2656,N_2435);
nor U3891 (N_3891,N_2956,N_2450);
nand U3892 (N_3892,N_2228,N_2082);
or U3893 (N_3893,N_2153,N_2129);
and U3894 (N_3894,N_2475,N_2544);
or U3895 (N_3895,N_2281,N_2596);
nand U3896 (N_3896,N_2169,N_2352);
nand U3897 (N_3897,N_2841,N_2024);
nand U3898 (N_3898,N_2477,N_2774);
nand U3899 (N_3899,N_2622,N_2051);
nor U3900 (N_3900,N_2617,N_2717);
xor U3901 (N_3901,N_2166,N_2396);
nand U3902 (N_3902,N_2350,N_2868);
or U3903 (N_3903,N_2982,N_2796);
xnor U3904 (N_3904,N_2038,N_2205);
and U3905 (N_3905,N_2645,N_2437);
xnor U3906 (N_3906,N_2337,N_2752);
xor U3907 (N_3907,N_2119,N_2310);
or U3908 (N_3908,N_2605,N_2810);
or U3909 (N_3909,N_2921,N_2671);
xnor U3910 (N_3910,N_2592,N_2394);
or U3911 (N_3911,N_2484,N_2234);
or U3912 (N_3912,N_2490,N_2949);
or U3913 (N_3913,N_2593,N_2057);
or U3914 (N_3914,N_2531,N_2702);
xor U3915 (N_3915,N_2090,N_2766);
nor U3916 (N_3916,N_2529,N_2982);
nand U3917 (N_3917,N_2798,N_2681);
and U3918 (N_3918,N_2486,N_2916);
xor U3919 (N_3919,N_2966,N_2433);
xnor U3920 (N_3920,N_2355,N_2844);
nor U3921 (N_3921,N_2314,N_2211);
nor U3922 (N_3922,N_2217,N_2736);
or U3923 (N_3923,N_2836,N_2973);
xnor U3924 (N_3924,N_2297,N_2101);
nor U3925 (N_3925,N_2704,N_2872);
nor U3926 (N_3926,N_2800,N_2965);
nand U3927 (N_3927,N_2046,N_2895);
nand U3928 (N_3928,N_2776,N_2523);
nand U3929 (N_3929,N_2991,N_2931);
xnor U3930 (N_3930,N_2419,N_2783);
xor U3931 (N_3931,N_2207,N_2853);
nor U3932 (N_3932,N_2991,N_2171);
and U3933 (N_3933,N_2658,N_2342);
xnor U3934 (N_3934,N_2406,N_2358);
xor U3935 (N_3935,N_2487,N_2766);
or U3936 (N_3936,N_2200,N_2575);
and U3937 (N_3937,N_2250,N_2673);
nand U3938 (N_3938,N_2193,N_2819);
nand U3939 (N_3939,N_2963,N_2888);
and U3940 (N_3940,N_2415,N_2640);
nand U3941 (N_3941,N_2177,N_2793);
or U3942 (N_3942,N_2336,N_2070);
xnor U3943 (N_3943,N_2520,N_2370);
or U3944 (N_3944,N_2888,N_2975);
nand U3945 (N_3945,N_2023,N_2910);
nand U3946 (N_3946,N_2505,N_2641);
and U3947 (N_3947,N_2082,N_2632);
and U3948 (N_3948,N_2083,N_2813);
or U3949 (N_3949,N_2391,N_2031);
xor U3950 (N_3950,N_2249,N_2581);
and U3951 (N_3951,N_2255,N_2316);
xor U3952 (N_3952,N_2987,N_2405);
and U3953 (N_3953,N_2218,N_2328);
or U3954 (N_3954,N_2597,N_2480);
nand U3955 (N_3955,N_2334,N_2227);
and U3956 (N_3956,N_2407,N_2226);
and U3957 (N_3957,N_2434,N_2364);
or U3958 (N_3958,N_2099,N_2413);
xor U3959 (N_3959,N_2746,N_2140);
xnor U3960 (N_3960,N_2253,N_2335);
or U3961 (N_3961,N_2021,N_2782);
xor U3962 (N_3962,N_2749,N_2781);
nand U3963 (N_3963,N_2020,N_2317);
or U3964 (N_3964,N_2940,N_2943);
or U3965 (N_3965,N_2604,N_2319);
or U3966 (N_3966,N_2572,N_2179);
nor U3967 (N_3967,N_2017,N_2324);
nand U3968 (N_3968,N_2471,N_2482);
or U3969 (N_3969,N_2347,N_2557);
nand U3970 (N_3970,N_2475,N_2323);
nand U3971 (N_3971,N_2245,N_2349);
xor U3972 (N_3972,N_2379,N_2282);
and U3973 (N_3973,N_2927,N_2484);
or U3974 (N_3974,N_2799,N_2369);
nand U3975 (N_3975,N_2079,N_2481);
nor U3976 (N_3976,N_2779,N_2537);
and U3977 (N_3977,N_2561,N_2714);
and U3978 (N_3978,N_2679,N_2309);
and U3979 (N_3979,N_2976,N_2550);
or U3980 (N_3980,N_2695,N_2901);
or U3981 (N_3981,N_2578,N_2890);
or U3982 (N_3982,N_2368,N_2025);
nor U3983 (N_3983,N_2403,N_2124);
xor U3984 (N_3984,N_2427,N_2284);
or U3985 (N_3985,N_2585,N_2128);
and U3986 (N_3986,N_2197,N_2117);
xor U3987 (N_3987,N_2884,N_2234);
and U3988 (N_3988,N_2759,N_2505);
or U3989 (N_3989,N_2255,N_2329);
xor U3990 (N_3990,N_2749,N_2954);
or U3991 (N_3991,N_2894,N_2802);
and U3992 (N_3992,N_2949,N_2603);
nand U3993 (N_3993,N_2777,N_2883);
nor U3994 (N_3994,N_2640,N_2101);
nor U3995 (N_3995,N_2274,N_2163);
and U3996 (N_3996,N_2830,N_2384);
xnor U3997 (N_3997,N_2491,N_2982);
nor U3998 (N_3998,N_2233,N_2045);
nand U3999 (N_3999,N_2921,N_2684);
nor U4000 (N_4000,N_3573,N_3727);
nand U4001 (N_4001,N_3480,N_3147);
and U4002 (N_4002,N_3347,N_3964);
xnor U4003 (N_4003,N_3708,N_3926);
nor U4004 (N_4004,N_3261,N_3114);
and U4005 (N_4005,N_3850,N_3288);
nor U4006 (N_4006,N_3344,N_3748);
nand U4007 (N_4007,N_3403,N_3284);
nand U4008 (N_4008,N_3343,N_3503);
or U4009 (N_4009,N_3691,N_3022);
and U4010 (N_4010,N_3671,N_3747);
nor U4011 (N_4011,N_3552,N_3351);
nand U4012 (N_4012,N_3101,N_3064);
xor U4013 (N_4013,N_3120,N_3137);
or U4014 (N_4014,N_3061,N_3297);
nor U4015 (N_4015,N_3650,N_3085);
or U4016 (N_4016,N_3198,N_3566);
and U4017 (N_4017,N_3400,N_3913);
nor U4018 (N_4018,N_3544,N_3067);
or U4019 (N_4019,N_3981,N_3482);
or U4020 (N_4020,N_3464,N_3791);
xor U4021 (N_4021,N_3001,N_3592);
or U4022 (N_4022,N_3232,N_3595);
xor U4023 (N_4023,N_3349,N_3947);
nor U4024 (N_4024,N_3522,N_3455);
xor U4025 (N_4025,N_3607,N_3336);
nor U4026 (N_4026,N_3366,N_3923);
nor U4027 (N_4027,N_3654,N_3514);
nand U4028 (N_4028,N_3800,N_3183);
and U4029 (N_4029,N_3688,N_3760);
nor U4030 (N_4030,N_3167,N_3775);
nand U4031 (N_4031,N_3585,N_3192);
and U4032 (N_4032,N_3833,N_3849);
xnor U4033 (N_4033,N_3524,N_3195);
and U4034 (N_4034,N_3541,N_3104);
nand U4035 (N_4035,N_3009,N_3633);
and U4036 (N_4036,N_3015,N_3393);
and U4037 (N_4037,N_3058,N_3793);
nand U4038 (N_4038,N_3672,N_3720);
or U4039 (N_4039,N_3334,N_3606);
nand U4040 (N_4040,N_3243,N_3837);
and U4041 (N_4041,N_3971,N_3270);
or U4042 (N_4042,N_3094,N_3008);
xnor U4043 (N_4043,N_3123,N_3630);
and U4044 (N_4044,N_3483,N_3076);
or U4045 (N_4045,N_3941,N_3286);
nand U4046 (N_4046,N_3012,N_3276);
nor U4047 (N_4047,N_3726,N_3025);
nand U4048 (N_4048,N_3485,N_3581);
xor U4049 (N_4049,N_3516,N_3081);
xor U4050 (N_4050,N_3899,N_3239);
nor U4051 (N_4051,N_3486,N_3365);
xnor U4052 (N_4052,N_3471,N_3865);
and U4053 (N_4053,N_3829,N_3171);
or U4054 (N_4054,N_3624,N_3704);
nand U4055 (N_4055,N_3262,N_3035);
nand U4056 (N_4056,N_3901,N_3756);
nand U4057 (N_4057,N_3282,N_3465);
or U4058 (N_4058,N_3152,N_3869);
and U4059 (N_4059,N_3433,N_3037);
xor U4060 (N_4060,N_3616,N_3158);
xnor U4061 (N_4061,N_3130,N_3538);
or U4062 (N_4062,N_3567,N_3718);
or U4063 (N_4063,N_3359,N_3223);
nand U4064 (N_4064,N_3303,N_3583);
or U4065 (N_4065,N_3325,N_3976);
and U4066 (N_4066,N_3499,N_3445);
or U4067 (N_4067,N_3294,N_3354);
and U4068 (N_4068,N_3319,N_3342);
and U4069 (N_4069,N_3231,N_3597);
nand U4070 (N_4070,N_3109,N_3017);
xor U4071 (N_4071,N_3222,N_3838);
nor U4072 (N_4072,N_3315,N_3690);
and U4073 (N_4073,N_3089,N_3611);
nor U4074 (N_4074,N_3204,N_3646);
and U4075 (N_4075,N_3280,N_3373);
xnor U4076 (N_4076,N_3874,N_3535);
or U4077 (N_4077,N_3221,N_3982);
nand U4078 (N_4078,N_3780,N_3448);
and U4079 (N_4079,N_3519,N_3052);
nand U4080 (N_4080,N_3186,N_3033);
and U4081 (N_4081,N_3752,N_3735);
nor U4082 (N_4082,N_3555,N_3125);
xnor U4083 (N_4083,N_3554,N_3233);
or U4084 (N_4084,N_3041,N_3134);
nor U4085 (N_4085,N_3447,N_3574);
xor U4086 (N_4086,N_3117,N_3989);
and U4087 (N_4087,N_3924,N_3778);
and U4088 (N_4088,N_3978,N_3897);
and U4089 (N_4089,N_3238,N_3316);
and U4090 (N_4090,N_3677,N_3371);
or U4091 (N_4091,N_3864,N_3938);
xor U4092 (N_4092,N_3478,N_3802);
or U4093 (N_4093,N_3467,N_3749);
or U4094 (N_4094,N_3593,N_3868);
nor U4095 (N_4095,N_3281,N_3449);
and U4096 (N_4096,N_3235,N_3405);
nand U4097 (N_4097,N_3438,N_3504);
or U4098 (N_4098,N_3220,N_3859);
and U4099 (N_4099,N_3717,N_3951);
or U4100 (N_4100,N_3248,N_3863);
or U4101 (N_4101,N_3434,N_3569);
or U4102 (N_4102,N_3757,N_3796);
nand U4103 (N_4103,N_3830,N_3200);
nor U4104 (N_4104,N_3072,N_3598);
nand U4105 (N_4105,N_3429,N_3783);
nand U4106 (N_4106,N_3182,N_3181);
nand U4107 (N_4107,N_3754,N_3875);
and U4108 (N_4108,N_3350,N_3475);
and U4109 (N_4109,N_3087,N_3695);
nand U4110 (N_4110,N_3962,N_3259);
and U4111 (N_4111,N_3827,N_3384);
or U4112 (N_4112,N_3651,N_3391);
xnor U4113 (N_4113,N_3051,N_3534);
or U4114 (N_4114,N_3702,N_3550);
xor U4115 (N_4115,N_3229,N_3338);
nor U4116 (N_4116,N_3804,N_3715);
nand U4117 (N_4117,N_3902,N_3249);
nor U4118 (N_4118,N_3030,N_3410);
or U4119 (N_4119,N_3662,N_3188);
xor U4120 (N_4120,N_3579,N_3339);
and U4121 (N_4121,N_3782,N_3692);
xnor U4122 (N_4122,N_3386,N_3431);
and U4123 (N_4123,N_3330,N_3210);
xor U4124 (N_4124,N_3424,N_3494);
xnor U4125 (N_4125,N_3224,N_3664);
xor U4126 (N_4126,N_3096,N_3716);
nand U4127 (N_4127,N_3712,N_3241);
nor U4128 (N_4128,N_3785,N_3044);
and U4129 (N_4129,N_3591,N_3111);
nor U4130 (N_4130,N_3866,N_3568);
or U4131 (N_4131,N_3641,N_3149);
and U4132 (N_4132,N_3142,N_3847);
nand U4133 (N_4133,N_3961,N_3640);
nor U4134 (N_4134,N_3685,N_3675);
nand U4135 (N_4135,N_3059,N_3387);
nand U4136 (N_4136,N_3832,N_3549);
and U4137 (N_4137,N_3011,N_3290);
nor U4138 (N_4138,N_3614,N_3762);
or U4139 (N_4139,N_3027,N_3751);
or U4140 (N_4140,N_3329,N_3605);
nand U4141 (N_4141,N_3040,N_3098);
or U4142 (N_4142,N_3036,N_3031);
nand U4143 (N_4143,N_3217,N_3079);
nor U4144 (N_4144,N_3257,N_3407);
nand U4145 (N_4145,N_3417,N_3604);
nand U4146 (N_4146,N_3620,N_3670);
and U4147 (N_4147,N_3644,N_3584);
xnor U4148 (N_4148,N_3856,N_3308);
or U4149 (N_4149,N_3808,N_3187);
or U4150 (N_4150,N_3103,N_3054);
nand U4151 (N_4151,N_3537,N_3794);
nand U4152 (N_4152,N_3296,N_3132);
xnor U4153 (N_4153,N_3673,N_3457);
nor U4154 (N_4154,N_3996,N_3706);
and U4155 (N_4155,N_3985,N_3444);
nor U4156 (N_4156,N_3805,N_3102);
or U4157 (N_4157,N_3967,N_3007);
or U4158 (N_4158,N_3321,N_3881);
nand U4159 (N_4159,N_3416,N_3841);
nand U4160 (N_4160,N_3769,N_3994);
or U4161 (N_4161,N_3974,N_3307);
xor U4162 (N_4162,N_3713,N_3674);
nand U4163 (N_4163,N_3189,N_3678);
and U4164 (N_4164,N_3264,N_3157);
and U4165 (N_4165,N_3473,N_3698);
and U4166 (N_4166,N_3118,N_3043);
nor U4167 (N_4167,N_3355,N_3122);
or U4168 (N_4168,N_3199,N_3969);
nand U4169 (N_4169,N_3739,N_3732);
nor U4170 (N_4170,N_3172,N_3470);
and U4171 (N_4171,N_3430,N_3601);
and U4172 (N_4172,N_3090,N_3379);
nor U4173 (N_4173,N_3218,N_3441);
nand U4174 (N_4174,N_3068,N_3385);
nand U4175 (N_4175,N_3244,N_3669);
or U4176 (N_4176,N_3358,N_3986);
nand U4177 (N_4177,N_3487,N_3993);
and U4178 (N_4178,N_3759,N_3860);
nor U4179 (N_4179,N_3828,N_3943);
and U4180 (N_4180,N_3415,N_3053);
xor U4181 (N_4181,N_3046,N_3772);
or U4182 (N_4182,N_3163,N_3177);
nand U4183 (N_4183,N_3495,N_3460);
or U4184 (N_4184,N_3419,N_3806);
nor U4185 (N_4185,N_3689,N_3298);
and U4186 (N_4186,N_3705,N_3942);
and U4187 (N_4187,N_3959,N_3477);
xnor U4188 (N_4188,N_3013,N_3446);
nor U4189 (N_4189,N_3932,N_3839);
nor U4190 (N_4190,N_3144,N_3882);
or U4191 (N_4191,N_3742,N_3723);
and U4192 (N_4192,N_3397,N_3944);
nor U4193 (N_4193,N_3505,N_3439);
nand U4194 (N_4194,N_3469,N_3703);
xor U4195 (N_4195,N_3092,N_3107);
nor U4196 (N_4196,N_3211,N_3411);
xor U4197 (N_4197,N_3071,N_3602);
or U4198 (N_4198,N_3452,N_3062);
and U4199 (N_4199,N_3139,N_3202);
or U4200 (N_4200,N_3907,N_3528);
and U4201 (N_4201,N_3443,N_3631);
nand U4202 (N_4202,N_3219,N_3572);
xnor U4203 (N_4203,N_3375,N_3225);
nand U4204 (N_4204,N_3639,N_3159);
xor U4205 (N_4205,N_3625,N_3075);
and U4206 (N_4206,N_3617,N_3966);
xnor U4207 (N_4207,N_3888,N_3658);
nand U4208 (N_4208,N_3842,N_3911);
nand U4209 (N_4209,N_3065,N_3401);
or U4210 (N_4210,N_3813,N_3694);
nand U4211 (N_4211,N_3077,N_3594);
nor U4212 (N_4212,N_3547,N_3771);
nor U4213 (N_4213,N_3816,N_3861);
xor U4214 (N_4214,N_3110,N_3176);
nor U4215 (N_4215,N_3809,N_3684);
or U4216 (N_4216,N_3073,N_3164);
and U4217 (N_4217,N_3180,N_3468);
xnor U4218 (N_4218,N_3738,N_3790);
or U4219 (N_4219,N_3984,N_3545);
or U4220 (N_4220,N_3655,N_3255);
nor U4221 (N_4221,N_3958,N_3807);
or U4222 (N_4222,N_3636,N_3922);
and U4223 (N_4223,N_3965,N_3454);
nor U4224 (N_4224,N_3332,N_3234);
xor U4225 (N_4225,N_3878,N_3484);
or U4226 (N_4226,N_3895,N_3948);
xnor U4227 (N_4227,N_3879,N_3408);
and U4228 (N_4228,N_3214,N_3877);
nand U4229 (N_4229,N_3283,N_3275);
xnor U4230 (N_4230,N_3331,N_3663);
nor U4231 (N_4231,N_3596,N_3287);
and U4232 (N_4232,N_3770,N_3175);
nor U4233 (N_4233,N_3954,N_3437);
nor U4234 (N_4234,N_3333,N_3803);
and U4235 (N_4235,N_3588,N_3997);
nand U4236 (N_4236,N_3462,N_3766);
nor U4237 (N_4237,N_3208,N_3786);
nor U4238 (N_4238,N_3896,N_3776);
xnor U4239 (N_4239,N_3666,N_3404);
xnor U4240 (N_4240,N_3173,N_3014);
nand U4241 (N_4241,N_3661,N_3196);
nor U4242 (N_4242,N_3817,N_3721);
nand U4243 (N_4243,N_3378,N_3129);
nand U4244 (N_4244,N_3362,N_3843);
nand U4245 (N_4245,N_3546,N_3736);
xor U4246 (N_4246,N_3936,N_3292);
and U4247 (N_4247,N_3696,N_3836);
or U4248 (N_4248,N_3066,N_3042);
or U4249 (N_4249,N_3931,N_3493);
and U4250 (N_4250,N_3975,N_3131);
nor U4251 (N_4251,N_3459,N_3299);
xnor U4252 (N_4252,N_3872,N_3920);
xnor U4253 (N_4253,N_3435,N_3532);
nor U4254 (N_4254,N_3768,N_3600);
nand U4255 (N_4255,N_3069,N_3876);
and U4256 (N_4256,N_3983,N_3300);
xnor U4257 (N_4257,N_3151,N_3517);
xor U4258 (N_4258,N_3921,N_3615);
or U4259 (N_4259,N_3491,N_3548);
xor U4260 (N_4260,N_3680,N_3972);
nand U4261 (N_4261,N_3097,N_3100);
xor U4262 (N_4262,N_3165,N_3973);
or U4263 (N_4263,N_3587,N_3267);
and U4264 (N_4264,N_3070,N_3178);
and U4265 (N_4265,N_3203,N_3621);
nor U4266 (N_4266,N_3019,N_3140);
nor U4267 (N_4267,N_3979,N_3657);
xnor U4268 (N_4268,N_3571,N_3511);
nand U4269 (N_4269,N_3010,N_3610);
nand U4270 (N_4270,N_3256,N_3057);
nand U4271 (N_4271,N_3258,N_3145);
xnor U4272 (N_4272,N_3635,N_3016);
or U4273 (N_4273,N_3949,N_3476);
and U4274 (N_4274,N_3834,N_3360);
nor U4275 (N_4275,N_3274,N_3905);
nand U4276 (N_4276,N_3518,N_3753);
nor U4277 (N_4277,N_3285,N_3987);
or U4278 (N_4278,N_3953,N_3002);
nand U4279 (N_4279,N_3466,N_3278);
or U4280 (N_4280,N_3853,N_3789);
nand U4281 (N_4281,N_3337,N_3939);
nor U4282 (N_4282,N_3481,N_3247);
or U4283 (N_4283,N_3521,N_3508);
or U4284 (N_4284,N_3492,N_3724);
or U4285 (N_4285,N_3626,N_3489);
and U4286 (N_4286,N_3370,N_3091);
xor U4287 (N_4287,N_3113,N_3867);
xnor U4288 (N_4288,N_3216,N_3909);
or U4289 (N_4289,N_3099,N_3647);
or U4290 (N_4290,N_3324,N_3764);
or U4291 (N_4291,N_3741,N_3798);
or U4292 (N_4292,N_3341,N_3472);
and U4293 (N_4293,N_3078,N_3908);
xnor U4294 (N_4294,N_3266,N_3925);
nor U4295 (N_4295,N_3507,N_3686);
nor U4296 (N_4296,N_3840,N_3364);
and U4297 (N_4297,N_3810,N_3029);
xor U4298 (N_4298,N_3496,N_3613);
xor U4299 (N_4299,N_3682,N_3020);
nor U4300 (N_4300,N_3004,N_3348);
xnor U4301 (N_4301,N_3245,N_3612);
xnor U4302 (N_4302,N_3719,N_3918);
xor U4303 (N_4303,N_3711,N_3930);
and U4304 (N_4304,N_3021,N_3995);
nor U4305 (N_4305,N_3525,N_3729);
nand U4306 (N_4306,N_3999,N_3381);
and U4307 (N_4307,N_3442,N_3426);
or U4308 (N_4308,N_3826,N_3609);
or U4309 (N_4309,N_3858,N_3461);
nor U4310 (N_4310,N_3160,N_3819);
or U4311 (N_4311,N_3784,N_3127);
and U4312 (N_4312,N_3056,N_3302);
nor U4313 (N_4313,N_3880,N_3251);
or U4314 (N_4314,N_3761,N_3005);
or U4315 (N_4315,N_3374,N_3561);
and U4316 (N_4316,N_3787,N_3055);
nand U4317 (N_4317,N_3520,N_3265);
xnor U4318 (N_4318,N_3990,N_3095);
or U4319 (N_4319,N_3291,N_3855);
nor U4320 (N_4320,N_3904,N_3138);
nand U4321 (N_4321,N_3335,N_3559);
xor U4322 (N_4322,N_3318,N_3952);
nand U4323 (N_4323,N_3889,N_3083);
nor U4324 (N_4324,N_3980,N_3844);
or U4325 (N_4325,N_3575,N_3553);
or U4326 (N_4326,N_3295,N_3795);
or U4327 (N_4327,N_3937,N_3676);
nor U4328 (N_4328,N_3821,N_3490);
xor U4329 (N_4329,N_3523,N_3873);
and U4330 (N_4330,N_3313,N_3389);
nand U4331 (N_4331,N_3608,N_3565);
or U4332 (N_4332,N_3629,N_3818);
nand U4333 (N_4333,N_3088,N_3557);
xnor U4334 (N_4334,N_3825,N_3136);
and U4335 (N_4335,N_3246,N_3279);
and U4336 (N_4336,N_3734,N_3352);
or U4337 (N_4337,N_3835,N_3121);
nand U4338 (N_4338,N_3506,N_3309);
or U4339 (N_4339,N_3126,N_3693);
nor U4340 (N_4340,N_3701,N_3133);
and U4341 (N_4341,N_3003,N_3831);
nor U4342 (N_4342,N_3150,N_3311);
and U4343 (N_4343,N_3420,N_3394);
nor U4344 (N_4344,N_3193,N_3846);
nand U4345 (N_4345,N_3060,N_3363);
xnor U4346 (N_4346,N_3322,N_3038);
and U4347 (N_4347,N_3562,N_3082);
nand U4348 (N_4348,N_3627,N_3201);
nand U4349 (N_4349,N_3515,N_3935);
or U4350 (N_4350,N_3722,N_3240);
xnor U4351 (N_4351,N_3968,N_3892);
xor U4352 (N_4352,N_3166,N_3432);
nor U4353 (N_4353,N_3665,N_3327);
xor U4354 (N_4354,N_3209,N_3268);
nand U4355 (N_4355,N_3032,N_3618);
nand U4356 (N_4356,N_3632,N_3540);
or U4357 (N_4357,N_3148,N_3578);
xor U4358 (N_4358,N_3206,N_3250);
and U4359 (N_4359,N_3084,N_3227);
and U4360 (N_4360,N_3305,N_3928);
nor U4361 (N_4361,N_3028,N_3707);
nor U4362 (N_4362,N_3765,N_3049);
or U4363 (N_4363,N_3425,N_3854);
and U4364 (N_4364,N_3950,N_3306);
xor U4365 (N_4365,N_3513,N_3603);
nand U4366 (N_4366,N_3412,N_3498);
xnor U4367 (N_4367,N_3891,N_3380);
xor U4368 (N_4368,N_3301,N_3992);
and U4369 (N_4369,N_3745,N_3851);
xor U4370 (N_4370,N_3115,N_3326);
nor U4371 (N_4371,N_3773,N_3758);
and U4372 (N_4372,N_3230,N_3599);
nand U4373 (N_4373,N_3893,N_3169);
nand U4374 (N_4374,N_3755,N_3212);
or U4375 (N_4375,N_3155,N_3822);
or U4376 (N_4376,N_3509,N_3414);
and U4377 (N_4377,N_3699,N_3582);
nand U4378 (N_4378,N_3733,N_3638);
and U4379 (N_4379,N_3543,N_3048);
nor U4380 (N_4380,N_3047,N_3197);
xor U4381 (N_4381,N_3497,N_3356);
xnor U4382 (N_4382,N_3643,N_3558);
and U4383 (N_4383,N_3887,N_3940);
xnor U4384 (N_4384,N_3919,N_3914);
nor U4385 (N_4385,N_3746,N_3645);
nor U4386 (N_4386,N_3141,N_3927);
nor U4387 (N_4387,N_3273,N_3915);
nor U4388 (N_4388,N_3080,N_3501);
or U4389 (N_4389,N_3293,N_3185);
and U4390 (N_4390,N_3906,N_3656);
or U4391 (N_4391,N_3890,N_3576);
xnor U4392 (N_4392,N_3886,N_3812);
and U4393 (N_4393,N_3026,N_3709);
nor U4394 (N_4394,N_3564,N_3777);
nand U4395 (N_4395,N_3289,N_3551);
nor U4396 (N_4396,N_3310,N_3112);
nand U4397 (N_4397,N_3395,N_3668);
nor U4398 (N_4398,N_3642,N_3399);
nand U4399 (N_4399,N_3063,N_3667);
or U4400 (N_4400,N_3074,N_3988);
nor U4401 (N_4401,N_3254,N_3413);
and U4402 (N_4402,N_3884,N_3590);
and U4403 (N_4403,N_3418,N_3086);
nand U4404 (N_4404,N_3916,N_3767);
xor U4405 (N_4405,N_3153,N_3710);
nand U4406 (N_4406,N_3398,N_3116);
or U4407 (N_4407,N_3406,N_3955);
xnor U4408 (N_4408,N_3731,N_3502);
nand U4409 (N_4409,N_3162,N_3191);
and U4410 (N_4410,N_3228,N_3253);
or U4411 (N_4411,N_3168,N_3367);
xor U4412 (N_4412,N_3570,N_3623);
xor U4413 (N_4413,N_3361,N_3006);
xor U4414 (N_4414,N_3527,N_3402);
and U4415 (N_4415,N_3883,N_3392);
nand U4416 (N_4416,N_3945,N_3563);
or U4417 (N_4417,N_3589,N_3423);
xnor U4418 (N_4418,N_3119,N_3346);
xor U4419 (N_4419,N_3143,N_3124);
nand U4420 (N_4420,N_3660,N_3900);
or U4421 (N_4421,N_3215,N_3637);
xor U4422 (N_4422,N_3422,N_3500);
nor U4423 (N_4423,N_3312,N_3269);
nor U4424 (N_4424,N_3372,N_3530);
xor U4425 (N_4425,N_3377,N_3533);
and U4426 (N_4426,N_3237,N_3531);
nand U4427 (N_4427,N_3252,N_3845);
or U4428 (N_4428,N_3050,N_3910);
or U4429 (N_4429,N_3421,N_3536);
and U4430 (N_4430,N_3488,N_3529);
nor U4431 (N_4431,N_3763,N_3912);
nor U4432 (N_4432,N_3453,N_3263);
nor U4433 (N_4433,N_3871,N_3045);
and U4434 (N_4434,N_3862,N_3190);
xnor U4435 (N_4435,N_3236,N_3560);
or U4436 (N_4436,N_3382,N_3368);
nor U4437 (N_4437,N_3396,N_3146);
nor U4438 (N_4438,N_3474,N_3797);
and U4439 (N_4439,N_3106,N_3323);
xor U4440 (N_4440,N_3648,N_3857);
nand U4441 (N_4441,N_3376,N_3799);
and U4442 (N_4442,N_3357,N_3328);
nor U4443 (N_4443,N_3314,N_3304);
xnor U4444 (N_4444,N_3619,N_3934);
nand U4445 (N_4445,N_3135,N_3659);
xor U4446 (N_4446,N_3622,N_3801);
or U4447 (N_4447,N_3450,N_3929);
nor U4448 (N_4448,N_3815,N_3510);
and U4449 (N_4449,N_3226,N_3207);
nand U4450 (N_4450,N_3779,N_3458);
xor U4451 (N_4451,N_3023,N_3652);
nor U4452 (N_4452,N_3156,N_3811);
nor U4453 (N_4453,N_3714,N_3440);
nor U4454 (N_4454,N_3260,N_3039);
and U4455 (N_4455,N_3687,N_3653);
xnor U4456 (N_4456,N_3024,N_3586);
nand U4457 (N_4457,N_3272,N_3018);
and U4458 (N_4458,N_3681,N_3409);
nand U4459 (N_4459,N_3577,N_3194);
and U4460 (N_4460,N_3957,N_3898);
or U4461 (N_4461,N_3427,N_3728);
or U4462 (N_4462,N_3730,N_3539);
xnor U4463 (N_4463,N_3823,N_3774);
nand U4464 (N_4464,N_3700,N_3242);
and U4465 (N_4465,N_3317,N_3743);
or U4466 (N_4466,N_3034,N_3456);
or U4467 (N_4467,N_3277,N_3824);
or U4468 (N_4468,N_3184,N_3428);
nand U4469 (N_4469,N_3814,N_3960);
xnor U4470 (N_4470,N_3956,N_3820);
or U4471 (N_4471,N_3963,N_3345);
and U4472 (N_4472,N_3991,N_3161);
xnor U4473 (N_4473,N_3970,N_3383);
nand U4474 (N_4474,N_3885,N_3894);
or U4475 (N_4475,N_3000,N_3744);
nand U4476 (N_4476,N_3998,N_3105);
nor U4477 (N_4477,N_3463,N_3128);
nor U4478 (N_4478,N_3390,N_3781);
and U4479 (N_4479,N_3679,N_3792);
nand U4480 (N_4480,N_3512,N_3271);
nand U4481 (N_4481,N_3634,N_3946);
nand U4482 (N_4482,N_3388,N_3542);
nor U4483 (N_4483,N_3628,N_3369);
xor U4484 (N_4484,N_3737,N_3649);
nor U4485 (N_4485,N_3340,N_3108);
nor U4486 (N_4486,N_3205,N_3320);
and U4487 (N_4487,N_3977,N_3093);
nand U4488 (N_4488,N_3697,N_3154);
nand U4489 (N_4489,N_3451,N_3870);
or U4490 (N_4490,N_3848,N_3170);
and U4491 (N_4491,N_3740,N_3580);
nor U4492 (N_4492,N_3526,N_3750);
nand U4493 (N_4493,N_3788,N_3917);
or U4494 (N_4494,N_3725,N_3436);
nor U4495 (N_4495,N_3174,N_3179);
nand U4496 (N_4496,N_3479,N_3933);
or U4497 (N_4497,N_3353,N_3556);
or U4498 (N_4498,N_3852,N_3683);
and U4499 (N_4499,N_3213,N_3903);
nand U4500 (N_4500,N_3816,N_3392);
nand U4501 (N_4501,N_3988,N_3246);
nor U4502 (N_4502,N_3510,N_3415);
nor U4503 (N_4503,N_3289,N_3409);
nand U4504 (N_4504,N_3116,N_3993);
nor U4505 (N_4505,N_3495,N_3853);
or U4506 (N_4506,N_3834,N_3296);
nand U4507 (N_4507,N_3696,N_3073);
or U4508 (N_4508,N_3432,N_3479);
xnor U4509 (N_4509,N_3446,N_3272);
and U4510 (N_4510,N_3812,N_3393);
nor U4511 (N_4511,N_3840,N_3975);
or U4512 (N_4512,N_3098,N_3626);
nor U4513 (N_4513,N_3326,N_3186);
nand U4514 (N_4514,N_3454,N_3260);
nor U4515 (N_4515,N_3618,N_3303);
nand U4516 (N_4516,N_3046,N_3283);
and U4517 (N_4517,N_3839,N_3824);
nor U4518 (N_4518,N_3558,N_3958);
xnor U4519 (N_4519,N_3500,N_3921);
and U4520 (N_4520,N_3029,N_3694);
and U4521 (N_4521,N_3231,N_3721);
nand U4522 (N_4522,N_3448,N_3096);
xnor U4523 (N_4523,N_3630,N_3733);
and U4524 (N_4524,N_3028,N_3462);
nor U4525 (N_4525,N_3454,N_3024);
and U4526 (N_4526,N_3052,N_3687);
nor U4527 (N_4527,N_3148,N_3368);
or U4528 (N_4528,N_3507,N_3326);
or U4529 (N_4529,N_3197,N_3780);
nor U4530 (N_4530,N_3784,N_3839);
xnor U4531 (N_4531,N_3457,N_3006);
nor U4532 (N_4532,N_3647,N_3824);
xor U4533 (N_4533,N_3036,N_3953);
or U4534 (N_4534,N_3679,N_3385);
nand U4535 (N_4535,N_3522,N_3341);
xnor U4536 (N_4536,N_3596,N_3182);
nand U4537 (N_4537,N_3207,N_3761);
nor U4538 (N_4538,N_3662,N_3132);
xor U4539 (N_4539,N_3686,N_3433);
and U4540 (N_4540,N_3667,N_3246);
xor U4541 (N_4541,N_3695,N_3047);
and U4542 (N_4542,N_3408,N_3901);
xnor U4543 (N_4543,N_3824,N_3642);
nor U4544 (N_4544,N_3472,N_3482);
nor U4545 (N_4545,N_3230,N_3037);
nand U4546 (N_4546,N_3146,N_3230);
or U4547 (N_4547,N_3850,N_3600);
and U4548 (N_4548,N_3969,N_3046);
xnor U4549 (N_4549,N_3644,N_3666);
xnor U4550 (N_4550,N_3011,N_3878);
nand U4551 (N_4551,N_3088,N_3436);
or U4552 (N_4552,N_3201,N_3083);
nor U4553 (N_4553,N_3013,N_3880);
nor U4554 (N_4554,N_3537,N_3886);
nor U4555 (N_4555,N_3725,N_3598);
nand U4556 (N_4556,N_3171,N_3922);
or U4557 (N_4557,N_3130,N_3838);
xor U4558 (N_4558,N_3550,N_3292);
and U4559 (N_4559,N_3338,N_3608);
xor U4560 (N_4560,N_3262,N_3242);
nor U4561 (N_4561,N_3339,N_3374);
xor U4562 (N_4562,N_3421,N_3591);
xnor U4563 (N_4563,N_3806,N_3008);
xnor U4564 (N_4564,N_3022,N_3731);
and U4565 (N_4565,N_3359,N_3409);
xnor U4566 (N_4566,N_3271,N_3022);
xor U4567 (N_4567,N_3078,N_3192);
and U4568 (N_4568,N_3828,N_3586);
nor U4569 (N_4569,N_3715,N_3473);
and U4570 (N_4570,N_3985,N_3365);
nand U4571 (N_4571,N_3019,N_3825);
or U4572 (N_4572,N_3196,N_3517);
nor U4573 (N_4573,N_3754,N_3467);
nand U4574 (N_4574,N_3346,N_3103);
or U4575 (N_4575,N_3956,N_3109);
or U4576 (N_4576,N_3056,N_3994);
and U4577 (N_4577,N_3732,N_3615);
xnor U4578 (N_4578,N_3250,N_3968);
nand U4579 (N_4579,N_3718,N_3345);
or U4580 (N_4580,N_3106,N_3899);
and U4581 (N_4581,N_3810,N_3785);
nor U4582 (N_4582,N_3922,N_3579);
or U4583 (N_4583,N_3163,N_3741);
xor U4584 (N_4584,N_3392,N_3489);
xnor U4585 (N_4585,N_3744,N_3813);
xnor U4586 (N_4586,N_3949,N_3140);
xor U4587 (N_4587,N_3393,N_3670);
nor U4588 (N_4588,N_3471,N_3413);
and U4589 (N_4589,N_3162,N_3940);
nor U4590 (N_4590,N_3084,N_3776);
nor U4591 (N_4591,N_3300,N_3601);
xnor U4592 (N_4592,N_3765,N_3526);
nor U4593 (N_4593,N_3396,N_3881);
xnor U4594 (N_4594,N_3057,N_3250);
and U4595 (N_4595,N_3570,N_3215);
and U4596 (N_4596,N_3331,N_3077);
and U4597 (N_4597,N_3822,N_3464);
nand U4598 (N_4598,N_3349,N_3652);
nand U4599 (N_4599,N_3035,N_3239);
nor U4600 (N_4600,N_3201,N_3174);
or U4601 (N_4601,N_3716,N_3784);
and U4602 (N_4602,N_3238,N_3507);
or U4603 (N_4603,N_3037,N_3503);
xnor U4604 (N_4604,N_3109,N_3339);
xnor U4605 (N_4605,N_3999,N_3823);
or U4606 (N_4606,N_3933,N_3216);
xor U4607 (N_4607,N_3359,N_3917);
or U4608 (N_4608,N_3822,N_3962);
or U4609 (N_4609,N_3753,N_3052);
xnor U4610 (N_4610,N_3462,N_3191);
nor U4611 (N_4611,N_3767,N_3726);
nor U4612 (N_4612,N_3222,N_3398);
xor U4613 (N_4613,N_3437,N_3555);
nor U4614 (N_4614,N_3712,N_3156);
and U4615 (N_4615,N_3310,N_3435);
nor U4616 (N_4616,N_3487,N_3356);
or U4617 (N_4617,N_3420,N_3005);
nor U4618 (N_4618,N_3696,N_3798);
nor U4619 (N_4619,N_3647,N_3905);
nor U4620 (N_4620,N_3090,N_3151);
and U4621 (N_4621,N_3757,N_3690);
and U4622 (N_4622,N_3963,N_3179);
or U4623 (N_4623,N_3856,N_3457);
nor U4624 (N_4624,N_3704,N_3429);
xor U4625 (N_4625,N_3843,N_3589);
nand U4626 (N_4626,N_3941,N_3658);
nand U4627 (N_4627,N_3000,N_3595);
and U4628 (N_4628,N_3122,N_3091);
xor U4629 (N_4629,N_3926,N_3551);
or U4630 (N_4630,N_3141,N_3826);
and U4631 (N_4631,N_3273,N_3737);
and U4632 (N_4632,N_3767,N_3276);
or U4633 (N_4633,N_3899,N_3331);
xor U4634 (N_4634,N_3563,N_3663);
nor U4635 (N_4635,N_3149,N_3873);
xor U4636 (N_4636,N_3770,N_3256);
xnor U4637 (N_4637,N_3321,N_3351);
xnor U4638 (N_4638,N_3814,N_3532);
and U4639 (N_4639,N_3901,N_3611);
nand U4640 (N_4640,N_3319,N_3847);
nand U4641 (N_4641,N_3523,N_3823);
nand U4642 (N_4642,N_3905,N_3058);
or U4643 (N_4643,N_3789,N_3486);
or U4644 (N_4644,N_3876,N_3262);
nor U4645 (N_4645,N_3849,N_3105);
nand U4646 (N_4646,N_3215,N_3074);
nor U4647 (N_4647,N_3618,N_3346);
nand U4648 (N_4648,N_3639,N_3340);
xnor U4649 (N_4649,N_3718,N_3537);
nor U4650 (N_4650,N_3365,N_3272);
nand U4651 (N_4651,N_3440,N_3612);
nand U4652 (N_4652,N_3512,N_3107);
and U4653 (N_4653,N_3271,N_3131);
nor U4654 (N_4654,N_3616,N_3805);
nand U4655 (N_4655,N_3908,N_3585);
and U4656 (N_4656,N_3645,N_3561);
xor U4657 (N_4657,N_3711,N_3704);
and U4658 (N_4658,N_3985,N_3001);
and U4659 (N_4659,N_3263,N_3384);
or U4660 (N_4660,N_3055,N_3740);
and U4661 (N_4661,N_3259,N_3419);
nand U4662 (N_4662,N_3852,N_3787);
and U4663 (N_4663,N_3158,N_3043);
nor U4664 (N_4664,N_3949,N_3835);
nor U4665 (N_4665,N_3403,N_3871);
nor U4666 (N_4666,N_3930,N_3018);
or U4667 (N_4667,N_3365,N_3068);
or U4668 (N_4668,N_3101,N_3796);
nand U4669 (N_4669,N_3860,N_3424);
nand U4670 (N_4670,N_3205,N_3827);
or U4671 (N_4671,N_3770,N_3740);
nand U4672 (N_4672,N_3135,N_3424);
and U4673 (N_4673,N_3665,N_3971);
xnor U4674 (N_4674,N_3093,N_3688);
nand U4675 (N_4675,N_3493,N_3006);
nand U4676 (N_4676,N_3609,N_3951);
xor U4677 (N_4677,N_3349,N_3041);
nor U4678 (N_4678,N_3262,N_3557);
nand U4679 (N_4679,N_3542,N_3054);
nand U4680 (N_4680,N_3389,N_3605);
nor U4681 (N_4681,N_3034,N_3530);
or U4682 (N_4682,N_3384,N_3323);
or U4683 (N_4683,N_3606,N_3712);
and U4684 (N_4684,N_3092,N_3405);
nand U4685 (N_4685,N_3605,N_3782);
or U4686 (N_4686,N_3289,N_3896);
nand U4687 (N_4687,N_3060,N_3867);
xor U4688 (N_4688,N_3990,N_3456);
or U4689 (N_4689,N_3308,N_3654);
or U4690 (N_4690,N_3766,N_3824);
or U4691 (N_4691,N_3229,N_3060);
nor U4692 (N_4692,N_3323,N_3338);
and U4693 (N_4693,N_3606,N_3039);
xor U4694 (N_4694,N_3941,N_3810);
nor U4695 (N_4695,N_3105,N_3113);
nand U4696 (N_4696,N_3798,N_3110);
nand U4697 (N_4697,N_3035,N_3002);
nand U4698 (N_4698,N_3355,N_3516);
xor U4699 (N_4699,N_3727,N_3654);
or U4700 (N_4700,N_3934,N_3834);
and U4701 (N_4701,N_3560,N_3333);
and U4702 (N_4702,N_3318,N_3794);
and U4703 (N_4703,N_3631,N_3298);
xor U4704 (N_4704,N_3666,N_3414);
or U4705 (N_4705,N_3736,N_3958);
nand U4706 (N_4706,N_3180,N_3326);
or U4707 (N_4707,N_3032,N_3820);
xnor U4708 (N_4708,N_3665,N_3535);
or U4709 (N_4709,N_3541,N_3670);
nand U4710 (N_4710,N_3093,N_3268);
nand U4711 (N_4711,N_3043,N_3605);
xnor U4712 (N_4712,N_3581,N_3132);
nor U4713 (N_4713,N_3503,N_3430);
and U4714 (N_4714,N_3306,N_3787);
or U4715 (N_4715,N_3984,N_3939);
and U4716 (N_4716,N_3218,N_3817);
or U4717 (N_4717,N_3807,N_3766);
nor U4718 (N_4718,N_3058,N_3667);
and U4719 (N_4719,N_3537,N_3834);
or U4720 (N_4720,N_3506,N_3575);
and U4721 (N_4721,N_3679,N_3730);
nor U4722 (N_4722,N_3112,N_3238);
or U4723 (N_4723,N_3082,N_3260);
nand U4724 (N_4724,N_3387,N_3107);
nand U4725 (N_4725,N_3362,N_3147);
nand U4726 (N_4726,N_3431,N_3372);
xnor U4727 (N_4727,N_3089,N_3433);
nand U4728 (N_4728,N_3003,N_3233);
or U4729 (N_4729,N_3141,N_3971);
or U4730 (N_4730,N_3008,N_3929);
nand U4731 (N_4731,N_3029,N_3818);
nand U4732 (N_4732,N_3794,N_3183);
and U4733 (N_4733,N_3634,N_3761);
nor U4734 (N_4734,N_3050,N_3471);
nand U4735 (N_4735,N_3330,N_3548);
or U4736 (N_4736,N_3020,N_3108);
nor U4737 (N_4737,N_3048,N_3934);
or U4738 (N_4738,N_3141,N_3246);
and U4739 (N_4739,N_3094,N_3736);
or U4740 (N_4740,N_3849,N_3329);
xnor U4741 (N_4741,N_3531,N_3249);
or U4742 (N_4742,N_3204,N_3327);
or U4743 (N_4743,N_3278,N_3017);
and U4744 (N_4744,N_3190,N_3735);
and U4745 (N_4745,N_3212,N_3605);
xnor U4746 (N_4746,N_3412,N_3011);
and U4747 (N_4747,N_3871,N_3906);
xor U4748 (N_4748,N_3257,N_3724);
nand U4749 (N_4749,N_3671,N_3444);
xnor U4750 (N_4750,N_3105,N_3342);
and U4751 (N_4751,N_3328,N_3585);
or U4752 (N_4752,N_3066,N_3845);
nor U4753 (N_4753,N_3383,N_3086);
xnor U4754 (N_4754,N_3127,N_3563);
and U4755 (N_4755,N_3642,N_3187);
and U4756 (N_4756,N_3200,N_3140);
xor U4757 (N_4757,N_3465,N_3456);
or U4758 (N_4758,N_3702,N_3798);
nand U4759 (N_4759,N_3506,N_3039);
nand U4760 (N_4760,N_3788,N_3222);
xor U4761 (N_4761,N_3687,N_3738);
nor U4762 (N_4762,N_3593,N_3753);
or U4763 (N_4763,N_3560,N_3929);
nand U4764 (N_4764,N_3902,N_3769);
xor U4765 (N_4765,N_3939,N_3548);
and U4766 (N_4766,N_3714,N_3262);
xnor U4767 (N_4767,N_3564,N_3587);
xor U4768 (N_4768,N_3797,N_3586);
or U4769 (N_4769,N_3469,N_3026);
nor U4770 (N_4770,N_3284,N_3704);
xor U4771 (N_4771,N_3681,N_3188);
nor U4772 (N_4772,N_3784,N_3077);
xor U4773 (N_4773,N_3721,N_3708);
nor U4774 (N_4774,N_3604,N_3096);
nand U4775 (N_4775,N_3748,N_3331);
nand U4776 (N_4776,N_3115,N_3595);
or U4777 (N_4777,N_3437,N_3700);
xnor U4778 (N_4778,N_3725,N_3754);
nor U4779 (N_4779,N_3699,N_3072);
or U4780 (N_4780,N_3649,N_3741);
or U4781 (N_4781,N_3336,N_3492);
xor U4782 (N_4782,N_3939,N_3073);
nand U4783 (N_4783,N_3345,N_3318);
xnor U4784 (N_4784,N_3251,N_3988);
and U4785 (N_4785,N_3826,N_3173);
or U4786 (N_4786,N_3916,N_3815);
xor U4787 (N_4787,N_3018,N_3191);
xor U4788 (N_4788,N_3155,N_3617);
nand U4789 (N_4789,N_3921,N_3664);
nor U4790 (N_4790,N_3958,N_3435);
nand U4791 (N_4791,N_3084,N_3470);
xor U4792 (N_4792,N_3850,N_3214);
and U4793 (N_4793,N_3605,N_3611);
xnor U4794 (N_4794,N_3157,N_3420);
or U4795 (N_4795,N_3707,N_3857);
nand U4796 (N_4796,N_3972,N_3799);
or U4797 (N_4797,N_3294,N_3205);
nand U4798 (N_4798,N_3958,N_3421);
nor U4799 (N_4799,N_3004,N_3059);
xnor U4800 (N_4800,N_3688,N_3034);
nor U4801 (N_4801,N_3267,N_3509);
nor U4802 (N_4802,N_3645,N_3045);
nand U4803 (N_4803,N_3331,N_3407);
nand U4804 (N_4804,N_3224,N_3334);
xnor U4805 (N_4805,N_3131,N_3843);
and U4806 (N_4806,N_3377,N_3330);
xor U4807 (N_4807,N_3602,N_3033);
or U4808 (N_4808,N_3064,N_3203);
and U4809 (N_4809,N_3550,N_3217);
nor U4810 (N_4810,N_3932,N_3841);
nor U4811 (N_4811,N_3595,N_3429);
xor U4812 (N_4812,N_3051,N_3023);
xnor U4813 (N_4813,N_3284,N_3262);
and U4814 (N_4814,N_3329,N_3821);
and U4815 (N_4815,N_3985,N_3801);
or U4816 (N_4816,N_3027,N_3959);
nand U4817 (N_4817,N_3860,N_3658);
and U4818 (N_4818,N_3834,N_3626);
xor U4819 (N_4819,N_3244,N_3164);
nand U4820 (N_4820,N_3309,N_3251);
and U4821 (N_4821,N_3760,N_3632);
and U4822 (N_4822,N_3734,N_3520);
nor U4823 (N_4823,N_3293,N_3459);
and U4824 (N_4824,N_3981,N_3315);
nor U4825 (N_4825,N_3289,N_3541);
nor U4826 (N_4826,N_3725,N_3252);
or U4827 (N_4827,N_3900,N_3052);
nand U4828 (N_4828,N_3038,N_3542);
nand U4829 (N_4829,N_3406,N_3032);
nor U4830 (N_4830,N_3661,N_3718);
xor U4831 (N_4831,N_3267,N_3254);
xor U4832 (N_4832,N_3418,N_3599);
nand U4833 (N_4833,N_3394,N_3006);
or U4834 (N_4834,N_3173,N_3802);
xor U4835 (N_4835,N_3742,N_3259);
xor U4836 (N_4836,N_3592,N_3019);
nand U4837 (N_4837,N_3592,N_3032);
and U4838 (N_4838,N_3987,N_3680);
xnor U4839 (N_4839,N_3795,N_3380);
nor U4840 (N_4840,N_3304,N_3948);
nor U4841 (N_4841,N_3387,N_3270);
nand U4842 (N_4842,N_3091,N_3403);
and U4843 (N_4843,N_3884,N_3378);
xnor U4844 (N_4844,N_3949,N_3959);
and U4845 (N_4845,N_3911,N_3867);
nand U4846 (N_4846,N_3902,N_3247);
nand U4847 (N_4847,N_3985,N_3784);
and U4848 (N_4848,N_3031,N_3509);
and U4849 (N_4849,N_3108,N_3577);
and U4850 (N_4850,N_3794,N_3418);
nor U4851 (N_4851,N_3424,N_3981);
and U4852 (N_4852,N_3135,N_3846);
xor U4853 (N_4853,N_3745,N_3544);
nor U4854 (N_4854,N_3674,N_3568);
and U4855 (N_4855,N_3396,N_3601);
nor U4856 (N_4856,N_3094,N_3151);
or U4857 (N_4857,N_3549,N_3849);
nand U4858 (N_4858,N_3209,N_3042);
xor U4859 (N_4859,N_3923,N_3078);
xnor U4860 (N_4860,N_3695,N_3038);
nand U4861 (N_4861,N_3510,N_3547);
nand U4862 (N_4862,N_3428,N_3171);
nor U4863 (N_4863,N_3755,N_3385);
and U4864 (N_4864,N_3727,N_3338);
nor U4865 (N_4865,N_3598,N_3438);
xor U4866 (N_4866,N_3562,N_3412);
nand U4867 (N_4867,N_3164,N_3227);
or U4868 (N_4868,N_3094,N_3010);
xor U4869 (N_4869,N_3490,N_3480);
and U4870 (N_4870,N_3118,N_3995);
nand U4871 (N_4871,N_3524,N_3916);
xnor U4872 (N_4872,N_3749,N_3994);
nand U4873 (N_4873,N_3827,N_3034);
and U4874 (N_4874,N_3833,N_3265);
nor U4875 (N_4875,N_3623,N_3347);
nand U4876 (N_4876,N_3103,N_3935);
xor U4877 (N_4877,N_3596,N_3002);
nand U4878 (N_4878,N_3135,N_3710);
xor U4879 (N_4879,N_3283,N_3920);
or U4880 (N_4880,N_3288,N_3006);
xnor U4881 (N_4881,N_3904,N_3366);
xnor U4882 (N_4882,N_3765,N_3779);
nand U4883 (N_4883,N_3128,N_3635);
nand U4884 (N_4884,N_3221,N_3209);
or U4885 (N_4885,N_3891,N_3259);
nand U4886 (N_4886,N_3280,N_3819);
nand U4887 (N_4887,N_3520,N_3904);
and U4888 (N_4888,N_3737,N_3580);
xor U4889 (N_4889,N_3131,N_3334);
nor U4890 (N_4890,N_3804,N_3955);
and U4891 (N_4891,N_3859,N_3735);
xor U4892 (N_4892,N_3487,N_3359);
nor U4893 (N_4893,N_3772,N_3230);
nand U4894 (N_4894,N_3405,N_3905);
or U4895 (N_4895,N_3333,N_3433);
and U4896 (N_4896,N_3279,N_3653);
nor U4897 (N_4897,N_3365,N_3970);
and U4898 (N_4898,N_3604,N_3236);
xor U4899 (N_4899,N_3460,N_3086);
nor U4900 (N_4900,N_3169,N_3589);
nor U4901 (N_4901,N_3133,N_3259);
and U4902 (N_4902,N_3263,N_3849);
nand U4903 (N_4903,N_3468,N_3450);
nand U4904 (N_4904,N_3268,N_3181);
or U4905 (N_4905,N_3264,N_3904);
nand U4906 (N_4906,N_3847,N_3881);
xnor U4907 (N_4907,N_3920,N_3393);
or U4908 (N_4908,N_3552,N_3506);
xor U4909 (N_4909,N_3861,N_3676);
or U4910 (N_4910,N_3999,N_3897);
nand U4911 (N_4911,N_3264,N_3984);
and U4912 (N_4912,N_3375,N_3975);
nand U4913 (N_4913,N_3372,N_3625);
xor U4914 (N_4914,N_3922,N_3489);
or U4915 (N_4915,N_3692,N_3785);
nand U4916 (N_4916,N_3126,N_3583);
nor U4917 (N_4917,N_3042,N_3205);
or U4918 (N_4918,N_3699,N_3572);
xor U4919 (N_4919,N_3718,N_3758);
nor U4920 (N_4920,N_3220,N_3255);
xnor U4921 (N_4921,N_3379,N_3678);
and U4922 (N_4922,N_3367,N_3752);
xnor U4923 (N_4923,N_3169,N_3356);
xor U4924 (N_4924,N_3034,N_3278);
and U4925 (N_4925,N_3638,N_3645);
xor U4926 (N_4926,N_3793,N_3461);
nor U4927 (N_4927,N_3939,N_3874);
nand U4928 (N_4928,N_3537,N_3277);
nor U4929 (N_4929,N_3722,N_3804);
xor U4930 (N_4930,N_3387,N_3034);
xnor U4931 (N_4931,N_3878,N_3934);
nor U4932 (N_4932,N_3428,N_3501);
and U4933 (N_4933,N_3300,N_3217);
nor U4934 (N_4934,N_3545,N_3960);
nor U4935 (N_4935,N_3127,N_3332);
and U4936 (N_4936,N_3194,N_3271);
or U4937 (N_4937,N_3973,N_3866);
or U4938 (N_4938,N_3868,N_3650);
and U4939 (N_4939,N_3002,N_3504);
nand U4940 (N_4940,N_3726,N_3540);
nor U4941 (N_4941,N_3965,N_3350);
nand U4942 (N_4942,N_3951,N_3493);
and U4943 (N_4943,N_3235,N_3451);
or U4944 (N_4944,N_3925,N_3407);
nor U4945 (N_4945,N_3015,N_3603);
xor U4946 (N_4946,N_3390,N_3800);
nor U4947 (N_4947,N_3985,N_3332);
nor U4948 (N_4948,N_3877,N_3847);
xnor U4949 (N_4949,N_3842,N_3316);
xnor U4950 (N_4950,N_3958,N_3365);
nand U4951 (N_4951,N_3486,N_3725);
nand U4952 (N_4952,N_3871,N_3743);
nand U4953 (N_4953,N_3576,N_3220);
xor U4954 (N_4954,N_3095,N_3258);
xor U4955 (N_4955,N_3240,N_3743);
nor U4956 (N_4956,N_3114,N_3334);
xnor U4957 (N_4957,N_3450,N_3379);
or U4958 (N_4958,N_3331,N_3469);
nand U4959 (N_4959,N_3003,N_3919);
and U4960 (N_4960,N_3821,N_3884);
xor U4961 (N_4961,N_3615,N_3284);
xnor U4962 (N_4962,N_3032,N_3461);
nor U4963 (N_4963,N_3241,N_3499);
and U4964 (N_4964,N_3553,N_3651);
and U4965 (N_4965,N_3492,N_3449);
nor U4966 (N_4966,N_3531,N_3221);
nand U4967 (N_4967,N_3868,N_3194);
nand U4968 (N_4968,N_3976,N_3119);
nand U4969 (N_4969,N_3597,N_3166);
and U4970 (N_4970,N_3122,N_3927);
xnor U4971 (N_4971,N_3327,N_3736);
or U4972 (N_4972,N_3503,N_3608);
nor U4973 (N_4973,N_3841,N_3905);
and U4974 (N_4974,N_3127,N_3343);
nor U4975 (N_4975,N_3948,N_3011);
xnor U4976 (N_4976,N_3165,N_3425);
or U4977 (N_4977,N_3457,N_3825);
nand U4978 (N_4978,N_3441,N_3102);
xor U4979 (N_4979,N_3633,N_3107);
nand U4980 (N_4980,N_3820,N_3627);
nor U4981 (N_4981,N_3053,N_3560);
nand U4982 (N_4982,N_3550,N_3140);
and U4983 (N_4983,N_3782,N_3678);
nand U4984 (N_4984,N_3254,N_3015);
xor U4985 (N_4985,N_3969,N_3447);
nand U4986 (N_4986,N_3800,N_3267);
and U4987 (N_4987,N_3631,N_3660);
and U4988 (N_4988,N_3837,N_3185);
nor U4989 (N_4989,N_3091,N_3505);
xor U4990 (N_4990,N_3275,N_3560);
nand U4991 (N_4991,N_3512,N_3695);
nand U4992 (N_4992,N_3780,N_3633);
or U4993 (N_4993,N_3235,N_3780);
nand U4994 (N_4994,N_3478,N_3024);
xor U4995 (N_4995,N_3121,N_3457);
nor U4996 (N_4996,N_3757,N_3718);
nor U4997 (N_4997,N_3374,N_3311);
and U4998 (N_4998,N_3054,N_3480);
or U4999 (N_4999,N_3731,N_3442);
and U5000 (N_5000,N_4528,N_4107);
xor U5001 (N_5001,N_4064,N_4870);
nand U5002 (N_5002,N_4799,N_4193);
or U5003 (N_5003,N_4411,N_4535);
nand U5004 (N_5004,N_4735,N_4301);
or U5005 (N_5005,N_4942,N_4075);
and U5006 (N_5006,N_4484,N_4050);
nand U5007 (N_5007,N_4544,N_4212);
nor U5008 (N_5008,N_4290,N_4277);
nand U5009 (N_5009,N_4747,N_4200);
xnor U5010 (N_5010,N_4332,N_4917);
nor U5011 (N_5011,N_4732,N_4131);
or U5012 (N_5012,N_4828,N_4175);
nor U5013 (N_5013,N_4328,N_4974);
and U5014 (N_5014,N_4526,N_4871);
xor U5015 (N_5015,N_4310,N_4795);
and U5016 (N_5016,N_4319,N_4598);
nand U5017 (N_5017,N_4971,N_4842);
nand U5018 (N_5018,N_4282,N_4731);
or U5019 (N_5019,N_4936,N_4533);
nand U5020 (N_5020,N_4362,N_4684);
nor U5021 (N_5021,N_4932,N_4509);
xor U5022 (N_5022,N_4632,N_4173);
nand U5023 (N_5023,N_4367,N_4771);
nand U5024 (N_5024,N_4647,N_4990);
nand U5025 (N_5025,N_4079,N_4292);
nor U5026 (N_5026,N_4057,N_4089);
nor U5027 (N_5027,N_4389,N_4439);
nand U5028 (N_5028,N_4031,N_4849);
or U5029 (N_5029,N_4046,N_4124);
nand U5030 (N_5030,N_4404,N_4233);
and U5031 (N_5031,N_4984,N_4775);
or U5032 (N_5032,N_4368,N_4262);
and U5033 (N_5033,N_4369,N_4495);
nand U5034 (N_5034,N_4905,N_4896);
xor U5035 (N_5035,N_4739,N_4510);
nor U5036 (N_5036,N_4016,N_4946);
or U5037 (N_5037,N_4000,N_4225);
or U5038 (N_5038,N_4140,N_4630);
or U5039 (N_5039,N_4792,N_4185);
and U5040 (N_5040,N_4530,N_4980);
xnor U5041 (N_5041,N_4897,N_4551);
or U5042 (N_5042,N_4023,N_4336);
or U5043 (N_5043,N_4348,N_4229);
or U5044 (N_5044,N_4375,N_4916);
nand U5045 (N_5045,N_4621,N_4355);
xnor U5046 (N_5046,N_4431,N_4654);
and U5047 (N_5047,N_4283,N_4781);
xor U5048 (N_5048,N_4489,N_4014);
or U5049 (N_5049,N_4331,N_4009);
and U5050 (N_5050,N_4467,N_4851);
xor U5051 (N_5051,N_4545,N_4094);
or U5052 (N_5052,N_4278,N_4886);
nor U5053 (N_5053,N_4762,N_4958);
or U5054 (N_5054,N_4561,N_4424);
and U5055 (N_5055,N_4539,N_4496);
xnor U5056 (N_5056,N_4227,N_4318);
and U5057 (N_5057,N_4821,N_4253);
and U5058 (N_5058,N_4127,N_4977);
and U5059 (N_5059,N_4201,N_4214);
or U5060 (N_5060,N_4710,N_4714);
xor U5061 (N_5061,N_4479,N_4125);
xor U5062 (N_5062,N_4066,N_4119);
nor U5063 (N_5063,N_4087,N_4835);
or U5064 (N_5064,N_4970,N_4593);
or U5065 (N_5065,N_4867,N_4651);
xor U5066 (N_5066,N_4091,N_4542);
and U5067 (N_5067,N_4302,N_4888);
nor U5068 (N_5068,N_4706,N_4846);
nor U5069 (N_5069,N_4002,N_4737);
xor U5070 (N_5070,N_4478,N_4092);
or U5071 (N_5071,N_4191,N_4518);
and U5072 (N_5072,N_4720,N_4939);
nand U5073 (N_5073,N_4655,N_4215);
nand U5074 (N_5074,N_4707,N_4379);
nor U5075 (N_5075,N_4752,N_4251);
or U5076 (N_5076,N_4156,N_4248);
or U5077 (N_5077,N_4725,N_4987);
nor U5078 (N_5078,N_4117,N_4448);
xor U5079 (N_5079,N_4113,N_4402);
or U5080 (N_5080,N_4620,N_4801);
and U5081 (N_5081,N_4154,N_4171);
xnor U5082 (N_5082,N_4826,N_4427);
nor U5083 (N_5083,N_4388,N_4321);
nand U5084 (N_5084,N_4182,N_4605);
xor U5085 (N_5085,N_4144,N_4232);
xnor U5086 (N_5086,N_4883,N_4837);
xnor U5087 (N_5087,N_4062,N_4037);
nand U5088 (N_5088,N_4054,N_4220);
and U5089 (N_5089,N_4341,N_4433);
nand U5090 (N_5090,N_4281,N_4093);
nor U5091 (N_5091,N_4418,N_4419);
and U5092 (N_5092,N_4931,N_4679);
nor U5093 (N_5093,N_4158,N_4122);
xnor U5094 (N_5094,N_4941,N_4636);
and U5095 (N_5095,N_4920,N_4738);
xnor U5096 (N_5096,N_4488,N_4757);
nand U5097 (N_5097,N_4996,N_4614);
or U5098 (N_5098,N_4698,N_4020);
and U5099 (N_5099,N_4449,N_4635);
xnor U5100 (N_5100,N_4678,N_4934);
nand U5101 (N_5101,N_4500,N_4390);
nor U5102 (N_5102,N_4574,N_4250);
nand U5103 (N_5103,N_4568,N_4313);
nand U5104 (N_5104,N_4070,N_4805);
and U5105 (N_5105,N_4299,N_4219);
or U5106 (N_5106,N_4653,N_4718);
nand U5107 (N_5107,N_4203,N_4656);
nor U5108 (N_5108,N_4257,N_4398);
nand U5109 (N_5109,N_4863,N_4463);
xnor U5110 (N_5110,N_4541,N_4470);
nor U5111 (N_5111,N_4013,N_4428);
xnor U5112 (N_5112,N_4516,N_4802);
nand U5113 (N_5113,N_4855,N_4506);
or U5114 (N_5114,N_4962,N_4167);
and U5115 (N_5115,N_4026,N_4329);
nor U5116 (N_5116,N_4304,N_4242);
nor U5117 (N_5117,N_4162,N_4715);
or U5118 (N_5118,N_4546,N_4733);
nand U5119 (N_5119,N_4447,N_4041);
nor U5120 (N_5120,N_4777,N_4454);
xor U5121 (N_5121,N_4157,N_4004);
or U5122 (N_5122,N_4322,N_4314);
nor U5123 (N_5123,N_4213,N_4692);
xor U5124 (N_5124,N_4284,N_4058);
nand U5125 (N_5125,N_4475,N_4114);
and U5126 (N_5126,N_4882,N_4409);
nor U5127 (N_5127,N_4554,N_4661);
nand U5128 (N_5128,N_4256,N_4384);
xor U5129 (N_5129,N_4817,N_4323);
nor U5130 (N_5130,N_4074,N_4560);
or U5131 (N_5131,N_4021,N_4856);
and U5132 (N_5132,N_4688,N_4209);
or U5133 (N_5133,N_4523,N_4986);
nor U5134 (N_5134,N_4105,N_4935);
and U5135 (N_5135,N_4702,N_4435);
nand U5136 (N_5136,N_4921,N_4100);
nand U5137 (N_5137,N_4018,N_4206);
and U5138 (N_5138,N_4778,N_4394);
and U5139 (N_5139,N_4749,N_4950);
or U5140 (N_5140,N_4838,N_4315);
nand U5141 (N_5141,N_4880,N_4690);
and U5142 (N_5142,N_4640,N_4589);
and U5143 (N_5143,N_4132,N_4112);
xnor U5144 (N_5144,N_4729,N_4503);
nand U5145 (N_5145,N_4486,N_4176);
nand U5146 (N_5146,N_4972,N_4997);
nand U5147 (N_5147,N_4174,N_4343);
and U5148 (N_5148,N_4774,N_4249);
nand U5149 (N_5149,N_4755,N_4421);
and U5150 (N_5150,N_4618,N_4907);
nor U5151 (N_5151,N_4833,N_4859);
and U5152 (N_5152,N_4810,N_4443);
nand U5153 (N_5153,N_4334,N_4955);
nand U5154 (N_5154,N_4045,N_4150);
nand U5155 (N_5155,N_4342,N_4832);
nand U5156 (N_5156,N_4116,N_4204);
nor U5157 (N_5157,N_4773,N_4269);
xor U5158 (N_5158,N_4121,N_4383);
nand U5159 (N_5159,N_4337,N_4584);
xor U5160 (N_5160,N_4964,N_4722);
xor U5161 (N_5161,N_4401,N_4245);
nand U5162 (N_5162,N_4730,N_4371);
or U5163 (N_5163,N_4104,N_4994);
or U5164 (N_5164,N_4999,N_4827);
xor U5165 (N_5165,N_4413,N_4874);
nor U5166 (N_5166,N_4288,N_4627);
nand U5167 (N_5167,N_4216,N_4396);
nor U5168 (N_5168,N_4060,N_4571);
nand U5169 (N_5169,N_4989,N_4316);
or U5170 (N_5170,N_4712,N_4207);
nor U5171 (N_5171,N_4196,N_4280);
xnor U5172 (N_5172,N_4937,N_4668);
nand U5173 (N_5173,N_4407,N_4746);
nor U5174 (N_5174,N_4978,N_4527);
or U5175 (N_5175,N_4370,N_4569);
nor U5176 (N_5176,N_4345,N_4436);
and U5177 (N_5177,N_4538,N_4149);
or U5178 (N_5178,N_4078,N_4294);
xnor U5179 (N_5179,N_4759,N_4643);
nor U5180 (N_5180,N_4812,N_4155);
nand U5181 (N_5181,N_4291,N_4263);
or U5182 (N_5182,N_4459,N_4372);
nand U5183 (N_5183,N_4289,N_4457);
nor U5184 (N_5184,N_4273,N_4128);
or U5185 (N_5185,N_4548,N_4797);
nor U5186 (N_5186,N_4965,N_4634);
nand U5187 (N_5187,N_4866,N_4638);
xnor U5188 (N_5188,N_4068,N_4432);
nor U5189 (N_5189,N_4160,N_4596);
xnor U5190 (N_5190,N_4308,N_4953);
xnor U5191 (N_5191,N_4648,N_4344);
nand U5192 (N_5192,N_4864,N_4504);
and U5193 (N_5193,N_4639,N_4307);
xor U5194 (N_5194,N_4611,N_4850);
and U5195 (N_5195,N_4721,N_4887);
and U5196 (N_5196,N_4052,N_4352);
or U5197 (N_5197,N_4194,N_4951);
xor U5198 (N_5198,N_4386,N_4034);
xor U5199 (N_5199,N_4255,N_4268);
xnor U5200 (N_5200,N_4305,N_4782);
and U5201 (N_5201,N_4005,N_4453);
or U5202 (N_5202,N_4086,N_4858);
nand U5203 (N_5203,N_4208,N_4025);
xnor U5204 (N_5204,N_4550,N_4303);
xnor U5205 (N_5205,N_4685,N_4734);
and U5206 (N_5206,N_4873,N_4487);
xnor U5207 (N_5207,N_4531,N_4403);
and U5208 (N_5208,N_4673,N_4320);
or U5209 (N_5209,N_4945,N_4039);
nand U5210 (N_5210,N_4082,N_4293);
and U5211 (N_5211,N_4210,N_4133);
nand U5212 (N_5212,N_4297,N_4152);
or U5213 (N_5213,N_4456,N_4575);
or U5214 (N_5214,N_4241,N_4683);
nor U5215 (N_5215,N_4508,N_4565);
nor U5216 (N_5216,N_4780,N_4361);
nand U5217 (N_5217,N_4236,N_4163);
nor U5218 (N_5218,N_4577,N_4222);
and U5219 (N_5219,N_4415,N_4146);
or U5220 (N_5220,N_4736,N_4134);
nor U5221 (N_5221,N_4750,N_4099);
nand U5222 (N_5222,N_4480,N_4686);
xor U5223 (N_5223,N_4406,N_4552);
nand U5224 (N_5224,N_4813,N_4948);
or U5225 (N_5225,N_4553,N_4108);
or U5226 (N_5226,N_4754,N_4143);
xor U5227 (N_5227,N_4033,N_4366);
nand U5228 (N_5228,N_4701,N_4011);
or U5229 (N_5229,N_4695,N_4359);
nor U5230 (N_5230,N_4603,N_4434);
and U5231 (N_5231,N_4633,N_4032);
and U5232 (N_5232,N_4335,N_4547);
nor U5233 (N_5233,N_4915,N_4615);
or U5234 (N_5234,N_4061,N_4854);
nand U5235 (N_5235,N_4610,N_4392);
or U5236 (N_5236,N_4377,N_4471);
nand U5237 (N_5237,N_4898,N_4324);
nand U5238 (N_5238,N_4363,N_4665);
nand U5239 (N_5239,N_4260,N_4816);
and U5240 (N_5240,N_4499,N_4875);
and U5241 (N_5241,N_4505,N_4689);
and U5242 (N_5242,N_4968,N_4556);
nor U5243 (N_5243,N_4764,N_4161);
nand U5244 (N_5244,N_4581,N_4072);
nand U5245 (N_5245,N_4741,N_4326);
nand U5246 (N_5246,N_4783,N_4514);
nand U5247 (N_5247,N_4520,N_4085);
nand U5248 (N_5248,N_4010,N_4599);
or U5249 (N_5249,N_4501,N_4008);
and U5250 (N_5250,N_4385,N_4007);
nor U5251 (N_5251,N_4834,N_4272);
nand U5252 (N_5252,N_4266,N_4472);
and U5253 (N_5253,N_4847,N_4682);
or U5254 (N_5254,N_4376,N_4609);
nand U5255 (N_5255,N_4769,N_4420);
or U5256 (N_5256,N_4617,N_4878);
xor U5257 (N_5257,N_4286,N_4024);
xor U5258 (N_5258,N_4613,N_4794);
nand U5259 (N_5259,N_4270,N_4889);
nor U5260 (N_5260,N_4814,N_4306);
or U5261 (N_5261,N_4570,N_4482);
nand U5262 (N_5262,N_4267,N_4728);
xnor U5263 (N_5263,N_4462,N_4006);
or U5264 (N_5264,N_4562,N_4481);
nand U5265 (N_5265,N_4669,N_4468);
or U5266 (N_5266,N_4566,N_4612);
nor U5267 (N_5267,N_4136,N_4490);
nand U5268 (N_5268,N_4238,N_4954);
nand U5269 (N_5269,N_4360,N_4914);
xor U5270 (N_5270,N_4559,N_4658);
xor U5271 (N_5271,N_4819,N_4895);
xnor U5272 (N_5272,N_4590,N_4139);
and U5273 (N_5273,N_4164,N_4199);
xnor U5274 (N_5274,N_4694,N_4903);
or U5275 (N_5275,N_4374,N_4412);
and U5276 (N_5276,N_4626,N_4317);
xnor U5277 (N_5277,N_4804,N_4624);
nand U5278 (N_5278,N_4606,N_4600);
nand U5279 (N_5279,N_4758,N_4081);
nand U5280 (N_5280,N_4029,N_4271);
xnor U5281 (N_5281,N_4727,N_4660);
nor U5282 (N_5282,N_4170,N_4998);
or U5283 (N_5283,N_4397,N_4993);
nand U5284 (N_5284,N_4697,N_4927);
or U5285 (N_5285,N_4586,N_4857);
xnor U5286 (N_5286,N_4035,N_4616);
and U5287 (N_5287,N_4168,N_4126);
nand U5288 (N_5288,N_4800,N_4373);
or U5289 (N_5289,N_4441,N_4038);
xor U5290 (N_5290,N_4988,N_4549);
nor U5291 (N_5291,N_4423,N_4925);
nand U5292 (N_5292,N_4952,N_4844);
xor U5293 (N_5293,N_4451,N_4153);
nor U5294 (N_5294,N_4760,N_4346);
nor U5295 (N_5295,N_4221,N_4963);
nor U5296 (N_5296,N_4090,N_4142);
nor U5297 (N_5297,N_4521,N_4666);
and U5298 (N_5298,N_4400,N_4159);
xnor U5299 (N_5299,N_4452,N_4576);
xnor U5300 (N_5300,N_4027,N_4726);
nand U5301 (N_5301,N_4298,N_4073);
nor U5302 (N_5302,N_4492,N_4218);
xnor U5303 (N_5303,N_4195,N_4865);
and U5304 (N_5304,N_4525,N_4943);
or U5305 (N_5305,N_4675,N_4637);
nand U5306 (N_5306,N_4455,N_4340);
xnor U5307 (N_5307,N_4354,N_4976);
xor U5308 (N_5308,N_4776,N_4077);
nand U5309 (N_5309,N_4169,N_4223);
nor U5310 (N_5310,N_4391,N_4130);
nor U5311 (N_5311,N_4098,N_4664);
nor U5312 (N_5312,N_4017,N_4183);
nand U5313 (N_5313,N_4900,N_4312);
nor U5314 (N_5314,N_4186,N_4476);
nand U5315 (N_5315,N_4123,N_4350);
nand U5316 (N_5316,N_4069,N_4822);
or U5317 (N_5317,N_4879,N_4982);
or U5318 (N_5318,N_4497,N_4843);
nor U5319 (N_5319,N_4908,N_4330);
and U5320 (N_5320,N_4719,N_4949);
nand U5321 (N_5321,N_4519,N_4217);
or U5322 (N_5322,N_4180,N_4894);
xnor U5323 (N_5323,N_4101,N_4680);
and U5324 (N_5324,N_4043,N_4422);
or U5325 (N_5325,N_4437,N_4237);
xor U5326 (N_5326,N_4744,N_4458);
and U5327 (N_5327,N_4670,N_4940);
or U5328 (N_5328,N_4557,N_4309);
nor U5329 (N_5329,N_4166,N_4063);
and U5330 (N_5330,N_4876,N_4469);
nor U5331 (N_5331,N_4790,N_4957);
nand U5332 (N_5332,N_4071,N_4172);
or U5333 (N_5333,N_4440,N_4053);
nor U5334 (N_5334,N_4608,N_4691);
xor U5335 (N_5335,N_4923,N_4973);
xor U5336 (N_5336,N_4483,N_4338);
nand U5337 (N_5337,N_4646,N_4198);
xnor U5338 (N_5338,N_4587,N_4959);
and U5339 (N_5339,N_4244,N_4364);
and U5340 (N_5340,N_4625,N_4667);
or U5341 (N_5341,N_4147,N_4788);
nand U5342 (N_5342,N_4051,N_4770);
or U5343 (N_5343,N_4408,N_4365);
nand U5344 (N_5344,N_4912,N_4967);
and U5345 (N_5345,N_4387,N_4573);
nand U5346 (N_5346,N_4485,N_4507);
nor U5347 (N_5347,N_4595,N_4787);
or U5348 (N_5348,N_4239,N_4189);
and U5349 (N_5349,N_4823,N_4202);
and U5350 (N_5350,N_4382,N_4891);
nand U5351 (N_5351,N_4477,N_4929);
nand U5352 (N_5352,N_4188,N_4899);
xor U5353 (N_5353,N_4681,N_4096);
nor U5354 (N_5354,N_4676,N_4275);
or U5355 (N_5355,N_4522,N_4243);
nand U5356 (N_5356,N_4818,N_4055);
and U5357 (N_5357,N_4784,N_4474);
nand U5358 (N_5358,N_4532,N_4111);
nand U5359 (N_5359,N_4177,N_4141);
or U5360 (N_5360,N_4264,N_4502);
or U5361 (N_5361,N_4567,N_4393);
nand U5362 (N_5362,N_4724,N_4279);
xor U5363 (N_5363,N_4181,N_4926);
nor U5364 (N_5364,N_4913,N_4930);
and U5365 (N_5365,N_4657,N_4036);
nand U5366 (N_5366,N_4641,N_4911);
nand U5367 (N_5367,N_4713,N_4353);
or U5368 (N_5368,N_4357,N_4430);
and U5369 (N_5369,N_4743,N_4687);
or U5370 (N_5370,N_4740,N_4498);
xor U5371 (N_5371,N_4869,N_4840);
and U5372 (N_5372,N_4426,N_4659);
or U5373 (N_5373,N_4700,N_4966);
nand U5374 (N_5374,N_4644,N_4347);
nor U5375 (N_5375,N_4751,N_4517);
nor U5376 (N_5376,N_4247,N_4022);
nand U5377 (N_5377,N_4956,N_4473);
nor U5378 (N_5378,N_4138,N_4806);
or U5379 (N_5379,N_4356,N_4534);
and U5380 (N_5380,N_4325,N_4597);
xnor U5381 (N_5381,N_4704,N_4056);
nand U5382 (N_5382,N_4830,N_4672);
or U5383 (N_5383,N_4358,N_4872);
nand U5384 (N_5384,N_4265,N_4540);
or U5385 (N_5385,N_4578,N_4829);
nor U5386 (N_5386,N_4919,N_4761);
xnor U5387 (N_5387,N_4230,N_4494);
nor U5388 (N_5388,N_4811,N_4555);
nand U5389 (N_5389,N_4572,N_4803);
and U5390 (N_5390,N_4622,N_4042);
xnor U5391 (N_5391,N_4228,N_4028);
xnor U5392 (N_5392,N_4118,N_4148);
nand U5393 (N_5393,N_4327,N_4395);
and U5394 (N_5394,N_4461,N_4095);
and U5395 (N_5395,N_4960,N_4645);
nor U5396 (N_5396,N_4197,N_4991);
nand U5397 (N_5397,N_4466,N_4493);
xor U5398 (N_5398,N_4115,N_4861);
xor U5399 (N_5399,N_4088,N_4261);
nor U5400 (N_5400,N_4080,N_4629);
nor U5401 (N_5401,N_4604,N_4444);
xnor U5402 (N_5402,N_4465,N_4287);
nand U5403 (N_5403,N_4097,N_4594);
or U5404 (N_5404,N_4992,N_4120);
nor U5405 (N_5405,N_4512,N_4602);
xnor U5406 (N_5406,N_4258,N_4254);
xnor U5407 (N_5407,N_4129,N_4145);
nand U5408 (N_5408,N_4807,N_4786);
nand U5409 (N_5409,N_4065,N_4893);
nor U5410 (N_5410,N_4563,N_4179);
nor U5411 (N_5411,N_4717,N_4748);
nor U5412 (N_5412,N_4579,N_4076);
nor U5413 (N_5413,N_4592,N_4924);
nand U5414 (N_5414,N_4848,N_4909);
nand U5415 (N_5415,N_4333,N_4631);
nor U5416 (N_5416,N_4445,N_4623);
nand U5417 (N_5417,N_4723,N_4607);
nand U5418 (N_5418,N_4947,N_4184);
nand U5419 (N_5419,N_4785,N_4137);
or U5420 (N_5420,N_4853,N_4106);
and U5421 (N_5421,N_4693,N_4979);
nor U5422 (N_5422,N_4711,N_4414);
and U5423 (N_5423,N_4151,N_4663);
nand U5424 (N_5424,N_4938,N_4588);
nor U5425 (N_5425,N_4928,N_4235);
or U5426 (N_5426,N_4628,N_4580);
or U5427 (N_5427,N_4015,N_4049);
nand U5428 (N_5428,N_4083,N_4791);
nand U5429 (N_5429,N_4902,N_4652);
and U5430 (N_5430,N_4862,N_4558);
xnor U5431 (N_5431,N_4001,N_4524);
nand U5432 (N_5432,N_4793,N_4918);
or U5433 (N_5433,N_4378,N_4809);
or U5434 (N_5434,N_4852,N_4564);
nor U5435 (N_5435,N_4300,N_4696);
or U5436 (N_5436,N_4351,N_4906);
nor U5437 (N_5437,N_4399,N_4981);
nor U5438 (N_5438,N_4178,N_4767);
nand U5439 (N_5439,N_4808,N_4234);
and U5440 (N_5440,N_4619,N_4190);
xnor U5441 (N_5441,N_4276,N_4048);
or U5442 (N_5442,N_4380,N_4815);
xnor U5443 (N_5443,N_4044,N_4019);
nand U5444 (N_5444,N_4529,N_4825);
xor U5445 (N_5445,N_4969,N_4904);
nand U5446 (N_5446,N_4796,N_4933);
nor U5447 (N_5447,N_4311,N_4885);
nand U5448 (N_5448,N_4513,N_4922);
or U5449 (N_5449,N_4030,N_4779);
or U5450 (N_5450,N_4798,N_4841);
nand U5451 (N_5451,N_4429,N_4716);
xor U5452 (N_5452,N_4884,N_4836);
nand U5453 (N_5453,N_4464,N_4084);
or U5454 (N_5454,N_4766,N_4789);
nor U5455 (N_5455,N_4425,N_4491);
nand U5456 (N_5456,N_4768,N_4601);
nor U5457 (N_5457,N_4662,N_4642);
nand U5458 (N_5458,N_4410,N_4831);
xnor U5459 (N_5459,N_4583,N_4881);
or U5460 (N_5460,N_4003,N_4585);
nand U5461 (N_5461,N_4860,N_4446);
xor U5462 (N_5462,N_4753,N_4416);
nand U5463 (N_5463,N_4677,N_4824);
nor U5464 (N_5464,N_4868,N_4187);
xnor U5465 (N_5465,N_4205,N_4059);
or U5466 (N_5466,N_4983,N_4438);
nor U5467 (N_5467,N_4109,N_4820);
and U5468 (N_5468,N_4582,N_4274);
nand U5469 (N_5469,N_4450,N_4047);
nor U5470 (N_5470,N_4910,N_4224);
or U5471 (N_5471,N_4192,N_4240);
xor U5472 (N_5472,N_4763,N_4537);
and U5473 (N_5473,N_4995,N_4349);
or U5474 (N_5474,N_4961,N_4442);
nand U5475 (N_5475,N_4975,N_4296);
and U5476 (N_5476,N_4252,N_4649);
and U5477 (N_5477,N_4742,N_4405);
xnor U5478 (N_5478,N_4135,N_4745);
nor U5479 (N_5479,N_4839,N_4103);
nand U5480 (N_5480,N_4515,N_4417);
xor U5481 (N_5481,N_4339,N_4165);
and U5482 (N_5482,N_4511,N_4765);
nand U5483 (N_5483,N_4102,N_4259);
or U5484 (N_5484,N_4709,N_4012);
or U5485 (N_5485,N_4543,N_4536);
or U5486 (N_5486,N_4460,N_4231);
nor U5487 (N_5487,N_4890,N_4067);
or U5488 (N_5488,N_4040,N_4772);
and U5489 (N_5489,N_4703,N_4671);
nor U5490 (N_5490,N_4285,N_4699);
xor U5491 (N_5491,N_4845,N_4944);
nor U5492 (N_5492,N_4892,N_4650);
and U5493 (N_5493,N_4708,N_4985);
xnor U5494 (N_5494,N_4877,N_4226);
nand U5495 (N_5495,N_4591,N_4705);
nand U5496 (N_5496,N_4295,N_4674);
xor U5497 (N_5497,N_4211,N_4901);
nand U5498 (N_5498,N_4381,N_4756);
nor U5499 (N_5499,N_4246,N_4110);
xor U5500 (N_5500,N_4528,N_4032);
or U5501 (N_5501,N_4026,N_4145);
or U5502 (N_5502,N_4890,N_4589);
nor U5503 (N_5503,N_4079,N_4621);
and U5504 (N_5504,N_4676,N_4600);
or U5505 (N_5505,N_4275,N_4737);
nor U5506 (N_5506,N_4639,N_4602);
and U5507 (N_5507,N_4339,N_4278);
nor U5508 (N_5508,N_4500,N_4982);
xnor U5509 (N_5509,N_4144,N_4606);
nor U5510 (N_5510,N_4094,N_4791);
or U5511 (N_5511,N_4033,N_4987);
nor U5512 (N_5512,N_4483,N_4473);
xnor U5513 (N_5513,N_4253,N_4467);
nor U5514 (N_5514,N_4847,N_4612);
and U5515 (N_5515,N_4240,N_4405);
or U5516 (N_5516,N_4551,N_4442);
nand U5517 (N_5517,N_4322,N_4103);
nand U5518 (N_5518,N_4478,N_4662);
xor U5519 (N_5519,N_4369,N_4817);
xor U5520 (N_5520,N_4440,N_4680);
xor U5521 (N_5521,N_4673,N_4176);
and U5522 (N_5522,N_4591,N_4538);
xor U5523 (N_5523,N_4613,N_4340);
nand U5524 (N_5524,N_4856,N_4470);
nor U5525 (N_5525,N_4170,N_4073);
and U5526 (N_5526,N_4242,N_4430);
nor U5527 (N_5527,N_4236,N_4382);
and U5528 (N_5528,N_4000,N_4340);
nand U5529 (N_5529,N_4297,N_4949);
and U5530 (N_5530,N_4660,N_4005);
or U5531 (N_5531,N_4105,N_4577);
nor U5532 (N_5532,N_4603,N_4644);
nand U5533 (N_5533,N_4346,N_4668);
nand U5534 (N_5534,N_4879,N_4028);
nand U5535 (N_5535,N_4121,N_4600);
xor U5536 (N_5536,N_4055,N_4935);
nand U5537 (N_5537,N_4334,N_4479);
nand U5538 (N_5538,N_4681,N_4905);
xor U5539 (N_5539,N_4761,N_4233);
nor U5540 (N_5540,N_4836,N_4838);
and U5541 (N_5541,N_4850,N_4350);
and U5542 (N_5542,N_4079,N_4075);
xor U5543 (N_5543,N_4691,N_4647);
nor U5544 (N_5544,N_4057,N_4098);
and U5545 (N_5545,N_4008,N_4794);
or U5546 (N_5546,N_4978,N_4482);
or U5547 (N_5547,N_4939,N_4656);
and U5548 (N_5548,N_4961,N_4114);
xor U5549 (N_5549,N_4202,N_4116);
nor U5550 (N_5550,N_4146,N_4196);
xnor U5551 (N_5551,N_4088,N_4500);
xnor U5552 (N_5552,N_4746,N_4326);
and U5553 (N_5553,N_4078,N_4387);
and U5554 (N_5554,N_4694,N_4881);
or U5555 (N_5555,N_4910,N_4621);
nor U5556 (N_5556,N_4461,N_4541);
nor U5557 (N_5557,N_4238,N_4353);
nand U5558 (N_5558,N_4194,N_4526);
and U5559 (N_5559,N_4475,N_4683);
or U5560 (N_5560,N_4600,N_4730);
or U5561 (N_5561,N_4281,N_4035);
xnor U5562 (N_5562,N_4005,N_4335);
or U5563 (N_5563,N_4906,N_4933);
nor U5564 (N_5564,N_4862,N_4071);
and U5565 (N_5565,N_4896,N_4037);
and U5566 (N_5566,N_4192,N_4959);
nand U5567 (N_5567,N_4454,N_4437);
xor U5568 (N_5568,N_4114,N_4946);
or U5569 (N_5569,N_4154,N_4739);
and U5570 (N_5570,N_4360,N_4824);
or U5571 (N_5571,N_4360,N_4212);
xor U5572 (N_5572,N_4107,N_4771);
xnor U5573 (N_5573,N_4795,N_4377);
xor U5574 (N_5574,N_4068,N_4547);
xor U5575 (N_5575,N_4674,N_4301);
or U5576 (N_5576,N_4449,N_4303);
nand U5577 (N_5577,N_4358,N_4445);
and U5578 (N_5578,N_4136,N_4272);
xnor U5579 (N_5579,N_4192,N_4588);
and U5580 (N_5580,N_4296,N_4468);
nand U5581 (N_5581,N_4498,N_4693);
nand U5582 (N_5582,N_4572,N_4690);
nand U5583 (N_5583,N_4993,N_4082);
or U5584 (N_5584,N_4089,N_4644);
xor U5585 (N_5585,N_4459,N_4685);
nand U5586 (N_5586,N_4619,N_4546);
or U5587 (N_5587,N_4763,N_4755);
xnor U5588 (N_5588,N_4266,N_4240);
nor U5589 (N_5589,N_4263,N_4888);
or U5590 (N_5590,N_4578,N_4953);
and U5591 (N_5591,N_4593,N_4352);
nor U5592 (N_5592,N_4165,N_4908);
and U5593 (N_5593,N_4516,N_4578);
nand U5594 (N_5594,N_4660,N_4714);
nor U5595 (N_5595,N_4342,N_4293);
and U5596 (N_5596,N_4209,N_4532);
and U5597 (N_5597,N_4700,N_4049);
and U5598 (N_5598,N_4628,N_4296);
and U5599 (N_5599,N_4064,N_4801);
nand U5600 (N_5600,N_4323,N_4220);
nor U5601 (N_5601,N_4462,N_4740);
and U5602 (N_5602,N_4711,N_4291);
nor U5603 (N_5603,N_4357,N_4656);
nand U5604 (N_5604,N_4672,N_4995);
xor U5605 (N_5605,N_4837,N_4717);
nor U5606 (N_5606,N_4054,N_4427);
xor U5607 (N_5607,N_4833,N_4388);
xnor U5608 (N_5608,N_4316,N_4652);
or U5609 (N_5609,N_4864,N_4176);
nor U5610 (N_5610,N_4370,N_4677);
or U5611 (N_5611,N_4693,N_4820);
xor U5612 (N_5612,N_4830,N_4701);
or U5613 (N_5613,N_4335,N_4143);
xnor U5614 (N_5614,N_4007,N_4193);
nor U5615 (N_5615,N_4145,N_4677);
nor U5616 (N_5616,N_4175,N_4344);
or U5617 (N_5617,N_4178,N_4289);
or U5618 (N_5618,N_4405,N_4816);
xor U5619 (N_5619,N_4007,N_4648);
nor U5620 (N_5620,N_4208,N_4844);
nand U5621 (N_5621,N_4947,N_4589);
or U5622 (N_5622,N_4304,N_4572);
xor U5623 (N_5623,N_4356,N_4421);
xnor U5624 (N_5624,N_4450,N_4802);
or U5625 (N_5625,N_4981,N_4240);
and U5626 (N_5626,N_4985,N_4231);
or U5627 (N_5627,N_4436,N_4022);
xor U5628 (N_5628,N_4254,N_4356);
xor U5629 (N_5629,N_4164,N_4197);
and U5630 (N_5630,N_4364,N_4196);
or U5631 (N_5631,N_4242,N_4801);
and U5632 (N_5632,N_4939,N_4396);
xor U5633 (N_5633,N_4932,N_4114);
or U5634 (N_5634,N_4349,N_4173);
nand U5635 (N_5635,N_4978,N_4214);
xor U5636 (N_5636,N_4183,N_4730);
nand U5637 (N_5637,N_4305,N_4461);
or U5638 (N_5638,N_4469,N_4643);
xnor U5639 (N_5639,N_4922,N_4647);
or U5640 (N_5640,N_4870,N_4985);
nand U5641 (N_5641,N_4229,N_4536);
or U5642 (N_5642,N_4549,N_4474);
nor U5643 (N_5643,N_4650,N_4139);
xnor U5644 (N_5644,N_4837,N_4215);
xor U5645 (N_5645,N_4243,N_4406);
nor U5646 (N_5646,N_4916,N_4225);
nand U5647 (N_5647,N_4814,N_4056);
xnor U5648 (N_5648,N_4014,N_4266);
nand U5649 (N_5649,N_4996,N_4055);
nor U5650 (N_5650,N_4699,N_4951);
or U5651 (N_5651,N_4123,N_4268);
nand U5652 (N_5652,N_4164,N_4134);
nor U5653 (N_5653,N_4642,N_4432);
xnor U5654 (N_5654,N_4713,N_4827);
and U5655 (N_5655,N_4933,N_4617);
xnor U5656 (N_5656,N_4818,N_4554);
and U5657 (N_5657,N_4537,N_4433);
nor U5658 (N_5658,N_4284,N_4494);
xor U5659 (N_5659,N_4202,N_4226);
and U5660 (N_5660,N_4265,N_4724);
or U5661 (N_5661,N_4117,N_4101);
or U5662 (N_5662,N_4674,N_4199);
nor U5663 (N_5663,N_4440,N_4429);
xor U5664 (N_5664,N_4868,N_4174);
nor U5665 (N_5665,N_4006,N_4981);
nand U5666 (N_5666,N_4388,N_4172);
and U5667 (N_5667,N_4564,N_4655);
or U5668 (N_5668,N_4042,N_4291);
or U5669 (N_5669,N_4864,N_4187);
or U5670 (N_5670,N_4879,N_4209);
or U5671 (N_5671,N_4064,N_4497);
xor U5672 (N_5672,N_4975,N_4929);
and U5673 (N_5673,N_4513,N_4881);
nand U5674 (N_5674,N_4559,N_4530);
nand U5675 (N_5675,N_4148,N_4692);
nor U5676 (N_5676,N_4222,N_4175);
and U5677 (N_5677,N_4828,N_4285);
or U5678 (N_5678,N_4208,N_4685);
nor U5679 (N_5679,N_4570,N_4624);
and U5680 (N_5680,N_4351,N_4276);
and U5681 (N_5681,N_4906,N_4229);
nor U5682 (N_5682,N_4260,N_4179);
nand U5683 (N_5683,N_4471,N_4737);
nand U5684 (N_5684,N_4477,N_4021);
and U5685 (N_5685,N_4589,N_4815);
or U5686 (N_5686,N_4231,N_4472);
nor U5687 (N_5687,N_4641,N_4217);
xor U5688 (N_5688,N_4934,N_4530);
and U5689 (N_5689,N_4930,N_4870);
nor U5690 (N_5690,N_4482,N_4883);
nor U5691 (N_5691,N_4632,N_4278);
nand U5692 (N_5692,N_4901,N_4171);
or U5693 (N_5693,N_4885,N_4067);
nor U5694 (N_5694,N_4948,N_4334);
or U5695 (N_5695,N_4176,N_4479);
nand U5696 (N_5696,N_4230,N_4504);
nand U5697 (N_5697,N_4479,N_4643);
xnor U5698 (N_5698,N_4900,N_4201);
or U5699 (N_5699,N_4471,N_4489);
nand U5700 (N_5700,N_4731,N_4589);
or U5701 (N_5701,N_4887,N_4752);
nand U5702 (N_5702,N_4138,N_4262);
xor U5703 (N_5703,N_4743,N_4158);
nor U5704 (N_5704,N_4783,N_4941);
nor U5705 (N_5705,N_4023,N_4122);
and U5706 (N_5706,N_4473,N_4355);
nand U5707 (N_5707,N_4241,N_4373);
and U5708 (N_5708,N_4230,N_4212);
or U5709 (N_5709,N_4049,N_4795);
nand U5710 (N_5710,N_4036,N_4076);
or U5711 (N_5711,N_4455,N_4625);
nor U5712 (N_5712,N_4353,N_4153);
nand U5713 (N_5713,N_4893,N_4480);
xnor U5714 (N_5714,N_4461,N_4349);
nand U5715 (N_5715,N_4793,N_4114);
xnor U5716 (N_5716,N_4260,N_4683);
nor U5717 (N_5717,N_4885,N_4182);
xnor U5718 (N_5718,N_4166,N_4649);
xor U5719 (N_5719,N_4603,N_4237);
or U5720 (N_5720,N_4962,N_4654);
and U5721 (N_5721,N_4982,N_4246);
or U5722 (N_5722,N_4882,N_4060);
nand U5723 (N_5723,N_4433,N_4897);
nor U5724 (N_5724,N_4984,N_4853);
nor U5725 (N_5725,N_4903,N_4867);
or U5726 (N_5726,N_4647,N_4441);
or U5727 (N_5727,N_4219,N_4802);
nand U5728 (N_5728,N_4631,N_4892);
and U5729 (N_5729,N_4953,N_4152);
nor U5730 (N_5730,N_4358,N_4428);
or U5731 (N_5731,N_4516,N_4856);
or U5732 (N_5732,N_4797,N_4032);
or U5733 (N_5733,N_4700,N_4883);
and U5734 (N_5734,N_4933,N_4916);
or U5735 (N_5735,N_4915,N_4895);
nand U5736 (N_5736,N_4993,N_4985);
and U5737 (N_5737,N_4037,N_4235);
xor U5738 (N_5738,N_4430,N_4137);
or U5739 (N_5739,N_4049,N_4392);
nor U5740 (N_5740,N_4039,N_4365);
nand U5741 (N_5741,N_4484,N_4367);
and U5742 (N_5742,N_4491,N_4567);
nor U5743 (N_5743,N_4594,N_4154);
nand U5744 (N_5744,N_4052,N_4130);
xnor U5745 (N_5745,N_4251,N_4858);
and U5746 (N_5746,N_4460,N_4187);
or U5747 (N_5747,N_4174,N_4119);
or U5748 (N_5748,N_4741,N_4522);
xor U5749 (N_5749,N_4661,N_4680);
or U5750 (N_5750,N_4085,N_4882);
nand U5751 (N_5751,N_4523,N_4322);
nand U5752 (N_5752,N_4818,N_4573);
and U5753 (N_5753,N_4998,N_4693);
nand U5754 (N_5754,N_4056,N_4842);
nor U5755 (N_5755,N_4399,N_4849);
and U5756 (N_5756,N_4753,N_4519);
nor U5757 (N_5757,N_4299,N_4360);
xnor U5758 (N_5758,N_4508,N_4992);
and U5759 (N_5759,N_4962,N_4399);
nand U5760 (N_5760,N_4309,N_4088);
xor U5761 (N_5761,N_4323,N_4625);
nand U5762 (N_5762,N_4945,N_4277);
nor U5763 (N_5763,N_4654,N_4334);
xnor U5764 (N_5764,N_4246,N_4862);
xor U5765 (N_5765,N_4080,N_4537);
xor U5766 (N_5766,N_4802,N_4572);
or U5767 (N_5767,N_4547,N_4549);
nor U5768 (N_5768,N_4289,N_4781);
xnor U5769 (N_5769,N_4872,N_4196);
nand U5770 (N_5770,N_4545,N_4271);
or U5771 (N_5771,N_4211,N_4485);
nor U5772 (N_5772,N_4396,N_4404);
xnor U5773 (N_5773,N_4630,N_4609);
nor U5774 (N_5774,N_4504,N_4218);
nand U5775 (N_5775,N_4843,N_4261);
xnor U5776 (N_5776,N_4384,N_4083);
nand U5777 (N_5777,N_4828,N_4976);
nand U5778 (N_5778,N_4417,N_4002);
nor U5779 (N_5779,N_4437,N_4812);
nor U5780 (N_5780,N_4892,N_4695);
or U5781 (N_5781,N_4860,N_4255);
nand U5782 (N_5782,N_4249,N_4737);
and U5783 (N_5783,N_4674,N_4403);
nand U5784 (N_5784,N_4679,N_4782);
nor U5785 (N_5785,N_4149,N_4456);
or U5786 (N_5786,N_4591,N_4968);
and U5787 (N_5787,N_4018,N_4056);
nor U5788 (N_5788,N_4969,N_4680);
nor U5789 (N_5789,N_4480,N_4648);
or U5790 (N_5790,N_4542,N_4811);
and U5791 (N_5791,N_4877,N_4967);
xor U5792 (N_5792,N_4842,N_4090);
and U5793 (N_5793,N_4381,N_4978);
and U5794 (N_5794,N_4420,N_4650);
and U5795 (N_5795,N_4548,N_4733);
and U5796 (N_5796,N_4516,N_4612);
xnor U5797 (N_5797,N_4634,N_4385);
and U5798 (N_5798,N_4434,N_4365);
nor U5799 (N_5799,N_4032,N_4016);
or U5800 (N_5800,N_4981,N_4172);
nand U5801 (N_5801,N_4910,N_4870);
nand U5802 (N_5802,N_4854,N_4989);
xnor U5803 (N_5803,N_4318,N_4941);
or U5804 (N_5804,N_4493,N_4302);
nand U5805 (N_5805,N_4975,N_4388);
or U5806 (N_5806,N_4970,N_4558);
nand U5807 (N_5807,N_4861,N_4469);
or U5808 (N_5808,N_4049,N_4538);
nand U5809 (N_5809,N_4872,N_4328);
nor U5810 (N_5810,N_4994,N_4572);
xnor U5811 (N_5811,N_4341,N_4376);
nor U5812 (N_5812,N_4047,N_4949);
or U5813 (N_5813,N_4165,N_4167);
nand U5814 (N_5814,N_4655,N_4992);
nand U5815 (N_5815,N_4163,N_4868);
xnor U5816 (N_5816,N_4586,N_4990);
xnor U5817 (N_5817,N_4826,N_4159);
xor U5818 (N_5818,N_4292,N_4378);
xor U5819 (N_5819,N_4376,N_4677);
nand U5820 (N_5820,N_4259,N_4852);
nor U5821 (N_5821,N_4471,N_4996);
and U5822 (N_5822,N_4513,N_4063);
and U5823 (N_5823,N_4298,N_4899);
or U5824 (N_5824,N_4642,N_4066);
nor U5825 (N_5825,N_4542,N_4428);
nand U5826 (N_5826,N_4834,N_4483);
nand U5827 (N_5827,N_4846,N_4368);
and U5828 (N_5828,N_4116,N_4685);
nand U5829 (N_5829,N_4581,N_4760);
and U5830 (N_5830,N_4444,N_4862);
xnor U5831 (N_5831,N_4579,N_4904);
or U5832 (N_5832,N_4702,N_4511);
and U5833 (N_5833,N_4573,N_4325);
and U5834 (N_5834,N_4815,N_4175);
xnor U5835 (N_5835,N_4672,N_4443);
xor U5836 (N_5836,N_4429,N_4593);
xor U5837 (N_5837,N_4465,N_4518);
nor U5838 (N_5838,N_4584,N_4920);
and U5839 (N_5839,N_4770,N_4784);
xnor U5840 (N_5840,N_4985,N_4617);
nand U5841 (N_5841,N_4916,N_4376);
xnor U5842 (N_5842,N_4224,N_4346);
xnor U5843 (N_5843,N_4177,N_4772);
and U5844 (N_5844,N_4853,N_4999);
or U5845 (N_5845,N_4887,N_4532);
nand U5846 (N_5846,N_4498,N_4927);
and U5847 (N_5847,N_4949,N_4838);
nor U5848 (N_5848,N_4329,N_4985);
nand U5849 (N_5849,N_4640,N_4182);
xnor U5850 (N_5850,N_4728,N_4615);
nor U5851 (N_5851,N_4341,N_4146);
nor U5852 (N_5852,N_4882,N_4460);
nand U5853 (N_5853,N_4175,N_4457);
or U5854 (N_5854,N_4309,N_4363);
nand U5855 (N_5855,N_4148,N_4514);
xnor U5856 (N_5856,N_4468,N_4387);
nor U5857 (N_5857,N_4733,N_4768);
nand U5858 (N_5858,N_4532,N_4361);
nor U5859 (N_5859,N_4280,N_4095);
nand U5860 (N_5860,N_4279,N_4949);
nor U5861 (N_5861,N_4214,N_4857);
or U5862 (N_5862,N_4395,N_4675);
or U5863 (N_5863,N_4829,N_4591);
nand U5864 (N_5864,N_4575,N_4402);
or U5865 (N_5865,N_4160,N_4658);
or U5866 (N_5866,N_4834,N_4879);
nor U5867 (N_5867,N_4415,N_4686);
or U5868 (N_5868,N_4259,N_4529);
nand U5869 (N_5869,N_4159,N_4790);
xnor U5870 (N_5870,N_4817,N_4007);
nand U5871 (N_5871,N_4904,N_4010);
nor U5872 (N_5872,N_4233,N_4467);
nor U5873 (N_5873,N_4270,N_4682);
xnor U5874 (N_5874,N_4466,N_4437);
or U5875 (N_5875,N_4426,N_4764);
xnor U5876 (N_5876,N_4035,N_4047);
xnor U5877 (N_5877,N_4434,N_4855);
or U5878 (N_5878,N_4391,N_4924);
and U5879 (N_5879,N_4702,N_4068);
xor U5880 (N_5880,N_4446,N_4288);
xnor U5881 (N_5881,N_4374,N_4064);
nand U5882 (N_5882,N_4950,N_4583);
nand U5883 (N_5883,N_4199,N_4429);
nand U5884 (N_5884,N_4455,N_4683);
and U5885 (N_5885,N_4986,N_4216);
nand U5886 (N_5886,N_4874,N_4456);
or U5887 (N_5887,N_4571,N_4575);
nand U5888 (N_5888,N_4610,N_4032);
xor U5889 (N_5889,N_4351,N_4927);
and U5890 (N_5890,N_4642,N_4762);
xnor U5891 (N_5891,N_4103,N_4568);
or U5892 (N_5892,N_4247,N_4004);
nor U5893 (N_5893,N_4627,N_4409);
xor U5894 (N_5894,N_4755,N_4220);
nand U5895 (N_5895,N_4113,N_4684);
and U5896 (N_5896,N_4183,N_4120);
and U5897 (N_5897,N_4840,N_4075);
xnor U5898 (N_5898,N_4160,N_4816);
nand U5899 (N_5899,N_4582,N_4655);
nor U5900 (N_5900,N_4809,N_4630);
nor U5901 (N_5901,N_4830,N_4562);
xnor U5902 (N_5902,N_4022,N_4694);
nor U5903 (N_5903,N_4895,N_4710);
and U5904 (N_5904,N_4572,N_4504);
xor U5905 (N_5905,N_4977,N_4939);
nor U5906 (N_5906,N_4533,N_4570);
nor U5907 (N_5907,N_4483,N_4843);
xor U5908 (N_5908,N_4230,N_4087);
xnor U5909 (N_5909,N_4435,N_4009);
nand U5910 (N_5910,N_4809,N_4417);
nand U5911 (N_5911,N_4464,N_4575);
and U5912 (N_5912,N_4651,N_4225);
xnor U5913 (N_5913,N_4452,N_4740);
xor U5914 (N_5914,N_4884,N_4549);
and U5915 (N_5915,N_4907,N_4178);
nand U5916 (N_5916,N_4132,N_4353);
nand U5917 (N_5917,N_4134,N_4168);
nor U5918 (N_5918,N_4445,N_4807);
nor U5919 (N_5919,N_4640,N_4588);
xor U5920 (N_5920,N_4121,N_4922);
or U5921 (N_5921,N_4327,N_4364);
nand U5922 (N_5922,N_4033,N_4510);
xor U5923 (N_5923,N_4188,N_4782);
xor U5924 (N_5924,N_4136,N_4383);
xor U5925 (N_5925,N_4145,N_4162);
or U5926 (N_5926,N_4575,N_4009);
xor U5927 (N_5927,N_4835,N_4684);
and U5928 (N_5928,N_4730,N_4513);
and U5929 (N_5929,N_4839,N_4871);
and U5930 (N_5930,N_4115,N_4004);
nand U5931 (N_5931,N_4922,N_4285);
or U5932 (N_5932,N_4544,N_4723);
and U5933 (N_5933,N_4228,N_4512);
and U5934 (N_5934,N_4078,N_4833);
xor U5935 (N_5935,N_4128,N_4141);
and U5936 (N_5936,N_4035,N_4859);
and U5937 (N_5937,N_4986,N_4712);
and U5938 (N_5938,N_4823,N_4564);
and U5939 (N_5939,N_4967,N_4089);
xnor U5940 (N_5940,N_4419,N_4712);
or U5941 (N_5941,N_4088,N_4526);
nor U5942 (N_5942,N_4700,N_4380);
nand U5943 (N_5943,N_4862,N_4808);
nor U5944 (N_5944,N_4456,N_4754);
or U5945 (N_5945,N_4043,N_4550);
or U5946 (N_5946,N_4959,N_4377);
and U5947 (N_5947,N_4581,N_4967);
or U5948 (N_5948,N_4141,N_4435);
or U5949 (N_5949,N_4168,N_4824);
or U5950 (N_5950,N_4040,N_4261);
nand U5951 (N_5951,N_4334,N_4554);
and U5952 (N_5952,N_4065,N_4969);
and U5953 (N_5953,N_4618,N_4563);
and U5954 (N_5954,N_4469,N_4098);
or U5955 (N_5955,N_4595,N_4544);
and U5956 (N_5956,N_4939,N_4274);
nand U5957 (N_5957,N_4245,N_4768);
xnor U5958 (N_5958,N_4907,N_4182);
and U5959 (N_5959,N_4928,N_4507);
xor U5960 (N_5960,N_4758,N_4020);
and U5961 (N_5961,N_4934,N_4985);
or U5962 (N_5962,N_4129,N_4554);
nand U5963 (N_5963,N_4129,N_4832);
nor U5964 (N_5964,N_4525,N_4908);
and U5965 (N_5965,N_4711,N_4822);
and U5966 (N_5966,N_4142,N_4275);
xor U5967 (N_5967,N_4128,N_4680);
nand U5968 (N_5968,N_4791,N_4516);
nand U5969 (N_5969,N_4211,N_4432);
xor U5970 (N_5970,N_4112,N_4637);
and U5971 (N_5971,N_4734,N_4916);
nor U5972 (N_5972,N_4345,N_4494);
or U5973 (N_5973,N_4090,N_4831);
xor U5974 (N_5974,N_4564,N_4292);
xnor U5975 (N_5975,N_4018,N_4637);
nor U5976 (N_5976,N_4741,N_4963);
and U5977 (N_5977,N_4160,N_4916);
xor U5978 (N_5978,N_4861,N_4087);
or U5979 (N_5979,N_4186,N_4109);
nand U5980 (N_5980,N_4697,N_4987);
xor U5981 (N_5981,N_4716,N_4034);
nand U5982 (N_5982,N_4114,N_4935);
nand U5983 (N_5983,N_4869,N_4971);
and U5984 (N_5984,N_4942,N_4109);
xor U5985 (N_5985,N_4513,N_4180);
xnor U5986 (N_5986,N_4035,N_4549);
xor U5987 (N_5987,N_4659,N_4178);
xor U5988 (N_5988,N_4400,N_4822);
and U5989 (N_5989,N_4727,N_4968);
nor U5990 (N_5990,N_4384,N_4262);
nand U5991 (N_5991,N_4080,N_4194);
or U5992 (N_5992,N_4024,N_4826);
and U5993 (N_5993,N_4814,N_4977);
or U5994 (N_5994,N_4668,N_4990);
or U5995 (N_5995,N_4785,N_4401);
or U5996 (N_5996,N_4772,N_4477);
nand U5997 (N_5997,N_4840,N_4995);
nand U5998 (N_5998,N_4944,N_4900);
and U5999 (N_5999,N_4417,N_4870);
xnor U6000 (N_6000,N_5895,N_5846);
nor U6001 (N_6001,N_5556,N_5486);
nor U6002 (N_6002,N_5521,N_5044);
and U6003 (N_6003,N_5661,N_5926);
xnor U6004 (N_6004,N_5387,N_5997);
nor U6005 (N_6005,N_5698,N_5314);
or U6006 (N_6006,N_5467,N_5214);
nor U6007 (N_6007,N_5810,N_5254);
or U6008 (N_6008,N_5774,N_5751);
nor U6009 (N_6009,N_5909,N_5550);
or U6010 (N_6010,N_5931,N_5206);
nor U6011 (N_6011,N_5872,N_5617);
or U6012 (N_6012,N_5109,N_5445);
or U6013 (N_6013,N_5442,N_5938);
or U6014 (N_6014,N_5527,N_5407);
nand U6015 (N_6015,N_5058,N_5220);
nor U6016 (N_6016,N_5136,N_5611);
nand U6017 (N_6017,N_5284,N_5596);
nor U6018 (N_6018,N_5197,N_5885);
nor U6019 (N_6019,N_5838,N_5686);
or U6020 (N_6020,N_5884,N_5719);
nor U6021 (N_6021,N_5945,N_5697);
or U6022 (N_6022,N_5340,N_5615);
or U6023 (N_6023,N_5776,N_5302);
nor U6024 (N_6024,N_5976,N_5180);
and U6025 (N_6025,N_5127,N_5813);
nor U6026 (N_6026,N_5273,N_5770);
nor U6027 (N_6027,N_5444,N_5033);
or U6028 (N_6028,N_5419,N_5211);
xor U6029 (N_6029,N_5785,N_5979);
and U6030 (N_6030,N_5786,N_5683);
xnor U6031 (N_6031,N_5417,N_5173);
nor U6032 (N_6032,N_5261,N_5236);
and U6033 (N_6033,N_5218,N_5692);
xor U6034 (N_6034,N_5803,N_5944);
and U6035 (N_6035,N_5122,N_5729);
nand U6036 (N_6036,N_5981,N_5231);
or U6037 (N_6037,N_5753,N_5565);
xnor U6038 (N_6038,N_5933,N_5608);
nor U6039 (N_6039,N_5539,N_5124);
xor U6040 (N_6040,N_5987,N_5942);
nor U6041 (N_6041,N_5735,N_5963);
and U6042 (N_6042,N_5098,N_5577);
nor U6043 (N_6043,N_5534,N_5061);
nor U6044 (N_6044,N_5456,N_5282);
nor U6045 (N_6045,N_5506,N_5923);
or U6046 (N_6046,N_5269,N_5916);
nand U6047 (N_6047,N_5425,N_5102);
or U6048 (N_6048,N_5929,N_5319);
nor U6049 (N_6049,N_5087,N_5907);
and U6050 (N_6050,N_5429,N_5154);
or U6051 (N_6051,N_5705,N_5734);
nand U6052 (N_6052,N_5537,N_5393);
nand U6053 (N_6053,N_5966,N_5941);
nand U6054 (N_6054,N_5754,N_5675);
or U6055 (N_6055,N_5679,N_5263);
xor U6056 (N_6056,N_5583,N_5247);
nand U6057 (N_6057,N_5993,N_5003);
nor U6058 (N_6058,N_5581,N_5355);
or U6059 (N_6059,N_5213,N_5348);
xnor U6060 (N_6060,N_5050,N_5170);
xnor U6061 (N_6061,N_5439,N_5210);
nor U6062 (N_6062,N_5175,N_5833);
xor U6063 (N_6063,N_5763,N_5051);
xor U6064 (N_6064,N_5742,N_5094);
or U6065 (N_6065,N_5315,N_5322);
or U6066 (N_6066,N_5317,N_5682);
xor U6067 (N_6067,N_5318,N_5092);
nor U6068 (N_6068,N_5112,N_5497);
nor U6069 (N_6069,N_5186,N_5009);
nand U6070 (N_6070,N_5202,N_5538);
xnor U6071 (N_6071,N_5825,N_5347);
nand U6072 (N_6072,N_5835,N_5890);
nor U6073 (N_6073,N_5925,N_5164);
or U6074 (N_6074,N_5035,N_5715);
or U6075 (N_6075,N_5612,N_5396);
xor U6076 (N_6076,N_5081,N_5181);
xnor U6077 (N_6077,N_5519,N_5666);
xor U6078 (N_6078,N_5057,N_5755);
nand U6079 (N_6079,N_5491,N_5409);
nor U6080 (N_6080,N_5034,N_5451);
xor U6081 (N_6081,N_5352,N_5073);
and U6082 (N_6082,N_5485,N_5333);
or U6083 (N_6083,N_5784,N_5634);
and U6084 (N_6084,N_5054,N_5182);
xor U6085 (N_6085,N_5310,N_5790);
and U6086 (N_6086,N_5732,N_5921);
xnor U6087 (N_6087,N_5829,N_5176);
nor U6088 (N_6088,N_5511,N_5896);
xor U6089 (N_6089,N_5727,N_5305);
nand U6090 (N_6090,N_5541,N_5465);
nand U6091 (N_6091,N_5149,N_5660);
xnor U6092 (N_6092,N_5607,N_5168);
nor U6093 (N_6093,N_5240,N_5914);
xor U6094 (N_6094,N_5496,N_5591);
nand U6095 (N_6095,N_5723,N_5163);
and U6096 (N_6096,N_5398,N_5857);
nor U6097 (N_6097,N_5104,N_5958);
xor U6098 (N_6098,N_5466,N_5276);
xor U6099 (N_6099,N_5584,N_5039);
or U6100 (N_6100,N_5648,N_5426);
xnor U6101 (N_6101,N_5069,N_5851);
xor U6102 (N_6102,N_5649,N_5593);
nand U6103 (N_6103,N_5960,N_5128);
nand U6104 (N_6104,N_5381,N_5939);
nor U6105 (N_6105,N_5085,N_5971);
nor U6106 (N_6106,N_5344,N_5244);
xnor U6107 (N_6107,N_5821,N_5133);
nand U6108 (N_6108,N_5817,N_5903);
nand U6109 (N_6109,N_5765,N_5811);
and U6110 (N_6110,N_5863,N_5476);
nor U6111 (N_6111,N_5684,N_5889);
or U6112 (N_6112,N_5870,N_5038);
and U6113 (N_6113,N_5015,N_5222);
and U6114 (N_6114,N_5190,N_5516);
nor U6115 (N_6115,N_5056,N_5037);
and U6116 (N_6116,N_5695,N_5012);
nor U6117 (N_6117,N_5594,N_5329);
nor U6118 (N_6118,N_5200,N_5052);
nand U6119 (N_6119,N_5234,N_5001);
nand U6120 (N_6120,N_5191,N_5880);
nand U6121 (N_6121,N_5739,N_5948);
xnor U6122 (N_6122,N_5874,N_5303);
nand U6123 (N_6123,N_5005,N_5494);
nor U6124 (N_6124,N_5459,N_5716);
nand U6125 (N_6125,N_5915,N_5659);
xor U6126 (N_6126,N_5778,N_5865);
xor U6127 (N_6127,N_5363,N_5408);
nand U6128 (N_6128,N_5399,N_5287);
or U6129 (N_6129,N_5126,N_5826);
nor U6130 (N_6130,N_5858,N_5959);
xnor U6131 (N_6131,N_5510,N_5422);
or U6132 (N_6132,N_5132,N_5994);
nor U6133 (N_6133,N_5414,N_5225);
or U6134 (N_6134,N_5131,N_5194);
or U6135 (N_6135,N_5327,N_5654);
nor U6136 (N_6136,N_5328,N_5791);
xnor U6137 (N_6137,N_5193,N_5554);
nor U6138 (N_6138,N_5637,N_5837);
xnor U6139 (N_6139,N_5733,N_5908);
or U6140 (N_6140,N_5828,N_5843);
xnor U6141 (N_6141,N_5504,N_5088);
nor U6142 (N_6142,N_5452,N_5349);
and U6143 (N_6143,N_5571,N_5670);
nand U6144 (N_6144,N_5805,N_5120);
nor U6145 (N_6145,N_5443,N_5717);
or U6146 (N_6146,N_5326,N_5324);
or U6147 (N_6147,N_5954,N_5405);
or U6148 (N_6148,N_5397,N_5582);
xnor U6149 (N_6149,N_5892,N_5301);
nand U6150 (N_6150,N_5762,N_5410);
and U6151 (N_6151,N_5059,N_5802);
xor U6152 (N_6152,N_5421,N_5067);
nor U6153 (N_6153,N_5470,N_5157);
and U6154 (N_6154,N_5590,N_5226);
and U6155 (N_6155,N_5970,N_5990);
nand U6156 (N_6156,N_5553,N_5246);
nand U6157 (N_6157,N_5650,N_5949);
and U6158 (N_6158,N_5002,N_5080);
nand U6159 (N_6159,N_5882,N_5875);
xor U6160 (N_6160,N_5866,N_5557);
and U6161 (N_6161,N_5573,N_5713);
xor U6162 (N_6162,N_5325,N_5091);
or U6163 (N_6163,N_5824,N_5125);
or U6164 (N_6164,N_5711,N_5687);
and U6165 (N_6165,N_5673,N_5975);
xnor U6166 (N_6166,N_5106,N_5148);
or U6167 (N_6167,N_5464,N_5375);
nor U6168 (N_6168,N_5580,N_5576);
and U6169 (N_6169,N_5783,N_5512);
and U6170 (N_6170,N_5487,N_5374);
nor U6171 (N_6171,N_5313,N_5674);
xnor U6172 (N_6172,N_5855,N_5748);
nand U6173 (N_6173,N_5271,N_5701);
or U6174 (N_6174,N_5499,N_5007);
and U6175 (N_6175,N_5894,N_5691);
or U6176 (N_6176,N_5545,N_5049);
nor U6177 (N_6177,N_5587,N_5555);
or U6178 (N_6178,N_5390,N_5878);
nand U6179 (N_6179,N_5598,N_5747);
xnor U6180 (N_6180,N_5699,N_5888);
nand U6181 (N_6181,N_5201,N_5804);
and U6182 (N_6182,N_5588,N_5524);
nor U6183 (N_6183,N_5901,N_5657);
xor U6184 (N_6184,N_5841,N_5794);
or U6185 (N_6185,N_5710,N_5570);
nand U6186 (N_6186,N_5281,N_5533);
xor U6187 (N_6187,N_5529,N_5620);
and U6188 (N_6188,N_5307,N_5296);
and U6189 (N_6189,N_5740,N_5178);
and U6190 (N_6190,N_5292,N_5707);
or U6191 (N_6191,N_5101,N_5902);
xnor U6192 (N_6192,N_5083,N_5130);
or U6193 (N_6193,N_5071,N_5547);
nand U6194 (N_6194,N_5394,N_5940);
and U6195 (N_6195,N_5346,N_5469);
or U6196 (N_6196,N_5980,N_5066);
nand U6197 (N_6197,N_5773,N_5391);
nand U6198 (N_6198,N_5043,N_5230);
and U6199 (N_6199,N_5886,N_5638);
nor U6200 (N_6200,N_5946,N_5262);
or U6201 (N_6201,N_5165,N_5782);
and U6202 (N_6202,N_5664,N_5291);
nor U6203 (N_6203,N_5830,N_5455);
and U6204 (N_6204,N_5252,N_5256);
nand U6205 (N_6205,N_5517,N_5241);
nor U6206 (N_6206,N_5141,N_5248);
nor U6207 (N_6207,N_5224,N_5432);
xor U6208 (N_6208,N_5105,N_5074);
or U6209 (N_6209,N_5883,N_5392);
nand U6210 (N_6210,N_5653,N_5140);
nor U6211 (N_6211,N_5063,N_5046);
and U6212 (N_6212,N_5293,N_5471);
nor U6213 (N_6213,N_5192,N_5472);
nand U6214 (N_6214,N_5306,N_5336);
nand U6215 (N_6215,N_5227,N_5482);
nand U6216 (N_6216,N_5532,N_5750);
and U6217 (N_6217,N_5647,N_5635);
and U6218 (N_6218,N_5369,N_5280);
nor U6219 (N_6219,N_5977,N_5450);
and U6220 (N_6220,N_5599,N_5428);
xor U6221 (N_6221,N_5152,N_5366);
nor U6222 (N_6222,N_5278,N_5334);
and U6223 (N_6223,N_5943,N_5367);
and U6224 (N_6224,N_5379,N_5984);
xor U6225 (N_6225,N_5676,N_5242);
and U6226 (N_6226,N_5536,N_5503);
or U6227 (N_6227,N_5279,N_5730);
xnor U6228 (N_6228,N_5749,N_5481);
nand U6229 (N_6229,N_5458,N_5437);
xor U6230 (N_6230,N_5703,N_5669);
nor U6231 (N_6231,N_5245,N_5911);
and U6232 (N_6232,N_5642,N_5021);
or U6233 (N_6233,N_5509,N_5142);
nor U6234 (N_6234,N_5139,N_5010);
xnor U6235 (N_6235,N_5341,N_5042);
nor U6236 (N_6236,N_5989,N_5800);
xor U6237 (N_6237,N_5304,N_5289);
or U6238 (N_6238,N_5849,N_5853);
xor U6239 (N_6239,N_5361,N_5223);
and U6240 (N_6240,N_5834,N_5342);
or U6241 (N_6241,N_5400,N_5714);
xor U6242 (N_6242,N_5075,N_5771);
nand U6243 (N_6243,N_5881,N_5688);
nand U6244 (N_6244,N_5696,N_5619);
and U6245 (N_6245,N_5665,N_5431);
nand U6246 (N_6246,N_5077,N_5845);
or U6247 (N_6247,N_5277,N_5158);
and U6248 (N_6248,N_5160,N_5258);
and U6249 (N_6249,N_5370,N_5119);
and U6250 (N_6250,N_5718,N_5275);
xnor U6251 (N_6251,N_5685,N_5045);
xnor U6252 (N_6252,N_5973,N_5072);
nor U6253 (N_6253,N_5099,N_5060);
nand U6254 (N_6254,N_5483,N_5951);
or U6255 (N_6255,N_5053,N_5474);
xnor U6256 (N_6256,N_5298,N_5383);
nand U6257 (N_6257,N_5135,N_5871);
nand U6258 (N_6258,N_5016,N_5781);
nor U6259 (N_6259,N_5873,N_5462);
or U6260 (N_6260,N_5427,N_5253);
and U6261 (N_6261,N_5116,N_5836);
nand U6262 (N_6262,N_5952,N_5842);
and U6263 (N_6263,N_5048,N_5508);
nor U6264 (N_6264,N_5726,N_5779);
and U6265 (N_6265,N_5562,N_5420);
nand U6266 (N_6266,N_5531,N_5636);
and U6267 (N_6267,N_5295,N_5632);
xor U6268 (N_6268,N_5702,N_5115);
nor U6269 (N_6269,N_5025,N_5932);
or U6270 (N_6270,N_5887,N_5561);
and U6271 (N_6271,N_5799,N_5935);
or U6272 (N_6272,N_5910,N_5528);
nand U6273 (N_6273,N_5758,N_5772);
nand U6274 (N_6274,N_5460,N_5560);
xnor U6275 (N_6275,N_5377,N_5237);
nor U6276 (N_6276,N_5103,N_5195);
nor U6277 (N_6277,N_5618,N_5566);
and U6278 (N_6278,N_5530,N_5068);
nand U6279 (N_6279,N_5622,N_5725);
and U6280 (N_6280,N_5283,N_5546);
xnor U6281 (N_6281,N_5793,N_5600);
nand U6282 (N_6282,N_5548,N_5905);
and U6283 (N_6283,N_5693,N_5238);
and U6284 (N_6284,N_5756,N_5143);
and U6285 (N_6285,N_5655,N_5300);
nand U6286 (N_6286,N_5498,N_5264);
nand U6287 (N_6287,N_5609,N_5672);
or U6288 (N_6288,N_5578,N_5912);
and U6289 (N_6289,N_5311,N_5339);
xor U6290 (N_6290,N_5967,N_5720);
and U6291 (N_6291,N_5513,N_5917);
nand U6292 (N_6292,N_5449,N_5331);
or U6293 (N_6293,N_5257,N_5402);
and U6294 (N_6294,N_5171,N_5645);
nand U6295 (N_6295,N_5731,N_5024);
nand U6296 (N_6296,N_5757,N_5386);
xor U6297 (N_6297,N_5243,N_5436);
nor U6298 (N_6298,N_5475,N_5188);
nor U6299 (N_6299,N_5232,N_5898);
nand U6300 (N_6300,N_5368,N_5815);
or U6301 (N_6301,N_5639,N_5014);
xnor U6302 (N_6302,N_5123,N_5177);
and U6303 (N_6303,N_5026,N_5183);
nor U6304 (N_6304,N_5961,N_5265);
and U6305 (N_6305,N_5070,N_5076);
nor U6306 (N_6306,N_5543,N_5260);
nand U6307 (N_6307,N_5752,N_5614);
nor U6308 (N_6308,N_5797,N_5671);
and U6309 (N_6309,N_5274,N_5228);
nand U6310 (N_6310,N_5575,N_5505);
nand U6311 (N_6311,N_5928,N_5589);
or U6312 (N_6312,N_5924,N_5996);
and U6313 (N_6313,N_5216,N_5544);
nor U6314 (N_6314,N_5032,N_5096);
nor U6315 (N_6315,N_5864,N_5477);
nor U6316 (N_6316,N_5345,N_5934);
nor U6317 (N_6317,N_5623,N_5605);
nor U6318 (N_6318,N_5259,N_5029);
xnor U6319 (N_6319,N_5658,N_5041);
and U6320 (N_6320,N_5953,N_5854);
xor U6321 (N_6321,N_5272,N_5606);
or U6322 (N_6322,N_5167,N_5904);
and U6323 (N_6323,N_5415,N_5055);
nor U6324 (N_6324,N_5962,N_5767);
or U6325 (N_6325,N_5522,N_5964);
or U6326 (N_6326,N_5332,N_5484);
nand U6327 (N_6327,N_5205,N_5360);
nand U6328 (N_6328,N_5288,N_5930);
nor U6329 (N_6329,N_5356,N_5551);
or U6330 (N_6330,N_5988,N_5820);
nand U6331 (N_6331,N_5681,N_5919);
nor U6332 (N_6332,N_5113,N_5249);
nor U6333 (N_6333,N_5488,N_5891);
xnor U6334 (N_6334,N_5831,N_5760);
and U6335 (N_6335,N_5359,N_5769);
xnor U6336 (N_6336,N_5798,N_5019);
nand U6337 (N_6337,N_5184,N_5848);
nand U6338 (N_6338,N_5625,N_5114);
and U6339 (N_6339,N_5816,N_5983);
and U6340 (N_6340,N_5978,N_5108);
nand U6341 (N_6341,N_5229,N_5985);
nor U6342 (N_6342,N_5489,N_5761);
and U6343 (N_6343,N_5312,N_5385);
or U6344 (N_6344,N_5011,N_5166);
and U6345 (N_6345,N_5204,N_5362);
or U6346 (N_6346,N_5795,N_5473);
nor U6347 (N_6347,N_5198,N_5656);
nor U6348 (N_6348,N_5266,N_5100);
or U6349 (N_6349,N_5906,N_5233);
xnor U6350 (N_6350,N_5372,N_5937);
or U6351 (N_6351,N_5129,N_5780);
xor U6352 (N_6352,N_5461,N_5633);
nand U6353 (N_6353,N_5741,N_5823);
and U6354 (N_6354,N_5592,N_5086);
xnor U6355 (N_6355,N_5564,N_5540);
xor U6356 (N_6356,N_5239,N_5364);
or U6357 (N_6357,N_5006,N_5972);
and U6358 (N_6358,N_5089,N_5627);
xor U6359 (N_6359,N_5809,N_5646);
and U6360 (N_6360,N_5630,N_5084);
nor U6361 (N_6361,N_5376,N_5031);
xnor U6362 (N_6362,N_5955,N_5667);
xnor U6363 (N_6363,N_5861,N_5468);
or U6364 (N_6364,N_5255,N_5523);
xnor U6365 (N_6365,N_5365,N_5144);
nor U6366 (N_6366,N_5023,N_5968);
xor U6367 (N_6367,N_5913,N_5950);
xor U6368 (N_6368,N_5065,N_5172);
nand U6369 (N_6369,N_5117,N_5788);
nand U6370 (N_6370,N_5535,N_5169);
and U6371 (N_6371,N_5900,N_5185);
and U6372 (N_6372,N_5563,N_5179);
xor U6373 (N_6373,N_5789,N_5027);
nor U6374 (N_6374,N_5559,N_5212);
nor U6375 (N_6375,N_5722,N_5728);
nor U6376 (N_6376,N_5161,N_5738);
nor U6377 (N_6377,N_5013,N_5764);
nand U6378 (N_6378,N_5746,N_5744);
nor U6379 (N_6379,N_5777,N_5062);
xor U6380 (N_6380,N_5447,N_5500);
and U6381 (N_6381,N_5574,N_5680);
xor U6382 (N_6382,N_5207,N_5957);
nor U6383 (N_6383,N_5189,N_5330);
and U6384 (N_6384,N_5146,N_5004);
xnor U6385 (N_6385,N_5208,N_5268);
xor U6386 (N_6386,N_5640,N_5787);
and U6387 (N_6387,N_5595,N_5965);
nor U6388 (N_6388,N_5411,N_5601);
nand U6389 (N_6389,N_5812,N_5401);
and U6390 (N_6390,N_5706,N_5792);
or U6391 (N_6391,N_5852,N_5338);
nand U6392 (N_6392,N_5187,N_5867);
xnor U6393 (N_6393,N_5663,N_5585);
nand U6394 (N_6394,N_5737,N_5478);
nand U6395 (N_6395,N_5251,N_5579);
nand U6396 (N_6396,N_5353,N_5371);
nand U6397 (N_6397,N_5412,N_5947);
and U6398 (N_6398,N_5388,N_5413);
xor U6399 (N_6399,N_5441,N_5424);
and U6400 (N_6400,N_5221,N_5991);
nand U6401 (N_6401,N_5927,N_5479);
and U6402 (N_6402,N_5869,N_5626);
or U6403 (N_6403,N_5350,N_5678);
and U6404 (N_6404,N_5203,N_5294);
nor U6405 (N_6405,N_5597,N_5982);
or U6406 (N_6406,N_5631,N_5712);
nand U6407 (N_6407,N_5518,N_5378);
and U6408 (N_6408,N_5406,N_5807);
nand U6409 (N_6409,N_5416,N_5299);
or U6410 (N_6410,N_5520,N_5453);
nand U6411 (N_6411,N_5549,N_5270);
xnor U6412 (N_6412,N_5433,N_5724);
nand U6413 (N_6413,N_5602,N_5613);
nor U6414 (N_6414,N_5492,N_5457);
nor U6415 (N_6415,N_5111,N_5490);
nor U6416 (N_6416,N_5876,N_5986);
xor U6417 (N_6417,N_5309,N_5709);
nand U6418 (N_6418,N_5493,N_5155);
nor U6419 (N_6419,N_5999,N_5423);
nand U6420 (N_6420,N_5859,N_5542);
or U6421 (N_6421,N_5879,N_5357);
and U6422 (N_6422,N_5215,N_5047);
and U6423 (N_6423,N_5604,N_5616);
nor U6424 (N_6424,N_5078,N_5028);
xnor U6425 (N_6425,N_5651,N_5569);
nor U6426 (N_6426,N_5862,N_5819);
xnor U6427 (N_6427,N_5138,N_5775);
nand U6428 (N_6428,N_5877,N_5847);
nand U6429 (N_6429,N_5150,N_5286);
xnor U6430 (N_6430,N_5093,N_5694);
nor U6431 (N_6431,N_5335,N_5480);
xor U6432 (N_6432,N_5082,N_5384);
and U6433 (N_6433,N_5174,N_5463);
xnor U6434 (N_6434,N_5404,N_5844);
or U6435 (N_6435,N_5354,N_5525);
and U6436 (N_6436,N_5814,N_5118);
nand U6437 (N_6437,N_5822,N_5893);
xnor U6438 (N_6438,N_5389,N_5801);
xnor U6439 (N_6439,N_5808,N_5868);
nand U6440 (N_6440,N_5438,N_5850);
and U6441 (N_6441,N_5358,N_5121);
nor U6442 (N_6442,N_5316,N_5827);
and U6443 (N_6443,N_5700,N_5454);
and U6444 (N_6444,N_5250,N_5022);
xnor U6445 (N_6445,N_5156,N_5107);
or U6446 (N_6446,N_5162,N_5759);
nand U6447 (N_6447,N_5558,N_5514);
and U6448 (N_6448,N_5662,N_5323);
nand U6449 (N_6449,N_5677,N_5403);
nor U6450 (N_6450,N_5736,N_5690);
or U6451 (N_6451,N_5017,N_5818);
or U6452 (N_6452,N_5796,N_5446);
nand U6453 (N_6453,N_5382,N_5217);
or U6454 (N_6454,N_5806,N_5766);
xor U6455 (N_6455,N_5064,N_5992);
and U6456 (N_6456,N_5153,N_5643);
or U6457 (N_6457,N_5095,N_5147);
and U6458 (N_6458,N_5434,N_5721);
and U6459 (N_6459,N_5918,N_5308);
nor U6460 (N_6460,N_5418,N_5159);
and U6461 (N_6461,N_5936,N_5708);
xnor U6462 (N_6462,N_5145,N_5235);
or U6463 (N_6463,N_5448,N_5008);
nor U6464 (N_6464,N_5267,N_5219);
nand U6465 (N_6465,N_5285,N_5297);
nand U6466 (N_6466,N_5768,N_5343);
xor U6467 (N_6467,N_5652,N_5290);
xnor U6468 (N_6468,N_5196,N_5097);
or U6469 (N_6469,N_5974,N_5897);
xor U6470 (N_6470,N_5495,N_5743);
and U6471 (N_6471,N_5832,N_5586);
nor U6472 (N_6472,N_5572,N_5840);
nand U6473 (N_6473,N_5199,N_5137);
nor U6474 (N_6474,N_5502,N_5430);
and U6475 (N_6475,N_5079,N_5320);
xor U6476 (N_6476,N_5969,N_5040);
nor U6477 (N_6477,N_5603,N_5435);
nand U6478 (N_6478,N_5020,N_5624);
nand U6479 (N_6479,N_5380,N_5110);
and U6480 (N_6480,N_5860,N_5956);
and U6481 (N_6481,N_5018,N_5526);
and U6482 (N_6482,N_5641,N_5628);
and U6483 (N_6483,N_5515,N_5995);
and U6484 (N_6484,N_5030,N_5610);
nor U6485 (N_6485,N_5899,N_5507);
nor U6486 (N_6486,N_5567,N_5440);
or U6487 (N_6487,N_5209,N_5704);
nand U6488 (N_6488,N_5036,N_5000);
xor U6489 (N_6489,N_5151,N_5668);
nand U6490 (N_6490,N_5337,N_5373);
nor U6491 (N_6491,N_5644,N_5090);
nand U6492 (N_6492,N_5621,N_5552);
xor U6493 (N_6493,N_5689,N_5922);
and U6494 (N_6494,N_5321,N_5856);
xor U6495 (N_6495,N_5920,N_5568);
nand U6496 (N_6496,N_5501,N_5134);
or U6497 (N_6497,N_5395,N_5745);
and U6498 (N_6498,N_5351,N_5629);
nor U6499 (N_6499,N_5839,N_5998);
or U6500 (N_6500,N_5721,N_5260);
and U6501 (N_6501,N_5592,N_5806);
nand U6502 (N_6502,N_5716,N_5257);
nor U6503 (N_6503,N_5503,N_5542);
nor U6504 (N_6504,N_5265,N_5010);
nor U6505 (N_6505,N_5826,N_5472);
nand U6506 (N_6506,N_5564,N_5095);
nand U6507 (N_6507,N_5128,N_5434);
or U6508 (N_6508,N_5084,N_5553);
and U6509 (N_6509,N_5215,N_5233);
or U6510 (N_6510,N_5835,N_5671);
xor U6511 (N_6511,N_5360,N_5544);
xnor U6512 (N_6512,N_5582,N_5836);
xnor U6513 (N_6513,N_5141,N_5936);
nor U6514 (N_6514,N_5489,N_5600);
xor U6515 (N_6515,N_5068,N_5602);
nand U6516 (N_6516,N_5845,N_5473);
nand U6517 (N_6517,N_5095,N_5072);
nor U6518 (N_6518,N_5240,N_5869);
nor U6519 (N_6519,N_5248,N_5161);
and U6520 (N_6520,N_5261,N_5785);
nor U6521 (N_6521,N_5689,N_5496);
or U6522 (N_6522,N_5957,N_5829);
nand U6523 (N_6523,N_5859,N_5246);
and U6524 (N_6524,N_5965,N_5760);
and U6525 (N_6525,N_5964,N_5182);
or U6526 (N_6526,N_5670,N_5067);
and U6527 (N_6527,N_5222,N_5284);
nor U6528 (N_6528,N_5992,N_5689);
and U6529 (N_6529,N_5567,N_5934);
nand U6530 (N_6530,N_5127,N_5964);
xnor U6531 (N_6531,N_5601,N_5522);
nor U6532 (N_6532,N_5457,N_5237);
and U6533 (N_6533,N_5030,N_5393);
or U6534 (N_6534,N_5227,N_5656);
and U6535 (N_6535,N_5334,N_5837);
and U6536 (N_6536,N_5979,N_5802);
nand U6537 (N_6537,N_5795,N_5998);
or U6538 (N_6538,N_5666,N_5155);
nand U6539 (N_6539,N_5071,N_5290);
or U6540 (N_6540,N_5892,N_5123);
nand U6541 (N_6541,N_5284,N_5534);
nand U6542 (N_6542,N_5844,N_5815);
xor U6543 (N_6543,N_5916,N_5308);
nor U6544 (N_6544,N_5189,N_5412);
and U6545 (N_6545,N_5291,N_5411);
nand U6546 (N_6546,N_5700,N_5198);
nor U6547 (N_6547,N_5537,N_5283);
nor U6548 (N_6548,N_5589,N_5324);
nand U6549 (N_6549,N_5065,N_5073);
or U6550 (N_6550,N_5752,N_5162);
nor U6551 (N_6551,N_5123,N_5115);
xor U6552 (N_6552,N_5667,N_5933);
nand U6553 (N_6553,N_5331,N_5427);
xnor U6554 (N_6554,N_5947,N_5384);
and U6555 (N_6555,N_5228,N_5602);
nor U6556 (N_6556,N_5207,N_5149);
xnor U6557 (N_6557,N_5919,N_5455);
xnor U6558 (N_6558,N_5111,N_5892);
nor U6559 (N_6559,N_5025,N_5066);
nor U6560 (N_6560,N_5835,N_5263);
xnor U6561 (N_6561,N_5175,N_5529);
nor U6562 (N_6562,N_5867,N_5502);
nand U6563 (N_6563,N_5104,N_5258);
nor U6564 (N_6564,N_5302,N_5495);
nor U6565 (N_6565,N_5210,N_5396);
nand U6566 (N_6566,N_5215,N_5309);
and U6567 (N_6567,N_5248,N_5881);
and U6568 (N_6568,N_5768,N_5874);
nor U6569 (N_6569,N_5675,N_5204);
nor U6570 (N_6570,N_5923,N_5312);
or U6571 (N_6571,N_5421,N_5737);
and U6572 (N_6572,N_5920,N_5531);
nand U6573 (N_6573,N_5176,N_5972);
and U6574 (N_6574,N_5340,N_5803);
and U6575 (N_6575,N_5507,N_5940);
or U6576 (N_6576,N_5291,N_5105);
or U6577 (N_6577,N_5442,N_5137);
nand U6578 (N_6578,N_5051,N_5296);
nand U6579 (N_6579,N_5346,N_5516);
nand U6580 (N_6580,N_5486,N_5899);
nand U6581 (N_6581,N_5866,N_5602);
xor U6582 (N_6582,N_5859,N_5871);
nand U6583 (N_6583,N_5103,N_5353);
nand U6584 (N_6584,N_5168,N_5029);
xnor U6585 (N_6585,N_5070,N_5944);
nand U6586 (N_6586,N_5440,N_5667);
xnor U6587 (N_6587,N_5370,N_5574);
nor U6588 (N_6588,N_5973,N_5954);
xor U6589 (N_6589,N_5420,N_5132);
nand U6590 (N_6590,N_5699,N_5505);
and U6591 (N_6591,N_5222,N_5902);
or U6592 (N_6592,N_5677,N_5376);
and U6593 (N_6593,N_5035,N_5439);
and U6594 (N_6594,N_5518,N_5388);
nand U6595 (N_6595,N_5669,N_5817);
xnor U6596 (N_6596,N_5553,N_5817);
nor U6597 (N_6597,N_5823,N_5829);
nand U6598 (N_6598,N_5561,N_5664);
xnor U6599 (N_6599,N_5470,N_5739);
nor U6600 (N_6600,N_5443,N_5092);
or U6601 (N_6601,N_5662,N_5774);
nand U6602 (N_6602,N_5394,N_5398);
or U6603 (N_6603,N_5612,N_5784);
or U6604 (N_6604,N_5507,N_5602);
xor U6605 (N_6605,N_5367,N_5910);
nor U6606 (N_6606,N_5437,N_5227);
xor U6607 (N_6607,N_5317,N_5769);
and U6608 (N_6608,N_5643,N_5299);
and U6609 (N_6609,N_5473,N_5829);
and U6610 (N_6610,N_5353,N_5519);
nor U6611 (N_6611,N_5169,N_5247);
and U6612 (N_6612,N_5458,N_5410);
and U6613 (N_6613,N_5553,N_5996);
nor U6614 (N_6614,N_5654,N_5291);
and U6615 (N_6615,N_5957,N_5171);
or U6616 (N_6616,N_5022,N_5787);
nand U6617 (N_6617,N_5496,N_5983);
or U6618 (N_6618,N_5774,N_5564);
or U6619 (N_6619,N_5270,N_5796);
or U6620 (N_6620,N_5626,N_5098);
nor U6621 (N_6621,N_5605,N_5359);
and U6622 (N_6622,N_5736,N_5838);
or U6623 (N_6623,N_5012,N_5378);
xnor U6624 (N_6624,N_5185,N_5091);
or U6625 (N_6625,N_5882,N_5907);
nor U6626 (N_6626,N_5122,N_5164);
nand U6627 (N_6627,N_5521,N_5010);
nor U6628 (N_6628,N_5442,N_5177);
nor U6629 (N_6629,N_5423,N_5178);
xor U6630 (N_6630,N_5727,N_5314);
xor U6631 (N_6631,N_5459,N_5036);
and U6632 (N_6632,N_5241,N_5744);
or U6633 (N_6633,N_5197,N_5695);
nand U6634 (N_6634,N_5799,N_5603);
and U6635 (N_6635,N_5880,N_5754);
and U6636 (N_6636,N_5707,N_5071);
or U6637 (N_6637,N_5726,N_5934);
nand U6638 (N_6638,N_5082,N_5938);
nor U6639 (N_6639,N_5901,N_5094);
nor U6640 (N_6640,N_5222,N_5349);
and U6641 (N_6641,N_5041,N_5880);
nand U6642 (N_6642,N_5355,N_5419);
or U6643 (N_6643,N_5173,N_5992);
or U6644 (N_6644,N_5527,N_5226);
nand U6645 (N_6645,N_5287,N_5469);
or U6646 (N_6646,N_5087,N_5118);
and U6647 (N_6647,N_5860,N_5510);
xor U6648 (N_6648,N_5810,N_5890);
nor U6649 (N_6649,N_5446,N_5875);
nor U6650 (N_6650,N_5964,N_5172);
and U6651 (N_6651,N_5144,N_5069);
xnor U6652 (N_6652,N_5479,N_5417);
or U6653 (N_6653,N_5852,N_5210);
xnor U6654 (N_6654,N_5619,N_5090);
and U6655 (N_6655,N_5697,N_5696);
or U6656 (N_6656,N_5650,N_5769);
nand U6657 (N_6657,N_5607,N_5944);
and U6658 (N_6658,N_5315,N_5587);
xnor U6659 (N_6659,N_5031,N_5853);
nor U6660 (N_6660,N_5069,N_5624);
xnor U6661 (N_6661,N_5464,N_5158);
xnor U6662 (N_6662,N_5012,N_5271);
and U6663 (N_6663,N_5988,N_5812);
or U6664 (N_6664,N_5099,N_5245);
nor U6665 (N_6665,N_5229,N_5659);
nor U6666 (N_6666,N_5192,N_5575);
or U6667 (N_6667,N_5444,N_5293);
nand U6668 (N_6668,N_5738,N_5974);
or U6669 (N_6669,N_5884,N_5872);
and U6670 (N_6670,N_5809,N_5656);
or U6671 (N_6671,N_5604,N_5244);
nand U6672 (N_6672,N_5343,N_5340);
or U6673 (N_6673,N_5127,N_5675);
and U6674 (N_6674,N_5493,N_5118);
and U6675 (N_6675,N_5519,N_5981);
nor U6676 (N_6676,N_5478,N_5536);
or U6677 (N_6677,N_5523,N_5842);
or U6678 (N_6678,N_5285,N_5907);
xnor U6679 (N_6679,N_5943,N_5656);
nand U6680 (N_6680,N_5082,N_5826);
nand U6681 (N_6681,N_5689,N_5618);
or U6682 (N_6682,N_5044,N_5863);
and U6683 (N_6683,N_5207,N_5141);
nor U6684 (N_6684,N_5496,N_5185);
nand U6685 (N_6685,N_5930,N_5136);
xnor U6686 (N_6686,N_5746,N_5335);
and U6687 (N_6687,N_5142,N_5654);
xnor U6688 (N_6688,N_5625,N_5622);
or U6689 (N_6689,N_5216,N_5792);
nand U6690 (N_6690,N_5368,N_5571);
nor U6691 (N_6691,N_5295,N_5435);
xnor U6692 (N_6692,N_5463,N_5172);
nand U6693 (N_6693,N_5272,N_5128);
xor U6694 (N_6694,N_5504,N_5212);
xor U6695 (N_6695,N_5656,N_5440);
nor U6696 (N_6696,N_5200,N_5886);
nor U6697 (N_6697,N_5867,N_5604);
nand U6698 (N_6698,N_5310,N_5877);
xnor U6699 (N_6699,N_5045,N_5605);
nand U6700 (N_6700,N_5239,N_5837);
xnor U6701 (N_6701,N_5684,N_5371);
or U6702 (N_6702,N_5806,N_5469);
nor U6703 (N_6703,N_5790,N_5804);
and U6704 (N_6704,N_5201,N_5189);
nand U6705 (N_6705,N_5827,N_5603);
or U6706 (N_6706,N_5311,N_5609);
nand U6707 (N_6707,N_5486,N_5629);
and U6708 (N_6708,N_5163,N_5298);
xor U6709 (N_6709,N_5121,N_5583);
xor U6710 (N_6710,N_5742,N_5312);
nor U6711 (N_6711,N_5353,N_5113);
nor U6712 (N_6712,N_5727,N_5687);
or U6713 (N_6713,N_5323,N_5558);
and U6714 (N_6714,N_5989,N_5941);
and U6715 (N_6715,N_5013,N_5515);
and U6716 (N_6716,N_5404,N_5132);
xor U6717 (N_6717,N_5557,N_5656);
nor U6718 (N_6718,N_5568,N_5616);
xor U6719 (N_6719,N_5219,N_5200);
and U6720 (N_6720,N_5738,N_5570);
or U6721 (N_6721,N_5430,N_5927);
xor U6722 (N_6722,N_5214,N_5356);
nand U6723 (N_6723,N_5321,N_5445);
nand U6724 (N_6724,N_5884,N_5689);
nor U6725 (N_6725,N_5957,N_5096);
or U6726 (N_6726,N_5883,N_5559);
or U6727 (N_6727,N_5067,N_5974);
and U6728 (N_6728,N_5932,N_5198);
nand U6729 (N_6729,N_5838,N_5121);
xnor U6730 (N_6730,N_5503,N_5022);
nand U6731 (N_6731,N_5560,N_5656);
nor U6732 (N_6732,N_5259,N_5158);
xor U6733 (N_6733,N_5623,N_5632);
xnor U6734 (N_6734,N_5491,N_5213);
xnor U6735 (N_6735,N_5162,N_5192);
nor U6736 (N_6736,N_5259,N_5361);
xnor U6737 (N_6737,N_5024,N_5877);
nand U6738 (N_6738,N_5902,N_5714);
nor U6739 (N_6739,N_5386,N_5985);
nor U6740 (N_6740,N_5197,N_5723);
or U6741 (N_6741,N_5014,N_5655);
and U6742 (N_6742,N_5380,N_5104);
nand U6743 (N_6743,N_5677,N_5028);
or U6744 (N_6744,N_5494,N_5487);
and U6745 (N_6745,N_5850,N_5786);
nor U6746 (N_6746,N_5673,N_5388);
and U6747 (N_6747,N_5832,N_5654);
nand U6748 (N_6748,N_5939,N_5559);
nor U6749 (N_6749,N_5058,N_5413);
nor U6750 (N_6750,N_5425,N_5312);
or U6751 (N_6751,N_5629,N_5125);
nand U6752 (N_6752,N_5690,N_5373);
nand U6753 (N_6753,N_5854,N_5304);
nor U6754 (N_6754,N_5799,N_5428);
nor U6755 (N_6755,N_5668,N_5078);
and U6756 (N_6756,N_5512,N_5191);
and U6757 (N_6757,N_5727,N_5379);
and U6758 (N_6758,N_5556,N_5855);
and U6759 (N_6759,N_5438,N_5842);
nor U6760 (N_6760,N_5264,N_5688);
xnor U6761 (N_6761,N_5524,N_5804);
nor U6762 (N_6762,N_5455,N_5367);
and U6763 (N_6763,N_5237,N_5328);
nor U6764 (N_6764,N_5610,N_5700);
or U6765 (N_6765,N_5328,N_5496);
or U6766 (N_6766,N_5887,N_5545);
nor U6767 (N_6767,N_5852,N_5665);
or U6768 (N_6768,N_5570,N_5019);
and U6769 (N_6769,N_5679,N_5278);
or U6770 (N_6770,N_5695,N_5156);
nand U6771 (N_6771,N_5945,N_5065);
nor U6772 (N_6772,N_5425,N_5599);
nand U6773 (N_6773,N_5911,N_5475);
and U6774 (N_6774,N_5287,N_5477);
nand U6775 (N_6775,N_5587,N_5524);
xor U6776 (N_6776,N_5960,N_5468);
xnor U6777 (N_6777,N_5200,N_5120);
xor U6778 (N_6778,N_5417,N_5281);
nor U6779 (N_6779,N_5892,N_5677);
or U6780 (N_6780,N_5139,N_5599);
xnor U6781 (N_6781,N_5718,N_5790);
and U6782 (N_6782,N_5225,N_5550);
and U6783 (N_6783,N_5837,N_5058);
nand U6784 (N_6784,N_5195,N_5041);
nor U6785 (N_6785,N_5417,N_5312);
or U6786 (N_6786,N_5804,N_5982);
nor U6787 (N_6787,N_5315,N_5894);
nor U6788 (N_6788,N_5045,N_5757);
nand U6789 (N_6789,N_5788,N_5341);
and U6790 (N_6790,N_5157,N_5174);
nor U6791 (N_6791,N_5382,N_5618);
or U6792 (N_6792,N_5403,N_5852);
nand U6793 (N_6793,N_5914,N_5569);
nor U6794 (N_6794,N_5595,N_5416);
nor U6795 (N_6795,N_5584,N_5031);
or U6796 (N_6796,N_5628,N_5929);
and U6797 (N_6797,N_5614,N_5318);
and U6798 (N_6798,N_5052,N_5145);
nand U6799 (N_6799,N_5984,N_5497);
xnor U6800 (N_6800,N_5972,N_5054);
or U6801 (N_6801,N_5894,N_5926);
xnor U6802 (N_6802,N_5041,N_5290);
xor U6803 (N_6803,N_5071,N_5987);
xnor U6804 (N_6804,N_5807,N_5051);
nor U6805 (N_6805,N_5946,N_5876);
nor U6806 (N_6806,N_5732,N_5987);
xor U6807 (N_6807,N_5419,N_5676);
nor U6808 (N_6808,N_5996,N_5192);
nand U6809 (N_6809,N_5057,N_5514);
and U6810 (N_6810,N_5535,N_5628);
xor U6811 (N_6811,N_5133,N_5086);
or U6812 (N_6812,N_5635,N_5257);
xnor U6813 (N_6813,N_5219,N_5077);
nand U6814 (N_6814,N_5343,N_5140);
nand U6815 (N_6815,N_5143,N_5952);
or U6816 (N_6816,N_5932,N_5118);
and U6817 (N_6817,N_5894,N_5445);
xor U6818 (N_6818,N_5937,N_5553);
nor U6819 (N_6819,N_5149,N_5599);
or U6820 (N_6820,N_5837,N_5179);
and U6821 (N_6821,N_5611,N_5398);
nand U6822 (N_6822,N_5281,N_5678);
nor U6823 (N_6823,N_5019,N_5281);
xnor U6824 (N_6824,N_5063,N_5039);
nor U6825 (N_6825,N_5702,N_5899);
nor U6826 (N_6826,N_5528,N_5392);
or U6827 (N_6827,N_5595,N_5898);
nor U6828 (N_6828,N_5548,N_5168);
and U6829 (N_6829,N_5558,N_5145);
xor U6830 (N_6830,N_5630,N_5892);
or U6831 (N_6831,N_5439,N_5693);
nor U6832 (N_6832,N_5749,N_5338);
nor U6833 (N_6833,N_5055,N_5407);
or U6834 (N_6834,N_5730,N_5406);
nor U6835 (N_6835,N_5603,N_5727);
or U6836 (N_6836,N_5967,N_5435);
and U6837 (N_6837,N_5860,N_5889);
and U6838 (N_6838,N_5009,N_5755);
or U6839 (N_6839,N_5912,N_5308);
and U6840 (N_6840,N_5151,N_5366);
xnor U6841 (N_6841,N_5559,N_5619);
nand U6842 (N_6842,N_5403,N_5860);
xnor U6843 (N_6843,N_5944,N_5498);
nand U6844 (N_6844,N_5349,N_5403);
nor U6845 (N_6845,N_5940,N_5335);
nor U6846 (N_6846,N_5748,N_5142);
nor U6847 (N_6847,N_5016,N_5473);
xor U6848 (N_6848,N_5357,N_5334);
nor U6849 (N_6849,N_5653,N_5069);
nor U6850 (N_6850,N_5261,N_5166);
nand U6851 (N_6851,N_5189,N_5453);
nand U6852 (N_6852,N_5812,N_5231);
xor U6853 (N_6853,N_5421,N_5131);
and U6854 (N_6854,N_5189,N_5707);
and U6855 (N_6855,N_5237,N_5441);
nand U6856 (N_6856,N_5955,N_5152);
and U6857 (N_6857,N_5889,N_5563);
or U6858 (N_6858,N_5904,N_5092);
xnor U6859 (N_6859,N_5206,N_5827);
and U6860 (N_6860,N_5612,N_5628);
xnor U6861 (N_6861,N_5175,N_5407);
or U6862 (N_6862,N_5036,N_5336);
nor U6863 (N_6863,N_5707,N_5924);
xor U6864 (N_6864,N_5140,N_5017);
or U6865 (N_6865,N_5267,N_5402);
nor U6866 (N_6866,N_5765,N_5541);
or U6867 (N_6867,N_5166,N_5141);
nand U6868 (N_6868,N_5385,N_5566);
nand U6869 (N_6869,N_5240,N_5482);
nor U6870 (N_6870,N_5315,N_5256);
or U6871 (N_6871,N_5827,N_5508);
nand U6872 (N_6872,N_5120,N_5922);
nor U6873 (N_6873,N_5600,N_5780);
and U6874 (N_6874,N_5706,N_5114);
and U6875 (N_6875,N_5818,N_5736);
nand U6876 (N_6876,N_5748,N_5226);
and U6877 (N_6877,N_5197,N_5593);
xor U6878 (N_6878,N_5164,N_5313);
or U6879 (N_6879,N_5662,N_5108);
and U6880 (N_6880,N_5296,N_5935);
or U6881 (N_6881,N_5640,N_5062);
nor U6882 (N_6882,N_5288,N_5016);
or U6883 (N_6883,N_5212,N_5409);
and U6884 (N_6884,N_5109,N_5176);
xnor U6885 (N_6885,N_5335,N_5100);
xnor U6886 (N_6886,N_5538,N_5227);
and U6887 (N_6887,N_5441,N_5337);
xnor U6888 (N_6888,N_5813,N_5872);
or U6889 (N_6889,N_5398,N_5228);
or U6890 (N_6890,N_5545,N_5557);
and U6891 (N_6891,N_5390,N_5267);
and U6892 (N_6892,N_5228,N_5008);
or U6893 (N_6893,N_5015,N_5976);
nor U6894 (N_6894,N_5392,N_5942);
xnor U6895 (N_6895,N_5494,N_5402);
or U6896 (N_6896,N_5051,N_5390);
and U6897 (N_6897,N_5452,N_5832);
nand U6898 (N_6898,N_5724,N_5979);
nand U6899 (N_6899,N_5982,N_5890);
and U6900 (N_6900,N_5114,N_5482);
xor U6901 (N_6901,N_5208,N_5838);
nand U6902 (N_6902,N_5790,N_5579);
and U6903 (N_6903,N_5799,N_5313);
xor U6904 (N_6904,N_5326,N_5116);
nand U6905 (N_6905,N_5341,N_5032);
xor U6906 (N_6906,N_5281,N_5607);
or U6907 (N_6907,N_5066,N_5062);
or U6908 (N_6908,N_5460,N_5237);
and U6909 (N_6909,N_5897,N_5574);
xnor U6910 (N_6910,N_5719,N_5948);
or U6911 (N_6911,N_5658,N_5780);
xnor U6912 (N_6912,N_5667,N_5049);
and U6913 (N_6913,N_5188,N_5121);
nand U6914 (N_6914,N_5342,N_5424);
or U6915 (N_6915,N_5264,N_5127);
and U6916 (N_6916,N_5251,N_5291);
nand U6917 (N_6917,N_5278,N_5297);
nand U6918 (N_6918,N_5078,N_5018);
nor U6919 (N_6919,N_5216,N_5841);
nand U6920 (N_6920,N_5983,N_5361);
and U6921 (N_6921,N_5342,N_5802);
nand U6922 (N_6922,N_5071,N_5063);
nand U6923 (N_6923,N_5512,N_5917);
xnor U6924 (N_6924,N_5620,N_5025);
and U6925 (N_6925,N_5481,N_5364);
or U6926 (N_6926,N_5567,N_5462);
or U6927 (N_6927,N_5227,N_5899);
and U6928 (N_6928,N_5196,N_5480);
or U6929 (N_6929,N_5957,N_5791);
xnor U6930 (N_6930,N_5671,N_5819);
and U6931 (N_6931,N_5039,N_5638);
xnor U6932 (N_6932,N_5086,N_5081);
xor U6933 (N_6933,N_5493,N_5922);
and U6934 (N_6934,N_5782,N_5855);
or U6935 (N_6935,N_5303,N_5982);
or U6936 (N_6936,N_5949,N_5815);
and U6937 (N_6937,N_5653,N_5960);
xnor U6938 (N_6938,N_5326,N_5491);
or U6939 (N_6939,N_5186,N_5382);
and U6940 (N_6940,N_5220,N_5640);
nand U6941 (N_6941,N_5382,N_5996);
or U6942 (N_6942,N_5603,N_5505);
nor U6943 (N_6943,N_5762,N_5631);
nor U6944 (N_6944,N_5966,N_5351);
nor U6945 (N_6945,N_5270,N_5833);
nand U6946 (N_6946,N_5006,N_5143);
and U6947 (N_6947,N_5097,N_5000);
xor U6948 (N_6948,N_5907,N_5403);
and U6949 (N_6949,N_5356,N_5090);
or U6950 (N_6950,N_5590,N_5106);
or U6951 (N_6951,N_5136,N_5189);
xnor U6952 (N_6952,N_5597,N_5353);
nand U6953 (N_6953,N_5535,N_5243);
xor U6954 (N_6954,N_5615,N_5048);
xor U6955 (N_6955,N_5540,N_5234);
or U6956 (N_6956,N_5234,N_5106);
nand U6957 (N_6957,N_5060,N_5483);
or U6958 (N_6958,N_5788,N_5778);
and U6959 (N_6959,N_5437,N_5545);
or U6960 (N_6960,N_5877,N_5755);
and U6961 (N_6961,N_5874,N_5963);
or U6962 (N_6962,N_5876,N_5062);
nor U6963 (N_6963,N_5897,N_5550);
nor U6964 (N_6964,N_5682,N_5342);
nor U6965 (N_6965,N_5020,N_5191);
xor U6966 (N_6966,N_5387,N_5078);
and U6967 (N_6967,N_5571,N_5967);
or U6968 (N_6968,N_5208,N_5885);
xor U6969 (N_6969,N_5930,N_5845);
nand U6970 (N_6970,N_5451,N_5540);
nand U6971 (N_6971,N_5452,N_5916);
xnor U6972 (N_6972,N_5904,N_5334);
nor U6973 (N_6973,N_5853,N_5623);
or U6974 (N_6974,N_5243,N_5734);
and U6975 (N_6975,N_5270,N_5830);
and U6976 (N_6976,N_5466,N_5950);
nor U6977 (N_6977,N_5798,N_5463);
xnor U6978 (N_6978,N_5948,N_5992);
and U6979 (N_6979,N_5226,N_5677);
xnor U6980 (N_6980,N_5999,N_5845);
nand U6981 (N_6981,N_5470,N_5405);
or U6982 (N_6982,N_5050,N_5214);
nor U6983 (N_6983,N_5393,N_5072);
and U6984 (N_6984,N_5274,N_5015);
xor U6985 (N_6985,N_5379,N_5214);
xor U6986 (N_6986,N_5716,N_5867);
nand U6987 (N_6987,N_5231,N_5624);
or U6988 (N_6988,N_5131,N_5814);
or U6989 (N_6989,N_5391,N_5173);
or U6990 (N_6990,N_5856,N_5705);
and U6991 (N_6991,N_5522,N_5726);
nand U6992 (N_6992,N_5607,N_5662);
xnor U6993 (N_6993,N_5694,N_5804);
nor U6994 (N_6994,N_5392,N_5004);
nand U6995 (N_6995,N_5406,N_5432);
or U6996 (N_6996,N_5200,N_5797);
or U6997 (N_6997,N_5444,N_5593);
xnor U6998 (N_6998,N_5220,N_5995);
or U6999 (N_6999,N_5203,N_5070);
or U7000 (N_7000,N_6201,N_6974);
nand U7001 (N_7001,N_6569,N_6587);
xor U7002 (N_7002,N_6849,N_6314);
nand U7003 (N_7003,N_6066,N_6609);
nand U7004 (N_7004,N_6038,N_6144);
xnor U7005 (N_7005,N_6394,N_6619);
or U7006 (N_7006,N_6866,N_6082);
nor U7007 (N_7007,N_6488,N_6355);
nand U7008 (N_7008,N_6207,N_6597);
and U7009 (N_7009,N_6812,N_6432);
nor U7010 (N_7010,N_6362,N_6146);
nand U7011 (N_7011,N_6834,N_6854);
nor U7012 (N_7012,N_6745,N_6277);
nor U7013 (N_7013,N_6899,N_6100);
nand U7014 (N_7014,N_6228,N_6474);
and U7015 (N_7015,N_6536,N_6612);
xnor U7016 (N_7016,N_6115,N_6708);
or U7017 (N_7017,N_6097,N_6752);
or U7018 (N_7018,N_6252,N_6946);
or U7019 (N_7019,N_6811,N_6683);
nor U7020 (N_7020,N_6578,N_6672);
and U7021 (N_7021,N_6200,N_6271);
nor U7022 (N_7022,N_6731,N_6113);
nor U7023 (N_7023,N_6724,N_6225);
and U7024 (N_7024,N_6985,N_6903);
or U7025 (N_7025,N_6922,N_6361);
xnor U7026 (N_7026,N_6127,N_6570);
nand U7027 (N_7027,N_6810,N_6494);
xor U7028 (N_7028,N_6801,N_6472);
and U7029 (N_7029,N_6136,N_6171);
xnor U7030 (N_7030,N_6017,N_6084);
and U7031 (N_7031,N_6514,N_6935);
xor U7032 (N_7032,N_6580,N_6680);
and U7033 (N_7033,N_6101,N_6936);
nor U7034 (N_7034,N_6546,N_6965);
and U7035 (N_7035,N_6908,N_6738);
or U7036 (N_7036,N_6972,N_6729);
or U7037 (N_7037,N_6143,N_6697);
nor U7038 (N_7038,N_6463,N_6667);
nand U7039 (N_7039,N_6960,N_6205);
nand U7040 (N_7040,N_6382,N_6033);
and U7041 (N_7041,N_6184,N_6118);
nand U7042 (N_7042,N_6349,N_6210);
nor U7043 (N_7043,N_6885,N_6178);
nand U7044 (N_7044,N_6319,N_6088);
nor U7045 (N_7045,N_6600,N_6458);
and U7046 (N_7046,N_6691,N_6336);
xor U7047 (N_7047,N_6931,N_6828);
xnor U7048 (N_7048,N_6313,N_6878);
nand U7049 (N_7049,N_6119,N_6354);
nor U7050 (N_7050,N_6071,N_6288);
xor U7051 (N_7051,N_6401,N_6552);
nand U7052 (N_7052,N_6913,N_6495);
nor U7053 (N_7053,N_6021,N_6593);
xor U7054 (N_7054,N_6562,N_6303);
xor U7055 (N_7055,N_6340,N_6765);
and U7056 (N_7056,N_6383,N_6756);
nand U7057 (N_7057,N_6864,N_6169);
xnor U7058 (N_7058,N_6278,N_6186);
or U7059 (N_7059,N_6841,N_6995);
nor U7060 (N_7060,N_6705,N_6821);
nor U7061 (N_7061,N_6945,N_6190);
nand U7062 (N_7062,N_6296,N_6188);
or U7063 (N_7063,N_6116,N_6723);
xor U7064 (N_7064,N_6370,N_6852);
and U7065 (N_7065,N_6457,N_6187);
or U7066 (N_7066,N_6363,N_6490);
and U7067 (N_7067,N_6316,N_6962);
xnor U7068 (N_7068,N_6531,N_6709);
xnor U7069 (N_7069,N_6895,N_6846);
or U7070 (N_7070,N_6031,N_6543);
or U7071 (N_7071,N_6439,N_6125);
xor U7072 (N_7072,N_6628,N_6173);
or U7073 (N_7073,N_6876,N_6371);
or U7074 (N_7074,N_6964,N_6501);
or U7075 (N_7075,N_6845,N_6627);
nor U7076 (N_7076,N_6838,N_6427);
and U7077 (N_7077,N_6366,N_6389);
xor U7078 (N_7078,N_6663,N_6180);
or U7079 (N_7079,N_6437,N_6605);
xor U7080 (N_7080,N_6504,N_6727);
nand U7081 (N_7081,N_6689,N_6179);
nor U7082 (N_7082,N_6739,N_6121);
xor U7083 (N_7083,N_6684,N_6994);
nor U7084 (N_7084,N_6796,N_6331);
nor U7085 (N_7085,N_6424,N_6728);
nand U7086 (N_7086,N_6741,N_6557);
xor U7087 (N_7087,N_6860,N_6137);
or U7088 (N_7088,N_6454,N_6615);
or U7089 (N_7089,N_6134,N_6231);
nand U7090 (N_7090,N_6699,N_6284);
nor U7091 (N_7091,N_6817,N_6568);
xor U7092 (N_7092,N_6259,N_6075);
and U7093 (N_7093,N_6668,N_6999);
nand U7094 (N_7094,N_6268,N_6461);
and U7095 (N_7095,N_6435,N_6926);
xnor U7096 (N_7096,N_6819,N_6286);
nand U7097 (N_7097,N_6011,N_6932);
and U7098 (N_7098,N_6620,N_6692);
or U7099 (N_7099,N_6799,N_6820);
nand U7100 (N_7100,N_6132,N_6548);
or U7101 (N_7101,N_6093,N_6338);
or U7102 (N_7102,N_6792,N_6662);
nor U7103 (N_7103,N_6090,N_6248);
or U7104 (N_7104,N_6954,N_6760);
nand U7105 (N_7105,N_6197,N_6884);
or U7106 (N_7106,N_6446,N_6123);
and U7107 (N_7107,N_6526,N_6152);
xnor U7108 (N_7108,N_6714,N_6001);
nor U7109 (N_7109,N_6824,N_6560);
xor U7110 (N_7110,N_6577,N_6579);
nand U7111 (N_7111,N_6258,N_6014);
or U7112 (N_7112,N_6287,N_6279);
nor U7113 (N_7113,N_6487,N_6528);
and U7114 (N_7114,N_6292,N_6897);
and U7115 (N_7115,N_6106,N_6216);
nand U7116 (N_7116,N_6540,N_6039);
or U7117 (N_7117,N_6256,N_6584);
or U7118 (N_7118,N_6914,N_6696);
and U7119 (N_7119,N_6889,N_6112);
and U7120 (N_7120,N_6059,N_6640);
or U7121 (N_7121,N_6529,N_6986);
xor U7122 (N_7122,N_6372,N_6069);
xnor U7123 (N_7123,N_6721,N_6212);
nand U7124 (N_7124,N_6678,N_6245);
nand U7125 (N_7125,N_6720,N_6227);
nor U7126 (N_7126,N_6676,N_6533);
or U7127 (N_7127,N_6153,N_6334);
xor U7128 (N_7128,N_6520,N_6208);
xnor U7129 (N_7129,N_6920,N_6462);
xor U7130 (N_7130,N_6753,N_6309);
nand U7131 (N_7131,N_6428,N_6639);
or U7132 (N_7132,N_6503,N_6912);
nor U7133 (N_7133,N_6892,N_6734);
xor U7134 (N_7134,N_6433,N_6596);
nor U7135 (N_7135,N_6235,N_6744);
nand U7136 (N_7136,N_6464,N_6452);
xor U7137 (N_7137,N_6673,N_6657);
nand U7138 (N_7138,N_6213,N_6358);
and U7139 (N_7139,N_6966,N_6471);
nor U7140 (N_7140,N_6545,N_6440);
nor U7141 (N_7141,N_6702,N_6388);
nor U7142 (N_7142,N_6157,N_6660);
and U7143 (N_7143,N_6040,N_6633);
nor U7144 (N_7144,N_6484,N_6698);
nor U7145 (N_7145,N_6110,N_6839);
xnor U7146 (N_7146,N_6230,N_6614);
xor U7147 (N_7147,N_6426,N_6594);
and U7148 (N_7148,N_6055,N_6324);
and U7149 (N_7149,N_6390,N_6583);
nand U7150 (N_7150,N_6675,N_6374);
and U7151 (N_7151,N_6518,N_6911);
nor U7152 (N_7152,N_6505,N_6647);
nand U7153 (N_7153,N_6131,N_6567);
nand U7154 (N_7154,N_6516,N_6599);
nand U7155 (N_7155,N_6951,N_6151);
nand U7156 (N_7156,N_6274,N_6666);
xor U7157 (N_7157,N_6209,N_6996);
and U7158 (N_7158,N_6735,N_6750);
nand U7159 (N_7159,N_6233,N_6621);
and U7160 (N_7160,N_6393,N_6322);
xor U7161 (N_7161,N_6757,N_6513);
nand U7162 (N_7162,N_6430,N_6973);
or U7163 (N_7163,N_6351,N_6875);
or U7164 (N_7164,N_6802,N_6970);
nor U7165 (N_7165,N_6403,N_6681);
nand U7166 (N_7166,N_6510,N_6581);
xnor U7167 (N_7167,N_6664,N_6805);
or U7168 (N_7168,N_6242,N_6105);
xor U7169 (N_7169,N_6375,N_6145);
xor U7170 (N_7170,N_6498,N_6489);
or U7171 (N_7171,N_6079,N_6298);
nand U7172 (N_7172,N_6019,N_6166);
nand U7173 (N_7173,N_6421,N_6719);
xnor U7174 (N_7174,N_6880,N_6299);
nor U7175 (N_7175,N_6831,N_6645);
or U7176 (N_7176,N_6434,N_6833);
nand U7177 (N_7177,N_6006,N_6005);
nand U7178 (N_7178,N_6671,N_6641);
and U7179 (N_7179,N_6783,N_6400);
nand U7180 (N_7180,N_6669,N_6991);
and U7181 (N_7181,N_6122,N_6422);
and U7182 (N_7182,N_6527,N_6195);
xnor U7183 (N_7183,N_6301,N_6626);
nand U7184 (N_7184,N_6532,N_6413);
xnor U7185 (N_7185,N_6830,N_6058);
or U7186 (N_7186,N_6406,N_6335);
nor U7187 (N_7187,N_6992,N_6193);
xor U7188 (N_7188,N_6764,N_6873);
and U7189 (N_7189,N_6653,N_6141);
and U7190 (N_7190,N_6930,N_6979);
nand U7191 (N_7191,N_6343,N_6679);
and U7192 (N_7192,N_6982,N_6987);
or U7193 (N_7193,N_6002,N_6191);
nor U7194 (N_7194,N_6969,N_6823);
nand U7195 (N_7195,N_6900,N_6417);
nand U7196 (N_7196,N_6337,N_6718);
or U7197 (N_7197,N_6219,N_6547);
nor U7198 (N_7198,N_6323,N_6674);
xor U7199 (N_7199,N_6923,N_6257);
or U7200 (N_7200,N_6565,N_6246);
or U7201 (N_7201,N_6704,N_6089);
nand U7202 (N_7202,N_6350,N_6469);
nor U7203 (N_7203,N_6402,N_6163);
nor U7204 (N_7204,N_6412,N_6953);
xor U7205 (N_7205,N_6077,N_6238);
xnor U7206 (N_7206,N_6008,N_6826);
nor U7207 (N_7207,N_6176,N_6386);
and U7208 (N_7208,N_6018,N_6070);
or U7209 (N_7209,N_6007,N_6120);
or U7210 (N_7210,N_6870,N_6524);
xor U7211 (N_7211,N_6326,N_6263);
and U7212 (N_7212,N_6815,N_6445);
and U7213 (N_7213,N_6379,N_6825);
nor U7214 (N_7214,N_6194,N_6384);
xor U7215 (N_7215,N_6816,N_6478);
nor U7216 (N_7216,N_6539,N_6407);
nand U7217 (N_7217,N_6293,N_6789);
xor U7218 (N_7218,N_6726,N_6598);
xnor U7219 (N_7219,N_6637,N_6650);
nor U7220 (N_7220,N_6102,N_6538);
and U7221 (N_7221,N_6218,N_6978);
or U7222 (N_7222,N_6273,N_6352);
and U7223 (N_7223,N_6509,N_6881);
and U7224 (N_7224,N_6677,N_6921);
xnor U7225 (N_7225,N_6555,N_6595);
nor U7226 (N_7226,N_6010,N_6096);
and U7227 (N_7227,N_6177,N_6665);
nor U7228 (N_7228,N_6712,N_6281);
nand U7229 (N_7229,N_6778,N_6061);
nor U7230 (N_7230,N_6170,N_6850);
nand U7231 (N_7231,N_6133,N_6499);
xnor U7232 (N_7232,N_6015,N_6138);
and U7233 (N_7233,N_6081,N_6837);
and U7234 (N_7234,N_6043,N_6332);
nand U7235 (N_7235,N_6943,N_6981);
xnor U7236 (N_7236,N_6732,N_6453);
xnor U7237 (N_7237,N_6198,N_6758);
and U7238 (N_7238,N_6196,N_6185);
or U7239 (N_7239,N_6203,N_6217);
or U7240 (N_7240,N_6302,N_6717);
nand U7241 (N_7241,N_6780,N_6571);
nor U7242 (N_7242,N_6874,N_6104);
or U7243 (N_7243,N_6763,N_6941);
xor U7244 (N_7244,N_6243,N_6103);
nand U7245 (N_7245,N_6859,N_6420);
nand U7246 (N_7246,N_6586,N_6976);
xnor U7247 (N_7247,N_6333,N_6901);
xor U7248 (N_7248,N_6575,N_6749);
nor U7249 (N_7249,N_6861,N_6894);
nand U7250 (N_7250,N_6507,N_6648);
xor U7251 (N_7251,N_6512,N_6211);
xor U7252 (N_7252,N_6632,N_6848);
xnor U7253 (N_7253,N_6775,N_6057);
nand U7254 (N_7254,N_6130,N_6500);
xnor U7255 (N_7255,N_6768,N_6020);
nor U7256 (N_7256,N_6787,N_6346);
xor U7257 (N_7257,N_6856,N_6441);
xnor U7258 (N_7258,N_6730,N_6624);
and U7259 (N_7259,N_6294,N_6934);
or U7260 (N_7260,N_6843,N_6751);
xnor U7261 (N_7261,N_6927,N_6634);
or U7262 (N_7262,N_6016,N_6162);
xnor U7263 (N_7263,N_6431,N_6686);
and U7264 (N_7264,N_6161,N_6916);
nor U7265 (N_7265,N_6036,N_6755);
or U7266 (N_7266,N_6521,N_6267);
xor U7267 (N_7267,N_6502,N_6658);
xnor U7268 (N_7268,N_6491,N_6013);
nor U7269 (N_7269,N_6415,N_6553);
or U7270 (N_7270,N_6904,N_6638);
xnor U7271 (N_7271,N_6782,N_6442);
nor U7272 (N_7272,N_6844,N_6327);
xor U7273 (N_7273,N_6618,N_6554);
or U7274 (N_7274,N_6047,N_6906);
nand U7275 (N_7275,N_6592,N_6154);
or U7276 (N_7276,N_6998,N_6392);
or U7277 (N_7277,N_6736,N_6940);
nor U7278 (N_7278,N_6467,N_6305);
nand U7279 (N_7279,N_6168,N_6492);
xor U7280 (N_7280,N_6290,N_6050);
nand U7281 (N_7281,N_6344,N_6202);
xor U7282 (N_7282,N_6221,N_6308);
xnor U7283 (N_7283,N_6054,N_6387);
or U7284 (N_7284,N_6476,N_6771);
nor U7285 (N_7285,N_6380,N_6670);
nand U7286 (N_7286,N_6167,N_6601);
or U7287 (N_7287,N_6032,N_6397);
and U7288 (N_7288,N_6368,N_6591);
and U7289 (N_7289,N_6456,N_6073);
nor U7290 (N_7290,N_6952,N_6646);
xor U7291 (N_7291,N_6888,N_6297);
and U7292 (N_7292,N_6949,N_6049);
nand U7293 (N_7293,N_6902,N_6147);
or U7294 (N_7294,N_6865,N_6784);
nand U7295 (N_7295,N_6409,N_6360);
or U7296 (N_7296,N_6944,N_6947);
xnor U7297 (N_7297,N_6264,N_6416);
and U7298 (N_7298,N_6530,N_6656);
nand U7299 (N_7299,N_6980,N_6408);
nor U7300 (N_7300,N_6482,N_6522);
nor U7301 (N_7301,N_6740,N_6030);
nor U7302 (N_7302,N_6385,N_6239);
or U7303 (N_7303,N_6369,N_6270);
nand U7304 (N_7304,N_6321,N_6448);
nor U7305 (N_7305,N_6939,N_6206);
nor U7306 (N_7306,N_6269,N_6291);
nor U7307 (N_7307,N_6304,N_6769);
or U7308 (N_7308,N_6318,N_6808);
xor U7309 (N_7309,N_6000,N_6788);
nand U7310 (N_7310,N_6260,N_6480);
and U7311 (N_7311,N_6687,N_6928);
nor U7312 (N_7312,N_6156,N_6139);
nor U7313 (N_7313,N_6485,N_6181);
or U7314 (N_7314,N_6710,N_6087);
and U7315 (N_7315,N_6142,N_6465);
nand U7316 (N_7316,N_6777,N_6247);
or U7317 (N_7317,N_6023,N_6971);
nand U7318 (N_7318,N_6051,N_6045);
xnor U7319 (N_7319,N_6542,N_6517);
xor U7320 (N_7320,N_6929,N_6479);
nand U7321 (N_7321,N_6265,N_6429);
nor U7322 (N_7322,N_6779,N_6887);
or U7323 (N_7323,N_6715,N_6857);
xnor U7324 (N_7324,N_6357,N_6411);
nor U7325 (N_7325,N_6182,N_6655);
or U7326 (N_7326,N_6942,N_6958);
xnor U7327 (N_7327,N_6898,N_6086);
or U7328 (N_7328,N_6048,N_6128);
nand U7329 (N_7329,N_6255,N_6470);
or U7330 (N_7330,N_6737,N_6649);
nand U7331 (N_7331,N_6872,N_6549);
nand U7332 (N_7332,N_6004,N_6395);
xor U7333 (N_7333,N_6042,N_6391);
and U7334 (N_7334,N_6983,N_6716);
nand U7335 (N_7335,N_6933,N_6907);
xor U7336 (N_7336,N_6094,N_6695);
and U7337 (N_7337,N_6604,N_6289);
and U7338 (N_7338,N_6251,N_6317);
xor U7339 (N_7339,N_6266,N_6244);
nand U7340 (N_7340,N_6091,N_6607);
and U7341 (N_7341,N_6525,N_6558);
nand U7342 (N_7342,N_6468,N_6977);
and U7343 (N_7343,N_6064,N_6481);
xnor U7344 (N_7344,N_6842,N_6766);
nand U7345 (N_7345,N_6204,N_6272);
or U7346 (N_7346,N_6827,N_6652);
xnor U7347 (N_7347,N_6012,N_6886);
or U7348 (N_7348,N_6993,N_6083);
or U7349 (N_7349,N_6642,N_6871);
nand U7350 (N_7350,N_6438,N_6742);
nor U7351 (N_7351,N_6956,N_6688);
xor U7352 (N_7352,N_6192,N_6910);
nor U7353 (N_7353,N_6046,N_6328);
xor U7354 (N_7354,N_6114,N_6067);
xor U7355 (N_7355,N_6798,N_6813);
nand U7356 (N_7356,N_6229,N_6785);
nand U7357 (N_7357,N_6800,N_6330);
and U7358 (N_7358,N_6155,N_6585);
nor U7359 (N_7359,N_6795,N_6353);
nor U7360 (N_7360,N_6733,N_6475);
or U7361 (N_7361,N_6711,N_6148);
nor U7362 (N_7362,N_6781,N_6616);
nor U7363 (N_7363,N_6589,N_6867);
xnor U7364 (N_7364,N_6034,N_6280);
xor U7365 (N_7365,N_6832,N_6804);
nor U7366 (N_7366,N_6603,N_6300);
nand U7367 (N_7367,N_6561,N_6028);
and U7368 (N_7368,N_6572,N_6232);
nor U7369 (N_7369,N_6451,N_6224);
and U7370 (N_7370,N_6312,N_6635);
nand U7371 (N_7371,N_6822,N_6793);
nor U7372 (N_7372,N_6925,N_6611);
nand U7373 (N_7373,N_6356,N_6172);
nor U7374 (N_7374,N_6713,N_6275);
nor U7375 (N_7375,N_6065,N_6025);
nor U7376 (N_7376,N_6905,N_6342);
xnor U7377 (N_7377,N_6078,N_6541);
or U7378 (N_7378,N_6165,N_6877);
or U7379 (N_7379,N_6563,N_6701);
nor U7380 (N_7380,N_6997,N_6534);
nand U7381 (N_7381,N_6234,N_6938);
or U7382 (N_7382,N_6636,N_6035);
or U7383 (N_7383,N_6550,N_6261);
or U7384 (N_7384,N_6746,N_6215);
nand U7385 (N_7385,N_6809,N_6590);
or U7386 (N_7386,N_6341,N_6968);
nor U7387 (N_7387,N_6836,N_6044);
nor U7388 (N_7388,N_6535,N_6307);
or U7389 (N_7389,N_6918,N_6365);
and U7390 (N_7390,N_6582,N_6556);
nand U7391 (N_7391,N_6449,N_6606);
nor U7392 (N_7392,N_6311,N_6770);
or U7393 (N_7393,N_6685,N_6450);
and U7394 (N_7394,N_6226,N_6282);
nand U7395 (N_7395,N_6851,N_6347);
xor U7396 (N_7396,N_6483,N_6060);
xor U7397 (N_7397,N_6074,N_6310);
and U7398 (N_7398,N_6117,N_6348);
xnor U7399 (N_7399,N_6486,N_6378);
and U7400 (N_7400,N_6948,N_6419);
nand U7401 (N_7401,N_6359,N_6963);
and U7402 (N_7402,N_6644,N_6460);
xor U7403 (N_7403,N_6630,N_6791);
and U7404 (N_7404,N_6706,N_6773);
nand U7405 (N_7405,N_6092,N_6608);
nor U7406 (N_7406,N_6703,N_6099);
or U7407 (N_7407,N_6855,N_6984);
or U7408 (N_7408,N_6975,N_6436);
or U7409 (N_7409,N_6772,N_6544);
and U7410 (N_7410,N_6220,N_6937);
xor U7411 (N_7411,N_6126,N_6806);
nand U7412 (N_7412,N_6576,N_6329);
nand U7413 (N_7413,N_6869,N_6283);
or U7414 (N_7414,N_6957,N_6829);
xor U7415 (N_7415,N_6896,N_6276);
nor U7416 (N_7416,N_6803,N_6573);
xnor U7417 (N_7417,N_6241,N_6108);
nand U7418 (N_7418,N_6654,N_6062);
nand U7419 (N_7419,N_6443,N_6214);
xor U7420 (N_7420,N_6262,N_6041);
nor U7421 (N_7421,N_6022,N_6423);
or U7422 (N_7422,N_6858,N_6661);
nand U7423 (N_7423,N_6250,N_6508);
nand U7424 (N_7424,N_6707,N_6891);
nand U7425 (N_7425,N_6790,N_6915);
and U7426 (N_7426,N_6853,N_6882);
or U7427 (N_7427,N_6497,N_6519);
and U7428 (N_7428,N_6748,N_6240);
or U7429 (N_7429,N_6295,N_6694);
nor U7430 (N_7430,N_6722,N_6767);
nand U7431 (N_7431,N_6072,N_6418);
or U7432 (N_7432,N_6919,N_6140);
or U7433 (N_7433,N_6523,N_6135);
nand U7434 (N_7434,N_6863,N_6818);
and U7435 (N_7435,N_6076,N_6414);
nand U7436 (N_7436,N_6690,N_6774);
nor U7437 (N_7437,N_6236,N_6659);
nand U7438 (N_7438,N_6098,N_6222);
xnor U7439 (N_7439,N_6990,N_6367);
nor U7440 (N_7440,N_6399,N_6003);
and U7441 (N_7441,N_6564,N_6610);
or U7442 (N_7442,N_6223,N_6325);
nor U7443 (N_7443,N_6183,N_6339);
nand U7444 (N_7444,N_6024,N_6080);
or U7445 (N_7445,N_6743,N_6381);
and U7446 (N_7446,N_6879,N_6794);
nor U7447 (N_7447,N_6477,N_6455);
xor U7448 (N_7448,N_6959,N_6373);
nor U7449 (N_7449,N_6754,N_6149);
or U7450 (N_7450,N_6693,N_6063);
xnor U7451 (N_7451,N_6776,N_6700);
or U7452 (N_7452,N_6364,N_6009);
xnor U7453 (N_7453,N_6164,N_6053);
and U7454 (N_7454,N_6835,N_6883);
nor U7455 (N_7455,N_6566,N_6315);
nor U7456 (N_7456,N_6506,N_6629);
xnor U7457 (N_7457,N_6559,N_6909);
nor U7458 (N_7458,N_6989,N_6924);
nor U7459 (N_7459,N_6345,N_6249);
or U7460 (N_7460,N_6761,N_6306);
nor U7461 (N_7461,N_6955,N_6253);
xnor U7462 (N_7462,N_6320,N_6551);
and U7463 (N_7463,N_6961,N_6496);
and U7464 (N_7464,N_6068,N_6029);
or U7465 (N_7465,N_6537,N_6158);
nor U7466 (N_7466,N_6160,N_6613);
nor U7467 (N_7467,N_6868,N_6199);
and U7468 (N_7468,N_6376,N_6651);
nor U7469 (N_7469,N_6159,N_6396);
and U7470 (N_7470,N_6175,N_6515);
and U7471 (N_7471,N_6631,N_6237);
nand U7472 (N_7472,N_6950,N_6285);
xor U7473 (N_7473,N_6052,N_6967);
or U7474 (N_7474,N_6410,N_6814);
xnor U7475 (N_7475,N_6027,N_6444);
or U7476 (N_7476,N_6493,N_6890);
nor U7477 (N_7477,N_6189,N_6447);
and U7478 (N_7478,N_6174,N_6124);
and U7479 (N_7479,N_6377,N_6404);
nor U7480 (N_7480,N_6807,N_6797);
nand U7481 (N_7481,N_6840,N_6107);
and U7482 (N_7482,N_6623,N_6095);
and U7483 (N_7483,N_6425,N_6847);
nor U7484 (N_7484,N_6085,N_6762);
and U7485 (N_7485,N_6150,N_6466);
xnor U7486 (N_7486,N_6398,N_6617);
or U7487 (N_7487,N_6511,N_6602);
xor U7488 (N_7488,N_6405,N_6893);
nor U7489 (N_7489,N_6026,N_6473);
or U7490 (N_7490,N_6588,N_6643);
xnor U7491 (N_7491,N_6056,N_6862);
and U7492 (N_7492,N_6254,N_6129);
or U7493 (N_7493,N_6917,N_6037);
nand U7494 (N_7494,N_6625,N_6747);
and U7495 (N_7495,N_6725,N_6622);
nand U7496 (N_7496,N_6459,N_6111);
nand U7497 (N_7497,N_6574,N_6682);
xnor U7498 (N_7498,N_6109,N_6988);
nor U7499 (N_7499,N_6759,N_6786);
or U7500 (N_7500,N_6584,N_6353);
nand U7501 (N_7501,N_6449,N_6274);
and U7502 (N_7502,N_6506,N_6947);
or U7503 (N_7503,N_6286,N_6022);
or U7504 (N_7504,N_6270,N_6150);
or U7505 (N_7505,N_6045,N_6286);
or U7506 (N_7506,N_6469,N_6405);
nor U7507 (N_7507,N_6838,N_6697);
and U7508 (N_7508,N_6435,N_6485);
or U7509 (N_7509,N_6617,N_6481);
nand U7510 (N_7510,N_6840,N_6310);
nand U7511 (N_7511,N_6571,N_6692);
nor U7512 (N_7512,N_6846,N_6361);
xnor U7513 (N_7513,N_6618,N_6183);
xnor U7514 (N_7514,N_6973,N_6247);
and U7515 (N_7515,N_6012,N_6142);
nand U7516 (N_7516,N_6823,N_6765);
xnor U7517 (N_7517,N_6299,N_6697);
xnor U7518 (N_7518,N_6465,N_6946);
and U7519 (N_7519,N_6025,N_6181);
nor U7520 (N_7520,N_6579,N_6133);
nand U7521 (N_7521,N_6122,N_6670);
or U7522 (N_7522,N_6817,N_6342);
nor U7523 (N_7523,N_6615,N_6779);
and U7524 (N_7524,N_6137,N_6635);
and U7525 (N_7525,N_6895,N_6205);
xnor U7526 (N_7526,N_6267,N_6899);
or U7527 (N_7527,N_6728,N_6747);
nor U7528 (N_7528,N_6362,N_6244);
nand U7529 (N_7529,N_6052,N_6775);
nand U7530 (N_7530,N_6898,N_6945);
nand U7531 (N_7531,N_6959,N_6238);
and U7532 (N_7532,N_6148,N_6017);
nand U7533 (N_7533,N_6612,N_6879);
nor U7534 (N_7534,N_6324,N_6719);
nand U7535 (N_7535,N_6374,N_6029);
nand U7536 (N_7536,N_6453,N_6086);
and U7537 (N_7537,N_6744,N_6930);
xnor U7538 (N_7538,N_6868,N_6413);
xor U7539 (N_7539,N_6313,N_6712);
nand U7540 (N_7540,N_6381,N_6882);
xor U7541 (N_7541,N_6227,N_6986);
nor U7542 (N_7542,N_6075,N_6221);
nand U7543 (N_7543,N_6091,N_6369);
nor U7544 (N_7544,N_6904,N_6283);
nor U7545 (N_7545,N_6178,N_6427);
nor U7546 (N_7546,N_6055,N_6555);
nor U7547 (N_7547,N_6697,N_6530);
xnor U7548 (N_7548,N_6463,N_6744);
and U7549 (N_7549,N_6750,N_6005);
xor U7550 (N_7550,N_6012,N_6363);
or U7551 (N_7551,N_6791,N_6591);
and U7552 (N_7552,N_6574,N_6553);
nand U7553 (N_7553,N_6469,N_6465);
nor U7554 (N_7554,N_6499,N_6801);
and U7555 (N_7555,N_6645,N_6817);
nor U7556 (N_7556,N_6902,N_6094);
nor U7557 (N_7557,N_6429,N_6433);
and U7558 (N_7558,N_6635,N_6483);
xor U7559 (N_7559,N_6135,N_6131);
or U7560 (N_7560,N_6018,N_6429);
and U7561 (N_7561,N_6569,N_6952);
or U7562 (N_7562,N_6320,N_6577);
nor U7563 (N_7563,N_6210,N_6799);
xnor U7564 (N_7564,N_6933,N_6428);
and U7565 (N_7565,N_6330,N_6194);
or U7566 (N_7566,N_6567,N_6868);
nor U7567 (N_7567,N_6288,N_6214);
nor U7568 (N_7568,N_6567,N_6141);
nand U7569 (N_7569,N_6404,N_6700);
nor U7570 (N_7570,N_6951,N_6456);
nand U7571 (N_7571,N_6884,N_6970);
xor U7572 (N_7572,N_6481,N_6704);
xor U7573 (N_7573,N_6814,N_6337);
or U7574 (N_7574,N_6959,N_6745);
or U7575 (N_7575,N_6259,N_6322);
xnor U7576 (N_7576,N_6107,N_6376);
and U7577 (N_7577,N_6524,N_6410);
nand U7578 (N_7578,N_6758,N_6843);
xnor U7579 (N_7579,N_6292,N_6490);
and U7580 (N_7580,N_6543,N_6809);
nand U7581 (N_7581,N_6489,N_6384);
xnor U7582 (N_7582,N_6460,N_6354);
or U7583 (N_7583,N_6704,N_6079);
nand U7584 (N_7584,N_6753,N_6355);
nand U7585 (N_7585,N_6768,N_6169);
nand U7586 (N_7586,N_6846,N_6771);
nor U7587 (N_7587,N_6463,N_6673);
and U7588 (N_7588,N_6438,N_6824);
xnor U7589 (N_7589,N_6424,N_6949);
nor U7590 (N_7590,N_6705,N_6216);
or U7591 (N_7591,N_6752,N_6906);
and U7592 (N_7592,N_6965,N_6599);
nand U7593 (N_7593,N_6789,N_6967);
nand U7594 (N_7594,N_6425,N_6843);
nor U7595 (N_7595,N_6600,N_6558);
or U7596 (N_7596,N_6323,N_6504);
nor U7597 (N_7597,N_6151,N_6578);
nand U7598 (N_7598,N_6535,N_6601);
and U7599 (N_7599,N_6887,N_6865);
xor U7600 (N_7600,N_6262,N_6237);
or U7601 (N_7601,N_6420,N_6172);
nor U7602 (N_7602,N_6748,N_6208);
nand U7603 (N_7603,N_6675,N_6467);
xor U7604 (N_7604,N_6960,N_6994);
xor U7605 (N_7605,N_6885,N_6079);
and U7606 (N_7606,N_6230,N_6725);
nand U7607 (N_7607,N_6573,N_6109);
nand U7608 (N_7608,N_6487,N_6879);
nand U7609 (N_7609,N_6234,N_6979);
xnor U7610 (N_7610,N_6090,N_6490);
xnor U7611 (N_7611,N_6739,N_6451);
nand U7612 (N_7612,N_6993,N_6243);
nand U7613 (N_7613,N_6687,N_6048);
nand U7614 (N_7614,N_6079,N_6245);
nor U7615 (N_7615,N_6124,N_6231);
and U7616 (N_7616,N_6742,N_6179);
xor U7617 (N_7617,N_6732,N_6000);
and U7618 (N_7618,N_6635,N_6563);
and U7619 (N_7619,N_6958,N_6168);
nand U7620 (N_7620,N_6102,N_6485);
nand U7621 (N_7621,N_6654,N_6868);
and U7622 (N_7622,N_6134,N_6496);
and U7623 (N_7623,N_6658,N_6692);
xnor U7624 (N_7624,N_6969,N_6664);
nor U7625 (N_7625,N_6548,N_6510);
nor U7626 (N_7626,N_6578,N_6649);
or U7627 (N_7627,N_6882,N_6801);
or U7628 (N_7628,N_6501,N_6300);
nor U7629 (N_7629,N_6194,N_6772);
nand U7630 (N_7630,N_6833,N_6506);
and U7631 (N_7631,N_6388,N_6082);
nand U7632 (N_7632,N_6205,N_6851);
xor U7633 (N_7633,N_6268,N_6568);
xnor U7634 (N_7634,N_6127,N_6973);
nand U7635 (N_7635,N_6053,N_6773);
and U7636 (N_7636,N_6571,N_6377);
nand U7637 (N_7637,N_6492,N_6769);
xnor U7638 (N_7638,N_6575,N_6457);
nor U7639 (N_7639,N_6103,N_6852);
xor U7640 (N_7640,N_6957,N_6590);
xnor U7641 (N_7641,N_6426,N_6313);
or U7642 (N_7642,N_6629,N_6041);
and U7643 (N_7643,N_6287,N_6629);
nand U7644 (N_7644,N_6801,N_6096);
nor U7645 (N_7645,N_6431,N_6166);
and U7646 (N_7646,N_6645,N_6102);
nor U7647 (N_7647,N_6407,N_6668);
and U7648 (N_7648,N_6261,N_6173);
or U7649 (N_7649,N_6052,N_6039);
xor U7650 (N_7650,N_6466,N_6433);
or U7651 (N_7651,N_6567,N_6486);
nor U7652 (N_7652,N_6377,N_6291);
xnor U7653 (N_7653,N_6947,N_6178);
or U7654 (N_7654,N_6645,N_6821);
xnor U7655 (N_7655,N_6076,N_6304);
nand U7656 (N_7656,N_6928,N_6019);
nand U7657 (N_7657,N_6407,N_6012);
xnor U7658 (N_7658,N_6212,N_6767);
nor U7659 (N_7659,N_6338,N_6091);
xnor U7660 (N_7660,N_6674,N_6418);
nand U7661 (N_7661,N_6399,N_6839);
or U7662 (N_7662,N_6220,N_6070);
nand U7663 (N_7663,N_6464,N_6336);
xor U7664 (N_7664,N_6487,N_6007);
or U7665 (N_7665,N_6826,N_6695);
nand U7666 (N_7666,N_6117,N_6456);
xor U7667 (N_7667,N_6022,N_6383);
or U7668 (N_7668,N_6042,N_6788);
xor U7669 (N_7669,N_6629,N_6712);
nor U7670 (N_7670,N_6016,N_6349);
and U7671 (N_7671,N_6179,N_6030);
and U7672 (N_7672,N_6735,N_6785);
nor U7673 (N_7673,N_6497,N_6359);
or U7674 (N_7674,N_6399,N_6521);
nand U7675 (N_7675,N_6071,N_6983);
or U7676 (N_7676,N_6029,N_6774);
or U7677 (N_7677,N_6645,N_6290);
xnor U7678 (N_7678,N_6657,N_6811);
or U7679 (N_7679,N_6602,N_6789);
nor U7680 (N_7680,N_6964,N_6412);
nor U7681 (N_7681,N_6334,N_6575);
xor U7682 (N_7682,N_6353,N_6014);
nand U7683 (N_7683,N_6478,N_6975);
nor U7684 (N_7684,N_6385,N_6339);
or U7685 (N_7685,N_6072,N_6923);
and U7686 (N_7686,N_6232,N_6001);
or U7687 (N_7687,N_6084,N_6316);
nand U7688 (N_7688,N_6531,N_6285);
xor U7689 (N_7689,N_6096,N_6965);
and U7690 (N_7690,N_6949,N_6815);
and U7691 (N_7691,N_6591,N_6715);
and U7692 (N_7692,N_6282,N_6783);
nand U7693 (N_7693,N_6067,N_6941);
nand U7694 (N_7694,N_6348,N_6192);
xnor U7695 (N_7695,N_6972,N_6005);
xor U7696 (N_7696,N_6238,N_6341);
or U7697 (N_7697,N_6449,N_6187);
and U7698 (N_7698,N_6977,N_6276);
nor U7699 (N_7699,N_6719,N_6895);
nor U7700 (N_7700,N_6678,N_6029);
nor U7701 (N_7701,N_6036,N_6215);
nor U7702 (N_7702,N_6039,N_6982);
nand U7703 (N_7703,N_6005,N_6471);
nand U7704 (N_7704,N_6334,N_6809);
and U7705 (N_7705,N_6574,N_6412);
nand U7706 (N_7706,N_6481,N_6102);
xnor U7707 (N_7707,N_6431,N_6064);
and U7708 (N_7708,N_6858,N_6926);
nor U7709 (N_7709,N_6383,N_6099);
and U7710 (N_7710,N_6492,N_6081);
and U7711 (N_7711,N_6140,N_6162);
xor U7712 (N_7712,N_6193,N_6730);
or U7713 (N_7713,N_6928,N_6854);
nand U7714 (N_7714,N_6428,N_6807);
nand U7715 (N_7715,N_6094,N_6803);
and U7716 (N_7716,N_6885,N_6543);
nand U7717 (N_7717,N_6118,N_6514);
nand U7718 (N_7718,N_6624,N_6973);
xor U7719 (N_7719,N_6197,N_6807);
nand U7720 (N_7720,N_6336,N_6870);
xor U7721 (N_7721,N_6155,N_6913);
xor U7722 (N_7722,N_6460,N_6870);
nand U7723 (N_7723,N_6863,N_6061);
nor U7724 (N_7724,N_6251,N_6940);
nor U7725 (N_7725,N_6283,N_6180);
or U7726 (N_7726,N_6188,N_6480);
or U7727 (N_7727,N_6025,N_6504);
nor U7728 (N_7728,N_6676,N_6375);
xnor U7729 (N_7729,N_6635,N_6656);
or U7730 (N_7730,N_6176,N_6576);
and U7731 (N_7731,N_6195,N_6876);
and U7732 (N_7732,N_6804,N_6194);
nor U7733 (N_7733,N_6669,N_6211);
nor U7734 (N_7734,N_6770,N_6160);
and U7735 (N_7735,N_6597,N_6708);
xnor U7736 (N_7736,N_6686,N_6948);
or U7737 (N_7737,N_6452,N_6077);
nor U7738 (N_7738,N_6887,N_6824);
xnor U7739 (N_7739,N_6507,N_6186);
and U7740 (N_7740,N_6256,N_6132);
and U7741 (N_7741,N_6643,N_6687);
xnor U7742 (N_7742,N_6992,N_6352);
nand U7743 (N_7743,N_6691,N_6555);
nor U7744 (N_7744,N_6911,N_6380);
nor U7745 (N_7745,N_6977,N_6589);
and U7746 (N_7746,N_6355,N_6228);
nor U7747 (N_7747,N_6063,N_6356);
xnor U7748 (N_7748,N_6794,N_6308);
xnor U7749 (N_7749,N_6240,N_6294);
nor U7750 (N_7750,N_6391,N_6959);
and U7751 (N_7751,N_6085,N_6569);
or U7752 (N_7752,N_6281,N_6920);
nor U7753 (N_7753,N_6119,N_6266);
nand U7754 (N_7754,N_6387,N_6497);
and U7755 (N_7755,N_6997,N_6490);
or U7756 (N_7756,N_6250,N_6948);
or U7757 (N_7757,N_6382,N_6781);
nand U7758 (N_7758,N_6129,N_6036);
nand U7759 (N_7759,N_6737,N_6132);
or U7760 (N_7760,N_6908,N_6986);
xnor U7761 (N_7761,N_6929,N_6225);
and U7762 (N_7762,N_6771,N_6371);
nor U7763 (N_7763,N_6587,N_6203);
nand U7764 (N_7764,N_6129,N_6595);
and U7765 (N_7765,N_6744,N_6756);
nand U7766 (N_7766,N_6924,N_6229);
nand U7767 (N_7767,N_6027,N_6016);
or U7768 (N_7768,N_6795,N_6992);
nor U7769 (N_7769,N_6384,N_6998);
nor U7770 (N_7770,N_6401,N_6957);
and U7771 (N_7771,N_6391,N_6015);
nand U7772 (N_7772,N_6319,N_6811);
nand U7773 (N_7773,N_6237,N_6246);
nor U7774 (N_7774,N_6302,N_6191);
or U7775 (N_7775,N_6244,N_6813);
xor U7776 (N_7776,N_6743,N_6823);
xnor U7777 (N_7777,N_6201,N_6206);
and U7778 (N_7778,N_6833,N_6166);
and U7779 (N_7779,N_6902,N_6336);
or U7780 (N_7780,N_6663,N_6744);
xor U7781 (N_7781,N_6295,N_6065);
or U7782 (N_7782,N_6961,N_6022);
nand U7783 (N_7783,N_6678,N_6694);
xor U7784 (N_7784,N_6856,N_6533);
nand U7785 (N_7785,N_6997,N_6945);
and U7786 (N_7786,N_6635,N_6009);
and U7787 (N_7787,N_6602,N_6722);
and U7788 (N_7788,N_6588,N_6916);
or U7789 (N_7789,N_6477,N_6354);
or U7790 (N_7790,N_6158,N_6452);
and U7791 (N_7791,N_6314,N_6057);
or U7792 (N_7792,N_6484,N_6359);
nor U7793 (N_7793,N_6262,N_6790);
nor U7794 (N_7794,N_6231,N_6161);
nor U7795 (N_7795,N_6629,N_6430);
and U7796 (N_7796,N_6308,N_6331);
xor U7797 (N_7797,N_6822,N_6176);
and U7798 (N_7798,N_6936,N_6824);
nand U7799 (N_7799,N_6683,N_6782);
nor U7800 (N_7800,N_6851,N_6549);
nand U7801 (N_7801,N_6407,N_6492);
nor U7802 (N_7802,N_6948,N_6699);
xor U7803 (N_7803,N_6836,N_6723);
xor U7804 (N_7804,N_6832,N_6418);
nand U7805 (N_7805,N_6920,N_6632);
nor U7806 (N_7806,N_6426,N_6223);
and U7807 (N_7807,N_6944,N_6445);
nor U7808 (N_7808,N_6148,N_6699);
xor U7809 (N_7809,N_6797,N_6198);
or U7810 (N_7810,N_6558,N_6651);
nor U7811 (N_7811,N_6533,N_6346);
xnor U7812 (N_7812,N_6654,N_6664);
or U7813 (N_7813,N_6533,N_6144);
nand U7814 (N_7814,N_6735,N_6035);
and U7815 (N_7815,N_6005,N_6256);
nor U7816 (N_7816,N_6342,N_6212);
xnor U7817 (N_7817,N_6467,N_6213);
or U7818 (N_7818,N_6955,N_6504);
nand U7819 (N_7819,N_6811,N_6529);
and U7820 (N_7820,N_6272,N_6725);
nand U7821 (N_7821,N_6298,N_6871);
nor U7822 (N_7822,N_6879,N_6415);
nor U7823 (N_7823,N_6362,N_6723);
nand U7824 (N_7824,N_6799,N_6886);
nor U7825 (N_7825,N_6432,N_6427);
or U7826 (N_7826,N_6888,N_6217);
or U7827 (N_7827,N_6704,N_6272);
nand U7828 (N_7828,N_6273,N_6320);
nor U7829 (N_7829,N_6380,N_6102);
nand U7830 (N_7830,N_6304,N_6320);
xor U7831 (N_7831,N_6318,N_6297);
or U7832 (N_7832,N_6764,N_6371);
nand U7833 (N_7833,N_6673,N_6560);
or U7834 (N_7834,N_6244,N_6292);
xor U7835 (N_7835,N_6574,N_6825);
xnor U7836 (N_7836,N_6585,N_6815);
nand U7837 (N_7837,N_6985,N_6029);
nand U7838 (N_7838,N_6882,N_6856);
nand U7839 (N_7839,N_6277,N_6954);
xor U7840 (N_7840,N_6613,N_6203);
xnor U7841 (N_7841,N_6893,N_6913);
and U7842 (N_7842,N_6536,N_6179);
and U7843 (N_7843,N_6910,N_6441);
nand U7844 (N_7844,N_6719,N_6527);
or U7845 (N_7845,N_6405,N_6601);
nand U7846 (N_7846,N_6941,N_6454);
nand U7847 (N_7847,N_6719,N_6176);
xor U7848 (N_7848,N_6222,N_6544);
nor U7849 (N_7849,N_6663,N_6667);
xor U7850 (N_7850,N_6875,N_6356);
nor U7851 (N_7851,N_6259,N_6720);
and U7852 (N_7852,N_6281,N_6239);
or U7853 (N_7853,N_6882,N_6063);
and U7854 (N_7854,N_6931,N_6380);
nor U7855 (N_7855,N_6790,N_6836);
nor U7856 (N_7856,N_6907,N_6749);
nand U7857 (N_7857,N_6981,N_6907);
nor U7858 (N_7858,N_6357,N_6121);
or U7859 (N_7859,N_6100,N_6835);
or U7860 (N_7860,N_6821,N_6230);
xor U7861 (N_7861,N_6808,N_6849);
and U7862 (N_7862,N_6783,N_6329);
nor U7863 (N_7863,N_6636,N_6429);
nand U7864 (N_7864,N_6425,N_6490);
and U7865 (N_7865,N_6303,N_6672);
and U7866 (N_7866,N_6777,N_6026);
nand U7867 (N_7867,N_6068,N_6065);
nand U7868 (N_7868,N_6176,N_6875);
and U7869 (N_7869,N_6547,N_6484);
or U7870 (N_7870,N_6943,N_6702);
xnor U7871 (N_7871,N_6462,N_6788);
or U7872 (N_7872,N_6921,N_6885);
xnor U7873 (N_7873,N_6785,N_6617);
and U7874 (N_7874,N_6917,N_6019);
and U7875 (N_7875,N_6688,N_6378);
and U7876 (N_7876,N_6389,N_6381);
nand U7877 (N_7877,N_6195,N_6536);
nor U7878 (N_7878,N_6974,N_6265);
and U7879 (N_7879,N_6457,N_6525);
nand U7880 (N_7880,N_6645,N_6364);
and U7881 (N_7881,N_6955,N_6361);
xor U7882 (N_7882,N_6373,N_6966);
xnor U7883 (N_7883,N_6017,N_6034);
or U7884 (N_7884,N_6086,N_6004);
nand U7885 (N_7885,N_6089,N_6508);
or U7886 (N_7886,N_6067,N_6218);
xor U7887 (N_7887,N_6590,N_6141);
or U7888 (N_7888,N_6101,N_6555);
or U7889 (N_7889,N_6839,N_6760);
or U7890 (N_7890,N_6532,N_6296);
nand U7891 (N_7891,N_6845,N_6826);
xnor U7892 (N_7892,N_6680,N_6871);
nor U7893 (N_7893,N_6740,N_6647);
xor U7894 (N_7894,N_6964,N_6469);
nor U7895 (N_7895,N_6218,N_6296);
nand U7896 (N_7896,N_6948,N_6025);
or U7897 (N_7897,N_6012,N_6905);
nor U7898 (N_7898,N_6059,N_6512);
nand U7899 (N_7899,N_6558,N_6135);
and U7900 (N_7900,N_6955,N_6829);
or U7901 (N_7901,N_6058,N_6182);
nor U7902 (N_7902,N_6994,N_6232);
or U7903 (N_7903,N_6875,N_6446);
nor U7904 (N_7904,N_6885,N_6039);
nand U7905 (N_7905,N_6899,N_6763);
or U7906 (N_7906,N_6553,N_6258);
and U7907 (N_7907,N_6483,N_6813);
xor U7908 (N_7908,N_6012,N_6510);
or U7909 (N_7909,N_6301,N_6034);
nor U7910 (N_7910,N_6309,N_6671);
nand U7911 (N_7911,N_6021,N_6014);
nor U7912 (N_7912,N_6895,N_6460);
and U7913 (N_7913,N_6694,N_6348);
and U7914 (N_7914,N_6769,N_6525);
and U7915 (N_7915,N_6238,N_6916);
nand U7916 (N_7916,N_6295,N_6135);
nand U7917 (N_7917,N_6022,N_6121);
xor U7918 (N_7918,N_6948,N_6297);
nand U7919 (N_7919,N_6335,N_6045);
or U7920 (N_7920,N_6263,N_6362);
nor U7921 (N_7921,N_6256,N_6493);
or U7922 (N_7922,N_6278,N_6178);
xnor U7923 (N_7923,N_6246,N_6985);
and U7924 (N_7924,N_6967,N_6760);
nand U7925 (N_7925,N_6445,N_6295);
or U7926 (N_7926,N_6506,N_6560);
nor U7927 (N_7927,N_6043,N_6763);
or U7928 (N_7928,N_6478,N_6751);
xnor U7929 (N_7929,N_6115,N_6521);
and U7930 (N_7930,N_6788,N_6994);
and U7931 (N_7931,N_6923,N_6061);
or U7932 (N_7932,N_6541,N_6874);
nand U7933 (N_7933,N_6824,N_6591);
nand U7934 (N_7934,N_6414,N_6916);
nand U7935 (N_7935,N_6287,N_6303);
xor U7936 (N_7936,N_6319,N_6583);
nand U7937 (N_7937,N_6635,N_6740);
and U7938 (N_7938,N_6238,N_6580);
nor U7939 (N_7939,N_6323,N_6456);
or U7940 (N_7940,N_6160,N_6768);
xor U7941 (N_7941,N_6986,N_6962);
nand U7942 (N_7942,N_6638,N_6481);
nor U7943 (N_7943,N_6671,N_6344);
nand U7944 (N_7944,N_6191,N_6520);
nand U7945 (N_7945,N_6949,N_6024);
nor U7946 (N_7946,N_6846,N_6684);
and U7947 (N_7947,N_6135,N_6415);
nor U7948 (N_7948,N_6398,N_6985);
xor U7949 (N_7949,N_6666,N_6396);
xnor U7950 (N_7950,N_6723,N_6326);
nor U7951 (N_7951,N_6236,N_6203);
nand U7952 (N_7952,N_6653,N_6802);
nor U7953 (N_7953,N_6105,N_6378);
and U7954 (N_7954,N_6068,N_6816);
or U7955 (N_7955,N_6795,N_6111);
and U7956 (N_7956,N_6021,N_6994);
xnor U7957 (N_7957,N_6170,N_6260);
or U7958 (N_7958,N_6268,N_6918);
or U7959 (N_7959,N_6113,N_6094);
and U7960 (N_7960,N_6213,N_6339);
or U7961 (N_7961,N_6043,N_6961);
nand U7962 (N_7962,N_6116,N_6740);
nor U7963 (N_7963,N_6970,N_6011);
nor U7964 (N_7964,N_6364,N_6662);
nor U7965 (N_7965,N_6722,N_6676);
nand U7966 (N_7966,N_6317,N_6333);
or U7967 (N_7967,N_6774,N_6343);
or U7968 (N_7968,N_6721,N_6760);
nand U7969 (N_7969,N_6790,N_6755);
nor U7970 (N_7970,N_6464,N_6326);
xor U7971 (N_7971,N_6841,N_6028);
or U7972 (N_7972,N_6092,N_6272);
xnor U7973 (N_7973,N_6582,N_6446);
nor U7974 (N_7974,N_6087,N_6046);
nand U7975 (N_7975,N_6435,N_6616);
or U7976 (N_7976,N_6217,N_6305);
nand U7977 (N_7977,N_6114,N_6334);
and U7978 (N_7978,N_6044,N_6972);
xor U7979 (N_7979,N_6940,N_6499);
nor U7980 (N_7980,N_6221,N_6084);
or U7981 (N_7981,N_6496,N_6871);
nand U7982 (N_7982,N_6817,N_6107);
nand U7983 (N_7983,N_6304,N_6174);
or U7984 (N_7984,N_6128,N_6575);
or U7985 (N_7985,N_6124,N_6552);
nor U7986 (N_7986,N_6287,N_6627);
xor U7987 (N_7987,N_6144,N_6544);
xnor U7988 (N_7988,N_6800,N_6419);
or U7989 (N_7989,N_6642,N_6664);
and U7990 (N_7990,N_6197,N_6193);
nand U7991 (N_7991,N_6680,N_6210);
or U7992 (N_7992,N_6101,N_6777);
or U7993 (N_7993,N_6226,N_6867);
and U7994 (N_7994,N_6602,N_6807);
xor U7995 (N_7995,N_6614,N_6583);
or U7996 (N_7996,N_6836,N_6018);
nand U7997 (N_7997,N_6173,N_6423);
nor U7998 (N_7998,N_6726,N_6261);
and U7999 (N_7999,N_6289,N_6493);
nand U8000 (N_8000,N_7046,N_7528);
and U8001 (N_8001,N_7229,N_7183);
and U8002 (N_8002,N_7757,N_7732);
nor U8003 (N_8003,N_7271,N_7615);
nor U8004 (N_8004,N_7403,N_7614);
and U8005 (N_8005,N_7177,N_7690);
or U8006 (N_8006,N_7034,N_7659);
nor U8007 (N_8007,N_7423,N_7079);
nor U8008 (N_8008,N_7936,N_7838);
nor U8009 (N_8009,N_7344,N_7716);
and U8010 (N_8010,N_7182,N_7485);
nor U8011 (N_8011,N_7374,N_7415);
or U8012 (N_8012,N_7579,N_7536);
xnor U8013 (N_8013,N_7147,N_7882);
and U8014 (N_8014,N_7026,N_7376);
xor U8015 (N_8015,N_7245,N_7860);
nor U8016 (N_8016,N_7808,N_7259);
nor U8017 (N_8017,N_7653,N_7152);
or U8018 (N_8018,N_7915,N_7181);
or U8019 (N_8019,N_7360,N_7404);
nor U8020 (N_8020,N_7981,N_7512);
and U8021 (N_8021,N_7207,N_7749);
nor U8022 (N_8022,N_7569,N_7684);
or U8023 (N_8023,N_7622,N_7924);
or U8024 (N_8024,N_7298,N_7371);
xnor U8025 (N_8025,N_7351,N_7879);
or U8026 (N_8026,N_7567,N_7267);
nand U8027 (N_8027,N_7115,N_7347);
xnor U8028 (N_8028,N_7580,N_7297);
nor U8029 (N_8029,N_7209,N_7912);
nand U8030 (N_8030,N_7167,N_7558);
and U8031 (N_8031,N_7178,N_7726);
xor U8032 (N_8032,N_7102,N_7332);
nor U8033 (N_8033,N_7846,N_7644);
and U8034 (N_8034,N_7392,N_7244);
xnor U8035 (N_8035,N_7434,N_7414);
nor U8036 (N_8036,N_7138,N_7765);
and U8037 (N_8037,N_7467,N_7055);
xnor U8038 (N_8038,N_7847,N_7497);
xnor U8039 (N_8039,N_7225,N_7288);
xor U8040 (N_8040,N_7907,N_7424);
or U8041 (N_8041,N_7294,N_7247);
nand U8042 (N_8042,N_7545,N_7352);
xor U8043 (N_8043,N_7648,N_7903);
and U8044 (N_8044,N_7228,N_7979);
xnor U8045 (N_8045,N_7353,N_7672);
or U8046 (N_8046,N_7469,N_7830);
xor U8047 (N_8047,N_7557,N_7792);
or U8048 (N_8048,N_7998,N_7215);
or U8049 (N_8049,N_7880,N_7354);
or U8050 (N_8050,N_7463,N_7108);
and U8051 (N_8051,N_7511,N_7693);
xnor U8052 (N_8052,N_7285,N_7787);
and U8053 (N_8053,N_7211,N_7823);
xnor U8054 (N_8054,N_7443,N_7649);
nor U8055 (N_8055,N_7427,N_7238);
or U8056 (N_8056,N_7118,N_7123);
nand U8057 (N_8057,N_7121,N_7277);
and U8058 (N_8058,N_7893,N_7875);
xnor U8059 (N_8059,N_7717,N_7296);
and U8060 (N_8060,N_7196,N_7212);
nor U8061 (N_8061,N_7052,N_7180);
or U8062 (N_8062,N_7368,N_7170);
nor U8063 (N_8063,N_7464,N_7542);
nand U8064 (N_8064,N_7494,N_7287);
nand U8065 (N_8065,N_7074,N_7521);
nor U8066 (N_8066,N_7194,N_7772);
and U8067 (N_8067,N_7411,N_7987);
xnor U8068 (N_8068,N_7687,N_7728);
xor U8069 (N_8069,N_7894,N_7016);
or U8070 (N_8070,N_7933,N_7375);
xnor U8071 (N_8071,N_7843,N_7759);
nor U8072 (N_8072,N_7793,N_7361);
nor U8073 (N_8073,N_7175,N_7327);
nand U8074 (N_8074,N_7665,N_7931);
and U8075 (N_8075,N_7852,N_7646);
and U8076 (N_8076,N_7989,N_7002);
nand U8077 (N_8077,N_7281,N_7145);
and U8078 (N_8078,N_7543,N_7519);
nand U8079 (N_8079,N_7509,N_7030);
nor U8080 (N_8080,N_7642,N_7635);
and U8081 (N_8081,N_7734,N_7518);
or U8082 (N_8082,N_7921,N_7533);
or U8083 (N_8083,N_7539,N_7025);
or U8084 (N_8084,N_7286,N_7553);
or U8085 (N_8085,N_7559,N_7746);
or U8086 (N_8086,N_7675,N_7794);
nand U8087 (N_8087,N_7337,N_7457);
and U8088 (N_8088,N_7663,N_7962);
and U8089 (N_8089,N_7205,N_7389);
and U8090 (N_8090,N_7428,N_7733);
xnor U8091 (N_8091,N_7791,N_7061);
nor U8092 (N_8092,N_7764,N_7397);
and U8093 (N_8093,N_7219,N_7527);
nand U8094 (N_8094,N_7010,N_7340);
nand U8095 (N_8095,N_7314,N_7012);
or U8096 (N_8096,N_7949,N_7249);
or U8097 (N_8097,N_7032,N_7654);
xor U8098 (N_8098,N_7839,N_7199);
or U8099 (N_8099,N_7942,N_7508);
xor U8100 (N_8100,N_7948,N_7097);
nor U8101 (N_8101,N_7813,N_7562);
nor U8102 (N_8102,N_7279,N_7187);
xnor U8103 (N_8103,N_7163,N_7722);
nor U8104 (N_8104,N_7956,N_7438);
and U8105 (N_8105,N_7982,N_7947);
or U8106 (N_8106,N_7779,N_7385);
or U8107 (N_8107,N_7645,N_7867);
nor U8108 (N_8108,N_7240,N_7261);
xnor U8109 (N_8109,N_7117,N_7554);
and U8110 (N_8110,N_7643,N_7574);
or U8111 (N_8111,N_7017,N_7439);
xnor U8112 (N_8112,N_7070,N_7520);
nand U8113 (N_8113,N_7076,N_7381);
nor U8114 (N_8114,N_7563,N_7627);
and U8115 (N_8115,N_7999,N_7022);
nor U8116 (N_8116,N_7141,N_7262);
nand U8117 (N_8117,N_7573,N_7695);
xor U8118 (N_8118,N_7977,N_7328);
and U8119 (N_8119,N_7590,N_7681);
and U8120 (N_8120,N_7253,N_7930);
nand U8121 (N_8121,N_7561,N_7005);
nand U8122 (N_8122,N_7081,N_7243);
or U8123 (N_8123,N_7971,N_7383);
or U8124 (N_8124,N_7172,N_7831);
xor U8125 (N_8125,N_7782,N_7738);
nor U8126 (N_8126,N_7700,N_7587);
nand U8127 (N_8127,N_7384,N_7284);
nor U8128 (N_8128,N_7668,N_7278);
or U8129 (N_8129,N_7448,N_7776);
or U8130 (N_8130,N_7318,N_7682);
or U8131 (N_8131,N_7471,N_7293);
nor U8132 (N_8132,N_7817,N_7393);
nor U8133 (N_8133,N_7719,N_7869);
and U8134 (N_8134,N_7781,N_7596);
nand U8135 (N_8135,N_7116,N_7767);
or U8136 (N_8136,N_7067,N_7300);
xor U8137 (N_8137,N_7689,N_7953);
nor U8138 (N_8138,N_7083,N_7446);
nand U8139 (N_8139,N_7832,N_7641);
xor U8140 (N_8140,N_7816,N_7904);
or U8141 (N_8141,N_7315,N_7686);
nor U8142 (N_8142,N_7110,N_7727);
xor U8143 (N_8143,N_7378,N_7593);
nor U8144 (N_8144,N_7242,N_7203);
nor U8145 (N_8145,N_7217,N_7739);
xor U8146 (N_8146,N_7698,N_7221);
nor U8147 (N_8147,N_7155,N_7822);
nand U8148 (N_8148,N_7068,N_7410);
xor U8149 (N_8149,N_7537,N_7866);
nand U8150 (N_8150,N_7946,N_7650);
nor U8151 (N_8151,N_7507,N_7872);
xnor U8152 (N_8152,N_7707,N_7576);
or U8153 (N_8153,N_7131,N_7608);
and U8154 (N_8154,N_7906,N_7958);
nand U8155 (N_8155,N_7699,N_7185);
xnor U8156 (N_8156,N_7692,N_7619);
xnor U8157 (N_8157,N_7120,N_7861);
nand U8158 (N_8158,N_7575,N_7900);
xor U8159 (N_8159,N_7156,N_7235);
and U8160 (N_8160,N_7640,N_7339);
and U8161 (N_8161,N_7623,N_7957);
nand U8162 (N_8162,N_7320,N_7134);
or U8163 (N_8163,N_7685,N_7132);
xnor U8164 (N_8164,N_7701,N_7041);
nor U8165 (N_8165,N_7112,N_7342);
nand U8166 (N_8166,N_7788,N_7369);
nand U8167 (N_8167,N_7317,N_7283);
and U8168 (N_8168,N_7015,N_7011);
and U8169 (N_8169,N_7054,N_7826);
nand U8170 (N_8170,N_7657,N_7829);
nor U8171 (N_8171,N_7268,N_7988);
nor U8172 (N_8172,N_7819,N_7548);
nand U8173 (N_8173,N_7600,N_7835);
and U8174 (N_8174,N_7963,N_7857);
xor U8175 (N_8175,N_7892,N_7925);
and U8176 (N_8176,N_7720,N_7150);
and U8177 (N_8177,N_7673,N_7955);
or U8178 (N_8178,N_7555,N_7127);
nor U8179 (N_8179,N_7671,N_7472);
nor U8180 (N_8180,N_7790,N_7263);
xor U8181 (N_8181,N_7935,N_7321);
nand U8182 (N_8182,N_7252,N_7395);
nor U8183 (N_8183,N_7871,N_7870);
and U8184 (N_8184,N_7616,N_7544);
and U8185 (N_8185,N_7876,N_7483);
or U8186 (N_8186,N_7095,N_7799);
xor U8187 (N_8187,N_7612,N_7997);
nor U8188 (N_8188,N_7858,N_7157);
nand U8189 (N_8189,N_7085,N_7394);
xor U8190 (N_8190,N_7639,N_7908);
or U8191 (N_8191,N_7996,N_7807);
xnor U8192 (N_8192,N_7809,N_7059);
nor U8193 (N_8193,N_7887,N_7431);
nand U8194 (N_8194,N_7168,N_7056);
and U8195 (N_8195,N_7018,N_7477);
and U8196 (N_8196,N_7230,N_7609);
and U8197 (N_8197,N_7223,N_7101);
or U8198 (N_8198,N_7160,N_7350);
nor U8199 (N_8199,N_7902,N_7753);
and U8200 (N_8200,N_7454,N_7552);
or U8201 (N_8201,N_7966,N_7938);
and U8202 (N_8202,N_7125,N_7824);
xnor U8203 (N_8203,N_7868,N_7578);
and U8204 (N_8204,N_7197,N_7346);
and U8205 (N_8205,N_7628,N_7096);
or U8206 (N_8206,N_7380,N_7401);
and U8207 (N_8207,N_7149,N_7420);
and U8208 (N_8208,N_7250,N_7091);
and U8209 (N_8209,N_7198,N_7571);
nor U8210 (N_8210,N_7304,N_7677);
or U8211 (N_8211,N_7432,N_7007);
or U8212 (N_8212,N_7363,N_7481);
and U8213 (N_8213,N_7541,N_7724);
xnor U8214 (N_8214,N_7031,N_7291);
xnor U8215 (N_8215,N_7975,N_7331);
and U8216 (N_8216,N_7128,N_7610);
xor U8217 (N_8217,N_7430,N_7366);
nand U8218 (N_8218,N_7456,N_7001);
or U8219 (N_8219,N_7305,N_7918);
or U8220 (N_8220,N_7451,N_7206);
nand U8221 (N_8221,N_7029,N_7744);
and U8222 (N_8222,N_7992,N_7549);
nand U8223 (N_8223,N_7402,N_7784);
xor U8224 (N_8224,N_7064,N_7863);
or U8225 (N_8225,N_7633,N_7773);
and U8226 (N_8226,N_7489,N_7986);
xor U8227 (N_8227,N_7154,N_7950);
and U8228 (N_8228,N_7421,N_7737);
nand U8229 (N_8229,N_7660,N_7877);
nor U8230 (N_8230,N_7522,N_7714);
or U8231 (N_8231,N_7934,N_7943);
nor U8232 (N_8232,N_7967,N_7124);
and U8233 (N_8233,N_7637,N_7264);
and U8234 (N_8234,N_7103,N_7873);
nor U8235 (N_8235,N_7276,N_7445);
nor U8236 (N_8236,N_7334,N_7043);
xor U8237 (N_8237,N_7422,N_7683);
xor U8238 (N_8238,N_7752,N_7195);
and U8239 (N_8239,N_7617,N_7591);
and U8240 (N_8240,N_7329,N_7704);
nand U8241 (N_8241,N_7778,N_7419);
nand U8242 (N_8242,N_7504,N_7362);
or U8243 (N_8243,N_7038,N_7258);
nand U8244 (N_8244,N_7179,N_7437);
and U8245 (N_8245,N_7308,N_7336);
nand U8246 (N_8246,N_7510,N_7820);
nor U8247 (N_8247,N_7801,N_7019);
and U8248 (N_8248,N_7176,N_7740);
nor U8249 (N_8249,N_7592,N_7771);
nand U8250 (N_8250,N_7670,N_7540);
nand U8251 (N_8251,N_7914,N_7234);
nor U8252 (N_8252,N_7406,N_7917);
xor U8253 (N_8253,N_7078,N_7983);
nor U8254 (N_8254,N_7532,N_7324);
or U8255 (N_8255,N_7881,N_7488);
nor U8256 (N_8256,N_7845,N_7222);
nor U8257 (N_8257,N_7850,N_7502);
xor U8258 (N_8258,N_7564,N_7239);
nor U8259 (N_8259,N_7028,N_7373);
xnor U8260 (N_8260,N_7100,N_7390);
nor U8261 (N_8261,N_7530,N_7503);
nor U8262 (N_8262,N_7656,N_7306);
xnor U8263 (N_8263,N_7629,N_7758);
xor U8264 (N_8264,N_7595,N_7516);
nand U8265 (N_8265,N_7444,N_7452);
or U8266 (N_8266,N_7429,N_7498);
or U8267 (N_8267,N_7747,N_7370);
nand U8268 (N_8268,N_7715,N_7275);
nand U8269 (N_8269,N_7073,N_7137);
xnor U8270 (N_8270,N_7224,N_7743);
nor U8271 (N_8271,N_7534,N_7400);
nor U8272 (N_8272,N_7135,N_7634);
nor U8273 (N_8273,N_7589,N_7486);
nor U8274 (N_8274,N_7356,N_7084);
nand U8275 (N_8275,N_7796,N_7413);
and U8276 (N_8276,N_7696,N_7333);
nand U8277 (N_8277,N_7661,N_7805);
nor U8278 (N_8278,N_7674,N_7923);
and U8279 (N_8279,N_7077,N_7804);
xnor U8280 (N_8280,N_7256,N_7775);
xnor U8281 (N_8281,N_7251,N_7289);
nor U8282 (N_8282,N_7647,N_7878);
or U8283 (N_8283,N_7531,N_7789);
nand U8284 (N_8284,N_7736,N_7037);
nor U8285 (N_8285,N_7898,N_7080);
nor U8286 (N_8286,N_7325,N_7470);
xnor U8287 (N_8287,N_7468,N_7349);
nor U8288 (N_8288,N_7377,N_7697);
and U8289 (N_8289,N_7322,N_7087);
nand U8290 (N_8290,N_7144,N_7856);
or U8291 (N_8291,N_7550,N_7785);
nor U8292 (N_8292,N_7895,N_7844);
and U8293 (N_8293,N_7780,N_7425);
xnor U8294 (N_8294,N_7009,N_7114);
xnor U8295 (N_8295,N_7761,N_7260);
nor U8296 (N_8296,N_7631,N_7802);
and U8297 (N_8297,N_7313,N_7756);
and U8298 (N_8298,N_7597,N_7940);
or U8299 (N_8299,N_7113,N_7514);
nor U8300 (N_8300,N_7409,N_7777);
and U8301 (N_8301,N_7754,N_7570);
xor U8302 (N_8302,N_7216,N_7237);
and U8303 (N_8303,N_7526,N_7301);
or U8304 (N_8304,N_7712,N_7556);
nand U8305 (N_8305,N_7506,N_7006);
and U8306 (N_8306,N_7797,N_7048);
nor U8307 (N_8307,N_7505,N_7500);
and U8308 (N_8308,N_7226,N_7618);
xor U8309 (N_8309,N_7770,N_7093);
nor U8310 (N_8310,N_7343,N_7399);
and U8311 (N_8311,N_7841,N_7270);
or U8312 (N_8312,N_7466,N_7937);
nor U8313 (N_8313,N_7105,N_7326);
and U8314 (N_8314,N_7063,N_7786);
nor U8315 (N_8315,N_7450,N_7236);
xor U8316 (N_8316,N_7365,N_7932);
nand U8317 (N_8317,N_7825,N_7960);
nand U8318 (N_8318,N_7538,N_7513);
nor U8319 (N_8319,N_7367,N_7441);
and U8320 (N_8320,N_7458,N_7435);
xor U8321 (N_8321,N_7227,N_7192);
and U8322 (N_8322,N_7920,N_7969);
and U8323 (N_8323,N_7952,N_7638);
or U8324 (N_8324,N_7964,N_7899);
nand U8325 (N_8325,N_7694,N_7651);
or U8326 (N_8326,N_7040,N_7072);
or U8327 (N_8327,N_7926,N_7916);
xor U8328 (N_8328,N_7711,N_7652);
xor U8329 (N_8329,N_7584,N_7929);
nor U8330 (N_8330,N_7581,N_7345);
nand U8331 (N_8331,N_7042,N_7834);
nor U8332 (N_8332,N_7848,N_7143);
and U8333 (N_8333,N_7515,N_7828);
and U8334 (N_8334,N_7763,N_7136);
xnor U8335 (N_8335,N_7594,N_7440);
nand U8336 (N_8336,N_7171,N_7951);
nand U8337 (N_8337,N_7849,N_7139);
nor U8338 (N_8338,N_7184,N_7233);
xor U8339 (N_8339,N_7082,N_7751);
and U8340 (N_8340,N_7529,N_7388);
xor U8341 (N_8341,N_7173,N_7525);
xnor U8342 (N_8342,N_7624,N_7416);
xor U8343 (N_8343,N_7330,N_7161);
or U8344 (N_8344,N_7050,N_7044);
or U8345 (N_8345,N_7473,N_7023);
or U8346 (N_8346,N_7910,N_7436);
nand U8347 (N_8347,N_7153,N_7968);
or U8348 (N_8348,N_7057,N_7658);
nor U8349 (N_8349,N_7386,N_7051);
or U8350 (N_8350,N_7919,N_7970);
or U8351 (N_8351,N_7299,N_7391);
xor U8352 (N_8352,N_7387,N_7396);
nand U8353 (N_8353,N_7680,N_7210);
nand U8354 (N_8354,N_7755,N_7107);
or U8355 (N_8355,N_7257,N_7295);
or U8356 (N_8356,N_7547,N_7664);
xor U8357 (N_8357,N_7418,N_7109);
nand U8358 (N_8358,N_7478,N_7027);
nand U8359 (N_8359,N_7142,N_7162);
nor U8360 (N_8360,N_7604,N_7071);
xnor U8361 (N_8361,N_7146,N_7821);
nand U8362 (N_8362,N_7060,N_7837);
or U8363 (N_8363,N_7721,N_7311);
nand U8364 (N_8364,N_7985,N_7836);
nand U8365 (N_8365,N_7408,N_7723);
xor U8366 (N_8366,N_7667,N_7959);
and U8367 (N_8367,N_7220,N_7620);
xor U8368 (N_8368,N_7901,N_7272);
and U8369 (N_8369,N_7282,N_7407);
nand U8370 (N_8370,N_7292,N_7523);
and U8371 (N_8371,N_7735,N_7524);
and U8372 (N_8372,N_7455,N_7165);
nand U8373 (N_8373,N_7598,N_7566);
nand U8374 (N_8374,N_7862,N_7851);
nand U8375 (N_8375,N_7588,N_7214);
xnor U8376 (N_8376,N_7461,N_7750);
and U8377 (N_8377,N_7883,N_7748);
nor U8378 (N_8378,N_7274,N_7355);
nor U8379 (N_8379,N_7688,N_7200);
or U8380 (N_8380,N_7348,N_7889);
or U8381 (N_8381,N_7086,N_7607);
or U8382 (N_8382,N_7021,N_7874);
xor U8383 (N_8383,N_7290,N_7066);
and U8384 (N_8384,N_7405,N_7812);
nor U8385 (N_8385,N_7913,N_7583);
or U8386 (N_8386,N_7577,N_7246);
and U8387 (N_8387,N_7709,N_7491);
xor U8388 (N_8388,N_7191,N_7842);
nor U8389 (N_8389,N_7853,N_7104);
or U8390 (N_8390,N_7316,N_7742);
xor U8391 (N_8391,N_7762,N_7398);
and U8392 (N_8392,N_7897,N_7449);
or U8393 (N_8393,N_7495,N_7188);
or U8394 (N_8394,N_7599,N_7855);
xnor U8395 (N_8395,N_7961,N_7568);
nand U8396 (N_8396,N_7013,N_7859);
and U8397 (N_8397,N_7241,N_7335);
and U8398 (N_8398,N_7803,N_7075);
or U8399 (N_8399,N_7218,N_7159);
nand U8400 (N_8400,N_7815,N_7372);
nor U8401 (N_8401,N_7814,N_7703);
nand U8402 (N_8402,N_7586,N_7069);
xnor U8403 (N_8403,N_7280,N_7922);
and U8404 (N_8404,N_7730,N_7189);
nor U8405 (N_8405,N_7119,N_7885);
nand U8406 (N_8406,N_7731,N_7047);
and U8407 (N_8407,N_7725,N_7896);
xnor U8408 (N_8408,N_7613,N_7254);
or U8409 (N_8409,N_7800,N_7482);
and U8410 (N_8410,N_7053,N_7760);
or U8411 (N_8411,N_7944,N_7669);
nand U8412 (N_8412,N_7158,N_7148);
or U8413 (N_8413,N_7312,N_7140);
or U8414 (N_8414,N_7049,N_7480);
or U8415 (N_8415,N_7718,N_7357);
or U8416 (N_8416,N_7954,N_7662);
and U8417 (N_8417,N_7231,N_7106);
xnor U8418 (N_8418,N_7062,N_7601);
nand U8419 (N_8419,N_7585,N_7706);
nor U8420 (N_8420,N_7008,N_7768);
nor U8421 (N_8421,N_7169,N_7213);
or U8422 (N_8422,N_7323,N_7033);
and U8423 (N_8423,N_7493,N_7603);
nand U8424 (N_8424,N_7713,N_7766);
nor U8425 (N_8425,N_7827,N_7462);
nand U8426 (N_8426,N_7991,N_7941);
and U8427 (N_8427,N_7995,N_7993);
and U8428 (N_8428,N_7490,N_7965);
nor U8429 (N_8429,N_7465,N_7433);
xor U8430 (N_8430,N_7605,N_7572);
and U8431 (N_8431,N_7004,N_7678);
nand U8432 (N_8432,N_7978,N_7806);
xnor U8433 (N_8433,N_7499,N_7460);
or U8434 (N_8434,N_7891,N_7621);
nor U8435 (N_8435,N_7302,N_7338);
nand U8436 (N_8436,N_7492,N_7798);
xor U8437 (N_8437,N_7774,N_7865);
xor U8438 (N_8438,N_7984,N_7447);
nand U8439 (N_8439,N_7928,N_7783);
or U8440 (N_8440,N_7045,N_7269);
nand U8441 (N_8441,N_7098,N_7810);
and U8442 (N_8442,N_7412,N_7129);
nor U8443 (N_8443,N_7164,N_7560);
or U8444 (N_8444,N_7632,N_7020);
nor U8445 (N_8445,N_7174,N_7626);
or U8446 (N_8446,N_7795,N_7729);
and U8447 (N_8447,N_7190,N_7551);
xnor U8448 (N_8448,N_7702,N_7602);
nand U8449 (N_8449,N_7973,N_7636);
xnor U8450 (N_8450,N_7255,N_7840);
nor U8451 (N_8451,N_7201,N_7151);
nand U8452 (N_8452,N_7035,N_7442);
nor U8453 (N_8453,N_7310,N_7036);
nand U8454 (N_8454,N_7990,N_7939);
and U8455 (N_8455,N_7111,N_7024);
nand U8456 (N_8456,N_7625,N_7089);
nand U8457 (N_8457,N_7382,N_7122);
nand U8458 (N_8458,N_7501,N_7945);
xor U8459 (N_8459,N_7976,N_7058);
nor U8460 (N_8460,N_7705,N_7232);
nand U8461 (N_8461,N_7911,N_7359);
nor U8462 (N_8462,N_7606,N_7303);
nor U8463 (N_8463,N_7565,N_7833);
nor U8464 (N_8464,N_7090,N_7248);
xnor U8465 (N_8465,N_7341,N_7905);
or U8466 (N_8466,N_7204,N_7358);
nor U8467 (N_8467,N_7890,N_7884);
nand U8468 (N_8468,N_7487,N_7546);
xnor U8469 (N_8469,N_7474,N_7888);
xor U8470 (N_8470,N_7479,N_7092);
nand U8471 (N_8471,N_7186,N_7708);
xor U8472 (N_8472,N_7741,N_7691);
nand U8473 (N_8473,N_7273,N_7000);
or U8474 (N_8474,N_7611,N_7065);
and U8475 (N_8475,N_7417,N_7676);
nor U8476 (N_8476,N_7193,N_7854);
or U8477 (N_8477,N_7811,N_7769);
and U8478 (N_8478,N_7517,N_7133);
xor U8479 (N_8479,N_7014,N_7582);
xor U8480 (N_8480,N_7459,N_7094);
nand U8481 (N_8481,N_7994,N_7364);
xor U8482 (N_8482,N_7909,N_7655);
xnor U8483 (N_8483,N_7130,N_7972);
nor U8484 (N_8484,N_7099,N_7710);
xor U8485 (N_8485,N_7476,N_7679);
xor U8486 (N_8486,N_7309,N_7927);
xnor U8487 (N_8487,N_7475,N_7265);
and U8488 (N_8488,N_7484,N_7630);
xnor U8489 (N_8489,N_7535,N_7126);
or U8490 (N_8490,N_7864,N_7319);
nor U8491 (N_8491,N_7426,N_7208);
nor U8492 (N_8492,N_7166,N_7745);
xor U8493 (N_8493,N_7666,N_7974);
nor U8494 (N_8494,N_7266,N_7088);
xnor U8495 (N_8495,N_7453,N_7003);
xor U8496 (N_8496,N_7496,N_7039);
or U8497 (N_8497,N_7379,N_7818);
nand U8498 (N_8498,N_7202,N_7307);
xor U8499 (N_8499,N_7886,N_7980);
and U8500 (N_8500,N_7392,N_7837);
xnor U8501 (N_8501,N_7760,N_7401);
nor U8502 (N_8502,N_7036,N_7851);
nand U8503 (N_8503,N_7752,N_7228);
nor U8504 (N_8504,N_7251,N_7023);
and U8505 (N_8505,N_7729,N_7316);
or U8506 (N_8506,N_7741,N_7278);
nor U8507 (N_8507,N_7403,N_7747);
or U8508 (N_8508,N_7034,N_7962);
nand U8509 (N_8509,N_7718,N_7518);
xor U8510 (N_8510,N_7136,N_7355);
or U8511 (N_8511,N_7818,N_7653);
nor U8512 (N_8512,N_7197,N_7261);
or U8513 (N_8513,N_7078,N_7990);
nand U8514 (N_8514,N_7426,N_7537);
xnor U8515 (N_8515,N_7038,N_7316);
and U8516 (N_8516,N_7221,N_7875);
and U8517 (N_8517,N_7243,N_7313);
xnor U8518 (N_8518,N_7078,N_7804);
nand U8519 (N_8519,N_7900,N_7920);
and U8520 (N_8520,N_7804,N_7239);
or U8521 (N_8521,N_7713,N_7582);
xnor U8522 (N_8522,N_7096,N_7846);
nand U8523 (N_8523,N_7284,N_7713);
nand U8524 (N_8524,N_7456,N_7075);
or U8525 (N_8525,N_7013,N_7821);
xnor U8526 (N_8526,N_7741,N_7195);
xor U8527 (N_8527,N_7556,N_7214);
or U8528 (N_8528,N_7303,N_7998);
or U8529 (N_8529,N_7847,N_7246);
nor U8530 (N_8530,N_7528,N_7273);
and U8531 (N_8531,N_7580,N_7133);
nand U8532 (N_8532,N_7200,N_7731);
nor U8533 (N_8533,N_7009,N_7413);
nand U8534 (N_8534,N_7249,N_7696);
nor U8535 (N_8535,N_7747,N_7900);
and U8536 (N_8536,N_7614,N_7277);
or U8537 (N_8537,N_7095,N_7147);
and U8538 (N_8538,N_7733,N_7935);
or U8539 (N_8539,N_7895,N_7836);
and U8540 (N_8540,N_7382,N_7028);
or U8541 (N_8541,N_7194,N_7665);
and U8542 (N_8542,N_7554,N_7691);
nor U8543 (N_8543,N_7715,N_7906);
nor U8544 (N_8544,N_7757,N_7764);
xnor U8545 (N_8545,N_7788,N_7134);
or U8546 (N_8546,N_7461,N_7365);
xnor U8547 (N_8547,N_7664,N_7288);
nor U8548 (N_8548,N_7896,N_7479);
nand U8549 (N_8549,N_7967,N_7658);
xor U8550 (N_8550,N_7888,N_7783);
nor U8551 (N_8551,N_7669,N_7300);
xnor U8552 (N_8552,N_7741,N_7356);
xor U8553 (N_8553,N_7918,N_7109);
xor U8554 (N_8554,N_7954,N_7740);
xnor U8555 (N_8555,N_7614,N_7399);
nor U8556 (N_8556,N_7250,N_7950);
and U8557 (N_8557,N_7299,N_7161);
nor U8558 (N_8558,N_7218,N_7538);
and U8559 (N_8559,N_7547,N_7911);
xnor U8560 (N_8560,N_7244,N_7106);
nand U8561 (N_8561,N_7783,N_7125);
nor U8562 (N_8562,N_7968,N_7104);
xor U8563 (N_8563,N_7386,N_7763);
nor U8564 (N_8564,N_7859,N_7275);
or U8565 (N_8565,N_7570,N_7763);
nor U8566 (N_8566,N_7155,N_7952);
nand U8567 (N_8567,N_7204,N_7694);
xor U8568 (N_8568,N_7168,N_7405);
xnor U8569 (N_8569,N_7284,N_7427);
xor U8570 (N_8570,N_7382,N_7653);
nand U8571 (N_8571,N_7090,N_7790);
xnor U8572 (N_8572,N_7857,N_7327);
nand U8573 (N_8573,N_7517,N_7421);
nor U8574 (N_8574,N_7754,N_7947);
or U8575 (N_8575,N_7482,N_7784);
nor U8576 (N_8576,N_7085,N_7994);
nand U8577 (N_8577,N_7124,N_7680);
or U8578 (N_8578,N_7768,N_7940);
or U8579 (N_8579,N_7095,N_7442);
or U8580 (N_8580,N_7210,N_7700);
or U8581 (N_8581,N_7090,N_7308);
and U8582 (N_8582,N_7315,N_7116);
xnor U8583 (N_8583,N_7628,N_7741);
nand U8584 (N_8584,N_7232,N_7489);
nor U8585 (N_8585,N_7861,N_7402);
and U8586 (N_8586,N_7239,N_7630);
nand U8587 (N_8587,N_7669,N_7745);
nor U8588 (N_8588,N_7960,N_7013);
nand U8589 (N_8589,N_7079,N_7022);
and U8590 (N_8590,N_7806,N_7509);
nor U8591 (N_8591,N_7833,N_7599);
nor U8592 (N_8592,N_7925,N_7567);
nor U8593 (N_8593,N_7461,N_7696);
or U8594 (N_8594,N_7284,N_7821);
nand U8595 (N_8595,N_7743,N_7932);
or U8596 (N_8596,N_7939,N_7332);
xnor U8597 (N_8597,N_7124,N_7053);
nand U8598 (N_8598,N_7400,N_7515);
or U8599 (N_8599,N_7171,N_7421);
nand U8600 (N_8600,N_7921,N_7336);
and U8601 (N_8601,N_7887,N_7842);
and U8602 (N_8602,N_7519,N_7038);
nand U8603 (N_8603,N_7516,N_7914);
nand U8604 (N_8604,N_7650,N_7314);
nor U8605 (N_8605,N_7726,N_7825);
and U8606 (N_8606,N_7653,N_7299);
xnor U8607 (N_8607,N_7047,N_7805);
or U8608 (N_8608,N_7231,N_7602);
xnor U8609 (N_8609,N_7035,N_7904);
and U8610 (N_8610,N_7103,N_7478);
nor U8611 (N_8611,N_7524,N_7698);
or U8612 (N_8612,N_7193,N_7454);
xnor U8613 (N_8613,N_7173,N_7167);
or U8614 (N_8614,N_7321,N_7987);
and U8615 (N_8615,N_7139,N_7189);
or U8616 (N_8616,N_7252,N_7211);
nand U8617 (N_8617,N_7193,N_7040);
xor U8618 (N_8618,N_7485,N_7644);
xor U8619 (N_8619,N_7569,N_7185);
xnor U8620 (N_8620,N_7617,N_7186);
and U8621 (N_8621,N_7028,N_7854);
nor U8622 (N_8622,N_7056,N_7641);
xor U8623 (N_8623,N_7833,N_7316);
nand U8624 (N_8624,N_7533,N_7667);
nand U8625 (N_8625,N_7318,N_7246);
xor U8626 (N_8626,N_7932,N_7752);
and U8627 (N_8627,N_7724,N_7645);
xor U8628 (N_8628,N_7103,N_7973);
nor U8629 (N_8629,N_7007,N_7131);
and U8630 (N_8630,N_7436,N_7090);
or U8631 (N_8631,N_7834,N_7177);
nor U8632 (N_8632,N_7567,N_7726);
nand U8633 (N_8633,N_7879,N_7441);
or U8634 (N_8634,N_7299,N_7272);
and U8635 (N_8635,N_7489,N_7672);
and U8636 (N_8636,N_7847,N_7949);
nand U8637 (N_8637,N_7507,N_7480);
nand U8638 (N_8638,N_7047,N_7958);
or U8639 (N_8639,N_7365,N_7406);
nand U8640 (N_8640,N_7007,N_7295);
xnor U8641 (N_8641,N_7225,N_7751);
or U8642 (N_8642,N_7702,N_7650);
xor U8643 (N_8643,N_7760,N_7388);
nand U8644 (N_8644,N_7345,N_7612);
nor U8645 (N_8645,N_7160,N_7097);
or U8646 (N_8646,N_7309,N_7534);
nor U8647 (N_8647,N_7487,N_7130);
xnor U8648 (N_8648,N_7553,N_7247);
nand U8649 (N_8649,N_7303,N_7567);
nand U8650 (N_8650,N_7115,N_7061);
or U8651 (N_8651,N_7250,N_7135);
nand U8652 (N_8652,N_7113,N_7466);
nor U8653 (N_8653,N_7148,N_7474);
nor U8654 (N_8654,N_7405,N_7135);
nor U8655 (N_8655,N_7501,N_7951);
and U8656 (N_8656,N_7704,N_7174);
xor U8657 (N_8657,N_7080,N_7820);
nand U8658 (N_8658,N_7976,N_7061);
and U8659 (N_8659,N_7012,N_7516);
and U8660 (N_8660,N_7720,N_7951);
or U8661 (N_8661,N_7136,N_7183);
or U8662 (N_8662,N_7362,N_7396);
nor U8663 (N_8663,N_7600,N_7148);
or U8664 (N_8664,N_7210,N_7793);
nand U8665 (N_8665,N_7690,N_7039);
xor U8666 (N_8666,N_7622,N_7617);
and U8667 (N_8667,N_7003,N_7999);
and U8668 (N_8668,N_7722,N_7331);
nor U8669 (N_8669,N_7605,N_7690);
xnor U8670 (N_8670,N_7159,N_7037);
and U8671 (N_8671,N_7739,N_7736);
nand U8672 (N_8672,N_7696,N_7540);
and U8673 (N_8673,N_7261,N_7763);
xor U8674 (N_8674,N_7980,N_7889);
and U8675 (N_8675,N_7340,N_7004);
or U8676 (N_8676,N_7358,N_7354);
xor U8677 (N_8677,N_7785,N_7435);
nor U8678 (N_8678,N_7128,N_7661);
or U8679 (N_8679,N_7002,N_7382);
xnor U8680 (N_8680,N_7294,N_7504);
and U8681 (N_8681,N_7133,N_7457);
or U8682 (N_8682,N_7920,N_7203);
nor U8683 (N_8683,N_7470,N_7592);
xnor U8684 (N_8684,N_7662,N_7203);
or U8685 (N_8685,N_7971,N_7913);
or U8686 (N_8686,N_7500,N_7285);
or U8687 (N_8687,N_7451,N_7283);
nor U8688 (N_8688,N_7464,N_7525);
or U8689 (N_8689,N_7830,N_7159);
xor U8690 (N_8690,N_7343,N_7783);
and U8691 (N_8691,N_7378,N_7864);
nor U8692 (N_8692,N_7442,N_7939);
nand U8693 (N_8693,N_7113,N_7359);
or U8694 (N_8694,N_7874,N_7793);
xor U8695 (N_8695,N_7337,N_7123);
nor U8696 (N_8696,N_7709,N_7057);
nor U8697 (N_8697,N_7718,N_7811);
and U8698 (N_8698,N_7257,N_7816);
nand U8699 (N_8699,N_7267,N_7335);
nor U8700 (N_8700,N_7106,N_7501);
xnor U8701 (N_8701,N_7420,N_7361);
or U8702 (N_8702,N_7937,N_7119);
nor U8703 (N_8703,N_7140,N_7708);
or U8704 (N_8704,N_7140,N_7898);
nand U8705 (N_8705,N_7406,N_7836);
or U8706 (N_8706,N_7511,N_7946);
nor U8707 (N_8707,N_7157,N_7801);
or U8708 (N_8708,N_7782,N_7844);
nor U8709 (N_8709,N_7000,N_7252);
nand U8710 (N_8710,N_7978,N_7640);
or U8711 (N_8711,N_7540,N_7926);
or U8712 (N_8712,N_7633,N_7498);
nor U8713 (N_8713,N_7628,N_7359);
nand U8714 (N_8714,N_7588,N_7023);
xnor U8715 (N_8715,N_7142,N_7734);
xor U8716 (N_8716,N_7100,N_7693);
or U8717 (N_8717,N_7807,N_7135);
xnor U8718 (N_8718,N_7821,N_7260);
or U8719 (N_8719,N_7626,N_7526);
and U8720 (N_8720,N_7600,N_7908);
or U8721 (N_8721,N_7338,N_7491);
nor U8722 (N_8722,N_7951,N_7366);
or U8723 (N_8723,N_7822,N_7171);
nand U8724 (N_8724,N_7412,N_7960);
xnor U8725 (N_8725,N_7740,N_7248);
or U8726 (N_8726,N_7163,N_7359);
and U8727 (N_8727,N_7898,N_7688);
or U8728 (N_8728,N_7811,N_7287);
or U8729 (N_8729,N_7759,N_7813);
or U8730 (N_8730,N_7210,N_7354);
or U8731 (N_8731,N_7150,N_7380);
nand U8732 (N_8732,N_7750,N_7833);
or U8733 (N_8733,N_7637,N_7550);
and U8734 (N_8734,N_7423,N_7773);
nand U8735 (N_8735,N_7852,N_7848);
nand U8736 (N_8736,N_7847,N_7791);
xor U8737 (N_8737,N_7612,N_7710);
nor U8738 (N_8738,N_7289,N_7655);
or U8739 (N_8739,N_7429,N_7923);
nor U8740 (N_8740,N_7596,N_7187);
and U8741 (N_8741,N_7930,N_7074);
nand U8742 (N_8742,N_7773,N_7052);
or U8743 (N_8743,N_7471,N_7545);
xor U8744 (N_8744,N_7355,N_7382);
or U8745 (N_8745,N_7761,N_7228);
and U8746 (N_8746,N_7631,N_7409);
or U8747 (N_8747,N_7360,N_7846);
xnor U8748 (N_8748,N_7901,N_7827);
nor U8749 (N_8749,N_7149,N_7380);
xnor U8750 (N_8750,N_7157,N_7431);
nand U8751 (N_8751,N_7062,N_7437);
and U8752 (N_8752,N_7436,N_7275);
or U8753 (N_8753,N_7658,N_7188);
xor U8754 (N_8754,N_7273,N_7600);
or U8755 (N_8755,N_7032,N_7980);
and U8756 (N_8756,N_7038,N_7208);
or U8757 (N_8757,N_7515,N_7725);
or U8758 (N_8758,N_7721,N_7173);
or U8759 (N_8759,N_7166,N_7991);
or U8760 (N_8760,N_7104,N_7513);
nor U8761 (N_8761,N_7551,N_7458);
nor U8762 (N_8762,N_7510,N_7110);
nand U8763 (N_8763,N_7884,N_7339);
and U8764 (N_8764,N_7178,N_7735);
or U8765 (N_8765,N_7284,N_7342);
xor U8766 (N_8766,N_7874,N_7660);
nand U8767 (N_8767,N_7079,N_7938);
nand U8768 (N_8768,N_7625,N_7798);
and U8769 (N_8769,N_7606,N_7285);
nand U8770 (N_8770,N_7442,N_7291);
nor U8771 (N_8771,N_7084,N_7675);
nand U8772 (N_8772,N_7123,N_7413);
and U8773 (N_8773,N_7648,N_7010);
nand U8774 (N_8774,N_7426,N_7467);
or U8775 (N_8775,N_7499,N_7593);
and U8776 (N_8776,N_7058,N_7866);
or U8777 (N_8777,N_7947,N_7814);
nor U8778 (N_8778,N_7240,N_7016);
nor U8779 (N_8779,N_7724,N_7626);
nand U8780 (N_8780,N_7521,N_7086);
xor U8781 (N_8781,N_7079,N_7290);
and U8782 (N_8782,N_7572,N_7335);
or U8783 (N_8783,N_7191,N_7376);
nor U8784 (N_8784,N_7973,N_7429);
nor U8785 (N_8785,N_7248,N_7997);
nor U8786 (N_8786,N_7866,N_7696);
or U8787 (N_8787,N_7719,N_7631);
nand U8788 (N_8788,N_7243,N_7673);
nand U8789 (N_8789,N_7129,N_7071);
or U8790 (N_8790,N_7229,N_7037);
xnor U8791 (N_8791,N_7252,N_7488);
nand U8792 (N_8792,N_7332,N_7797);
nor U8793 (N_8793,N_7055,N_7315);
or U8794 (N_8794,N_7991,N_7017);
xor U8795 (N_8795,N_7118,N_7025);
nand U8796 (N_8796,N_7972,N_7898);
and U8797 (N_8797,N_7299,N_7808);
nor U8798 (N_8798,N_7375,N_7081);
or U8799 (N_8799,N_7320,N_7372);
or U8800 (N_8800,N_7662,N_7455);
nand U8801 (N_8801,N_7750,N_7698);
nor U8802 (N_8802,N_7579,N_7352);
nor U8803 (N_8803,N_7181,N_7930);
xnor U8804 (N_8804,N_7113,N_7198);
nor U8805 (N_8805,N_7733,N_7720);
nor U8806 (N_8806,N_7044,N_7634);
xor U8807 (N_8807,N_7382,N_7221);
or U8808 (N_8808,N_7536,N_7273);
nor U8809 (N_8809,N_7783,N_7467);
nand U8810 (N_8810,N_7176,N_7465);
nand U8811 (N_8811,N_7468,N_7257);
xnor U8812 (N_8812,N_7548,N_7666);
nor U8813 (N_8813,N_7596,N_7151);
and U8814 (N_8814,N_7223,N_7483);
nor U8815 (N_8815,N_7879,N_7904);
xnor U8816 (N_8816,N_7241,N_7798);
or U8817 (N_8817,N_7988,N_7403);
or U8818 (N_8818,N_7544,N_7426);
nor U8819 (N_8819,N_7737,N_7538);
and U8820 (N_8820,N_7877,N_7348);
nor U8821 (N_8821,N_7901,N_7908);
or U8822 (N_8822,N_7885,N_7102);
nor U8823 (N_8823,N_7908,N_7284);
or U8824 (N_8824,N_7171,N_7565);
xor U8825 (N_8825,N_7050,N_7913);
nand U8826 (N_8826,N_7478,N_7556);
nor U8827 (N_8827,N_7498,N_7782);
or U8828 (N_8828,N_7848,N_7991);
xor U8829 (N_8829,N_7767,N_7599);
nand U8830 (N_8830,N_7123,N_7777);
nor U8831 (N_8831,N_7827,N_7431);
or U8832 (N_8832,N_7312,N_7464);
nand U8833 (N_8833,N_7475,N_7127);
and U8834 (N_8834,N_7018,N_7191);
xor U8835 (N_8835,N_7369,N_7901);
and U8836 (N_8836,N_7977,N_7664);
or U8837 (N_8837,N_7851,N_7024);
and U8838 (N_8838,N_7204,N_7765);
or U8839 (N_8839,N_7525,N_7121);
and U8840 (N_8840,N_7495,N_7609);
or U8841 (N_8841,N_7687,N_7567);
and U8842 (N_8842,N_7959,N_7123);
or U8843 (N_8843,N_7385,N_7118);
nor U8844 (N_8844,N_7624,N_7707);
nor U8845 (N_8845,N_7761,N_7353);
and U8846 (N_8846,N_7895,N_7397);
or U8847 (N_8847,N_7479,N_7004);
xnor U8848 (N_8848,N_7215,N_7015);
nor U8849 (N_8849,N_7890,N_7109);
or U8850 (N_8850,N_7121,N_7687);
xor U8851 (N_8851,N_7855,N_7648);
nor U8852 (N_8852,N_7213,N_7081);
xnor U8853 (N_8853,N_7979,N_7836);
nand U8854 (N_8854,N_7826,N_7557);
or U8855 (N_8855,N_7274,N_7177);
or U8856 (N_8856,N_7622,N_7268);
or U8857 (N_8857,N_7040,N_7101);
and U8858 (N_8858,N_7599,N_7513);
and U8859 (N_8859,N_7440,N_7055);
and U8860 (N_8860,N_7750,N_7276);
nor U8861 (N_8861,N_7848,N_7110);
or U8862 (N_8862,N_7071,N_7534);
xnor U8863 (N_8863,N_7297,N_7293);
or U8864 (N_8864,N_7853,N_7193);
or U8865 (N_8865,N_7698,N_7069);
nor U8866 (N_8866,N_7307,N_7186);
nor U8867 (N_8867,N_7271,N_7849);
and U8868 (N_8868,N_7742,N_7313);
and U8869 (N_8869,N_7394,N_7450);
nand U8870 (N_8870,N_7993,N_7779);
nand U8871 (N_8871,N_7748,N_7561);
nand U8872 (N_8872,N_7976,N_7585);
nor U8873 (N_8873,N_7444,N_7762);
xnor U8874 (N_8874,N_7906,N_7953);
or U8875 (N_8875,N_7268,N_7983);
nand U8876 (N_8876,N_7293,N_7910);
nor U8877 (N_8877,N_7273,N_7383);
nand U8878 (N_8878,N_7069,N_7539);
and U8879 (N_8879,N_7444,N_7167);
or U8880 (N_8880,N_7050,N_7134);
and U8881 (N_8881,N_7668,N_7877);
and U8882 (N_8882,N_7114,N_7932);
nor U8883 (N_8883,N_7646,N_7817);
xor U8884 (N_8884,N_7176,N_7528);
nand U8885 (N_8885,N_7427,N_7504);
xor U8886 (N_8886,N_7776,N_7378);
or U8887 (N_8887,N_7549,N_7376);
or U8888 (N_8888,N_7517,N_7341);
nor U8889 (N_8889,N_7843,N_7716);
xor U8890 (N_8890,N_7453,N_7566);
and U8891 (N_8891,N_7729,N_7382);
and U8892 (N_8892,N_7307,N_7554);
nand U8893 (N_8893,N_7436,N_7581);
or U8894 (N_8894,N_7740,N_7661);
nor U8895 (N_8895,N_7384,N_7864);
and U8896 (N_8896,N_7244,N_7911);
or U8897 (N_8897,N_7462,N_7914);
nor U8898 (N_8898,N_7736,N_7412);
or U8899 (N_8899,N_7667,N_7601);
or U8900 (N_8900,N_7355,N_7631);
xnor U8901 (N_8901,N_7654,N_7659);
nand U8902 (N_8902,N_7926,N_7504);
xor U8903 (N_8903,N_7000,N_7027);
nor U8904 (N_8904,N_7995,N_7928);
nor U8905 (N_8905,N_7806,N_7064);
or U8906 (N_8906,N_7017,N_7304);
nand U8907 (N_8907,N_7974,N_7159);
xnor U8908 (N_8908,N_7169,N_7202);
or U8909 (N_8909,N_7772,N_7294);
and U8910 (N_8910,N_7121,N_7718);
or U8911 (N_8911,N_7234,N_7461);
or U8912 (N_8912,N_7149,N_7446);
nand U8913 (N_8913,N_7324,N_7540);
nor U8914 (N_8914,N_7835,N_7253);
nor U8915 (N_8915,N_7924,N_7948);
and U8916 (N_8916,N_7741,N_7228);
nor U8917 (N_8917,N_7050,N_7898);
xor U8918 (N_8918,N_7013,N_7634);
nand U8919 (N_8919,N_7711,N_7834);
xnor U8920 (N_8920,N_7089,N_7306);
nand U8921 (N_8921,N_7583,N_7836);
and U8922 (N_8922,N_7651,N_7537);
or U8923 (N_8923,N_7854,N_7211);
nor U8924 (N_8924,N_7638,N_7161);
xor U8925 (N_8925,N_7154,N_7514);
and U8926 (N_8926,N_7196,N_7003);
nand U8927 (N_8927,N_7999,N_7127);
or U8928 (N_8928,N_7818,N_7004);
nor U8929 (N_8929,N_7709,N_7606);
nand U8930 (N_8930,N_7008,N_7353);
nand U8931 (N_8931,N_7876,N_7485);
or U8932 (N_8932,N_7285,N_7566);
nor U8933 (N_8933,N_7430,N_7469);
or U8934 (N_8934,N_7459,N_7181);
or U8935 (N_8935,N_7301,N_7635);
or U8936 (N_8936,N_7982,N_7403);
xor U8937 (N_8937,N_7706,N_7234);
or U8938 (N_8938,N_7587,N_7973);
xnor U8939 (N_8939,N_7863,N_7316);
or U8940 (N_8940,N_7178,N_7704);
nor U8941 (N_8941,N_7352,N_7892);
or U8942 (N_8942,N_7832,N_7130);
and U8943 (N_8943,N_7256,N_7092);
nor U8944 (N_8944,N_7123,N_7655);
nor U8945 (N_8945,N_7716,N_7876);
and U8946 (N_8946,N_7685,N_7631);
xor U8947 (N_8947,N_7817,N_7888);
nand U8948 (N_8948,N_7183,N_7860);
nor U8949 (N_8949,N_7698,N_7878);
xor U8950 (N_8950,N_7502,N_7879);
xnor U8951 (N_8951,N_7876,N_7785);
or U8952 (N_8952,N_7300,N_7725);
nand U8953 (N_8953,N_7617,N_7631);
or U8954 (N_8954,N_7199,N_7360);
xnor U8955 (N_8955,N_7600,N_7462);
xor U8956 (N_8956,N_7507,N_7681);
nand U8957 (N_8957,N_7215,N_7428);
xor U8958 (N_8958,N_7443,N_7535);
or U8959 (N_8959,N_7225,N_7271);
nor U8960 (N_8960,N_7260,N_7127);
nor U8961 (N_8961,N_7702,N_7833);
nor U8962 (N_8962,N_7238,N_7204);
and U8963 (N_8963,N_7596,N_7961);
and U8964 (N_8964,N_7154,N_7442);
nor U8965 (N_8965,N_7637,N_7374);
nand U8966 (N_8966,N_7435,N_7251);
nand U8967 (N_8967,N_7915,N_7091);
xnor U8968 (N_8968,N_7561,N_7230);
or U8969 (N_8969,N_7342,N_7320);
and U8970 (N_8970,N_7309,N_7561);
or U8971 (N_8971,N_7109,N_7402);
nor U8972 (N_8972,N_7513,N_7149);
or U8973 (N_8973,N_7097,N_7047);
nand U8974 (N_8974,N_7024,N_7980);
nor U8975 (N_8975,N_7946,N_7184);
xnor U8976 (N_8976,N_7797,N_7084);
nor U8977 (N_8977,N_7795,N_7754);
and U8978 (N_8978,N_7587,N_7920);
or U8979 (N_8979,N_7380,N_7454);
xnor U8980 (N_8980,N_7294,N_7450);
and U8981 (N_8981,N_7885,N_7359);
xor U8982 (N_8982,N_7955,N_7914);
nor U8983 (N_8983,N_7256,N_7337);
nor U8984 (N_8984,N_7251,N_7034);
and U8985 (N_8985,N_7405,N_7584);
or U8986 (N_8986,N_7243,N_7161);
or U8987 (N_8987,N_7650,N_7364);
and U8988 (N_8988,N_7897,N_7973);
nand U8989 (N_8989,N_7317,N_7640);
nor U8990 (N_8990,N_7529,N_7512);
nand U8991 (N_8991,N_7280,N_7255);
nand U8992 (N_8992,N_7919,N_7271);
or U8993 (N_8993,N_7411,N_7639);
xnor U8994 (N_8994,N_7366,N_7315);
nor U8995 (N_8995,N_7517,N_7638);
nor U8996 (N_8996,N_7688,N_7767);
nand U8997 (N_8997,N_7746,N_7969);
nand U8998 (N_8998,N_7969,N_7422);
nor U8999 (N_8999,N_7692,N_7491);
nand U9000 (N_9000,N_8155,N_8839);
xnor U9001 (N_9001,N_8660,N_8154);
nor U9002 (N_9002,N_8417,N_8787);
and U9003 (N_9003,N_8567,N_8906);
nand U9004 (N_9004,N_8962,N_8815);
xnor U9005 (N_9005,N_8497,N_8427);
or U9006 (N_9006,N_8079,N_8745);
nor U9007 (N_9007,N_8283,N_8621);
nor U9008 (N_9008,N_8960,N_8425);
or U9009 (N_9009,N_8101,N_8186);
nand U9010 (N_9010,N_8534,N_8844);
xnor U9011 (N_9011,N_8050,N_8359);
xor U9012 (N_9012,N_8580,N_8727);
and U9013 (N_9013,N_8366,N_8560);
or U9014 (N_9014,N_8975,N_8995);
and U9015 (N_9015,N_8742,N_8877);
nor U9016 (N_9016,N_8349,N_8119);
and U9017 (N_9017,N_8686,N_8615);
nand U9018 (N_9018,N_8765,N_8584);
and U9019 (N_9019,N_8950,N_8315);
nand U9020 (N_9020,N_8990,N_8077);
or U9021 (N_9021,N_8299,N_8099);
nor U9022 (N_9022,N_8360,N_8638);
nand U9023 (N_9023,N_8432,N_8625);
nand U9024 (N_9024,N_8460,N_8258);
and U9025 (N_9025,N_8313,N_8056);
xnor U9026 (N_9026,N_8536,N_8134);
or U9027 (N_9027,N_8164,N_8715);
xnor U9028 (N_9028,N_8256,N_8393);
and U9029 (N_9029,N_8949,N_8856);
nor U9030 (N_9030,N_8821,N_8792);
or U9031 (N_9031,N_8097,N_8306);
xnor U9032 (N_9032,N_8019,N_8448);
and U9033 (N_9033,N_8802,N_8798);
xnor U9034 (N_9034,N_8545,N_8649);
xor U9035 (N_9035,N_8233,N_8945);
xor U9036 (N_9036,N_8185,N_8923);
nor U9037 (N_9037,N_8200,N_8702);
or U9038 (N_9038,N_8531,N_8132);
nand U9039 (N_9039,N_8518,N_8231);
or U9040 (N_9040,N_8896,N_8805);
or U9041 (N_9041,N_8537,N_8958);
xnor U9042 (N_9042,N_8812,N_8407);
nand U9043 (N_9043,N_8522,N_8160);
xor U9044 (N_9044,N_8635,N_8043);
and U9045 (N_9045,N_8972,N_8287);
or U9046 (N_9046,N_8373,N_8936);
nand U9047 (N_9047,N_8281,N_8309);
xor U9048 (N_9048,N_8161,N_8398);
and U9049 (N_9049,N_8888,N_8098);
nand U9050 (N_9050,N_8706,N_8796);
nand U9051 (N_9051,N_8627,N_8644);
and U9052 (N_9052,N_8709,N_8198);
or U9053 (N_9053,N_8435,N_8211);
nor U9054 (N_9054,N_8314,N_8948);
and U9055 (N_9055,N_8140,N_8903);
or U9056 (N_9056,N_8130,N_8719);
nor U9057 (N_9057,N_8254,N_8403);
and U9058 (N_9058,N_8919,N_8981);
or U9059 (N_9059,N_8251,N_8933);
nor U9060 (N_9060,N_8540,N_8003);
nand U9061 (N_9061,N_8480,N_8380);
or U9062 (N_9062,N_8129,N_8870);
nand U9063 (N_9063,N_8110,N_8670);
or U9064 (N_9064,N_8645,N_8546);
xnor U9065 (N_9065,N_8671,N_8012);
or U9066 (N_9066,N_8769,N_8612);
xor U9067 (N_9067,N_8117,N_8004);
nand U9068 (N_9068,N_8467,N_8901);
or U9069 (N_9069,N_8152,N_8339);
and U9070 (N_9070,N_8147,N_8983);
and U9071 (N_9071,N_8951,N_8886);
xnor U9072 (N_9072,N_8109,N_8293);
or U9073 (N_9073,N_8663,N_8883);
and U9074 (N_9074,N_8298,N_8089);
xnor U9075 (N_9075,N_8102,N_8723);
nor U9076 (N_9076,N_8803,N_8630);
nand U9077 (N_9077,N_8464,N_8419);
or U9078 (N_9078,N_8711,N_8224);
and U9079 (N_9079,N_8956,N_8512);
and U9080 (N_9080,N_8178,N_8561);
nor U9081 (N_9081,N_8874,N_8639);
and U9082 (N_9082,N_8494,N_8850);
nand U9083 (N_9083,N_8086,N_8684);
nand U9084 (N_9084,N_8397,N_8613);
or U9085 (N_9085,N_8876,N_8107);
or U9086 (N_9086,N_8106,N_8409);
and U9087 (N_9087,N_8898,N_8405);
and U9088 (N_9088,N_8288,N_8520);
or U9089 (N_9089,N_8880,N_8559);
xor U9090 (N_9090,N_8875,N_8683);
xor U9091 (N_9091,N_8624,N_8761);
or U9092 (N_9092,N_8857,N_8925);
nand U9093 (N_9093,N_8291,N_8661);
or U9094 (N_9094,N_8666,N_8776);
or U9095 (N_9095,N_8731,N_8895);
and U9096 (N_9096,N_8368,N_8450);
xor U9097 (N_9097,N_8093,N_8087);
or U9098 (N_9098,N_8694,N_8230);
and U9099 (N_9099,N_8234,N_8810);
nor U9100 (N_9100,N_8966,N_8685);
and U9101 (N_9101,N_8263,N_8381);
nor U9102 (N_9102,N_8378,N_8357);
or U9103 (N_9103,N_8169,N_8626);
xnor U9104 (N_9104,N_8307,N_8817);
or U9105 (N_9105,N_8406,N_8979);
or U9106 (N_9106,N_8400,N_8150);
nand U9107 (N_9107,N_8597,N_8506);
nor U9108 (N_9108,N_8111,N_8245);
nor U9109 (N_9109,N_8005,N_8121);
or U9110 (N_9110,N_8328,N_8402);
or U9111 (N_9111,N_8565,N_8182);
nor U9112 (N_9112,N_8693,N_8734);
nor U9113 (N_9113,N_8066,N_8461);
nand U9114 (N_9114,N_8940,N_8992);
xnor U9115 (N_9115,N_8733,N_8551);
or U9116 (N_9116,N_8372,N_8415);
and U9117 (N_9117,N_8083,N_8327);
nor U9118 (N_9118,N_8801,N_8300);
nor U9119 (N_9119,N_8015,N_8146);
nand U9120 (N_9120,N_8773,N_8371);
nor U9121 (N_9121,N_8189,N_8569);
or U9122 (N_9122,N_8984,N_8541);
or U9123 (N_9123,N_8481,N_8302);
xnor U9124 (N_9124,N_8843,N_8595);
xnor U9125 (N_9125,N_8193,N_8241);
nor U9126 (N_9126,N_8814,N_8092);
xor U9127 (N_9127,N_8764,N_8500);
and U9128 (N_9128,N_8637,N_8775);
xor U9129 (N_9129,N_8548,N_8179);
and U9130 (N_9130,N_8934,N_8082);
or U9131 (N_9131,N_8633,N_8504);
and U9132 (N_9132,N_8355,N_8038);
nor U9133 (N_9133,N_8042,N_8159);
nand U9134 (N_9134,N_8701,N_8851);
nand U9135 (N_9135,N_8599,N_8552);
or U9136 (N_9136,N_8620,N_8730);
nor U9137 (N_9137,N_8205,N_8474);
and U9138 (N_9138,N_8413,N_8045);
and U9139 (N_9139,N_8112,N_8505);
nor U9140 (N_9140,N_8157,N_8104);
and U9141 (N_9141,N_8519,N_8310);
xnor U9142 (N_9142,N_8891,N_8404);
and U9143 (N_9143,N_8434,N_8369);
and U9144 (N_9144,N_8757,N_8301);
xnor U9145 (N_9145,N_8067,N_8203);
xnor U9146 (N_9146,N_8459,N_8037);
nand U9147 (N_9147,N_8980,N_8333);
or U9148 (N_9148,N_8214,N_8695);
xnor U9149 (N_9149,N_8652,N_8704);
xnor U9150 (N_9150,N_8503,N_8566);
nand U9151 (N_9151,N_8501,N_8705);
nor U9152 (N_9152,N_8549,N_8657);
and U9153 (N_9153,N_8384,N_8240);
nor U9154 (N_9154,N_8041,N_8879);
and U9155 (N_9155,N_8399,N_8837);
xor U9156 (N_9156,N_8659,N_8974);
and U9157 (N_9157,N_8768,N_8953);
nand U9158 (N_9158,N_8465,N_8232);
and U9159 (N_9159,N_8141,N_8353);
nand U9160 (N_9160,N_8676,N_8331);
xnor U9161 (N_9161,N_8887,N_8517);
nor U9162 (N_9162,N_8242,N_8064);
xor U9163 (N_9163,N_8462,N_8063);
or U9164 (N_9164,N_8847,N_8445);
xor U9165 (N_9165,N_8364,N_8148);
xnor U9166 (N_9166,N_8350,N_8912);
nor U9167 (N_9167,N_8323,N_8303);
and U9168 (N_9168,N_8866,N_8526);
and U9169 (N_9169,N_8678,N_8908);
xor U9170 (N_9170,N_8304,N_8859);
and U9171 (N_9171,N_8215,N_8721);
nand U9172 (N_9172,N_8662,N_8585);
and U9173 (N_9173,N_8564,N_8578);
nor U9174 (N_9174,N_8123,N_8894);
and U9175 (N_9175,N_8954,N_8818);
nand U9176 (N_9176,N_8910,N_8167);
nand U9177 (N_9177,N_8862,N_8216);
nand U9178 (N_9178,N_8763,N_8065);
or U9179 (N_9179,N_8834,N_8848);
and U9180 (N_9180,N_8691,N_8095);
xor U9181 (N_9181,N_8744,N_8884);
nand U9182 (N_9182,N_8292,N_8316);
nand U9183 (N_9183,N_8591,N_8618);
and U9184 (N_9184,N_8819,N_8790);
xor U9185 (N_9185,N_8555,N_8498);
nor U9186 (N_9186,N_8777,N_8736);
nand U9187 (N_9187,N_8478,N_8999);
nor U9188 (N_9188,N_8345,N_8139);
xor U9189 (N_9189,N_8424,N_8516);
and U9190 (N_9190,N_8458,N_8668);
xor U9191 (N_9191,N_8100,N_8690);
nand U9192 (N_9192,N_8664,N_8982);
or U9193 (N_9193,N_8493,N_8689);
or U9194 (N_9194,N_8680,N_8260);
and U9195 (N_9195,N_8062,N_8492);
xor U9196 (N_9196,N_8348,N_8563);
and U9197 (N_9197,N_8008,N_8539);
or U9198 (N_9198,N_8998,N_8344);
or U9199 (N_9199,N_8845,N_8971);
xnor U9200 (N_9200,N_8014,N_8320);
nor U9201 (N_9201,N_8718,N_8162);
nor U9202 (N_9202,N_8282,N_8988);
xor U9203 (N_9203,N_8249,N_8743);
nor U9204 (N_9204,N_8656,N_8437);
nor U9205 (N_9205,N_8396,N_8024);
nand U9206 (N_9206,N_8085,N_8277);
nand U9207 (N_9207,N_8643,N_8813);
xnor U9208 (N_9208,N_8330,N_8806);
or U9209 (N_9209,N_8917,N_8124);
nand U9210 (N_9210,N_8290,N_8515);
nor U9211 (N_9211,N_8025,N_8412);
and U9212 (N_9212,N_8527,N_8658);
or U9213 (N_9213,N_8881,N_8033);
nor U9214 (N_9214,N_8446,N_8408);
xor U9215 (N_9215,N_8379,N_8672);
nand U9216 (N_9216,N_8495,N_8909);
and U9217 (N_9217,N_8453,N_8236);
or U9218 (N_9218,N_8782,N_8700);
nor U9219 (N_9219,N_8809,N_8811);
nand U9220 (N_9220,N_8017,N_8210);
and U9221 (N_9221,N_8907,N_8554);
and U9222 (N_9222,N_8514,N_8778);
xor U9223 (N_9223,N_8825,N_8133);
or U9224 (N_9224,N_8994,N_8677);
nand U9225 (N_9225,N_8616,N_8284);
xnor U9226 (N_9226,N_8502,N_8737);
and U9227 (N_9227,N_8930,N_8352);
xnor U9228 (N_9228,N_8918,N_8867);
or U9229 (N_9229,N_8305,N_8755);
or U9230 (N_9230,N_8206,N_8795);
xnor U9231 (N_9231,N_8321,N_8385);
xnor U9232 (N_9232,N_8807,N_8028);
nor U9233 (N_9233,N_8108,N_8416);
nor U9234 (N_9234,N_8854,N_8929);
or U9235 (N_9235,N_8257,N_8196);
or U9236 (N_9236,N_8892,N_8222);
xnor U9237 (N_9237,N_8931,N_8275);
xor U9238 (N_9238,N_8319,N_8968);
nand U9239 (N_9239,N_8921,N_8893);
xnor U9240 (N_9240,N_8212,N_8529);
and U9241 (N_9241,N_8758,N_8034);
and U9242 (N_9242,N_8955,N_8836);
and U9243 (N_9243,N_8568,N_8596);
nand U9244 (N_9244,N_8278,N_8127);
xnor U9245 (N_9245,N_8872,N_8838);
nand U9246 (N_9246,N_8927,N_8080);
xor U9247 (N_9247,N_8528,N_8835);
or U9248 (N_9248,N_8970,N_8911);
nor U9249 (N_9249,N_8722,N_8963);
nand U9250 (N_9250,N_8606,N_8010);
xor U9251 (N_9251,N_8728,N_8588);
xnor U9252 (N_9252,N_8829,N_8675);
nand U9253 (N_9253,N_8830,N_8897);
and U9254 (N_9254,N_8267,N_8717);
or U9255 (N_9255,N_8439,N_8090);
or U9256 (N_9256,N_8128,N_8882);
and U9257 (N_9257,N_8174,N_8126);
xor U9258 (N_9258,N_8376,N_8036);
nand U9259 (N_9259,N_8197,N_8273);
and U9260 (N_9260,N_8105,N_8421);
and U9261 (N_9261,N_8928,N_8573);
nand U9262 (N_9262,N_8991,N_8272);
nor U9263 (N_9263,N_8674,N_8716);
or U9264 (N_9264,N_8032,N_8748);
or U9265 (N_9265,N_8158,N_8422);
or U9266 (N_9266,N_8786,N_8952);
nand U9267 (N_9267,N_8570,N_8482);
or U9268 (N_9268,N_8967,N_8058);
nand U9269 (N_9269,N_8899,N_8989);
nor U9270 (N_9270,N_8122,N_8131);
or U9271 (N_9271,N_8781,N_8508);
or U9272 (N_9272,N_8858,N_8617);
xor U9273 (N_9273,N_8873,N_8280);
xnor U9274 (N_9274,N_8833,N_8783);
nor U9275 (N_9275,N_8852,N_8070);
and U9276 (N_9276,N_8013,N_8423);
nor U9277 (N_9277,N_8871,N_8523);
nor U9278 (N_9278,N_8044,N_8039);
nor U9279 (N_9279,N_8828,N_8078);
nor U9280 (N_9280,N_8442,N_8285);
and U9281 (N_9281,N_8392,N_8239);
nand U9282 (N_9282,N_8227,N_8673);
nand U9283 (N_9283,N_8264,N_8754);
nand U9284 (N_9284,N_8027,N_8246);
or U9285 (N_9285,N_8749,N_8342);
nor U9286 (N_9286,N_8740,N_8204);
nand U9287 (N_9287,N_8978,N_8456);
xnor U9288 (N_9288,N_8430,N_8542);
xor U9289 (N_9289,N_8029,N_8746);
nor U9290 (N_9290,N_8387,N_8476);
nand U9291 (N_9291,N_8779,N_8286);
nor U9292 (N_9292,N_8634,N_8996);
nand U9293 (N_9293,N_8023,N_8395);
or U9294 (N_9294,N_8325,N_8985);
and U9295 (N_9295,N_8558,N_8472);
nand U9296 (N_9296,N_8855,N_8143);
or U9297 (N_9297,N_8006,N_8324);
and U9298 (N_9298,N_8347,N_8729);
and U9299 (N_9299,N_8863,N_8831);
nor U9300 (N_9300,N_8195,N_8488);
xor U9301 (N_9301,N_8521,N_8269);
nand U9302 (N_9302,N_8337,N_8900);
nor U9303 (N_9303,N_8173,N_8712);
nand U9304 (N_9304,N_8444,N_8221);
nand U9305 (N_9305,N_8669,N_8832);
xnor U9306 (N_9306,N_8218,N_8125);
or U9307 (N_9307,N_8804,N_8868);
nand U9308 (N_9308,N_8466,N_8594);
or U9309 (N_9309,N_8646,N_8068);
nand U9310 (N_9310,N_8361,N_8388);
xnor U9311 (N_9311,N_8581,N_8589);
xor U9312 (N_9312,N_8180,N_8496);
or U9313 (N_9313,N_8753,N_8391);
xor U9314 (N_9314,N_8153,N_8470);
or U9315 (N_9315,N_8961,N_8115);
or U9316 (N_9316,N_8270,N_8084);
xnor U9317 (N_9317,N_8438,N_8681);
or U9318 (N_9318,N_8279,N_8760);
nand U9319 (N_9319,N_8149,N_8553);
nand U9320 (N_9320,N_8394,N_8338);
or U9321 (N_9321,N_8688,N_8619);
or U9322 (N_9322,N_8904,N_8329);
or U9323 (N_9323,N_8969,N_8827);
xor U9324 (N_9324,N_8640,N_8145);
or U9325 (N_9325,N_8168,N_8650);
xnor U9326 (N_9326,N_8081,N_8808);
or U9327 (N_9327,N_8418,N_8060);
or U9328 (N_9328,N_8603,N_8046);
or U9329 (N_9329,N_8920,N_8454);
and U9330 (N_9330,N_8252,N_8411);
and U9331 (N_9331,N_8374,N_8053);
xnor U9332 (N_9332,N_8648,N_8433);
xor U9333 (N_9333,N_8294,N_8860);
nand U9334 (N_9334,N_8166,N_8049);
nor U9335 (N_9335,N_8274,N_8532);
xnor U9336 (N_9336,N_8605,N_8343);
xor U9337 (N_9337,N_8924,N_8601);
or U9338 (N_9338,N_8785,N_8118);
xnor U9339 (N_9339,N_8336,N_8171);
nor U9340 (N_9340,N_8295,N_8572);
or U9341 (N_9341,N_8370,N_8579);
xor U9342 (N_9342,N_8362,N_8363);
and U9343 (N_9343,N_8889,N_8946);
nand U9344 (N_9344,N_8271,N_8268);
and U9345 (N_9345,N_8944,N_8055);
and U9346 (N_9346,N_8312,N_8696);
or U9347 (N_9347,N_8199,N_8181);
nand U9348 (N_9348,N_8842,N_8987);
xnor U9349 (N_9349,N_8217,N_8047);
nand U9350 (N_9350,N_8018,N_8297);
xnor U9351 (N_9351,N_8582,N_8943);
and U9352 (N_9352,N_8219,N_8071);
or U9353 (N_9353,N_8020,N_8750);
or U9354 (N_9354,N_8608,N_8759);
xnor U9355 (N_9355,N_8993,N_8797);
xor U9356 (N_9356,N_8317,N_8151);
xor U9357 (N_9357,N_8220,N_8163);
nor U9358 (N_9358,N_8698,N_8692);
nor U9359 (N_9359,N_8976,N_8590);
and U9360 (N_9360,N_8610,N_8266);
nand U9361 (N_9361,N_8926,N_8641);
nand U9362 (N_9362,N_8440,N_8826);
nand U9363 (N_9363,N_8187,N_8375);
and U9364 (N_9364,N_8367,N_8751);
and U9365 (N_9365,N_8841,N_8959);
and U9366 (N_9366,N_8441,N_8007);
or U9367 (N_9367,N_8544,N_8452);
nand U9368 (N_9368,N_8530,N_8642);
or U9369 (N_9369,N_8864,N_8799);
nor U9370 (N_9370,N_8138,N_8977);
xnor U9371 (N_9371,N_8586,N_8513);
and U9372 (N_9372,N_8631,N_8651);
nand U9373 (N_9373,N_8598,N_8451);
nor U9374 (N_9374,N_8401,N_8935);
nor U9375 (N_9375,N_8964,N_8774);
xnor U9376 (N_9376,N_8471,N_8194);
xnor U9377 (N_9377,N_8484,N_8244);
or U9378 (N_9378,N_8655,N_8176);
nand U9379 (N_9379,N_8449,N_8575);
xor U9380 (N_9380,N_8913,N_8547);
nor U9381 (N_9381,N_8600,N_8628);
nand U9382 (N_9382,N_8784,N_8697);
and U9383 (N_9383,N_8410,N_8426);
nand U9384 (N_9384,N_8846,N_8747);
nand U9385 (N_9385,N_8550,N_8072);
or U9386 (N_9386,N_8136,N_8986);
or U9387 (N_9387,N_8524,N_8469);
nand U9388 (N_9388,N_8475,N_8890);
and U9389 (N_9389,N_8762,N_8223);
or U9390 (N_9390,N_8885,N_8243);
nand U9391 (N_9391,N_8389,N_8687);
nor U9392 (N_9392,N_8209,N_8714);
or U9393 (N_9393,N_8172,N_8069);
xor U9394 (N_9394,N_8035,N_8490);
or U9395 (N_9395,N_8915,N_8738);
nand U9396 (N_9396,N_8334,N_8226);
nor U9397 (N_9397,N_8247,N_8483);
xor U9398 (N_9398,N_8120,N_8011);
nor U9399 (N_9399,N_8499,N_8094);
and U9400 (N_9400,N_8351,N_8739);
or U9401 (N_9401,N_8365,N_8823);
or U9402 (N_9402,N_8800,N_8191);
nor U9403 (N_9403,N_8647,N_8574);
xnor U9404 (N_9404,N_8116,N_8009);
nand U9405 (N_9405,N_8791,N_8562);
xnor U9406 (N_9406,N_8665,N_8507);
or U9407 (N_9407,N_8604,N_8447);
nor U9408 (N_9408,N_8390,N_8766);
and U9409 (N_9409,N_8142,N_8473);
nand U9410 (N_9410,N_8489,N_8965);
or U9411 (N_9411,N_8144,N_8725);
and U9412 (N_9412,N_8061,N_8708);
nand U9413 (N_9413,N_8074,N_8679);
nand U9414 (N_9414,N_8477,N_8623);
nor U9415 (N_9415,N_8543,N_8535);
nand U9416 (N_9416,N_8629,N_8040);
xnor U9417 (N_9417,N_8853,N_8113);
nand U9418 (N_9418,N_8332,N_8510);
nand U9419 (N_9419,N_8820,N_8436);
xor U9420 (N_9420,N_8724,N_8703);
xor U9421 (N_9421,N_8238,N_8188);
and U9422 (N_9422,N_8228,N_8772);
or U9423 (N_9423,N_8824,N_8103);
nor U9424 (N_9424,N_8822,N_8485);
or U9425 (N_9425,N_8609,N_8816);
and U9426 (N_9426,N_8253,N_8431);
and U9427 (N_9427,N_8622,N_8016);
nand U9428 (N_9428,N_8941,N_8052);
xnor U9429 (N_9429,N_8756,N_8255);
nor U9430 (N_9430,N_8326,N_8096);
and U9431 (N_9431,N_8031,N_8261);
or U9432 (N_9432,N_8914,N_8576);
nor U9433 (N_9433,N_8420,N_8849);
xnor U9434 (N_9434,N_8030,N_8593);
or U9435 (N_9435,N_8571,N_8201);
or U9436 (N_9436,N_8752,N_8607);
nor U9437 (N_9437,N_8021,N_8611);
nor U9438 (N_9438,N_8468,N_8289);
or U9439 (N_9439,N_8794,N_8296);
nor U9440 (N_9440,N_8533,N_8184);
or U9441 (N_9441,N_8937,N_8491);
or U9442 (N_9442,N_8707,N_8577);
nor U9443 (N_9443,N_8377,N_8356);
nand U9444 (N_9444,N_8457,N_8383);
or U9445 (N_9445,N_8865,N_8770);
or U9446 (N_9446,N_8051,N_8048);
nand U9447 (N_9447,N_8957,N_8878);
and U9448 (N_9448,N_8636,N_8156);
xnor U9449 (N_9449,N_8793,N_8973);
or U9450 (N_9450,N_8905,N_8177);
or U9451 (N_9451,N_8190,N_8509);
and U9452 (N_9452,N_8443,N_8054);
or U9453 (N_9453,N_8091,N_8340);
nand U9454 (N_9454,N_8932,N_8207);
xor U9455 (N_9455,N_8308,N_8354);
or U9456 (N_9456,N_8780,N_8059);
xnor U9457 (N_9457,N_8699,N_8869);
xor U9458 (N_9458,N_8479,N_8248);
xnor U9459 (N_9459,N_8208,N_8902);
or U9460 (N_9460,N_8183,N_8713);
or U9461 (N_9461,N_8259,N_8000);
and U9462 (N_9462,N_8455,N_8225);
and U9463 (N_9463,N_8997,N_8587);
or U9464 (N_9464,N_8486,N_8653);
nor U9465 (N_9465,N_8026,N_8382);
xor U9466 (N_9466,N_8592,N_8463);
xor U9467 (N_9467,N_8654,N_8916);
and U9468 (N_9468,N_8861,N_8358);
nand U9469 (N_9469,N_8076,N_8237);
and U9470 (N_9470,N_8202,N_8726);
nor U9471 (N_9471,N_8732,N_8947);
nor U9472 (N_9472,N_8583,N_8002);
and U9473 (N_9473,N_8938,N_8192);
or U9474 (N_9474,N_8114,N_8318);
nor U9475 (N_9475,N_8557,N_8942);
or U9476 (N_9476,N_8429,N_8922);
nand U9477 (N_9477,N_8170,N_8073);
nand U9478 (N_9478,N_8614,N_8341);
xor U9479 (N_9479,N_8735,N_8428);
nor U9480 (N_9480,N_8602,N_8556);
and U9481 (N_9481,N_8767,N_8632);
and U9482 (N_9482,N_8667,N_8022);
xnor U9483 (N_9483,N_8939,N_8414);
nor U9484 (N_9484,N_8311,N_8165);
xnor U9485 (N_9485,N_8771,N_8250);
xnor U9486 (N_9486,N_8741,N_8088);
nor U9487 (N_9487,N_8525,N_8057);
or U9488 (N_9488,N_8135,N_8511);
and U9489 (N_9489,N_8487,N_8710);
nor U9490 (N_9490,N_8538,N_8386);
nor U9491 (N_9491,N_8720,N_8335);
and U9492 (N_9492,N_8175,N_8265);
and U9493 (N_9493,N_8001,N_8789);
nor U9494 (N_9494,N_8235,N_8840);
xor U9495 (N_9495,N_8137,N_8276);
xor U9496 (N_9496,N_8229,N_8682);
xnor U9497 (N_9497,N_8346,N_8322);
nor U9498 (N_9498,N_8075,N_8213);
nand U9499 (N_9499,N_8788,N_8262);
and U9500 (N_9500,N_8581,N_8953);
nor U9501 (N_9501,N_8775,N_8362);
and U9502 (N_9502,N_8179,N_8719);
and U9503 (N_9503,N_8777,N_8880);
or U9504 (N_9504,N_8739,N_8515);
xor U9505 (N_9505,N_8734,N_8653);
and U9506 (N_9506,N_8612,N_8699);
and U9507 (N_9507,N_8358,N_8464);
nand U9508 (N_9508,N_8174,N_8707);
nand U9509 (N_9509,N_8352,N_8084);
xor U9510 (N_9510,N_8015,N_8393);
xor U9511 (N_9511,N_8122,N_8423);
nand U9512 (N_9512,N_8634,N_8193);
xor U9513 (N_9513,N_8045,N_8519);
xnor U9514 (N_9514,N_8132,N_8060);
xor U9515 (N_9515,N_8595,N_8844);
or U9516 (N_9516,N_8849,N_8918);
and U9517 (N_9517,N_8550,N_8509);
and U9518 (N_9518,N_8072,N_8885);
and U9519 (N_9519,N_8840,N_8122);
xnor U9520 (N_9520,N_8706,N_8897);
nand U9521 (N_9521,N_8001,N_8876);
xor U9522 (N_9522,N_8713,N_8053);
or U9523 (N_9523,N_8008,N_8354);
xnor U9524 (N_9524,N_8148,N_8639);
or U9525 (N_9525,N_8626,N_8129);
nand U9526 (N_9526,N_8375,N_8482);
xor U9527 (N_9527,N_8574,N_8665);
xor U9528 (N_9528,N_8600,N_8570);
nand U9529 (N_9529,N_8208,N_8176);
and U9530 (N_9530,N_8862,N_8632);
or U9531 (N_9531,N_8214,N_8288);
nand U9532 (N_9532,N_8276,N_8434);
or U9533 (N_9533,N_8757,N_8117);
nand U9534 (N_9534,N_8663,N_8876);
or U9535 (N_9535,N_8950,N_8560);
or U9536 (N_9536,N_8064,N_8814);
xor U9537 (N_9537,N_8612,N_8764);
or U9538 (N_9538,N_8501,N_8273);
or U9539 (N_9539,N_8895,N_8537);
or U9540 (N_9540,N_8962,N_8170);
nand U9541 (N_9541,N_8068,N_8915);
xor U9542 (N_9542,N_8010,N_8265);
nor U9543 (N_9543,N_8324,N_8383);
nand U9544 (N_9544,N_8175,N_8617);
and U9545 (N_9545,N_8361,N_8446);
nand U9546 (N_9546,N_8831,N_8879);
xor U9547 (N_9547,N_8827,N_8982);
or U9548 (N_9548,N_8155,N_8843);
xor U9549 (N_9549,N_8963,N_8176);
nor U9550 (N_9550,N_8363,N_8100);
and U9551 (N_9551,N_8135,N_8246);
nor U9552 (N_9552,N_8011,N_8731);
and U9553 (N_9553,N_8792,N_8527);
nand U9554 (N_9554,N_8566,N_8109);
nor U9555 (N_9555,N_8442,N_8181);
and U9556 (N_9556,N_8518,N_8184);
xnor U9557 (N_9557,N_8806,N_8083);
nor U9558 (N_9558,N_8340,N_8806);
nor U9559 (N_9559,N_8453,N_8149);
xnor U9560 (N_9560,N_8730,N_8256);
nand U9561 (N_9561,N_8017,N_8364);
nand U9562 (N_9562,N_8545,N_8123);
nor U9563 (N_9563,N_8194,N_8223);
nor U9564 (N_9564,N_8122,N_8922);
xnor U9565 (N_9565,N_8795,N_8495);
nor U9566 (N_9566,N_8045,N_8811);
xor U9567 (N_9567,N_8522,N_8706);
or U9568 (N_9568,N_8056,N_8659);
nand U9569 (N_9569,N_8264,N_8824);
nor U9570 (N_9570,N_8625,N_8928);
and U9571 (N_9571,N_8224,N_8116);
or U9572 (N_9572,N_8528,N_8417);
nand U9573 (N_9573,N_8485,N_8083);
nor U9574 (N_9574,N_8498,N_8840);
nor U9575 (N_9575,N_8060,N_8932);
or U9576 (N_9576,N_8033,N_8784);
nor U9577 (N_9577,N_8521,N_8281);
nor U9578 (N_9578,N_8466,N_8470);
xor U9579 (N_9579,N_8258,N_8352);
nor U9580 (N_9580,N_8897,N_8484);
and U9581 (N_9581,N_8802,N_8520);
xnor U9582 (N_9582,N_8457,N_8346);
or U9583 (N_9583,N_8536,N_8921);
nand U9584 (N_9584,N_8566,N_8338);
nand U9585 (N_9585,N_8159,N_8804);
xor U9586 (N_9586,N_8972,N_8945);
and U9587 (N_9587,N_8846,N_8254);
and U9588 (N_9588,N_8848,N_8139);
nor U9589 (N_9589,N_8996,N_8409);
nor U9590 (N_9590,N_8306,N_8835);
and U9591 (N_9591,N_8809,N_8414);
nor U9592 (N_9592,N_8176,N_8429);
nor U9593 (N_9593,N_8442,N_8870);
and U9594 (N_9594,N_8563,N_8421);
nand U9595 (N_9595,N_8736,N_8207);
nor U9596 (N_9596,N_8624,N_8546);
nand U9597 (N_9597,N_8436,N_8870);
xnor U9598 (N_9598,N_8287,N_8311);
xnor U9599 (N_9599,N_8022,N_8134);
nor U9600 (N_9600,N_8215,N_8257);
nor U9601 (N_9601,N_8958,N_8892);
xor U9602 (N_9602,N_8276,N_8649);
nand U9603 (N_9603,N_8090,N_8175);
or U9604 (N_9604,N_8250,N_8539);
or U9605 (N_9605,N_8247,N_8979);
nand U9606 (N_9606,N_8119,N_8632);
nand U9607 (N_9607,N_8405,N_8887);
and U9608 (N_9608,N_8228,N_8771);
nand U9609 (N_9609,N_8569,N_8183);
and U9610 (N_9610,N_8060,N_8728);
or U9611 (N_9611,N_8541,N_8968);
nand U9612 (N_9612,N_8789,N_8790);
xor U9613 (N_9613,N_8580,N_8013);
or U9614 (N_9614,N_8884,N_8794);
xor U9615 (N_9615,N_8975,N_8320);
xor U9616 (N_9616,N_8439,N_8844);
nand U9617 (N_9617,N_8333,N_8442);
nand U9618 (N_9618,N_8024,N_8967);
xor U9619 (N_9619,N_8484,N_8707);
and U9620 (N_9620,N_8912,N_8954);
nand U9621 (N_9621,N_8540,N_8345);
nand U9622 (N_9622,N_8198,N_8523);
nor U9623 (N_9623,N_8577,N_8696);
or U9624 (N_9624,N_8469,N_8048);
and U9625 (N_9625,N_8724,N_8013);
or U9626 (N_9626,N_8576,N_8615);
nand U9627 (N_9627,N_8253,N_8938);
xor U9628 (N_9628,N_8250,N_8367);
and U9629 (N_9629,N_8366,N_8647);
nand U9630 (N_9630,N_8706,N_8611);
nor U9631 (N_9631,N_8571,N_8194);
nand U9632 (N_9632,N_8577,N_8119);
or U9633 (N_9633,N_8889,N_8279);
or U9634 (N_9634,N_8581,N_8182);
nand U9635 (N_9635,N_8965,N_8132);
nand U9636 (N_9636,N_8822,N_8617);
nand U9637 (N_9637,N_8234,N_8933);
or U9638 (N_9638,N_8739,N_8147);
or U9639 (N_9639,N_8437,N_8689);
nand U9640 (N_9640,N_8903,N_8598);
nand U9641 (N_9641,N_8189,N_8206);
nor U9642 (N_9642,N_8484,N_8183);
nor U9643 (N_9643,N_8318,N_8501);
and U9644 (N_9644,N_8649,N_8588);
xnor U9645 (N_9645,N_8518,N_8581);
nor U9646 (N_9646,N_8562,N_8232);
xnor U9647 (N_9647,N_8873,N_8751);
and U9648 (N_9648,N_8254,N_8525);
nor U9649 (N_9649,N_8299,N_8868);
nand U9650 (N_9650,N_8026,N_8573);
xnor U9651 (N_9651,N_8644,N_8476);
nor U9652 (N_9652,N_8614,N_8456);
or U9653 (N_9653,N_8621,N_8402);
nor U9654 (N_9654,N_8366,N_8733);
or U9655 (N_9655,N_8104,N_8474);
nand U9656 (N_9656,N_8688,N_8512);
nor U9657 (N_9657,N_8705,N_8890);
or U9658 (N_9658,N_8734,N_8004);
nor U9659 (N_9659,N_8552,N_8263);
xor U9660 (N_9660,N_8423,N_8602);
xor U9661 (N_9661,N_8017,N_8056);
xor U9662 (N_9662,N_8941,N_8862);
and U9663 (N_9663,N_8194,N_8967);
nand U9664 (N_9664,N_8336,N_8373);
xnor U9665 (N_9665,N_8913,N_8516);
nand U9666 (N_9666,N_8181,N_8015);
and U9667 (N_9667,N_8369,N_8017);
nand U9668 (N_9668,N_8076,N_8183);
or U9669 (N_9669,N_8387,N_8114);
nand U9670 (N_9670,N_8898,N_8850);
xor U9671 (N_9671,N_8652,N_8791);
or U9672 (N_9672,N_8222,N_8702);
or U9673 (N_9673,N_8026,N_8714);
and U9674 (N_9674,N_8955,N_8597);
and U9675 (N_9675,N_8523,N_8904);
or U9676 (N_9676,N_8462,N_8649);
xnor U9677 (N_9677,N_8171,N_8143);
nor U9678 (N_9678,N_8837,N_8040);
nor U9679 (N_9679,N_8371,N_8055);
nor U9680 (N_9680,N_8676,N_8266);
nor U9681 (N_9681,N_8610,N_8776);
or U9682 (N_9682,N_8051,N_8589);
nor U9683 (N_9683,N_8677,N_8807);
and U9684 (N_9684,N_8333,N_8629);
or U9685 (N_9685,N_8345,N_8172);
xor U9686 (N_9686,N_8745,N_8651);
nand U9687 (N_9687,N_8416,N_8312);
and U9688 (N_9688,N_8868,N_8333);
or U9689 (N_9689,N_8322,N_8587);
nand U9690 (N_9690,N_8196,N_8787);
and U9691 (N_9691,N_8161,N_8910);
nand U9692 (N_9692,N_8255,N_8375);
nand U9693 (N_9693,N_8402,N_8349);
and U9694 (N_9694,N_8481,N_8963);
or U9695 (N_9695,N_8614,N_8272);
nor U9696 (N_9696,N_8702,N_8703);
and U9697 (N_9697,N_8539,N_8716);
nand U9698 (N_9698,N_8656,N_8653);
or U9699 (N_9699,N_8716,N_8005);
nand U9700 (N_9700,N_8616,N_8574);
xnor U9701 (N_9701,N_8951,N_8264);
and U9702 (N_9702,N_8138,N_8525);
nand U9703 (N_9703,N_8821,N_8007);
xnor U9704 (N_9704,N_8298,N_8652);
nand U9705 (N_9705,N_8316,N_8927);
nor U9706 (N_9706,N_8006,N_8712);
xnor U9707 (N_9707,N_8394,N_8840);
nor U9708 (N_9708,N_8534,N_8970);
and U9709 (N_9709,N_8588,N_8263);
xnor U9710 (N_9710,N_8378,N_8810);
nor U9711 (N_9711,N_8779,N_8088);
nand U9712 (N_9712,N_8495,N_8003);
and U9713 (N_9713,N_8262,N_8777);
and U9714 (N_9714,N_8494,N_8100);
nor U9715 (N_9715,N_8206,N_8806);
and U9716 (N_9716,N_8023,N_8898);
nor U9717 (N_9717,N_8503,N_8274);
and U9718 (N_9718,N_8145,N_8043);
xnor U9719 (N_9719,N_8276,N_8328);
nand U9720 (N_9720,N_8030,N_8542);
nand U9721 (N_9721,N_8780,N_8185);
xnor U9722 (N_9722,N_8068,N_8840);
nand U9723 (N_9723,N_8771,N_8565);
or U9724 (N_9724,N_8606,N_8743);
nand U9725 (N_9725,N_8002,N_8706);
nor U9726 (N_9726,N_8805,N_8176);
or U9727 (N_9727,N_8655,N_8856);
and U9728 (N_9728,N_8185,N_8207);
xor U9729 (N_9729,N_8183,N_8617);
xor U9730 (N_9730,N_8986,N_8369);
nor U9731 (N_9731,N_8955,N_8171);
nor U9732 (N_9732,N_8979,N_8789);
nor U9733 (N_9733,N_8711,N_8644);
nand U9734 (N_9734,N_8940,N_8711);
and U9735 (N_9735,N_8922,N_8110);
and U9736 (N_9736,N_8450,N_8792);
or U9737 (N_9737,N_8570,N_8233);
nand U9738 (N_9738,N_8628,N_8410);
nand U9739 (N_9739,N_8854,N_8102);
xor U9740 (N_9740,N_8609,N_8464);
or U9741 (N_9741,N_8892,N_8019);
and U9742 (N_9742,N_8315,N_8903);
xor U9743 (N_9743,N_8530,N_8348);
or U9744 (N_9744,N_8325,N_8878);
or U9745 (N_9745,N_8908,N_8270);
nand U9746 (N_9746,N_8808,N_8103);
and U9747 (N_9747,N_8897,N_8188);
nor U9748 (N_9748,N_8175,N_8212);
nand U9749 (N_9749,N_8417,N_8145);
or U9750 (N_9750,N_8981,N_8333);
and U9751 (N_9751,N_8091,N_8005);
xnor U9752 (N_9752,N_8034,N_8499);
nand U9753 (N_9753,N_8719,N_8467);
xnor U9754 (N_9754,N_8622,N_8397);
nand U9755 (N_9755,N_8774,N_8386);
nor U9756 (N_9756,N_8108,N_8712);
nor U9757 (N_9757,N_8096,N_8909);
xor U9758 (N_9758,N_8619,N_8637);
and U9759 (N_9759,N_8431,N_8584);
and U9760 (N_9760,N_8161,N_8344);
nand U9761 (N_9761,N_8100,N_8956);
or U9762 (N_9762,N_8230,N_8030);
or U9763 (N_9763,N_8359,N_8123);
xor U9764 (N_9764,N_8875,N_8951);
nand U9765 (N_9765,N_8938,N_8662);
nand U9766 (N_9766,N_8309,N_8300);
nand U9767 (N_9767,N_8655,N_8604);
nor U9768 (N_9768,N_8692,N_8522);
and U9769 (N_9769,N_8398,N_8755);
and U9770 (N_9770,N_8097,N_8423);
nand U9771 (N_9771,N_8031,N_8174);
nand U9772 (N_9772,N_8942,N_8865);
and U9773 (N_9773,N_8273,N_8756);
xor U9774 (N_9774,N_8527,N_8755);
xor U9775 (N_9775,N_8174,N_8408);
nand U9776 (N_9776,N_8625,N_8593);
nand U9777 (N_9777,N_8878,N_8079);
nor U9778 (N_9778,N_8290,N_8263);
nand U9779 (N_9779,N_8013,N_8608);
nand U9780 (N_9780,N_8635,N_8662);
and U9781 (N_9781,N_8059,N_8481);
or U9782 (N_9782,N_8014,N_8102);
xnor U9783 (N_9783,N_8146,N_8565);
nand U9784 (N_9784,N_8321,N_8874);
xor U9785 (N_9785,N_8108,N_8142);
nor U9786 (N_9786,N_8162,N_8846);
nor U9787 (N_9787,N_8983,N_8663);
and U9788 (N_9788,N_8353,N_8233);
nor U9789 (N_9789,N_8559,N_8843);
or U9790 (N_9790,N_8579,N_8176);
nand U9791 (N_9791,N_8329,N_8221);
nor U9792 (N_9792,N_8850,N_8577);
and U9793 (N_9793,N_8123,N_8588);
and U9794 (N_9794,N_8073,N_8489);
nand U9795 (N_9795,N_8872,N_8858);
or U9796 (N_9796,N_8219,N_8349);
and U9797 (N_9797,N_8631,N_8605);
xnor U9798 (N_9798,N_8981,N_8279);
xor U9799 (N_9799,N_8439,N_8478);
xnor U9800 (N_9800,N_8566,N_8339);
or U9801 (N_9801,N_8626,N_8633);
nand U9802 (N_9802,N_8161,N_8318);
nand U9803 (N_9803,N_8286,N_8326);
nor U9804 (N_9804,N_8549,N_8889);
nand U9805 (N_9805,N_8578,N_8493);
nand U9806 (N_9806,N_8043,N_8611);
or U9807 (N_9807,N_8965,N_8506);
nor U9808 (N_9808,N_8464,N_8996);
nor U9809 (N_9809,N_8173,N_8418);
xnor U9810 (N_9810,N_8851,N_8466);
xor U9811 (N_9811,N_8887,N_8506);
nor U9812 (N_9812,N_8269,N_8717);
xor U9813 (N_9813,N_8851,N_8252);
nor U9814 (N_9814,N_8602,N_8499);
xor U9815 (N_9815,N_8264,N_8106);
nand U9816 (N_9816,N_8603,N_8964);
and U9817 (N_9817,N_8430,N_8048);
nand U9818 (N_9818,N_8412,N_8386);
or U9819 (N_9819,N_8854,N_8669);
nand U9820 (N_9820,N_8550,N_8796);
nand U9821 (N_9821,N_8656,N_8021);
or U9822 (N_9822,N_8833,N_8143);
nand U9823 (N_9823,N_8858,N_8491);
xor U9824 (N_9824,N_8679,N_8099);
nand U9825 (N_9825,N_8211,N_8311);
or U9826 (N_9826,N_8464,N_8199);
nor U9827 (N_9827,N_8166,N_8679);
nor U9828 (N_9828,N_8562,N_8037);
nor U9829 (N_9829,N_8477,N_8034);
nor U9830 (N_9830,N_8776,N_8313);
or U9831 (N_9831,N_8182,N_8031);
nor U9832 (N_9832,N_8293,N_8010);
nor U9833 (N_9833,N_8180,N_8158);
xor U9834 (N_9834,N_8852,N_8236);
xnor U9835 (N_9835,N_8373,N_8203);
or U9836 (N_9836,N_8715,N_8181);
or U9837 (N_9837,N_8098,N_8018);
nor U9838 (N_9838,N_8205,N_8295);
xor U9839 (N_9839,N_8018,N_8955);
xor U9840 (N_9840,N_8825,N_8731);
nand U9841 (N_9841,N_8436,N_8511);
nor U9842 (N_9842,N_8440,N_8284);
nor U9843 (N_9843,N_8496,N_8297);
and U9844 (N_9844,N_8490,N_8781);
nand U9845 (N_9845,N_8673,N_8395);
or U9846 (N_9846,N_8912,N_8194);
and U9847 (N_9847,N_8065,N_8821);
or U9848 (N_9848,N_8234,N_8594);
or U9849 (N_9849,N_8394,N_8967);
nand U9850 (N_9850,N_8551,N_8012);
or U9851 (N_9851,N_8029,N_8149);
nand U9852 (N_9852,N_8478,N_8753);
xor U9853 (N_9853,N_8745,N_8719);
or U9854 (N_9854,N_8843,N_8005);
nand U9855 (N_9855,N_8564,N_8924);
and U9856 (N_9856,N_8522,N_8556);
and U9857 (N_9857,N_8967,N_8917);
and U9858 (N_9858,N_8846,N_8213);
xnor U9859 (N_9859,N_8496,N_8238);
and U9860 (N_9860,N_8083,N_8080);
or U9861 (N_9861,N_8846,N_8119);
and U9862 (N_9862,N_8390,N_8109);
and U9863 (N_9863,N_8239,N_8621);
nand U9864 (N_9864,N_8846,N_8644);
nor U9865 (N_9865,N_8783,N_8791);
or U9866 (N_9866,N_8074,N_8508);
or U9867 (N_9867,N_8810,N_8201);
nand U9868 (N_9868,N_8888,N_8277);
and U9869 (N_9869,N_8004,N_8991);
nand U9870 (N_9870,N_8819,N_8468);
nor U9871 (N_9871,N_8136,N_8210);
nand U9872 (N_9872,N_8746,N_8311);
or U9873 (N_9873,N_8546,N_8631);
nand U9874 (N_9874,N_8578,N_8844);
nand U9875 (N_9875,N_8110,N_8855);
nor U9876 (N_9876,N_8698,N_8706);
and U9877 (N_9877,N_8959,N_8426);
or U9878 (N_9878,N_8461,N_8922);
and U9879 (N_9879,N_8734,N_8477);
xnor U9880 (N_9880,N_8506,N_8571);
nor U9881 (N_9881,N_8623,N_8578);
nand U9882 (N_9882,N_8255,N_8240);
or U9883 (N_9883,N_8192,N_8977);
nand U9884 (N_9884,N_8482,N_8543);
or U9885 (N_9885,N_8723,N_8204);
nor U9886 (N_9886,N_8841,N_8849);
and U9887 (N_9887,N_8569,N_8674);
nand U9888 (N_9888,N_8699,N_8299);
and U9889 (N_9889,N_8907,N_8608);
or U9890 (N_9890,N_8347,N_8133);
nand U9891 (N_9891,N_8113,N_8281);
or U9892 (N_9892,N_8952,N_8800);
and U9893 (N_9893,N_8753,N_8895);
and U9894 (N_9894,N_8472,N_8917);
nand U9895 (N_9895,N_8913,N_8543);
nor U9896 (N_9896,N_8657,N_8808);
or U9897 (N_9897,N_8299,N_8114);
nand U9898 (N_9898,N_8919,N_8311);
or U9899 (N_9899,N_8534,N_8659);
and U9900 (N_9900,N_8525,N_8571);
and U9901 (N_9901,N_8378,N_8256);
nand U9902 (N_9902,N_8520,N_8994);
and U9903 (N_9903,N_8068,N_8675);
or U9904 (N_9904,N_8526,N_8666);
nor U9905 (N_9905,N_8043,N_8301);
xnor U9906 (N_9906,N_8796,N_8931);
nor U9907 (N_9907,N_8446,N_8012);
nand U9908 (N_9908,N_8941,N_8714);
and U9909 (N_9909,N_8702,N_8776);
and U9910 (N_9910,N_8197,N_8449);
nor U9911 (N_9911,N_8002,N_8280);
nand U9912 (N_9912,N_8627,N_8617);
or U9913 (N_9913,N_8605,N_8030);
xor U9914 (N_9914,N_8072,N_8147);
nor U9915 (N_9915,N_8384,N_8269);
xor U9916 (N_9916,N_8895,N_8072);
nor U9917 (N_9917,N_8023,N_8144);
or U9918 (N_9918,N_8940,N_8158);
nor U9919 (N_9919,N_8610,N_8631);
and U9920 (N_9920,N_8641,N_8541);
nand U9921 (N_9921,N_8972,N_8045);
or U9922 (N_9922,N_8756,N_8248);
nor U9923 (N_9923,N_8571,N_8048);
xor U9924 (N_9924,N_8081,N_8781);
nor U9925 (N_9925,N_8994,N_8210);
or U9926 (N_9926,N_8219,N_8755);
and U9927 (N_9927,N_8981,N_8590);
and U9928 (N_9928,N_8174,N_8091);
and U9929 (N_9929,N_8843,N_8319);
nor U9930 (N_9930,N_8449,N_8259);
and U9931 (N_9931,N_8049,N_8005);
xor U9932 (N_9932,N_8614,N_8962);
or U9933 (N_9933,N_8842,N_8941);
nor U9934 (N_9934,N_8976,N_8352);
nor U9935 (N_9935,N_8721,N_8048);
nand U9936 (N_9936,N_8834,N_8824);
nor U9937 (N_9937,N_8140,N_8167);
or U9938 (N_9938,N_8507,N_8985);
or U9939 (N_9939,N_8165,N_8058);
nor U9940 (N_9940,N_8263,N_8069);
nand U9941 (N_9941,N_8654,N_8992);
and U9942 (N_9942,N_8928,N_8977);
and U9943 (N_9943,N_8347,N_8768);
nand U9944 (N_9944,N_8472,N_8895);
and U9945 (N_9945,N_8278,N_8404);
and U9946 (N_9946,N_8044,N_8235);
nand U9947 (N_9947,N_8285,N_8846);
xor U9948 (N_9948,N_8672,N_8772);
nor U9949 (N_9949,N_8367,N_8338);
or U9950 (N_9950,N_8741,N_8654);
nor U9951 (N_9951,N_8216,N_8201);
or U9952 (N_9952,N_8867,N_8193);
xnor U9953 (N_9953,N_8255,N_8557);
xor U9954 (N_9954,N_8600,N_8684);
and U9955 (N_9955,N_8756,N_8978);
or U9956 (N_9956,N_8656,N_8848);
and U9957 (N_9957,N_8813,N_8678);
nor U9958 (N_9958,N_8280,N_8860);
nand U9959 (N_9959,N_8171,N_8933);
or U9960 (N_9960,N_8579,N_8838);
or U9961 (N_9961,N_8875,N_8466);
nand U9962 (N_9962,N_8749,N_8249);
nand U9963 (N_9963,N_8644,N_8936);
xor U9964 (N_9964,N_8876,N_8720);
or U9965 (N_9965,N_8347,N_8482);
nand U9966 (N_9966,N_8687,N_8641);
xor U9967 (N_9967,N_8951,N_8451);
or U9968 (N_9968,N_8751,N_8283);
or U9969 (N_9969,N_8875,N_8241);
xnor U9970 (N_9970,N_8419,N_8117);
and U9971 (N_9971,N_8593,N_8014);
nor U9972 (N_9972,N_8793,N_8547);
nor U9973 (N_9973,N_8944,N_8323);
or U9974 (N_9974,N_8763,N_8700);
xor U9975 (N_9975,N_8284,N_8326);
xor U9976 (N_9976,N_8747,N_8635);
xnor U9977 (N_9977,N_8100,N_8271);
nor U9978 (N_9978,N_8975,N_8626);
xor U9979 (N_9979,N_8472,N_8307);
xor U9980 (N_9980,N_8777,N_8312);
xor U9981 (N_9981,N_8510,N_8272);
nor U9982 (N_9982,N_8568,N_8227);
or U9983 (N_9983,N_8069,N_8928);
or U9984 (N_9984,N_8570,N_8176);
and U9985 (N_9985,N_8812,N_8022);
nand U9986 (N_9986,N_8189,N_8257);
xnor U9987 (N_9987,N_8508,N_8571);
or U9988 (N_9988,N_8287,N_8181);
nor U9989 (N_9989,N_8755,N_8031);
nor U9990 (N_9990,N_8793,N_8159);
nor U9991 (N_9991,N_8465,N_8188);
xnor U9992 (N_9992,N_8860,N_8455);
and U9993 (N_9993,N_8446,N_8331);
xnor U9994 (N_9994,N_8018,N_8240);
or U9995 (N_9995,N_8854,N_8653);
or U9996 (N_9996,N_8137,N_8828);
or U9997 (N_9997,N_8062,N_8693);
nor U9998 (N_9998,N_8938,N_8183);
nand U9999 (N_9999,N_8079,N_8818);
and U10000 (N_10000,N_9044,N_9035);
or U10001 (N_10001,N_9352,N_9291);
nand U10002 (N_10002,N_9506,N_9161);
nand U10003 (N_10003,N_9400,N_9608);
nor U10004 (N_10004,N_9524,N_9290);
nand U10005 (N_10005,N_9888,N_9060);
nor U10006 (N_10006,N_9926,N_9149);
and U10007 (N_10007,N_9979,N_9756);
nor U10008 (N_10008,N_9542,N_9385);
or U10009 (N_10009,N_9374,N_9207);
and U10010 (N_10010,N_9558,N_9763);
and U10011 (N_10011,N_9118,N_9719);
xnor U10012 (N_10012,N_9484,N_9805);
or U10013 (N_10013,N_9139,N_9544);
nand U10014 (N_10014,N_9194,N_9783);
nor U10015 (N_10015,N_9659,N_9618);
xnor U10016 (N_10016,N_9178,N_9096);
xnor U10017 (N_10017,N_9319,N_9577);
and U10018 (N_10018,N_9933,N_9058);
and U10019 (N_10019,N_9799,N_9968);
nor U10020 (N_10020,N_9476,N_9419);
nor U10021 (N_10021,N_9731,N_9960);
and U10022 (N_10022,N_9499,N_9620);
nor U10023 (N_10023,N_9737,N_9257);
or U10024 (N_10024,N_9985,N_9367);
nor U10025 (N_10025,N_9582,N_9706);
nand U10026 (N_10026,N_9029,N_9231);
nor U10027 (N_10027,N_9376,N_9741);
nor U10028 (N_10028,N_9022,N_9898);
xnor U10029 (N_10029,N_9510,N_9301);
and U10030 (N_10030,N_9818,N_9609);
and U10031 (N_10031,N_9346,N_9769);
nand U10032 (N_10032,N_9403,N_9165);
or U10033 (N_10033,N_9736,N_9974);
and U10034 (N_10034,N_9028,N_9622);
and U10035 (N_10035,N_9759,N_9148);
xor U10036 (N_10036,N_9122,N_9417);
nor U10037 (N_10037,N_9869,N_9481);
nor U10038 (N_10038,N_9503,N_9964);
nand U10039 (N_10039,N_9535,N_9611);
and U10040 (N_10040,N_9652,N_9594);
nand U10041 (N_10041,N_9619,N_9184);
nor U10042 (N_10042,N_9021,N_9976);
or U10043 (N_10043,N_9552,N_9851);
nor U10044 (N_10044,N_9893,N_9754);
xor U10045 (N_10045,N_9463,N_9802);
xor U10046 (N_10046,N_9935,N_9088);
and U10047 (N_10047,N_9091,N_9863);
xnor U10048 (N_10048,N_9639,N_9950);
nand U10049 (N_10049,N_9697,N_9886);
nand U10050 (N_10050,N_9437,N_9342);
nand U10051 (N_10051,N_9186,N_9293);
xor U10052 (N_10052,N_9331,N_9540);
and U10053 (N_10053,N_9525,N_9292);
xnor U10054 (N_10054,N_9930,N_9114);
or U10055 (N_10055,N_9171,N_9948);
or U10056 (N_10056,N_9313,N_9341);
xor U10057 (N_10057,N_9444,N_9682);
nor U10058 (N_10058,N_9547,N_9738);
nand U10059 (N_10059,N_9823,N_9792);
nor U10060 (N_10060,N_9046,N_9045);
nor U10061 (N_10061,N_9730,N_9065);
or U10062 (N_10062,N_9461,N_9879);
or U10063 (N_10063,N_9143,N_9026);
nor U10064 (N_10064,N_9664,N_9732);
nand U10065 (N_10065,N_9214,N_9631);
nand U10066 (N_10066,N_9339,N_9438);
nor U10067 (N_10067,N_9151,N_9453);
nand U10068 (N_10068,N_9702,N_9614);
nor U10069 (N_10069,N_9877,N_9066);
nand U10070 (N_10070,N_9193,N_9435);
xnor U10071 (N_10071,N_9366,N_9222);
nand U10072 (N_10072,N_9883,N_9982);
nor U10073 (N_10073,N_9031,N_9857);
nand U10074 (N_10074,N_9358,N_9523);
xor U10075 (N_10075,N_9955,N_9472);
or U10076 (N_10076,N_9800,N_9746);
xnor U10077 (N_10077,N_9971,N_9003);
xor U10078 (N_10078,N_9957,N_9519);
or U10079 (N_10079,N_9309,N_9545);
and U10080 (N_10080,N_9905,N_9534);
or U10081 (N_10081,N_9873,N_9345);
nand U10082 (N_10082,N_9602,N_9870);
or U10083 (N_10083,N_9267,N_9915);
xnor U10084 (N_10084,N_9777,N_9686);
nand U10085 (N_10085,N_9679,N_9411);
nor U10086 (N_10086,N_9943,N_9755);
or U10087 (N_10087,N_9793,N_9043);
or U10088 (N_10088,N_9491,N_9150);
or U10089 (N_10089,N_9703,N_9928);
xnor U10090 (N_10090,N_9610,N_9642);
nor U10091 (N_10091,N_9827,N_9215);
nor U10092 (N_10092,N_9418,N_9287);
and U10093 (N_10093,N_9593,N_9439);
nor U10094 (N_10094,N_9784,N_9571);
nand U10095 (N_10095,N_9729,N_9424);
nor U10096 (N_10096,N_9647,N_9271);
and U10097 (N_10097,N_9744,N_9742);
or U10098 (N_10098,N_9906,N_9182);
nor U10099 (N_10099,N_9504,N_9489);
and U10100 (N_10100,N_9468,N_9349);
nor U10101 (N_10101,N_9655,N_9170);
or U10102 (N_10102,N_9913,N_9087);
and U10103 (N_10103,N_9621,N_9520);
nor U10104 (N_10104,N_9543,N_9392);
nand U10105 (N_10105,N_9138,N_9634);
and U10106 (N_10106,N_9762,N_9590);
or U10107 (N_10107,N_9006,N_9064);
nor U10108 (N_10108,N_9104,N_9350);
and U10109 (N_10109,N_9377,N_9255);
nor U10110 (N_10110,N_9119,N_9597);
and U10111 (N_10111,N_9187,N_9954);
nand U10112 (N_10112,N_9401,N_9852);
and U10113 (N_10113,N_9426,N_9651);
and U10114 (N_10114,N_9123,N_9166);
or U10115 (N_10115,N_9821,N_9557);
or U10116 (N_10116,N_9268,N_9383);
xnor U10117 (N_10117,N_9183,N_9497);
or U10118 (N_10118,N_9208,N_9764);
or U10119 (N_10119,N_9717,N_9202);
and U10120 (N_10120,N_9250,N_9917);
and U10121 (N_10121,N_9430,N_9623);
nand U10122 (N_10122,N_9889,N_9724);
xor U10123 (N_10123,N_9692,N_9097);
nand U10124 (N_10124,N_9939,N_9600);
or U10125 (N_10125,N_9455,N_9284);
xor U10126 (N_10126,N_9993,N_9113);
and U10127 (N_10127,N_9226,N_9042);
xnor U10128 (N_10128,N_9727,N_9080);
nand U10129 (N_10129,N_9130,N_9953);
and U10130 (N_10130,N_9705,N_9887);
xor U10131 (N_10131,N_9258,N_9630);
and U10132 (N_10132,N_9711,N_9036);
xor U10133 (N_10133,N_9074,N_9279);
nor U10134 (N_10134,N_9308,N_9371);
xnor U10135 (N_10135,N_9106,N_9340);
xnor U10136 (N_10136,N_9030,N_9062);
nand U10137 (N_10137,N_9740,N_9266);
and U10138 (N_10138,N_9512,N_9635);
nor U10139 (N_10139,N_9452,N_9919);
and U10140 (N_10140,N_9568,N_9613);
xnor U10141 (N_10141,N_9563,N_9837);
nand U10142 (N_10142,N_9422,N_9154);
nor U10143 (N_10143,N_9068,N_9945);
or U10144 (N_10144,N_9361,N_9517);
nand U10145 (N_10145,N_9907,N_9144);
or U10146 (N_10146,N_9265,N_9332);
or U10147 (N_10147,N_9561,N_9606);
and U10148 (N_10148,N_9910,N_9522);
or U10149 (N_10149,N_9567,N_9248);
or U10150 (N_10150,N_9728,N_9270);
nor U10151 (N_10151,N_9989,N_9205);
xnor U10152 (N_10152,N_9809,N_9120);
xnor U10153 (N_10153,N_9644,N_9766);
or U10154 (N_10154,N_9177,N_9082);
nand U10155 (N_10155,N_9500,N_9688);
and U10156 (N_10156,N_9986,N_9896);
or U10157 (N_10157,N_9861,N_9531);
nor U10158 (N_10158,N_9903,N_9019);
nand U10159 (N_10159,N_9718,N_9211);
xnor U10160 (N_10160,N_9908,N_9856);
or U10161 (N_10161,N_9244,N_9956);
or U10162 (N_10162,N_9918,N_9372);
nor U10163 (N_10163,N_9078,N_9431);
xor U10164 (N_10164,N_9174,N_9236);
and U10165 (N_10165,N_9607,N_9768);
xor U10166 (N_10166,N_9318,N_9053);
nand U10167 (N_10167,N_9946,N_9115);
and U10168 (N_10168,N_9774,N_9427);
xor U10169 (N_10169,N_9232,N_9395);
or U10170 (N_10170,N_9428,N_9480);
nor U10171 (N_10171,N_9810,N_9798);
nand U10172 (N_10172,N_9402,N_9460);
nand U10173 (N_10173,N_9627,N_9537);
xnor U10174 (N_10174,N_9983,N_9160);
xnor U10175 (N_10175,N_9456,N_9882);
nor U10176 (N_10176,N_9009,N_9116);
nor U10177 (N_10177,N_9677,N_9575);
or U10178 (N_10178,N_9826,N_9146);
and U10179 (N_10179,N_9787,N_9722);
nand U10180 (N_10180,N_9312,N_9824);
or U10181 (N_10181,N_9599,N_9192);
or U10182 (N_10182,N_9649,N_9854);
nand U10183 (N_10183,N_9325,N_9197);
xnor U10184 (N_10184,N_9147,N_9018);
nand U10185 (N_10185,N_9834,N_9498);
and U10186 (N_10186,N_9334,N_9942);
nor U10187 (N_10187,N_9434,N_9382);
or U10188 (N_10188,N_9526,N_9344);
nand U10189 (N_10189,N_9663,N_9761);
nor U10190 (N_10190,N_9176,N_9351);
nor U10191 (N_10191,N_9335,N_9962);
nor U10192 (N_10192,N_9758,N_9085);
or U10193 (N_10193,N_9583,N_9548);
and U10194 (N_10194,N_9155,N_9038);
xor U10195 (N_10195,N_9254,N_9289);
nand U10196 (N_10196,N_9820,N_9733);
or U10197 (N_10197,N_9714,N_9923);
and U10198 (N_10198,N_9041,N_9675);
or U10199 (N_10199,N_9264,N_9572);
and U10200 (N_10200,N_9513,N_9328);
or U10201 (N_10201,N_9716,N_9363);
nor U10202 (N_10202,N_9134,N_9140);
nor U10203 (N_10203,N_9734,N_9128);
or U10204 (N_10204,N_9885,N_9788);
and U10205 (N_10205,N_9218,N_9391);
or U10206 (N_10206,N_9704,N_9855);
or U10207 (N_10207,N_9396,N_9812);
or U10208 (N_10208,N_9375,N_9816);
nand U10209 (N_10209,N_9099,N_9315);
xnor U10210 (N_10210,N_9587,N_9813);
nand U10211 (N_10211,N_9860,N_9646);
nand U10212 (N_10212,N_9121,N_9189);
or U10213 (N_10213,N_9574,N_9598);
nand U10214 (N_10214,N_9604,N_9937);
nor U10215 (N_10215,N_9234,N_9486);
nor U10216 (N_10216,N_9168,N_9237);
nor U10217 (N_10217,N_9735,N_9507);
nand U10218 (N_10218,N_9063,N_9242);
nand U10219 (N_10219,N_9451,N_9014);
nor U10220 (N_10220,N_9090,N_9839);
or U10221 (N_10221,N_9348,N_9829);
nand U10222 (N_10222,N_9201,N_9836);
and U10223 (N_10223,N_9680,N_9076);
xor U10224 (N_10224,N_9164,N_9551);
and U10225 (N_10225,N_9589,N_9696);
xor U10226 (N_10226,N_9892,N_9111);
or U10227 (N_10227,N_9089,N_9102);
nor U10228 (N_10228,N_9317,N_9083);
nand U10229 (N_10229,N_9853,N_9238);
nand U10230 (N_10230,N_9409,N_9676);
nor U10231 (N_10231,N_9566,N_9387);
and U10232 (N_10232,N_9353,N_9162);
nor U10233 (N_10233,N_9715,N_9681);
xnor U10234 (N_10234,N_9327,N_9198);
and U10235 (N_10235,N_9748,N_9797);
or U10236 (N_10236,N_9112,N_9934);
and U10237 (N_10237,N_9093,N_9591);
nor U10238 (N_10238,N_9040,N_9720);
xor U10239 (N_10239,N_9286,N_9263);
nand U10240 (N_10240,N_9054,N_9808);
and U10241 (N_10241,N_9016,N_9700);
or U10242 (N_10242,N_9546,N_9467);
nand U10243 (N_10243,N_9878,N_9378);
and U10244 (N_10244,N_9752,N_9920);
nand U10245 (N_10245,N_9458,N_9479);
or U10246 (N_10246,N_9025,N_9811);
xnor U10247 (N_10247,N_9921,N_9273);
xnor U10248 (N_10248,N_9636,N_9588);
nand U10249 (N_10249,N_9012,N_9145);
nor U10250 (N_10250,N_9277,N_9753);
nor U10251 (N_10251,N_9767,N_9098);
nand U10252 (N_10252,N_9894,N_9880);
or U10253 (N_10253,N_9423,N_9533);
xnor U10254 (N_10254,N_9141,N_9927);
or U10255 (N_10255,N_9295,N_9413);
or U10256 (N_10256,N_9010,N_9180);
nand U10257 (N_10257,N_9336,N_9743);
xnor U10258 (N_10258,N_9240,N_9629);
or U10259 (N_10259,N_9429,N_9819);
nor U10260 (N_10260,N_9890,N_9477);
and U10261 (N_10261,N_9388,N_9092);
xor U10262 (N_10262,N_9555,N_9450);
nor U10263 (N_10263,N_9586,N_9624);
nor U10264 (N_10264,N_9970,N_9550);
nand U10265 (N_10265,N_9446,N_9305);
or U10266 (N_10266,N_9306,N_9159);
nor U10267 (N_10267,N_9801,N_9984);
and U10268 (N_10268,N_9781,N_9457);
nand U10269 (N_10269,N_9039,N_9219);
nand U10270 (N_10270,N_9471,N_9601);
nor U10271 (N_10271,N_9658,N_9389);
xor U10272 (N_10272,N_9640,N_9033);
nand U10273 (N_10273,N_9195,N_9911);
or U10274 (N_10274,N_9108,N_9807);
xnor U10275 (N_10275,N_9868,N_9084);
nand U10276 (N_10276,N_9669,N_9838);
or U10277 (N_10277,N_9296,N_9532);
xor U10278 (N_10278,N_9069,N_9490);
and U10279 (N_10279,N_9408,N_9488);
nand U10280 (N_10280,N_9924,N_9881);
and U10281 (N_10281,N_9803,N_9963);
nand U10282 (N_10282,N_9390,N_9280);
nor U10283 (N_10283,N_9210,N_9225);
nor U10284 (N_10284,N_9929,N_9127);
or U10285 (N_10285,N_9343,N_9991);
and U10286 (N_10286,N_9081,N_9684);
nor U10287 (N_10287,N_9354,N_9661);
nor U10288 (N_10288,N_9188,N_9482);
and U10289 (N_10289,N_9052,N_9274);
and U10290 (N_10290,N_9698,N_9657);
nor U10291 (N_10291,N_9191,N_9282);
nor U10292 (N_10292,N_9951,N_9131);
nor U10293 (N_10293,N_9830,N_9645);
xnor U10294 (N_10294,N_9002,N_9831);
nand U10295 (N_10295,N_9355,N_9245);
xnor U10296 (N_10296,N_9961,N_9771);
nand U10297 (N_10297,N_9612,N_9478);
or U10298 (N_10298,N_9515,N_9508);
nand U10299 (N_10299,N_9721,N_9023);
nor U10300 (N_10300,N_9780,N_9360);
xor U10301 (N_10301,N_9433,N_9379);
nand U10302 (N_10302,N_9605,N_9185);
xor U10303 (N_10303,N_9569,N_9220);
and U10304 (N_10304,N_9158,N_9157);
xnor U10305 (N_10305,N_9005,N_9253);
xor U10306 (N_10306,N_9959,N_9017);
nor U10307 (N_10307,N_9673,N_9322);
and U10308 (N_10308,N_9814,N_9656);
nor U10309 (N_10309,N_9199,N_9474);
xnor U10310 (N_10310,N_9776,N_9668);
and U10311 (N_10311,N_9032,N_9665);
nor U10312 (N_10312,N_9056,N_9678);
nor U10313 (N_10313,N_9978,N_9901);
nand U10314 (N_10314,N_9283,N_9393);
and U10315 (N_10315,N_9048,N_9230);
and U10316 (N_10316,N_9632,N_9107);
nor U10317 (N_10317,N_9848,N_9502);
nand U10318 (N_10318,N_9285,N_9726);
xor U10319 (N_10319,N_9008,N_9135);
or U10320 (N_10320,N_9394,N_9573);
nand U10321 (N_10321,N_9603,N_9633);
and U10322 (N_10322,N_9496,N_9440);
nor U10323 (N_10323,N_9027,N_9259);
or U10324 (N_10324,N_9077,N_9037);
xnor U10325 (N_10325,N_9299,N_9007);
xor U10326 (N_10326,N_9055,N_9384);
nor U10327 (N_10327,N_9224,N_9916);
nand U10328 (N_10328,N_9615,N_9994);
nor U10329 (N_10329,N_9772,N_9203);
or U10330 (N_10330,N_9136,N_9712);
nand U10331 (N_10331,N_9338,N_9415);
xnor U10332 (N_10332,N_9368,N_9835);
or U10333 (N_10333,N_9420,N_9804);
or U10334 (N_10334,N_9685,N_9163);
and U10335 (N_10335,N_9674,N_9778);
or U10336 (N_10336,N_9850,N_9973);
and U10337 (N_10337,N_9323,N_9725);
nor U10338 (N_10338,N_9337,N_9739);
or U10339 (N_10339,N_9447,N_9443);
nand U10340 (N_10340,N_9874,N_9321);
or U10341 (N_10341,N_9859,N_9235);
and U10342 (N_10342,N_9966,N_9079);
xor U10343 (N_10343,N_9637,N_9936);
nand U10344 (N_10344,N_9297,N_9847);
nand U10345 (N_10345,N_9204,N_9667);
nor U10346 (N_10346,N_9223,N_9660);
or U10347 (N_10347,N_9528,N_9152);
and U10348 (N_10348,N_9683,N_9272);
nor U10349 (N_10349,N_9316,N_9708);
nor U10350 (N_10350,N_9100,N_9747);
and U10351 (N_10351,N_9213,N_9672);
xor U10352 (N_10352,N_9539,N_9228);
nand U10353 (N_10353,N_9981,N_9579);
or U10354 (N_10354,N_9485,N_9521);
or U10355 (N_10355,N_9239,N_9904);
nand U10356 (N_10356,N_9047,N_9536);
nor U10357 (N_10357,N_9173,N_9559);
xor U10358 (N_10358,N_9181,N_9990);
and U10359 (N_10359,N_9051,N_9749);
and U10360 (N_10360,N_9330,N_9364);
or U10361 (N_10361,N_9365,N_9790);
and U10362 (N_10362,N_9445,N_9796);
and U10363 (N_10363,N_9570,N_9845);
and U10364 (N_10364,N_9262,N_9750);
nand U10365 (N_10365,N_9462,N_9487);
or U10366 (N_10366,N_9779,N_9483);
xnor U10367 (N_10367,N_9866,N_9822);
xor U10368 (N_10368,N_9011,N_9695);
nor U10369 (N_10369,N_9581,N_9564);
and U10370 (N_10370,N_9243,N_9965);
nor U10371 (N_10371,N_9549,N_9333);
or U10372 (N_10372,N_9662,N_9397);
xnor U10373 (N_10373,N_9862,N_9817);
nor U10374 (N_10374,N_9212,N_9687);
nand U10375 (N_10375,N_9884,N_9404);
or U10376 (N_10376,N_9126,N_9129);
or U10377 (N_10377,N_9584,N_9710);
and U10378 (N_10378,N_9105,N_9626);
or U10379 (N_10379,N_9641,N_9464);
xor U10380 (N_10380,N_9307,N_9132);
nand U10381 (N_10381,N_9061,N_9441);
nor U10382 (N_10382,N_9900,N_9849);
xor U10383 (N_10383,N_9459,N_9169);
nor U10384 (N_10384,N_9745,N_9858);
and U10385 (N_10385,N_9909,N_9565);
xor U10386 (N_10386,N_9897,N_9142);
nand U10387 (N_10387,N_9997,N_9405);
and U10388 (N_10388,N_9380,N_9465);
and U10389 (N_10389,N_9925,N_9914);
nor U10390 (N_10390,N_9101,N_9992);
xor U10391 (N_10391,N_9454,N_9175);
xor U10392 (N_10392,N_9806,N_9511);
and U10393 (N_10393,N_9560,N_9891);
and U10394 (N_10394,N_9416,N_9691);
xor U10395 (N_10395,N_9252,N_9693);
xor U10396 (N_10396,N_9757,N_9643);
or U10397 (N_10397,N_9596,N_9514);
nor U10398 (N_10398,N_9554,N_9944);
nand U10399 (N_10399,N_9947,N_9495);
nand U10400 (N_10400,N_9311,N_9095);
xnor U10401 (N_10401,N_9494,N_9251);
nor U10402 (N_10402,N_9050,N_9556);
nand U10403 (N_10403,N_9247,N_9867);
and U10404 (N_10404,N_9980,N_9931);
xnor U10405 (N_10405,N_9386,N_9406);
xor U10406 (N_10406,N_9751,N_9723);
or U10407 (N_10407,N_9124,N_9329);
or U10408 (N_10408,N_9833,N_9421);
xor U10409 (N_10409,N_9190,N_9785);
or U10410 (N_10410,N_9617,N_9701);
xnor U10411 (N_10411,N_9999,N_9425);
nor U10412 (N_10412,N_9059,N_9094);
or U10413 (N_10413,N_9690,N_9576);
nor U10414 (N_10414,N_9276,N_9932);
xor U10415 (N_10415,N_9024,N_9398);
or U10416 (N_10416,N_9902,N_9899);
nor U10417 (N_10417,N_9977,N_9541);
nor U10418 (N_10418,N_9449,N_9671);
nor U10419 (N_10419,N_9269,N_9288);
or U10420 (N_10420,N_9109,N_9347);
xor U10421 (N_10421,N_9412,N_9470);
and U10422 (N_10422,N_9689,N_9509);
and U10423 (N_10423,N_9302,N_9000);
xor U10424 (N_10424,N_9020,N_9310);
nand U10425 (N_10425,N_9246,N_9842);
nand U10426 (N_10426,N_9770,N_9473);
or U10427 (N_10427,N_9324,N_9057);
xor U10428 (N_10428,N_9357,N_9125);
or U10429 (N_10429,N_9530,N_9998);
or U10430 (N_10430,N_9527,N_9529);
or U10431 (N_10431,N_9103,N_9713);
or U10432 (N_10432,N_9941,N_9256);
and U10433 (N_10433,N_9261,N_9278);
nor U10434 (N_10434,N_9049,N_9013);
nand U10435 (N_10435,N_9004,N_9791);
nor U10436 (N_10436,N_9650,N_9967);
nor U10437 (N_10437,N_9369,N_9843);
or U10438 (N_10438,N_9875,N_9407);
nor U10439 (N_10439,N_9775,N_9585);
nand U10440 (N_10440,N_9410,N_9206);
nor U10441 (N_10441,N_9815,N_9912);
xor U10442 (N_10442,N_9072,N_9553);
or U10443 (N_10443,N_9709,N_9628);
xor U10444 (N_10444,N_9249,N_9616);
nand U10445 (N_10445,N_9760,N_9825);
xnor U10446 (N_10446,N_9872,N_9949);
nor U10447 (N_10447,N_9217,N_9216);
nor U10448 (N_10448,N_9865,N_9281);
nand U10449 (N_10449,N_9493,N_9492);
nand U10450 (N_10450,N_9015,N_9969);
xor U10451 (N_10451,N_9995,N_9876);
nor U10452 (N_10452,N_9233,N_9840);
xnor U10453 (N_10453,N_9356,N_9795);
or U10454 (N_10454,N_9846,N_9832);
nand U10455 (N_10455,N_9694,N_9260);
nand U10456 (N_10456,N_9275,N_9699);
or U10457 (N_10457,N_9469,N_9153);
and U10458 (N_10458,N_9172,N_9314);
nand U10459 (N_10459,N_9958,N_9304);
xnor U10460 (N_10460,N_9070,N_9179);
and U10461 (N_10461,N_9987,N_9294);
xor U10462 (N_10462,N_9209,N_9200);
and U10463 (N_10463,N_9595,N_9938);
and U10464 (N_10464,N_9653,N_9466);
nor U10465 (N_10465,N_9505,N_9518);
nor U10466 (N_10466,N_9414,N_9996);
xnor U10467 (N_10467,N_9789,N_9298);
nor U10468 (N_10468,N_9075,N_9229);
and U10469 (N_10469,N_9562,N_9516);
and U10470 (N_10470,N_9670,N_9073);
nand U10471 (N_10471,N_9001,N_9196);
or U10472 (N_10472,N_9654,N_9436);
nor U10473 (N_10473,N_9844,N_9975);
or U10474 (N_10474,N_9501,N_9864);
nor U10475 (N_10475,N_9156,N_9373);
and U10476 (N_10476,N_9241,N_9359);
and U10477 (N_10477,N_9666,N_9110);
or U10478 (N_10478,N_9786,N_9638);
xor U10479 (N_10479,N_9320,N_9841);
or U10480 (N_10480,N_9972,N_9580);
and U10481 (N_10481,N_9117,N_9578);
and U10482 (N_10482,N_9828,N_9362);
xnor U10483 (N_10483,N_9625,N_9167);
or U10484 (N_10484,N_9773,N_9399);
and U10485 (N_10485,N_9988,N_9086);
and U10486 (N_10486,N_9782,N_9034);
nand U10487 (N_10487,N_9442,N_9538);
nor U10488 (N_10488,N_9475,N_9432);
or U10489 (N_10489,N_9300,N_9940);
xnor U10490 (N_10490,N_9707,N_9592);
or U10491 (N_10491,N_9765,N_9922);
and U10492 (N_10492,N_9370,N_9071);
or U10493 (N_10493,N_9227,N_9895);
nand U10494 (N_10494,N_9133,N_9871);
or U10495 (N_10495,N_9137,N_9067);
or U10496 (N_10496,N_9221,N_9303);
nor U10497 (N_10497,N_9794,N_9952);
nor U10498 (N_10498,N_9381,N_9648);
xnor U10499 (N_10499,N_9448,N_9326);
nand U10500 (N_10500,N_9229,N_9093);
nor U10501 (N_10501,N_9742,N_9824);
or U10502 (N_10502,N_9681,N_9048);
and U10503 (N_10503,N_9733,N_9922);
nor U10504 (N_10504,N_9558,N_9357);
xnor U10505 (N_10505,N_9888,N_9634);
nor U10506 (N_10506,N_9764,N_9898);
xor U10507 (N_10507,N_9752,N_9539);
xnor U10508 (N_10508,N_9799,N_9152);
and U10509 (N_10509,N_9725,N_9571);
or U10510 (N_10510,N_9570,N_9276);
and U10511 (N_10511,N_9348,N_9752);
or U10512 (N_10512,N_9245,N_9839);
and U10513 (N_10513,N_9592,N_9843);
xor U10514 (N_10514,N_9108,N_9262);
nor U10515 (N_10515,N_9256,N_9615);
and U10516 (N_10516,N_9690,N_9305);
nand U10517 (N_10517,N_9160,N_9960);
and U10518 (N_10518,N_9463,N_9258);
nand U10519 (N_10519,N_9111,N_9423);
and U10520 (N_10520,N_9339,N_9663);
nor U10521 (N_10521,N_9913,N_9304);
or U10522 (N_10522,N_9922,N_9916);
xnor U10523 (N_10523,N_9995,N_9960);
nand U10524 (N_10524,N_9200,N_9472);
nand U10525 (N_10525,N_9070,N_9428);
xor U10526 (N_10526,N_9965,N_9152);
nor U10527 (N_10527,N_9852,N_9632);
and U10528 (N_10528,N_9297,N_9694);
xnor U10529 (N_10529,N_9166,N_9465);
or U10530 (N_10530,N_9049,N_9078);
and U10531 (N_10531,N_9776,N_9614);
xnor U10532 (N_10532,N_9409,N_9166);
xnor U10533 (N_10533,N_9195,N_9143);
nor U10534 (N_10534,N_9163,N_9479);
xnor U10535 (N_10535,N_9046,N_9784);
nand U10536 (N_10536,N_9853,N_9011);
and U10537 (N_10537,N_9506,N_9748);
xnor U10538 (N_10538,N_9776,N_9479);
and U10539 (N_10539,N_9145,N_9046);
and U10540 (N_10540,N_9518,N_9822);
nor U10541 (N_10541,N_9940,N_9533);
nor U10542 (N_10542,N_9082,N_9124);
xnor U10543 (N_10543,N_9052,N_9980);
xor U10544 (N_10544,N_9256,N_9149);
nand U10545 (N_10545,N_9525,N_9889);
or U10546 (N_10546,N_9988,N_9020);
nand U10547 (N_10547,N_9519,N_9985);
nor U10548 (N_10548,N_9855,N_9497);
nand U10549 (N_10549,N_9112,N_9951);
xor U10550 (N_10550,N_9695,N_9101);
nand U10551 (N_10551,N_9294,N_9417);
nor U10552 (N_10552,N_9901,N_9401);
or U10553 (N_10553,N_9627,N_9940);
and U10554 (N_10554,N_9555,N_9024);
xor U10555 (N_10555,N_9537,N_9391);
nand U10556 (N_10556,N_9681,N_9008);
nor U10557 (N_10557,N_9350,N_9133);
xnor U10558 (N_10558,N_9300,N_9448);
xor U10559 (N_10559,N_9257,N_9274);
nor U10560 (N_10560,N_9786,N_9874);
or U10561 (N_10561,N_9984,N_9363);
xnor U10562 (N_10562,N_9399,N_9801);
nor U10563 (N_10563,N_9101,N_9181);
nor U10564 (N_10564,N_9109,N_9483);
and U10565 (N_10565,N_9230,N_9273);
and U10566 (N_10566,N_9172,N_9584);
nor U10567 (N_10567,N_9439,N_9094);
nor U10568 (N_10568,N_9095,N_9475);
and U10569 (N_10569,N_9241,N_9259);
or U10570 (N_10570,N_9754,N_9494);
nand U10571 (N_10571,N_9932,N_9153);
and U10572 (N_10572,N_9525,N_9320);
and U10573 (N_10573,N_9963,N_9682);
nand U10574 (N_10574,N_9817,N_9709);
nand U10575 (N_10575,N_9684,N_9996);
nor U10576 (N_10576,N_9236,N_9635);
xor U10577 (N_10577,N_9747,N_9961);
or U10578 (N_10578,N_9135,N_9013);
and U10579 (N_10579,N_9709,N_9922);
nand U10580 (N_10580,N_9507,N_9681);
and U10581 (N_10581,N_9914,N_9737);
nor U10582 (N_10582,N_9946,N_9040);
xnor U10583 (N_10583,N_9302,N_9487);
nand U10584 (N_10584,N_9060,N_9730);
nand U10585 (N_10585,N_9612,N_9500);
xor U10586 (N_10586,N_9421,N_9025);
nor U10587 (N_10587,N_9968,N_9635);
nand U10588 (N_10588,N_9951,N_9354);
nand U10589 (N_10589,N_9430,N_9596);
nand U10590 (N_10590,N_9743,N_9154);
or U10591 (N_10591,N_9782,N_9150);
xor U10592 (N_10592,N_9523,N_9640);
or U10593 (N_10593,N_9739,N_9771);
nand U10594 (N_10594,N_9689,N_9476);
nor U10595 (N_10595,N_9730,N_9933);
or U10596 (N_10596,N_9150,N_9590);
xnor U10597 (N_10597,N_9440,N_9686);
and U10598 (N_10598,N_9912,N_9414);
or U10599 (N_10599,N_9982,N_9919);
nand U10600 (N_10600,N_9095,N_9543);
or U10601 (N_10601,N_9464,N_9441);
nor U10602 (N_10602,N_9617,N_9375);
nand U10603 (N_10603,N_9049,N_9073);
and U10604 (N_10604,N_9714,N_9764);
and U10605 (N_10605,N_9197,N_9878);
or U10606 (N_10606,N_9170,N_9154);
nor U10607 (N_10607,N_9426,N_9372);
nand U10608 (N_10608,N_9939,N_9651);
xnor U10609 (N_10609,N_9611,N_9791);
or U10610 (N_10610,N_9882,N_9895);
and U10611 (N_10611,N_9056,N_9482);
nor U10612 (N_10612,N_9214,N_9891);
nor U10613 (N_10613,N_9997,N_9605);
or U10614 (N_10614,N_9730,N_9127);
and U10615 (N_10615,N_9481,N_9279);
or U10616 (N_10616,N_9377,N_9334);
nand U10617 (N_10617,N_9724,N_9141);
and U10618 (N_10618,N_9956,N_9229);
nand U10619 (N_10619,N_9874,N_9414);
nand U10620 (N_10620,N_9990,N_9009);
xnor U10621 (N_10621,N_9943,N_9881);
nand U10622 (N_10622,N_9052,N_9938);
nand U10623 (N_10623,N_9763,N_9530);
nor U10624 (N_10624,N_9247,N_9043);
or U10625 (N_10625,N_9240,N_9252);
xor U10626 (N_10626,N_9784,N_9618);
and U10627 (N_10627,N_9033,N_9944);
nand U10628 (N_10628,N_9838,N_9148);
nor U10629 (N_10629,N_9996,N_9307);
nor U10630 (N_10630,N_9090,N_9122);
or U10631 (N_10631,N_9050,N_9270);
nor U10632 (N_10632,N_9268,N_9995);
xor U10633 (N_10633,N_9216,N_9060);
and U10634 (N_10634,N_9075,N_9931);
or U10635 (N_10635,N_9139,N_9133);
xnor U10636 (N_10636,N_9038,N_9384);
nor U10637 (N_10637,N_9409,N_9174);
and U10638 (N_10638,N_9007,N_9822);
and U10639 (N_10639,N_9352,N_9110);
nor U10640 (N_10640,N_9106,N_9348);
nand U10641 (N_10641,N_9331,N_9307);
nand U10642 (N_10642,N_9436,N_9715);
nand U10643 (N_10643,N_9625,N_9711);
or U10644 (N_10644,N_9742,N_9886);
nor U10645 (N_10645,N_9619,N_9052);
and U10646 (N_10646,N_9369,N_9236);
and U10647 (N_10647,N_9539,N_9481);
nor U10648 (N_10648,N_9346,N_9687);
xor U10649 (N_10649,N_9616,N_9803);
xnor U10650 (N_10650,N_9638,N_9554);
or U10651 (N_10651,N_9712,N_9682);
nand U10652 (N_10652,N_9460,N_9789);
xor U10653 (N_10653,N_9259,N_9627);
xnor U10654 (N_10654,N_9204,N_9910);
xnor U10655 (N_10655,N_9700,N_9689);
and U10656 (N_10656,N_9293,N_9524);
nand U10657 (N_10657,N_9205,N_9785);
and U10658 (N_10658,N_9770,N_9579);
or U10659 (N_10659,N_9416,N_9865);
nand U10660 (N_10660,N_9040,N_9043);
or U10661 (N_10661,N_9942,N_9423);
nor U10662 (N_10662,N_9770,N_9550);
and U10663 (N_10663,N_9775,N_9917);
and U10664 (N_10664,N_9590,N_9024);
and U10665 (N_10665,N_9811,N_9551);
nor U10666 (N_10666,N_9598,N_9179);
nor U10667 (N_10667,N_9406,N_9550);
xnor U10668 (N_10668,N_9924,N_9298);
nand U10669 (N_10669,N_9130,N_9424);
and U10670 (N_10670,N_9633,N_9884);
and U10671 (N_10671,N_9186,N_9318);
and U10672 (N_10672,N_9002,N_9591);
or U10673 (N_10673,N_9578,N_9830);
nor U10674 (N_10674,N_9253,N_9055);
nor U10675 (N_10675,N_9779,N_9285);
nor U10676 (N_10676,N_9211,N_9151);
and U10677 (N_10677,N_9844,N_9698);
or U10678 (N_10678,N_9467,N_9592);
nand U10679 (N_10679,N_9161,N_9688);
nand U10680 (N_10680,N_9347,N_9247);
nand U10681 (N_10681,N_9406,N_9418);
xor U10682 (N_10682,N_9315,N_9152);
and U10683 (N_10683,N_9107,N_9616);
nand U10684 (N_10684,N_9257,N_9150);
xor U10685 (N_10685,N_9305,N_9114);
and U10686 (N_10686,N_9909,N_9083);
xnor U10687 (N_10687,N_9635,N_9952);
xnor U10688 (N_10688,N_9591,N_9964);
nor U10689 (N_10689,N_9876,N_9954);
and U10690 (N_10690,N_9701,N_9783);
nor U10691 (N_10691,N_9749,N_9733);
nor U10692 (N_10692,N_9688,N_9626);
and U10693 (N_10693,N_9580,N_9759);
or U10694 (N_10694,N_9391,N_9670);
nand U10695 (N_10695,N_9993,N_9879);
or U10696 (N_10696,N_9674,N_9034);
nor U10697 (N_10697,N_9925,N_9803);
and U10698 (N_10698,N_9391,N_9897);
or U10699 (N_10699,N_9172,N_9292);
nand U10700 (N_10700,N_9430,N_9829);
or U10701 (N_10701,N_9334,N_9601);
or U10702 (N_10702,N_9909,N_9969);
and U10703 (N_10703,N_9296,N_9878);
nand U10704 (N_10704,N_9362,N_9069);
nand U10705 (N_10705,N_9661,N_9375);
or U10706 (N_10706,N_9900,N_9371);
and U10707 (N_10707,N_9787,N_9115);
or U10708 (N_10708,N_9811,N_9218);
and U10709 (N_10709,N_9179,N_9786);
and U10710 (N_10710,N_9047,N_9673);
or U10711 (N_10711,N_9532,N_9928);
nor U10712 (N_10712,N_9688,N_9341);
xnor U10713 (N_10713,N_9241,N_9171);
nor U10714 (N_10714,N_9815,N_9226);
xor U10715 (N_10715,N_9249,N_9869);
nand U10716 (N_10716,N_9971,N_9457);
nand U10717 (N_10717,N_9391,N_9942);
xor U10718 (N_10718,N_9964,N_9674);
nand U10719 (N_10719,N_9060,N_9826);
or U10720 (N_10720,N_9937,N_9811);
nand U10721 (N_10721,N_9152,N_9354);
nand U10722 (N_10722,N_9280,N_9379);
or U10723 (N_10723,N_9725,N_9511);
or U10724 (N_10724,N_9552,N_9700);
or U10725 (N_10725,N_9841,N_9691);
nor U10726 (N_10726,N_9043,N_9637);
nor U10727 (N_10727,N_9280,N_9462);
nor U10728 (N_10728,N_9698,N_9509);
nand U10729 (N_10729,N_9846,N_9683);
xnor U10730 (N_10730,N_9046,N_9760);
nor U10731 (N_10731,N_9198,N_9160);
nor U10732 (N_10732,N_9745,N_9969);
xor U10733 (N_10733,N_9093,N_9026);
or U10734 (N_10734,N_9802,N_9173);
and U10735 (N_10735,N_9280,N_9249);
xnor U10736 (N_10736,N_9472,N_9499);
nand U10737 (N_10737,N_9359,N_9568);
xor U10738 (N_10738,N_9323,N_9841);
or U10739 (N_10739,N_9897,N_9090);
or U10740 (N_10740,N_9461,N_9777);
nand U10741 (N_10741,N_9908,N_9377);
xnor U10742 (N_10742,N_9284,N_9131);
nand U10743 (N_10743,N_9299,N_9192);
nor U10744 (N_10744,N_9378,N_9197);
or U10745 (N_10745,N_9495,N_9878);
xor U10746 (N_10746,N_9945,N_9581);
xnor U10747 (N_10747,N_9976,N_9235);
or U10748 (N_10748,N_9913,N_9799);
nor U10749 (N_10749,N_9663,N_9766);
nand U10750 (N_10750,N_9585,N_9168);
nor U10751 (N_10751,N_9241,N_9121);
xnor U10752 (N_10752,N_9330,N_9379);
nand U10753 (N_10753,N_9294,N_9482);
nor U10754 (N_10754,N_9329,N_9860);
and U10755 (N_10755,N_9929,N_9278);
nor U10756 (N_10756,N_9648,N_9822);
or U10757 (N_10757,N_9647,N_9178);
nand U10758 (N_10758,N_9616,N_9202);
or U10759 (N_10759,N_9091,N_9040);
nand U10760 (N_10760,N_9327,N_9259);
xor U10761 (N_10761,N_9660,N_9902);
and U10762 (N_10762,N_9916,N_9082);
or U10763 (N_10763,N_9623,N_9589);
nand U10764 (N_10764,N_9156,N_9955);
nor U10765 (N_10765,N_9659,N_9976);
nand U10766 (N_10766,N_9299,N_9444);
and U10767 (N_10767,N_9965,N_9479);
nand U10768 (N_10768,N_9433,N_9341);
or U10769 (N_10769,N_9412,N_9795);
nand U10770 (N_10770,N_9933,N_9000);
and U10771 (N_10771,N_9171,N_9760);
or U10772 (N_10772,N_9083,N_9462);
and U10773 (N_10773,N_9984,N_9337);
nand U10774 (N_10774,N_9381,N_9784);
xor U10775 (N_10775,N_9531,N_9938);
and U10776 (N_10776,N_9859,N_9425);
xnor U10777 (N_10777,N_9612,N_9396);
nand U10778 (N_10778,N_9984,N_9375);
and U10779 (N_10779,N_9155,N_9170);
and U10780 (N_10780,N_9962,N_9748);
and U10781 (N_10781,N_9872,N_9542);
and U10782 (N_10782,N_9367,N_9139);
or U10783 (N_10783,N_9009,N_9622);
nor U10784 (N_10784,N_9252,N_9496);
nor U10785 (N_10785,N_9428,N_9201);
xor U10786 (N_10786,N_9497,N_9702);
nand U10787 (N_10787,N_9246,N_9595);
or U10788 (N_10788,N_9519,N_9872);
and U10789 (N_10789,N_9722,N_9801);
and U10790 (N_10790,N_9079,N_9332);
nor U10791 (N_10791,N_9783,N_9030);
or U10792 (N_10792,N_9759,N_9257);
and U10793 (N_10793,N_9231,N_9496);
xnor U10794 (N_10794,N_9635,N_9048);
xnor U10795 (N_10795,N_9786,N_9033);
and U10796 (N_10796,N_9245,N_9231);
and U10797 (N_10797,N_9062,N_9017);
nand U10798 (N_10798,N_9194,N_9761);
nor U10799 (N_10799,N_9144,N_9838);
nor U10800 (N_10800,N_9008,N_9447);
and U10801 (N_10801,N_9726,N_9011);
xor U10802 (N_10802,N_9182,N_9471);
or U10803 (N_10803,N_9372,N_9246);
nand U10804 (N_10804,N_9458,N_9124);
nor U10805 (N_10805,N_9550,N_9489);
xor U10806 (N_10806,N_9877,N_9663);
and U10807 (N_10807,N_9000,N_9085);
and U10808 (N_10808,N_9840,N_9441);
nor U10809 (N_10809,N_9678,N_9058);
or U10810 (N_10810,N_9275,N_9015);
or U10811 (N_10811,N_9427,N_9983);
and U10812 (N_10812,N_9937,N_9906);
or U10813 (N_10813,N_9335,N_9690);
xor U10814 (N_10814,N_9707,N_9744);
or U10815 (N_10815,N_9460,N_9151);
nor U10816 (N_10816,N_9163,N_9427);
nor U10817 (N_10817,N_9991,N_9551);
xor U10818 (N_10818,N_9414,N_9316);
nor U10819 (N_10819,N_9300,N_9416);
and U10820 (N_10820,N_9524,N_9653);
nor U10821 (N_10821,N_9522,N_9753);
nand U10822 (N_10822,N_9854,N_9943);
or U10823 (N_10823,N_9478,N_9868);
and U10824 (N_10824,N_9436,N_9086);
and U10825 (N_10825,N_9555,N_9273);
nor U10826 (N_10826,N_9211,N_9222);
nand U10827 (N_10827,N_9142,N_9705);
and U10828 (N_10828,N_9258,N_9724);
and U10829 (N_10829,N_9519,N_9323);
or U10830 (N_10830,N_9609,N_9969);
nor U10831 (N_10831,N_9998,N_9824);
xnor U10832 (N_10832,N_9505,N_9694);
xnor U10833 (N_10833,N_9576,N_9203);
nand U10834 (N_10834,N_9287,N_9515);
nor U10835 (N_10835,N_9699,N_9412);
xnor U10836 (N_10836,N_9886,N_9872);
and U10837 (N_10837,N_9178,N_9378);
or U10838 (N_10838,N_9166,N_9566);
xor U10839 (N_10839,N_9886,N_9270);
and U10840 (N_10840,N_9243,N_9454);
xnor U10841 (N_10841,N_9921,N_9773);
nand U10842 (N_10842,N_9998,N_9660);
and U10843 (N_10843,N_9789,N_9847);
xnor U10844 (N_10844,N_9066,N_9757);
nand U10845 (N_10845,N_9961,N_9823);
and U10846 (N_10846,N_9158,N_9068);
nor U10847 (N_10847,N_9368,N_9082);
nor U10848 (N_10848,N_9043,N_9895);
or U10849 (N_10849,N_9646,N_9196);
and U10850 (N_10850,N_9132,N_9890);
xnor U10851 (N_10851,N_9444,N_9655);
or U10852 (N_10852,N_9521,N_9483);
or U10853 (N_10853,N_9920,N_9562);
xnor U10854 (N_10854,N_9598,N_9419);
xnor U10855 (N_10855,N_9981,N_9240);
nor U10856 (N_10856,N_9796,N_9836);
nand U10857 (N_10857,N_9634,N_9982);
or U10858 (N_10858,N_9315,N_9578);
nand U10859 (N_10859,N_9132,N_9175);
and U10860 (N_10860,N_9296,N_9629);
and U10861 (N_10861,N_9337,N_9110);
and U10862 (N_10862,N_9082,N_9169);
nor U10863 (N_10863,N_9034,N_9606);
nor U10864 (N_10864,N_9030,N_9876);
nand U10865 (N_10865,N_9035,N_9723);
and U10866 (N_10866,N_9140,N_9332);
xor U10867 (N_10867,N_9277,N_9111);
nor U10868 (N_10868,N_9778,N_9449);
nand U10869 (N_10869,N_9186,N_9742);
nor U10870 (N_10870,N_9873,N_9365);
xnor U10871 (N_10871,N_9855,N_9259);
nand U10872 (N_10872,N_9050,N_9565);
nand U10873 (N_10873,N_9061,N_9899);
nor U10874 (N_10874,N_9653,N_9815);
nand U10875 (N_10875,N_9684,N_9328);
and U10876 (N_10876,N_9423,N_9130);
nor U10877 (N_10877,N_9336,N_9143);
xor U10878 (N_10878,N_9155,N_9987);
xor U10879 (N_10879,N_9608,N_9403);
and U10880 (N_10880,N_9506,N_9080);
or U10881 (N_10881,N_9044,N_9421);
and U10882 (N_10882,N_9581,N_9663);
nand U10883 (N_10883,N_9264,N_9152);
nand U10884 (N_10884,N_9760,N_9064);
nor U10885 (N_10885,N_9693,N_9080);
xor U10886 (N_10886,N_9644,N_9865);
xor U10887 (N_10887,N_9211,N_9861);
nand U10888 (N_10888,N_9309,N_9280);
xnor U10889 (N_10889,N_9886,N_9541);
nor U10890 (N_10890,N_9923,N_9206);
or U10891 (N_10891,N_9910,N_9439);
xnor U10892 (N_10892,N_9222,N_9990);
and U10893 (N_10893,N_9682,N_9353);
nor U10894 (N_10894,N_9010,N_9587);
and U10895 (N_10895,N_9718,N_9279);
or U10896 (N_10896,N_9007,N_9779);
nor U10897 (N_10897,N_9252,N_9473);
nand U10898 (N_10898,N_9531,N_9556);
nand U10899 (N_10899,N_9177,N_9233);
nand U10900 (N_10900,N_9277,N_9843);
nand U10901 (N_10901,N_9139,N_9347);
nor U10902 (N_10902,N_9203,N_9123);
nand U10903 (N_10903,N_9875,N_9818);
or U10904 (N_10904,N_9642,N_9925);
or U10905 (N_10905,N_9788,N_9769);
xor U10906 (N_10906,N_9916,N_9002);
or U10907 (N_10907,N_9466,N_9591);
nand U10908 (N_10908,N_9496,N_9432);
nor U10909 (N_10909,N_9081,N_9846);
xnor U10910 (N_10910,N_9782,N_9976);
xor U10911 (N_10911,N_9945,N_9369);
xor U10912 (N_10912,N_9062,N_9738);
nor U10913 (N_10913,N_9635,N_9863);
or U10914 (N_10914,N_9451,N_9617);
or U10915 (N_10915,N_9626,N_9179);
nand U10916 (N_10916,N_9422,N_9448);
and U10917 (N_10917,N_9440,N_9468);
or U10918 (N_10918,N_9597,N_9527);
nor U10919 (N_10919,N_9961,N_9499);
and U10920 (N_10920,N_9887,N_9607);
xor U10921 (N_10921,N_9585,N_9583);
nand U10922 (N_10922,N_9631,N_9332);
xor U10923 (N_10923,N_9429,N_9939);
xor U10924 (N_10924,N_9736,N_9051);
xnor U10925 (N_10925,N_9971,N_9785);
and U10926 (N_10926,N_9195,N_9004);
nand U10927 (N_10927,N_9974,N_9049);
nor U10928 (N_10928,N_9818,N_9707);
nand U10929 (N_10929,N_9284,N_9719);
xnor U10930 (N_10930,N_9515,N_9111);
or U10931 (N_10931,N_9965,N_9176);
nor U10932 (N_10932,N_9401,N_9147);
xnor U10933 (N_10933,N_9273,N_9166);
nor U10934 (N_10934,N_9979,N_9514);
or U10935 (N_10935,N_9750,N_9382);
or U10936 (N_10936,N_9269,N_9742);
nor U10937 (N_10937,N_9387,N_9227);
nand U10938 (N_10938,N_9950,N_9187);
nor U10939 (N_10939,N_9297,N_9036);
and U10940 (N_10940,N_9606,N_9401);
nor U10941 (N_10941,N_9931,N_9593);
nor U10942 (N_10942,N_9823,N_9051);
nand U10943 (N_10943,N_9482,N_9243);
nor U10944 (N_10944,N_9545,N_9865);
and U10945 (N_10945,N_9228,N_9572);
or U10946 (N_10946,N_9799,N_9763);
nand U10947 (N_10947,N_9321,N_9961);
and U10948 (N_10948,N_9331,N_9620);
xor U10949 (N_10949,N_9264,N_9529);
and U10950 (N_10950,N_9071,N_9980);
xnor U10951 (N_10951,N_9032,N_9614);
xor U10952 (N_10952,N_9752,N_9202);
xor U10953 (N_10953,N_9528,N_9038);
or U10954 (N_10954,N_9217,N_9015);
and U10955 (N_10955,N_9013,N_9259);
xor U10956 (N_10956,N_9939,N_9761);
and U10957 (N_10957,N_9737,N_9552);
xor U10958 (N_10958,N_9797,N_9218);
and U10959 (N_10959,N_9284,N_9417);
and U10960 (N_10960,N_9348,N_9776);
nand U10961 (N_10961,N_9082,N_9387);
or U10962 (N_10962,N_9447,N_9762);
nand U10963 (N_10963,N_9026,N_9800);
or U10964 (N_10964,N_9723,N_9536);
nand U10965 (N_10965,N_9140,N_9180);
xnor U10966 (N_10966,N_9656,N_9323);
nand U10967 (N_10967,N_9753,N_9526);
and U10968 (N_10968,N_9875,N_9473);
nand U10969 (N_10969,N_9568,N_9081);
xor U10970 (N_10970,N_9706,N_9980);
and U10971 (N_10971,N_9861,N_9041);
xnor U10972 (N_10972,N_9286,N_9152);
nor U10973 (N_10973,N_9913,N_9541);
or U10974 (N_10974,N_9181,N_9427);
nor U10975 (N_10975,N_9772,N_9923);
xnor U10976 (N_10976,N_9367,N_9714);
and U10977 (N_10977,N_9462,N_9726);
xor U10978 (N_10978,N_9292,N_9077);
nand U10979 (N_10979,N_9340,N_9406);
nand U10980 (N_10980,N_9783,N_9627);
or U10981 (N_10981,N_9250,N_9900);
nand U10982 (N_10982,N_9939,N_9852);
or U10983 (N_10983,N_9424,N_9488);
nand U10984 (N_10984,N_9657,N_9673);
xnor U10985 (N_10985,N_9805,N_9473);
nor U10986 (N_10986,N_9963,N_9727);
or U10987 (N_10987,N_9611,N_9259);
nor U10988 (N_10988,N_9993,N_9803);
and U10989 (N_10989,N_9814,N_9606);
and U10990 (N_10990,N_9965,N_9815);
nor U10991 (N_10991,N_9764,N_9011);
nand U10992 (N_10992,N_9702,N_9291);
xor U10993 (N_10993,N_9865,N_9771);
nor U10994 (N_10994,N_9766,N_9233);
nand U10995 (N_10995,N_9865,N_9681);
nand U10996 (N_10996,N_9906,N_9738);
and U10997 (N_10997,N_9315,N_9609);
xnor U10998 (N_10998,N_9488,N_9399);
and U10999 (N_10999,N_9759,N_9089);
and U11000 (N_11000,N_10111,N_10010);
and U11001 (N_11001,N_10237,N_10796);
nor U11002 (N_11002,N_10361,N_10159);
xor U11003 (N_11003,N_10340,N_10858);
nor U11004 (N_11004,N_10203,N_10472);
or U11005 (N_11005,N_10549,N_10216);
and U11006 (N_11006,N_10798,N_10025);
nand U11007 (N_11007,N_10628,N_10031);
xor U11008 (N_11008,N_10615,N_10117);
nand U11009 (N_11009,N_10270,N_10248);
or U11010 (N_11010,N_10105,N_10928);
nor U11011 (N_11011,N_10589,N_10144);
nor U11012 (N_11012,N_10879,N_10433);
or U11013 (N_11013,N_10902,N_10636);
and U11014 (N_11014,N_10817,N_10689);
nor U11015 (N_11015,N_10850,N_10767);
or U11016 (N_11016,N_10480,N_10322);
and U11017 (N_11017,N_10191,N_10383);
and U11018 (N_11018,N_10417,N_10753);
nand U11019 (N_11019,N_10476,N_10369);
nand U11020 (N_11020,N_10202,N_10640);
xnor U11021 (N_11021,N_10930,N_10471);
nor U11022 (N_11022,N_10974,N_10279);
nand U11023 (N_11023,N_10030,N_10052);
and U11024 (N_11024,N_10578,N_10418);
or U11025 (N_11025,N_10944,N_10698);
nor U11026 (N_11026,N_10092,N_10244);
nand U11027 (N_11027,N_10078,N_10326);
and U11028 (N_11028,N_10941,N_10680);
and U11029 (N_11029,N_10749,N_10014);
or U11030 (N_11030,N_10797,N_10574);
xor U11031 (N_11031,N_10392,N_10286);
xnor U11032 (N_11032,N_10423,N_10960);
and U11033 (N_11033,N_10327,N_10737);
or U11034 (N_11034,N_10234,N_10422);
xnor U11035 (N_11035,N_10544,N_10353);
xor U11036 (N_11036,N_10534,N_10835);
xnor U11037 (N_11037,N_10171,N_10603);
and U11038 (N_11038,N_10722,N_10212);
nand U11039 (N_11039,N_10613,N_10996);
and U11040 (N_11040,N_10242,N_10320);
or U11041 (N_11041,N_10464,N_10355);
xnor U11042 (N_11042,N_10696,N_10830);
or U11043 (N_11043,N_10806,N_10113);
xor U11044 (N_11044,N_10412,N_10182);
xor U11045 (N_11045,N_10185,N_10344);
or U11046 (N_11046,N_10739,N_10206);
nand U11047 (N_11047,N_10087,N_10913);
xor U11048 (N_11048,N_10477,N_10091);
nand U11049 (N_11049,N_10110,N_10961);
nand U11050 (N_11050,N_10661,N_10777);
and U11051 (N_11051,N_10108,N_10955);
and U11052 (N_11052,N_10540,N_10588);
and U11053 (N_11053,N_10964,N_10535);
xor U11054 (N_11054,N_10808,N_10844);
xnor U11055 (N_11055,N_10869,N_10484);
nor U11056 (N_11056,N_10848,N_10559);
nor U11057 (N_11057,N_10932,N_10395);
or U11058 (N_11058,N_10391,N_10311);
xnor U11059 (N_11059,N_10424,N_10720);
or U11060 (N_11060,N_10623,N_10569);
or U11061 (N_11061,N_10883,N_10498);
or U11062 (N_11062,N_10599,N_10576);
and U11063 (N_11063,N_10218,N_10328);
nor U11064 (N_11064,N_10300,N_10343);
xor U11065 (N_11065,N_10250,N_10884);
nor U11066 (N_11066,N_10297,N_10730);
and U11067 (N_11067,N_10290,N_10004);
or U11068 (N_11068,N_10033,N_10750);
nand U11069 (N_11069,N_10979,N_10790);
or U11070 (N_11070,N_10943,N_10192);
xnor U11071 (N_11071,N_10019,N_10106);
nor U11072 (N_11072,N_10653,N_10826);
and U11073 (N_11073,N_10204,N_10533);
and U11074 (N_11074,N_10444,N_10304);
xor U11075 (N_11075,N_10002,N_10123);
or U11076 (N_11076,N_10952,N_10449);
xor U11077 (N_11077,N_10462,N_10566);
and U11078 (N_11078,N_10688,N_10428);
or U11079 (N_11079,N_10421,N_10219);
or U11080 (N_11080,N_10445,N_10515);
or U11081 (N_11081,N_10855,N_10673);
and U11082 (N_11082,N_10824,N_10486);
xnor U11083 (N_11083,N_10415,N_10781);
or U11084 (N_11084,N_10315,N_10906);
and U11085 (N_11085,N_10289,N_10865);
or U11086 (N_11086,N_10926,N_10363);
and U11087 (N_11087,N_10898,N_10285);
nand U11088 (N_11088,N_10592,N_10061);
xor U11089 (N_11089,N_10939,N_10651);
and U11090 (N_11090,N_10537,N_10342);
xnor U11091 (N_11091,N_10551,N_10312);
xor U11092 (N_11092,N_10775,N_10836);
nor U11093 (N_11093,N_10145,N_10741);
and U11094 (N_11094,N_10512,N_10178);
nand U11095 (N_11095,N_10230,N_10450);
nand U11096 (N_11096,N_10893,N_10772);
and U11097 (N_11097,N_10481,N_10530);
and U11098 (N_11098,N_10213,N_10600);
nor U11099 (N_11099,N_10210,N_10849);
and U11100 (N_11100,N_10972,N_10347);
nand U11101 (N_11101,N_10725,N_10090);
nand U11102 (N_11102,N_10967,N_10080);
xnor U11103 (N_11103,N_10372,N_10126);
nand U11104 (N_11104,N_10882,N_10293);
nand U11105 (N_11105,N_10359,N_10973);
xnor U11106 (N_11106,N_10716,N_10067);
nand U11107 (N_11107,N_10971,N_10135);
or U11108 (N_11108,N_10310,N_10386);
nor U11109 (N_11109,N_10241,N_10558);
nand U11110 (N_11110,N_10438,N_10325);
nand U11111 (N_11111,N_10373,N_10682);
and U11112 (N_11112,N_10503,N_10583);
or U11113 (N_11113,N_10497,N_10130);
nor U11114 (N_11114,N_10041,N_10837);
and U11115 (N_11115,N_10128,N_10866);
xor U11116 (N_11116,N_10246,N_10282);
or U11117 (N_11117,N_10571,N_10520);
nand U11118 (N_11118,N_10499,N_10873);
nand U11119 (N_11119,N_10389,N_10400);
nor U11120 (N_11120,N_10454,N_10924);
nor U11121 (N_11121,N_10747,N_10114);
nor U11122 (N_11122,N_10949,N_10658);
and U11123 (N_11123,N_10733,N_10555);
or U11124 (N_11124,N_10055,N_10194);
nor U11125 (N_11125,N_10984,N_10137);
nand U11126 (N_11126,N_10693,N_10351);
or U11127 (N_11127,N_10341,N_10431);
nor U11128 (N_11128,N_10662,N_10319);
nor U11129 (N_11129,N_10860,N_10539);
or U11130 (N_11130,N_10907,N_10985);
nand U11131 (N_11131,N_10629,N_10280);
or U11132 (N_11132,N_10547,N_10316);
nor U11133 (N_11133,N_10235,N_10474);
and U11134 (N_11134,N_10645,N_10803);
nor U11135 (N_11135,N_10761,N_10604);
nor U11136 (N_11136,N_10633,N_10022);
and U11137 (N_11137,N_10337,N_10575);
xor U11138 (N_11138,N_10525,N_10005);
xnor U11139 (N_11139,N_10077,N_10610);
and U11140 (N_11140,N_10778,N_10771);
or U11141 (N_11141,N_10068,N_10129);
or U11142 (N_11142,N_10915,N_10073);
nor U11143 (N_11143,N_10841,N_10284);
nand U11144 (N_11144,N_10043,N_10085);
or U11145 (N_11145,N_10082,N_10365);
nand U11146 (N_11146,N_10488,N_10265);
and U11147 (N_11147,N_10697,N_10845);
and U11148 (N_11148,N_10452,N_10529);
or U11149 (N_11149,N_10189,N_10644);
or U11150 (N_11150,N_10190,N_10614);
xnor U11151 (N_11151,N_10787,N_10788);
xnor U11152 (N_11152,N_10795,N_10469);
or U11153 (N_11153,N_10362,N_10147);
nor U11154 (N_11154,N_10302,N_10938);
and U11155 (N_11155,N_10443,N_10671);
and U11156 (N_11156,N_10721,N_10382);
and U11157 (N_11157,N_10686,N_10839);
xor U11158 (N_11158,N_10088,N_10397);
nor U11159 (N_11159,N_10852,N_10232);
and U11160 (N_11160,N_10442,N_10874);
and U11161 (N_11161,N_10903,N_10231);
xor U11162 (N_11162,N_10692,N_10676);
xor U11163 (N_11163,N_10862,N_10070);
or U11164 (N_11164,N_10263,N_10148);
or U11165 (N_11165,N_10141,N_10097);
and U11166 (N_11166,N_10880,N_10139);
nand U11167 (N_11167,N_10398,N_10485);
and U11168 (N_11168,N_10724,N_10475);
nand U11169 (N_11169,N_10410,N_10306);
xor U11170 (N_11170,N_10158,N_10799);
xor U11171 (N_11171,N_10098,N_10630);
and U11172 (N_11172,N_10162,N_10872);
xnor U11173 (N_11173,N_10432,N_10018);
nor U11174 (N_11174,N_10674,N_10995);
xor U11175 (N_11175,N_10649,N_10871);
or U11176 (N_11176,N_10762,N_10809);
nor U11177 (N_11177,N_10101,N_10396);
xor U11178 (N_11178,N_10179,N_10063);
nand U11179 (N_11179,N_10193,N_10140);
nor U11180 (N_11180,N_10991,N_10208);
or U11181 (N_11181,N_10483,N_10657);
xnor U11182 (N_11182,N_10152,N_10196);
nand U11183 (N_11183,N_10313,N_10407);
xor U11184 (N_11184,N_10411,N_10460);
xnor U11185 (N_11185,N_10380,N_10046);
nand U11186 (N_11186,N_10958,N_10201);
xnor U11187 (N_11187,N_10729,N_10586);
nand U11188 (N_11188,N_10997,N_10954);
nor U11189 (N_11189,N_10699,N_10274);
nand U11190 (N_11190,N_10172,N_10524);
nor U11191 (N_11191,N_10511,N_10582);
and U11192 (N_11192,N_10492,N_10023);
xnor U11193 (N_11193,N_10329,N_10983);
xnor U11194 (N_11194,N_10805,N_10681);
nand U11195 (N_11195,N_10323,N_10794);
nand U11196 (N_11196,N_10367,N_10715);
xnor U11197 (N_11197,N_10160,N_10154);
or U11198 (N_11198,N_10800,N_10542);
nor U11199 (N_11199,N_10834,N_10783);
and U11200 (N_11200,N_10277,N_10695);
nand U11201 (N_11201,N_10816,N_10829);
nand U11202 (N_11202,N_10912,N_10595);
xnor U11203 (N_11203,N_10252,N_10264);
nor U11204 (N_11204,N_10822,N_10751);
or U11205 (N_11205,N_10931,N_10027);
or U11206 (N_11206,N_10157,N_10670);
and U11207 (N_11207,N_10935,N_10665);
xor U11208 (N_11208,N_10593,N_10032);
xor U11209 (N_11209,N_10028,N_10654);
and U11210 (N_11210,N_10173,N_10732);
or U11211 (N_11211,N_10261,N_10756);
or U11212 (N_11212,N_10707,N_10044);
xor U11213 (N_11213,N_10434,N_10408);
and U11214 (N_11214,N_10121,N_10255);
nand U11215 (N_11215,N_10186,N_10000);
and U11216 (N_11216,N_10220,N_10618);
and U11217 (N_11217,N_10217,N_10099);
or U11218 (N_11218,N_10426,N_10647);
nand U11219 (N_11219,N_10006,N_10580);
xnor U11220 (N_11220,N_10049,N_10929);
or U11221 (N_11221,N_10225,N_10769);
xor U11222 (N_11222,N_10050,N_10562);
xor U11223 (N_11223,N_10587,N_10403);
nor U11224 (N_11224,N_10755,N_10458);
or U11225 (N_11225,N_10891,N_10532);
or U11226 (N_11226,N_10057,N_10040);
and U11227 (N_11227,N_10296,N_10885);
nand U11228 (N_11228,N_10393,N_10299);
xor U11229 (N_11229,N_10222,N_10768);
or U11230 (N_11230,N_10249,N_10784);
xor U11231 (N_11231,N_10635,N_10251);
nor U11232 (N_11232,N_10550,N_10287);
or U11233 (N_11233,N_10621,N_10664);
xor U11234 (N_11234,N_10840,N_10786);
nand U11235 (N_11235,N_10714,N_10919);
xor U11236 (N_11236,N_10655,N_10161);
xnor U11237 (N_11237,N_10905,N_10863);
nor U11238 (N_11238,N_10205,N_10404);
nor U11239 (N_11239,N_10276,N_10197);
or U11240 (N_11240,N_10861,N_10993);
or U11241 (N_11241,N_10272,N_10356);
and U11242 (N_11242,N_10667,N_10058);
xor U11243 (N_11243,N_10591,N_10579);
nor U11244 (N_11244,N_10451,N_10336);
or U11245 (N_11245,N_10473,N_10009);
nor U11246 (N_11246,N_10727,N_10598);
nand U11247 (N_11247,N_10508,N_10151);
xor U11248 (N_11248,N_10870,N_10745);
xor U11249 (N_11249,N_10703,N_10112);
and U11250 (N_11250,N_10490,N_10823);
and U11251 (N_11251,N_10257,N_10447);
or U11252 (N_11252,N_10414,N_10076);
nand U11253 (N_11253,N_10744,N_10992);
xor U11254 (N_11254,N_10352,N_10243);
and U11255 (N_11255,N_10086,N_10305);
nor U11256 (N_11256,N_10233,N_10740);
and U11257 (N_11257,N_10999,N_10368);
or U11258 (N_11258,N_10896,N_10666);
nor U11259 (N_11259,N_10072,N_10318);
nand U11260 (N_11260,N_10224,N_10229);
nand U11261 (N_11261,N_10887,N_10959);
and U11262 (N_11262,N_10247,N_10510);
xor U11263 (N_11263,N_10791,N_10927);
xnor U11264 (N_11264,N_10564,N_10487);
and U11265 (N_11265,N_10789,N_10911);
and U11266 (N_11266,N_10910,N_10782);
nor U11267 (N_11267,N_10897,N_10597);
or U11268 (N_11268,N_10026,N_10986);
nor U11269 (N_11269,N_10001,N_10275);
nand U11270 (N_11270,N_10262,N_10890);
nor U11271 (N_11271,N_10970,N_10053);
xor U11272 (N_11272,N_10461,N_10760);
nand U11273 (N_11273,N_10093,N_10214);
nor U11274 (N_11274,N_10626,N_10734);
and U11275 (N_11275,N_10301,N_10228);
and U11276 (N_11276,N_10536,N_10625);
nor U11277 (N_11277,N_10138,N_10675);
xnor U11278 (N_11278,N_10560,N_10440);
nor U11279 (N_11279,N_10641,N_10399);
or U11280 (N_11280,N_10051,N_10843);
or U11281 (N_11281,N_10254,N_10075);
nand U11282 (N_11282,N_10677,N_10375);
and U11283 (N_11283,N_10115,N_10008);
and U11284 (N_11284,N_10377,N_10917);
nand U11285 (N_11285,N_10493,N_10268);
or U11286 (N_11286,N_10925,N_10267);
and U11287 (N_11287,N_10556,N_10209);
xor U11288 (N_11288,N_10916,N_10062);
nand U11289 (N_11289,N_10757,N_10457);
nand U11290 (N_11290,N_10853,N_10543);
nand U11291 (N_11291,N_10705,N_10495);
xnor U11292 (N_11292,N_10184,N_10831);
or U11293 (N_11293,N_10687,N_10012);
and U11294 (N_11294,N_10521,N_10283);
nand U11295 (N_11295,N_10957,N_10933);
nor U11296 (N_11296,N_10846,N_10468);
and U11297 (N_11297,N_10909,N_10708);
and U11298 (N_11298,N_10669,N_10642);
and U11299 (N_11299,N_10709,N_10812);
and U11300 (N_11300,N_10020,N_10357);
nor U11301 (N_11301,N_10859,N_10616);
xor U11302 (N_11302,N_10281,N_10940);
and U11303 (N_11303,N_10548,N_10465);
nand U11304 (N_11304,N_10684,N_10828);
and U11305 (N_11305,N_10854,N_10420);
xnor U11306 (N_11306,N_10785,N_10968);
nand U11307 (N_11307,N_10758,N_10198);
nor U11308 (N_11308,N_10446,N_10015);
or U11309 (N_11309,N_10253,N_10934);
xor U11310 (N_11310,N_10333,N_10385);
xor U11311 (N_11311,N_10491,N_10672);
nand U11312 (N_11312,N_10164,N_10016);
xor U11313 (N_11313,N_10726,N_10617);
or U11314 (N_11314,N_10131,N_10109);
and U11315 (N_11315,N_10683,N_10719);
or U11316 (N_11316,N_10314,N_10379);
or U11317 (N_11317,N_10700,N_10565);
xor U11318 (N_11318,N_10723,N_10605);
and U11319 (N_11319,N_10064,N_10042);
xor U11320 (N_11320,N_10466,N_10429);
nor U11321 (N_11321,N_10436,N_10266);
xnor U11322 (N_11322,N_10168,N_10288);
xor U11323 (N_11323,N_10563,N_10011);
and U11324 (N_11324,N_10814,N_10338);
nand U11325 (N_11325,N_10833,N_10942);
and U11326 (N_11326,N_10013,N_10779);
nand U11327 (N_11327,N_10561,N_10608);
nand U11328 (N_11328,N_10083,N_10081);
nand U11329 (N_11329,N_10624,N_10066);
or U11330 (N_11330,N_10260,N_10679);
xnor U11331 (N_11331,N_10975,N_10153);
nor U11332 (N_11332,N_10923,N_10427);
and U11333 (N_11333,N_10065,N_10573);
nor U11334 (N_11334,N_10951,N_10619);
or U11335 (N_11335,N_10036,N_10962);
xnor U11336 (N_11336,N_10948,N_10136);
or U11337 (N_11337,N_10811,N_10308);
or U11338 (N_11338,N_10743,N_10394);
xnor U11339 (N_11339,N_10663,N_10611);
and U11340 (N_11340,N_10646,N_10609);
or U11341 (N_11341,N_10994,N_10878);
nor U11342 (N_11342,N_10346,N_10819);
nand U11343 (N_11343,N_10501,N_10425);
nand U11344 (N_11344,N_10764,N_10736);
nand U11345 (N_11345,N_10505,N_10701);
nand U11346 (N_11346,N_10376,N_10378);
or U11347 (N_11347,N_10084,N_10594);
nand U11348 (N_11348,N_10691,N_10601);
nor U11349 (N_11349,N_10572,N_10345);
or U11350 (N_11350,N_10401,N_10731);
or U11351 (N_11351,N_10102,N_10079);
and U11352 (N_11352,N_10133,N_10045);
nand U11353 (N_11353,N_10119,N_10867);
nand U11354 (N_11354,N_10978,N_10374);
xnor U11355 (N_11355,N_10459,N_10419);
nand U11356 (N_11356,N_10792,N_10335);
nand U11357 (N_11357,N_10409,N_10364);
xnor U11358 (N_11358,N_10895,N_10331);
nor U11359 (N_11359,N_10478,N_10069);
or U11360 (N_11360,N_10226,N_10437);
nand U11361 (N_11361,N_10095,N_10766);
xnor U11362 (N_11362,N_10528,N_10349);
nand U11363 (N_11363,N_10966,N_10965);
nand U11364 (N_11364,N_10856,N_10504);
nand U11365 (N_11365,N_10463,N_10238);
nand U11366 (N_11366,N_10034,N_10953);
xor U11367 (N_11367,N_10039,N_10292);
xor U11368 (N_11368,N_10514,N_10513);
xnor U11369 (N_11369,N_10339,N_10384);
and U11370 (N_11370,N_10763,N_10711);
and U11371 (N_11371,N_10754,N_10522);
nor U11372 (N_11372,N_10712,N_10652);
or U11373 (N_11373,N_10988,N_10236);
nand U11374 (N_11374,N_10195,N_10494);
nor U11375 (N_11375,N_10746,N_10294);
nand U11376 (N_11376,N_10980,N_10321);
xor U11377 (N_11377,N_10825,N_10334);
or U11378 (N_11378,N_10937,N_10581);
and U11379 (N_11379,N_10188,N_10908);
xor U11380 (N_11380,N_10324,N_10413);
nand U11381 (N_11381,N_10567,N_10538);
nor U11382 (N_11382,N_10877,N_10632);
or U11383 (N_11383,N_10875,N_10489);
or U11384 (N_11384,N_10557,N_10441);
nand U11385 (N_11385,N_10899,N_10143);
and U11386 (N_11386,N_10998,N_10024);
or U11387 (N_11387,N_10029,N_10596);
nor U11388 (N_11388,N_10804,N_10273);
xor U11389 (N_11389,N_10969,N_10470);
nor U11390 (N_11390,N_10659,N_10060);
or U11391 (N_11391,N_10259,N_10456);
or U11392 (N_11392,N_10627,N_10602);
or U11393 (N_11393,N_10183,N_10388);
nand U11394 (N_11394,N_10668,N_10295);
nand U11395 (N_11395,N_10568,N_10718);
or U11396 (N_11396,N_10634,N_10821);
nand U11397 (N_11397,N_10832,N_10134);
xnor U11398 (N_11398,N_10759,N_10370);
or U11399 (N_11399,N_10527,N_10155);
or U11400 (N_11400,N_10765,N_10947);
and U11401 (N_11401,N_10976,N_10650);
nor U11402 (N_11402,N_10163,N_10150);
xnor U11403 (N_11403,N_10793,N_10735);
or U11404 (N_11404,N_10227,N_10606);
nand U11405 (N_11405,N_10348,N_10054);
or U11406 (N_11406,N_10059,N_10207);
nor U11407 (N_11407,N_10554,N_10223);
nand U11408 (N_11408,N_10620,N_10774);
nand U11409 (N_11409,N_10502,N_10118);
nand U11410 (N_11410,N_10922,N_10801);
nor U11411 (N_11411,N_10981,N_10936);
xnor U11412 (N_11412,N_10309,N_10678);
and U11413 (N_11413,N_10914,N_10813);
and U11414 (N_11414,N_10950,N_10330);
nand U11415 (N_11415,N_10851,N_10156);
and U11416 (N_11416,N_10094,N_10888);
xor U11417 (N_11417,N_10256,N_10728);
nand U11418 (N_11418,N_10546,N_10694);
nor U11419 (N_11419,N_10946,N_10876);
and U11420 (N_11420,N_10802,N_10815);
nor U11421 (N_11421,N_10584,N_10071);
nor U11422 (N_11422,N_10531,N_10149);
nand U11423 (N_11423,N_10577,N_10982);
and U11424 (N_11424,N_10738,N_10142);
xor U11425 (N_11425,N_10901,N_10245);
nand U11426 (N_11426,N_10945,N_10643);
and U11427 (N_11427,N_10430,N_10035);
nand U11428 (N_11428,N_10211,N_10176);
xnor U11429 (N_11429,N_10387,N_10350);
or U11430 (N_11430,N_10169,N_10406);
nand U11431 (N_11431,N_10631,N_10639);
xnor U11432 (N_11432,N_10089,N_10107);
nand U11433 (N_11433,N_10298,N_10713);
or U11434 (N_11434,N_10990,N_10904);
or U11435 (N_11435,N_10748,N_10167);
or U11436 (N_11436,N_10900,N_10240);
and U11437 (N_11437,N_10048,N_10977);
nand U11438 (N_11438,N_10810,N_10607);
or U11439 (N_11439,N_10637,N_10100);
nor U11440 (N_11440,N_10047,N_10056);
and U11441 (N_11441,N_10989,N_10199);
nand U11442 (N_11442,N_10770,N_10889);
and U11443 (N_11443,N_10366,N_10455);
xor U11444 (N_11444,N_10007,N_10405);
nand U11445 (N_11445,N_10170,N_10818);
or U11446 (N_11446,N_10200,N_10660);
xnor U11447 (N_11447,N_10921,N_10892);
or U11448 (N_11448,N_10706,N_10622);
nand U11449 (N_11449,N_10710,N_10165);
nand U11450 (N_11450,N_10125,N_10827);
or U11451 (N_11451,N_10506,N_10881);
or U11452 (N_11452,N_10479,N_10552);
xor U11453 (N_11453,N_10122,N_10180);
nand U11454 (N_11454,N_10894,N_10868);
nand U11455 (N_11455,N_10500,N_10752);
or U11456 (N_11456,N_10120,N_10857);
xor U11457 (N_11457,N_10656,N_10271);
and U11458 (N_11458,N_10017,N_10685);
xor U11459 (N_11459,N_10003,N_10104);
nor U11460 (N_11460,N_10402,N_10453);
nor U11461 (N_11461,N_10354,N_10864);
or U11462 (N_11462,N_10371,N_10585);
nand U11463 (N_11463,N_10358,N_10074);
nor U11464 (N_11464,N_10303,N_10987);
nor U11465 (N_11465,N_10612,N_10518);
or U11466 (N_11466,N_10590,N_10291);
xor U11467 (N_11467,N_10381,N_10776);
and U11468 (N_11468,N_10842,N_10742);
and U11469 (N_11469,N_10096,N_10448);
or U11470 (N_11470,N_10416,N_10127);
nand U11471 (N_11471,N_10918,N_10038);
nor U11472 (N_11472,N_10239,N_10648);
nor U11473 (N_11473,N_10482,N_10963);
xor U11474 (N_11474,N_10702,N_10116);
or U11475 (N_11475,N_10526,N_10439);
nand U11476 (N_11476,N_10435,N_10807);
or U11477 (N_11477,N_10146,N_10269);
and U11478 (N_11478,N_10545,N_10780);
and U11479 (N_11479,N_10509,N_10517);
xor U11480 (N_11480,N_10177,N_10317);
nor U11481 (N_11481,N_10496,N_10773);
nand U11482 (N_11482,N_10174,N_10175);
or U11483 (N_11483,N_10181,N_10956);
xor U11484 (N_11484,N_10886,N_10278);
and U11485 (N_11485,N_10507,N_10541);
and U11486 (N_11486,N_10221,N_10553);
nand U11487 (N_11487,N_10332,N_10166);
or U11488 (N_11488,N_10519,N_10307);
and U11489 (N_11489,N_10103,N_10704);
xnor U11490 (N_11490,N_10690,N_10820);
or U11491 (N_11491,N_10920,N_10187);
nand U11492 (N_11492,N_10037,N_10847);
or U11493 (N_11493,N_10467,N_10516);
xnor U11494 (N_11494,N_10717,N_10021);
nor U11495 (N_11495,N_10638,N_10570);
and U11496 (N_11496,N_10258,N_10523);
nor U11497 (N_11497,N_10124,N_10215);
and U11498 (N_11498,N_10390,N_10132);
or U11499 (N_11499,N_10360,N_10838);
nand U11500 (N_11500,N_10097,N_10452);
xor U11501 (N_11501,N_10939,N_10729);
or U11502 (N_11502,N_10965,N_10336);
or U11503 (N_11503,N_10985,N_10028);
and U11504 (N_11504,N_10877,N_10732);
xnor U11505 (N_11505,N_10037,N_10107);
and U11506 (N_11506,N_10657,N_10497);
nor U11507 (N_11507,N_10204,N_10138);
and U11508 (N_11508,N_10064,N_10114);
nor U11509 (N_11509,N_10964,N_10528);
nor U11510 (N_11510,N_10454,N_10721);
or U11511 (N_11511,N_10859,N_10047);
xnor U11512 (N_11512,N_10949,N_10609);
nor U11513 (N_11513,N_10382,N_10006);
nand U11514 (N_11514,N_10835,N_10276);
nand U11515 (N_11515,N_10740,N_10710);
nand U11516 (N_11516,N_10157,N_10037);
xor U11517 (N_11517,N_10099,N_10489);
and U11518 (N_11518,N_10407,N_10128);
xor U11519 (N_11519,N_10989,N_10522);
xor U11520 (N_11520,N_10560,N_10746);
nor U11521 (N_11521,N_10448,N_10863);
nand U11522 (N_11522,N_10813,N_10163);
or U11523 (N_11523,N_10743,N_10337);
or U11524 (N_11524,N_10810,N_10935);
nand U11525 (N_11525,N_10216,N_10480);
or U11526 (N_11526,N_10022,N_10366);
nor U11527 (N_11527,N_10774,N_10145);
nor U11528 (N_11528,N_10676,N_10632);
xor U11529 (N_11529,N_10002,N_10610);
xnor U11530 (N_11530,N_10487,N_10418);
nand U11531 (N_11531,N_10107,N_10256);
nor U11532 (N_11532,N_10853,N_10224);
xnor U11533 (N_11533,N_10389,N_10762);
and U11534 (N_11534,N_10774,N_10804);
or U11535 (N_11535,N_10149,N_10536);
and U11536 (N_11536,N_10605,N_10718);
or U11537 (N_11537,N_10860,N_10703);
nand U11538 (N_11538,N_10159,N_10400);
nor U11539 (N_11539,N_10431,N_10826);
nor U11540 (N_11540,N_10747,N_10323);
and U11541 (N_11541,N_10666,N_10532);
xnor U11542 (N_11542,N_10923,N_10470);
xor U11543 (N_11543,N_10809,N_10325);
xor U11544 (N_11544,N_10994,N_10047);
xor U11545 (N_11545,N_10838,N_10020);
or U11546 (N_11546,N_10444,N_10681);
xnor U11547 (N_11547,N_10301,N_10497);
and U11548 (N_11548,N_10181,N_10701);
nor U11549 (N_11549,N_10227,N_10488);
and U11550 (N_11550,N_10718,N_10229);
and U11551 (N_11551,N_10117,N_10836);
and U11552 (N_11552,N_10847,N_10418);
or U11553 (N_11553,N_10647,N_10525);
nand U11554 (N_11554,N_10310,N_10224);
xnor U11555 (N_11555,N_10328,N_10671);
nand U11556 (N_11556,N_10250,N_10966);
and U11557 (N_11557,N_10029,N_10247);
nor U11558 (N_11558,N_10096,N_10681);
and U11559 (N_11559,N_10498,N_10707);
nand U11560 (N_11560,N_10750,N_10665);
xnor U11561 (N_11561,N_10858,N_10600);
and U11562 (N_11562,N_10183,N_10977);
and U11563 (N_11563,N_10479,N_10159);
nor U11564 (N_11564,N_10226,N_10676);
or U11565 (N_11565,N_10995,N_10027);
and U11566 (N_11566,N_10073,N_10676);
and U11567 (N_11567,N_10878,N_10381);
nand U11568 (N_11568,N_10210,N_10561);
xnor U11569 (N_11569,N_10136,N_10776);
nor U11570 (N_11570,N_10946,N_10090);
nor U11571 (N_11571,N_10501,N_10875);
or U11572 (N_11572,N_10927,N_10790);
xnor U11573 (N_11573,N_10540,N_10508);
nand U11574 (N_11574,N_10381,N_10108);
xor U11575 (N_11575,N_10701,N_10948);
nand U11576 (N_11576,N_10898,N_10681);
xor U11577 (N_11577,N_10700,N_10770);
nand U11578 (N_11578,N_10588,N_10016);
and U11579 (N_11579,N_10344,N_10843);
and U11580 (N_11580,N_10013,N_10286);
nor U11581 (N_11581,N_10870,N_10635);
or U11582 (N_11582,N_10673,N_10937);
and U11583 (N_11583,N_10549,N_10076);
or U11584 (N_11584,N_10869,N_10851);
nand U11585 (N_11585,N_10012,N_10070);
and U11586 (N_11586,N_10539,N_10180);
xor U11587 (N_11587,N_10402,N_10915);
and U11588 (N_11588,N_10881,N_10315);
or U11589 (N_11589,N_10063,N_10417);
nor U11590 (N_11590,N_10579,N_10915);
or U11591 (N_11591,N_10993,N_10307);
xnor U11592 (N_11592,N_10113,N_10796);
nand U11593 (N_11593,N_10214,N_10222);
or U11594 (N_11594,N_10491,N_10894);
or U11595 (N_11595,N_10896,N_10417);
or U11596 (N_11596,N_10742,N_10442);
xnor U11597 (N_11597,N_10094,N_10278);
xnor U11598 (N_11598,N_10290,N_10183);
nand U11599 (N_11599,N_10193,N_10430);
nand U11600 (N_11600,N_10178,N_10002);
and U11601 (N_11601,N_10304,N_10366);
xnor U11602 (N_11602,N_10062,N_10178);
and U11603 (N_11603,N_10946,N_10288);
or U11604 (N_11604,N_10384,N_10959);
nand U11605 (N_11605,N_10864,N_10736);
xnor U11606 (N_11606,N_10850,N_10197);
nand U11607 (N_11607,N_10111,N_10519);
and U11608 (N_11608,N_10741,N_10285);
or U11609 (N_11609,N_10495,N_10270);
xnor U11610 (N_11610,N_10396,N_10265);
and U11611 (N_11611,N_10778,N_10356);
nor U11612 (N_11612,N_10646,N_10708);
and U11613 (N_11613,N_10853,N_10686);
xnor U11614 (N_11614,N_10074,N_10707);
and U11615 (N_11615,N_10350,N_10140);
or U11616 (N_11616,N_10222,N_10265);
or U11617 (N_11617,N_10548,N_10271);
nor U11618 (N_11618,N_10347,N_10371);
nand U11619 (N_11619,N_10375,N_10647);
xor U11620 (N_11620,N_10163,N_10676);
and U11621 (N_11621,N_10716,N_10109);
and U11622 (N_11622,N_10684,N_10980);
nand U11623 (N_11623,N_10172,N_10596);
and U11624 (N_11624,N_10823,N_10563);
or U11625 (N_11625,N_10330,N_10124);
nor U11626 (N_11626,N_10021,N_10598);
xor U11627 (N_11627,N_10809,N_10127);
nand U11628 (N_11628,N_10604,N_10426);
nand U11629 (N_11629,N_10262,N_10133);
xor U11630 (N_11630,N_10499,N_10571);
and U11631 (N_11631,N_10070,N_10628);
and U11632 (N_11632,N_10382,N_10377);
nand U11633 (N_11633,N_10066,N_10620);
and U11634 (N_11634,N_10589,N_10898);
xor U11635 (N_11635,N_10445,N_10062);
nand U11636 (N_11636,N_10463,N_10930);
nand U11637 (N_11637,N_10988,N_10370);
and U11638 (N_11638,N_10377,N_10422);
nand U11639 (N_11639,N_10202,N_10327);
xor U11640 (N_11640,N_10555,N_10479);
or U11641 (N_11641,N_10538,N_10681);
or U11642 (N_11642,N_10866,N_10238);
xor U11643 (N_11643,N_10669,N_10334);
and U11644 (N_11644,N_10450,N_10822);
xnor U11645 (N_11645,N_10680,N_10898);
or U11646 (N_11646,N_10809,N_10367);
nor U11647 (N_11647,N_10820,N_10628);
xor U11648 (N_11648,N_10799,N_10411);
nand U11649 (N_11649,N_10462,N_10397);
and U11650 (N_11650,N_10345,N_10963);
and U11651 (N_11651,N_10996,N_10825);
or U11652 (N_11652,N_10160,N_10480);
xor U11653 (N_11653,N_10545,N_10971);
or U11654 (N_11654,N_10296,N_10108);
and U11655 (N_11655,N_10754,N_10413);
xor U11656 (N_11656,N_10281,N_10259);
nor U11657 (N_11657,N_10026,N_10876);
xor U11658 (N_11658,N_10245,N_10842);
xor U11659 (N_11659,N_10847,N_10250);
nor U11660 (N_11660,N_10580,N_10728);
or U11661 (N_11661,N_10993,N_10296);
xor U11662 (N_11662,N_10530,N_10453);
xor U11663 (N_11663,N_10698,N_10999);
xnor U11664 (N_11664,N_10472,N_10571);
xnor U11665 (N_11665,N_10223,N_10810);
or U11666 (N_11666,N_10554,N_10275);
and U11667 (N_11667,N_10560,N_10289);
nor U11668 (N_11668,N_10165,N_10557);
xor U11669 (N_11669,N_10217,N_10944);
nor U11670 (N_11670,N_10414,N_10401);
xnor U11671 (N_11671,N_10689,N_10185);
and U11672 (N_11672,N_10920,N_10909);
xnor U11673 (N_11673,N_10444,N_10319);
nor U11674 (N_11674,N_10453,N_10008);
nor U11675 (N_11675,N_10692,N_10006);
and U11676 (N_11676,N_10395,N_10034);
nor U11677 (N_11677,N_10710,N_10879);
nor U11678 (N_11678,N_10353,N_10650);
nor U11679 (N_11679,N_10007,N_10450);
and U11680 (N_11680,N_10639,N_10030);
xor U11681 (N_11681,N_10022,N_10398);
nor U11682 (N_11682,N_10006,N_10277);
and U11683 (N_11683,N_10385,N_10566);
nand U11684 (N_11684,N_10741,N_10872);
or U11685 (N_11685,N_10498,N_10124);
xor U11686 (N_11686,N_10493,N_10606);
nand U11687 (N_11687,N_10859,N_10833);
or U11688 (N_11688,N_10157,N_10981);
xnor U11689 (N_11689,N_10984,N_10430);
nor U11690 (N_11690,N_10484,N_10642);
nor U11691 (N_11691,N_10536,N_10147);
and U11692 (N_11692,N_10375,N_10143);
nand U11693 (N_11693,N_10057,N_10133);
and U11694 (N_11694,N_10462,N_10945);
nor U11695 (N_11695,N_10738,N_10579);
and U11696 (N_11696,N_10789,N_10229);
nor U11697 (N_11697,N_10007,N_10156);
xnor U11698 (N_11698,N_10489,N_10501);
and U11699 (N_11699,N_10424,N_10785);
or U11700 (N_11700,N_10364,N_10317);
nand U11701 (N_11701,N_10959,N_10293);
nand U11702 (N_11702,N_10335,N_10182);
and U11703 (N_11703,N_10163,N_10674);
xnor U11704 (N_11704,N_10052,N_10767);
and U11705 (N_11705,N_10441,N_10150);
nand U11706 (N_11706,N_10517,N_10265);
nor U11707 (N_11707,N_10280,N_10740);
nor U11708 (N_11708,N_10746,N_10315);
or U11709 (N_11709,N_10294,N_10270);
and U11710 (N_11710,N_10466,N_10632);
nand U11711 (N_11711,N_10675,N_10377);
nor U11712 (N_11712,N_10367,N_10936);
and U11713 (N_11713,N_10877,N_10917);
or U11714 (N_11714,N_10048,N_10698);
nor U11715 (N_11715,N_10501,N_10513);
nor U11716 (N_11716,N_10977,N_10009);
or U11717 (N_11717,N_10034,N_10266);
nand U11718 (N_11718,N_10629,N_10785);
nand U11719 (N_11719,N_10497,N_10818);
nor U11720 (N_11720,N_10634,N_10967);
xor U11721 (N_11721,N_10912,N_10563);
or U11722 (N_11722,N_10992,N_10681);
nand U11723 (N_11723,N_10656,N_10426);
nand U11724 (N_11724,N_10660,N_10927);
and U11725 (N_11725,N_10396,N_10337);
or U11726 (N_11726,N_10225,N_10571);
nand U11727 (N_11727,N_10388,N_10338);
nand U11728 (N_11728,N_10828,N_10340);
or U11729 (N_11729,N_10193,N_10155);
xnor U11730 (N_11730,N_10313,N_10795);
and U11731 (N_11731,N_10796,N_10991);
and U11732 (N_11732,N_10744,N_10043);
nand U11733 (N_11733,N_10560,N_10631);
nor U11734 (N_11734,N_10823,N_10436);
or U11735 (N_11735,N_10882,N_10611);
xor U11736 (N_11736,N_10865,N_10559);
nor U11737 (N_11737,N_10281,N_10638);
or U11738 (N_11738,N_10494,N_10326);
or U11739 (N_11739,N_10604,N_10376);
and U11740 (N_11740,N_10195,N_10701);
xnor U11741 (N_11741,N_10596,N_10916);
and U11742 (N_11742,N_10396,N_10223);
or U11743 (N_11743,N_10381,N_10913);
and U11744 (N_11744,N_10889,N_10276);
xor U11745 (N_11745,N_10352,N_10276);
and U11746 (N_11746,N_10084,N_10425);
nor U11747 (N_11747,N_10152,N_10113);
or U11748 (N_11748,N_10727,N_10063);
and U11749 (N_11749,N_10849,N_10820);
and U11750 (N_11750,N_10081,N_10950);
and U11751 (N_11751,N_10261,N_10490);
and U11752 (N_11752,N_10469,N_10969);
xor U11753 (N_11753,N_10317,N_10811);
and U11754 (N_11754,N_10773,N_10956);
nor U11755 (N_11755,N_10370,N_10747);
xnor U11756 (N_11756,N_10368,N_10294);
or U11757 (N_11757,N_10764,N_10576);
xor U11758 (N_11758,N_10577,N_10553);
or U11759 (N_11759,N_10515,N_10944);
and U11760 (N_11760,N_10880,N_10907);
nor U11761 (N_11761,N_10095,N_10694);
xor U11762 (N_11762,N_10735,N_10804);
nand U11763 (N_11763,N_10284,N_10156);
nor U11764 (N_11764,N_10106,N_10613);
nor U11765 (N_11765,N_10884,N_10569);
xor U11766 (N_11766,N_10304,N_10404);
xor U11767 (N_11767,N_10146,N_10358);
nand U11768 (N_11768,N_10087,N_10428);
nand U11769 (N_11769,N_10300,N_10067);
nor U11770 (N_11770,N_10836,N_10580);
or U11771 (N_11771,N_10290,N_10777);
nand U11772 (N_11772,N_10953,N_10005);
nand U11773 (N_11773,N_10647,N_10378);
xor U11774 (N_11774,N_10283,N_10284);
or U11775 (N_11775,N_10891,N_10995);
and U11776 (N_11776,N_10673,N_10497);
nand U11777 (N_11777,N_10487,N_10671);
or U11778 (N_11778,N_10724,N_10410);
nor U11779 (N_11779,N_10033,N_10189);
and U11780 (N_11780,N_10439,N_10615);
nand U11781 (N_11781,N_10645,N_10635);
xor U11782 (N_11782,N_10086,N_10930);
xnor U11783 (N_11783,N_10943,N_10774);
or U11784 (N_11784,N_10276,N_10530);
nor U11785 (N_11785,N_10062,N_10792);
nor U11786 (N_11786,N_10766,N_10858);
xnor U11787 (N_11787,N_10336,N_10412);
nand U11788 (N_11788,N_10494,N_10062);
and U11789 (N_11789,N_10936,N_10419);
xnor U11790 (N_11790,N_10567,N_10095);
xor U11791 (N_11791,N_10065,N_10721);
xnor U11792 (N_11792,N_10313,N_10383);
or U11793 (N_11793,N_10266,N_10010);
nand U11794 (N_11794,N_10337,N_10334);
xor U11795 (N_11795,N_10713,N_10721);
xnor U11796 (N_11796,N_10071,N_10948);
nor U11797 (N_11797,N_10714,N_10629);
nand U11798 (N_11798,N_10784,N_10148);
nor U11799 (N_11799,N_10083,N_10789);
and U11800 (N_11800,N_10886,N_10865);
nand U11801 (N_11801,N_10489,N_10174);
nor U11802 (N_11802,N_10846,N_10363);
and U11803 (N_11803,N_10042,N_10274);
and U11804 (N_11804,N_10094,N_10668);
xor U11805 (N_11805,N_10895,N_10037);
xor U11806 (N_11806,N_10421,N_10776);
nor U11807 (N_11807,N_10398,N_10215);
xnor U11808 (N_11808,N_10956,N_10571);
or U11809 (N_11809,N_10685,N_10248);
nor U11810 (N_11810,N_10938,N_10206);
nand U11811 (N_11811,N_10765,N_10480);
nor U11812 (N_11812,N_10661,N_10605);
or U11813 (N_11813,N_10085,N_10517);
xnor U11814 (N_11814,N_10994,N_10446);
nand U11815 (N_11815,N_10006,N_10263);
xor U11816 (N_11816,N_10058,N_10008);
and U11817 (N_11817,N_10866,N_10284);
nand U11818 (N_11818,N_10233,N_10696);
xor U11819 (N_11819,N_10221,N_10917);
and U11820 (N_11820,N_10420,N_10631);
nor U11821 (N_11821,N_10833,N_10858);
nand U11822 (N_11822,N_10521,N_10513);
or U11823 (N_11823,N_10785,N_10766);
nor U11824 (N_11824,N_10602,N_10282);
or U11825 (N_11825,N_10878,N_10523);
xor U11826 (N_11826,N_10780,N_10681);
and U11827 (N_11827,N_10030,N_10099);
or U11828 (N_11828,N_10361,N_10216);
and U11829 (N_11829,N_10462,N_10351);
xor U11830 (N_11830,N_10702,N_10051);
xor U11831 (N_11831,N_10673,N_10329);
xnor U11832 (N_11832,N_10746,N_10052);
nor U11833 (N_11833,N_10643,N_10805);
nand U11834 (N_11834,N_10290,N_10502);
xor U11835 (N_11835,N_10523,N_10343);
nand U11836 (N_11836,N_10937,N_10172);
or U11837 (N_11837,N_10049,N_10685);
nand U11838 (N_11838,N_10910,N_10693);
and U11839 (N_11839,N_10738,N_10907);
or U11840 (N_11840,N_10576,N_10451);
xnor U11841 (N_11841,N_10453,N_10097);
or U11842 (N_11842,N_10653,N_10188);
or U11843 (N_11843,N_10527,N_10030);
or U11844 (N_11844,N_10608,N_10574);
nand U11845 (N_11845,N_10490,N_10392);
and U11846 (N_11846,N_10496,N_10252);
and U11847 (N_11847,N_10782,N_10646);
nor U11848 (N_11848,N_10467,N_10675);
or U11849 (N_11849,N_10121,N_10312);
nand U11850 (N_11850,N_10755,N_10528);
nand U11851 (N_11851,N_10454,N_10927);
nor U11852 (N_11852,N_10733,N_10505);
nand U11853 (N_11853,N_10571,N_10404);
and U11854 (N_11854,N_10755,N_10293);
and U11855 (N_11855,N_10078,N_10941);
xor U11856 (N_11856,N_10498,N_10945);
nor U11857 (N_11857,N_10222,N_10941);
nor U11858 (N_11858,N_10527,N_10738);
nand U11859 (N_11859,N_10532,N_10728);
or U11860 (N_11860,N_10157,N_10746);
nor U11861 (N_11861,N_10280,N_10157);
nand U11862 (N_11862,N_10002,N_10442);
xnor U11863 (N_11863,N_10965,N_10557);
and U11864 (N_11864,N_10339,N_10698);
nand U11865 (N_11865,N_10112,N_10438);
xnor U11866 (N_11866,N_10918,N_10818);
or U11867 (N_11867,N_10236,N_10148);
or U11868 (N_11868,N_10746,N_10249);
and U11869 (N_11869,N_10555,N_10177);
nor U11870 (N_11870,N_10559,N_10047);
or U11871 (N_11871,N_10723,N_10996);
xor U11872 (N_11872,N_10755,N_10988);
or U11873 (N_11873,N_10288,N_10429);
nand U11874 (N_11874,N_10077,N_10557);
and U11875 (N_11875,N_10907,N_10051);
and U11876 (N_11876,N_10593,N_10719);
nor U11877 (N_11877,N_10612,N_10879);
or U11878 (N_11878,N_10742,N_10666);
xnor U11879 (N_11879,N_10210,N_10565);
xor U11880 (N_11880,N_10945,N_10664);
nor U11881 (N_11881,N_10142,N_10395);
and U11882 (N_11882,N_10983,N_10475);
nor U11883 (N_11883,N_10644,N_10655);
nand U11884 (N_11884,N_10462,N_10822);
nor U11885 (N_11885,N_10623,N_10815);
xnor U11886 (N_11886,N_10391,N_10224);
or U11887 (N_11887,N_10981,N_10399);
and U11888 (N_11888,N_10386,N_10998);
or U11889 (N_11889,N_10346,N_10202);
and U11890 (N_11890,N_10266,N_10159);
or U11891 (N_11891,N_10925,N_10515);
or U11892 (N_11892,N_10355,N_10263);
nand U11893 (N_11893,N_10672,N_10032);
nor U11894 (N_11894,N_10841,N_10694);
or U11895 (N_11895,N_10668,N_10709);
and U11896 (N_11896,N_10065,N_10487);
nor U11897 (N_11897,N_10640,N_10528);
nor U11898 (N_11898,N_10928,N_10325);
xnor U11899 (N_11899,N_10181,N_10897);
and U11900 (N_11900,N_10529,N_10685);
nor U11901 (N_11901,N_10407,N_10371);
xor U11902 (N_11902,N_10656,N_10755);
nor U11903 (N_11903,N_10323,N_10339);
or U11904 (N_11904,N_10341,N_10314);
or U11905 (N_11905,N_10956,N_10207);
or U11906 (N_11906,N_10997,N_10904);
xnor U11907 (N_11907,N_10865,N_10409);
or U11908 (N_11908,N_10625,N_10804);
and U11909 (N_11909,N_10759,N_10389);
nand U11910 (N_11910,N_10653,N_10195);
xnor U11911 (N_11911,N_10468,N_10771);
and U11912 (N_11912,N_10978,N_10342);
or U11913 (N_11913,N_10326,N_10275);
or U11914 (N_11914,N_10291,N_10200);
nand U11915 (N_11915,N_10099,N_10310);
nand U11916 (N_11916,N_10703,N_10019);
xnor U11917 (N_11917,N_10561,N_10292);
or U11918 (N_11918,N_10582,N_10250);
xor U11919 (N_11919,N_10515,N_10384);
and U11920 (N_11920,N_10318,N_10810);
or U11921 (N_11921,N_10701,N_10381);
xor U11922 (N_11922,N_10426,N_10004);
or U11923 (N_11923,N_10245,N_10909);
or U11924 (N_11924,N_10878,N_10863);
xor U11925 (N_11925,N_10264,N_10458);
xor U11926 (N_11926,N_10602,N_10646);
nand U11927 (N_11927,N_10926,N_10385);
xor U11928 (N_11928,N_10654,N_10936);
nand U11929 (N_11929,N_10380,N_10990);
or U11930 (N_11930,N_10659,N_10932);
nor U11931 (N_11931,N_10549,N_10321);
nand U11932 (N_11932,N_10540,N_10306);
nor U11933 (N_11933,N_10161,N_10971);
nand U11934 (N_11934,N_10961,N_10536);
nor U11935 (N_11935,N_10652,N_10942);
and U11936 (N_11936,N_10415,N_10837);
nand U11937 (N_11937,N_10135,N_10931);
nor U11938 (N_11938,N_10329,N_10786);
nor U11939 (N_11939,N_10364,N_10519);
and U11940 (N_11940,N_10586,N_10153);
nor U11941 (N_11941,N_10682,N_10238);
nand U11942 (N_11942,N_10172,N_10872);
nand U11943 (N_11943,N_10996,N_10013);
xnor U11944 (N_11944,N_10354,N_10578);
and U11945 (N_11945,N_10967,N_10950);
and U11946 (N_11946,N_10159,N_10217);
or U11947 (N_11947,N_10724,N_10734);
or U11948 (N_11948,N_10224,N_10564);
nand U11949 (N_11949,N_10134,N_10600);
nand U11950 (N_11950,N_10374,N_10220);
nand U11951 (N_11951,N_10832,N_10906);
xor U11952 (N_11952,N_10539,N_10753);
nor U11953 (N_11953,N_10477,N_10441);
and U11954 (N_11954,N_10297,N_10738);
nor U11955 (N_11955,N_10728,N_10122);
and U11956 (N_11956,N_10591,N_10973);
xor U11957 (N_11957,N_10533,N_10863);
nor U11958 (N_11958,N_10220,N_10173);
nand U11959 (N_11959,N_10491,N_10796);
or U11960 (N_11960,N_10222,N_10491);
xor U11961 (N_11961,N_10782,N_10225);
nand U11962 (N_11962,N_10611,N_10531);
xor U11963 (N_11963,N_10511,N_10245);
or U11964 (N_11964,N_10596,N_10432);
nor U11965 (N_11965,N_10898,N_10678);
or U11966 (N_11966,N_10049,N_10394);
xnor U11967 (N_11967,N_10984,N_10583);
or U11968 (N_11968,N_10890,N_10981);
or U11969 (N_11969,N_10273,N_10453);
nand U11970 (N_11970,N_10574,N_10506);
nor U11971 (N_11971,N_10051,N_10195);
nand U11972 (N_11972,N_10742,N_10654);
xnor U11973 (N_11973,N_10155,N_10914);
xnor U11974 (N_11974,N_10636,N_10673);
xor U11975 (N_11975,N_10412,N_10919);
or U11976 (N_11976,N_10426,N_10110);
nor U11977 (N_11977,N_10039,N_10858);
nand U11978 (N_11978,N_10207,N_10844);
nor U11979 (N_11979,N_10440,N_10404);
or U11980 (N_11980,N_10829,N_10739);
nand U11981 (N_11981,N_10587,N_10104);
nand U11982 (N_11982,N_10802,N_10723);
nand U11983 (N_11983,N_10119,N_10586);
or U11984 (N_11984,N_10762,N_10679);
and U11985 (N_11985,N_10538,N_10795);
xor U11986 (N_11986,N_10317,N_10603);
xor U11987 (N_11987,N_10504,N_10771);
nand U11988 (N_11988,N_10990,N_10585);
or U11989 (N_11989,N_10791,N_10649);
or U11990 (N_11990,N_10158,N_10194);
and U11991 (N_11991,N_10147,N_10203);
or U11992 (N_11992,N_10826,N_10037);
or U11993 (N_11993,N_10368,N_10438);
xor U11994 (N_11994,N_10409,N_10247);
nand U11995 (N_11995,N_10469,N_10283);
nor U11996 (N_11996,N_10278,N_10732);
xnor U11997 (N_11997,N_10831,N_10352);
or U11998 (N_11998,N_10148,N_10770);
or U11999 (N_11999,N_10307,N_10731);
or U12000 (N_12000,N_11124,N_11739);
and U12001 (N_12001,N_11647,N_11291);
and U12002 (N_12002,N_11755,N_11621);
or U12003 (N_12003,N_11051,N_11322);
nand U12004 (N_12004,N_11513,N_11725);
nor U12005 (N_12005,N_11552,N_11980);
xor U12006 (N_12006,N_11366,N_11344);
nand U12007 (N_12007,N_11446,N_11556);
xor U12008 (N_12008,N_11610,N_11274);
nand U12009 (N_12009,N_11220,N_11460);
nand U12010 (N_12010,N_11862,N_11211);
nor U12011 (N_12011,N_11597,N_11903);
xnor U12012 (N_12012,N_11927,N_11848);
or U12013 (N_12013,N_11428,N_11228);
and U12014 (N_12014,N_11063,N_11112);
xor U12015 (N_12015,N_11675,N_11512);
and U12016 (N_12016,N_11880,N_11649);
nand U12017 (N_12017,N_11243,N_11297);
xor U12018 (N_12018,N_11449,N_11716);
xnor U12019 (N_12019,N_11642,N_11855);
xor U12020 (N_12020,N_11518,N_11204);
nand U12021 (N_12021,N_11607,N_11227);
and U12022 (N_12022,N_11666,N_11008);
nand U12023 (N_12023,N_11863,N_11343);
nor U12024 (N_12024,N_11439,N_11559);
nor U12025 (N_12025,N_11713,N_11194);
xor U12026 (N_12026,N_11507,N_11492);
nor U12027 (N_12027,N_11192,N_11686);
or U12028 (N_12028,N_11009,N_11674);
xor U12029 (N_12029,N_11979,N_11362);
or U12030 (N_12030,N_11892,N_11662);
xnor U12031 (N_12031,N_11265,N_11270);
xnor U12032 (N_12032,N_11949,N_11741);
xnor U12033 (N_12033,N_11942,N_11570);
nand U12034 (N_12034,N_11305,N_11854);
or U12035 (N_12035,N_11829,N_11723);
nand U12036 (N_12036,N_11074,N_11193);
nor U12037 (N_12037,N_11865,N_11718);
xnor U12038 (N_12038,N_11972,N_11622);
or U12039 (N_12039,N_11083,N_11497);
or U12040 (N_12040,N_11263,N_11921);
and U12041 (N_12041,N_11669,N_11434);
xor U12042 (N_12042,N_11920,N_11812);
nand U12043 (N_12043,N_11959,N_11054);
nor U12044 (N_12044,N_11525,N_11625);
and U12045 (N_12045,N_11711,N_11318);
or U12046 (N_12046,N_11715,N_11637);
nor U12047 (N_12047,N_11990,N_11103);
nor U12048 (N_12048,N_11698,N_11350);
xor U12049 (N_12049,N_11751,N_11514);
xnor U12050 (N_12050,N_11731,N_11822);
or U12051 (N_12051,N_11692,N_11538);
and U12052 (N_12052,N_11729,N_11244);
nand U12053 (N_12053,N_11239,N_11445);
nand U12054 (N_12054,N_11911,N_11548);
xnor U12055 (N_12055,N_11567,N_11250);
or U12056 (N_12056,N_11913,N_11383);
nand U12057 (N_12057,N_11037,N_11053);
or U12058 (N_12058,N_11140,N_11502);
nand U12059 (N_12059,N_11437,N_11640);
nor U12060 (N_12060,N_11129,N_11163);
xnor U12061 (N_12061,N_11029,N_11050);
and U12062 (N_12062,N_11233,N_11550);
nand U12063 (N_12063,N_11984,N_11299);
xor U12064 (N_12064,N_11832,N_11749);
or U12065 (N_12065,N_11876,N_11837);
and U12066 (N_12066,N_11255,N_11499);
and U12067 (N_12067,N_11064,N_11365);
nor U12068 (N_12068,N_11402,N_11369);
and U12069 (N_12069,N_11300,N_11438);
and U12070 (N_12070,N_11310,N_11352);
xor U12071 (N_12071,N_11648,N_11150);
xor U12072 (N_12072,N_11826,N_11221);
xnor U12073 (N_12073,N_11728,N_11405);
xor U12074 (N_12074,N_11230,N_11056);
or U12075 (N_12075,N_11278,N_11836);
and U12076 (N_12076,N_11116,N_11934);
xnor U12077 (N_12077,N_11041,N_11632);
xor U12078 (N_12078,N_11209,N_11973);
or U12079 (N_12079,N_11092,N_11391);
nor U12080 (N_12080,N_11823,N_11996);
xnor U12081 (N_12081,N_11667,N_11450);
xnor U12082 (N_12082,N_11453,N_11014);
xor U12083 (N_12083,N_11787,N_11598);
nand U12084 (N_12084,N_11146,N_11722);
and U12085 (N_12085,N_11483,N_11178);
and U12086 (N_12086,N_11771,N_11670);
or U12087 (N_12087,N_11821,N_11432);
nor U12088 (N_12088,N_11135,N_11073);
xnor U12089 (N_12089,N_11997,N_11816);
nand U12090 (N_12090,N_11646,N_11912);
and U12091 (N_12091,N_11440,N_11868);
xnor U12092 (N_12092,N_11746,N_11526);
nand U12093 (N_12093,N_11482,N_11561);
xor U12094 (N_12094,N_11045,N_11824);
nor U12095 (N_12095,N_11010,N_11825);
xor U12096 (N_12096,N_11149,N_11078);
nor U12097 (N_12097,N_11815,N_11409);
nor U12098 (N_12098,N_11510,N_11386);
nor U12099 (N_12099,N_11264,N_11191);
or U12100 (N_12100,N_11448,N_11423);
nand U12101 (N_12101,N_11447,N_11701);
xor U12102 (N_12102,N_11136,N_11605);
nand U12103 (N_12103,N_11871,N_11313);
nand U12104 (N_12104,N_11631,N_11864);
or U12105 (N_12105,N_11267,N_11321);
and U12106 (N_12106,N_11212,N_11102);
nor U12107 (N_12107,N_11852,N_11748);
xnor U12108 (N_12108,N_11909,N_11775);
or U12109 (N_12109,N_11006,N_11473);
and U12110 (N_12110,N_11065,N_11072);
and U12111 (N_12111,N_11677,N_11375);
nand U12112 (N_12112,N_11390,N_11442);
nor U12113 (N_12113,N_11800,N_11047);
nor U12114 (N_12114,N_11364,N_11097);
xnor U12115 (N_12115,N_11043,N_11897);
xnor U12116 (N_12116,N_11882,N_11184);
nand U12117 (N_12117,N_11120,N_11841);
or U12118 (N_12118,N_11324,N_11218);
and U12119 (N_12119,N_11700,N_11060);
nand U12120 (N_12120,N_11470,N_11726);
and U12121 (N_12121,N_11315,N_11123);
or U12122 (N_12122,N_11738,N_11340);
nand U12123 (N_12123,N_11298,N_11081);
nor U12124 (N_12124,N_11842,N_11472);
xnor U12125 (N_12125,N_11501,N_11110);
nor U12126 (N_12126,N_11888,N_11544);
nand U12127 (N_12127,N_11576,N_11828);
xnor U12128 (N_12128,N_11680,N_11554);
xor U12129 (N_12129,N_11515,N_11049);
nand U12130 (N_12130,N_11186,N_11183);
or U12131 (N_12131,N_11735,N_11287);
nand U12132 (N_12132,N_11813,N_11196);
and U12133 (N_12133,N_11777,N_11090);
nor U12134 (N_12134,N_11595,N_11866);
and U12135 (N_12135,N_11020,N_11965);
nand U12136 (N_12136,N_11633,N_11190);
nor U12137 (N_12137,N_11033,N_11985);
and U12138 (N_12138,N_11207,N_11469);
xor U12139 (N_12139,N_11847,N_11144);
and U12140 (N_12140,N_11283,N_11705);
nand U12141 (N_12141,N_11969,N_11917);
nor U12142 (N_12142,N_11257,N_11275);
or U12143 (N_12143,N_11484,N_11603);
or U12144 (N_12144,N_11232,N_11883);
or U12145 (N_12145,N_11736,N_11519);
xor U12146 (N_12146,N_11948,N_11328);
or U12147 (N_12147,N_11983,N_11306);
or U12148 (N_12148,N_11334,N_11893);
xnor U12149 (N_12149,N_11346,N_11976);
xor U12150 (N_12150,N_11148,N_11634);
or U12151 (N_12151,N_11914,N_11947);
and U12152 (N_12152,N_11377,N_11466);
and U12153 (N_12153,N_11704,N_11480);
and U12154 (N_12154,N_11485,N_11793);
nor U12155 (N_12155,N_11012,N_11487);
nand U12156 (N_12156,N_11034,N_11489);
nand U12157 (N_12157,N_11319,N_11424);
or U12158 (N_12158,N_11796,N_11960);
and U12159 (N_12159,N_11881,N_11908);
or U12160 (N_12160,N_11467,N_11496);
and U12161 (N_12161,N_11215,N_11898);
nand U12162 (N_12162,N_11774,N_11651);
nor U12163 (N_12163,N_11989,N_11293);
nand U12164 (N_12164,N_11696,N_11400);
xnor U12165 (N_12165,N_11582,N_11879);
xnor U12166 (N_12166,N_11999,N_11189);
nor U12167 (N_12167,N_11853,N_11187);
xnor U12168 (N_12168,N_11312,N_11106);
and U12169 (N_12169,N_11229,N_11644);
nor U12170 (N_12170,N_11660,N_11134);
or U12171 (N_12171,N_11180,N_11523);
and U12172 (N_12172,N_11981,N_11062);
xnor U12173 (N_12173,N_11536,N_11994);
nor U12174 (N_12174,N_11630,N_11753);
xnor U12175 (N_12175,N_11403,N_11331);
or U12176 (N_12176,N_11543,N_11727);
nand U12177 (N_12177,N_11673,N_11130);
xor U12178 (N_12178,N_11262,N_11923);
nand U12179 (N_12179,N_11356,N_11046);
or U12180 (N_12180,N_11918,N_11431);
nand U12181 (N_12181,N_11742,N_11583);
nor U12182 (N_12182,N_11370,N_11203);
or U12183 (N_12183,N_11117,N_11922);
nand U12184 (N_12184,N_11546,N_11814);
nand U12185 (N_12185,N_11943,N_11664);
and U12186 (N_12186,N_11145,N_11977);
nor U12187 (N_12187,N_11689,N_11153);
or U12188 (N_12188,N_11584,N_11127);
and U12189 (N_12189,N_11950,N_11810);
nor U12190 (N_12190,N_11587,N_11817);
nand U12191 (N_12191,N_11613,N_11846);
or U12192 (N_12192,N_11011,N_11137);
or U12193 (N_12193,N_11174,N_11463);
and U12194 (N_12194,N_11441,N_11216);
nand U12195 (N_12195,N_11872,N_11374);
nor U12196 (N_12196,N_11131,N_11084);
nand U12197 (N_12197,N_11296,N_11007);
nor U12198 (N_12198,N_11833,N_11044);
and U12199 (N_12199,N_11733,N_11776);
nor U12200 (N_12200,N_11158,N_11167);
nand U12201 (N_12201,N_11650,N_11363);
nand U12202 (N_12202,N_11085,N_11075);
xnor U12203 (N_12203,N_11429,N_11253);
and U12204 (N_12204,N_11724,N_11294);
or U12205 (N_12205,N_11773,N_11258);
or U12206 (N_12206,N_11557,N_11966);
or U12207 (N_12207,N_11867,N_11925);
nand U12208 (N_12208,N_11618,N_11122);
or U12209 (N_12209,N_11798,N_11138);
or U12210 (N_12210,N_11845,N_11500);
and U12211 (N_12211,N_11659,N_11024);
or U12212 (N_12212,N_11332,N_11185);
nor U12213 (N_12213,N_11381,N_11268);
and U12214 (N_12214,N_11353,N_11978);
xor U12215 (N_12215,N_11671,N_11308);
or U12216 (N_12216,N_11104,N_11427);
nand U12217 (N_12217,N_11417,N_11993);
or U12218 (N_12218,N_11048,N_11139);
nand U12219 (N_12219,N_11916,N_11589);
or U12220 (N_12220,N_11170,N_11354);
xor U12221 (N_12221,N_11577,N_11697);
nand U12222 (N_12222,N_11961,N_11132);
or U12223 (N_12223,N_11379,N_11367);
nor U12224 (N_12224,N_11086,N_11844);
xnor U12225 (N_12225,N_11133,N_11182);
and U12226 (N_12226,N_11373,N_11719);
nor U12227 (N_12227,N_11802,N_11387);
and U12228 (N_12228,N_11799,N_11330);
xor U12229 (N_12229,N_11763,N_11069);
and U12230 (N_12230,N_11068,N_11404);
nor U12231 (N_12231,N_11804,N_11752);
xor U12232 (N_12232,N_11475,N_11658);
or U12233 (N_12233,N_11778,N_11080);
nand U12234 (N_12234,N_11341,N_11693);
xor U12235 (N_12235,N_11702,N_11685);
and U12236 (N_12236,N_11504,N_11626);
and U12237 (N_12237,N_11540,N_11309);
nand U12238 (N_12238,N_11682,N_11172);
nand U12239 (N_12239,N_11433,N_11099);
or U12240 (N_12240,N_11498,N_11225);
xor U12241 (N_12241,N_11477,N_11430);
and U12242 (N_12242,N_11358,N_11160);
or U12243 (N_12243,N_11936,N_11592);
and U12244 (N_12244,N_11780,N_11986);
xnor U12245 (N_12245,N_11506,N_11668);
nand U12246 (N_12246,N_11851,N_11858);
and U12247 (N_12247,N_11517,N_11179);
nand U12248 (N_12248,N_11290,N_11089);
nor U12249 (N_12249,N_11412,N_11039);
nand U12250 (N_12250,N_11581,N_11590);
or U12251 (N_12251,N_11260,N_11884);
nor U12252 (N_12252,N_11326,N_11143);
nor U12253 (N_12253,N_11171,N_11935);
and U12254 (N_12254,N_11602,N_11076);
xor U12255 (N_12255,N_11026,N_11820);
or U12256 (N_12256,N_11141,N_11964);
and U12257 (N_12257,N_11388,N_11574);
xnor U12258 (N_12258,N_11055,N_11380);
nor U12259 (N_12259,N_11838,N_11712);
xnor U12260 (N_12260,N_11114,N_11995);
xnor U12261 (N_12261,N_11198,N_11806);
nand U12262 (N_12262,N_11563,N_11407);
xnor U12263 (N_12263,N_11952,N_11962);
or U12264 (N_12264,N_11443,N_11242);
or U12265 (N_12265,N_11474,N_11119);
nor U12266 (N_12266,N_11571,N_11240);
nor U12267 (N_12267,N_11740,N_11645);
nand U12268 (N_12268,N_11545,N_11732);
nand U12269 (N_12269,N_11461,N_11077);
or U12270 (N_12270,N_11121,N_11615);
and U12271 (N_12271,N_11394,N_11772);
nor U12272 (N_12272,N_11468,N_11398);
xor U12273 (N_12273,N_11537,N_11285);
nand U12274 (N_12274,N_11079,N_11125);
or U12275 (N_12275,N_11929,N_11451);
nor U12276 (N_12276,N_11527,N_11347);
or U12277 (N_12277,N_11524,N_11811);
xnor U12278 (N_12278,N_11565,N_11834);
and U12279 (N_12279,N_11560,N_11491);
nand U12280 (N_12280,N_11486,N_11805);
nor U12281 (N_12281,N_11765,N_11195);
xnor U12282 (N_12282,N_11788,N_11154);
or U12283 (N_12283,N_11159,N_11691);
nor U12284 (N_12284,N_11038,N_11493);
and U12285 (N_12285,N_11945,N_11663);
or U12286 (N_12286,N_11809,N_11606);
or U12287 (N_12287,N_11717,N_11249);
xnor U12288 (N_12288,N_11569,N_11345);
nor U12289 (N_12289,N_11769,N_11594);
and U12290 (N_12290,N_11338,N_11385);
nand U12291 (N_12291,N_11902,N_11494);
and U12292 (N_12292,N_11316,N_11396);
nand U12293 (N_12293,N_11311,N_11416);
xnor U12294 (N_12294,N_11176,N_11455);
and U12295 (N_12295,N_11588,N_11408);
or U12296 (N_12296,N_11454,N_11052);
and U12297 (N_12297,N_11436,N_11789);
and U12298 (N_12298,N_11707,N_11444);
xnor U12299 (N_12299,N_11004,N_11988);
xor U12300 (N_12300,N_11357,N_11600);
nand U12301 (N_12301,N_11992,N_11505);
nor U12302 (N_12302,N_11295,N_11568);
and U12303 (N_12303,N_11015,N_11681);
nor U12304 (N_12304,N_11259,N_11720);
and U12305 (N_12305,N_11213,N_11784);
and U12306 (N_12306,N_11181,N_11688);
nor U12307 (N_12307,N_11002,N_11155);
or U12308 (N_12308,N_11878,N_11635);
xnor U12309 (N_12309,N_11877,N_11779);
xor U12310 (N_12310,N_11827,N_11653);
and U12311 (N_12311,N_11040,N_11998);
and U12312 (N_12312,N_11478,N_11614);
or U12313 (N_12313,N_11819,N_11027);
nor U12314 (N_12314,N_11302,N_11803);
or U12315 (N_12315,N_11957,N_11111);
nand U12316 (N_12316,N_11933,N_11458);
nor U12317 (N_12317,N_11395,N_11005);
nor U12318 (N_12318,N_11757,N_11529);
nor U12319 (N_12319,N_11756,N_11292);
and U12320 (N_12320,N_11906,N_11406);
or U12321 (N_12321,N_11591,N_11797);
or U12322 (N_12322,N_11737,N_11217);
or U12323 (N_12323,N_11869,N_11573);
or U12324 (N_12324,N_11284,N_11231);
and U12325 (N_12325,N_11608,N_11282);
nor U12326 (N_12326,N_11036,N_11564);
nand U12327 (N_12327,N_11169,N_11508);
nor U12328 (N_12328,N_11730,N_11251);
or U12329 (N_12329,N_11128,N_11638);
and U12330 (N_12330,N_11082,N_11162);
or U12331 (N_12331,N_11744,N_11109);
xor U12332 (N_12332,N_11413,N_11580);
nand U12333 (N_12333,N_11747,N_11401);
nand U12334 (N_12334,N_11035,N_11206);
nor U12335 (N_12335,N_11899,N_11094);
or U12336 (N_12336,N_11360,N_11967);
or U12337 (N_12337,N_11910,N_11987);
and U12338 (N_12338,N_11223,N_11585);
xnor U12339 (N_12339,N_11411,N_11210);
xor U12340 (N_12340,N_11767,N_11522);
and U12341 (N_12341,N_11839,N_11017);
nand U12342 (N_12342,N_11954,N_11320);
xnor U12343 (N_12343,N_11889,N_11279);
or U12344 (N_12344,N_11021,N_11703);
and U12345 (N_12345,N_11951,N_11013);
or U12346 (N_12346,N_11059,N_11425);
nor U12347 (N_12347,N_11261,N_11539);
nand U12348 (N_12348,N_11932,N_11435);
and U12349 (N_12349,N_11547,N_11963);
or U12350 (N_12350,N_11070,N_11678);
xor U12351 (N_12351,N_11553,N_11907);
and U12352 (N_12352,N_11471,N_11792);
nor U12353 (N_12353,N_11241,N_11870);
and U12354 (N_12354,N_11214,N_11672);
nor U12355 (N_12355,N_11654,N_11378);
nand U12356 (N_12356,N_11327,N_11107);
xnor U12357 (N_12357,N_11721,N_11875);
xnor U12358 (N_12358,N_11157,N_11426);
or U12359 (N_12359,N_11419,N_11481);
nor U12360 (N_12360,N_11894,N_11801);
xnor U12361 (N_12361,N_11071,N_11452);
nand U12362 (N_12362,N_11246,N_11224);
nand U12363 (N_12363,N_11323,N_11376);
xor U12364 (N_12364,N_11115,N_11530);
nand U12365 (N_12365,N_11937,N_11277);
nor U12366 (N_12366,N_11641,N_11028);
and U12367 (N_12367,N_11333,N_11915);
or U12368 (N_12368,N_11359,N_11679);
nand U12369 (N_12369,N_11782,N_11843);
nor U12370 (N_12370,N_11890,N_11745);
xnor U12371 (N_12371,N_11301,N_11549);
nand U12372 (N_12372,N_11096,N_11562);
nor U12373 (N_12373,N_11555,N_11859);
nand U12374 (N_12374,N_11687,N_11465);
and U12375 (N_12375,N_11256,N_11337);
nor U12376 (N_12376,N_11355,N_11339);
xor U12377 (N_12377,N_11205,N_11349);
or U12378 (N_12378,N_11612,N_11414);
nand U12379 (N_12379,N_11891,N_11930);
nand U12380 (N_12380,N_11904,N_11532);
and U12381 (N_12381,N_11415,N_11629);
nor U12382 (N_12382,N_11520,N_11286);
or U12383 (N_12383,N_11156,N_11113);
nand U12384 (N_12384,N_11105,N_11147);
or U12385 (N_12385,N_11768,N_11652);
nor U12386 (N_12386,N_11503,N_11410);
and U12387 (N_12387,N_11535,N_11760);
and U12388 (N_12388,N_11329,N_11371);
xnor U12389 (N_12389,N_11860,N_11939);
and U12390 (N_12390,N_11273,N_11617);
or U12391 (N_12391,N_11226,N_11289);
xor U12392 (N_12392,N_11857,N_11770);
nand U12393 (N_12393,N_11420,N_11269);
xnor U12394 (N_12394,N_11032,N_11558);
xor U12395 (N_12395,N_11766,N_11236);
or U12396 (N_12396,N_11057,N_11968);
xor U12397 (N_12397,N_11247,N_11786);
nor U12398 (N_12398,N_11151,N_11066);
nor U12399 (N_12399,N_11095,N_11271);
or U12400 (N_12400,N_11542,N_11975);
or U12401 (N_12401,N_11188,N_11807);
and U12402 (N_12402,N_11831,N_11946);
xnor U12403 (N_12403,N_11656,N_11609);
xor U12404 (N_12404,N_11101,N_11579);
or U12405 (N_12405,N_11885,N_11022);
or U12406 (N_12406,N_11165,N_11761);
nand U12407 (N_12407,N_11616,N_11657);
xnor U12408 (N_12408,N_11361,N_11706);
xnor U12409 (N_12409,N_11676,N_11699);
and U12410 (N_12410,N_11222,N_11238);
nand U12411 (N_12411,N_11905,N_11288);
nor U12412 (N_12412,N_11785,N_11762);
and U12413 (N_12413,N_11783,N_11516);
xnor U12414 (N_12414,N_11457,N_11087);
and U12415 (N_12415,N_11694,N_11245);
xor U12416 (N_12416,N_11991,N_11709);
nand U12417 (N_12417,N_11901,N_11197);
nor U12418 (N_12418,N_11368,N_11208);
and U12419 (N_12419,N_11000,N_11808);
xor U12420 (N_12420,N_11714,N_11509);
and U12421 (N_12421,N_11202,N_11665);
xnor U12422 (N_12422,N_11953,N_11091);
xnor U12423 (N_12423,N_11304,N_11382);
nor U12424 (N_12424,N_11025,N_11058);
xor U12425 (N_12425,N_11325,N_11276);
or U12426 (N_12426,N_11931,N_11955);
or U12427 (N_12427,N_11272,N_11620);
or U12428 (N_12428,N_11303,N_11623);
or U12429 (N_12429,N_11490,N_11849);
nand U12430 (N_12430,N_11734,N_11593);
nand U12431 (N_12431,N_11164,N_11759);
and U12432 (N_12432,N_11200,N_11201);
nand U12433 (N_12433,N_11126,N_11578);
xnor U12434 (N_12434,N_11750,N_11886);
nand U12435 (N_12435,N_11791,N_11142);
and U12436 (N_12436,N_11393,N_11627);
nor U12437 (N_12437,N_11690,N_11237);
or U12438 (N_12438,N_11840,N_11521);
nand U12439 (N_12439,N_11684,N_11397);
nor U12440 (N_12440,N_11944,N_11611);
nand U12441 (N_12441,N_11511,N_11575);
or U12442 (N_12442,N_11604,N_11314);
nor U12443 (N_12443,N_11234,N_11896);
nand U12444 (N_12444,N_11266,N_11166);
and U12445 (N_12445,N_11177,N_11235);
nor U12446 (N_12446,N_11422,N_11683);
nand U12447 (N_12447,N_11456,N_11018);
and U12448 (N_12448,N_11372,N_11531);
and U12449 (N_12449,N_11956,N_11118);
nor U12450 (N_12450,N_11958,N_11941);
or U12451 (N_12451,N_11534,N_11317);
nand U12452 (N_12452,N_11342,N_11900);
nor U12453 (N_12453,N_11850,N_11152);
nand U12454 (N_12454,N_11795,N_11919);
nor U12455 (N_12455,N_11459,N_11175);
xnor U12456 (N_12456,N_11030,N_11794);
xnor U12457 (N_12457,N_11108,N_11348);
and U12458 (N_12458,N_11533,N_11541);
and U12459 (N_12459,N_11219,N_11572);
nor U12460 (N_12460,N_11861,N_11248);
xnor U12461 (N_12461,N_11088,N_11399);
and U12462 (N_12462,N_11061,N_11974);
nand U12463 (N_12463,N_11016,N_11856);
nor U12464 (N_12464,N_11421,N_11488);
nand U12465 (N_12465,N_11924,N_11601);
nand U12466 (N_12466,N_11479,N_11926);
and U12467 (N_12467,N_11093,N_11464);
nor U12468 (N_12468,N_11661,N_11495);
xnor U12469 (N_12469,N_11351,N_11695);
nor U12470 (N_12470,N_11835,N_11336);
and U12471 (N_12471,N_11874,N_11281);
or U12472 (N_12472,N_11003,N_11940);
nand U12473 (N_12473,N_11476,N_11280);
nand U12474 (N_12474,N_11001,N_11528);
xnor U12475 (N_12475,N_11818,N_11586);
or U12476 (N_12476,N_11982,N_11970);
nand U12477 (N_12477,N_11710,N_11636);
and U12478 (N_12478,N_11418,N_11971);
and U12479 (N_12479,N_11655,N_11599);
nor U12480 (N_12480,N_11873,N_11067);
nor U12481 (N_12481,N_11628,N_11335);
and U12482 (N_12482,N_11830,N_11252);
and U12483 (N_12483,N_11643,N_11384);
nand U12484 (N_12484,N_11254,N_11639);
xnor U12485 (N_12485,N_11392,N_11938);
nor U12486 (N_12486,N_11019,N_11566);
or U12487 (N_12487,N_11462,N_11596);
nand U12488 (N_12488,N_11743,N_11764);
and U12489 (N_12489,N_11624,N_11199);
or U12490 (N_12490,N_11098,N_11389);
xnor U12491 (N_12491,N_11708,N_11307);
and U12492 (N_12492,N_11790,N_11042);
and U12493 (N_12493,N_11619,N_11758);
and U12494 (N_12494,N_11173,N_11887);
xnor U12495 (N_12495,N_11023,N_11895);
nor U12496 (N_12496,N_11551,N_11754);
nor U12497 (N_12497,N_11928,N_11100);
nor U12498 (N_12498,N_11161,N_11031);
or U12499 (N_12499,N_11781,N_11168);
nor U12500 (N_12500,N_11353,N_11661);
nand U12501 (N_12501,N_11913,N_11237);
nor U12502 (N_12502,N_11514,N_11095);
nor U12503 (N_12503,N_11127,N_11177);
nor U12504 (N_12504,N_11180,N_11371);
or U12505 (N_12505,N_11210,N_11201);
or U12506 (N_12506,N_11308,N_11306);
nand U12507 (N_12507,N_11099,N_11751);
xnor U12508 (N_12508,N_11683,N_11975);
nand U12509 (N_12509,N_11932,N_11061);
nand U12510 (N_12510,N_11869,N_11764);
or U12511 (N_12511,N_11281,N_11453);
and U12512 (N_12512,N_11359,N_11741);
nor U12513 (N_12513,N_11207,N_11130);
nand U12514 (N_12514,N_11084,N_11831);
nor U12515 (N_12515,N_11081,N_11838);
and U12516 (N_12516,N_11155,N_11678);
and U12517 (N_12517,N_11156,N_11042);
or U12518 (N_12518,N_11546,N_11705);
and U12519 (N_12519,N_11505,N_11121);
nor U12520 (N_12520,N_11211,N_11681);
nand U12521 (N_12521,N_11221,N_11369);
and U12522 (N_12522,N_11664,N_11025);
nand U12523 (N_12523,N_11716,N_11615);
xor U12524 (N_12524,N_11382,N_11923);
nor U12525 (N_12525,N_11620,N_11170);
nor U12526 (N_12526,N_11950,N_11235);
nor U12527 (N_12527,N_11490,N_11881);
nand U12528 (N_12528,N_11762,N_11218);
or U12529 (N_12529,N_11522,N_11078);
nand U12530 (N_12530,N_11385,N_11690);
and U12531 (N_12531,N_11163,N_11194);
nand U12532 (N_12532,N_11197,N_11443);
xnor U12533 (N_12533,N_11168,N_11606);
nand U12534 (N_12534,N_11657,N_11558);
xor U12535 (N_12535,N_11556,N_11107);
and U12536 (N_12536,N_11786,N_11997);
nand U12537 (N_12537,N_11046,N_11483);
nand U12538 (N_12538,N_11560,N_11075);
nor U12539 (N_12539,N_11789,N_11125);
nand U12540 (N_12540,N_11690,N_11948);
nor U12541 (N_12541,N_11727,N_11968);
and U12542 (N_12542,N_11336,N_11885);
or U12543 (N_12543,N_11701,N_11319);
nand U12544 (N_12544,N_11285,N_11199);
nand U12545 (N_12545,N_11821,N_11920);
xnor U12546 (N_12546,N_11405,N_11018);
nor U12547 (N_12547,N_11153,N_11546);
nand U12548 (N_12548,N_11387,N_11759);
nand U12549 (N_12549,N_11220,N_11958);
nor U12550 (N_12550,N_11170,N_11880);
or U12551 (N_12551,N_11691,N_11706);
nor U12552 (N_12552,N_11081,N_11053);
and U12553 (N_12553,N_11178,N_11531);
xnor U12554 (N_12554,N_11460,N_11964);
xnor U12555 (N_12555,N_11341,N_11785);
nor U12556 (N_12556,N_11553,N_11555);
and U12557 (N_12557,N_11659,N_11390);
xnor U12558 (N_12558,N_11565,N_11460);
nand U12559 (N_12559,N_11364,N_11904);
and U12560 (N_12560,N_11839,N_11840);
nor U12561 (N_12561,N_11986,N_11038);
or U12562 (N_12562,N_11520,N_11431);
xor U12563 (N_12563,N_11191,N_11042);
and U12564 (N_12564,N_11758,N_11199);
or U12565 (N_12565,N_11630,N_11393);
nand U12566 (N_12566,N_11998,N_11388);
nor U12567 (N_12567,N_11710,N_11618);
or U12568 (N_12568,N_11882,N_11586);
nor U12569 (N_12569,N_11134,N_11128);
and U12570 (N_12570,N_11455,N_11548);
nor U12571 (N_12571,N_11292,N_11796);
xnor U12572 (N_12572,N_11637,N_11433);
xor U12573 (N_12573,N_11159,N_11363);
and U12574 (N_12574,N_11397,N_11728);
nand U12575 (N_12575,N_11128,N_11448);
or U12576 (N_12576,N_11006,N_11860);
nor U12577 (N_12577,N_11144,N_11602);
nand U12578 (N_12578,N_11909,N_11673);
xnor U12579 (N_12579,N_11077,N_11945);
or U12580 (N_12580,N_11714,N_11325);
and U12581 (N_12581,N_11409,N_11217);
xnor U12582 (N_12582,N_11358,N_11953);
or U12583 (N_12583,N_11221,N_11057);
nor U12584 (N_12584,N_11562,N_11619);
or U12585 (N_12585,N_11286,N_11213);
and U12586 (N_12586,N_11367,N_11710);
xor U12587 (N_12587,N_11559,N_11415);
nand U12588 (N_12588,N_11392,N_11141);
xnor U12589 (N_12589,N_11675,N_11585);
and U12590 (N_12590,N_11165,N_11920);
and U12591 (N_12591,N_11515,N_11604);
nor U12592 (N_12592,N_11042,N_11086);
xnor U12593 (N_12593,N_11923,N_11305);
nand U12594 (N_12594,N_11006,N_11110);
or U12595 (N_12595,N_11866,N_11771);
nor U12596 (N_12596,N_11188,N_11592);
or U12597 (N_12597,N_11190,N_11157);
or U12598 (N_12598,N_11048,N_11363);
nor U12599 (N_12599,N_11530,N_11297);
xnor U12600 (N_12600,N_11723,N_11967);
nor U12601 (N_12601,N_11188,N_11324);
nand U12602 (N_12602,N_11756,N_11091);
nand U12603 (N_12603,N_11332,N_11482);
and U12604 (N_12604,N_11074,N_11458);
xor U12605 (N_12605,N_11029,N_11669);
xor U12606 (N_12606,N_11193,N_11150);
xnor U12607 (N_12607,N_11409,N_11856);
xnor U12608 (N_12608,N_11964,N_11642);
xor U12609 (N_12609,N_11149,N_11526);
nor U12610 (N_12610,N_11363,N_11111);
or U12611 (N_12611,N_11465,N_11056);
and U12612 (N_12612,N_11633,N_11165);
and U12613 (N_12613,N_11732,N_11407);
nor U12614 (N_12614,N_11778,N_11372);
or U12615 (N_12615,N_11110,N_11796);
or U12616 (N_12616,N_11847,N_11869);
nor U12617 (N_12617,N_11083,N_11035);
nand U12618 (N_12618,N_11872,N_11844);
or U12619 (N_12619,N_11512,N_11053);
or U12620 (N_12620,N_11180,N_11893);
nor U12621 (N_12621,N_11002,N_11332);
xnor U12622 (N_12622,N_11572,N_11045);
and U12623 (N_12623,N_11566,N_11877);
nand U12624 (N_12624,N_11170,N_11602);
or U12625 (N_12625,N_11511,N_11033);
xnor U12626 (N_12626,N_11129,N_11729);
or U12627 (N_12627,N_11763,N_11110);
and U12628 (N_12628,N_11456,N_11402);
and U12629 (N_12629,N_11412,N_11092);
nor U12630 (N_12630,N_11271,N_11757);
xnor U12631 (N_12631,N_11859,N_11964);
and U12632 (N_12632,N_11638,N_11901);
nand U12633 (N_12633,N_11995,N_11729);
nor U12634 (N_12634,N_11498,N_11239);
nand U12635 (N_12635,N_11574,N_11591);
nor U12636 (N_12636,N_11566,N_11560);
and U12637 (N_12637,N_11939,N_11851);
xor U12638 (N_12638,N_11943,N_11756);
nand U12639 (N_12639,N_11162,N_11973);
nand U12640 (N_12640,N_11951,N_11219);
xor U12641 (N_12641,N_11168,N_11844);
or U12642 (N_12642,N_11869,N_11777);
nand U12643 (N_12643,N_11611,N_11683);
xor U12644 (N_12644,N_11809,N_11684);
nand U12645 (N_12645,N_11584,N_11189);
xor U12646 (N_12646,N_11281,N_11988);
nand U12647 (N_12647,N_11729,N_11571);
nand U12648 (N_12648,N_11168,N_11359);
xnor U12649 (N_12649,N_11441,N_11693);
or U12650 (N_12650,N_11489,N_11923);
or U12651 (N_12651,N_11760,N_11914);
or U12652 (N_12652,N_11250,N_11659);
and U12653 (N_12653,N_11850,N_11719);
xor U12654 (N_12654,N_11022,N_11238);
nor U12655 (N_12655,N_11635,N_11086);
or U12656 (N_12656,N_11973,N_11149);
nand U12657 (N_12657,N_11728,N_11719);
nand U12658 (N_12658,N_11359,N_11630);
nand U12659 (N_12659,N_11558,N_11612);
xnor U12660 (N_12660,N_11013,N_11056);
and U12661 (N_12661,N_11190,N_11689);
nand U12662 (N_12662,N_11016,N_11432);
or U12663 (N_12663,N_11337,N_11563);
and U12664 (N_12664,N_11958,N_11120);
or U12665 (N_12665,N_11304,N_11465);
nor U12666 (N_12666,N_11803,N_11650);
nand U12667 (N_12667,N_11132,N_11455);
nor U12668 (N_12668,N_11078,N_11331);
or U12669 (N_12669,N_11540,N_11114);
nor U12670 (N_12670,N_11046,N_11636);
and U12671 (N_12671,N_11553,N_11921);
and U12672 (N_12672,N_11154,N_11362);
and U12673 (N_12673,N_11834,N_11348);
and U12674 (N_12674,N_11521,N_11388);
and U12675 (N_12675,N_11276,N_11936);
or U12676 (N_12676,N_11360,N_11100);
xnor U12677 (N_12677,N_11900,N_11527);
xnor U12678 (N_12678,N_11721,N_11400);
and U12679 (N_12679,N_11288,N_11962);
nor U12680 (N_12680,N_11796,N_11413);
and U12681 (N_12681,N_11773,N_11165);
xor U12682 (N_12682,N_11666,N_11442);
nor U12683 (N_12683,N_11161,N_11171);
or U12684 (N_12684,N_11731,N_11668);
and U12685 (N_12685,N_11048,N_11217);
nor U12686 (N_12686,N_11755,N_11929);
nor U12687 (N_12687,N_11147,N_11724);
xnor U12688 (N_12688,N_11411,N_11256);
nor U12689 (N_12689,N_11052,N_11333);
xor U12690 (N_12690,N_11455,N_11805);
and U12691 (N_12691,N_11250,N_11157);
nor U12692 (N_12692,N_11850,N_11427);
or U12693 (N_12693,N_11893,N_11010);
and U12694 (N_12694,N_11780,N_11103);
and U12695 (N_12695,N_11113,N_11103);
xor U12696 (N_12696,N_11241,N_11940);
or U12697 (N_12697,N_11017,N_11752);
or U12698 (N_12698,N_11687,N_11566);
nor U12699 (N_12699,N_11076,N_11682);
or U12700 (N_12700,N_11835,N_11413);
nand U12701 (N_12701,N_11369,N_11932);
nor U12702 (N_12702,N_11581,N_11626);
nor U12703 (N_12703,N_11522,N_11981);
nor U12704 (N_12704,N_11574,N_11600);
nand U12705 (N_12705,N_11788,N_11163);
nor U12706 (N_12706,N_11561,N_11325);
and U12707 (N_12707,N_11896,N_11341);
or U12708 (N_12708,N_11768,N_11395);
nor U12709 (N_12709,N_11395,N_11596);
or U12710 (N_12710,N_11479,N_11108);
nand U12711 (N_12711,N_11891,N_11908);
and U12712 (N_12712,N_11271,N_11225);
nand U12713 (N_12713,N_11764,N_11971);
nand U12714 (N_12714,N_11575,N_11605);
nand U12715 (N_12715,N_11803,N_11489);
xor U12716 (N_12716,N_11776,N_11518);
xnor U12717 (N_12717,N_11845,N_11083);
or U12718 (N_12718,N_11817,N_11879);
nand U12719 (N_12719,N_11137,N_11445);
nand U12720 (N_12720,N_11185,N_11843);
nor U12721 (N_12721,N_11672,N_11527);
and U12722 (N_12722,N_11666,N_11448);
and U12723 (N_12723,N_11964,N_11085);
or U12724 (N_12724,N_11125,N_11732);
xnor U12725 (N_12725,N_11998,N_11080);
xor U12726 (N_12726,N_11735,N_11654);
and U12727 (N_12727,N_11541,N_11202);
or U12728 (N_12728,N_11613,N_11593);
xor U12729 (N_12729,N_11022,N_11013);
and U12730 (N_12730,N_11151,N_11661);
nand U12731 (N_12731,N_11854,N_11000);
or U12732 (N_12732,N_11925,N_11015);
xnor U12733 (N_12733,N_11038,N_11443);
and U12734 (N_12734,N_11689,N_11422);
and U12735 (N_12735,N_11386,N_11364);
or U12736 (N_12736,N_11689,N_11433);
and U12737 (N_12737,N_11627,N_11773);
or U12738 (N_12738,N_11177,N_11173);
xnor U12739 (N_12739,N_11097,N_11206);
or U12740 (N_12740,N_11194,N_11362);
or U12741 (N_12741,N_11796,N_11453);
nor U12742 (N_12742,N_11448,N_11578);
nand U12743 (N_12743,N_11229,N_11151);
nor U12744 (N_12744,N_11035,N_11174);
nand U12745 (N_12745,N_11227,N_11078);
nor U12746 (N_12746,N_11723,N_11860);
nand U12747 (N_12747,N_11297,N_11119);
nand U12748 (N_12748,N_11758,N_11544);
nand U12749 (N_12749,N_11477,N_11062);
or U12750 (N_12750,N_11192,N_11799);
or U12751 (N_12751,N_11962,N_11453);
nor U12752 (N_12752,N_11911,N_11814);
nand U12753 (N_12753,N_11717,N_11901);
or U12754 (N_12754,N_11056,N_11753);
and U12755 (N_12755,N_11917,N_11506);
nand U12756 (N_12756,N_11619,N_11474);
nor U12757 (N_12757,N_11846,N_11540);
and U12758 (N_12758,N_11768,N_11247);
xor U12759 (N_12759,N_11025,N_11842);
or U12760 (N_12760,N_11924,N_11739);
xor U12761 (N_12761,N_11811,N_11928);
xor U12762 (N_12762,N_11654,N_11486);
or U12763 (N_12763,N_11865,N_11021);
and U12764 (N_12764,N_11025,N_11885);
xnor U12765 (N_12765,N_11780,N_11551);
and U12766 (N_12766,N_11451,N_11395);
nand U12767 (N_12767,N_11581,N_11031);
xnor U12768 (N_12768,N_11768,N_11417);
nand U12769 (N_12769,N_11912,N_11957);
nand U12770 (N_12770,N_11491,N_11029);
and U12771 (N_12771,N_11343,N_11920);
and U12772 (N_12772,N_11584,N_11333);
nor U12773 (N_12773,N_11440,N_11595);
xnor U12774 (N_12774,N_11668,N_11404);
nor U12775 (N_12775,N_11877,N_11424);
nand U12776 (N_12776,N_11183,N_11283);
and U12777 (N_12777,N_11756,N_11610);
and U12778 (N_12778,N_11369,N_11175);
nor U12779 (N_12779,N_11504,N_11992);
or U12780 (N_12780,N_11672,N_11739);
nand U12781 (N_12781,N_11760,N_11932);
or U12782 (N_12782,N_11192,N_11685);
nand U12783 (N_12783,N_11198,N_11919);
nand U12784 (N_12784,N_11775,N_11980);
nand U12785 (N_12785,N_11688,N_11793);
xor U12786 (N_12786,N_11627,N_11475);
nor U12787 (N_12787,N_11793,N_11341);
or U12788 (N_12788,N_11882,N_11363);
nor U12789 (N_12789,N_11150,N_11289);
or U12790 (N_12790,N_11425,N_11910);
nand U12791 (N_12791,N_11434,N_11241);
nand U12792 (N_12792,N_11230,N_11772);
xor U12793 (N_12793,N_11920,N_11679);
and U12794 (N_12794,N_11731,N_11728);
nand U12795 (N_12795,N_11095,N_11048);
xnor U12796 (N_12796,N_11338,N_11420);
or U12797 (N_12797,N_11392,N_11376);
xnor U12798 (N_12798,N_11240,N_11642);
or U12799 (N_12799,N_11149,N_11811);
and U12800 (N_12800,N_11848,N_11847);
xor U12801 (N_12801,N_11305,N_11403);
nand U12802 (N_12802,N_11380,N_11354);
xor U12803 (N_12803,N_11201,N_11514);
and U12804 (N_12804,N_11165,N_11913);
nor U12805 (N_12805,N_11212,N_11321);
nor U12806 (N_12806,N_11255,N_11603);
or U12807 (N_12807,N_11759,N_11015);
nor U12808 (N_12808,N_11184,N_11007);
xor U12809 (N_12809,N_11941,N_11879);
or U12810 (N_12810,N_11559,N_11060);
or U12811 (N_12811,N_11380,N_11677);
xnor U12812 (N_12812,N_11604,N_11489);
nor U12813 (N_12813,N_11968,N_11299);
or U12814 (N_12814,N_11852,N_11209);
and U12815 (N_12815,N_11607,N_11125);
nor U12816 (N_12816,N_11411,N_11684);
or U12817 (N_12817,N_11428,N_11111);
nor U12818 (N_12818,N_11115,N_11610);
nor U12819 (N_12819,N_11632,N_11024);
nand U12820 (N_12820,N_11051,N_11370);
and U12821 (N_12821,N_11196,N_11440);
nor U12822 (N_12822,N_11673,N_11950);
or U12823 (N_12823,N_11939,N_11739);
nand U12824 (N_12824,N_11313,N_11128);
xnor U12825 (N_12825,N_11983,N_11223);
and U12826 (N_12826,N_11266,N_11150);
xnor U12827 (N_12827,N_11875,N_11626);
nor U12828 (N_12828,N_11005,N_11342);
or U12829 (N_12829,N_11268,N_11410);
nor U12830 (N_12830,N_11431,N_11037);
nor U12831 (N_12831,N_11564,N_11003);
and U12832 (N_12832,N_11141,N_11870);
xor U12833 (N_12833,N_11487,N_11156);
and U12834 (N_12834,N_11618,N_11989);
or U12835 (N_12835,N_11684,N_11705);
nand U12836 (N_12836,N_11110,N_11287);
and U12837 (N_12837,N_11310,N_11193);
nor U12838 (N_12838,N_11316,N_11661);
and U12839 (N_12839,N_11220,N_11310);
nand U12840 (N_12840,N_11934,N_11110);
xnor U12841 (N_12841,N_11314,N_11849);
nor U12842 (N_12842,N_11316,N_11786);
xor U12843 (N_12843,N_11031,N_11893);
nor U12844 (N_12844,N_11235,N_11894);
or U12845 (N_12845,N_11181,N_11094);
nand U12846 (N_12846,N_11980,N_11291);
nor U12847 (N_12847,N_11214,N_11637);
or U12848 (N_12848,N_11987,N_11920);
nor U12849 (N_12849,N_11675,N_11807);
nand U12850 (N_12850,N_11799,N_11024);
nor U12851 (N_12851,N_11210,N_11873);
nor U12852 (N_12852,N_11237,N_11678);
or U12853 (N_12853,N_11024,N_11124);
and U12854 (N_12854,N_11022,N_11781);
nor U12855 (N_12855,N_11705,N_11120);
xor U12856 (N_12856,N_11081,N_11687);
nand U12857 (N_12857,N_11245,N_11252);
xor U12858 (N_12858,N_11297,N_11561);
and U12859 (N_12859,N_11176,N_11884);
xnor U12860 (N_12860,N_11844,N_11098);
or U12861 (N_12861,N_11175,N_11268);
and U12862 (N_12862,N_11985,N_11045);
xor U12863 (N_12863,N_11496,N_11607);
or U12864 (N_12864,N_11096,N_11935);
xnor U12865 (N_12865,N_11877,N_11267);
nand U12866 (N_12866,N_11841,N_11040);
nor U12867 (N_12867,N_11976,N_11885);
xnor U12868 (N_12868,N_11178,N_11659);
nand U12869 (N_12869,N_11690,N_11229);
and U12870 (N_12870,N_11562,N_11035);
nor U12871 (N_12871,N_11359,N_11373);
xnor U12872 (N_12872,N_11413,N_11717);
nand U12873 (N_12873,N_11483,N_11878);
nor U12874 (N_12874,N_11020,N_11206);
nand U12875 (N_12875,N_11469,N_11750);
xor U12876 (N_12876,N_11236,N_11145);
nand U12877 (N_12877,N_11576,N_11743);
xor U12878 (N_12878,N_11489,N_11707);
or U12879 (N_12879,N_11437,N_11939);
nand U12880 (N_12880,N_11561,N_11259);
nor U12881 (N_12881,N_11819,N_11695);
nor U12882 (N_12882,N_11664,N_11870);
nand U12883 (N_12883,N_11531,N_11715);
nand U12884 (N_12884,N_11541,N_11276);
xor U12885 (N_12885,N_11930,N_11761);
nand U12886 (N_12886,N_11662,N_11986);
nor U12887 (N_12887,N_11091,N_11448);
nor U12888 (N_12888,N_11999,N_11308);
nand U12889 (N_12889,N_11566,N_11272);
xnor U12890 (N_12890,N_11066,N_11385);
nand U12891 (N_12891,N_11136,N_11248);
nor U12892 (N_12892,N_11004,N_11011);
nor U12893 (N_12893,N_11087,N_11846);
or U12894 (N_12894,N_11367,N_11178);
xor U12895 (N_12895,N_11248,N_11700);
or U12896 (N_12896,N_11602,N_11520);
nand U12897 (N_12897,N_11116,N_11023);
xor U12898 (N_12898,N_11117,N_11351);
xor U12899 (N_12899,N_11717,N_11544);
xnor U12900 (N_12900,N_11692,N_11522);
xor U12901 (N_12901,N_11472,N_11709);
nand U12902 (N_12902,N_11071,N_11713);
xor U12903 (N_12903,N_11030,N_11373);
nor U12904 (N_12904,N_11612,N_11644);
and U12905 (N_12905,N_11951,N_11065);
nand U12906 (N_12906,N_11523,N_11191);
xor U12907 (N_12907,N_11406,N_11075);
nor U12908 (N_12908,N_11365,N_11605);
and U12909 (N_12909,N_11141,N_11624);
nor U12910 (N_12910,N_11041,N_11496);
nand U12911 (N_12911,N_11454,N_11584);
nand U12912 (N_12912,N_11075,N_11480);
and U12913 (N_12913,N_11264,N_11972);
nor U12914 (N_12914,N_11766,N_11446);
nand U12915 (N_12915,N_11722,N_11425);
xnor U12916 (N_12916,N_11792,N_11027);
nor U12917 (N_12917,N_11993,N_11565);
or U12918 (N_12918,N_11342,N_11416);
and U12919 (N_12919,N_11612,N_11956);
and U12920 (N_12920,N_11136,N_11575);
or U12921 (N_12921,N_11501,N_11504);
and U12922 (N_12922,N_11866,N_11779);
nand U12923 (N_12923,N_11784,N_11177);
or U12924 (N_12924,N_11821,N_11458);
xor U12925 (N_12925,N_11288,N_11136);
xnor U12926 (N_12926,N_11783,N_11641);
nor U12927 (N_12927,N_11177,N_11958);
nor U12928 (N_12928,N_11186,N_11252);
nor U12929 (N_12929,N_11540,N_11758);
nor U12930 (N_12930,N_11238,N_11467);
or U12931 (N_12931,N_11977,N_11167);
nor U12932 (N_12932,N_11242,N_11200);
nand U12933 (N_12933,N_11100,N_11380);
xor U12934 (N_12934,N_11565,N_11624);
nor U12935 (N_12935,N_11990,N_11621);
or U12936 (N_12936,N_11727,N_11168);
and U12937 (N_12937,N_11154,N_11919);
xnor U12938 (N_12938,N_11434,N_11634);
nor U12939 (N_12939,N_11903,N_11772);
nor U12940 (N_12940,N_11289,N_11883);
nand U12941 (N_12941,N_11958,N_11257);
and U12942 (N_12942,N_11506,N_11504);
or U12943 (N_12943,N_11347,N_11456);
and U12944 (N_12944,N_11465,N_11786);
or U12945 (N_12945,N_11193,N_11375);
xor U12946 (N_12946,N_11430,N_11109);
or U12947 (N_12947,N_11996,N_11894);
nand U12948 (N_12948,N_11610,N_11309);
xor U12949 (N_12949,N_11251,N_11371);
xnor U12950 (N_12950,N_11333,N_11343);
xor U12951 (N_12951,N_11931,N_11340);
and U12952 (N_12952,N_11370,N_11577);
nor U12953 (N_12953,N_11132,N_11165);
nand U12954 (N_12954,N_11003,N_11674);
nand U12955 (N_12955,N_11255,N_11752);
nand U12956 (N_12956,N_11822,N_11209);
nand U12957 (N_12957,N_11365,N_11633);
and U12958 (N_12958,N_11660,N_11126);
nand U12959 (N_12959,N_11601,N_11134);
nand U12960 (N_12960,N_11037,N_11794);
xor U12961 (N_12961,N_11015,N_11261);
nor U12962 (N_12962,N_11059,N_11653);
nand U12963 (N_12963,N_11745,N_11140);
nand U12964 (N_12964,N_11318,N_11398);
and U12965 (N_12965,N_11918,N_11081);
nand U12966 (N_12966,N_11487,N_11399);
nor U12967 (N_12967,N_11997,N_11964);
or U12968 (N_12968,N_11795,N_11495);
nor U12969 (N_12969,N_11479,N_11161);
nor U12970 (N_12970,N_11220,N_11894);
nand U12971 (N_12971,N_11268,N_11378);
or U12972 (N_12972,N_11480,N_11484);
nor U12973 (N_12973,N_11107,N_11860);
or U12974 (N_12974,N_11493,N_11822);
nor U12975 (N_12975,N_11728,N_11697);
nand U12976 (N_12976,N_11307,N_11352);
xor U12977 (N_12977,N_11732,N_11008);
nand U12978 (N_12978,N_11902,N_11215);
nor U12979 (N_12979,N_11993,N_11140);
and U12980 (N_12980,N_11715,N_11510);
and U12981 (N_12981,N_11574,N_11570);
or U12982 (N_12982,N_11311,N_11348);
xor U12983 (N_12983,N_11012,N_11261);
nand U12984 (N_12984,N_11707,N_11512);
xnor U12985 (N_12985,N_11796,N_11605);
and U12986 (N_12986,N_11686,N_11724);
nor U12987 (N_12987,N_11138,N_11056);
or U12988 (N_12988,N_11401,N_11780);
nand U12989 (N_12989,N_11809,N_11726);
or U12990 (N_12990,N_11046,N_11247);
nand U12991 (N_12991,N_11177,N_11715);
xnor U12992 (N_12992,N_11047,N_11361);
xnor U12993 (N_12993,N_11666,N_11382);
and U12994 (N_12994,N_11079,N_11366);
xor U12995 (N_12995,N_11131,N_11378);
xor U12996 (N_12996,N_11689,N_11764);
nand U12997 (N_12997,N_11820,N_11398);
or U12998 (N_12998,N_11623,N_11063);
nor U12999 (N_12999,N_11525,N_11518);
nor U13000 (N_13000,N_12459,N_12834);
nand U13001 (N_13001,N_12288,N_12844);
nand U13002 (N_13002,N_12989,N_12967);
or U13003 (N_13003,N_12436,N_12871);
xor U13004 (N_13004,N_12371,N_12014);
nor U13005 (N_13005,N_12317,N_12074);
nor U13006 (N_13006,N_12617,N_12150);
or U13007 (N_13007,N_12772,N_12688);
and U13008 (N_13008,N_12455,N_12646);
or U13009 (N_13009,N_12940,N_12079);
nor U13010 (N_13010,N_12209,N_12846);
nor U13011 (N_13011,N_12979,N_12187);
or U13012 (N_13012,N_12765,N_12909);
and U13013 (N_13013,N_12190,N_12970);
nand U13014 (N_13014,N_12097,N_12193);
nor U13015 (N_13015,N_12867,N_12167);
and U13016 (N_13016,N_12432,N_12521);
or U13017 (N_13017,N_12286,N_12356);
or U13018 (N_13018,N_12959,N_12639);
nor U13019 (N_13019,N_12331,N_12069);
nand U13020 (N_13020,N_12489,N_12073);
or U13021 (N_13021,N_12121,N_12389);
and U13022 (N_13022,N_12166,N_12279);
or U13023 (N_13023,N_12610,N_12674);
xor U13024 (N_13024,N_12386,N_12008);
nand U13025 (N_13025,N_12434,N_12130);
or U13026 (N_13026,N_12559,N_12125);
nand U13027 (N_13027,N_12430,N_12025);
nor U13028 (N_13028,N_12128,N_12343);
xnor U13029 (N_13029,N_12315,N_12813);
xor U13030 (N_13030,N_12318,N_12786);
nand U13031 (N_13031,N_12024,N_12608);
nor U13032 (N_13032,N_12418,N_12974);
nand U13033 (N_13033,N_12466,N_12810);
or U13034 (N_13034,N_12872,N_12722);
nand U13035 (N_13035,N_12127,N_12376);
nand U13036 (N_13036,N_12023,N_12740);
and U13037 (N_13037,N_12769,N_12677);
and U13038 (N_13038,N_12754,N_12163);
or U13039 (N_13039,N_12523,N_12714);
xnor U13040 (N_13040,N_12388,N_12529);
nor U13041 (N_13041,N_12063,N_12986);
and U13042 (N_13042,N_12177,N_12732);
nor U13043 (N_13043,N_12377,N_12906);
nor U13044 (N_13044,N_12589,N_12304);
xnor U13045 (N_13045,N_12835,N_12435);
and U13046 (N_13046,N_12351,N_12933);
and U13047 (N_13047,N_12893,N_12445);
or U13048 (N_13048,N_12349,N_12293);
nor U13049 (N_13049,N_12486,N_12873);
xor U13050 (N_13050,N_12945,N_12483);
and U13051 (N_13051,N_12615,N_12464);
or U13052 (N_13052,N_12105,N_12258);
nor U13053 (N_13053,N_12492,N_12424);
xnor U13054 (N_13054,N_12977,N_12876);
or U13055 (N_13055,N_12325,N_12515);
nand U13056 (N_13056,N_12720,N_12509);
or U13057 (N_13057,N_12482,N_12021);
and U13058 (N_13058,N_12863,N_12238);
or U13059 (N_13059,N_12645,N_12660);
nand U13060 (N_13060,N_12973,N_12763);
xor U13061 (N_13061,N_12890,N_12273);
and U13062 (N_13062,N_12852,N_12228);
nand U13063 (N_13063,N_12067,N_12093);
and U13064 (N_13064,N_12943,N_12930);
nor U13065 (N_13065,N_12854,N_12172);
nand U13066 (N_13066,N_12691,N_12108);
nand U13067 (N_13067,N_12029,N_12045);
nand U13068 (N_13068,N_12874,N_12348);
nand U13069 (N_13069,N_12118,N_12707);
nand U13070 (N_13070,N_12946,N_12694);
and U13071 (N_13071,N_12632,N_12442);
xor U13072 (N_13072,N_12584,N_12923);
and U13073 (N_13073,N_12089,N_12953);
nor U13074 (N_13074,N_12672,N_12991);
or U13075 (N_13075,N_12947,N_12965);
nand U13076 (N_13076,N_12992,N_12746);
xor U13077 (N_13077,N_12247,N_12888);
and U13078 (N_13078,N_12282,N_12496);
xnor U13079 (N_13079,N_12058,N_12100);
and U13080 (N_13080,N_12295,N_12227);
and U13081 (N_13081,N_12107,N_12086);
nand U13082 (N_13082,N_12537,N_12360);
and U13083 (N_13083,N_12547,N_12636);
or U13084 (N_13084,N_12626,N_12091);
and U13085 (N_13085,N_12613,N_12160);
or U13086 (N_13086,N_12836,N_12422);
or U13087 (N_13087,N_12257,N_12594);
and U13088 (N_13088,N_12312,N_12679);
xnor U13089 (N_13089,N_12310,N_12218);
or U13090 (N_13090,N_12016,N_12503);
nand U13091 (N_13091,N_12805,N_12362);
or U13092 (N_13092,N_12733,N_12938);
xor U13093 (N_13093,N_12565,N_12548);
nand U13094 (N_13094,N_12598,N_12592);
xnor U13095 (N_13095,N_12781,N_12398);
xnor U13096 (N_13096,N_12819,N_12140);
nand U13097 (N_13097,N_12994,N_12614);
nand U13098 (N_13098,N_12178,N_12920);
and U13099 (N_13099,N_12612,N_12135);
nor U13100 (N_13100,N_12787,N_12124);
xor U13101 (N_13101,N_12400,N_12170);
and U13102 (N_13102,N_12018,N_12887);
or U13103 (N_13103,N_12477,N_12301);
or U13104 (N_13104,N_12937,N_12233);
and U13105 (N_13105,N_12364,N_12001);
or U13106 (N_13106,N_12568,N_12065);
or U13107 (N_13107,N_12651,N_12879);
xor U13108 (N_13108,N_12882,N_12320);
or U13109 (N_13109,N_12080,N_12927);
or U13110 (N_13110,N_12721,N_12062);
and U13111 (N_13111,N_12809,N_12028);
or U13112 (N_13112,N_12444,N_12112);
nor U13113 (N_13113,N_12984,N_12066);
xnor U13114 (N_13114,N_12750,N_12857);
nor U13115 (N_13115,N_12749,N_12499);
and U13116 (N_13116,N_12054,N_12072);
xnor U13117 (N_13117,N_12277,N_12043);
or U13118 (N_13118,N_12236,N_12372);
nor U13119 (N_13119,N_12302,N_12332);
nand U13120 (N_13120,N_12734,N_12294);
nand U13121 (N_13121,N_12159,N_12220);
nor U13122 (N_13122,N_12952,N_12420);
nor U13123 (N_13123,N_12534,N_12980);
nor U13124 (N_13124,N_12168,N_12189);
xor U13125 (N_13125,N_12131,N_12094);
or U13126 (N_13126,N_12602,N_12246);
nor U13127 (N_13127,N_12206,N_12911);
xnor U13128 (N_13128,N_12245,N_12510);
xor U13129 (N_13129,N_12768,N_12030);
nand U13130 (N_13130,N_12458,N_12048);
xnor U13131 (N_13131,N_12824,N_12794);
xor U13132 (N_13132,N_12078,N_12629);
or U13133 (N_13133,N_12725,N_12081);
nor U13134 (N_13134,N_12155,N_12950);
and U13135 (N_13135,N_12498,N_12531);
nor U13136 (N_13136,N_12902,N_12773);
or U13137 (N_13137,N_12962,N_12248);
nor U13138 (N_13138,N_12517,N_12524);
or U13139 (N_13139,N_12525,N_12745);
xor U13140 (N_13140,N_12151,N_12441);
or U13141 (N_13141,N_12268,N_12346);
nand U13142 (N_13142,N_12922,N_12514);
and U13143 (N_13143,N_12575,N_12801);
nand U13144 (N_13144,N_12504,N_12497);
and U13145 (N_13145,N_12657,N_12582);
nand U13146 (N_13146,N_12735,N_12068);
or U13147 (N_13147,N_12242,N_12821);
and U13148 (N_13148,N_12693,N_12505);
nand U13149 (N_13149,N_12174,N_12040);
nand U13150 (N_13150,N_12738,N_12713);
xnor U13151 (N_13151,N_12830,N_12410);
nor U13152 (N_13152,N_12433,N_12392);
or U13153 (N_13153,N_12766,N_12742);
nor U13154 (N_13154,N_12811,N_12676);
or U13155 (N_13155,N_12032,N_12196);
nor U13156 (N_13156,N_12240,N_12642);
or U13157 (N_13157,N_12143,N_12431);
or U13158 (N_13158,N_12051,N_12250);
nor U13159 (N_13159,N_12222,N_12931);
nor U13160 (N_13160,N_12269,N_12580);
and U13161 (N_13161,N_12491,N_12957);
nor U13162 (N_13162,N_12421,N_12387);
and U13163 (N_13163,N_12020,N_12638);
and U13164 (N_13164,N_12506,N_12280);
nor U13165 (N_13165,N_12005,N_12144);
nand U13166 (N_13166,N_12129,N_12481);
nor U13167 (N_13167,N_12415,N_12528);
and U13168 (N_13168,N_12347,N_12402);
nor U13169 (N_13169,N_12327,N_12982);
nand U13170 (N_13170,N_12955,N_12847);
xor U13171 (N_13171,N_12964,N_12000);
nand U13172 (N_13172,N_12208,N_12695);
or U13173 (N_13173,N_12539,N_12319);
and U13174 (N_13174,N_12335,N_12194);
and U13175 (N_13175,N_12285,N_12013);
nand U13176 (N_13176,N_12426,N_12554);
xnor U13177 (N_13177,N_12803,N_12535);
nor U13178 (N_13178,N_12485,N_12399);
or U13179 (N_13179,N_12244,N_12199);
or U13180 (N_13180,N_12156,N_12390);
xnor U13181 (N_13181,N_12487,N_12047);
and U13182 (N_13182,N_12900,N_12022);
nor U13183 (N_13183,N_12195,N_12833);
nand U13184 (N_13184,N_12479,N_12702);
nor U13185 (N_13185,N_12885,N_12493);
and U13186 (N_13186,N_12508,N_12184);
nor U13187 (N_13187,N_12814,N_12019);
xor U13188 (N_13188,N_12407,N_12292);
nand U13189 (N_13189,N_12126,N_12321);
nand U13190 (N_13190,N_12985,N_12717);
nand U13191 (N_13191,N_12684,N_12744);
xor U13192 (N_13192,N_12712,N_12858);
nor U13193 (N_13193,N_12404,N_12776);
and U13194 (N_13194,N_12624,N_12743);
and U13195 (N_13195,N_12186,N_12010);
and U13196 (N_13196,N_12255,N_12700);
nand U13197 (N_13197,N_12138,N_12842);
xnor U13198 (N_13198,N_12837,N_12755);
xnor U13199 (N_13199,N_12342,N_12604);
xor U13200 (N_13200,N_12012,N_12104);
and U13201 (N_13201,N_12035,N_12739);
nor U13202 (N_13202,N_12207,N_12061);
nor U13203 (N_13203,N_12549,N_12843);
nand U13204 (N_13204,N_12550,N_12411);
nand U13205 (N_13205,N_12116,N_12046);
nand U13206 (N_13206,N_12403,N_12033);
nand U13207 (N_13207,N_12910,N_12587);
nand U13208 (N_13208,N_12270,N_12782);
nor U13209 (N_13209,N_12800,N_12339);
or U13210 (N_13210,N_12928,N_12730);
nor U13211 (N_13211,N_12087,N_12899);
and U13212 (N_13212,N_12158,N_12203);
nand U13213 (N_13213,N_12494,N_12262);
or U13214 (N_13214,N_12103,N_12241);
nor U13215 (N_13215,N_12948,N_12380);
or U13216 (N_13216,N_12522,N_12903);
or U13217 (N_13217,N_12353,N_12818);
xnor U13218 (N_13218,N_12662,N_12059);
or U13219 (N_13219,N_12060,N_12469);
and U13220 (N_13220,N_12780,N_12289);
or U13221 (N_13221,N_12988,N_12309);
or U13222 (N_13222,N_12468,N_12077);
and U13223 (N_13223,N_12849,N_12221);
nand U13224 (N_13224,N_12519,N_12164);
xnor U13225 (N_13225,N_12741,N_12049);
nand U13226 (N_13226,N_12095,N_12394);
nand U13227 (N_13227,N_12748,N_12230);
nor U13228 (N_13228,N_12401,N_12098);
nor U13229 (N_13229,N_12188,N_12647);
xor U13230 (N_13230,N_12926,N_12284);
nand U13231 (N_13231,N_12179,N_12939);
or U13232 (N_13232,N_12460,N_12577);
nand U13233 (N_13233,N_12708,N_12239);
or U13234 (N_13234,N_12644,N_12832);
or U13235 (N_13235,N_12263,N_12884);
xnor U13236 (N_13236,N_12307,N_12042);
xor U13237 (N_13237,N_12605,N_12454);
nor U13238 (N_13238,N_12526,N_12113);
nor U13239 (N_13239,N_12572,N_12251);
and U13240 (N_13240,N_12202,N_12655);
or U13241 (N_13241,N_12929,N_12359);
nor U13242 (N_13242,N_12855,N_12419);
and U13243 (N_13243,N_12132,N_12070);
or U13244 (N_13244,N_12971,N_12588);
xor U13245 (N_13245,N_12696,N_12804);
nor U13246 (N_13246,N_12393,N_12681);
xor U13247 (N_13247,N_12234,N_12259);
or U13248 (N_13248,N_12663,N_12229);
nand U13249 (N_13249,N_12998,N_12231);
nor U13250 (N_13250,N_12664,N_12428);
and U13251 (N_13251,N_12341,N_12527);
xnor U13252 (N_13252,N_12115,N_12075);
and U13253 (N_13253,N_12999,N_12729);
nor U13254 (N_13254,N_12452,N_12011);
xor U13255 (N_13255,N_12057,N_12546);
and U13256 (N_13256,N_12266,N_12055);
or U13257 (N_13257,N_12366,N_12003);
or U13258 (N_13258,N_12542,N_12593);
and U13259 (N_13259,N_12275,N_12916);
nand U13260 (N_13260,N_12606,N_12567);
nor U13261 (N_13261,N_12328,N_12507);
and U13262 (N_13262,N_12137,N_12983);
nor U13263 (N_13263,N_12864,N_12774);
xnor U13264 (N_13264,N_12253,N_12976);
xnor U13265 (N_13265,N_12934,N_12449);
xnor U13266 (N_13266,N_12513,N_12840);
xor U13267 (N_13267,N_12495,N_12373);
or U13268 (N_13268,N_12566,N_12490);
or U13269 (N_13269,N_12978,N_12771);
nand U13270 (N_13270,N_12082,N_12648);
nor U13271 (N_13271,N_12039,N_12958);
or U13272 (N_13272,N_12185,N_12162);
or U13273 (N_13273,N_12017,N_12412);
and U13274 (N_13274,N_12026,N_12682);
or U13275 (N_13275,N_12053,N_12966);
xor U13276 (N_13276,N_12905,N_12789);
nand U13277 (N_13277,N_12261,N_12314);
xnor U13278 (N_13278,N_12281,N_12409);
nor U13279 (N_13279,N_12171,N_12471);
xnor U13280 (N_13280,N_12106,N_12050);
nand U13281 (N_13281,N_12395,N_12204);
or U13282 (N_13282,N_12564,N_12705);
nand U13283 (N_13283,N_12114,N_12201);
nand U13284 (N_13284,N_12555,N_12827);
or U13285 (N_13285,N_12904,N_12633);
xnor U13286 (N_13286,N_12627,N_12146);
nor U13287 (N_13287,N_12747,N_12429);
nand U13288 (N_13288,N_12601,N_12792);
nand U13289 (N_13289,N_12438,N_12191);
or U13290 (N_13290,N_12573,N_12668);
or U13291 (N_13291,N_12607,N_12272);
xnor U13292 (N_13292,N_12751,N_12340);
nand U13293 (N_13293,N_12044,N_12102);
or U13294 (N_13294,N_12894,N_12551);
xnor U13295 (N_13295,N_12853,N_12276);
nand U13296 (N_13296,N_12216,N_12862);
or U13297 (N_13297,N_12153,N_12678);
or U13298 (N_13298,N_12540,N_12583);
nor U13299 (N_13299,N_12192,N_12088);
and U13300 (N_13300,N_12440,N_12709);
or U13301 (N_13301,N_12793,N_12673);
or U13302 (N_13302,N_12635,N_12385);
or U13303 (N_13303,N_12161,N_12777);
xnor U13304 (N_13304,N_12149,N_12576);
nand U13305 (N_13305,N_12569,N_12267);
xnor U13306 (N_13306,N_12951,N_12297);
xnor U13307 (N_13307,N_12363,N_12456);
or U13308 (N_13308,N_12841,N_12532);
or U13309 (N_13309,N_12037,N_12993);
or U13310 (N_13310,N_12868,N_12384);
nor U13311 (N_13311,N_12649,N_12352);
or U13312 (N_13312,N_12512,N_12791);
xor U13313 (N_13313,N_12182,N_12715);
xnor U13314 (N_13314,N_12210,N_12071);
nor U13315 (N_13315,N_12806,N_12620);
nand U13316 (N_13316,N_12470,N_12052);
xor U13317 (N_13317,N_12439,N_12990);
or U13318 (N_13318,N_12880,N_12147);
or U13319 (N_13319,N_12690,N_12306);
xnor U13320 (N_13320,N_12446,N_12892);
and U13321 (N_13321,N_12912,N_12213);
nand U13322 (N_13322,N_12616,N_12981);
nor U13323 (N_13323,N_12680,N_12562);
nand U13324 (N_13324,N_12856,N_12585);
xor U13325 (N_13325,N_12311,N_12169);
xor U13326 (N_13326,N_12571,N_12232);
nand U13327 (N_13327,N_12084,N_12790);
xor U13328 (N_13328,N_12618,N_12543);
or U13329 (N_13329,N_12692,N_12807);
and U13330 (N_13330,N_12622,N_12101);
nor U13331 (N_13331,N_12578,N_12706);
nor U13332 (N_13332,N_12447,N_12932);
xnor U13333 (N_13333,N_12111,N_12536);
or U13334 (N_13334,N_12637,N_12226);
nand U13335 (N_13335,N_12139,N_12889);
xor U13336 (N_13336,N_12538,N_12689);
nand U13337 (N_13337,N_12368,N_12518);
and U13338 (N_13338,N_12064,N_12154);
nand U13339 (N_13339,N_12461,N_12784);
or U13340 (N_13340,N_12775,N_12041);
and U13341 (N_13341,N_12326,N_12961);
or U13342 (N_13342,N_12656,N_12558);
nor U13343 (N_13343,N_12731,N_12324);
xor U13344 (N_13344,N_12254,N_12181);
nor U13345 (N_13345,N_12628,N_12728);
xor U13346 (N_13346,N_12355,N_12770);
nand U13347 (N_13347,N_12703,N_12625);
and U13348 (N_13348,N_12623,N_12886);
and U13349 (N_13349,N_12756,N_12675);
or U13350 (N_13350,N_12848,N_12367);
and U13351 (N_13351,N_12704,N_12595);
and U13352 (N_13352,N_12278,N_12345);
xnor U13353 (N_13353,N_12724,N_12643);
xor U13354 (N_13354,N_12831,N_12370);
or U13355 (N_13355,N_12264,N_12375);
nand U13356 (N_13356,N_12451,N_12329);
and U13357 (N_13357,N_12076,N_12260);
or U13358 (N_13358,N_12785,N_12381);
nor U13359 (N_13359,N_12788,N_12472);
xnor U13360 (N_13360,N_12820,N_12133);
nand U13361 (N_13361,N_12736,N_12038);
nor U13362 (N_13362,N_12414,N_12300);
or U13363 (N_13363,N_12323,N_12453);
nand U13364 (N_13364,N_12249,N_12925);
nand U13365 (N_13365,N_12511,N_12015);
nand U13366 (N_13366,N_12009,N_12716);
nand U13367 (N_13367,N_12579,N_12090);
xnor U13368 (N_13368,N_12764,N_12850);
nor U13369 (N_13369,N_12563,N_12274);
nand U13370 (N_13370,N_12621,N_12305);
nand U13371 (N_13371,N_12619,N_12099);
and U13372 (N_13372,N_12223,N_12987);
and U13373 (N_13373,N_12574,N_12336);
nand U13374 (N_13374,N_12313,N_12463);
nor U13375 (N_13375,N_12596,N_12891);
and U13376 (N_13376,N_12557,N_12816);
or U13377 (N_13377,N_12176,N_12590);
xor U13378 (N_13378,N_12413,N_12205);
or U13379 (N_13379,N_12767,N_12896);
and U13380 (N_13380,N_12797,N_12500);
nand U13381 (N_13381,N_12779,N_12119);
and U13382 (N_13382,N_12802,N_12895);
nand U13383 (N_13383,N_12556,N_12936);
nand U13384 (N_13384,N_12611,N_12520);
or U13385 (N_13385,N_12036,N_12530);
nand U13386 (N_13386,N_12473,N_12711);
and U13387 (N_13387,N_12322,N_12671);
nand U13388 (N_13388,N_12180,N_12303);
or U13389 (N_13389,N_12183,N_12484);
or U13390 (N_13390,N_12443,N_12723);
nand U13391 (N_13391,N_12898,N_12669);
and U13392 (N_13392,N_12215,N_12397);
nand U13393 (N_13393,N_12173,N_12545);
nand U13394 (N_13394,N_12252,N_12283);
nand U13395 (N_13395,N_12737,N_12851);
and U13396 (N_13396,N_12027,N_12878);
nor U13397 (N_13397,N_12727,N_12365);
xnor U13398 (N_13398,N_12225,N_12369);
or U13399 (N_13399,N_12337,N_12609);
nor U13400 (N_13400,N_12865,N_12408);
nor U13401 (N_13401,N_12726,N_12997);
or U13402 (N_13402,N_12142,N_12901);
and U13403 (N_13403,N_12148,N_12007);
xnor U13404 (N_13404,N_12631,N_12815);
or U13405 (N_13405,N_12975,N_12652);
nor U13406 (N_13406,N_12561,N_12719);
and U13407 (N_13407,N_12759,N_12838);
or U13408 (N_13408,N_12686,N_12581);
xor U13409 (N_13409,N_12760,N_12913);
xor U13410 (N_13410,N_12197,N_12467);
nand U13411 (N_13411,N_12544,N_12870);
nor U13412 (N_13412,N_12996,N_12823);
or U13413 (N_13413,N_12425,N_12476);
and U13414 (N_13414,N_12416,N_12860);
and U13415 (N_13415,N_12591,N_12457);
nand U13416 (N_13416,N_12333,N_12718);
nor U13417 (N_13417,N_12214,N_12299);
and U13418 (N_13418,N_12271,N_12822);
or U13419 (N_13419,N_12552,N_12758);
or U13420 (N_13420,N_12211,N_12866);
or U13421 (N_13421,N_12883,N_12110);
nor U13422 (N_13422,N_12004,N_12031);
nand U13423 (N_13423,N_12560,N_12845);
or U13424 (N_13424,N_12963,N_12861);
or U13425 (N_13425,N_12212,N_12448);
and U13426 (N_13426,N_12480,N_12350);
nor U13427 (N_13427,N_12478,N_12956);
xnor U13428 (N_13428,N_12316,N_12501);
xnor U13429 (N_13429,N_12219,N_12437);
nor U13430 (N_13430,N_12995,N_12699);
and U13431 (N_13431,N_12761,N_12829);
nand U13432 (N_13432,N_12698,N_12600);
or U13433 (N_13433,N_12379,N_12122);
or U13434 (N_13434,N_12570,N_12915);
xor U13435 (N_13435,N_12917,N_12198);
or U13436 (N_13436,N_12907,N_12757);
and U13437 (N_13437,N_12145,N_12291);
nand U13438 (N_13438,N_12641,N_12488);
xor U13439 (N_13439,N_12083,N_12296);
nor U13440 (N_13440,N_12361,N_12200);
or U13441 (N_13441,N_12085,N_12808);
nand U13442 (N_13442,N_12960,N_12235);
xnor U13443 (N_13443,N_12897,N_12908);
and U13444 (N_13444,N_12117,N_12949);
nand U13445 (N_13445,N_12382,N_12374);
and U13446 (N_13446,N_12034,N_12541);
xor U13447 (N_13447,N_12175,N_12881);
xnor U13448 (N_13448,N_12465,N_12687);
xor U13449 (N_13449,N_12136,N_12599);
or U13450 (N_13450,N_12914,N_12634);
nand U13451 (N_13451,N_12092,N_12826);
nor U13452 (N_13452,N_12357,N_12290);
or U13453 (N_13453,N_12796,N_12683);
and U13454 (N_13454,N_12006,N_12330);
nand U13455 (N_13455,N_12877,N_12869);
xnor U13456 (N_13456,N_12654,N_12666);
or U13457 (N_13457,N_12391,N_12954);
nor U13458 (N_13458,N_12661,N_12096);
or U13459 (N_13459,N_12405,N_12002);
xnor U13460 (N_13460,N_12141,N_12056);
xor U13461 (N_13461,N_12224,N_12795);
nand U13462 (N_13462,N_12423,N_12653);
or U13463 (N_13463,N_12798,N_12640);
nand U13464 (N_13464,N_12338,N_12968);
nor U13465 (N_13465,N_12697,N_12685);
and U13466 (N_13466,N_12134,N_12354);
and U13467 (N_13467,N_12378,N_12817);
or U13468 (N_13468,N_12120,N_12217);
nand U13469 (N_13469,N_12859,N_12924);
nand U13470 (N_13470,N_12603,N_12701);
nor U13471 (N_13471,N_12553,N_12710);
xnor U13472 (N_13472,N_12237,N_12969);
xor U13473 (N_13473,N_12778,N_12533);
or U13474 (N_13474,N_12109,N_12935);
nand U13475 (N_13475,N_12243,N_12475);
nand U13476 (N_13476,N_12972,N_12650);
or U13477 (N_13477,N_12630,N_12396);
nor U13478 (N_13478,N_12670,N_12753);
or U13479 (N_13479,N_12502,N_12658);
nand U13480 (N_13480,N_12752,N_12918);
xnor U13481 (N_13481,N_12586,N_12875);
or U13482 (N_13482,N_12762,N_12123);
and U13483 (N_13483,N_12665,N_12919);
nor U13484 (N_13484,N_12165,N_12667);
nor U13485 (N_13485,N_12256,N_12157);
and U13486 (N_13486,N_12828,N_12921);
or U13487 (N_13487,N_12417,N_12659);
nand U13488 (N_13488,N_12344,N_12839);
nand U13489 (N_13489,N_12597,N_12783);
nand U13490 (N_13490,N_12825,N_12298);
xor U13491 (N_13491,N_12799,N_12942);
nand U13492 (N_13492,N_12516,N_12287);
nand U13493 (N_13493,N_12474,N_12265);
nor U13494 (N_13494,N_12812,N_12450);
nand U13495 (N_13495,N_12358,N_12308);
xnor U13496 (N_13496,N_12944,N_12462);
xnor U13497 (N_13497,N_12941,N_12427);
nor U13498 (N_13498,N_12383,N_12334);
xnor U13499 (N_13499,N_12406,N_12152);
and U13500 (N_13500,N_12551,N_12605);
and U13501 (N_13501,N_12306,N_12002);
nor U13502 (N_13502,N_12750,N_12938);
or U13503 (N_13503,N_12892,N_12748);
or U13504 (N_13504,N_12328,N_12019);
nor U13505 (N_13505,N_12698,N_12599);
nand U13506 (N_13506,N_12856,N_12937);
nor U13507 (N_13507,N_12348,N_12831);
nor U13508 (N_13508,N_12072,N_12258);
nor U13509 (N_13509,N_12173,N_12397);
nand U13510 (N_13510,N_12897,N_12928);
or U13511 (N_13511,N_12920,N_12080);
nor U13512 (N_13512,N_12673,N_12044);
and U13513 (N_13513,N_12672,N_12316);
xor U13514 (N_13514,N_12462,N_12604);
or U13515 (N_13515,N_12099,N_12415);
or U13516 (N_13516,N_12695,N_12389);
nor U13517 (N_13517,N_12281,N_12574);
nand U13518 (N_13518,N_12483,N_12550);
xor U13519 (N_13519,N_12904,N_12892);
and U13520 (N_13520,N_12837,N_12832);
and U13521 (N_13521,N_12861,N_12324);
nand U13522 (N_13522,N_12227,N_12398);
or U13523 (N_13523,N_12590,N_12201);
xor U13524 (N_13524,N_12803,N_12613);
and U13525 (N_13525,N_12454,N_12369);
xor U13526 (N_13526,N_12751,N_12060);
nor U13527 (N_13527,N_12755,N_12190);
and U13528 (N_13528,N_12068,N_12284);
nor U13529 (N_13529,N_12378,N_12159);
and U13530 (N_13530,N_12363,N_12825);
xnor U13531 (N_13531,N_12262,N_12146);
and U13532 (N_13532,N_12654,N_12091);
nand U13533 (N_13533,N_12500,N_12063);
nor U13534 (N_13534,N_12597,N_12527);
nand U13535 (N_13535,N_12076,N_12790);
or U13536 (N_13536,N_12922,N_12715);
xnor U13537 (N_13537,N_12770,N_12747);
nor U13538 (N_13538,N_12149,N_12575);
and U13539 (N_13539,N_12243,N_12101);
and U13540 (N_13540,N_12226,N_12959);
or U13541 (N_13541,N_12512,N_12459);
xor U13542 (N_13542,N_12037,N_12613);
or U13543 (N_13543,N_12678,N_12738);
nand U13544 (N_13544,N_12383,N_12375);
nor U13545 (N_13545,N_12604,N_12814);
nand U13546 (N_13546,N_12362,N_12022);
xor U13547 (N_13547,N_12713,N_12903);
or U13548 (N_13548,N_12464,N_12734);
and U13549 (N_13549,N_12049,N_12533);
and U13550 (N_13550,N_12341,N_12544);
and U13551 (N_13551,N_12862,N_12684);
nand U13552 (N_13552,N_12037,N_12127);
xor U13553 (N_13553,N_12631,N_12310);
nand U13554 (N_13554,N_12549,N_12519);
xor U13555 (N_13555,N_12102,N_12695);
and U13556 (N_13556,N_12781,N_12626);
and U13557 (N_13557,N_12695,N_12139);
xor U13558 (N_13558,N_12738,N_12851);
xnor U13559 (N_13559,N_12569,N_12195);
and U13560 (N_13560,N_12754,N_12257);
nand U13561 (N_13561,N_12707,N_12165);
xor U13562 (N_13562,N_12417,N_12279);
xnor U13563 (N_13563,N_12197,N_12837);
or U13564 (N_13564,N_12720,N_12984);
nand U13565 (N_13565,N_12445,N_12861);
or U13566 (N_13566,N_12460,N_12542);
and U13567 (N_13567,N_12743,N_12028);
nand U13568 (N_13568,N_12074,N_12105);
xnor U13569 (N_13569,N_12142,N_12210);
nand U13570 (N_13570,N_12628,N_12961);
nor U13571 (N_13571,N_12360,N_12046);
xor U13572 (N_13572,N_12663,N_12536);
xor U13573 (N_13573,N_12672,N_12527);
nor U13574 (N_13574,N_12475,N_12752);
xnor U13575 (N_13575,N_12737,N_12768);
or U13576 (N_13576,N_12679,N_12049);
nor U13577 (N_13577,N_12146,N_12803);
nor U13578 (N_13578,N_12408,N_12240);
and U13579 (N_13579,N_12967,N_12802);
xor U13580 (N_13580,N_12689,N_12739);
nor U13581 (N_13581,N_12590,N_12109);
nand U13582 (N_13582,N_12595,N_12396);
and U13583 (N_13583,N_12519,N_12783);
xnor U13584 (N_13584,N_12718,N_12853);
nor U13585 (N_13585,N_12072,N_12020);
nor U13586 (N_13586,N_12304,N_12921);
or U13587 (N_13587,N_12080,N_12694);
xor U13588 (N_13588,N_12990,N_12079);
and U13589 (N_13589,N_12501,N_12698);
nor U13590 (N_13590,N_12337,N_12150);
nand U13591 (N_13591,N_12164,N_12598);
nand U13592 (N_13592,N_12928,N_12318);
or U13593 (N_13593,N_12496,N_12151);
nor U13594 (N_13594,N_12095,N_12966);
and U13595 (N_13595,N_12955,N_12848);
nor U13596 (N_13596,N_12550,N_12699);
nor U13597 (N_13597,N_12267,N_12499);
or U13598 (N_13598,N_12725,N_12024);
and U13599 (N_13599,N_12526,N_12561);
nor U13600 (N_13600,N_12829,N_12198);
nor U13601 (N_13601,N_12084,N_12364);
nor U13602 (N_13602,N_12114,N_12616);
and U13603 (N_13603,N_12194,N_12724);
or U13604 (N_13604,N_12618,N_12144);
nand U13605 (N_13605,N_12066,N_12830);
nor U13606 (N_13606,N_12121,N_12838);
xor U13607 (N_13607,N_12761,N_12158);
xnor U13608 (N_13608,N_12540,N_12796);
or U13609 (N_13609,N_12087,N_12934);
xor U13610 (N_13610,N_12945,N_12160);
nor U13611 (N_13611,N_12559,N_12597);
or U13612 (N_13612,N_12381,N_12343);
nor U13613 (N_13613,N_12036,N_12843);
nor U13614 (N_13614,N_12027,N_12372);
and U13615 (N_13615,N_12162,N_12367);
and U13616 (N_13616,N_12893,N_12962);
nor U13617 (N_13617,N_12709,N_12295);
nor U13618 (N_13618,N_12273,N_12860);
xnor U13619 (N_13619,N_12461,N_12950);
nand U13620 (N_13620,N_12787,N_12404);
or U13621 (N_13621,N_12664,N_12971);
nand U13622 (N_13622,N_12525,N_12044);
xor U13623 (N_13623,N_12785,N_12185);
nand U13624 (N_13624,N_12074,N_12295);
or U13625 (N_13625,N_12644,N_12240);
nor U13626 (N_13626,N_12528,N_12177);
or U13627 (N_13627,N_12608,N_12335);
xor U13628 (N_13628,N_12490,N_12008);
nand U13629 (N_13629,N_12851,N_12139);
nor U13630 (N_13630,N_12827,N_12942);
xnor U13631 (N_13631,N_12277,N_12843);
nand U13632 (N_13632,N_12088,N_12164);
nor U13633 (N_13633,N_12330,N_12220);
nand U13634 (N_13634,N_12664,N_12715);
and U13635 (N_13635,N_12666,N_12219);
or U13636 (N_13636,N_12501,N_12854);
nor U13637 (N_13637,N_12133,N_12281);
or U13638 (N_13638,N_12860,N_12289);
xnor U13639 (N_13639,N_12697,N_12827);
nor U13640 (N_13640,N_12581,N_12011);
nand U13641 (N_13641,N_12966,N_12044);
nand U13642 (N_13642,N_12356,N_12348);
and U13643 (N_13643,N_12667,N_12934);
and U13644 (N_13644,N_12345,N_12831);
xnor U13645 (N_13645,N_12351,N_12879);
nand U13646 (N_13646,N_12796,N_12454);
or U13647 (N_13647,N_12374,N_12928);
xor U13648 (N_13648,N_12848,N_12821);
xnor U13649 (N_13649,N_12346,N_12677);
nand U13650 (N_13650,N_12479,N_12049);
xor U13651 (N_13651,N_12014,N_12378);
and U13652 (N_13652,N_12867,N_12721);
or U13653 (N_13653,N_12517,N_12352);
nand U13654 (N_13654,N_12590,N_12702);
nor U13655 (N_13655,N_12603,N_12393);
nor U13656 (N_13656,N_12895,N_12922);
or U13657 (N_13657,N_12149,N_12681);
or U13658 (N_13658,N_12554,N_12836);
or U13659 (N_13659,N_12882,N_12461);
nand U13660 (N_13660,N_12786,N_12613);
nand U13661 (N_13661,N_12114,N_12899);
nor U13662 (N_13662,N_12747,N_12622);
and U13663 (N_13663,N_12061,N_12228);
nor U13664 (N_13664,N_12525,N_12220);
or U13665 (N_13665,N_12037,N_12966);
nor U13666 (N_13666,N_12364,N_12267);
or U13667 (N_13667,N_12827,N_12037);
xor U13668 (N_13668,N_12498,N_12721);
xor U13669 (N_13669,N_12968,N_12515);
xnor U13670 (N_13670,N_12815,N_12992);
xnor U13671 (N_13671,N_12892,N_12597);
xor U13672 (N_13672,N_12054,N_12634);
xor U13673 (N_13673,N_12962,N_12135);
xnor U13674 (N_13674,N_12418,N_12099);
nor U13675 (N_13675,N_12231,N_12596);
xnor U13676 (N_13676,N_12829,N_12458);
nand U13677 (N_13677,N_12976,N_12409);
xor U13678 (N_13678,N_12207,N_12810);
nor U13679 (N_13679,N_12005,N_12380);
nor U13680 (N_13680,N_12741,N_12689);
nand U13681 (N_13681,N_12146,N_12870);
or U13682 (N_13682,N_12802,N_12535);
xor U13683 (N_13683,N_12977,N_12119);
xnor U13684 (N_13684,N_12332,N_12672);
xor U13685 (N_13685,N_12442,N_12133);
or U13686 (N_13686,N_12100,N_12034);
nor U13687 (N_13687,N_12979,N_12139);
nor U13688 (N_13688,N_12178,N_12237);
xnor U13689 (N_13689,N_12014,N_12955);
and U13690 (N_13690,N_12564,N_12658);
nor U13691 (N_13691,N_12931,N_12722);
or U13692 (N_13692,N_12570,N_12275);
nand U13693 (N_13693,N_12033,N_12738);
nor U13694 (N_13694,N_12594,N_12008);
and U13695 (N_13695,N_12273,N_12850);
nor U13696 (N_13696,N_12538,N_12887);
or U13697 (N_13697,N_12235,N_12949);
nor U13698 (N_13698,N_12281,N_12592);
nor U13699 (N_13699,N_12967,N_12181);
and U13700 (N_13700,N_12555,N_12029);
xor U13701 (N_13701,N_12506,N_12771);
or U13702 (N_13702,N_12435,N_12716);
nor U13703 (N_13703,N_12729,N_12664);
and U13704 (N_13704,N_12139,N_12637);
xor U13705 (N_13705,N_12496,N_12300);
nor U13706 (N_13706,N_12019,N_12796);
nor U13707 (N_13707,N_12757,N_12856);
or U13708 (N_13708,N_12323,N_12669);
and U13709 (N_13709,N_12594,N_12114);
nor U13710 (N_13710,N_12211,N_12837);
nor U13711 (N_13711,N_12187,N_12589);
nand U13712 (N_13712,N_12934,N_12553);
nor U13713 (N_13713,N_12209,N_12695);
or U13714 (N_13714,N_12299,N_12543);
xor U13715 (N_13715,N_12770,N_12168);
and U13716 (N_13716,N_12830,N_12822);
and U13717 (N_13717,N_12063,N_12878);
xor U13718 (N_13718,N_12320,N_12649);
or U13719 (N_13719,N_12326,N_12248);
nor U13720 (N_13720,N_12985,N_12681);
nand U13721 (N_13721,N_12279,N_12242);
or U13722 (N_13722,N_12987,N_12926);
and U13723 (N_13723,N_12828,N_12022);
nor U13724 (N_13724,N_12665,N_12553);
xnor U13725 (N_13725,N_12680,N_12442);
and U13726 (N_13726,N_12705,N_12969);
nor U13727 (N_13727,N_12271,N_12931);
or U13728 (N_13728,N_12380,N_12316);
xor U13729 (N_13729,N_12029,N_12727);
or U13730 (N_13730,N_12954,N_12638);
xnor U13731 (N_13731,N_12161,N_12606);
nand U13732 (N_13732,N_12531,N_12830);
xnor U13733 (N_13733,N_12424,N_12845);
nor U13734 (N_13734,N_12926,N_12540);
nand U13735 (N_13735,N_12156,N_12909);
nor U13736 (N_13736,N_12786,N_12219);
xor U13737 (N_13737,N_12553,N_12537);
nand U13738 (N_13738,N_12182,N_12574);
and U13739 (N_13739,N_12651,N_12296);
nand U13740 (N_13740,N_12368,N_12902);
xor U13741 (N_13741,N_12241,N_12362);
xnor U13742 (N_13742,N_12296,N_12533);
or U13743 (N_13743,N_12674,N_12229);
xor U13744 (N_13744,N_12096,N_12436);
xor U13745 (N_13745,N_12736,N_12728);
xnor U13746 (N_13746,N_12571,N_12427);
or U13747 (N_13747,N_12542,N_12984);
nor U13748 (N_13748,N_12416,N_12411);
nand U13749 (N_13749,N_12739,N_12089);
and U13750 (N_13750,N_12513,N_12032);
nand U13751 (N_13751,N_12621,N_12424);
and U13752 (N_13752,N_12685,N_12635);
nor U13753 (N_13753,N_12280,N_12307);
nor U13754 (N_13754,N_12422,N_12807);
nand U13755 (N_13755,N_12370,N_12634);
or U13756 (N_13756,N_12196,N_12831);
or U13757 (N_13757,N_12642,N_12490);
and U13758 (N_13758,N_12300,N_12837);
nor U13759 (N_13759,N_12480,N_12005);
nand U13760 (N_13760,N_12974,N_12362);
and U13761 (N_13761,N_12392,N_12851);
nor U13762 (N_13762,N_12732,N_12859);
nor U13763 (N_13763,N_12122,N_12373);
nor U13764 (N_13764,N_12211,N_12019);
or U13765 (N_13765,N_12502,N_12725);
nand U13766 (N_13766,N_12472,N_12318);
nor U13767 (N_13767,N_12468,N_12271);
nand U13768 (N_13768,N_12164,N_12014);
xnor U13769 (N_13769,N_12540,N_12507);
nand U13770 (N_13770,N_12207,N_12338);
and U13771 (N_13771,N_12297,N_12911);
xor U13772 (N_13772,N_12714,N_12744);
xnor U13773 (N_13773,N_12424,N_12331);
or U13774 (N_13774,N_12503,N_12741);
xnor U13775 (N_13775,N_12987,N_12791);
and U13776 (N_13776,N_12306,N_12909);
nor U13777 (N_13777,N_12158,N_12124);
nor U13778 (N_13778,N_12396,N_12708);
nor U13779 (N_13779,N_12475,N_12468);
xor U13780 (N_13780,N_12091,N_12356);
xnor U13781 (N_13781,N_12658,N_12279);
and U13782 (N_13782,N_12580,N_12994);
nand U13783 (N_13783,N_12185,N_12005);
or U13784 (N_13784,N_12085,N_12359);
xor U13785 (N_13785,N_12618,N_12440);
xor U13786 (N_13786,N_12198,N_12418);
and U13787 (N_13787,N_12228,N_12694);
nor U13788 (N_13788,N_12873,N_12786);
nor U13789 (N_13789,N_12042,N_12655);
or U13790 (N_13790,N_12135,N_12004);
and U13791 (N_13791,N_12723,N_12052);
nand U13792 (N_13792,N_12973,N_12571);
nor U13793 (N_13793,N_12310,N_12944);
nand U13794 (N_13794,N_12354,N_12128);
or U13795 (N_13795,N_12798,N_12491);
nor U13796 (N_13796,N_12912,N_12990);
xnor U13797 (N_13797,N_12980,N_12179);
and U13798 (N_13798,N_12503,N_12214);
or U13799 (N_13799,N_12466,N_12701);
nor U13800 (N_13800,N_12188,N_12662);
nor U13801 (N_13801,N_12305,N_12162);
nand U13802 (N_13802,N_12671,N_12268);
nand U13803 (N_13803,N_12692,N_12641);
xor U13804 (N_13804,N_12771,N_12053);
nand U13805 (N_13805,N_12548,N_12631);
nand U13806 (N_13806,N_12767,N_12579);
nand U13807 (N_13807,N_12543,N_12109);
nor U13808 (N_13808,N_12156,N_12140);
nand U13809 (N_13809,N_12833,N_12595);
nand U13810 (N_13810,N_12542,N_12839);
xnor U13811 (N_13811,N_12332,N_12575);
nor U13812 (N_13812,N_12886,N_12760);
xor U13813 (N_13813,N_12119,N_12714);
nand U13814 (N_13814,N_12683,N_12476);
nand U13815 (N_13815,N_12252,N_12770);
or U13816 (N_13816,N_12531,N_12638);
nand U13817 (N_13817,N_12700,N_12062);
xnor U13818 (N_13818,N_12500,N_12631);
and U13819 (N_13819,N_12855,N_12452);
or U13820 (N_13820,N_12100,N_12726);
xnor U13821 (N_13821,N_12122,N_12510);
or U13822 (N_13822,N_12720,N_12153);
or U13823 (N_13823,N_12403,N_12500);
and U13824 (N_13824,N_12130,N_12062);
nor U13825 (N_13825,N_12250,N_12148);
xor U13826 (N_13826,N_12343,N_12108);
nand U13827 (N_13827,N_12862,N_12505);
nor U13828 (N_13828,N_12879,N_12023);
and U13829 (N_13829,N_12692,N_12826);
or U13830 (N_13830,N_12380,N_12644);
nor U13831 (N_13831,N_12166,N_12993);
nor U13832 (N_13832,N_12876,N_12545);
or U13833 (N_13833,N_12400,N_12813);
nor U13834 (N_13834,N_12149,N_12437);
or U13835 (N_13835,N_12218,N_12441);
nor U13836 (N_13836,N_12402,N_12671);
nor U13837 (N_13837,N_12641,N_12934);
nor U13838 (N_13838,N_12199,N_12002);
nand U13839 (N_13839,N_12513,N_12164);
and U13840 (N_13840,N_12179,N_12194);
nand U13841 (N_13841,N_12066,N_12973);
nor U13842 (N_13842,N_12505,N_12155);
nor U13843 (N_13843,N_12526,N_12146);
xor U13844 (N_13844,N_12333,N_12624);
and U13845 (N_13845,N_12999,N_12976);
nor U13846 (N_13846,N_12545,N_12629);
nor U13847 (N_13847,N_12803,N_12587);
nand U13848 (N_13848,N_12509,N_12216);
and U13849 (N_13849,N_12411,N_12406);
xnor U13850 (N_13850,N_12288,N_12790);
xor U13851 (N_13851,N_12660,N_12947);
xnor U13852 (N_13852,N_12488,N_12178);
nand U13853 (N_13853,N_12273,N_12999);
xor U13854 (N_13854,N_12933,N_12330);
nor U13855 (N_13855,N_12505,N_12906);
xor U13856 (N_13856,N_12288,N_12156);
or U13857 (N_13857,N_12316,N_12108);
nand U13858 (N_13858,N_12204,N_12148);
xnor U13859 (N_13859,N_12911,N_12640);
xor U13860 (N_13860,N_12131,N_12154);
and U13861 (N_13861,N_12013,N_12577);
nor U13862 (N_13862,N_12440,N_12025);
xor U13863 (N_13863,N_12856,N_12158);
nand U13864 (N_13864,N_12987,N_12803);
nor U13865 (N_13865,N_12062,N_12020);
nor U13866 (N_13866,N_12114,N_12249);
xor U13867 (N_13867,N_12316,N_12277);
xor U13868 (N_13868,N_12192,N_12580);
or U13869 (N_13869,N_12093,N_12266);
nor U13870 (N_13870,N_12503,N_12545);
and U13871 (N_13871,N_12915,N_12278);
or U13872 (N_13872,N_12761,N_12919);
or U13873 (N_13873,N_12840,N_12043);
and U13874 (N_13874,N_12405,N_12618);
and U13875 (N_13875,N_12970,N_12858);
xor U13876 (N_13876,N_12186,N_12244);
xnor U13877 (N_13877,N_12937,N_12944);
and U13878 (N_13878,N_12062,N_12041);
nand U13879 (N_13879,N_12707,N_12510);
xnor U13880 (N_13880,N_12873,N_12772);
xnor U13881 (N_13881,N_12793,N_12193);
nand U13882 (N_13882,N_12999,N_12675);
nand U13883 (N_13883,N_12836,N_12231);
nand U13884 (N_13884,N_12934,N_12485);
nor U13885 (N_13885,N_12069,N_12583);
xor U13886 (N_13886,N_12983,N_12807);
nand U13887 (N_13887,N_12844,N_12811);
nor U13888 (N_13888,N_12720,N_12469);
or U13889 (N_13889,N_12925,N_12469);
xnor U13890 (N_13890,N_12501,N_12999);
nor U13891 (N_13891,N_12976,N_12021);
nand U13892 (N_13892,N_12339,N_12604);
and U13893 (N_13893,N_12576,N_12991);
nor U13894 (N_13894,N_12541,N_12404);
xnor U13895 (N_13895,N_12591,N_12075);
or U13896 (N_13896,N_12250,N_12872);
or U13897 (N_13897,N_12729,N_12649);
nand U13898 (N_13898,N_12435,N_12145);
and U13899 (N_13899,N_12941,N_12082);
xnor U13900 (N_13900,N_12456,N_12173);
and U13901 (N_13901,N_12119,N_12365);
or U13902 (N_13902,N_12419,N_12364);
xor U13903 (N_13903,N_12872,N_12246);
xor U13904 (N_13904,N_12575,N_12473);
nand U13905 (N_13905,N_12413,N_12526);
nand U13906 (N_13906,N_12772,N_12516);
xor U13907 (N_13907,N_12023,N_12339);
xor U13908 (N_13908,N_12765,N_12729);
or U13909 (N_13909,N_12720,N_12458);
nand U13910 (N_13910,N_12907,N_12110);
xnor U13911 (N_13911,N_12906,N_12562);
nand U13912 (N_13912,N_12343,N_12205);
xor U13913 (N_13913,N_12380,N_12393);
nand U13914 (N_13914,N_12769,N_12139);
nand U13915 (N_13915,N_12353,N_12138);
or U13916 (N_13916,N_12454,N_12800);
nand U13917 (N_13917,N_12390,N_12117);
or U13918 (N_13918,N_12904,N_12482);
nand U13919 (N_13919,N_12262,N_12960);
and U13920 (N_13920,N_12567,N_12692);
nand U13921 (N_13921,N_12603,N_12665);
or U13922 (N_13922,N_12722,N_12916);
and U13923 (N_13923,N_12182,N_12972);
or U13924 (N_13924,N_12195,N_12064);
nor U13925 (N_13925,N_12120,N_12984);
nor U13926 (N_13926,N_12861,N_12529);
nor U13927 (N_13927,N_12826,N_12698);
or U13928 (N_13928,N_12623,N_12780);
or U13929 (N_13929,N_12251,N_12586);
or U13930 (N_13930,N_12826,N_12262);
nand U13931 (N_13931,N_12198,N_12338);
nor U13932 (N_13932,N_12745,N_12985);
nand U13933 (N_13933,N_12848,N_12888);
or U13934 (N_13934,N_12888,N_12974);
nor U13935 (N_13935,N_12194,N_12009);
nand U13936 (N_13936,N_12220,N_12535);
and U13937 (N_13937,N_12476,N_12617);
xor U13938 (N_13938,N_12929,N_12217);
xor U13939 (N_13939,N_12777,N_12455);
nor U13940 (N_13940,N_12259,N_12716);
and U13941 (N_13941,N_12406,N_12581);
nand U13942 (N_13942,N_12045,N_12337);
nor U13943 (N_13943,N_12855,N_12250);
xor U13944 (N_13944,N_12660,N_12274);
nand U13945 (N_13945,N_12690,N_12046);
nor U13946 (N_13946,N_12170,N_12197);
or U13947 (N_13947,N_12367,N_12525);
and U13948 (N_13948,N_12534,N_12528);
or U13949 (N_13949,N_12433,N_12319);
and U13950 (N_13950,N_12082,N_12569);
nor U13951 (N_13951,N_12789,N_12682);
or U13952 (N_13952,N_12655,N_12964);
nand U13953 (N_13953,N_12596,N_12083);
nor U13954 (N_13954,N_12423,N_12114);
nor U13955 (N_13955,N_12015,N_12418);
nand U13956 (N_13956,N_12251,N_12434);
or U13957 (N_13957,N_12114,N_12725);
nor U13958 (N_13958,N_12328,N_12159);
and U13959 (N_13959,N_12004,N_12803);
nand U13960 (N_13960,N_12934,N_12353);
or U13961 (N_13961,N_12757,N_12941);
nor U13962 (N_13962,N_12889,N_12153);
and U13963 (N_13963,N_12974,N_12432);
xor U13964 (N_13964,N_12015,N_12319);
or U13965 (N_13965,N_12595,N_12113);
or U13966 (N_13966,N_12934,N_12600);
nand U13967 (N_13967,N_12474,N_12595);
nor U13968 (N_13968,N_12840,N_12755);
nor U13969 (N_13969,N_12422,N_12584);
nor U13970 (N_13970,N_12316,N_12305);
nor U13971 (N_13971,N_12445,N_12476);
or U13972 (N_13972,N_12303,N_12178);
xor U13973 (N_13973,N_12413,N_12778);
and U13974 (N_13974,N_12360,N_12991);
nor U13975 (N_13975,N_12307,N_12835);
and U13976 (N_13976,N_12710,N_12515);
xnor U13977 (N_13977,N_12916,N_12817);
nand U13978 (N_13978,N_12904,N_12748);
and U13979 (N_13979,N_12688,N_12268);
xnor U13980 (N_13980,N_12612,N_12641);
xnor U13981 (N_13981,N_12807,N_12131);
nor U13982 (N_13982,N_12287,N_12481);
and U13983 (N_13983,N_12787,N_12608);
xnor U13984 (N_13984,N_12156,N_12603);
nor U13985 (N_13985,N_12960,N_12202);
or U13986 (N_13986,N_12938,N_12649);
nand U13987 (N_13987,N_12862,N_12853);
nand U13988 (N_13988,N_12308,N_12363);
nand U13989 (N_13989,N_12599,N_12043);
nor U13990 (N_13990,N_12252,N_12079);
nor U13991 (N_13991,N_12223,N_12570);
or U13992 (N_13992,N_12950,N_12629);
and U13993 (N_13993,N_12046,N_12197);
nand U13994 (N_13994,N_12182,N_12212);
or U13995 (N_13995,N_12790,N_12799);
xnor U13996 (N_13996,N_12067,N_12241);
and U13997 (N_13997,N_12756,N_12554);
nand U13998 (N_13998,N_12975,N_12161);
nor U13999 (N_13999,N_12449,N_12100);
nand U14000 (N_14000,N_13517,N_13488);
nor U14001 (N_14001,N_13796,N_13417);
nand U14002 (N_14002,N_13861,N_13318);
nand U14003 (N_14003,N_13584,N_13332);
or U14004 (N_14004,N_13817,N_13610);
nand U14005 (N_14005,N_13745,N_13108);
and U14006 (N_14006,N_13766,N_13605);
nor U14007 (N_14007,N_13740,N_13991);
xnor U14008 (N_14008,N_13241,N_13525);
xor U14009 (N_14009,N_13988,N_13915);
and U14010 (N_14010,N_13254,N_13477);
and U14011 (N_14011,N_13048,N_13487);
and U14012 (N_14012,N_13963,N_13157);
xnor U14013 (N_14013,N_13039,N_13322);
and U14014 (N_14014,N_13936,N_13507);
or U14015 (N_14015,N_13981,N_13557);
and U14016 (N_14016,N_13177,N_13218);
nor U14017 (N_14017,N_13765,N_13213);
or U14018 (N_14018,N_13606,N_13815);
nor U14019 (N_14019,N_13669,N_13364);
nand U14020 (N_14020,N_13207,N_13801);
and U14021 (N_14021,N_13732,N_13920);
nand U14022 (N_14022,N_13104,N_13046);
nor U14023 (N_14023,N_13937,N_13164);
or U14024 (N_14024,N_13283,N_13800);
or U14025 (N_14025,N_13356,N_13686);
and U14026 (N_14026,N_13090,N_13343);
xor U14027 (N_14027,N_13200,N_13390);
or U14028 (N_14028,N_13060,N_13857);
nand U14029 (N_14029,N_13638,N_13186);
or U14030 (N_14030,N_13134,N_13107);
nor U14031 (N_14031,N_13274,N_13148);
nand U14032 (N_14032,N_13968,N_13337);
nand U14033 (N_14033,N_13158,N_13953);
nand U14034 (N_14034,N_13418,N_13630);
xor U14035 (N_14035,N_13054,N_13231);
or U14036 (N_14036,N_13537,N_13259);
or U14037 (N_14037,N_13497,N_13811);
xnor U14038 (N_14038,N_13550,N_13139);
nor U14039 (N_14039,N_13929,N_13722);
nor U14040 (N_14040,N_13210,N_13211);
xnor U14041 (N_14041,N_13633,N_13637);
or U14042 (N_14042,N_13085,N_13402);
or U14043 (N_14043,N_13240,N_13451);
xor U14044 (N_14044,N_13744,N_13273);
or U14045 (N_14045,N_13945,N_13999);
xor U14046 (N_14046,N_13018,N_13421);
or U14047 (N_14047,N_13217,N_13681);
and U14048 (N_14048,N_13966,N_13944);
nor U14049 (N_14049,N_13508,N_13179);
or U14050 (N_14050,N_13738,N_13142);
or U14051 (N_14051,N_13827,N_13196);
and U14052 (N_14052,N_13041,N_13710);
nor U14053 (N_14053,N_13394,N_13878);
and U14054 (N_14054,N_13871,N_13472);
and U14055 (N_14055,N_13187,N_13619);
nor U14056 (N_14056,N_13068,N_13327);
nand U14057 (N_14057,N_13132,N_13007);
and U14058 (N_14058,N_13830,N_13917);
xor U14059 (N_14059,N_13540,N_13400);
and U14060 (N_14060,N_13268,N_13987);
or U14061 (N_14061,N_13737,N_13731);
nor U14062 (N_14062,N_13263,N_13292);
nor U14063 (N_14063,N_13168,N_13795);
nor U14064 (N_14064,N_13647,N_13006);
and U14065 (N_14065,N_13693,N_13617);
or U14066 (N_14066,N_13869,N_13973);
xnor U14067 (N_14067,N_13499,N_13797);
xnor U14068 (N_14068,N_13805,N_13038);
nor U14069 (N_14069,N_13350,N_13432);
nand U14070 (N_14070,N_13596,N_13547);
or U14071 (N_14071,N_13354,N_13089);
or U14072 (N_14072,N_13904,N_13896);
nand U14073 (N_14073,N_13045,N_13082);
and U14074 (N_14074,N_13239,N_13062);
xor U14075 (N_14075,N_13438,N_13076);
nand U14076 (N_14076,N_13881,N_13473);
or U14077 (N_14077,N_13790,N_13339);
nor U14078 (N_14078,N_13246,N_13176);
nand U14079 (N_14079,N_13307,N_13956);
nand U14080 (N_14080,N_13426,N_13910);
or U14081 (N_14081,N_13951,N_13348);
and U14082 (N_14082,N_13236,N_13750);
and U14083 (N_14083,N_13919,N_13483);
or U14084 (N_14084,N_13078,N_13761);
or U14085 (N_14085,N_13194,N_13133);
or U14086 (N_14086,N_13478,N_13809);
and U14087 (N_14087,N_13719,N_13066);
or U14088 (N_14088,N_13304,N_13892);
nor U14089 (N_14089,N_13430,N_13276);
nand U14090 (N_14090,N_13579,N_13397);
and U14091 (N_14091,N_13728,N_13627);
nor U14092 (N_14092,N_13636,N_13126);
nand U14093 (N_14093,N_13026,N_13425);
and U14094 (N_14094,N_13688,N_13536);
nor U14095 (N_14095,N_13969,N_13293);
nor U14096 (N_14096,N_13852,N_13415);
or U14097 (N_14097,N_13564,N_13401);
and U14098 (N_14098,N_13768,N_13846);
nand U14099 (N_14099,N_13460,N_13812);
xor U14100 (N_14100,N_13371,N_13326);
nand U14101 (N_14101,N_13344,N_13664);
nor U14102 (N_14102,N_13144,N_13001);
xor U14103 (N_14103,N_13319,N_13404);
nand U14104 (N_14104,N_13206,N_13845);
xor U14105 (N_14105,N_13154,N_13734);
nand U14106 (N_14106,N_13823,N_13975);
or U14107 (N_14107,N_13109,N_13816);
or U14108 (N_14108,N_13569,N_13195);
and U14109 (N_14109,N_13172,N_13129);
nor U14110 (N_14110,N_13600,N_13872);
or U14111 (N_14111,N_13250,N_13361);
xor U14112 (N_14112,N_13625,N_13986);
or U14113 (N_14113,N_13767,N_13080);
and U14114 (N_14114,N_13465,N_13160);
xor U14115 (N_14115,N_13870,N_13383);
xnor U14116 (N_14116,N_13296,N_13754);
and U14117 (N_14117,N_13671,N_13924);
nor U14118 (N_14118,N_13373,N_13009);
and U14119 (N_14119,N_13709,N_13251);
and U14120 (N_14120,N_13716,N_13201);
or U14121 (N_14121,N_13715,N_13258);
nor U14122 (N_14122,N_13372,N_13175);
xnor U14123 (N_14123,N_13940,N_13559);
xnor U14124 (N_14124,N_13684,N_13786);
or U14125 (N_14125,N_13042,N_13355);
nor U14126 (N_14126,N_13612,N_13112);
or U14127 (N_14127,N_13762,N_13453);
or U14128 (N_14128,N_13285,N_13099);
and U14129 (N_14129,N_13959,N_13656);
nand U14130 (N_14130,N_13165,N_13952);
and U14131 (N_14131,N_13900,N_13860);
nor U14132 (N_14132,N_13444,N_13531);
or U14133 (N_14133,N_13275,N_13521);
nand U14134 (N_14134,N_13778,N_13242);
and U14135 (N_14135,N_13237,N_13169);
or U14136 (N_14136,N_13848,N_13065);
nor U14137 (N_14137,N_13663,N_13391);
nand U14138 (N_14138,N_13862,N_13808);
and U14139 (N_14139,N_13253,N_13198);
and U14140 (N_14140,N_13225,N_13149);
or U14141 (N_14141,N_13458,N_13594);
xor U14142 (N_14142,N_13689,N_13262);
nor U14143 (N_14143,N_13926,N_13931);
nand U14144 (N_14144,N_13083,N_13711);
or U14145 (N_14145,N_13943,N_13230);
or U14146 (N_14146,N_13985,N_13590);
nor U14147 (N_14147,N_13069,N_13049);
nand U14148 (N_14148,N_13529,N_13632);
xnor U14149 (N_14149,N_13958,N_13416);
xnor U14150 (N_14150,N_13515,N_13884);
xor U14151 (N_14151,N_13749,N_13270);
and U14152 (N_14152,N_13840,N_13803);
and U14153 (N_14153,N_13530,N_13983);
nand U14154 (N_14154,N_13466,N_13730);
nand U14155 (N_14155,N_13011,N_13675);
and U14156 (N_14156,N_13249,N_13777);
or U14157 (N_14157,N_13297,N_13310);
nor U14158 (N_14158,N_13654,N_13668);
nor U14159 (N_14159,N_13305,N_13114);
nand U14160 (N_14160,N_13101,N_13498);
xor U14161 (N_14161,N_13694,N_13272);
nor U14162 (N_14162,N_13159,N_13843);
or U14163 (N_14163,N_13311,N_13947);
nor U14164 (N_14164,N_13490,N_13533);
and U14165 (N_14165,N_13889,N_13696);
and U14166 (N_14166,N_13941,N_13500);
nor U14167 (N_14167,N_13994,N_13867);
xnor U14168 (N_14168,N_13829,N_13933);
or U14169 (N_14169,N_13202,N_13204);
and U14170 (N_14170,N_13482,N_13072);
nand U14171 (N_14171,N_13029,N_13491);
and U14172 (N_14172,N_13655,N_13161);
and U14173 (N_14173,N_13492,N_13174);
nor U14174 (N_14174,N_13727,N_13651);
xor U14175 (N_14175,N_13597,N_13171);
and U14176 (N_14176,N_13428,N_13601);
nor U14177 (N_14177,N_13431,N_13146);
or U14178 (N_14178,N_13087,N_13548);
xor U14179 (N_14179,N_13789,N_13347);
xnor U14180 (N_14180,N_13020,N_13094);
xnor U14181 (N_14181,N_13967,N_13756);
or U14182 (N_14182,N_13743,N_13475);
and U14183 (N_14183,N_13476,N_13692);
xor U14184 (N_14184,N_13395,N_13023);
and U14185 (N_14185,N_13027,N_13055);
or U14186 (N_14186,N_13102,N_13073);
and U14187 (N_14187,N_13015,N_13648);
nand U14188 (N_14188,N_13128,N_13123);
nor U14189 (N_14189,N_13323,N_13595);
nand U14190 (N_14190,N_13199,N_13984);
and U14191 (N_14191,N_13092,N_13505);
and U14192 (N_14192,N_13303,N_13593);
nand U14193 (N_14193,N_13289,N_13571);
or U14194 (N_14194,N_13459,N_13717);
nand U14195 (N_14195,N_13989,N_13676);
nand U14196 (N_14196,N_13858,N_13407);
xnor U14197 (N_14197,N_13036,N_13863);
nand U14198 (N_14198,N_13839,N_13316);
and U14199 (N_14199,N_13378,N_13427);
or U14200 (N_14200,N_13532,N_13554);
nand U14201 (N_14201,N_13935,N_13524);
nand U14202 (N_14202,N_13440,N_13971);
or U14203 (N_14203,N_13267,N_13489);
nor U14204 (N_14204,N_13992,N_13481);
nand U14205 (N_14205,N_13888,N_13124);
nor U14206 (N_14206,N_13622,N_13646);
and U14207 (N_14207,N_13660,N_13582);
or U14208 (N_14208,N_13847,N_13434);
nor U14209 (N_14209,N_13518,N_13188);
and U14210 (N_14210,N_13556,N_13064);
nand U14211 (N_14211,N_13704,N_13178);
nand U14212 (N_14212,N_13053,N_13785);
and U14213 (N_14213,N_13818,N_13781);
nor U14214 (N_14214,N_13315,N_13714);
or U14215 (N_14215,N_13257,N_13443);
xor U14216 (N_14216,N_13506,N_13494);
nor U14217 (N_14217,N_13927,N_13626);
and U14218 (N_14218,N_13718,N_13948);
xor U14219 (N_14219,N_13306,N_13567);
nor U14220 (N_14220,N_13770,N_13993);
xnor U14221 (N_14221,N_13370,N_13151);
nand U14222 (N_14222,N_13115,N_13442);
xnor U14223 (N_14223,N_13977,N_13523);
or U14224 (N_14224,N_13607,N_13613);
nor U14225 (N_14225,N_13726,N_13031);
or U14226 (N_14226,N_13914,N_13855);
nor U14227 (N_14227,N_13539,N_13598);
and U14228 (N_14228,N_13520,N_13368);
or U14229 (N_14229,N_13287,N_13030);
and U14230 (N_14230,N_13396,N_13534);
or U14231 (N_14231,N_13552,N_13098);
or U14232 (N_14232,N_13934,N_13995);
nand U14233 (N_14233,N_13649,N_13388);
xor U14234 (N_14234,N_13976,N_13997);
xor U14235 (N_14235,N_13615,N_13215);
nand U14236 (N_14236,N_13851,N_13614);
nor U14237 (N_14237,N_13553,N_13208);
and U14238 (N_14238,N_13185,N_13980);
or U14239 (N_14239,N_13224,N_13105);
and U14240 (N_14240,N_13116,N_13399);
xor U14241 (N_14241,N_13873,N_13844);
nand U14242 (N_14242,N_13897,N_13527);
nor U14243 (N_14243,N_13244,N_13712);
or U14244 (N_14244,N_13117,N_13592);
nor U14245 (N_14245,N_13783,N_13110);
nand U14246 (N_14246,N_13288,N_13555);
and U14247 (N_14247,N_13333,N_13903);
xor U14248 (N_14248,N_13760,N_13435);
nor U14249 (N_14249,N_13468,N_13377);
nand U14250 (N_14250,N_13358,N_13086);
or U14251 (N_14251,N_13752,N_13414);
and U14252 (N_14252,N_13720,N_13705);
xor U14253 (N_14253,N_13932,N_13898);
nand U14254 (N_14254,N_13227,N_13279);
xnor U14255 (N_14255,N_13155,N_13764);
and U14256 (N_14256,N_13683,N_13209);
or U14257 (N_14257,N_13173,N_13365);
or U14258 (N_14258,N_13005,N_13708);
and U14259 (N_14259,N_13526,N_13782);
nor U14260 (N_14260,N_13513,N_13831);
and U14261 (N_14261,N_13286,N_13616);
and U14262 (N_14262,N_13381,N_13403);
nand U14263 (N_14263,N_13561,N_13189);
xor U14264 (N_14264,N_13666,N_13100);
xnor U14265 (N_14265,N_13122,N_13970);
nor U14266 (N_14266,N_13658,N_13551);
nand U14267 (N_14267,N_13880,N_13152);
nand U14268 (N_14268,N_13854,N_13044);
or U14269 (N_14269,N_13150,N_13918);
and U14270 (N_14270,N_13883,N_13982);
and U14271 (N_14271,N_13012,N_13603);
nand U14272 (N_14272,N_13228,N_13670);
and U14273 (N_14273,N_13573,N_13560);
nand U14274 (N_14274,N_13939,N_13226);
or U14275 (N_14275,N_13794,N_13634);
nor U14276 (N_14276,N_13819,N_13216);
nor U14277 (N_14277,N_13212,N_13265);
or U14278 (N_14278,N_13890,N_13004);
and U14279 (N_14279,N_13504,N_13480);
xnor U14280 (N_14280,N_13759,N_13035);
or U14281 (N_14281,N_13763,N_13295);
and U14282 (N_14282,N_13037,N_13448);
nor U14283 (N_14283,N_13423,N_13868);
nand U14284 (N_14284,N_13894,N_13735);
xor U14285 (N_14285,N_13130,N_13503);
and U14286 (N_14286,N_13659,N_13446);
or U14287 (N_14287,N_13071,N_13779);
xor U14288 (N_14288,N_13853,N_13229);
nor U14289 (N_14289,N_13184,N_13366);
and U14290 (N_14290,N_13865,N_13181);
xnor U14291 (N_14291,N_13682,N_13901);
nor U14292 (N_14292,N_13909,N_13758);
xor U14293 (N_14293,N_13757,N_13799);
nor U14294 (N_14294,N_13885,N_13163);
xor U14295 (N_14295,N_13138,N_13784);
and U14296 (N_14296,N_13392,N_13429);
or U14297 (N_14297,N_13516,N_13197);
and U14298 (N_14298,N_13575,N_13538);
xnor U14299 (N_14299,N_13424,N_13056);
nand U14300 (N_14300,N_13641,N_13457);
nand U14301 (N_14301,N_13450,N_13814);
and U14302 (N_14302,N_13103,N_13893);
nor U14303 (N_14303,N_13070,N_13447);
xnor U14304 (N_14304,N_13271,N_13183);
xor U14305 (N_14305,N_13385,N_13156);
or U14306 (N_14306,N_13462,N_13528);
and U14307 (N_14307,N_13535,N_13923);
nor U14308 (N_14308,N_13807,N_13906);
and U14309 (N_14309,N_13203,N_13746);
xnor U14310 (N_14310,N_13410,N_13233);
and U14311 (N_14311,N_13574,N_13875);
nand U14312 (N_14312,N_13955,N_13628);
nand U14313 (N_14313,N_13850,N_13733);
and U14314 (N_14314,N_13581,N_13096);
or U14315 (N_14315,N_13695,N_13960);
xnor U14316 (N_14316,N_13609,N_13838);
nor U14317 (N_14317,N_13769,N_13585);
xnor U14318 (N_14318,N_13346,N_13887);
xnor U14319 (N_14319,N_13842,N_13170);
nand U14320 (N_14320,N_13820,N_13191);
nand U14321 (N_14321,N_13753,N_13841);
nor U14322 (N_14322,N_13057,N_13541);
nand U14323 (N_14323,N_13245,N_13962);
nor U14324 (N_14324,N_13008,N_13379);
nor U14325 (N_14325,N_13479,N_13545);
or U14326 (N_14326,N_13620,N_13136);
and U14327 (N_14327,N_13180,N_13234);
nand U14328 (N_14328,N_13357,N_13652);
nand U14329 (N_14329,N_13690,N_13665);
nor U14330 (N_14330,N_13905,N_13238);
or U14331 (N_14331,N_13514,N_13748);
nor U14332 (N_14332,N_13806,N_13353);
nor U14333 (N_14333,N_13672,N_13511);
nor U14334 (N_14334,N_13166,N_13463);
and U14335 (N_14335,N_13436,N_13602);
nor U14336 (N_14336,N_13393,N_13662);
xnor U14337 (N_14337,N_13911,N_13813);
xor U14338 (N_14338,N_13485,N_13502);
nand U14339 (N_14339,N_13467,N_13565);
nor U14340 (N_14340,N_13836,N_13495);
nand U14341 (N_14341,N_13580,N_13650);
or U14342 (N_14342,N_13736,N_13291);
or U14343 (N_14343,N_13810,N_13837);
nor U14344 (N_14344,N_13780,N_13512);
nor U14345 (N_14345,N_13328,N_13141);
xor U14346 (N_14346,N_13120,N_13624);
and U14347 (N_14347,N_13260,N_13859);
nand U14348 (N_14348,N_13111,N_13644);
nor U14349 (N_14349,N_13389,N_13701);
nor U14350 (N_14350,N_13050,N_13243);
or U14351 (N_14351,N_13773,N_13376);
nand U14352 (N_14352,N_13232,N_13412);
or U14353 (N_14353,N_13657,N_13127);
and U14354 (N_14354,N_13978,N_13587);
nand U14355 (N_14355,N_13570,N_13509);
nor U14356 (N_14356,N_13061,N_13033);
nor U14357 (N_14357,N_13010,N_13891);
nor U14358 (N_14358,N_13380,N_13879);
nor U14359 (N_14359,N_13949,N_13420);
nor U14360 (N_14360,N_13828,N_13546);
xnor U14361 (N_14361,N_13703,N_13063);
nor U14362 (N_14362,N_13367,N_13864);
and U14363 (N_14363,N_13729,N_13342);
or U14364 (N_14364,N_13996,N_13298);
nand U14365 (N_14365,N_13938,N_13586);
nor U14366 (N_14366,N_13334,N_13774);
and U14367 (N_14367,N_13034,N_13549);
and U14368 (N_14368,N_13832,N_13351);
or U14369 (N_14369,N_13882,N_13019);
or U14370 (N_14370,N_13685,N_13793);
nor U14371 (N_14371,N_13899,N_13916);
xor U14372 (N_14372,N_13566,N_13739);
xor U14373 (N_14373,N_13025,N_13974);
and U14374 (N_14374,N_13013,N_13252);
xnor U14375 (N_14375,N_13051,N_13247);
or U14376 (N_14376,N_13902,N_13331);
nor U14377 (N_14377,N_13886,N_13329);
or U14378 (N_14378,N_13445,N_13776);
xnor U14379 (N_14379,N_13470,N_13621);
and U14380 (N_14380,N_13058,N_13699);
and U14381 (N_14381,N_13577,N_13093);
and U14382 (N_14382,N_13826,N_13591);
and U14383 (N_14383,N_13433,N_13677);
or U14384 (N_14384,N_13091,N_13576);
nand U14385 (N_14385,N_13455,N_13266);
nor U14386 (N_14386,N_13639,N_13314);
nand U14387 (N_14387,N_13725,N_13235);
or U14388 (N_14388,N_13014,N_13798);
and U14389 (N_14389,N_13702,N_13723);
nand U14390 (N_14390,N_13834,N_13028);
or U14391 (N_14391,N_13017,N_13021);
nor U14392 (N_14392,N_13849,N_13484);
nor U14393 (N_14393,N_13653,N_13772);
and U14394 (N_14394,N_13280,N_13137);
nor U14395 (N_14395,N_13922,N_13724);
nand U14396 (N_14396,N_13349,N_13308);
nand U14397 (N_14397,N_13317,N_13707);
or U14398 (N_14398,N_13833,N_13441);
and U14399 (N_14399,N_13192,N_13925);
nand U14400 (N_14400,N_13409,N_13118);
nand U14401 (N_14401,N_13145,N_13930);
nor U14402 (N_14402,N_13856,N_13340);
xnor U14403 (N_14403,N_13697,N_13352);
nor U14404 (N_14404,N_13519,N_13698);
xor U14405 (N_14405,N_13335,N_13294);
and U14406 (N_14406,N_13946,N_13113);
or U14407 (N_14407,N_13928,N_13153);
or U14408 (N_14408,N_13486,N_13721);
xor U14409 (N_14409,N_13631,N_13713);
and U14410 (N_14410,N_13067,N_13387);
and U14411 (N_14411,N_13121,N_13755);
or U14412 (N_14412,N_13449,N_13398);
nor U14413 (N_14413,N_13075,N_13821);
nand U14414 (N_14414,N_13369,N_13588);
nor U14415 (N_14415,N_13277,N_13452);
nor U14416 (N_14416,N_13706,N_13413);
nand U14417 (N_14417,N_13804,N_13341);
and U14418 (N_14418,N_13255,N_13824);
or U14419 (N_14419,N_13119,N_13321);
xor U14420 (N_14420,N_13543,N_13406);
nor U14421 (N_14421,N_13261,N_13284);
xnor U14422 (N_14422,N_13667,N_13921);
and U14423 (N_14423,N_13700,N_13678);
or U14424 (N_14424,N_13248,N_13791);
nor U14425 (N_14425,N_13635,N_13077);
or U14426 (N_14426,N_13787,N_13162);
nor U14427 (N_14427,N_13691,N_13979);
xor U14428 (N_14428,N_13362,N_13493);
xnor U14429 (N_14429,N_13474,N_13792);
and U14430 (N_14430,N_13751,N_13583);
and U14431 (N_14431,N_13623,N_13360);
xnor U14432 (N_14432,N_13572,N_13679);
xnor U14433 (N_14433,N_13312,N_13954);
nor U14434 (N_14434,N_13106,N_13471);
or U14435 (N_14435,N_13167,N_13558);
xnor U14436 (N_14436,N_13950,N_13408);
and U14437 (N_14437,N_13264,N_13419);
or U14438 (N_14438,N_13325,N_13866);
or U14439 (N_14439,N_13299,N_13363);
nand U14440 (N_14440,N_13300,N_13895);
or U14441 (N_14441,N_13510,N_13741);
nand U14442 (N_14442,N_13147,N_13496);
or U14443 (N_14443,N_13747,N_13088);
or U14444 (N_14444,N_13282,N_13775);
nand U14445 (N_14445,N_13016,N_13190);
nor U14446 (N_14446,N_13411,N_13439);
and U14447 (N_14447,N_13674,N_13278);
xnor U14448 (N_14448,N_13220,N_13022);
nand U14449 (N_14449,N_13320,N_13386);
nand U14450 (N_14450,N_13290,N_13788);
nand U14451 (N_14451,N_13135,N_13269);
xnor U14452 (N_14452,N_13374,N_13084);
xnor U14453 (N_14453,N_13422,N_13384);
nor U14454 (N_14454,N_13382,N_13822);
and U14455 (N_14455,N_13223,N_13079);
or U14456 (N_14456,N_13052,N_13456);
nor U14457 (N_14457,N_13578,N_13522);
nand U14458 (N_14458,N_13043,N_13964);
nand U14459 (N_14459,N_13661,N_13125);
or U14460 (N_14460,N_13256,N_13542);
and U14461 (N_14461,N_13907,N_13338);
and U14462 (N_14462,N_13059,N_13501);
nor U14463 (N_14463,N_13643,N_13074);
nor U14464 (N_14464,N_13437,N_13345);
xor U14465 (N_14465,N_13568,N_13330);
nand U14466 (N_14466,N_13742,N_13143);
nand U14467 (N_14467,N_13281,N_13942);
or U14468 (N_14468,N_13040,N_13182);
xnor U14469 (N_14469,N_13642,N_13874);
and U14470 (N_14470,N_13095,N_13544);
nand U14471 (N_14471,N_13002,N_13618);
nor U14472 (N_14472,N_13313,N_13645);
nor U14473 (N_14473,N_13464,N_13219);
nand U14474 (N_14474,N_13990,N_13908);
xnor U14475 (N_14475,N_13205,N_13608);
xor U14476 (N_14476,N_13214,N_13131);
and U14477 (N_14477,N_13000,N_13825);
nand U14478 (N_14478,N_13302,N_13405);
or U14479 (N_14479,N_13221,N_13877);
or U14480 (N_14480,N_13562,N_13913);
and U14481 (N_14481,N_13097,N_13336);
or U14482 (N_14482,N_13301,N_13309);
or U14483 (N_14483,N_13461,N_13375);
nor U14484 (N_14484,N_13998,N_13563);
and U14485 (N_14485,N_13222,N_13469);
nand U14486 (N_14486,N_13640,N_13673);
nor U14487 (N_14487,N_13081,N_13835);
xor U14488 (N_14488,N_13599,N_13359);
and U14489 (N_14489,N_13003,N_13589);
nand U14490 (N_14490,N_13047,N_13629);
nor U14491 (N_14491,N_13611,N_13032);
nor U14492 (N_14492,N_13957,N_13802);
xnor U14493 (N_14493,N_13972,N_13771);
nand U14494 (N_14494,N_13193,N_13912);
and U14495 (N_14495,N_13961,N_13024);
xnor U14496 (N_14496,N_13140,N_13324);
xnor U14497 (N_14497,N_13965,N_13876);
and U14498 (N_14498,N_13680,N_13454);
nor U14499 (N_14499,N_13604,N_13687);
and U14500 (N_14500,N_13226,N_13478);
nand U14501 (N_14501,N_13943,N_13227);
nand U14502 (N_14502,N_13217,N_13078);
nand U14503 (N_14503,N_13376,N_13213);
and U14504 (N_14504,N_13040,N_13967);
xor U14505 (N_14505,N_13226,N_13534);
and U14506 (N_14506,N_13135,N_13374);
nand U14507 (N_14507,N_13779,N_13092);
nand U14508 (N_14508,N_13754,N_13377);
nor U14509 (N_14509,N_13669,N_13448);
nor U14510 (N_14510,N_13182,N_13234);
xor U14511 (N_14511,N_13330,N_13609);
and U14512 (N_14512,N_13617,N_13185);
nor U14513 (N_14513,N_13033,N_13193);
nor U14514 (N_14514,N_13887,N_13974);
and U14515 (N_14515,N_13469,N_13094);
nor U14516 (N_14516,N_13352,N_13180);
nand U14517 (N_14517,N_13227,N_13125);
nand U14518 (N_14518,N_13698,N_13347);
xor U14519 (N_14519,N_13687,N_13262);
nand U14520 (N_14520,N_13736,N_13036);
or U14521 (N_14521,N_13394,N_13259);
nor U14522 (N_14522,N_13232,N_13944);
nand U14523 (N_14523,N_13381,N_13499);
and U14524 (N_14524,N_13957,N_13287);
nor U14525 (N_14525,N_13258,N_13288);
nor U14526 (N_14526,N_13902,N_13645);
nand U14527 (N_14527,N_13046,N_13371);
nor U14528 (N_14528,N_13618,N_13398);
xnor U14529 (N_14529,N_13756,N_13440);
xnor U14530 (N_14530,N_13429,N_13391);
xnor U14531 (N_14531,N_13285,N_13168);
and U14532 (N_14532,N_13874,N_13996);
xor U14533 (N_14533,N_13725,N_13710);
xor U14534 (N_14534,N_13151,N_13107);
xor U14535 (N_14535,N_13923,N_13672);
nand U14536 (N_14536,N_13006,N_13349);
nor U14537 (N_14537,N_13469,N_13921);
or U14538 (N_14538,N_13306,N_13618);
and U14539 (N_14539,N_13689,N_13068);
nor U14540 (N_14540,N_13651,N_13511);
or U14541 (N_14541,N_13408,N_13865);
and U14542 (N_14542,N_13459,N_13868);
xor U14543 (N_14543,N_13521,N_13544);
nand U14544 (N_14544,N_13594,N_13722);
and U14545 (N_14545,N_13758,N_13858);
xnor U14546 (N_14546,N_13102,N_13020);
xor U14547 (N_14547,N_13362,N_13824);
or U14548 (N_14548,N_13656,N_13294);
nand U14549 (N_14549,N_13630,N_13032);
nor U14550 (N_14550,N_13222,N_13427);
and U14551 (N_14551,N_13247,N_13112);
nand U14552 (N_14552,N_13654,N_13170);
nor U14553 (N_14553,N_13818,N_13847);
nand U14554 (N_14554,N_13159,N_13809);
nor U14555 (N_14555,N_13794,N_13467);
and U14556 (N_14556,N_13959,N_13339);
xor U14557 (N_14557,N_13122,N_13327);
nand U14558 (N_14558,N_13955,N_13806);
nand U14559 (N_14559,N_13390,N_13722);
or U14560 (N_14560,N_13937,N_13463);
and U14561 (N_14561,N_13465,N_13386);
xor U14562 (N_14562,N_13506,N_13437);
or U14563 (N_14563,N_13769,N_13661);
nor U14564 (N_14564,N_13944,N_13719);
xnor U14565 (N_14565,N_13340,N_13153);
or U14566 (N_14566,N_13520,N_13104);
nand U14567 (N_14567,N_13449,N_13118);
xnor U14568 (N_14568,N_13303,N_13505);
or U14569 (N_14569,N_13454,N_13796);
and U14570 (N_14570,N_13389,N_13487);
nor U14571 (N_14571,N_13138,N_13441);
or U14572 (N_14572,N_13398,N_13996);
and U14573 (N_14573,N_13767,N_13444);
nand U14574 (N_14574,N_13277,N_13043);
nor U14575 (N_14575,N_13268,N_13823);
nor U14576 (N_14576,N_13003,N_13253);
nand U14577 (N_14577,N_13946,N_13468);
nand U14578 (N_14578,N_13924,N_13950);
xnor U14579 (N_14579,N_13562,N_13112);
xor U14580 (N_14580,N_13144,N_13708);
xor U14581 (N_14581,N_13898,N_13366);
nand U14582 (N_14582,N_13702,N_13405);
nor U14583 (N_14583,N_13479,N_13264);
xnor U14584 (N_14584,N_13455,N_13508);
nor U14585 (N_14585,N_13244,N_13157);
and U14586 (N_14586,N_13708,N_13608);
or U14587 (N_14587,N_13732,N_13803);
or U14588 (N_14588,N_13995,N_13110);
xor U14589 (N_14589,N_13400,N_13002);
xor U14590 (N_14590,N_13591,N_13463);
nand U14591 (N_14591,N_13990,N_13381);
nor U14592 (N_14592,N_13756,N_13306);
nand U14593 (N_14593,N_13661,N_13876);
or U14594 (N_14594,N_13526,N_13296);
nor U14595 (N_14595,N_13042,N_13979);
or U14596 (N_14596,N_13605,N_13745);
or U14597 (N_14597,N_13067,N_13328);
and U14598 (N_14598,N_13600,N_13998);
nand U14599 (N_14599,N_13719,N_13279);
nand U14600 (N_14600,N_13263,N_13852);
nand U14601 (N_14601,N_13370,N_13607);
and U14602 (N_14602,N_13976,N_13387);
nand U14603 (N_14603,N_13552,N_13916);
and U14604 (N_14604,N_13807,N_13077);
and U14605 (N_14605,N_13774,N_13591);
or U14606 (N_14606,N_13081,N_13797);
and U14607 (N_14607,N_13003,N_13646);
or U14608 (N_14608,N_13767,N_13449);
nor U14609 (N_14609,N_13270,N_13230);
and U14610 (N_14610,N_13705,N_13160);
or U14611 (N_14611,N_13386,N_13406);
xnor U14612 (N_14612,N_13385,N_13304);
or U14613 (N_14613,N_13941,N_13319);
and U14614 (N_14614,N_13595,N_13173);
nand U14615 (N_14615,N_13151,N_13275);
or U14616 (N_14616,N_13358,N_13453);
nor U14617 (N_14617,N_13921,N_13557);
or U14618 (N_14618,N_13291,N_13336);
xor U14619 (N_14619,N_13685,N_13989);
nor U14620 (N_14620,N_13869,N_13574);
xnor U14621 (N_14621,N_13108,N_13067);
or U14622 (N_14622,N_13969,N_13820);
xor U14623 (N_14623,N_13054,N_13603);
nor U14624 (N_14624,N_13675,N_13296);
nor U14625 (N_14625,N_13516,N_13298);
xnor U14626 (N_14626,N_13661,N_13849);
and U14627 (N_14627,N_13326,N_13886);
or U14628 (N_14628,N_13411,N_13720);
or U14629 (N_14629,N_13468,N_13891);
nand U14630 (N_14630,N_13060,N_13904);
nand U14631 (N_14631,N_13780,N_13112);
and U14632 (N_14632,N_13465,N_13657);
or U14633 (N_14633,N_13963,N_13131);
and U14634 (N_14634,N_13281,N_13543);
nand U14635 (N_14635,N_13339,N_13659);
and U14636 (N_14636,N_13999,N_13014);
nand U14637 (N_14637,N_13756,N_13664);
or U14638 (N_14638,N_13570,N_13406);
nor U14639 (N_14639,N_13139,N_13008);
and U14640 (N_14640,N_13805,N_13971);
or U14641 (N_14641,N_13908,N_13844);
nor U14642 (N_14642,N_13868,N_13871);
nor U14643 (N_14643,N_13840,N_13449);
nor U14644 (N_14644,N_13684,N_13101);
nor U14645 (N_14645,N_13359,N_13373);
or U14646 (N_14646,N_13367,N_13852);
or U14647 (N_14647,N_13138,N_13658);
or U14648 (N_14648,N_13919,N_13697);
xor U14649 (N_14649,N_13800,N_13928);
nand U14650 (N_14650,N_13431,N_13384);
and U14651 (N_14651,N_13204,N_13793);
nor U14652 (N_14652,N_13123,N_13986);
and U14653 (N_14653,N_13481,N_13996);
nand U14654 (N_14654,N_13198,N_13603);
nand U14655 (N_14655,N_13185,N_13739);
xor U14656 (N_14656,N_13824,N_13878);
nand U14657 (N_14657,N_13940,N_13781);
xor U14658 (N_14658,N_13114,N_13864);
nand U14659 (N_14659,N_13406,N_13498);
nand U14660 (N_14660,N_13495,N_13253);
nand U14661 (N_14661,N_13591,N_13646);
nor U14662 (N_14662,N_13930,N_13178);
or U14663 (N_14663,N_13797,N_13719);
nor U14664 (N_14664,N_13109,N_13888);
nor U14665 (N_14665,N_13077,N_13057);
nor U14666 (N_14666,N_13947,N_13643);
nor U14667 (N_14667,N_13005,N_13581);
xnor U14668 (N_14668,N_13029,N_13539);
nand U14669 (N_14669,N_13884,N_13487);
xnor U14670 (N_14670,N_13012,N_13091);
nor U14671 (N_14671,N_13295,N_13944);
nor U14672 (N_14672,N_13068,N_13727);
nor U14673 (N_14673,N_13022,N_13331);
or U14674 (N_14674,N_13619,N_13307);
nor U14675 (N_14675,N_13740,N_13427);
and U14676 (N_14676,N_13952,N_13459);
and U14677 (N_14677,N_13304,N_13227);
or U14678 (N_14678,N_13506,N_13479);
nor U14679 (N_14679,N_13309,N_13876);
or U14680 (N_14680,N_13904,N_13753);
nand U14681 (N_14681,N_13427,N_13781);
nor U14682 (N_14682,N_13086,N_13291);
nand U14683 (N_14683,N_13052,N_13926);
or U14684 (N_14684,N_13722,N_13699);
nand U14685 (N_14685,N_13999,N_13490);
nor U14686 (N_14686,N_13959,N_13401);
nor U14687 (N_14687,N_13829,N_13107);
nor U14688 (N_14688,N_13899,N_13150);
xor U14689 (N_14689,N_13943,N_13761);
nand U14690 (N_14690,N_13147,N_13230);
and U14691 (N_14691,N_13409,N_13096);
nor U14692 (N_14692,N_13517,N_13316);
or U14693 (N_14693,N_13648,N_13598);
and U14694 (N_14694,N_13724,N_13497);
nand U14695 (N_14695,N_13998,N_13412);
xnor U14696 (N_14696,N_13829,N_13088);
nor U14697 (N_14697,N_13162,N_13791);
nor U14698 (N_14698,N_13141,N_13018);
nor U14699 (N_14699,N_13684,N_13196);
or U14700 (N_14700,N_13137,N_13695);
or U14701 (N_14701,N_13520,N_13158);
xor U14702 (N_14702,N_13552,N_13139);
nor U14703 (N_14703,N_13660,N_13865);
xnor U14704 (N_14704,N_13142,N_13950);
xor U14705 (N_14705,N_13308,N_13671);
nor U14706 (N_14706,N_13242,N_13000);
nand U14707 (N_14707,N_13120,N_13440);
nor U14708 (N_14708,N_13705,N_13908);
and U14709 (N_14709,N_13364,N_13125);
xor U14710 (N_14710,N_13025,N_13456);
xnor U14711 (N_14711,N_13923,N_13083);
and U14712 (N_14712,N_13316,N_13222);
and U14713 (N_14713,N_13099,N_13368);
xor U14714 (N_14714,N_13140,N_13730);
xnor U14715 (N_14715,N_13688,N_13475);
nand U14716 (N_14716,N_13032,N_13564);
nand U14717 (N_14717,N_13849,N_13171);
xor U14718 (N_14718,N_13423,N_13397);
nor U14719 (N_14719,N_13666,N_13944);
xor U14720 (N_14720,N_13557,N_13844);
nand U14721 (N_14721,N_13549,N_13764);
nand U14722 (N_14722,N_13298,N_13737);
nand U14723 (N_14723,N_13857,N_13670);
or U14724 (N_14724,N_13782,N_13975);
xor U14725 (N_14725,N_13938,N_13365);
nand U14726 (N_14726,N_13851,N_13887);
nor U14727 (N_14727,N_13342,N_13870);
nand U14728 (N_14728,N_13205,N_13699);
and U14729 (N_14729,N_13513,N_13997);
or U14730 (N_14730,N_13109,N_13490);
or U14731 (N_14731,N_13384,N_13906);
nand U14732 (N_14732,N_13121,N_13569);
xor U14733 (N_14733,N_13772,N_13999);
nor U14734 (N_14734,N_13289,N_13531);
nor U14735 (N_14735,N_13074,N_13385);
nor U14736 (N_14736,N_13867,N_13232);
or U14737 (N_14737,N_13911,N_13694);
or U14738 (N_14738,N_13422,N_13467);
and U14739 (N_14739,N_13773,N_13813);
and U14740 (N_14740,N_13304,N_13823);
nor U14741 (N_14741,N_13840,N_13981);
or U14742 (N_14742,N_13854,N_13572);
or U14743 (N_14743,N_13219,N_13559);
xor U14744 (N_14744,N_13328,N_13834);
and U14745 (N_14745,N_13612,N_13332);
nand U14746 (N_14746,N_13431,N_13833);
or U14747 (N_14747,N_13373,N_13030);
xnor U14748 (N_14748,N_13453,N_13802);
or U14749 (N_14749,N_13406,N_13109);
and U14750 (N_14750,N_13338,N_13127);
or U14751 (N_14751,N_13354,N_13978);
nor U14752 (N_14752,N_13400,N_13061);
nor U14753 (N_14753,N_13086,N_13614);
nand U14754 (N_14754,N_13616,N_13533);
xnor U14755 (N_14755,N_13324,N_13207);
or U14756 (N_14756,N_13193,N_13895);
or U14757 (N_14757,N_13287,N_13552);
xor U14758 (N_14758,N_13498,N_13040);
nor U14759 (N_14759,N_13211,N_13498);
nand U14760 (N_14760,N_13723,N_13603);
and U14761 (N_14761,N_13470,N_13912);
nand U14762 (N_14762,N_13805,N_13250);
and U14763 (N_14763,N_13474,N_13418);
nor U14764 (N_14764,N_13210,N_13893);
xor U14765 (N_14765,N_13323,N_13871);
nor U14766 (N_14766,N_13279,N_13570);
xor U14767 (N_14767,N_13705,N_13599);
nand U14768 (N_14768,N_13964,N_13156);
nor U14769 (N_14769,N_13462,N_13400);
nor U14770 (N_14770,N_13281,N_13548);
nor U14771 (N_14771,N_13119,N_13426);
or U14772 (N_14772,N_13953,N_13884);
nor U14773 (N_14773,N_13009,N_13878);
or U14774 (N_14774,N_13351,N_13348);
and U14775 (N_14775,N_13415,N_13835);
xnor U14776 (N_14776,N_13125,N_13425);
nor U14777 (N_14777,N_13761,N_13400);
nand U14778 (N_14778,N_13431,N_13516);
nor U14779 (N_14779,N_13805,N_13856);
xnor U14780 (N_14780,N_13080,N_13232);
and U14781 (N_14781,N_13647,N_13030);
nand U14782 (N_14782,N_13799,N_13040);
or U14783 (N_14783,N_13878,N_13649);
and U14784 (N_14784,N_13983,N_13842);
or U14785 (N_14785,N_13449,N_13784);
nand U14786 (N_14786,N_13018,N_13612);
and U14787 (N_14787,N_13404,N_13548);
nor U14788 (N_14788,N_13479,N_13016);
xor U14789 (N_14789,N_13139,N_13874);
nand U14790 (N_14790,N_13409,N_13288);
nand U14791 (N_14791,N_13679,N_13464);
or U14792 (N_14792,N_13818,N_13589);
or U14793 (N_14793,N_13956,N_13125);
and U14794 (N_14794,N_13083,N_13109);
xor U14795 (N_14795,N_13456,N_13840);
and U14796 (N_14796,N_13406,N_13499);
nand U14797 (N_14797,N_13686,N_13108);
nand U14798 (N_14798,N_13520,N_13186);
or U14799 (N_14799,N_13436,N_13006);
or U14800 (N_14800,N_13832,N_13149);
or U14801 (N_14801,N_13387,N_13047);
nand U14802 (N_14802,N_13910,N_13030);
nand U14803 (N_14803,N_13356,N_13134);
nand U14804 (N_14804,N_13392,N_13342);
or U14805 (N_14805,N_13657,N_13680);
or U14806 (N_14806,N_13618,N_13334);
xnor U14807 (N_14807,N_13975,N_13143);
and U14808 (N_14808,N_13760,N_13527);
or U14809 (N_14809,N_13720,N_13195);
nand U14810 (N_14810,N_13456,N_13983);
and U14811 (N_14811,N_13197,N_13609);
nand U14812 (N_14812,N_13139,N_13328);
and U14813 (N_14813,N_13344,N_13383);
xor U14814 (N_14814,N_13064,N_13420);
or U14815 (N_14815,N_13546,N_13951);
xnor U14816 (N_14816,N_13791,N_13157);
nor U14817 (N_14817,N_13654,N_13028);
xnor U14818 (N_14818,N_13154,N_13122);
and U14819 (N_14819,N_13779,N_13083);
nand U14820 (N_14820,N_13664,N_13244);
or U14821 (N_14821,N_13156,N_13327);
nand U14822 (N_14822,N_13522,N_13975);
nand U14823 (N_14823,N_13527,N_13999);
xor U14824 (N_14824,N_13115,N_13273);
nand U14825 (N_14825,N_13466,N_13361);
or U14826 (N_14826,N_13165,N_13683);
nor U14827 (N_14827,N_13664,N_13054);
and U14828 (N_14828,N_13776,N_13828);
nand U14829 (N_14829,N_13587,N_13280);
nand U14830 (N_14830,N_13484,N_13810);
nor U14831 (N_14831,N_13326,N_13081);
nand U14832 (N_14832,N_13499,N_13562);
xor U14833 (N_14833,N_13695,N_13405);
or U14834 (N_14834,N_13124,N_13061);
xor U14835 (N_14835,N_13541,N_13431);
nand U14836 (N_14836,N_13146,N_13914);
or U14837 (N_14837,N_13496,N_13852);
nor U14838 (N_14838,N_13434,N_13909);
and U14839 (N_14839,N_13263,N_13889);
xnor U14840 (N_14840,N_13719,N_13711);
xor U14841 (N_14841,N_13550,N_13006);
nor U14842 (N_14842,N_13185,N_13652);
nand U14843 (N_14843,N_13121,N_13187);
xor U14844 (N_14844,N_13297,N_13044);
nand U14845 (N_14845,N_13622,N_13874);
nand U14846 (N_14846,N_13884,N_13875);
xnor U14847 (N_14847,N_13352,N_13177);
nor U14848 (N_14848,N_13300,N_13981);
or U14849 (N_14849,N_13414,N_13956);
nand U14850 (N_14850,N_13595,N_13138);
xnor U14851 (N_14851,N_13475,N_13289);
xor U14852 (N_14852,N_13748,N_13520);
nand U14853 (N_14853,N_13955,N_13726);
nand U14854 (N_14854,N_13970,N_13855);
or U14855 (N_14855,N_13851,N_13403);
or U14856 (N_14856,N_13555,N_13050);
nor U14857 (N_14857,N_13734,N_13239);
or U14858 (N_14858,N_13456,N_13690);
xor U14859 (N_14859,N_13058,N_13978);
nand U14860 (N_14860,N_13658,N_13347);
xnor U14861 (N_14861,N_13672,N_13237);
nand U14862 (N_14862,N_13521,N_13752);
nor U14863 (N_14863,N_13808,N_13286);
nand U14864 (N_14864,N_13015,N_13026);
nor U14865 (N_14865,N_13205,N_13297);
and U14866 (N_14866,N_13459,N_13797);
nor U14867 (N_14867,N_13232,N_13183);
xor U14868 (N_14868,N_13976,N_13356);
and U14869 (N_14869,N_13357,N_13774);
xnor U14870 (N_14870,N_13355,N_13026);
xnor U14871 (N_14871,N_13039,N_13238);
xor U14872 (N_14872,N_13942,N_13844);
and U14873 (N_14873,N_13087,N_13370);
nand U14874 (N_14874,N_13890,N_13449);
or U14875 (N_14875,N_13226,N_13715);
xnor U14876 (N_14876,N_13641,N_13290);
nand U14877 (N_14877,N_13492,N_13763);
and U14878 (N_14878,N_13028,N_13591);
xor U14879 (N_14879,N_13914,N_13805);
nor U14880 (N_14880,N_13534,N_13030);
nand U14881 (N_14881,N_13451,N_13061);
and U14882 (N_14882,N_13502,N_13175);
and U14883 (N_14883,N_13613,N_13616);
and U14884 (N_14884,N_13443,N_13267);
nand U14885 (N_14885,N_13648,N_13081);
or U14886 (N_14886,N_13258,N_13704);
nand U14887 (N_14887,N_13432,N_13800);
and U14888 (N_14888,N_13914,N_13575);
nor U14889 (N_14889,N_13594,N_13692);
xnor U14890 (N_14890,N_13497,N_13113);
and U14891 (N_14891,N_13154,N_13836);
and U14892 (N_14892,N_13994,N_13220);
and U14893 (N_14893,N_13925,N_13022);
nor U14894 (N_14894,N_13126,N_13817);
or U14895 (N_14895,N_13966,N_13393);
nor U14896 (N_14896,N_13943,N_13115);
or U14897 (N_14897,N_13440,N_13364);
or U14898 (N_14898,N_13796,N_13721);
nand U14899 (N_14899,N_13474,N_13832);
or U14900 (N_14900,N_13247,N_13651);
nand U14901 (N_14901,N_13274,N_13466);
or U14902 (N_14902,N_13220,N_13562);
or U14903 (N_14903,N_13683,N_13192);
nand U14904 (N_14904,N_13318,N_13949);
xor U14905 (N_14905,N_13865,N_13387);
nand U14906 (N_14906,N_13657,N_13330);
nor U14907 (N_14907,N_13250,N_13972);
or U14908 (N_14908,N_13110,N_13621);
nor U14909 (N_14909,N_13791,N_13086);
and U14910 (N_14910,N_13272,N_13050);
and U14911 (N_14911,N_13953,N_13271);
nor U14912 (N_14912,N_13981,N_13075);
and U14913 (N_14913,N_13271,N_13388);
nand U14914 (N_14914,N_13159,N_13509);
xnor U14915 (N_14915,N_13124,N_13164);
nand U14916 (N_14916,N_13275,N_13536);
nand U14917 (N_14917,N_13427,N_13805);
nor U14918 (N_14918,N_13307,N_13634);
and U14919 (N_14919,N_13921,N_13078);
nor U14920 (N_14920,N_13801,N_13673);
and U14921 (N_14921,N_13009,N_13789);
and U14922 (N_14922,N_13850,N_13139);
xnor U14923 (N_14923,N_13791,N_13610);
nand U14924 (N_14924,N_13290,N_13551);
nand U14925 (N_14925,N_13351,N_13982);
and U14926 (N_14926,N_13708,N_13716);
and U14927 (N_14927,N_13189,N_13862);
nor U14928 (N_14928,N_13349,N_13488);
xor U14929 (N_14929,N_13837,N_13289);
nor U14930 (N_14930,N_13098,N_13258);
and U14931 (N_14931,N_13238,N_13195);
and U14932 (N_14932,N_13524,N_13050);
nand U14933 (N_14933,N_13082,N_13254);
nand U14934 (N_14934,N_13799,N_13696);
xor U14935 (N_14935,N_13874,N_13160);
nor U14936 (N_14936,N_13552,N_13320);
nor U14937 (N_14937,N_13296,N_13678);
xnor U14938 (N_14938,N_13696,N_13422);
nand U14939 (N_14939,N_13111,N_13611);
or U14940 (N_14940,N_13801,N_13754);
and U14941 (N_14941,N_13304,N_13389);
xor U14942 (N_14942,N_13332,N_13222);
and U14943 (N_14943,N_13658,N_13651);
nand U14944 (N_14944,N_13452,N_13766);
nor U14945 (N_14945,N_13841,N_13347);
or U14946 (N_14946,N_13429,N_13641);
and U14947 (N_14947,N_13457,N_13885);
xor U14948 (N_14948,N_13604,N_13574);
and U14949 (N_14949,N_13350,N_13006);
nand U14950 (N_14950,N_13081,N_13465);
nand U14951 (N_14951,N_13766,N_13884);
nand U14952 (N_14952,N_13512,N_13807);
xnor U14953 (N_14953,N_13954,N_13401);
nor U14954 (N_14954,N_13116,N_13086);
xnor U14955 (N_14955,N_13314,N_13132);
and U14956 (N_14956,N_13135,N_13739);
nor U14957 (N_14957,N_13175,N_13926);
and U14958 (N_14958,N_13405,N_13950);
and U14959 (N_14959,N_13506,N_13052);
nand U14960 (N_14960,N_13997,N_13473);
or U14961 (N_14961,N_13554,N_13019);
xnor U14962 (N_14962,N_13745,N_13602);
nand U14963 (N_14963,N_13063,N_13510);
or U14964 (N_14964,N_13140,N_13887);
and U14965 (N_14965,N_13726,N_13262);
nand U14966 (N_14966,N_13068,N_13546);
nor U14967 (N_14967,N_13929,N_13174);
nand U14968 (N_14968,N_13630,N_13676);
nand U14969 (N_14969,N_13077,N_13285);
nand U14970 (N_14970,N_13031,N_13316);
or U14971 (N_14971,N_13253,N_13531);
nand U14972 (N_14972,N_13907,N_13366);
nor U14973 (N_14973,N_13510,N_13654);
or U14974 (N_14974,N_13381,N_13019);
and U14975 (N_14975,N_13976,N_13223);
or U14976 (N_14976,N_13166,N_13789);
nor U14977 (N_14977,N_13220,N_13047);
nor U14978 (N_14978,N_13096,N_13639);
and U14979 (N_14979,N_13971,N_13661);
or U14980 (N_14980,N_13402,N_13230);
or U14981 (N_14981,N_13873,N_13723);
and U14982 (N_14982,N_13030,N_13541);
xnor U14983 (N_14983,N_13842,N_13068);
xor U14984 (N_14984,N_13275,N_13424);
nand U14985 (N_14985,N_13286,N_13010);
xor U14986 (N_14986,N_13056,N_13537);
and U14987 (N_14987,N_13133,N_13564);
and U14988 (N_14988,N_13492,N_13197);
nand U14989 (N_14989,N_13821,N_13917);
nand U14990 (N_14990,N_13601,N_13215);
xor U14991 (N_14991,N_13175,N_13770);
and U14992 (N_14992,N_13851,N_13304);
or U14993 (N_14993,N_13605,N_13720);
and U14994 (N_14994,N_13023,N_13293);
and U14995 (N_14995,N_13996,N_13031);
nor U14996 (N_14996,N_13065,N_13952);
xnor U14997 (N_14997,N_13851,N_13785);
and U14998 (N_14998,N_13310,N_13143);
and U14999 (N_14999,N_13701,N_13721);
xnor U15000 (N_15000,N_14362,N_14988);
or U15001 (N_15001,N_14299,N_14238);
and U15002 (N_15002,N_14668,N_14703);
nor U15003 (N_15003,N_14459,N_14217);
nor U15004 (N_15004,N_14394,N_14442);
and U15005 (N_15005,N_14283,N_14875);
nor U15006 (N_15006,N_14794,N_14645);
nor U15007 (N_15007,N_14562,N_14034);
and U15008 (N_15008,N_14603,N_14734);
and U15009 (N_15009,N_14173,N_14010);
nand U15010 (N_15010,N_14975,N_14114);
nor U15011 (N_15011,N_14728,N_14111);
and U15012 (N_15012,N_14626,N_14029);
or U15013 (N_15013,N_14666,N_14829);
or U15014 (N_15014,N_14253,N_14190);
nor U15015 (N_15015,N_14554,N_14785);
and U15016 (N_15016,N_14431,N_14862);
nor U15017 (N_15017,N_14510,N_14376);
or U15018 (N_15018,N_14701,N_14230);
or U15019 (N_15019,N_14255,N_14392);
nand U15020 (N_15020,N_14891,N_14019);
and U15021 (N_15021,N_14078,N_14552);
nand U15022 (N_15022,N_14973,N_14610);
and U15023 (N_15023,N_14321,N_14850);
nand U15024 (N_15024,N_14699,N_14854);
nor U15025 (N_15025,N_14744,N_14476);
nand U15026 (N_15026,N_14528,N_14056);
and U15027 (N_15027,N_14006,N_14592);
nor U15028 (N_15028,N_14488,N_14355);
nor U15029 (N_15029,N_14767,N_14204);
or U15030 (N_15030,N_14531,N_14159);
or U15031 (N_15031,N_14541,N_14009);
nand U15032 (N_15032,N_14134,N_14293);
and U15033 (N_15033,N_14414,N_14315);
nand U15034 (N_15034,N_14583,N_14643);
xnor U15035 (N_15035,N_14187,N_14466);
xnor U15036 (N_15036,N_14967,N_14309);
xnor U15037 (N_15037,N_14537,N_14692);
xnor U15038 (N_15038,N_14427,N_14228);
nand U15039 (N_15039,N_14044,N_14695);
nor U15040 (N_15040,N_14193,N_14251);
nand U15041 (N_15041,N_14989,N_14103);
or U15042 (N_15042,N_14845,N_14132);
xnor U15043 (N_15043,N_14383,N_14840);
and U15044 (N_15044,N_14941,N_14005);
nor U15045 (N_15045,N_14121,N_14564);
or U15046 (N_15046,N_14671,N_14385);
or U15047 (N_15047,N_14259,N_14288);
and U15048 (N_15048,N_14836,N_14659);
or U15049 (N_15049,N_14826,N_14072);
nand U15050 (N_15050,N_14063,N_14742);
and U15051 (N_15051,N_14025,N_14735);
or U15052 (N_15052,N_14130,N_14038);
xor U15053 (N_15053,N_14558,N_14196);
nor U15054 (N_15054,N_14908,N_14194);
and U15055 (N_15055,N_14116,N_14573);
xnor U15056 (N_15056,N_14591,N_14675);
or U15057 (N_15057,N_14968,N_14422);
nor U15058 (N_15058,N_14195,N_14595);
nor U15059 (N_15059,N_14627,N_14687);
or U15060 (N_15060,N_14944,N_14706);
nand U15061 (N_15061,N_14389,N_14420);
nand U15062 (N_15062,N_14504,N_14873);
nand U15063 (N_15063,N_14447,N_14171);
or U15064 (N_15064,N_14921,N_14086);
nor U15065 (N_15065,N_14727,N_14100);
xor U15066 (N_15066,N_14756,N_14681);
or U15067 (N_15067,N_14048,N_14804);
and U15068 (N_15068,N_14249,N_14271);
nor U15069 (N_15069,N_14285,N_14887);
nand U15070 (N_15070,N_14018,N_14081);
nor U15071 (N_15071,N_14698,N_14185);
or U15072 (N_15072,N_14331,N_14515);
nand U15073 (N_15073,N_14502,N_14092);
or U15074 (N_15074,N_14684,N_14205);
xor U15075 (N_15075,N_14563,N_14013);
nand U15076 (N_15076,N_14227,N_14469);
or U15077 (N_15077,N_14015,N_14486);
nand U15078 (N_15078,N_14607,N_14158);
and U15079 (N_15079,N_14278,N_14885);
nor U15080 (N_15080,N_14039,N_14679);
or U15081 (N_15081,N_14032,N_14747);
and U15082 (N_15082,N_14404,N_14074);
and U15083 (N_15083,N_14880,N_14693);
nor U15084 (N_15084,N_14364,N_14323);
xor U15085 (N_15085,N_14677,N_14276);
or U15086 (N_15086,N_14306,N_14200);
nand U15087 (N_15087,N_14586,N_14443);
nand U15088 (N_15088,N_14184,N_14585);
nand U15089 (N_15089,N_14477,N_14865);
nand U15090 (N_15090,N_14341,N_14265);
xnor U15091 (N_15091,N_14898,N_14587);
nor U15092 (N_15092,N_14314,N_14770);
and U15093 (N_15093,N_14395,N_14648);
xnor U15094 (N_15094,N_14683,N_14464);
and U15095 (N_15095,N_14300,N_14805);
nor U15096 (N_15096,N_14042,N_14367);
or U15097 (N_15097,N_14233,N_14399);
or U15098 (N_15098,N_14670,N_14717);
xnor U15099 (N_15099,N_14709,N_14678);
xor U15100 (N_15100,N_14753,N_14872);
and U15101 (N_15101,N_14982,N_14538);
nor U15102 (N_15102,N_14590,N_14716);
or U15103 (N_15103,N_14485,N_14075);
and U15104 (N_15104,N_14738,N_14816);
nand U15105 (N_15105,N_14041,N_14214);
and U15106 (N_15106,N_14183,N_14848);
nor U15107 (N_15107,N_14802,N_14094);
and U15108 (N_15108,N_14417,N_14152);
xnor U15109 (N_15109,N_14370,N_14711);
or U15110 (N_15110,N_14943,N_14601);
nor U15111 (N_15111,N_14575,N_14867);
and U15112 (N_15112,N_14224,N_14823);
xor U15113 (N_15113,N_14962,N_14408);
nor U15114 (N_15114,N_14053,N_14932);
xnor U15115 (N_15115,N_14899,N_14553);
or U15116 (N_15116,N_14773,N_14388);
and U15117 (N_15117,N_14356,N_14297);
nor U15118 (N_15118,N_14234,N_14642);
and U15119 (N_15119,N_14567,N_14938);
nand U15120 (N_15120,N_14326,N_14798);
xnor U15121 (N_15121,N_14764,N_14062);
nor U15122 (N_15122,N_14954,N_14926);
nor U15123 (N_15123,N_14471,N_14030);
xor U15124 (N_15124,N_14223,N_14884);
and U15125 (N_15125,N_14107,N_14965);
xnor U15126 (N_15126,N_14813,N_14570);
or U15127 (N_15127,N_14170,N_14923);
and U15128 (N_15128,N_14858,N_14919);
xnor U15129 (N_15129,N_14952,N_14117);
or U15130 (N_15130,N_14572,N_14368);
and U15131 (N_15131,N_14410,N_14175);
nand U15132 (N_15132,N_14916,N_14128);
xor U15133 (N_15133,N_14914,N_14424);
xnor U15134 (N_15134,N_14058,N_14688);
or U15135 (N_15135,N_14113,N_14741);
and U15136 (N_15136,N_14219,N_14999);
and U15137 (N_15137,N_14256,N_14208);
nand U15138 (N_15138,N_14083,N_14868);
nand U15139 (N_15139,N_14400,N_14992);
nand U15140 (N_15140,N_14363,N_14815);
nor U15141 (N_15141,N_14778,N_14942);
or U15142 (N_15142,N_14977,N_14472);
and U15143 (N_15143,N_14149,N_14518);
or U15144 (N_15144,N_14596,N_14568);
nor U15145 (N_15145,N_14080,N_14661);
or U15146 (N_15146,N_14831,N_14345);
or U15147 (N_15147,N_14604,N_14147);
nand U15148 (N_15148,N_14281,N_14732);
nand U15149 (N_15149,N_14549,N_14165);
and U15150 (N_15150,N_14105,N_14754);
and U15151 (N_15151,N_14937,N_14237);
nand U15152 (N_15152,N_14245,N_14521);
nor U15153 (N_15153,N_14156,N_14386);
or U15154 (N_15154,N_14874,N_14526);
nor U15155 (N_15155,N_14857,N_14956);
or U15156 (N_15156,N_14883,N_14011);
nor U15157 (N_15157,N_14304,N_14786);
xor U15158 (N_15158,N_14972,N_14377);
and U15159 (N_15159,N_14261,N_14307);
or U15160 (N_15160,N_14847,N_14949);
or U15161 (N_15161,N_14310,N_14491);
nor U15162 (N_15162,N_14779,N_14799);
and U15163 (N_15163,N_14057,N_14536);
nand U15164 (N_15164,N_14373,N_14123);
xor U15165 (N_15165,N_14664,N_14654);
or U15166 (N_15166,N_14807,N_14461);
nor U15167 (N_15167,N_14933,N_14843);
or U15168 (N_15168,N_14220,N_14282);
nand U15169 (N_15169,N_14031,N_14320);
nor U15170 (N_15170,N_14723,N_14060);
or U15171 (N_15171,N_14674,N_14354);
nand U15172 (N_15172,N_14247,N_14133);
or U15173 (N_15173,N_14650,N_14012);
and U15174 (N_15174,N_14624,N_14448);
xor U15175 (N_15175,N_14896,N_14639);
nor U15176 (N_15176,N_14559,N_14555);
xnor U15177 (N_15177,N_14752,N_14468);
xnor U15178 (N_15178,N_14296,N_14758);
or U15179 (N_15179,N_14556,N_14174);
nor U15180 (N_15180,N_14361,N_14935);
and U15181 (N_15181,N_14811,N_14188);
nor U15182 (N_15182,N_14069,N_14222);
xnor U15183 (N_15183,N_14384,N_14743);
nor U15184 (N_15184,N_14463,N_14131);
and U15185 (N_15185,N_14917,N_14690);
or U15186 (N_15186,N_14425,N_14871);
xor U15187 (N_15187,N_14886,N_14007);
nand U15188 (N_15188,N_14700,N_14235);
nand U15189 (N_15189,N_14150,N_14109);
xor U15190 (N_15190,N_14474,N_14985);
nand U15191 (N_15191,N_14930,N_14533);
xor U15192 (N_15192,N_14763,N_14325);
and U15193 (N_15193,N_14339,N_14366);
xnor U15194 (N_15194,N_14998,N_14702);
xnor U15195 (N_15195,N_14046,N_14338);
or U15196 (N_15196,N_14279,N_14329);
nand U15197 (N_15197,N_14974,N_14598);
xor U15198 (N_15198,N_14498,N_14519);
nand U15199 (N_15199,N_14250,N_14082);
xor U15200 (N_15200,N_14911,N_14398);
or U15201 (N_15201,N_14569,N_14313);
nand U15202 (N_15202,N_14633,N_14691);
or U15203 (N_15203,N_14792,N_14878);
xnor U15204 (N_15204,N_14050,N_14902);
nand U15205 (N_15205,N_14396,N_14606);
nand U15206 (N_15206,N_14275,N_14202);
or U15207 (N_15207,N_14360,N_14008);
nor U15208 (N_15208,N_14907,N_14835);
or U15209 (N_15209,N_14451,N_14551);
or U15210 (N_15210,N_14856,N_14254);
xnor U15211 (N_15211,N_14168,N_14499);
or U15212 (N_15212,N_14182,N_14178);
and U15213 (N_15213,N_14284,N_14409);
or U15214 (N_15214,N_14163,N_14925);
nand U15215 (N_15215,N_14318,N_14393);
nor U15216 (N_15216,N_14808,N_14415);
xor U15217 (N_15217,N_14543,N_14242);
nor U15218 (N_15218,N_14291,N_14561);
nand U15219 (N_15219,N_14818,N_14017);
nand U15220 (N_15220,N_14506,N_14218);
or U15221 (N_15221,N_14828,N_14849);
and U15222 (N_15222,N_14277,N_14927);
and U15223 (N_15223,N_14176,N_14990);
or U15224 (N_15224,N_14494,N_14788);
nor U15225 (N_15225,N_14101,N_14001);
nor U15226 (N_15226,N_14820,N_14371);
and U15227 (N_15227,N_14768,N_14704);
or U15228 (N_15228,N_14881,N_14548);
nand U15229 (N_15229,N_14997,N_14433);
nor U15230 (N_15230,N_14746,N_14673);
xnor U15231 (N_15231,N_14895,N_14096);
xnor U15232 (N_15232,N_14330,N_14416);
nand U15233 (N_15233,N_14979,N_14324);
nand U15234 (N_15234,N_14232,N_14267);
xor U15235 (N_15235,N_14522,N_14390);
or U15236 (N_15236,N_14359,N_14656);
nor U15237 (N_15237,N_14003,N_14336);
xnor U15238 (N_15238,N_14516,N_14729);
and U15239 (N_15239,N_14697,N_14832);
or U15240 (N_15240,N_14369,N_14231);
nor U15241 (N_15241,N_14544,N_14508);
xor U15242 (N_15242,N_14397,N_14614);
xor U15243 (N_15243,N_14333,N_14167);
and U15244 (N_15244,N_14827,N_14920);
xor U15245 (N_15245,N_14120,N_14014);
nand U15246 (N_15246,N_14102,N_14118);
or U15247 (N_15247,N_14897,N_14566);
or U15248 (N_15248,N_14622,N_14458);
nor U15249 (N_15249,N_14412,N_14207);
nand U15250 (N_15250,N_14745,N_14421);
nor U15251 (N_15251,N_14093,N_14311);
xor U15252 (N_15252,N_14725,N_14157);
nand U15253 (N_15253,N_14966,N_14817);
or U15254 (N_15254,N_14636,N_14059);
nand U15255 (N_15255,N_14164,N_14721);
xnor U15256 (N_15256,N_14560,N_14667);
or U15257 (N_15257,N_14467,N_14658);
nand U15258 (N_15258,N_14091,N_14915);
xnor U15259 (N_15259,N_14489,N_14730);
xnor U15260 (N_15260,N_14672,N_14085);
and U15261 (N_15261,N_14576,N_14335);
xnor U15262 (N_15262,N_14181,N_14445);
nor U15263 (N_15263,N_14625,N_14628);
or U15264 (N_15264,N_14212,N_14160);
nand U15265 (N_15265,N_14210,N_14791);
or U15266 (N_15266,N_14248,N_14750);
xnor U15267 (N_15267,N_14180,N_14351);
nor U15268 (N_15268,N_14122,N_14470);
and U15269 (N_15269,N_14910,N_14795);
or U15270 (N_15270,N_14456,N_14064);
nand U15271 (N_15271,N_14715,N_14473);
and U15272 (N_15272,N_14144,N_14037);
nand U15273 (N_15273,N_14924,N_14381);
or U15274 (N_15274,N_14772,N_14162);
nor U15275 (N_15275,N_14405,N_14177);
nand U15276 (N_15276,N_14620,N_14138);
nor U15277 (N_15277,N_14951,N_14136);
xor U15278 (N_15278,N_14870,N_14580);
xnor U15279 (N_15279,N_14978,N_14146);
and U15280 (N_15280,N_14020,N_14026);
or U15281 (N_15281,N_14760,N_14577);
nand U15282 (N_15282,N_14446,N_14073);
xnor U15283 (N_15283,N_14615,N_14286);
nor U15284 (N_15284,N_14565,N_14452);
and U15285 (N_15285,N_14644,N_14024);
xnor U15286 (N_15286,N_14557,N_14199);
xnor U15287 (N_15287,N_14903,N_14864);
nor U15288 (N_15288,N_14027,N_14500);
nand U15289 (N_15289,N_14501,N_14757);
nand U15290 (N_15290,N_14269,N_14894);
xnor U15291 (N_15291,N_14953,N_14403);
nor U15292 (N_15292,N_14302,N_14525);
nor U15293 (N_15293,N_14514,N_14382);
nand U15294 (N_15294,N_14694,N_14976);
and U15295 (N_15295,N_14948,N_14995);
xor U15296 (N_15296,N_14774,N_14809);
nand U15297 (N_15297,N_14055,N_14344);
and U15298 (N_15298,N_14379,N_14240);
or U15299 (N_15299,N_14407,N_14731);
xor U15300 (N_15300,N_14274,N_14523);
nand U15301 (N_15301,N_14127,N_14819);
or U15302 (N_15302,N_14115,N_14124);
and U15303 (N_15303,N_14428,N_14334);
xor U15304 (N_15304,N_14539,N_14682);
nor U15305 (N_15305,N_14209,N_14104);
nor U15306 (N_15306,N_14509,N_14801);
or U15307 (N_15307,N_14766,N_14143);
nand U15308 (N_15308,N_14308,N_14912);
nand U15309 (N_15309,N_14593,N_14301);
nor U15310 (N_15310,N_14028,N_14655);
nand U15311 (N_15311,N_14071,N_14353);
xnor U15312 (N_15312,N_14800,N_14630);
nor U15313 (N_15313,N_14540,N_14478);
nor U15314 (N_15314,N_14051,N_14243);
xor U15315 (N_15315,N_14833,N_14928);
nor U15316 (N_15316,N_14892,N_14771);
nand U15317 (N_15317,N_14406,N_14787);
xor U15318 (N_15318,N_14838,N_14780);
nor U15319 (N_15319,N_14258,N_14350);
or U15320 (N_15320,N_14714,N_14505);
xor U15321 (N_15321,N_14618,N_14853);
or U15322 (N_15322,N_14969,N_14876);
nand U15323 (N_15323,N_14718,N_14068);
or U15324 (N_15324,N_14264,N_14260);
nor U15325 (N_15325,N_14439,N_14713);
xnor U15326 (N_15326,N_14890,N_14534);
and U15327 (N_15327,N_14939,N_14497);
nand U15328 (N_15328,N_14221,N_14043);
or U15329 (N_15329,N_14348,N_14947);
or U15330 (N_15330,N_14035,N_14426);
nand U15331 (N_15331,N_14273,N_14257);
and U15332 (N_15332,N_14934,N_14226);
xnor U15333 (N_15333,N_14151,N_14166);
nand U15334 (N_15334,N_14987,N_14705);
xor U15335 (N_15335,N_14419,N_14733);
nand U15336 (N_15336,N_14532,N_14783);
or U15337 (N_15337,N_14305,N_14841);
nand U15338 (N_15338,N_14453,N_14651);
nor U15339 (N_15339,N_14652,N_14550);
and U15340 (N_15340,N_14067,N_14112);
and U15341 (N_15341,N_14740,N_14430);
and U15342 (N_15342,N_14429,N_14287);
and U15343 (N_15343,N_14859,N_14378);
xor U15344 (N_15344,N_14803,N_14087);
nand U15345 (N_15345,N_14289,N_14004);
xor U15346 (N_15346,N_14981,N_14137);
or U15347 (N_15347,N_14629,N_14889);
and U15348 (N_15348,N_14996,N_14991);
nand U15349 (N_15349,N_14547,N_14946);
xnor U15350 (N_15350,N_14061,N_14810);
and U15351 (N_15351,N_14413,N_14436);
xnor U15352 (N_15352,N_14929,N_14696);
nor U15353 (N_15353,N_14759,N_14040);
and U15354 (N_15354,N_14686,N_14964);
and U15355 (N_15355,N_14179,N_14844);
nand U15356 (N_15356,N_14796,N_14052);
nand U15357 (N_15357,N_14597,N_14600);
nand U15358 (N_15358,N_14579,N_14877);
xor U15359 (N_15359,N_14342,N_14141);
or U15360 (N_15360,N_14825,N_14280);
nor U15361 (N_15361,N_14663,N_14527);
nand U15362 (N_15362,N_14822,N_14161);
nor U15363 (N_15363,N_14842,N_14680);
or U15364 (N_15364,N_14438,N_14047);
xnor U15365 (N_15365,N_14084,N_14244);
or U15366 (N_15366,N_14971,N_14045);
xor U15367 (N_15367,N_14140,N_14719);
xor U15368 (N_15368,N_14722,N_14483);
or U15369 (N_15369,N_14901,N_14649);
or U15370 (N_15370,N_14119,N_14511);
and U15371 (N_15371,N_14545,N_14814);
or U15372 (N_15372,N_14662,N_14513);
or U15373 (N_15373,N_14189,N_14391);
xor U15374 (N_15374,N_14021,N_14402);
or U15375 (N_15375,N_14099,N_14148);
xor U15376 (N_15376,N_14479,N_14748);
and U15377 (N_15377,N_14154,N_14669);
xnor U15378 (N_15378,N_14879,N_14077);
xor U15379 (N_15379,N_14215,N_14950);
nor U15380 (N_15380,N_14646,N_14749);
nand U15381 (N_15381,N_14186,N_14089);
or U15382 (N_15382,N_14507,N_14712);
nand U15383 (N_15383,N_14142,N_14322);
nand U15384 (N_15384,N_14777,N_14023);
nor U15385 (N_15385,N_14503,N_14098);
nand U15386 (N_15386,N_14905,N_14192);
or U15387 (N_15387,N_14198,N_14262);
nand U15388 (N_15388,N_14380,N_14460);
or U15389 (N_15389,N_14530,N_14613);
nand U15390 (N_15390,N_14839,N_14493);
nand U15391 (N_15391,N_14450,N_14837);
and U15392 (N_15392,N_14793,N_14882);
and U15393 (N_15393,N_14411,N_14432);
nand U15394 (N_15394,N_14957,N_14357);
nand U15395 (N_15395,N_14033,N_14036);
xor U15396 (N_15396,N_14524,N_14270);
nor U15397 (N_15397,N_14726,N_14578);
or U15398 (N_15398,N_14374,N_14108);
and U15399 (N_15399,N_14616,N_14961);
or U15400 (N_15400,N_14487,N_14888);
or U15401 (N_15401,N_14824,N_14863);
nor U15402 (N_15402,N_14789,N_14520);
xor U15403 (N_15403,N_14066,N_14762);
nor U15404 (N_15404,N_14710,N_14812);
and U15405 (N_15405,N_14936,N_14358);
nor U15406 (N_15406,N_14993,N_14172);
nor U15407 (N_15407,N_14866,N_14632);
or U15408 (N_15408,N_14784,N_14638);
nor U15409 (N_15409,N_14834,N_14761);
xnor U15410 (N_15410,N_14090,N_14401);
and U15411 (N_15411,N_14145,N_14736);
nor U15412 (N_15412,N_14455,N_14906);
or U15413 (N_15413,N_14016,N_14332);
xnor U15414 (N_15414,N_14959,N_14292);
nand U15415 (N_15415,N_14387,N_14676);
nor U15416 (N_15416,N_14640,N_14869);
or U15417 (N_15417,N_14197,N_14465);
nand U15418 (N_15418,N_14621,N_14707);
and U15419 (N_15419,N_14481,N_14303);
and U15420 (N_15420,N_14246,N_14855);
nor U15421 (N_15421,N_14135,N_14594);
or U15422 (N_15422,N_14316,N_14211);
and U15423 (N_15423,N_14480,N_14290);
nor U15424 (N_15424,N_14955,N_14529);
and U15425 (N_15425,N_14106,N_14125);
nand U15426 (N_15426,N_14931,N_14647);
and U15427 (N_15427,N_14846,N_14423);
or U15428 (N_15428,N_14317,N_14574);
and U15429 (N_15429,N_14904,N_14375);
or U15430 (N_15430,N_14994,N_14203);
xnor U15431 (N_15431,N_14913,N_14781);
nor U15432 (N_15432,N_14070,N_14437);
xor U15433 (N_15433,N_14191,N_14444);
and U15434 (N_15434,N_14076,N_14054);
and U15435 (N_15435,N_14236,N_14720);
or U15436 (N_15436,N_14724,N_14940);
nor U15437 (N_15437,N_14588,N_14918);
xnor U15438 (N_15438,N_14983,N_14599);
and U15439 (N_15439,N_14657,N_14206);
nor U15440 (N_15440,N_14328,N_14945);
or U15441 (N_15441,N_14272,N_14830);
nand U15442 (N_15442,N_14079,N_14457);
or U15443 (N_15443,N_14213,N_14900);
nor U15444 (N_15444,N_14980,N_14347);
and U15445 (N_15445,N_14637,N_14689);
nor U15446 (N_15446,N_14806,N_14861);
nor U15447 (N_15447,N_14685,N_14095);
nor U15448 (N_15448,N_14986,N_14797);
xor U15449 (N_15449,N_14776,N_14495);
nand U15450 (N_15450,N_14958,N_14435);
xnor U15451 (N_15451,N_14765,N_14263);
xor U15452 (N_15452,N_14860,N_14970);
and U15453 (N_15453,N_14343,N_14852);
or U15454 (N_15454,N_14337,N_14960);
nor U15455 (N_15455,N_14349,N_14110);
nand U15456 (N_15456,N_14441,N_14252);
nand U15457 (N_15457,N_14739,N_14984);
or U15458 (N_15458,N_14665,N_14631);
and U15459 (N_15459,N_14612,N_14660);
nand U15460 (N_15460,N_14582,N_14241);
and U15461 (N_15461,N_14609,N_14963);
or U15462 (N_15462,N_14319,N_14821);
nor U15463 (N_15463,N_14589,N_14295);
and U15464 (N_15464,N_14225,N_14434);
nor U15465 (N_15465,N_14312,N_14049);
xnor U15466 (N_15466,N_14169,N_14619);
and U15467 (N_15467,N_14546,N_14535);
or U15468 (N_15468,N_14893,N_14623);
nand U15469 (N_15469,N_14584,N_14126);
or U15470 (N_15470,N_14449,N_14571);
and U15471 (N_15471,N_14365,N_14216);
nand U15472 (N_15472,N_14229,N_14155);
nor U15473 (N_15473,N_14605,N_14352);
and U15474 (N_15474,N_14484,N_14139);
xor U15475 (N_15475,N_14440,N_14496);
xor U15476 (N_15476,N_14000,N_14088);
nor U15477 (N_15477,N_14708,N_14492);
nor U15478 (N_15478,N_14851,N_14490);
nor U15479 (N_15479,N_14608,N_14346);
xnor U15480 (N_15480,N_14475,N_14298);
and U15481 (N_15481,N_14581,N_14755);
and U15482 (N_15482,N_14641,N_14634);
or U15483 (N_15483,N_14909,N_14617);
or U15484 (N_15484,N_14454,N_14097);
nand U15485 (N_15485,N_14737,N_14653);
and U15486 (N_15486,N_14239,N_14418);
and U15487 (N_15487,N_14153,N_14751);
and U15488 (N_15488,N_14268,N_14002);
xnor U15489 (N_15489,N_14635,N_14482);
nand U15490 (N_15490,N_14340,N_14602);
or U15491 (N_15491,N_14790,N_14782);
and U15492 (N_15492,N_14769,N_14372);
xor U15493 (N_15493,N_14129,N_14065);
or U15494 (N_15494,N_14775,N_14922);
and U15495 (N_15495,N_14266,N_14512);
nor U15496 (N_15496,N_14462,N_14294);
nand U15497 (N_15497,N_14517,N_14327);
nor U15498 (N_15498,N_14201,N_14022);
or U15499 (N_15499,N_14611,N_14542);
nor U15500 (N_15500,N_14401,N_14049);
xor U15501 (N_15501,N_14784,N_14218);
xnor U15502 (N_15502,N_14186,N_14509);
or U15503 (N_15503,N_14304,N_14458);
nand U15504 (N_15504,N_14331,N_14741);
nor U15505 (N_15505,N_14400,N_14293);
or U15506 (N_15506,N_14339,N_14137);
or U15507 (N_15507,N_14883,N_14196);
and U15508 (N_15508,N_14639,N_14241);
nand U15509 (N_15509,N_14271,N_14157);
and U15510 (N_15510,N_14824,N_14182);
or U15511 (N_15511,N_14567,N_14906);
nor U15512 (N_15512,N_14596,N_14645);
xnor U15513 (N_15513,N_14185,N_14581);
or U15514 (N_15514,N_14857,N_14776);
nand U15515 (N_15515,N_14171,N_14255);
nand U15516 (N_15516,N_14632,N_14167);
nand U15517 (N_15517,N_14330,N_14548);
or U15518 (N_15518,N_14097,N_14312);
nor U15519 (N_15519,N_14393,N_14942);
nor U15520 (N_15520,N_14895,N_14989);
nor U15521 (N_15521,N_14606,N_14203);
xnor U15522 (N_15522,N_14727,N_14171);
nand U15523 (N_15523,N_14939,N_14088);
or U15524 (N_15524,N_14331,N_14000);
xor U15525 (N_15525,N_14639,N_14350);
nand U15526 (N_15526,N_14576,N_14067);
and U15527 (N_15527,N_14075,N_14518);
nand U15528 (N_15528,N_14166,N_14548);
and U15529 (N_15529,N_14635,N_14361);
or U15530 (N_15530,N_14790,N_14871);
nor U15531 (N_15531,N_14649,N_14738);
nor U15532 (N_15532,N_14360,N_14065);
nand U15533 (N_15533,N_14794,N_14738);
xor U15534 (N_15534,N_14984,N_14520);
nand U15535 (N_15535,N_14611,N_14660);
xor U15536 (N_15536,N_14624,N_14825);
or U15537 (N_15537,N_14761,N_14843);
or U15538 (N_15538,N_14385,N_14634);
nand U15539 (N_15539,N_14054,N_14469);
and U15540 (N_15540,N_14145,N_14348);
nor U15541 (N_15541,N_14355,N_14872);
and U15542 (N_15542,N_14011,N_14612);
nand U15543 (N_15543,N_14402,N_14777);
or U15544 (N_15544,N_14246,N_14113);
xor U15545 (N_15545,N_14106,N_14481);
nand U15546 (N_15546,N_14346,N_14906);
xnor U15547 (N_15547,N_14309,N_14063);
nor U15548 (N_15548,N_14527,N_14150);
or U15549 (N_15549,N_14518,N_14321);
or U15550 (N_15550,N_14269,N_14213);
xnor U15551 (N_15551,N_14728,N_14717);
or U15552 (N_15552,N_14323,N_14388);
xor U15553 (N_15553,N_14595,N_14504);
and U15554 (N_15554,N_14096,N_14768);
xnor U15555 (N_15555,N_14917,N_14913);
and U15556 (N_15556,N_14325,N_14578);
nand U15557 (N_15557,N_14742,N_14778);
nor U15558 (N_15558,N_14527,N_14472);
nor U15559 (N_15559,N_14234,N_14141);
xor U15560 (N_15560,N_14194,N_14512);
or U15561 (N_15561,N_14054,N_14014);
or U15562 (N_15562,N_14383,N_14813);
nor U15563 (N_15563,N_14432,N_14650);
or U15564 (N_15564,N_14686,N_14928);
or U15565 (N_15565,N_14391,N_14683);
nor U15566 (N_15566,N_14982,N_14229);
xnor U15567 (N_15567,N_14367,N_14261);
xnor U15568 (N_15568,N_14923,N_14740);
or U15569 (N_15569,N_14042,N_14062);
xor U15570 (N_15570,N_14752,N_14687);
nor U15571 (N_15571,N_14956,N_14280);
or U15572 (N_15572,N_14225,N_14852);
and U15573 (N_15573,N_14603,N_14328);
or U15574 (N_15574,N_14442,N_14695);
nand U15575 (N_15575,N_14481,N_14860);
nor U15576 (N_15576,N_14050,N_14957);
or U15577 (N_15577,N_14023,N_14260);
or U15578 (N_15578,N_14153,N_14320);
nor U15579 (N_15579,N_14889,N_14514);
nor U15580 (N_15580,N_14047,N_14437);
nor U15581 (N_15581,N_14739,N_14059);
nor U15582 (N_15582,N_14407,N_14686);
nor U15583 (N_15583,N_14888,N_14001);
nand U15584 (N_15584,N_14709,N_14570);
xnor U15585 (N_15585,N_14443,N_14076);
xor U15586 (N_15586,N_14827,N_14659);
and U15587 (N_15587,N_14798,N_14241);
or U15588 (N_15588,N_14963,N_14562);
or U15589 (N_15589,N_14619,N_14122);
or U15590 (N_15590,N_14065,N_14935);
nand U15591 (N_15591,N_14872,N_14996);
nand U15592 (N_15592,N_14841,N_14827);
nor U15593 (N_15593,N_14373,N_14855);
or U15594 (N_15594,N_14516,N_14937);
nand U15595 (N_15595,N_14749,N_14111);
xnor U15596 (N_15596,N_14367,N_14316);
nand U15597 (N_15597,N_14583,N_14567);
nor U15598 (N_15598,N_14756,N_14271);
xnor U15599 (N_15599,N_14841,N_14186);
or U15600 (N_15600,N_14920,N_14892);
nor U15601 (N_15601,N_14468,N_14378);
nand U15602 (N_15602,N_14335,N_14257);
xnor U15603 (N_15603,N_14092,N_14640);
or U15604 (N_15604,N_14839,N_14953);
nor U15605 (N_15605,N_14737,N_14704);
and U15606 (N_15606,N_14998,N_14693);
nor U15607 (N_15607,N_14132,N_14796);
nand U15608 (N_15608,N_14164,N_14841);
nand U15609 (N_15609,N_14797,N_14246);
and U15610 (N_15610,N_14567,N_14187);
nor U15611 (N_15611,N_14666,N_14131);
xnor U15612 (N_15612,N_14748,N_14155);
nor U15613 (N_15613,N_14777,N_14877);
and U15614 (N_15614,N_14711,N_14948);
nand U15615 (N_15615,N_14379,N_14407);
nor U15616 (N_15616,N_14310,N_14595);
nand U15617 (N_15617,N_14938,N_14583);
nand U15618 (N_15618,N_14391,N_14387);
and U15619 (N_15619,N_14376,N_14824);
xnor U15620 (N_15620,N_14712,N_14614);
xor U15621 (N_15621,N_14529,N_14493);
and U15622 (N_15622,N_14713,N_14478);
and U15623 (N_15623,N_14312,N_14833);
nor U15624 (N_15624,N_14189,N_14599);
xor U15625 (N_15625,N_14068,N_14290);
or U15626 (N_15626,N_14684,N_14950);
nand U15627 (N_15627,N_14078,N_14209);
nand U15628 (N_15628,N_14657,N_14008);
nor U15629 (N_15629,N_14980,N_14759);
nand U15630 (N_15630,N_14574,N_14969);
xnor U15631 (N_15631,N_14391,N_14463);
nor U15632 (N_15632,N_14301,N_14063);
or U15633 (N_15633,N_14330,N_14653);
xnor U15634 (N_15634,N_14199,N_14188);
nor U15635 (N_15635,N_14758,N_14092);
nor U15636 (N_15636,N_14917,N_14557);
nor U15637 (N_15637,N_14871,N_14942);
nor U15638 (N_15638,N_14514,N_14924);
nand U15639 (N_15639,N_14302,N_14972);
and U15640 (N_15640,N_14339,N_14302);
and U15641 (N_15641,N_14785,N_14225);
xor U15642 (N_15642,N_14846,N_14242);
xnor U15643 (N_15643,N_14507,N_14123);
nor U15644 (N_15644,N_14380,N_14566);
xor U15645 (N_15645,N_14039,N_14701);
nor U15646 (N_15646,N_14823,N_14245);
and U15647 (N_15647,N_14522,N_14527);
xnor U15648 (N_15648,N_14649,N_14980);
or U15649 (N_15649,N_14315,N_14533);
or U15650 (N_15650,N_14106,N_14715);
nand U15651 (N_15651,N_14466,N_14385);
or U15652 (N_15652,N_14637,N_14088);
and U15653 (N_15653,N_14803,N_14355);
xor U15654 (N_15654,N_14272,N_14511);
and U15655 (N_15655,N_14594,N_14873);
nor U15656 (N_15656,N_14842,N_14138);
xor U15657 (N_15657,N_14459,N_14747);
nand U15658 (N_15658,N_14172,N_14979);
and U15659 (N_15659,N_14111,N_14128);
or U15660 (N_15660,N_14319,N_14717);
nor U15661 (N_15661,N_14122,N_14684);
nand U15662 (N_15662,N_14132,N_14680);
and U15663 (N_15663,N_14122,N_14043);
xor U15664 (N_15664,N_14494,N_14288);
nor U15665 (N_15665,N_14961,N_14601);
nand U15666 (N_15666,N_14845,N_14661);
and U15667 (N_15667,N_14126,N_14587);
and U15668 (N_15668,N_14759,N_14465);
or U15669 (N_15669,N_14539,N_14162);
nand U15670 (N_15670,N_14194,N_14907);
nand U15671 (N_15671,N_14292,N_14668);
nor U15672 (N_15672,N_14964,N_14656);
nor U15673 (N_15673,N_14502,N_14499);
and U15674 (N_15674,N_14036,N_14671);
and U15675 (N_15675,N_14858,N_14819);
and U15676 (N_15676,N_14949,N_14194);
nand U15677 (N_15677,N_14039,N_14635);
nor U15678 (N_15678,N_14488,N_14209);
nand U15679 (N_15679,N_14189,N_14182);
and U15680 (N_15680,N_14384,N_14064);
nor U15681 (N_15681,N_14913,N_14918);
nor U15682 (N_15682,N_14154,N_14389);
nor U15683 (N_15683,N_14835,N_14422);
nand U15684 (N_15684,N_14362,N_14154);
xnor U15685 (N_15685,N_14087,N_14619);
and U15686 (N_15686,N_14410,N_14465);
nor U15687 (N_15687,N_14013,N_14929);
nor U15688 (N_15688,N_14414,N_14218);
nand U15689 (N_15689,N_14704,N_14937);
nand U15690 (N_15690,N_14103,N_14667);
nand U15691 (N_15691,N_14881,N_14898);
or U15692 (N_15692,N_14714,N_14718);
xnor U15693 (N_15693,N_14491,N_14331);
nor U15694 (N_15694,N_14280,N_14667);
nand U15695 (N_15695,N_14472,N_14330);
xnor U15696 (N_15696,N_14487,N_14971);
nand U15697 (N_15697,N_14910,N_14937);
xor U15698 (N_15698,N_14703,N_14754);
nor U15699 (N_15699,N_14567,N_14884);
xnor U15700 (N_15700,N_14064,N_14499);
and U15701 (N_15701,N_14500,N_14583);
nor U15702 (N_15702,N_14551,N_14196);
xnor U15703 (N_15703,N_14645,N_14608);
or U15704 (N_15704,N_14323,N_14067);
xnor U15705 (N_15705,N_14349,N_14015);
nor U15706 (N_15706,N_14000,N_14827);
or U15707 (N_15707,N_14219,N_14843);
nor U15708 (N_15708,N_14848,N_14304);
nand U15709 (N_15709,N_14470,N_14408);
xnor U15710 (N_15710,N_14315,N_14772);
or U15711 (N_15711,N_14109,N_14138);
or U15712 (N_15712,N_14070,N_14744);
or U15713 (N_15713,N_14735,N_14826);
and U15714 (N_15714,N_14509,N_14211);
and U15715 (N_15715,N_14583,N_14308);
and U15716 (N_15716,N_14124,N_14953);
nor U15717 (N_15717,N_14099,N_14478);
and U15718 (N_15718,N_14462,N_14617);
nor U15719 (N_15719,N_14163,N_14463);
xor U15720 (N_15720,N_14581,N_14832);
nand U15721 (N_15721,N_14985,N_14164);
or U15722 (N_15722,N_14223,N_14782);
and U15723 (N_15723,N_14311,N_14564);
nor U15724 (N_15724,N_14875,N_14425);
xor U15725 (N_15725,N_14716,N_14059);
xor U15726 (N_15726,N_14823,N_14235);
nor U15727 (N_15727,N_14203,N_14283);
nand U15728 (N_15728,N_14909,N_14309);
xnor U15729 (N_15729,N_14404,N_14448);
and U15730 (N_15730,N_14176,N_14697);
or U15731 (N_15731,N_14645,N_14976);
xor U15732 (N_15732,N_14804,N_14209);
and U15733 (N_15733,N_14021,N_14937);
and U15734 (N_15734,N_14475,N_14921);
nand U15735 (N_15735,N_14948,N_14998);
and U15736 (N_15736,N_14041,N_14336);
or U15737 (N_15737,N_14207,N_14257);
nand U15738 (N_15738,N_14816,N_14910);
nand U15739 (N_15739,N_14645,N_14567);
xnor U15740 (N_15740,N_14710,N_14108);
and U15741 (N_15741,N_14203,N_14371);
xnor U15742 (N_15742,N_14239,N_14002);
nand U15743 (N_15743,N_14035,N_14369);
xor U15744 (N_15744,N_14624,N_14957);
xnor U15745 (N_15745,N_14496,N_14502);
nor U15746 (N_15746,N_14580,N_14926);
and U15747 (N_15747,N_14704,N_14608);
xnor U15748 (N_15748,N_14189,N_14027);
xnor U15749 (N_15749,N_14257,N_14768);
xnor U15750 (N_15750,N_14887,N_14068);
or U15751 (N_15751,N_14210,N_14097);
xor U15752 (N_15752,N_14705,N_14948);
and U15753 (N_15753,N_14014,N_14763);
xnor U15754 (N_15754,N_14065,N_14929);
and U15755 (N_15755,N_14423,N_14347);
xnor U15756 (N_15756,N_14485,N_14218);
xnor U15757 (N_15757,N_14654,N_14090);
or U15758 (N_15758,N_14327,N_14399);
nand U15759 (N_15759,N_14439,N_14574);
nand U15760 (N_15760,N_14181,N_14725);
nand U15761 (N_15761,N_14284,N_14318);
xor U15762 (N_15762,N_14902,N_14797);
nor U15763 (N_15763,N_14842,N_14474);
nand U15764 (N_15764,N_14444,N_14543);
nand U15765 (N_15765,N_14331,N_14517);
or U15766 (N_15766,N_14571,N_14437);
nor U15767 (N_15767,N_14695,N_14615);
nand U15768 (N_15768,N_14675,N_14130);
nor U15769 (N_15769,N_14838,N_14063);
or U15770 (N_15770,N_14327,N_14960);
xor U15771 (N_15771,N_14353,N_14210);
xor U15772 (N_15772,N_14437,N_14178);
and U15773 (N_15773,N_14090,N_14482);
nand U15774 (N_15774,N_14655,N_14278);
nor U15775 (N_15775,N_14373,N_14266);
or U15776 (N_15776,N_14971,N_14787);
or U15777 (N_15777,N_14377,N_14054);
and U15778 (N_15778,N_14225,N_14729);
nand U15779 (N_15779,N_14048,N_14708);
and U15780 (N_15780,N_14826,N_14749);
xnor U15781 (N_15781,N_14557,N_14856);
xor U15782 (N_15782,N_14145,N_14551);
and U15783 (N_15783,N_14529,N_14185);
xnor U15784 (N_15784,N_14541,N_14250);
nor U15785 (N_15785,N_14568,N_14050);
nand U15786 (N_15786,N_14909,N_14416);
and U15787 (N_15787,N_14370,N_14329);
nand U15788 (N_15788,N_14780,N_14880);
and U15789 (N_15789,N_14999,N_14287);
or U15790 (N_15790,N_14129,N_14542);
nor U15791 (N_15791,N_14536,N_14701);
nor U15792 (N_15792,N_14960,N_14478);
or U15793 (N_15793,N_14307,N_14771);
xnor U15794 (N_15794,N_14047,N_14344);
or U15795 (N_15795,N_14151,N_14255);
and U15796 (N_15796,N_14689,N_14408);
xnor U15797 (N_15797,N_14019,N_14647);
nand U15798 (N_15798,N_14500,N_14882);
and U15799 (N_15799,N_14225,N_14127);
xnor U15800 (N_15800,N_14933,N_14552);
nand U15801 (N_15801,N_14430,N_14769);
nor U15802 (N_15802,N_14705,N_14669);
and U15803 (N_15803,N_14259,N_14846);
and U15804 (N_15804,N_14933,N_14540);
nand U15805 (N_15805,N_14678,N_14992);
nor U15806 (N_15806,N_14705,N_14801);
and U15807 (N_15807,N_14358,N_14485);
nand U15808 (N_15808,N_14791,N_14198);
and U15809 (N_15809,N_14928,N_14198);
or U15810 (N_15810,N_14216,N_14876);
xnor U15811 (N_15811,N_14752,N_14276);
nand U15812 (N_15812,N_14076,N_14274);
nor U15813 (N_15813,N_14603,N_14294);
xor U15814 (N_15814,N_14835,N_14694);
xor U15815 (N_15815,N_14433,N_14361);
nor U15816 (N_15816,N_14052,N_14054);
nand U15817 (N_15817,N_14999,N_14521);
or U15818 (N_15818,N_14314,N_14648);
xnor U15819 (N_15819,N_14357,N_14116);
nand U15820 (N_15820,N_14901,N_14685);
nor U15821 (N_15821,N_14894,N_14288);
and U15822 (N_15822,N_14010,N_14191);
xnor U15823 (N_15823,N_14432,N_14420);
or U15824 (N_15824,N_14708,N_14056);
and U15825 (N_15825,N_14530,N_14400);
xor U15826 (N_15826,N_14512,N_14383);
xnor U15827 (N_15827,N_14412,N_14594);
nor U15828 (N_15828,N_14968,N_14293);
xor U15829 (N_15829,N_14477,N_14852);
nor U15830 (N_15830,N_14383,N_14138);
nor U15831 (N_15831,N_14052,N_14117);
nand U15832 (N_15832,N_14682,N_14470);
or U15833 (N_15833,N_14059,N_14214);
nand U15834 (N_15834,N_14498,N_14367);
nand U15835 (N_15835,N_14154,N_14358);
xor U15836 (N_15836,N_14724,N_14836);
and U15837 (N_15837,N_14012,N_14955);
and U15838 (N_15838,N_14656,N_14319);
or U15839 (N_15839,N_14850,N_14656);
xnor U15840 (N_15840,N_14516,N_14534);
and U15841 (N_15841,N_14456,N_14473);
or U15842 (N_15842,N_14993,N_14130);
xnor U15843 (N_15843,N_14112,N_14496);
nand U15844 (N_15844,N_14787,N_14747);
xor U15845 (N_15845,N_14518,N_14563);
nand U15846 (N_15846,N_14272,N_14089);
xnor U15847 (N_15847,N_14608,N_14328);
nor U15848 (N_15848,N_14417,N_14928);
and U15849 (N_15849,N_14270,N_14530);
or U15850 (N_15850,N_14119,N_14617);
nand U15851 (N_15851,N_14863,N_14269);
or U15852 (N_15852,N_14797,N_14957);
and U15853 (N_15853,N_14951,N_14380);
and U15854 (N_15854,N_14689,N_14010);
nand U15855 (N_15855,N_14972,N_14362);
nor U15856 (N_15856,N_14852,N_14442);
nor U15857 (N_15857,N_14204,N_14335);
nor U15858 (N_15858,N_14226,N_14961);
or U15859 (N_15859,N_14959,N_14882);
xnor U15860 (N_15860,N_14777,N_14181);
xor U15861 (N_15861,N_14943,N_14354);
or U15862 (N_15862,N_14179,N_14812);
and U15863 (N_15863,N_14403,N_14627);
nand U15864 (N_15864,N_14833,N_14392);
xor U15865 (N_15865,N_14618,N_14454);
nand U15866 (N_15866,N_14952,N_14595);
and U15867 (N_15867,N_14793,N_14408);
and U15868 (N_15868,N_14139,N_14228);
xor U15869 (N_15869,N_14760,N_14902);
nor U15870 (N_15870,N_14630,N_14066);
or U15871 (N_15871,N_14473,N_14834);
xor U15872 (N_15872,N_14379,N_14721);
or U15873 (N_15873,N_14488,N_14356);
and U15874 (N_15874,N_14839,N_14200);
or U15875 (N_15875,N_14939,N_14580);
nand U15876 (N_15876,N_14029,N_14896);
nand U15877 (N_15877,N_14810,N_14307);
xnor U15878 (N_15878,N_14345,N_14252);
and U15879 (N_15879,N_14435,N_14469);
or U15880 (N_15880,N_14333,N_14055);
xor U15881 (N_15881,N_14139,N_14871);
xnor U15882 (N_15882,N_14389,N_14189);
nand U15883 (N_15883,N_14933,N_14254);
nand U15884 (N_15884,N_14353,N_14316);
or U15885 (N_15885,N_14648,N_14267);
nor U15886 (N_15886,N_14747,N_14610);
and U15887 (N_15887,N_14642,N_14606);
nor U15888 (N_15888,N_14588,N_14591);
and U15889 (N_15889,N_14417,N_14395);
and U15890 (N_15890,N_14719,N_14311);
nor U15891 (N_15891,N_14226,N_14921);
xnor U15892 (N_15892,N_14533,N_14402);
nand U15893 (N_15893,N_14477,N_14908);
nor U15894 (N_15894,N_14289,N_14731);
and U15895 (N_15895,N_14875,N_14665);
nor U15896 (N_15896,N_14893,N_14644);
xor U15897 (N_15897,N_14159,N_14355);
xor U15898 (N_15898,N_14748,N_14336);
or U15899 (N_15899,N_14118,N_14038);
xnor U15900 (N_15900,N_14814,N_14788);
xnor U15901 (N_15901,N_14456,N_14955);
and U15902 (N_15902,N_14132,N_14414);
xor U15903 (N_15903,N_14533,N_14829);
nor U15904 (N_15904,N_14679,N_14397);
xnor U15905 (N_15905,N_14316,N_14802);
and U15906 (N_15906,N_14174,N_14564);
nor U15907 (N_15907,N_14620,N_14287);
or U15908 (N_15908,N_14297,N_14058);
or U15909 (N_15909,N_14962,N_14063);
nand U15910 (N_15910,N_14401,N_14930);
and U15911 (N_15911,N_14116,N_14584);
and U15912 (N_15912,N_14546,N_14234);
nor U15913 (N_15913,N_14337,N_14886);
and U15914 (N_15914,N_14097,N_14045);
nand U15915 (N_15915,N_14409,N_14609);
xor U15916 (N_15916,N_14083,N_14364);
and U15917 (N_15917,N_14986,N_14185);
xnor U15918 (N_15918,N_14590,N_14913);
nor U15919 (N_15919,N_14808,N_14935);
nand U15920 (N_15920,N_14027,N_14680);
xor U15921 (N_15921,N_14587,N_14634);
nor U15922 (N_15922,N_14264,N_14789);
xor U15923 (N_15923,N_14268,N_14477);
xor U15924 (N_15924,N_14485,N_14342);
or U15925 (N_15925,N_14323,N_14663);
xor U15926 (N_15926,N_14970,N_14851);
nor U15927 (N_15927,N_14189,N_14497);
nor U15928 (N_15928,N_14550,N_14765);
xor U15929 (N_15929,N_14780,N_14395);
or U15930 (N_15930,N_14980,N_14791);
nand U15931 (N_15931,N_14661,N_14896);
and U15932 (N_15932,N_14030,N_14741);
and U15933 (N_15933,N_14228,N_14605);
or U15934 (N_15934,N_14433,N_14222);
nand U15935 (N_15935,N_14389,N_14752);
and U15936 (N_15936,N_14064,N_14161);
nor U15937 (N_15937,N_14742,N_14710);
or U15938 (N_15938,N_14070,N_14896);
or U15939 (N_15939,N_14003,N_14157);
nand U15940 (N_15940,N_14326,N_14411);
or U15941 (N_15941,N_14430,N_14089);
xnor U15942 (N_15942,N_14023,N_14607);
or U15943 (N_15943,N_14727,N_14938);
or U15944 (N_15944,N_14582,N_14502);
and U15945 (N_15945,N_14521,N_14059);
nand U15946 (N_15946,N_14423,N_14889);
xor U15947 (N_15947,N_14628,N_14306);
and U15948 (N_15948,N_14896,N_14627);
nor U15949 (N_15949,N_14678,N_14790);
nand U15950 (N_15950,N_14792,N_14628);
nor U15951 (N_15951,N_14828,N_14460);
or U15952 (N_15952,N_14968,N_14476);
xor U15953 (N_15953,N_14331,N_14131);
and U15954 (N_15954,N_14168,N_14803);
nor U15955 (N_15955,N_14423,N_14905);
and U15956 (N_15956,N_14772,N_14374);
nand U15957 (N_15957,N_14835,N_14435);
nor U15958 (N_15958,N_14367,N_14603);
or U15959 (N_15959,N_14531,N_14534);
nand U15960 (N_15960,N_14846,N_14995);
or U15961 (N_15961,N_14977,N_14028);
or U15962 (N_15962,N_14323,N_14441);
nand U15963 (N_15963,N_14642,N_14944);
nand U15964 (N_15964,N_14389,N_14155);
or U15965 (N_15965,N_14161,N_14788);
nand U15966 (N_15966,N_14583,N_14176);
nor U15967 (N_15967,N_14753,N_14042);
nand U15968 (N_15968,N_14650,N_14400);
and U15969 (N_15969,N_14724,N_14632);
and U15970 (N_15970,N_14520,N_14574);
nor U15971 (N_15971,N_14302,N_14040);
nand U15972 (N_15972,N_14200,N_14937);
xor U15973 (N_15973,N_14499,N_14867);
nand U15974 (N_15974,N_14503,N_14235);
nor U15975 (N_15975,N_14199,N_14139);
nor U15976 (N_15976,N_14878,N_14838);
xor U15977 (N_15977,N_14984,N_14684);
xnor U15978 (N_15978,N_14305,N_14545);
nor U15979 (N_15979,N_14376,N_14543);
and U15980 (N_15980,N_14140,N_14351);
and U15981 (N_15981,N_14890,N_14203);
and U15982 (N_15982,N_14741,N_14041);
nor U15983 (N_15983,N_14167,N_14161);
nand U15984 (N_15984,N_14756,N_14581);
and U15985 (N_15985,N_14906,N_14980);
or U15986 (N_15986,N_14967,N_14674);
or U15987 (N_15987,N_14063,N_14741);
or U15988 (N_15988,N_14376,N_14425);
and U15989 (N_15989,N_14874,N_14696);
or U15990 (N_15990,N_14832,N_14933);
nor U15991 (N_15991,N_14456,N_14450);
xor U15992 (N_15992,N_14357,N_14052);
nand U15993 (N_15993,N_14441,N_14696);
or U15994 (N_15994,N_14473,N_14538);
and U15995 (N_15995,N_14096,N_14670);
and U15996 (N_15996,N_14217,N_14154);
xor U15997 (N_15997,N_14580,N_14955);
nand U15998 (N_15998,N_14899,N_14013);
nand U15999 (N_15999,N_14534,N_14419);
nor U16000 (N_16000,N_15649,N_15028);
or U16001 (N_16001,N_15607,N_15755);
nor U16002 (N_16002,N_15447,N_15078);
nand U16003 (N_16003,N_15006,N_15105);
or U16004 (N_16004,N_15528,N_15308);
nand U16005 (N_16005,N_15323,N_15682);
xnor U16006 (N_16006,N_15088,N_15330);
or U16007 (N_16007,N_15773,N_15997);
and U16008 (N_16008,N_15551,N_15966);
and U16009 (N_16009,N_15871,N_15557);
or U16010 (N_16010,N_15146,N_15867);
nor U16011 (N_16011,N_15835,N_15362);
or U16012 (N_16012,N_15383,N_15374);
and U16013 (N_16013,N_15737,N_15222);
nand U16014 (N_16014,N_15510,N_15931);
nand U16015 (N_16015,N_15482,N_15377);
nand U16016 (N_16016,N_15511,N_15824);
nand U16017 (N_16017,N_15698,N_15556);
and U16018 (N_16018,N_15946,N_15788);
or U16019 (N_16019,N_15531,N_15672);
nand U16020 (N_16020,N_15422,N_15313);
or U16021 (N_16021,N_15353,N_15174);
nor U16022 (N_16022,N_15805,N_15483);
and U16023 (N_16023,N_15411,N_15999);
nor U16024 (N_16024,N_15332,N_15224);
nand U16025 (N_16025,N_15608,N_15303);
nor U16026 (N_16026,N_15387,N_15081);
nor U16027 (N_16027,N_15513,N_15667);
or U16028 (N_16028,N_15173,N_15991);
or U16029 (N_16029,N_15416,N_15256);
and U16030 (N_16030,N_15165,N_15379);
and U16031 (N_16031,N_15220,N_15590);
xnor U16032 (N_16032,N_15271,N_15123);
xnor U16033 (N_16033,N_15331,N_15978);
and U16034 (N_16034,N_15480,N_15525);
or U16035 (N_16035,N_15136,N_15106);
xor U16036 (N_16036,N_15104,N_15769);
and U16037 (N_16037,N_15240,N_15190);
nor U16038 (N_16038,N_15782,N_15428);
and U16039 (N_16039,N_15681,N_15650);
nor U16040 (N_16040,N_15077,N_15058);
or U16041 (N_16041,N_15318,N_15919);
nand U16042 (N_16042,N_15785,N_15098);
xnor U16043 (N_16043,N_15947,N_15490);
nand U16044 (N_16044,N_15524,N_15139);
xnor U16045 (N_16045,N_15301,N_15831);
nand U16046 (N_16046,N_15037,N_15419);
nor U16047 (N_16047,N_15679,N_15881);
and U16048 (N_16048,N_15237,N_15138);
nor U16049 (N_16049,N_15217,N_15870);
nand U16050 (N_16050,N_15904,N_15839);
nor U16051 (N_16051,N_15739,N_15656);
xor U16052 (N_16052,N_15235,N_15520);
and U16053 (N_16053,N_15215,N_15502);
or U16054 (N_16054,N_15474,N_15960);
nand U16055 (N_16055,N_15707,N_15726);
and U16056 (N_16056,N_15334,N_15521);
and U16057 (N_16057,N_15363,N_15924);
nand U16058 (N_16058,N_15748,N_15774);
nor U16059 (N_16059,N_15814,N_15856);
and U16060 (N_16060,N_15792,N_15840);
nand U16061 (N_16061,N_15963,N_15674);
nand U16062 (N_16062,N_15213,N_15514);
nor U16063 (N_16063,N_15722,N_15324);
and U16064 (N_16064,N_15024,N_15113);
xnor U16065 (N_16065,N_15427,N_15418);
or U16066 (N_16066,N_15336,N_15255);
or U16067 (N_16067,N_15749,N_15084);
nor U16068 (N_16068,N_15896,N_15654);
nand U16069 (N_16069,N_15056,N_15284);
or U16070 (N_16070,N_15412,N_15633);
nor U16071 (N_16071,N_15380,N_15048);
and U16072 (N_16072,N_15766,N_15397);
nor U16073 (N_16073,N_15877,N_15163);
or U16074 (N_16074,N_15593,N_15148);
nand U16075 (N_16075,N_15152,N_15075);
or U16076 (N_16076,N_15250,N_15600);
and U16077 (N_16077,N_15875,N_15697);
nand U16078 (N_16078,N_15503,N_15258);
xnor U16079 (N_16079,N_15478,N_15761);
nor U16080 (N_16080,N_15093,N_15144);
or U16081 (N_16081,N_15815,N_15309);
nand U16082 (N_16082,N_15276,N_15967);
and U16083 (N_16083,N_15598,N_15643);
nor U16084 (N_16084,N_15279,N_15920);
nand U16085 (N_16085,N_15696,N_15189);
xor U16086 (N_16086,N_15494,N_15818);
nand U16087 (N_16087,N_15929,N_15851);
nand U16088 (N_16088,N_15721,N_15927);
xor U16089 (N_16089,N_15245,N_15440);
and U16090 (N_16090,N_15197,N_15984);
or U16091 (N_16091,N_15689,N_15264);
nand U16092 (N_16092,N_15254,N_15372);
and U16093 (N_16093,N_15094,N_15351);
nor U16094 (N_16094,N_15114,N_15781);
or U16095 (N_16095,N_15054,N_15357);
or U16096 (N_16096,N_15122,N_15405);
nor U16097 (N_16097,N_15601,N_15089);
xor U16098 (N_16098,N_15631,N_15787);
and U16099 (N_16099,N_15652,N_15403);
or U16100 (N_16100,N_15670,N_15498);
nand U16101 (N_16101,N_15925,N_15425);
nor U16102 (N_16102,N_15901,N_15731);
and U16103 (N_16103,N_15622,N_15181);
and U16104 (N_16104,N_15062,N_15789);
and U16105 (N_16105,N_15985,N_15548);
nor U16106 (N_16106,N_15198,N_15472);
or U16107 (N_16107,N_15176,N_15708);
nand U16108 (N_16108,N_15434,N_15302);
nand U16109 (N_16109,N_15545,N_15050);
and U16110 (N_16110,N_15504,N_15897);
or U16111 (N_16111,N_15149,N_15025);
xnor U16112 (N_16112,N_15185,N_15981);
or U16113 (N_16113,N_15333,N_15147);
or U16114 (N_16114,N_15996,N_15571);
xor U16115 (N_16115,N_15687,N_15888);
nand U16116 (N_16116,N_15020,N_15116);
or U16117 (N_16117,N_15413,N_15141);
nor U16118 (N_16118,N_15164,N_15349);
nand U16119 (N_16119,N_15791,N_15690);
or U16120 (N_16120,N_15797,N_15779);
xnor U16121 (N_16121,N_15051,N_15120);
xor U16122 (N_16122,N_15311,N_15740);
or U16123 (N_16123,N_15068,N_15639);
xor U16124 (N_16124,N_15903,N_15407);
nand U16125 (N_16125,N_15004,N_15205);
and U16126 (N_16126,N_15424,N_15420);
or U16127 (N_16127,N_15591,N_15251);
nand U16128 (N_16128,N_15756,N_15270);
or U16129 (N_16129,N_15341,N_15400);
xor U16130 (N_16130,N_15874,N_15913);
xor U16131 (N_16131,N_15705,N_15854);
and U16132 (N_16132,N_15399,N_15073);
and U16133 (N_16133,N_15575,N_15476);
or U16134 (N_16134,N_15429,N_15908);
or U16135 (N_16135,N_15039,N_15325);
xor U16136 (N_16136,N_15530,N_15277);
and U16137 (N_16137,N_15227,N_15370);
nor U16138 (N_16138,N_15605,N_15312);
and U16139 (N_16139,N_15635,N_15793);
nand U16140 (N_16140,N_15828,N_15604);
or U16141 (N_16141,N_15768,N_15449);
and U16142 (N_16142,N_15486,N_15550);
nand U16143 (N_16143,N_15119,N_15415);
xor U16144 (N_16144,N_15445,N_15493);
nand U16145 (N_16145,N_15743,N_15041);
xnor U16146 (N_16146,N_15337,N_15365);
nand U16147 (N_16147,N_15950,N_15375);
or U16148 (N_16148,N_15975,N_15310);
or U16149 (N_16149,N_15944,N_15135);
xnor U16150 (N_16150,N_15653,N_15388);
xnor U16151 (N_16151,N_15547,N_15384);
and U16152 (N_16152,N_15853,N_15053);
nor U16153 (N_16153,N_15118,N_15408);
and U16154 (N_16154,N_15640,N_15448);
xor U16155 (N_16155,N_15491,N_15451);
xnor U16156 (N_16156,N_15281,N_15226);
xor U16157 (N_16157,N_15468,N_15023);
xor U16158 (N_16158,N_15659,N_15618);
or U16159 (N_16159,N_15001,N_15803);
and U16160 (N_16160,N_15012,N_15177);
and U16161 (N_16161,N_15130,N_15280);
or U16162 (N_16162,N_15910,N_15350);
nor U16163 (N_16163,N_15439,N_15942);
and U16164 (N_16164,N_15263,N_15868);
and U16165 (N_16165,N_15540,N_15988);
or U16166 (N_16166,N_15795,N_15560);
nor U16167 (N_16167,N_15460,N_15500);
nor U16168 (N_16168,N_15433,N_15579);
or U16169 (N_16169,N_15395,N_15907);
xnor U16170 (N_16170,N_15335,N_15225);
nor U16171 (N_16171,N_15770,N_15552);
xor U16172 (N_16172,N_15750,N_15275);
nand U16173 (N_16173,N_15783,N_15695);
xnor U16174 (N_16174,N_15466,N_15706);
nor U16175 (N_16175,N_15969,N_15732);
xor U16176 (N_16176,N_15059,N_15402);
nand U16177 (N_16177,N_15269,N_15352);
xnor U16178 (N_16178,N_15763,N_15542);
nand U16179 (N_16179,N_15668,N_15305);
or U16180 (N_16180,N_15872,N_15720);
and U16181 (N_16181,N_15716,N_15718);
and U16182 (N_16182,N_15693,N_15671);
xor U16183 (N_16183,N_15249,N_15047);
and U16184 (N_16184,N_15183,N_15565);
nor U16185 (N_16185,N_15293,N_15287);
nor U16186 (N_16186,N_15443,N_15206);
or U16187 (N_16187,N_15736,N_15473);
nand U16188 (N_16188,N_15481,N_15055);
nand U16189 (N_16189,N_15133,N_15949);
xnor U16190 (N_16190,N_15159,N_15848);
nand U16191 (N_16191,N_15369,N_15233);
and U16192 (N_16192,N_15188,N_15813);
nor U16193 (N_16193,N_15517,N_15994);
or U16194 (N_16194,N_15841,N_15317);
or U16195 (N_16195,N_15930,N_15583);
or U16196 (N_16196,N_15801,N_15112);
or U16197 (N_16197,N_15385,N_15961);
and U16198 (N_16198,N_15389,N_15862);
or U16199 (N_16199,N_15603,N_15728);
or U16200 (N_16200,N_15941,N_15321);
and U16201 (N_16201,N_15115,N_15137);
xnor U16202 (N_16202,N_15157,N_15328);
nor U16203 (N_16203,N_15409,N_15858);
xor U16204 (N_16204,N_15630,N_15817);
or U16205 (N_16205,N_15594,N_15035);
nor U16206 (N_16206,N_15034,N_15767);
nor U16207 (N_16207,N_15936,N_15134);
xor U16208 (N_16208,N_15200,N_15715);
nand U16209 (N_16209,N_15169,N_15285);
nor U16210 (N_16210,N_15691,N_15725);
xor U16211 (N_16211,N_15381,N_15762);
nor U16212 (N_16212,N_15734,N_15107);
xor U16213 (N_16213,N_15982,N_15757);
and U16214 (N_16214,N_15348,N_15660);
nor U16215 (N_16215,N_15121,N_15866);
xor U16216 (N_16216,N_15194,N_15912);
xor U16217 (N_16217,N_15760,N_15651);
xnor U16218 (N_16218,N_15515,N_15296);
nor U16219 (N_16219,N_15009,N_15290);
and U16220 (N_16220,N_15219,N_15299);
and U16221 (N_16221,N_15628,N_15602);
xor U16222 (N_16222,N_15017,N_15469);
xor U16223 (N_16223,N_15234,N_15849);
or U16224 (N_16224,N_15150,N_15532);
nor U16225 (N_16225,N_15678,N_15184);
or U16226 (N_16226,N_15989,N_15153);
nand U16227 (N_16227,N_15526,N_15446);
and U16228 (N_16228,N_15923,N_15329);
and U16229 (N_16229,N_15616,N_15090);
nand U16230 (N_16230,N_15005,N_15719);
nor U16231 (N_16231,N_15142,N_15562);
nand U16232 (N_16232,N_15980,N_15366);
nand U16233 (N_16233,N_15573,N_15778);
xnor U16234 (N_16234,N_15585,N_15692);
and U16235 (N_16235,N_15044,N_15800);
xor U16236 (N_16236,N_15228,N_15855);
nor U16237 (N_16237,N_15223,N_15257);
nor U16238 (N_16238,N_15555,N_15821);
nor U16239 (N_16239,N_15820,N_15661);
and U16240 (N_16240,N_15627,N_15968);
or U16241 (N_16241,N_15666,N_15906);
nor U16242 (N_16242,N_15236,N_15470);
nand U16243 (N_16243,N_15554,N_15995);
or U16244 (N_16244,N_15845,N_15117);
xnor U16245 (N_16245,N_15155,N_15100);
and U16246 (N_16246,N_15242,N_15209);
nand U16247 (N_16247,N_15764,N_15175);
nor U16248 (N_16248,N_15637,N_15536);
and U16249 (N_16249,N_15248,N_15799);
nand U16250 (N_16250,N_15216,N_15742);
xor U16251 (N_16251,N_15029,N_15648);
or U16252 (N_16252,N_15915,N_15027);
nand U16253 (N_16253,N_15192,N_15928);
nor U16254 (N_16254,N_15326,N_15124);
or U16255 (N_16255,N_15677,N_15902);
xor U16256 (N_16256,N_15373,N_15361);
and U16257 (N_16257,N_15570,N_15626);
and U16258 (N_16258,N_15066,N_15376);
nor U16259 (N_16259,N_15158,N_15645);
or U16260 (N_16260,N_15315,N_15431);
nor U16261 (N_16261,N_15834,N_15688);
nand U16262 (N_16262,N_15067,N_15426);
xnor U16263 (N_16263,N_15404,N_15683);
nor U16264 (N_16264,N_15771,N_15232);
or U16265 (N_16265,N_15878,N_15492);
or U16266 (N_16266,N_15452,N_15956);
nor U16267 (N_16267,N_15010,N_15092);
or U16268 (N_16268,N_15527,N_15979);
and U16269 (N_16269,N_15578,N_15684);
nand U16270 (N_16270,N_15109,N_15926);
and U16271 (N_16271,N_15702,N_15391);
xor U16272 (N_16272,N_15022,N_15806);
nor U16273 (N_16273,N_15441,N_15450);
nand U16274 (N_16274,N_15701,N_15421);
and U16275 (N_16275,N_15191,N_15561);
and U16276 (N_16276,N_15873,N_15355);
nand U16277 (N_16277,N_15955,N_15523);
or U16278 (N_16278,N_15247,N_15617);
xor U16279 (N_16279,N_15438,N_15809);
or U16280 (N_16280,N_15563,N_15614);
or U16281 (N_16281,N_15259,N_15040);
xor U16282 (N_16282,N_15751,N_15463);
and U16283 (N_16283,N_15162,N_15798);
and U16284 (N_16284,N_15143,N_15609);
nor U16285 (N_16285,N_15414,N_15647);
nand U16286 (N_16286,N_15951,N_15338);
nand U16287 (N_16287,N_15052,N_15916);
or U16288 (N_16288,N_15457,N_15266);
or U16289 (N_16289,N_15884,N_15125);
xor U16290 (N_16290,N_15595,N_15909);
and U16291 (N_16291,N_15599,N_15673);
xor U16292 (N_16292,N_15819,N_15241);
and U16293 (N_16293,N_15160,N_15364);
and U16294 (N_16294,N_15973,N_15156);
xnor U16295 (N_16295,N_15069,N_15586);
or U16296 (N_16296,N_15826,N_15072);
nand U16297 (N_16297,N_15529,N_15102);
and U16298 (N_16298,N_15099,N_15008);
xnor U16299 (N_16299,N_15295,N_15339);
nand U16300 (N_16300,N_15253,N_15998);
nor U16301 (N_16301,N_15442,N_15863);
or U16302 (N_16302,N_15300,N_15972);
and U16303 (N_16303,N_15892,N_15231);
nand U16304 (N_16304,N_15320,N_15852);
or U16305 (N_16305,N_15546,N_15816);
nand U16306 (N_16306,N_15880,N_15128);
nor U16307 (N_16307,N_15703,N_15087);
nor U16308 (N_16308,N_15566,N_15837);
nor U16309 (N_16309,N_15286,N_15417);
and U16310 (N_16310,N_15976,N_15914);
nand U16311 (N_16311,N_15905,N_15076);
nand U16312 (N_16312,N_15484,N_15161);
xnor U16313 (N_16313,N_15712,N_15581);
xnor U16314 (N_16314,N_15026,N_15918);
xnor U16315 (N_16315,N_15680,N_15857);
nor U16316 (N_16316,N_15045,N_15895);
and U16317 (N_16317,N_15990,N_15534);
or U16318 (N_16318,N_15744,N_15199);
nand U16319 (N_16319,N_15019,N_15790);
xnor U16320 (N_16320,N_15214,N_15836);
nand U16321 (N_16321,N_15611,N_15992);
nand U16322 (N_16322,N_15030,N_15103);
nand U16323 (N_16323,N_15516,N_15390);
and U16324 (N_16324,N_15596,N_15962);
or U16325 (N_16325,N_15606,N_15830);
nand U16326 (N_16326,N_15292,N_15393);
xor U16327 (N_16327,N_15340,N_15060);
or U16328 (N_16328,N_15876,N_15900);
and U16329 (N_16329,N_15274,N_15082);
or U16330 (N_16330,N_15230,N_15196);
or U16331 (N_16331,N_15735,N_15356);
or U16332 (N_16332,N_15584,N_15623);
or U16333 (N_16333,N_15031,N_15965);
nand U16334 (N_16334,N_15210,N_15489);
and U16335 (N_16335,N_15945,N_15487);
or U16336 (N_16336,N_15717,N_15347);
or U16337 (N_16337,N_15238,N_15278);
or U16338 (N_16338,N_15079,N_15610);
nand U16339 (N_16339,N_15638,N_15752);
xnor U16340 (N_16340,N_15589,N_15432);
or U16341 (N_16341,N_15987,N_15435);
nand U16342 (N_16342,N_15002,N_15784);
xor U16343 (N_16343,N_15453,N_15568);
xnor U16344 (N_16344,N_15657,N_15592);
nor U16345 (N_16345,N_15046,N_15580);
and U16346 (N_16346,N_15759,N_15479);
nand U16347 (N_16347,N_15057,N_15166);
nor U16348 (N_16348,N_15095,N_15675);
nor U16349 (N_16349,N_15083,N_15993);
xnor U16350 (N_16350,N_15268,N_15911);
nor U16351 (N_16351,N_15939,N_15894);
xor U16352 (N_16352,N_15890,N_15367);
nand U16353 (N_16353,N_15294,N_15850);
nand U16354 (N_16354,N_15319,N_15694);
nor U16355 (N_16355,N_15847,N_15537);
xnor U16356 (N_16356,N_15049,N_15632);
or U16357 (N_16357,N_15273,N_15015);
nor U16358 (N_16358,N_15179,N_15086);
and U16359 (N_16359,N_15108,N_15097);
nor U16360 (N_16360,N_15954,N_15288);
nor U16361 (N_16361,N_15043,N_15346);
nor U16362 (N_16362,N_15802,N_15260);
nor U16363 (N_16363,N_15170,N_15780);
nor U16364 (N_16364,N_15127,N_15378);
nand U16365 (N_16365,N_15467,N_15444);
nand U16366 (N_16366,N_15282,N_15953);
xnor U16367 (N_16367,N_15676,N_15859);
and U16368 (N_16368,N_15665,N_15304);
or U16369 (N_16369,N_15921,N_15459);
nor U16370 (N_16370,N_15506,N_15615);
nor U16371 (N_16371,N_15063,N_15741);
nor U16372 (N_16372,N_15252,N_15948);
xor U16373 (N_16373,N_15011,N_15934);
nand U16374 (N_16374,N_15832,N_15612);
nand U16375 (N_16375,N_15038,N_15182);
xor U16376 (N_16376,N_15983,N_15343);
nand U16377 (N_16377,N_15016,N_15382);
nand U16378 (N_16378,N_15344,N_15811);
nor U16379 (N_16379,N_15986,N_15297);
nand U16380 (N_16380,N_15882,N_15423);
xnor U16381 (N_16381,N_15624,N_15074);
or U16382 (N_16382,N_15714,N_15641);
or U16383 (N_16383,N_15488,N_15101);
xor U16384 (N_16384,N_15812,N_15619);
nor U16385 (N_16385,N_15723,N_15937);
xor U16386 (N_16386,N_15007,N_15202);
and U16387 (N_16387,N_15964,N_15359);
nor U16388 (N_16388,N_15110,N_15754);
and U16389 (N_16389,N_15777,N_15392);
xor U16390 (N_16390,N_15662,N_15574);
nand U16391 (N_16391,N_15709,N_15091);
or U16392 (N_16392,N_15634,N_15229);
nor U16393 (N_16393,N_15505,N_15132);
or U16394 (N_16394,N_15129,N_15471);
and U16395 (N_16395,N_15765,N_15410);
nor U16396 (N_16396,N_15558,N_15186);
and U16397 (N_16397,N_15401,N_15208);
nand U16398 (N_16398,N_15061,N_15265);
nor U16399 (N_16399,N_15246,N_15577);
nor U16400 (N_16400,N_15636,N_15456);
nand U16401 (N_16401,N_15239,N_15700);
xnor U16402 (N_16402,N_15396,N_15572);
or U16403 (N_16403,N_15746,N_15553);
xor U16404 (N_16404,N_15807,N_15933);
or U16405 (N_16405,N_15710,N_15733);
nor U16406 (N_16406,N_15512,N_15738);
nand U16407 (N_16407,N_15195,N_15111);
xnor U16408 (N_16408,N_15314,N_15977);
and U16409 (N_16409,N_15368,N_15518);
and U16410 (N_16410,N_15167,N_15458);
nand U16411 (N_16411,N_15727,N_15406);
and U16412 (N_16412,N_15283,N_15842);
and U16413 (N_16413,N_15663,N_15544);
or U16414 (N_16414,N_15316,N_15730);
xor U16415 (N_16415,N_15496,N_15014);
or U16416 (N_16416,N_15509,N_15204);
nor U16417 (N_16417,N_15891,N_15291);
nor U16418 (N_16418,N_15358,N_15940);
or U16419 (N_16419,N_15655,N_15776);
and U16420 (N_16420,N_15729,N_15629);
xor U16421 (N_16421,N_15971,N_15932);
nor U16422 (N_16422,N_15644,N_15685);
and U16423 (N_16423,N_15180,N_15898);
nand U16424 (N_16424,N_15151,N_15327);
or U16425 (N_16425,N_15065,N_15808);
and U16426 (N_16426,N_15935,N_15522);
nand U16427 (N_16427,N_15699,N_15211);
nand U16428 (N_16428,N_15064,N_15804);
and U16429 (N_16429,N_15794,N_15822);
xnor U16430 (N_16430,N_15462,N_15207);
or U16431 (N_16431,N_15436,N_15298);
nor U16432 (N_16432,N_15262,N_15243);
nand U16433 (N_16433,N_15597,N_15080);
xnor U16434 (N_16434,N_15454,N_15508);
xor U16435 (N_16435,N_15013,N_15885);
nor U16436 (N_16436,N_15272,N_15464);
xor U16437 (N_16437,N_15430,N_15549);
or U16438 (N_16438,N_15096,N_15032);
nand U16439 (N_16439,N_15796,N_15642);
nand U16440 (N_16440,N_15620,N_15203);
nand U16441 (N_16441,N_15786,N_15861);
xnor U16442 (N_16442,N_15477,N_15843);
and U16443 (N_16443,N_15864,N_15938);
xor U16444 (N_16444,N_15559,N_15846);
or U16445 (N_16445,N_15543,N_15974);
xor U16446 (N_16446,N_15865,N_15775);
nor U16447 (N_16447,N_15289,N_15261);
nand U16448 (N_16448,N_15070,N_15193);
or U16449 (N_16449,N_15922,N_15042);
nand U16450 (N_16450,N_15021,N_15587);
nor U16451 (N_16451,N_15686,N_15394);
nor U16452 (N_16452,N_15747,N_15533);
nor U16453 (N_16453,N_15519,N_15753);
and U16454 (N_16454,N_15507,N_15475);
xnor U16455 (N_16455,N_15582,N_15201);
nand U16456 (N_16456,N_15495,N_15669);
nor U16457 (N_16457,N_15307,N_15154);
and U16458 (N_16458,N_15172,N_15810);
xor U16459 (N_16459,N_15168,N_15386);
or U16460 (N_16460,N_15745,N_15567);
xnor U16461 (N_16461,N_15588,N_15625);
and U16462 (N_16462,N_15838,N_15646);
nor U16463 (N_16463,N_15085,N_15879);
xnor U16464 (N_16464,N_15957,N_15886);
nand U16465 (N_16465,N_15499,N_15036);
and U16466 (N_16466,N_15306,N_15126);
nor U16467 (N_16467,N_15943,N_15887);
nand U16468 (N_16468,N_15485,N_15033);
nor U16469 (N_16469,N_15003,N_15541);
and U16470 (N_16470,N_15825,N_15564);
nor U16471 (N_16471,N_15140,N_15018);
and U16472 (N_16472,N_15664,N_15711);
and U16473 (N_16473,N_15171,N_15218);
and U16474 (N_16474,N_15772,N_15461);
xor U16475 (N_16475,N_15959,N_15538);
xor U16476 (N_16476,N_15501,N_15354);
nand U16477 (N_16477,N_15000,N_15658);
xor U16478 (N_16478,N_15539,N_15244);
nor U16479 (N_16479,N_15958,N_15345);
xnor U16480 (N_16480,N_15371,N_15187);
nand U16481 (N_16481,N_15576,N_15398);
nand U16482 (N_16482,N_15221,N_15829);
or U16483 (N_16483,N_15704,N_15883);
or U16484 (N_16484,N_15535,N_15869);
and U16485 (N_16485,N_15758,N_15621);
nor U16486 (N_16486,N_15178,N_15823);
and U16487 (N_16487,N_15497,N_15613);
or U16488 (N_16488,N_15844,N_15827);
and U16489 (N_16489,N_15899,N_15724);
xnor U16490 (N_16490,N_15970,N_15860);
xor U16491 (N_16491,N_15569,N_15360);
nand U16492 (N_16492,N_15455,N_15342);
and U16493 (N_16493,N_15131,N_15322);
and U16494 (N_16494,N_15267,N_15952);
nand U16495 (N_16495,N_15833,N_15465);
nor U16496 (N_16496,N_15437,N_15212);
nor U16497 (N_16497,N_15893,N_15917);
or U16498 (N_16498,N_15713,N_15071);
nor U16499 (N_16499,N_15145,N_15889);
or U16500 (N_16500,N_15923,N_15573);
nand U16501 (N_16501,N_15248,N_15425);
or U16502 (N_16502,N_15628,N_15900);
and U16503 (N_16503,N_15083,N_15599);
nor U16504 (N_16504,N_15455,N_15369);
nor U16505 (N_16505,N_15466,N_15330);
or U16506 (N_16506,N_15739,N_15532);
xnor U16507 (N_16507,N_15712,N_15310);
xnor U16508 (N_16508,N_15512,N_15012);
nor U16509 (N_16509,N_15709,N_15794);
nand U16510 (N_16510,N_15168,N_15515);
nor U16511 (N_16511,N_15471,N_15397);
nor U16512 (N_16512,N_15722,N_15477);
nor U16513 (N_16513,N_15445,N_15840);
nor U16514 (N_16514,N_15185,N_15534);
nand U16515 (N_16515,N_15049,N_15118);
and U16516 (N_16516,N_15715,N_15245);
nand U16517 (N_16517,N_15907,N_15476);
nor U16518 (N_16518,N_15079,N_15446);
xnor U16519 (N_16519,N_15141,N_15011);
nor U16520 (N_16520,N_15120,N_15780);
nand U16521 (N_16521,N_15620,N_15501);
nor U16522 (N_16522,N_15735,N_15410);
or U16523 (N_16523,N_15976,N_15090);
or U16524 (N_16524,N_15537,N_15925);
xnor U16525 (N_16525,N_15486,N_15896);
nor U16526 (N_16526,N_15089,N_15298);
and U16527 (N_16527,N_15391,N_15014);
nor U16528 (N_16528,N_15893,N_15963);
nor U16529 (N_16529,N_15356,N_15145);
nor U16530 (N_16530,N_15122,N_15802);
xor U16531 (N_16531,N_15553,N_15286);
nor U16532 (N_16532,N_15665,N_15838);
nand U16533 (N_16533,N_15772,N_15274);
or U16534 (N_16534,N_15327,N_15851);
or U16535 (N_16535,N_15621,N_15973);
and U16536 (N_16536,N_15653,N_15582);
and U16537 (N_16537,N_15251,N_15378);
nand U16538 (N_16538,N_15248,N_15721);
xnor U16539 (N_16539,N_15869,N_15658);
nand U16540 (N_16540,N_15100,N_15666);
nand U16541 (N_16541,N_15474,N_15608);
nand U16542 (N_16542,N_15845,N_15835);
nor U16543 (N_16543,N_15547,N_15677);
and U16544 (N_16544,N_15297,N_15806);
xor U16545 (N_16545,N_15320,N_15690);
nor U16546 (N_16546,N_15110,N_15950);
nor U16547 (N_16547,N_15085,N_15686);
nand U16548 (N_16548,N_15205,N_15871);
nand U16549 (N_16549,N_15072,N_15150);
or U16550 (N_16550,N_15454,N_15720);
and U16551 (N_16551,N_15026,N_15533);
or U16552 (N_16552,N_15233,N_15071);
and U16553 (N_16553,N_15732,N_15237);
xnor U16554 (N_16554,N_15388,N_15861);
xnor U16555 (N_16555,N_15323,N_15332);
xnor U16556 (N_16556,N_15302,N_15697);
or U16557 (N_16557,N_15861,N_15792);
nand U16558 (N_16558,N_15137,N_15544);
nor U16559 (N_16559,N_15399,N_15085);
and U16560 (N_16560,N_15916,N_15358);
xnor U16561 (N_16561,N_15618,N_15712);
nand U16562 (N_16562,N_15187,N_15839);
and U16563 (N_16563,N_15353,N_15304);
or U16564 (N_16564,N_15460,N_15791);
nand U16565 (N_16565,N_15591,N_15780);
and U16566 (N_16566,N_15338,N_15679);
and U16567 (N_16567,N_15992,N_15559);
and U16568 (N_16568,N_15516,N_15407);
nand U16569 (N_16569,N_15648,N_15711);
nor U16570 (N_16570,N_15637,N_15235);
or U16571 (N_16571,N_15142,N_15651);
and U16572 (N_16572,N_15736,N_15400);
and U16573 (N_16573,N_15360,N_15183);
xor U16574 (N_16574,N_15946,N_15248);
or U16575 (N_16575,N_15023,N_15558);
xor U16576 (N_16576,N_15539,N_15029);
and U16577 (N_16577,N_15136,N_15941);
xor U16578 (N_16578,N_15762,N_15030);
or U16579 (N_16579,N_15605,N_15596);
xnor U16580 (N_16580,N_15312,N_15458);
nor U16581 (N_16581,N_15416,N_15680);
or U16582 (N_16582,N_15423,N_15472);
nand U16583 (N_16583,N_15907,N_15306);
xnor U16584 (N_16584,N_15243,N_15044);
nor U16585 (N_16585,N_15435,N_15495);
nand U16586 (N_16586,N_15189,N_15661);
xor U16587 (N_16587,N_15375,N_15131);
xor U16588 (N_16588,N_15925,N_15210);
nor U16589 (N_16589,N_15797,N_15219);
nor U16590 (N_16590,N_15883,N_15081);
and U16591 (N_16591,N_15864,N_15616);
and U16592 (N_16592,N_15338,N_15562);
xnor U16593 (N_16593,N_15889,N_15852);
or U16594 (N_16594,N_15955,N_15952);
nand U16595 (N_16595,N_15912,N_15190);
nand U16596 (N_16596,N_15158,N_15257);
xor U16597 (N_16597,N_15978,N_15608);
and U16598 (N_16598,N_15345,N_15492);
nand U16599 (N_16599,N_15254,N_15493);
or U16600 (N_16600,N_15736,N_15809);
or U16601 (N_16601,N_15392,N_15571);
and U16602 (N_16602,N_15016,N_15779);
or U16603 (N_16603,N_15464,N_15006);
xnor U16604 (N_16604,N_15948,N_15840);
nor U16605 (N_16605,N_15765,N_15088);
nor U16606 (N_16606,N_15767,N_15859);
xnor U16607 (N_16607,N_15210,N_15138);
and U16608 (N_16608,N_15556,N_15312);
nor U16609 (N_16609,N_15298,N_15783);
nor U16610 (N_16610,N_15868,N_15820);
nor U16611 (N_16611,N_15837,N_15099);
nor U16612 (N_16612,N_15625,N_15438);
and U16613 (N_16613,N_15418,N_15650);
nand U16614 (N_16614,N_15760,N_15470);
or U16615 (N_16615,N_15696,N_15086);
and U16616 (N_16616,N_15476,N_15635);
and U16617 (N_16617,N_15453,N_15426);
nor U16618 (N_16618,N_15589,N_15420);
nand U16619 (N_16619,N_15565,N_15743);
nand U16620 (N_16620,N_15157,N_15908);
nor U16621 (N_16621,N_15597,N_15241);
nor U16622 (N_16622,N_15114,N_15711);
xor U16623 (N_16623,N_15059,N_15067);
nor U16624 (N_16624,N_15996,N_15840);
nand U16625 (N_16625,N_15496,N_15697);
nor U16626 (N_16626,N_15234,N_15646);
xnor U16627 (N_16627,N_15534,N_15968);
xor U16628 (N_16628,N_15542,N_15089);
and U16629 (N_16629,N_15283,N_15821);
and U16630 (N_16630,N_15726,N_15767);
and U16631 (N_16631,N_15388,N_15009);
nand U16632 (N_16632,N_15959,N_15685);
nor U16633 (N_16633,N_15918,N_15946);
nor U16634 (N_16634,N_15934,N_15229);
and U16635 (N_16635,N_15258,N_15905);
nor U16636 (N_16636,N_15798,N_15501);
xnor U16637 (N_16637,N_15729,N_15031);
and U16638 (N_16638,N_15406,N_15313);
or U16639 (N_16639,N_15781,N_15008);
or U16640 (N_16640,N_15212,N_15419);
and U16641 (N_16641,N_15401,N_15092);
and U16642 (N_16642,N_15074,N_15221);
and U16643 (N_16643,N_15903,N_15791);
nand U16644 (N_16644,N_15292,N_15062);
nand U16645 (N_16645,N_15079,N_15679);
or U16646 (N_16646,N_15417,N_15280);
nand U16647 (N_16647,N_15138,N_15845);
nor U16648 (N_16648,N_15702,N_15930);
and U16649 (N_16649,N_15686,N_15187);
nand U16650 (N_16650,N_15970,N_15675);
nand U16651 (N_16651,N_15411,N_15791);
and U16652 (N_16652,N_15477,N_15508);
xnor U16653 (N_16653,N_15132,N_15046);
and U16654 (N_16654,N_15996,N_15100);
nand U16655 (N_16655,N_15088,N_15075);
or U16656 (N_16656,N_15493,N_15808);
xor U16657 (N_16657,N_15197,N_15880);
nand U16658 (N_16658,N_15797,N_15103);
and U16659 (N_16659,N_15846,N_15445);
nor U16660 (N_16660,N_15491,N_15754);
xnor U16661 (N_16661,N_15734,N_15027);
or U16662 (N_16662,N_15482,N_15119);
nor U16663 (N_16663,N_15645,N_15466);
nand U16664 (N_16664,N_15163,N_15702);
or U16665 (N_16665,N_15855,N_15070);
nand U16666 (N_16666,N_15795,N_15556);
and U16667 (N_16667,N_15866,N_15558);
or U16668 (N_16668,N_15051,N_15660);
nand U16669 (N_16669,N_15359,N_15388);
nand U16670 (N_16670,N_15710,N_15408);
nand U16671 (N_16671,N_15420,N_15239);
nand U16672 (N_16672,N_15793,N_15425);
or U16673 (N_16673,N_15747,N_15155);
xnor U16674 (N_16674,N_15904,N_15042);
nor U16675 (N_16675,N_15183,N_15169);
or U16676 (N_16676,N_15091,N_15331);
and U16677 (N_16677,N_15394,N_15867);
or U16678 (N_16678,N_15641,N_15799);
and U16679 (N_16679,N_15995,N_15735);
xor U16680 (N_16680,N_15734,N_15143);
nor U16681 (N_16681,N_15940,N_15073);
nor U16682 (N_16682,N_15929,N_15480);
nor U16683 (N_16683,N_15794,N_15166);
and U16684 (N_16684,N_15932,N_15520);
nor U16685 (N_16685,N_15951,N_15692);
and U16686 (N_16686,N_15326,N_15054);
nand U16687 (N_16687,N_15028,N_15273);
nand U16688 (N_16688,N_15133,N_15306);
nand U16689 (N_16689,N_15404,N_15006);
nor U16690 (N_16690,N_15892,N_15186);
xor U16691 (N_16691,N_15063,N_15089);
xor U16692 (N_16692,N_15821,N_15600);
nand U16693 (N_16693,N_15517,N_15848);
nor U16694 (N_16694,N_15009,N_15754);
or U16695 (N_16695,N_15071,N_15306);
nand U16696 (N_16696,N_15227,N_15279);
and U16697 (N_16697,N_15786,N_15580);
xor U16698 (N_16698,N_15023,N_15915);
or U16699 (N_16699,N_15504,N_15413);
xor U16700 (N_16700,N_15756,N_15819);
xnor U16701 (N_16701,N_15934,N_15912);
and U16702 (N_16702,N_15839,N_15675);
and U16703 (N_16703,N_15846,N_15066);
or U16704 (N_16704,N_15227,N_15748);
nand U16705 (N_16705,N_15888,N_15916);
nor U16706 (N_16706,N_15567,N_15391);
nand U16707 (N_16707,N_15481,N_15006);
and U16708 (N_16708,N_15280,N_15271);
nor U16709 (N_16709,N_15975,N_15644);
or U16710 (N_16710,N_15680,N_15206);
xor U16711 (N_16711,N_15527,N_15467);
nor U16712 (N_16712,N_15040,N_15017);
nand U16713 (N_16713,N_15985,N_15356);
or U16714 (N_16714,N_15042,N_15524);
and U16715 (N_16715,N_15307,N_15226);
or U16716 (N_16716,N_15411,N_15318);
xor U16717 (N_16717,N_15517,N_15103);
or U16718 (N_16718,N_15288,N_15017);
and U16719 (N_16719,N_15403,N_15515);
and U16720 (N_16720,N_15316,N_15160);
or U16721 (N_16721,N_15494,N_15019);
and U16722 (N_16722,N_15900,N_15370);
nor U16723 (N_16723,N_15574,N_15995);
and U16724 (N_16724,N_15943,N_15200);
nand U16725 (N_16725,N_15944,N_15349);
and U16726 (N_16726,N_15736,N_15707);
nor U16727 (N_16727,N_15945,N_15671);
nor U16728 (N_16728,N_15657,N_15030);
or U16729 (N_16729,N_15041,N_15882);
xnor U16730 (N_16730,N_15435,N_15224);
or U16731 (N_16731,N_15740,N_15092);
nand U16732 (N_16732,N_15984,N_15012);
and U16733 (N_16733,N_15809,N_15899);
or U16734 (N_16734,N_15291,N_15455);
and U16735 (N_16735,N_15166,N_15640);
nand U16736 (N_16736,N_15392,N_15237);
nor U16737 (N_16737,N_15430,N_15310);
xor U16738 (N_16738,N_15860,N_15688);
xnor U16739 (N_16739,N_15518,N_15475);
nor U16740 (N_16740,N_15332,N_15156);
nand U16741 (N_16741,N_15199,N_15327);
or U16742 (N_16742,N_15208,N_15071);
and U16743 (N_16743,N_15582,N_15853);
xnor U16744 (N_16744,N_15986,N_15816);
xnor U16745 (N_16745,N_15171,N_15114);
xnor U16746 (N_16746,N_15734,N_15235);
and U16747 (N_16747,N_15572,N_15463);
nor U16748 (N_16748,N_15211,N_15472);
or U16749 (N_16749,N_15416,N_15992);
nand U16750 (N_16750,N_15543,N_15456);
xnor U16751 (N_16751,N_15803,N_15632);
nand U16752 (N_16752,N_15726,N_15774);
nor U16753 (N_16753,N_15523,N_15916);
nor U16754 (N_16754,N_15520,N_15402);
and U16755 (N_16755,N_15887,N_15803);
and U16756 (N_16756,N_15250,N_15353);
xor U16757 (N_16757,N_15863,N_15926);
xor U16758 (N_16758,N_15920,N_15553);
xor U16759 (N_16759,N_15981,N_15144);
xnor U16760 (N_16760,N_15456,N_15064);
and U16761 (N_16761,N_15944,N_15188);
nor U16762 (N_16762,N_15451,N_15815);
and U16763 (N_16763,N_15412,N_15995);
and U16764 (N_16764,N_15750,N_15128);
xnor U16765 (N_16765,N_15037,N_15175);
and U16766 (N_16766,N_15401,N_15417);
nor U16767 (N_16767,N_15869,N_15115);
and U16768 (N_16768,N_15020,N_15462);
nor U16769 (N_16769,N_15923,N_15237);
and U16770 (N_16770,N_15520,N_15092);
xnor U16771 (N_16771,N_15647,N_15384);
nor U16772 (N_16772,N_15245,N_15173);
or U16773 (N_16773,N_15108,N_15185);
and U16774 (N_16774,N_15192,N_15585);
xor U16775 (N_16775,N_15972,N_15137);
xor U16776 (N_16776,N_15881,N_15701);
or U16777 (N_16777,N_15814,N_15733);
or U16778 (N_16778,N_15172,N_15921);
nor U16779 (N_16779,N_15653,N_15300);
xor U16780 (N_16780,N_15797,N_15296);
and U16781 (N_16781,N_15028,N_15463);
and U16782 (N_16782,N_15526,N_15881);
and U16783 (N_16783,N_15534,N_15323);
or U16784 (N_16784,N_15879,N_15853);
or U16785 (N_16785,N_15656,N_15677);
and U16786 (N_16786,N_15392,N_15609);
xnor U16787 (N_16787,N_15172,N_15851);
or U16788 (N_16788,N_15315,N_15959);
and U16789 (N_16789,N_15007,N_15411);
and U16790 (N_16790,N_15029,N_15419);
and U16791 (N_16791,N_15559,N_15453);
and U16792 (N_16792,N_15823,N_15917);
and U16793 (N_16793,N_15319,N_15912);
and U16794 (N_16794,N_15321,N_15572);
nand U16795 (N_16795,N_15985,N_15286);
nand U16796 (N_16796,N_15997,N_15826);
xnor U16797 (N_16797,N_15873,N_15339);
nand U16798 (N_16798,N_15823,N_15167);
and U16799 (N_16799,N_15416,N_15534);
nor U16800 (N_16800,N_15717,N_15445);
and U16801 (N_16801,N_15477,N_15233);
and U16802 (N_16802,N_15658,N_15094);
and U16803 (N_16803,N_15758,N_15372);
nor U16804 (N_16804,N_15131,N_15152);
nor U16805 (N_16805,N_15750,N_15114);
nor U16806 (N_16806,N_15857,N_15109);
nand U16807 (N_16807,N_15341,N_15703);
and U16808 (N_16808,N_15070,N_15875);
and U16809 (N_16809,N_15218,N_15688);
or U16810 (N_16810,N_15241,N_15529);
and U16811 (N_16811,N_15914,N_15307);
xor U16812 (N_16812,N_15044,N_15999);
nand U16813 (N_16813,N_15643,N_15756);
and U16814 (N_16814,N_15912,N_15480);
or U16815 (N_16815,N_15344,N_15976);
or U16816 (N_16816,N_15656,N_15569);
nor U16817 (N_16817,N_15829,N_15849);
and U16818 (N_16818,N_15367,N_15541);
nor U16819 (N_16819,N_15332,N_15438);
nand U16820 (N_16820,N_15071,N_15729);
and U16821 (N_16821,N_15601,N_15498);
and U16822 (N_16822,N_15968,N_15833);
nand U16823 (N_16823,N_15219,N_15967);
nand U16824 (N_16824,N_15807,N_15501);
or U16825 (N_16825,N_15864,N_15635);
or U16826 (N_16826,N_15971,N_15352);
or U16827 (N_16827,N_15430,N_15933);
xor U16828 (N_16828,N_15090,N_15517);
nand U16829 (N_16829,N_15140,N_15063);
nand U16830 (N_16830,N_15462,N_15069);
xnor U16831 (N_16831,N_15966,N_15858);
nand U16832 (N_16832,N_15069,N_15436);
nor U16833 (N_16833,N_15938,N_15455);
nor U16834 (N_16834,N_15698,N_15902);
nor U16835 (N_16835,N_15495,N_15843);
or U16836 (N_16836,N_15448,N_15564);
and U16837 (N_16837,N_15155,N_15454);
and U16838 (N_16838,N_15583,N_15590);
and U16839 (N_16839,N_15809,N_15898);
and U16840 (N_16840,N_15870,N_15853);
xnor U16841 (N_16841,N_15697,N_15191);
and U16842 (N_16842,N_15538,N_15243);
nor U16843 (N_16843,N_15430,N_15116);
or U16844 (N_16844,N_15429,N_15917);
or U16845 (N_16845,N_15533,N_15050);
xnor U16846 (N_16846,N_15194,N_15491);
nor U16847 (N_16847,N_15679,N_15326);
and U16848 (N_16848,N_15256,N_15102);
nand U16849 (N_16849,N_15618,N_15858);
or U16850 (N_16850,N_15302,N_15719);
xnor U16851 (N_16851,N_15886,N_15233);
xnor U16852 (N_16852,N_15515,N_15558);
nand U16853 (N_16853,N_15302,N_15263);
nand U16854 (N_16854,N_15039,N_15464);
and U16855 (N_16855,N_15897,N_15970);
nor U16856 (N_16856,N_15800,N_15968);
xor U16857 (N_16857,N_15202,N_15298);
nand U16858 (N_16858,N_15833,N_15536);
xnor U16859 (N_16859,N_15205,N_15156);
xor U16860 (N_16860,N_15597,N_15722);
xor U16861 (N_16861,N_15236,N_15953);
nor U16862 (N_16862,N_15330,N_15282);
xnor U16863 (N_16863,N_15577,N_15757);
nor U16864 (N_16864,N_15585,N_15793);
nor U16865 (N_16865,N_15814,N_15450);
nand U16866 (N_16866,N_15320,N_15848);
nor U16867 (N_16867,N_15231,N_15924);
xor U16868 (N_16868,N_15983,N_15674);
nand U16869 (N_16869,N_15740,N_15914);
and U16870 (N_16870,N_15499,N_15590);
xnor U16871 (N_16871,N_15148,N_15365);
and U16872 (N_16872,N_15421,N_15874);
or U16873 (N_16873,N_15238,N_15799);
nand U16874 (N_16874,N_15148,N_15420);
nand U16875 (N_16875,N_15783,N_15654);
xnor U16876 (N_16876,N_15558,N_15119);
xor U16877 (N_16877,N_15633,N_15677);
nand U16878 (N_16878,N_15890,N_15194);
xor U16879 (N_16879,N_15891,N_15077);
and U16880 (N_16880,N_15668,N_15360);
or U16881 (N_16881,N_15935,N_15215);
xnor U16882 (N_16882,N_15789,N_15139);
nor U16883 (N_16883,N_15209,N_15508);
nand U16884 (N_16884,N_15662,N_15380);
or U16885 (N_16885,N_15819,N_15680);
xnor U16886 (N_16886,N_15122,N_15765);
nand U16887 (N_16887,N_15676,N_15000);
xor U16888 (N_16888,N_15267,N_15857);
nor U16889 (N_16889,N_15334,N_15015);
xnor U16890 (N_16890,N_15590,N_15584);
xor U16891 (N_16891,N_15496,N_15329);
nor U16892 (N_16892,N_15496,N_15767);
or U16893 (N_16893,N_15851,N_15474);
xnor U16894 (N_16894,N_15583,N_15679);
nor U16895 (N_16895,N_15566,N_15319);
or U16896 (N_16896,N_15328,N_15060);
xnor U16897 (N_16897,N_15832,N_15467);
and U16898 (N_16898,N_15564,N_15907);
nand U16899 (N_16899,N_15694,N_15500);
nor U16900 (N_16900,N_15881,N_15015);
nor U16901 (N_16901,N_15496,N_15317);
xnor U16902 (N_16902,N_15986,N_15755);
nor U16903 (N_16903,N_15879,N_15046);
and U16904 (N_16904,N_15487,N_15890);
nor U16905 (N_16905,N_15303,N_15857);
nor U16906 (N_16906,N_15094,N_15113);
nand U16907 (N_16907,N_15710,N_15224);
xnor U16908 (N_16908,N_15065,N_15563);
nor U16909 (N_16909,N_15709,N_15344);
xor U16910 (N_16910,N_15638,N_15929);
nor U16911 (N_16911,N_15638,N_15827);
xnor U16912 (N_16912,N_15477,N_15823);
or U16913 (N_16913,N_15549,N_15463);
nand U16914 (N_16914,N_15417,N_15459);
nand U16915 (N_16915,N_15681,N_15398);
or U16916 (N_16916,N_15903,N_15984);
or U16917 (N_16917,N_15321,N_15566);
or U16918 (N_16918,N_15828,N_15508);
nand U16919 (N_16919,N_15166,N_15193);
and U16920 (N_16920,N_15731,N_15612);
or U16921 (N_16921,N_15995,N_15822);
nor U16922 (N_16922,N_15963,N_15952);
xor U16923 (N_16923,N_15722,N_15185);
nor U16924 (N_16924,N_15576,N_15160);
and U16925 (N_16925,N_15750,N_15373);
nor U16926 (N_16926,N_15209,N_15315);
nor U16927 (N_16927,N_15011,N_15810);
xor U16928 (N_16928,N_15376,N_15937);
xnor U16929 (N_16929,N_15557,N_15042);
nand U16930 (N_16930,N_15071,N_15239);
or U16931 (N_16931,N_15407,N_15853);
or U16932 (N_16932,N_15923,N_15409);
nand U16933 (N_16933,N_15362,N_15156);
nor U16934 (N_16934,N_15893,N_15157);
or U16935 (N_16935,N_15594,N_15159);
or U16936 (N_16936,N_15312,N_15986);
and U16937 (N_16937,N_15866,N_15091);
and U16938 (N_16938,N_15924,N_15370);
xnor U16939 (N_16939,N_15811,N_15703);
nor U16940 (N_16940,N_15348,N_15742);
nand U16941 (N_16941,N_15538,N_15219);
nor U16942 (N_16942,N_15989,N_15911);
or U16943 (N_16943,N_15322,N_15375);
and U16944 (N_16944,N_15692,N_15915);
xor U16945 (N_16945,N_15879,N_15014);
nand U16946 (N_16946,N_15443,N_15319);
nand U16947 (N_16947,N_15919,N_15745);
or U16948 (N_16948,N_15694,N_15587);
and U16949 (N_16949,N_15675,N_15976);
and U16950 (N_16950,N_15462,N_15213);
or U16951 (N_16951,N_15524,N_15716);
or U16952 (N_16952,N_15129,N_15999);
and U16953 (N_16953,N_15286,N_15113);
nand U16954 (N_16954,N_15663,N_15215);
or U16955 (N_16955,N_15631,N_15797);
and U16956 (N_16956,N_15848,N_15943);
or U16957 (N_16957,N_15022,N_15522);
xor U16958 (N_16958,N_15437,N_15714);
nor U16959 (N_16959,N_15678,N_15578);
nor U16960 (N_16960,N_15014,N_15578);
and U16961 (N_16961,N_15675,N_15296);
nor U16962 (N_16962,N_15684,N_15609);
nand U16963 (N_16963,N_15452,N_15685);
or U16964 (N_16964,N_15154,N_15840);
nor U16965 (N_16965,N_15208,N_15603);
and U16966 (N_16966,N_15993,N_15216);
xnor U16967 (N_16967,N_15725,N_15041);
or U16968 (N_16968,N_15982,N_15059);
or U16969 (N_16969,N_15060,N_15843);
xor U16970 (N_16970,N_15455,N_15461);
xnor U16971 (N_16971,N_15066,N_15776);
xor U16972 (N_16972,N_15649,N_15546);
and U16973 (N_16973,N_15699,N_15055);
or U16974 (N_16974,N_15758,N_15131);
nor U16975 (N_16975,N_15914,N_15393);
xor U16976 (N_16976,N_15846,N_15702);
or U16977 (N_16977,N_15969,N_15990);
nand U16978 (N_16978,N_15707,N_15346);
nor U16979 (N_16979,N_15343,N_15379);
nor U16980 (N_16980,N_15971,N_15486);
nor U16981 (N_16981,N_15923,N_15842);
nor U16982 (N_16982,N_15162,N_15690);
nand U16983 (N_16983,N_15095,N_15778);
xnor U16984 (N_16984,N_15118,N_15207);
and U16985 (N_16985,N_15380,N_15810);
nor U16986 (N_16986,N_15645,N_15476);
nand U16987 (N_16987,N_15025,N_15356);
nand U16988 (N_16988,N_15783,N_15450);
nand U16989 (N_16989,N_15212,N_15836);
xor U16990 (N_16990,N_15855,N_15847);
or U16991 (N_16991,N_15744,N_15657);
nor U16992 (N_16992,N_15441,N_15404);
and U16993 (N_16993,N_15002,N_15284);
or U16994 (N_16994,N_15673,N_15185);
nand U16995 (N_16995,N_15427,N_15903);
nand U16996 (N_16996,N_15543,N_15915);
nand U16997 (N_16997,N_15352,N_15053);
nand U16998 (N_16998,N_15541,N_15872);
nand U16999 (N_16999,N_15288,N_15743);
nor U17000 (N_17000,N_16554,N_16353);
or U17001 (N_17001,N_16146,N_16297);
xnor U17002 (N_17002,N_16153,N_16439);
and U17003 (N_17003,N_16056,N_16018);
and U17004 (N_17004,N_16227,N_16148);
xnor U17005 (N_17005,N_16071,N_16529);
nand U17006 (N_17006,N_16396,N_16995);
xnor U17007 (N_17007,N_16425,N_16285);
nand U17008 (N_17008,N_16670,N_16752);
xor U17009 (N_17009,N_16631,N_16026);
nand U17010 (N_17010,N_16009,N_16973);
nand U17011 (N_17011,N_16103,N_16940);
xor U17012 (N_17012,N_16731,N_16773);
nand U17013 (N_17013,N_16151,N_16900);
nand U17014 (N_17014,N_16790,N_16958);
or U17015 (N_17015,N_16339,N_16524);
nor U17016 (N_17016,N_16345,N_16219);
nor U17017 (N_17017,N_16022,N_16276);
nor U17018 (N_17018,N_16555,N_16216);
xnor U17019 (N_17019,N_16336,N_16901);
nor U17020 (N_17020,N_16804,N_16789);
or U17021 (N_17021,N_16762,N_16064);
xnor U17022 (N_17022,N_16992,N_16451);
or U17023 (N_17023,N_16122,N_16182);
or U17024 (N_17024,N_16570,N_16826);
nor U17025 (N_17025,N_16659,N_16728);
nor U17026 (N_17026,N_16539,N_16948);
nand U17027 (N_17027,N_16200,N_16473);
nor U17028 (N_17028,N_16419,N_16602);
and U17029 (N_17029,N_16431,N_16787);
nor U17030 (N_17030,N_16976,N_16552);
or U17031 (N_17031,N_16646,N_16880);
and U17032 (N_17032,N_16034,N_16202);
and U17033 (N_17033,N_16263,N_16145);
and U17034 (N_17034,N_16512,N_16622);
nor U17035 (N_17035,N_16126,N_16320);
nor U17036 (N_17036,N_16073,N_16831);
nand U17037 (N_17037,N_16447,N_16575);
or U17038 (N_17038,N_16290,N_16137);
xnor U17039 (N_17039,N_16315,N_16028);
or U17040 (N_17040,N_16993,N_16438);
or U17041 (N_17041,N_16326,N_16716);
nand U17042 (N_17042,N_16189,N_16070);
xor U17043 (N_17043,N_16489,N_16827);
xor U17044 (N_17044,N_16531,N_16635);
and U17045 (N_17045,N_16767,N_16763);
and U17046 (N_17046,N_16113,N_16400);
nor U17047 (N_17047,N_16371,N_16311);
xor U17048 (N_17048,N_16818,N_16382);
nand U17049 (N_17049,N_16803,N_16810);
nand U17050 (N_17050,N_16864,N_16820);
xnor U17051 (N_17051,N_16896,N_16696);
nand U17052 (N_17052,N_16463,N_16641);
nand U17053 (N_17053,N_16332,N_16292);
or U17054 (N_17054,N_16330,N_16185);
and U17055 (N_17055,N_16709,N_16015);
or U17056 (N_17056,N_16475,N_16576);
and U17057 (N_17057,N_16331,N_16746);
and U17058 (N_17058,N_16091,N_16893);
or U17059 (N_17059,N_16328,N_16538);
and U17060 (N_17060,N_16230,N_16727);
nand U17061 (N_17061,N_16847,N_16055);
nand U17062 (N_17062,N_16526,N_16777);
xor U17063 (N_17063,N_16933,N_16887);
nor U17064 (N_17064,N_16406,N_16164);
or U17065 (N_17065,N_16736,N_16180);
xnor U17066 (N_17066,N_16032,N_16037);
and U17067 (N_17067,N_16983,N_16193);
and U17068 (N_17068,N_16996,N_16249);
or U17069 (N_17069,N_16187,N_16490);
or U17070 (N_17070,N_16387,N_16742);
nor U17071 (N_17071,N_16421,N_16237);
nand U17072 (N_17072,N_16749,N_16944);
nor U17073 (N_17073,N_16344,N_16652);
nand U17074 (N_17074,N_16825,N_16204);
and U17075 (N_17075,N_16255,N_16945);
nand U17076 (N_17076,N_16444,N_16912);
or U17077 (N_17077,N_16318,N_16341);
or U17078 (N_17078,N_16160,N_16173);
nor U17079 (N_17079,N_16197,N_16136);
or U17080 (N_17080,N_16691,N_16250);
xor U17081 (N_17081,N_16981,N_16239);
or U17082 (N_17082,N_16074,N_16140);
and U17083 (N_17083,N_16050,N_16934);
nor U17084 (N_17084,N_16468,N_16523);
or U17085 (N_17085,N_16482,N_16288);
xor U17086 (N_17086,N_16618,N_16700);
xnor U17087 (N_17087,N_16929,N_16969);
nor U17088 (N_17088,N_16596,N_16205);
and U17089 (N_17089,N_16017,N_16726);
or U17090 (N_17090,N_16172,N_16747);
nor U17091 (N_17091,N_16310,N_16886);
nor U17092 (N_17092,N_16422,N_16395);
and U17093 (N_17093,N_16201,N_16918);
and U17094 (N_17094,N_16407,N_16319);
nor U17095 (N_17095,N_16333,N_16133);
or U17096 (N_17096,N_16066,N_16503);
or U17097 (N_17097,N_16874,N_16054);
and U17098 (N_17098,N_16838,N_16919);
and U17099 (N_17099,N_16356,N_16672);
and U17100 (N_17100,N_16351,N_16931);
and U17101 (N_17101,N_16540,N_16571);
nor U17102 (N_17102,N_16049,N_16008);
and U17103 (N_17103,N_16725,N_16279);
and U17104 (N_17104,N_16653,N_16678);
and U17105 (N_17105,N_16461,N_16507);
and U17106 (N_17106,N_16951,N_16980);
nor U17107 (N_17107,N_16184,N_16927);
nor U17108 (N_17108,N_16303,N_16433);
and U17109 (N_17109,N_16398,N_16513);
or U17110 (N_17110,N_16495,N_16355);
and U17111 (N_17111,N_16553,N_16680);
and U17112 (N_17112,N_16175,N_16590);
or U17113 (N_17113,N_16664,N_16624);
nand U17114 (N_17114,N_16634,N_16591);
nor U17115 (N_17115,N_16248,N_16761);
nand U17116 (N_17116,N_16440,N_16217);
nor U17117 (N_17117,N_16636,N_16010);
nor U17118 (N_17118,N_16785,N_16308);
nand U17119 (N_17119,N_16446,N_16102);
xor U17120 (N_17120,N_16480,N_16990);
xor U17121 (N_17121,N_16892,N_16501);
xnor U17122 (N_17122,N_16504,N_16774);
xnor U17123 (N_17123,N_16264,N_16242);
xnor U17124 (N_17124,N_16394,N_16615);
nand U17125 (N_17125,N_16967,N_16510);
xnor U17126 (N_17126,N_16915,N_16581);
or U17127 (N_17127,N_16645,N_16038);
nand U17128 (N_17128,N_16267,N_16417);
nor U17129 (N_17129,N_16956,N_16930);
and U17130 (N_17130,N_16844,N_16679);
xor U17131 (N_17131,N_16550,N_16284);
or U17132 (N_17132,N_16724,N_16890);
and U17133 (N_17133,N_16506,N_16152);
nand U17134 (N_17134,N_16100,N_16030);
and U17135 (N_17135,N_16542,N_16701);
and U17136 (N_17136,N_16648,N_16130);
or U17137 (N_17137,N_16706,N_16358);
and U17138 (N_17138,N_16003,N_16532);
xnor U17139 (N_17139,N_16920,N_16499);
and U17140 (N_17140,N_16690,N_16765);
or U17141 (N_17141,N_16220,N_16610);
nor U17142 (N_17142,N_16546,N_16595);
nor U17143 (N_17143,N_16748,N_16174);
and U17144 (N_17144,N_16138,N_16357);
or U17145 (N_17145,N_16042,N_16023);
xor U17146 (N_17146,N_16223,N_16085);
nor U17147 (N_17147,N_16535,N_16092);
nor U17148 (N_17148,N_16982,N_16637);
or U17149 (N_17149,N_16206,N_16380);
nor U17150 (N_17150,N_16077,N_16739);
nand U17151 (N_17151,N_16561,N_16278);
and U17152 (N_17152,N_16830,N_16608);
or U17153 (N_17153,N_16729,N_16271);
nor U17154 (N_17154,N_16177,N_16161);
xnor U17155 (N_17155,N_16083,N_16839);
nor U17156 (N_17156,N_16572,N_16514);
nor U17157 (N_17157,N_16817,N_16882);
nand U17158 (N_17158,N_16041,N_16178);
xnor U17159 (N_17159,N_16620,N_16655);
or U17160 (N_17160,N_16386,N_16587);
and U17161 (N_17161,N_16738,N_16462);
and U17162 (N_17162,N_16135,N_16006);
or U17163 (N_17163,N_16238,N_16094);
and U17164 (N_17164,N_16467,N_16883);
and U17165 (N_17165,N_16604,N_16335);
nor U17166 (N_17166,N_16031,N_16941);
nand U17167 (N_17167,N_16169,N_16585);
nand U17168 (N_17168,N_16340,N_16894);
nor U17169 (N_17169,N_16511,N_16361);
and U17170 (N_17170,N_16757,N_16708);
nand U17171 (N_17171,N_16589,N_16835);
xnor U17172 (N_17172,N_16811,N_16866);
nor U17173 (N_17173,N_16270,N_16955);
and U17174 (N_17174,N_16833,N_16671);
and U17175 (N_17175,N_16619,N_16296);
and U17176 (N_17176,N_16950,N_16115);
or U17177 (N_17177,N_16300,N_16801);
nor U17178 (N_17178,N_16159,N_16127);
or U17179 (N_17179,N_16280,N_16459);
nand U17180 (N_17180,N_16388,N_16856);
or U17181 (N_17181,N_16832,N_16621);
xnor U17182 (N_17182,N_16859,N_16316);
xnor U17183 (N_17183,N_16163,N_16287);
and U17184 (N_17184,N_16626,N_16128);
nor U17185 (N_17185,N_16409,N_16360);
nand U17186 (N_17186,N_16557,N_16998);
nor U17187 (N_17187,N_16011,N_16613);
nor U17188 (N_17188,N_16989,N_16381);
nor U17189 (N_17189,N_16517,N_16953);
or U17190 (N_17190,N_16377,N_16876);
nand U17191 (N_17191,N_16013,N_16656);
and U17192 (N_17192,N_16669,N_16594);
nor U17193 (N_17193,N_16067,N_16942);
and U17194 (N_17194,N_16014,N_16329);
nand U17195 (N_17195,N_16254,N_16821);
xor U17196 (N_17196,N_16843,N_16166);
nor U17197 (N_17197,N_16865,N_16578);
nand U17198 (N_17198,N_16661,N_16792);
xnor U17199 (N_17199,N_16347,N_16647);
and U17200 (N_17200,N_16699,N_16337);
or U17201 (N_17201,N_16500,N_16755);
and U17202 (N_17202,N_16798,N_16260);
xor U17203 (N_17203,N_16518,N_16564);
nor U17204 (N_17204,N_16171,N_16158);
or U17205 (N_17205,N_16449,N_16858);
nor U17206 (N_17206,N_16226,N_16586);
xnor U17207 (N_17207,N_16952,N_16283);
and U17208 (N_17208,N_16673,N_16805);
and U17209 (N_17209,N_16004,N_16663);
xor U17210 (N_17210,N_16860,N_16139);
nand U17211 (N_17211,N_16352,N_16403);
nor U17212 (N_17212,N_16027,N_16486);
xor U17213 (N_17213,N_16299,N_16640);
or U17214 (N_17214,N_16965,N_16836);
and U17215 (N_17215,N_16307,N_16881);
nand U17216 (N_17216,N_16232,N_16411);
nand U17217 (N_17217,N_16548,N_16134);
or U17218 (N_17218,N_16366,N_16806);
xor U17219 (N_17219,N_16213,N_16157);
nor U17220 (N_17220,N_16574,N_16852);
xor U17221 (N_17221,N_16854,N_16627);
or U17222 (N_17222,N_16051,N_16741);
nand U17223 (N_17223,N_16488,N_16666);
or U17224 (N_17224,N_16412,N_16991);
nand U17225 (N_17225,N_16743,N_16913);
nor U17226 (N_17226,N_16065,N_16099);
and U17227 (N_17227,N_16472,N_16947);
xnor U17228 (N_17228,N_16101,N_16252);
xnor U17229 (N_17229,N_16889,N_16362);
nor U17230 (N_17230,N_16460,N_16181);
nand U17231 (N_17231,N_16251,N_16273);
or U17232 (N_17232,N_16816,N_16730);
and U17233 (N_17233,N_16601,N_16520);
nor U17234 (N_17234,N_16457,N_16118);
nor U17235 (N_17235,N_16676,N_16917);
xor U17236 (N_17236,N_16932,N_16108);
and U17237 (N_17237,N_16001,N_16584);
or U17238 (N_17238,N_16110,N_16740);
xor U17239 (N_17239,N_16168,N_16390);
xnor U17240 (N_17240,N_16667,N_16002);
xnor U17241 (N_17241,N_16097,N_16611);
and U17242 (N_17242,N_16855,N_16095);
xor U17243 (N_17243,N_16734,N_16455);
nand U17244 (N_17244,N_16209,N_16350);
xnor U17245 (N_17245,N_16588,N_16089);
xnor U17246 (N_17246,N_16443,N_16946);
or U17247 (N_17247,N_16849,N_16788);
and U17248 (N_17248,N_16183,N_16176);
and U17249 (N_17249,N_16782,N_16985);
xnor U17250 (N_17250,N_16294,N_16598);
and U17251 (N_17251,N_16469,N_16221);
nor U17252 (N_17252,N_16878,N_16057);
or U17253 (N_17253,N_16541,N_16434);
nand U17254 (N_17254,N_16977,N_16418);
or U17255 (N_17255,N_16824,N_16132);
xor U17256 (N_17256,N_16819,N_16593);
and U17257 (N_17257,N_16979,N_16558);
xor U17258 (N_17258,N_16081,N_16420);
or U17259 (N_17259,N_16210,N_16685);
or U17260 (N_17260,N_16508,N_16605);
nand U17261 (N_17261,N_16428,N_16198);
nor U17262 (N_17262,N_16668,N_16649);
and U17263 (N_17263,N_16687,N_16314);
and U17264 (N_17264,N_16662,N_16046);
xnor U17265 (N_17265,N_16212,N_16907);
xnor U17266 (N_17266,N_16505,N_16104);
xnor U17267 (N_17267,N_16033,N_16978);
nor U17268 (N_17268,N_16342,N_16794);
nor U17269 (N_17269,N_16144,N_16938);
nand U17270 (N_17270,N_16426,N_16703);
or U17271 (N_17271,N_16231,N_16937);
nor U17272 (N_17272,N_16758,N_16705);
nand U17273 (N_17273,N_16987,N_16682);
nor U17274 (N_17274,N_16614,N_16921);
or U17275 (N_17275,N_16309,N_16293);
xor U17276 (N_17276,N_16846,N_16768);
nor U17277 (N_17277,N_16922,N_16246);
nor U17278 (N_17278,N_16391,N_16448);
nand U17279 (N_17279,N_16088,N_16630);
nand U17280 (N_17280,N_16441,N_16923);
nor U17281 (N_17281,N_16688,N_16963);
or U17282 (N_17282,N_16043,N_16650);
and U17283 (N_17283,N_16430,N_16474);
nor U17284 (N_17284,N_16207,N_16327);
or U17285 (N_17285,N_16502,N_16107);
nand U17286 (N_17286,N_16272,N_16975);
and U17287 (N_17287,N_16029,N_16954);
and U17288 (N_17288,N_16791,N_16891);
xor U17289 (N_17289,N_16215,N_16379);
xnor U17290 (N_17290,N_16566,N_16657);
and U17291 (N_17291,N_16737,N_16607);
nand U17292 (N_17292,N_16999,N_16754);
nor U17293 (N_17293,N_16317,N_16225);
or U17294 (N_17294,N_16909,N_16697);
xnor U17295 (N_17295,N_16733,N_16828);
or U17296 (N_17296,N_16735,N_16961);
and U17297 (N_17297,N_16643,N_16568);
xnor U17298 (N_17298,N_16483,N_16924);
or U17299 (N_17299,N_16036,N_16481);
xnor U17300 (N_17300,N_16665,N_16243);
or U17301 (N_17301,N_16905,N_16298);
or U17302 (N_17302,N_16949,N_16075);
and U17303 (N_17303,N_16496,N_16408);
and U17304 (N_17304,N_16367,N_16710);
xnor U17305 (N_17305,N_16244,N_16675);
or U17306 (N_17306,N_16632,N_16452);
and U17307 (N_17307,N_16879,N_16258);
xnor U17308 (N_17308,N_16111,N_16397);
or U17309 (N_17309,N_16764,N_16861);
nor U17310 (N_17310,N_16322,N_16974);
xor U17311 (N_17311,N_16484,N_16405);
or U17312 (N_17312,N_16808,N_16775);
nand U17313 (N_17313,N_16039,N_16208);
nor U17314 (N_17314,N_16052,N_16305);
and U17315 (N_17315,N_16402,N_16714);
nor U17316 (N_17316,N_16143,N_16393);
nand U17317 (N_17317,N_16616,N_16372);
or U17318 (N_17318,N_16131,N_16994);
nand U17319 (N_17319,N_16261,N_16125);
nor U17320 (N_17320,N_16378,N_16025);
and U17321 (N_17321,N_16556,N_16914);
and U17322 (N_17322,N_16848,N_16376);
or U17323 (N_17323,N_16304,N_16899);
and U17324 (N_17324,N_16536,N_16389);
and U17325 (N_17325,N_16257,N_16850);
or U17326 (N_17326,N_16612,N_16698);
nor U17327 (N_17327,N_16302,N_16109);
nand U17328 (N_17328,N_16800,N_16363);
nor U17329 (N_17329,N_16677,N_16245);
nand U17330 (N_17330,N_16119,N_16224);
nor U17331 (N_17331,N_16021,N_16903);
or U17332 (N_17332,N_16493,N_16877);
nand U17333 (N_17333,N_16779,N_16072);
or U17334 (N_17334,N_16943,N_16259);
nor U17335 (N_17335,N_16079,N_16123);
xor U17336 (N_17336,N_16962,N_16851);
xnor U17337 (N_17337,N_16162,N_16603);
nor U17338 (N_17338,N_16957,N_16241);
or U17339 (N_17339,N_16416,N_16718);
nand U17340 (N_17340,N_16684,N_16753);
nor U17341 (N_17341,N_16766,N_16809);
nand U17342 (N_17342,N_16707,N_16199);
xnor U17343 (N_17343,N_16970,N_16194);
or U17344 (N_17344,N_16984,N_16295);
and U17345 (N_17345,N_16547,N_16654);
or U17346 (N_17346,N_16888,N_16885);
and U17347 (N_17347,N_16410,N_16712);
nor U17348 (N_17348,N_16458,N_16549);
and U17349 (N_17349,N_16639,N_16823);
xor U17350 (N_17350,N_16498,N_16179);
xor U17351 (N_17351,N_16745,N_16732);
xor U17352 (N_17352,N_16229,N_16964);
xnor U17353 (N_17353,N_16165,N_16167);
and U17354 (N_17354,N_16926,N_16007);
or U17355 (N_17355,N_16516,N_16191);
or U17356 (N_17356,N_16150,N_16471);
xor U17357 (N_17357,N_16479,N_16580);
nor U17358 (N_17358,N_16609,N_16325);
or U17359 (N_17359,N_16721,N_16756);
nand U17360 (N_17360,N_16525,N_16062);
nand U17361 (N_17361,N_16904,N_16186);
xor U17362 (N_17362,N_16873,N_16658);
xnor U17363 (N_17363,N_16559,N_16369);
or U17364 (N_17364,N_16082,N_16060);
or U17365 (N_17365,N_16195,N_16203);
and U17366 (N_17366,N_16813,N_16573);
nor U17367 (N_17367,N_16569,N_16196);
nor U17368 (N_17368,N_16348,N_16870);
and U17369 (N_17369,N_16156,N_16384);
and U17370 (N_17370,N_16868,N_16744);
or U17371 (N_17371,N_16359,N_16491);
and U17372 (N_17372,N_16515,N_16098);
nor U17373 (N_17373,N_16413,N_16533);
xnor U17374 (N_17374,N_16911,N_16059);
or U17375 (N_17375,N_16247,N_16840);
nand U17376 (N_17376,N_16642,N_16863);
nor U17377 (N_17377,N_16770,N_16190);
or U17378 (N_17378,N_16597,N_16494);
and U17379 (N_17379,N_16582,N_16466);
nor U17380 (N_17380,N_16445,N_16759);
xor U17381 (N_17381,N_16218,N_16814);
xnor U17382 (N_17382,N_16427,N_16253);
or U17383 (N_17383,N_16374,N_16044);
xnor U17384 (N_17384,N_16385,N_16268);
xor U17385 (N_17385,N_16842,N_16783);
or U17386 (N_17386,N_16048,N_16214);
nand U17387 (N_17387,N_16117,N_16432);
nor U17388 (N_17388,N_16142,N_16796);
xnor U17389 (N_17389,N_16368,N_16236);
or U17390 (N_17390,N_16492,N_16769);
xnor U17391 (N_17391,N_16834,N_16005);
xor U17392 (N_17392,N_16338,N_16853);
nand U17393 (N_17393,N_16837,N_16509);
and U17394 (N_17394,N_16908,N_16124);
and U17395 (N_17395,N_16760,N_16289);
xnor U17396 (N_17396,N_16476,N_16829);
nand U17397 (N_17397,N_16414,N_16485);
nand U17398 (N_17398,N_16477,N_16528);
and U17399 (N_17399,N_16076,N_16155);
or U17400 (N_17400,N_16545,N_16935);
xor U17401 (N_17401,N_16149,N_16211);
nor U17402 (N_17402,N_16562,N_16644);
or U17403 (N_17403,N_16415,N_16960);
or U17404 (N_17404,N_16629,N_16660);
nand U17405 (N_17405,N_16781,N_16872);
nor U17406 (N_17406,N_16928,N_16024);
or U17407 (N_17407,N_16487,N_16936);
nor U17408 (N_17408,N_16857,N_16793);
nor U17409 (N_17409,N_16401,N_16544);
or U17410 (N_17410,N_16453,N_16623);
and U17411 (N_17411,N_16522,N_16988);
nand U17412 (N_17412,N_16392,N_16577);
nand U17413 (N_17413,N_16058,N_16600);
or U17414 (N_17414,N_16897,N_16711);
nand U17415 (N_17415,N_16959,N_16301);
nor U17416 (N_17416,N_16188,N_16147);
nand U17417 (N_17417,N_16871,N_16265);
or U17418 (N_17418,N_16228,N_16778);
nand U17419 (N_17419,N_16651,N_16365);
nor U17420 (N_17420,N_16751,N_16966);
nor U17421 (N_17421,N_16266,N_16465);
xor U17422 (N_17422,N_16799,N_16323);
and U17423 (N_17423,N_16105,N_16527);
and U17424 (N_17424,N_16807,N_16906);
xor U17425 (N_17425,N_16061,N_16086);
nand U17426 (N_17426,N_16862,N_16364);
nor U17427 (N_17427,N_16537,N_16939);
nor U17428 (N_17428,N_16141,N_16543);
xor U17429 (N_17429,N_16235,N_16638);
nor U17430 (N_17430,N_16715,N_16291);
nor U17431 (N_17431,N_16456,N_16772);
xnor U17432 (N_17432,N_16625,N_16628);
or U17433 (N_17433,N_16530,N_16429);
nand U17434 (N_17434,N_16093,N_16106);
or U17435 (N_17435,N_16567,N_16695);
nor U17436 (N_17436,N_16424,N_16016);
nor U17437 (N_17437,N_16012,N_16683);
nor U17438 (N_17438,N_16313,N_16812);
or U17439 (N_17439,N_16192,N_16343);
nor U17440 (N_17440,N_16563,N_16720);
nand U17441 (N_17441,N_16797,N_16884);
xnor U17442 (N_17442,N_16704,N_16080);
nor U17443 (N_17443,N_16442,N_16020);
xor U17444 (N_17444,N_16045,N_16497);
nand U17445 (N_17445,N_16233,N_16121);
or U17446 (N_17446,N_16269,N_16786);
nand U17447 (N_17447,N_16129,N_16702);
nor U17448 (N_17448,N_16599,N_16841);
nand U17449 (N_17449,N_16689,N_16565);
xor U17450 (N_17450,N_16053,N_16606);
and U17451 (N_17451,N_16717,N_16047);
xor U17452 (N_17452,N_16069,N_16277);
and U17453 (N_17453,N_16090,N_16399);
and U17454 (N_17454,N_16617,N_16423);
nor U17455 (N_17455,N_16321,N_16324);
xor U17456 (N_17456,N_16035,N_16120);
and U17457 (N_17457,N_16815,N_16114);
or U17458 (N_17458,N_16478,N_16713);
nand U17459 (N_17459,N_16349,N_16521);
xnor U17460 (N_17460,N_16282,N_16910);
nand U17461 (N_17461,N_16375,N_16454);
or U17462 (N_17462,N_16583,N_16776);
xor U17463 (N_17463,N_16040,N_16681);
or U17464 (N_17464,N_16968,N_16281);
nor U17465 (N_17465,N_16579,N_16000);
or U17466 (N_17466,N_16674,N_16154);
or U17467 (N_17467,N_16436,N_16470);
nor U17468 (N_17468,N_16898,N_16902);
nor U17469 (N_17469,N_16972,N_16869);
or U17470 (N_17470,N_16534,N_16997);
or U17471 (N_17471,N_16084,N_16802);
or U17472 (N_17472,N_16780,N_16519);
nor U17473 (N_17473,N_16986,N_16063);
xor U17474 (N_17474,N_16275,N_16222);
nand U17475 (N_17475,N_16719,N_16895);
nand U17476 (N_17476,N_16464,N_16822);
xnor U17477 (N_17477,N_16592,N_16686);
nand U17478 (N_17478,N_16256,N_16551);
or U17479 (N_17479,N_16240,N_16925);
or U17480 (N_17480,N_16383,N_16771);
nand U17481 (N_17481,N_16845,N_16723);
xnor U17482 (N_17482,N_16078,N_16795);
xor U17483 (N_17483,N_16334,N_16560);
and U17484 (N_17484,N_16262,N_16404);
nor U17485 (N_17485,N_16096,N_16068);
and U17486 (N_17486,N_16274,N_16867);
nor U17487 (N_17487,N_16087,N_16116);
nor U17488 (N_17488,N_16437,N_16306);
nor U17489 (N_17489,N_16354,N_16693);
nand U17490 (N_17490,N_16112,N_16234);
and U17491 (N_17491,N_16784,N_16633);
xnor U17492 (N_17492,N_16435,N_16019);
nor U17493 (N_17493,N_16346,N_16373);
or U17494 (N_17494,N_16722,N_16750);
xor U17495 (N_17495,N_16916,N_16286);
xnor U17496 (N_17496,N_16692,N_16694);
or U17497 (N_17497,N_16370,N_16875);
nor U17498 (N_17498,N_16312,N_16450);
and U17499 (N_17499,N_16170,N_16971);
nand U17500 (N_17500,N_16440,N_16458);
and U17501 (N_17501,N_16830,N_16631);
nor U17502 (N_17502,N_16311,N_16731);
nor U17503 (N_17503,N_16142,N_16892);
or U17504 (N_17504,N_16400,N_16254);
nor U17505 (N_17505,N_16968,N_16762);
nand U17506 (N_17506,N_16667,N_16534);
xor U17507 (N_17507,N_16137,N_16808);
and U17508 (N_17508,N_16116,N_16540);
nor U17509 (N_17509,N_16870,N_16411);
xor U17510 (N_17510,N_16802,N_16628);
or U17511 (N_17511,N_16700,N_16259);
and U17512 (N_17512,N_16852,N_16552);
or U17513 (N_17513,N_16294,N_16574);
nor U17514 (N_17514,N_16894,N_16441);
or U17515 (N_17515,N_16104,N_16033);
nor U17516 (N_17516,N_16502,N_16311);
xnor U17517 (N_17517,N_16975,N_16471);
nor U17518 (N_17518,N_16517,N_16395);
and U17519 (N_17519,N_16125,N_16422);
xor U17520 (N_17520,N_16522,N_16277);
or U17521 (N_17521,N_16816,N_16020);
or U17522 (N_17522,N_16844,N_16693);
and U17523 (N_17523,N_16770,N_16029);
nand U17524 (N_17524,N_16382,N_16454);
or U17525 (N_17525,N_16375,N_16982);
nand U17526 (N_17526,N_16191,N_16047);
and U17527 (N_17527,N_16951,N_16740);
xnor U17528 (N_17528,N_16750,N_16595);
xor U17529 (N_17529,N_16502,N_16069);
nand U17530 (N_17530,N_16147,N_16780);
and U17531 (N_17531,N_16831,N_16459);
and U17532 (N_17532,N_16301,N_16066);
nor U17533 (N_17533,N_16637,N_16926);
xor U17534 (N_17534,N_16382,N_16293);
nor U17535 (N_17535,N_16006,N_16560);
or U17536 (N_17536,N_16507,N_16205);
xnor U17537 (N_17537,N_16856,N_16723);
xnor U17538 (N_17538,N_16522,N_16567);
nor U17539 (N_17539,N_16896,N_16618);
nand U17540 (N_17540,N_16027,N_16758);
nand U17541 (N_17541,N_16271,N_16432);
xor U17542 (N_17542,N_16579,N_16154);
xnor U17543 (N_17543,N_16050,N_16667);
nand U17544 (N_17544,N_16045,N_16319);
nor U17545 (N_17545,N_16556,N_16621);
nor U17546 (N_17546,N_16554,N_16695);
nand U17547 (N_17547,N_16231,N_16899);
nand U17548 (N_17548,N_16445,N_16468);
or U17549 (N_17549,N_16335,N_16924);
or U17550 (N_17550,N_16438,N_16005);
and U17551 (N_17551,N_16250,N_16681);
or U17552 (N_17552,N_16789,N_16979);
nand U17553 (N_17553,N_16844,N_16079);
or U17554 (N_17554,N_16081,N_16085);
or U17555 (N_17555,N_16707,N_16192);
and U17556 (N_17556,N_16070,N_16058);
and U17557 (N_17557,N_16681,N_16651);
nor U17558 (N_17558,N_16938,N_16527);
or U17559 (N_17559,N_16721,N_16978);
xor U17560 (N_17560,N_16211,N_16204);
xor U17561 (N_17561,N_16578,N_16337);
nand U17562 (N_17562,N_16117,N_16743);
xnor U17563 (N_17563,N_16472,N_16251);
and U17564 (N_17564,N_16168,N_16203);
xor U17565 (N_17565,N_16383,N_16960);
nand U17566 (N_17566,N_16932,N_16297);
nor U17567 (N_17567,N_16219,N_16214);
nand U17568 (N_17568,N_16750,N_16768);
or U17569 (N_17569,N_16666,N_16648);
xor U17570 (N_17570,N_16439,N_16226);
or U17571 (N_17571,N_16981,N_16566);
nand U17572 (N_17572,N_16817,N_16703);
nand U17573 (N_17573,N_16356,N_16936);
xnor U17574 (N_17574,N_16877,N_16895);
nor U17575 (N_17575,N_16423,N_16044);
nor U17576 (N_17576,N_16925,N_16355);
nor U17577 (N_17577,N_16495,N_16999);
nand U17578 (N_17578,N_16204,N_16849);
or U17579 (N_17579,N_16176,N_16380);
and U17580 (N_17580,N_16430,N_16632);
nand U17581 (N_17581,N_16362,N_16698);
xor U17582 (N_17582,N_16191,N_16445);
nor U17583 (N_17583,N_16046,N_16146);
or U17584 (N_17584,N_16944,N_16494);
nand U17585 (N_17585,N_16155,N_16678);
and U17586 (N_17586,N_16452,N_16426);
nand U17587 (N_17587,N_16988,N_16218);
and U17588 (N_17588,N_16267,N_16782);
xor U17589 (N_17589,N_16542,N_16299);
nor U17590 (N_17590,N_16685,N_16268);
xor U17591 (N_17591,N_16333,N_16118);
nand U17592 (N_17592,N_16913,N_16378);
and U17593 (N_17593,N_16137,N_16985);
or U17594 (N_17594,N_16074,N_16429);
and U17595 (N_17595,N_16178,N_16864);
nand U17596 (N_17596,N_16834,N_16953);
nor U17597 (N_17597,N_16054,N_16502);
nand U17598 (N_17598,N_16982,N_16771);
nand U17599 (N_17599,N_16715,N_16609);
or U17600 (N_17600,N_16258,N_16781);
or U17601 (N_17601,N_16721,N_16119);
and U17602 (N_17602,N_16250,N_16816);
and U17603 (N_17603,N_16179,N_16051);
nor U17604 (N_17604,N_16480,N_16947);
and U17605 (N_17605,N_16411,N_16533);
or U17606 (N_17606,N_16319,N_16387);
xnor U17607 (N_17607,N_16815,N_16197);
and U17608 (N_17608,N_16686,N_16742);
nor U17609 (N_17609,N_16755,N_16362);
nand U17610 (N_17610,N_16376,N_16250);
and U17611 (N_17611,N_16054,N_16835);
xor U17612 (N_17612,N_16413,N_16848);
or U17613 (N_17613,N_16229,N_16727);
and U17614 (N_17614,N_16741,N_16506);
nand U17615 (N_17615,N_16115,N_16971);
nand U17616 (N_17616,N_16219,N_16802);
xor U17617 (N_17617,N_16181,N_16379);
nor U17618 (N_17618,N_16209,N_16511);
and U17619 (N_17619,N_16478,N_16184);
and U17620 (N_17620,N_16684,N_16232);
xor U17621 (N_17621,N_16241,N_16993);
nand U17622 (N_17622,N_16477,N_16330);
xor U17623 (N_17623,N_16697,N_16502);
and U17624 (N_17624,N_16347,N_16153);
or U17625 (N_17625,N_16799,N_16433);
xnor U17626 (N_17626,N_16873,N_16931);
xnor U17627 (N_17627,N_16795,N_16091);
nand U17628 (N_17628,N_16780,N_16551);
xnor U17629 (N_17629,N_16143,N_16024);
xor U17630 (N_17630,N_16825,N_16031);
nand U17631 (N_17631,N_16719,N_16247);
xor U17632 (N_17632,N_16746,N_16706);
or U17633 (N_17633,N_16492,N_16315);
or U17634 (N_17634,N_16546,N_16888);
and U17635 (N_17635,N_16473,N_16701);
and U17636 (N_17636,N_16452,N_16170);
xnor U17637 (N_17637,N_16393,N_16594);
nor U17638 (N_17638,N_16663,N_16489);
nor U17639 (N_17639,N_16672,N_16595);
and U17640 (N_17640,N_16138,N_16289);
nor U17641 (N_17641,N_16568,N_16853);
and U17642 (N_17642,N_16979,N_16202);
nand U17643 (N_17643,N_16429,N_16670);
xor U17644 (N_17644,N_16901,N_16132);
nor U17645 (N_17645,N_16228,N_16200);
xor U17646 (N_17646,N_16614,N_16334);
nand U17647 (N_17647,N_16332,N_16077);
and U17648 (N_17648,N_16404,N_16899);
nor U17649 (N_17649,N_16554,N_16615);
xnor U17650 (N_17650,N_16048,N_16343);
nor U17651 (N_17651,N_16626,N_16243);
nor U17652 (N_17652,N_16493,N_16045);
xor U17653 (N_17653,N_16498,N_16348);
or U17654 (N_17654,N_16285,N_16393);
and U17655 (N_17655,N_16288,N_16807);
xnor U17656 (N_17656,N_16302,N_16744);
or U17657 (N_17657,N_16210,N_16023);
nand U17658 (N_17658,N_16655,N_16510);
or U17659 (N_17659,N_16807,N_16155);
and U17660 (N_17660,N_16507,N_16246);
nand U17661 (N_17661,N_16193,N_16776);
or U17662 (N_17662,N_16827,N_16931);
nand U17663 (N_17663,N_16340,N_16194);
nor U17664 (N_17664,N_16298,N_16226);
or U17665 (N_17665,N_16596,N_16141);
or U17666 (N_17666,N_16271,N_16850);
and U17667 (N_17667,N_16145,N_16170);
and U17668 (N_17668,N_16551,N_16868);
nor U17669 (N_17669,N_16401,N_16804);
and U17670 (N_17670,N_16750,N_16935);
and U17671 (N_17671,N_16102,N_16253);
xor U17672 (N_17672,N_16755,N_16441);
or U17673 (N_17673,N_16066,N_16810);
and U17674 (N_17674,N_16534,N_16376);
and U17675 (N_17675,N_16025,N_16185);
nand U17676 (N_17676,N_16813,N_16177);
nor U17677 (N_17677,N_16062,N_16854);
nand U17678 (N_17678,N_16166,N_16956);
nand U17679 (N_17679,N_16491,N_16140);
nand U17680 (N_17680,N_16030,N_16308);
nand U17681 (N_17681,N_16704,N_16334);
or U17682 (N_17682,N_16362,N_16138);
nor U17683 (N_17683,N_16114,N_16675);
or U17684 (N_17684,N_16633,N_16070);
nor U17685 (N_17685,N_16350,N_16664);
nand U17686 (N_17686,N_16339,N_16533);
nand U17687 (N_17687,N_16863,N_16829);
and U17688 (N_17688,N_16585,N_16121);
nand U17689 (N_17689,N_16251,N_16360);
nor U17690 (N_17690,N_16422,N_16134);
and U17691 (N_17691,N_16012,N_16718);
or U17692 (N_17692,N_16272,N_16323);
xnor U17693 (N_17693,N_16735,N_16671);
nor U17694 (N_17694,N_16099,N_16722);
xnor U17695 (N_17695,N_16348,N_16596);
nand U17696 (N_17696,N_16975,N_16413);
nand U17697 (N_17697,N_16802,N_16978);
and U17698 (N_17698,N_16355,N_16048);
nor U17699 (N_17699,N_16233,N_16031);
nand U17700 (N_17700,N_16474,N_16124);
nor U17701 (N_17701,N_16976,N_16726);
or U17702 (N_17702,N_16883,N_16479);
nand U17703 (N_17703,N_16567,N_16369);
xor U17704 (N_17704,N_16323,N_16028);
nor U17705 (N_17705,N_16749,N_16332);
nor U17706 (N_17706,N_16655,N_16884);
nor U17707 (N_17707,N_16426,N_16394);
and U17708 (N_17708,N_16937,N_16496);
and U17709 (N_17709,N_16342,N_16038);
and U17710 (N_17710,N_16602,N_16756);
nor U17711 (N_17711,N_16997,N_16728);
nand U17712 (N_17712,N_16930,N_16087);
nor U17713 (N_17713,N_16998,N_16326);
nand U17714 (N_17714,N_16923,N_16576);
or U17715 (N_17715,N_16818,N_16718);
nor U17716 (N_17716,N_16664,N_16288);
xnor U17717 (N_17717,N_16534,N_16021);
nand U17718 (N_17718,N_16106,N_16863);
or U17719 (N_17719,N_16773,N_16870);
and U17720 (N_17720,N_16519,N_16229);
or U17721 (N_17721,N_16133,N_16029);
and U17722 (N_17722,N_16349,N_16043);
or U17723 (N_17723,N_16143,N_16116);
nand U17724 (N_17724,N_16369,N_16876);
nor U17725 (N_17725,N_16751,N_16697);
and U17726 (N_17726,N_16615,N_16318);
nor U17727 (N_17727,N_16975,N_16171);
nand U17728 (N_17728,N_16491,N_16610);
or U17729 (N_17729,N_16516,N_16584);
or U17730 (N_17730,N_16525,N_16173);
or U17731 (N_17731,N_16966,N_16489);
or U17732 (N_17732,N_16922,N_16853);
xnor U17733 (N_17733,N_16420,N_16787);
or U17734 (N_17734,N_16905,N_16997);
xor U17735 (N_17735,N_16770,N_16890);
xnor U17736 (N_17736,N_16160,N_16242);
nand U17737 (N_17737,N_16185,N_16677);
or U17738 (N_17738,N_16692,N_16345);
nor U17739 (N_17739,N_16170,N_16249);
and U17740 (N_17740,N_16795,N_16011);
or U17741 (N_17741,N_16169,N_16496);
and U17742 (N_17742,N_16112,N_16640);
nor U17743 (N_17743,N_16853,N_16821);
or U17744 (N_17744,N_16710,N_16804);
nand U17745 (N_17745,N_16561,N_16817);
and U17746 (N_17746,N_16918,N_16724);
or U17747 (N_17747,N_16966,N_16949);
or U17748 (N_17748,N_16213,N_16144);
xor U17749 (N_17749,N_16790,N_16216);
nand U17750 (N_17750,N_16058,N_16473);
or U17751 (N_17751,N_16224,N_16752);
or U17752 (N_17752,N_16379,N_16675);
nand U17753 (N_17753,N_16563,N_16528);
and U17754 (N_17754,N_16000,N_16342);
or U17755 (N_17755,N_16501,N_16301);
nor U17756 (N_17756,N_16948,N_16009);
and U17757 (N_17757,N_16502,N_16426);
and U17758 (N_17758,N_16297,N_16559);
nand U17759 (N_17759,N_16622,N_16316);
or U17760 (N_17760,N_16900,N_16621);
xor U17761 (N_17761,N_16530,N_16414);
nand U17762 (N_17762,N_16364,N_16637);
nand U17763 (N_17763,N_16390,N_16130);
and U17764 (N_17764,N_16430,N_16368);
xnor U17765 (N_17765,N_16169,N_16827);
nor U17766 (N_17766,N_16991,N_16431);
nand U17767 (N_17767,N_16739,N_16104);
and U17768 (N_17768,N_16659,N_16842);
and U17769 (N_17769,N_16486,N_16668);
nor U17770 (N_17770,N_16234,N_16568);
xor U17771 (N_17771,N_16865,N_16360);
and U17772 (N_17772,N_16350,N_16514);
and U17773 (N_17773,N_16710,N_16775);
nand U17774 (N_17774,N_16954,N_16231);
or U17775 (N_17775,N_16542,N_16987);
nand U17776 (N_17776,N_16629,N_16417);
xnor U17777 (N_17777,N_16503,N_16965);
nor U17778 (N_17778,N_16264,N_16706);
nor U17779 (N_17779,N_16429,N_16319);
or U17780 (N_17780,N_16136,N_16123);
xor U17781 (N_17781,N_16574,N_16936);
xnor U17782 (N_17782,N_16669,N_16817);
or U17783 (N_17783,N_16421,N_16675);
nand U17784 (N_17784,N_16340,N_16842);
nor U17785 (N_17785,N_16318,N_16235);
nor U17786 (N_17786,N_16292,N_16324);
nand U17787 (N_17787,N_16332,N_16775);
nor U17788 (N_17788,N_16833,N_16363);
xnor U17789 (N_17789,N_16218,N_16819);
nand U17790 (N_17790,N_16739,N_16553);
xor U17791 (N_17791,N_16484,N_16181);
nand U17792 (N_17792,N_16455,N_16467);
xor U17793 (N_17793,N_16239,N_16723);
nand U17794 (N_17794,N_16611,N_16654);
nor U17795 (N_17795,N_16068,N_16675);
or U17796 (N_17796,N_16715,N_16209);
nor U17797 (N_17797,N_16130,N_16192);
nand U17798 (N_17798,N_16206,N_16375);
or U17799 (N_17799,N_16925,N_16286);
and U17800 (N_17800,N_16078,N_16459);
xnor U17801 (N_17801,N_16920,N_16691);
nand U17802 (N_17802,N_16434,N_16433);
or U17803 (N_17803,N_16265,N_16650);
nand U17804 (N_17804,N_16508,N_16301);
or U17805 (N_17805,N_16362,N_16704);
nand U17806 (N_17806,N_16683,N_16974);
nand U17807 (N_17807,N_16574,N_16137);
and U17808 (N_17808,N_16355,N_16639);
xnor U17809 (N_17809,N_16926,N_16323);
xnor U17810 (N_17810,N_16741,N_16375);
nor U17811 (N_17811,N_16066,N_16234);
or U17812 (N_17812,N_16403,N_16027);
xnor U17813 (N_17813,N_16692,N_16895);
or U17814 (N_17814,N_16404,N_16747);
xor U17815 (N_17815,N_16953,N_16655);
nand U17816 (N_17816,N_16977,N_16493);
or U17817 (N_17817,N_16583,N_16526);
xor U17818 (N_17818,N_16110,N_16311);
or U17819 (N_17819,N_16729,N_16276);
nor U17820 (N_17820,N_16036,N_16102);
xor U17821 (N_17821,N_16384,N_16194);
nand U17822 (N_17822,N_16409,N_16025);
and U17823 (N_17823,N_16882,N_16964);
or U17824 (N_17824,N_16162,N_16288);
nor U17825 (N_17825,N_16563,N_16087);
or U17826 (N_17826,N_16344,N_16928);
nor U17827 (N_17827,N_16717,N_16943);
xor U17828 (N_17828,N_16153,N_16690);
or U17829 (N_17829,N_16189,N_16663);
and U17830 (N_17830,N_16205,N_16193);
or U17831 (N_17831,N_16395,N_16056);
and U17832 (N_17832,N_16881,N_16470);
nor U17833 (N_17833,N_16313,N_16485);
nor U17834 (N_17834,N_16874,N_16595);
and U17835 (N_17835,N_16739,N_16577);
nor U17836 (N_17836,N_16728,N_16182);
or U17837 (N_17837,N_16027,N_16040);
and U17838 (N_17838,N_16590,N_16581);
xnor U17839 (N_17839,N_16829,N_16713);
or U17840 (N_17840,N_16009,N_16990);
or U17841 (N_17841,N_16843,N_16323);
and U17842 (N_17842,N_16117,N_16019);
or U17843 (N_17843,N_16675,N_16799);
xor U17844 (N_17844,N_16989,N_16275);
or U17845 (N_17845,N_16870,N_16165);
and U17846 (N_17846,N_16874,N_16337);
nand U17847 (N_17847,N_16297,N_16119);
nand U17848 (N_17848,N_16715,N_16915);
nand U17849 (N_17849,N_16269,N_16384);
nor U17850 (N_17850,N_16520,N_16323);
nand U17851 (N_17851,N_16837,N_16976);
xor U17852 (N_17852,N_16772,N_16481);
nor U17853 (N_17853,N_16450,N_16203);
or U17854 (N_17854,N_16471,N_16957);
nor U17855 (N_17855,N_16538,N_16886);
or U17856 (N_17856,N_16740,N_16422);
xnor U17857 (N_17857,N_16917,N_16061);
nand U17858 (N_17858,N_16350,N_16219);
nand U17859 (N_17859,N_16135,N_16172);
or U17860 (N_17860,N_16560,N_16116);
and U17861 (N_17861,N_16466,N_16957);
nand U17862 (N_17862,N_16963,N_16257);
and U17863 (N_17863,N_16214,N_16770);
and U17864 (N_17864,N_16076,N_16135);
and U17865 (N_17865,N_16584,N_16088);
and U17866 (N_17866,N_16947,N_16614);
nor U17867 (N_17867,N_16066,N_16705);
nor U17868 (N_17868,N_16571,N_16392);
xor U17869 (N_17869,N_16818,N_16925);
nor U17870 (N_17870,N_16481,N_16291);
nand U17871 (N_17871,N_16850,N_16106);
nor U17872 (N_17872,N_16633,N_16922);
and U17873 (N_17873,N_16592,N_16982);
xnor U17874 (N_17874,N_16570,N_16806);
nor U17875 (N_17875,N_16843,N_16398);
nand U17876 (N_17876,N_16832,N_16983);
nor U17877 (N_17877,N_16416,N_16571);
and U17878 (N_17878,N_16021,N_16002);
nand U17879 (N_17879,N_16322,N_16144);
xor U17880 (N_17880,N_16964,N_16022);
nor U17881 (N_17881,N_16831,N_16248);
nand U17882 (N_17882,N_16165,N_16881);
and U17883 (N_17883,N_16399,N_16229);
or U17884 (N_17884,N_16774,N_16967);
nor U17885 (N_17885,N_16584,N_16057);
and U17886 (N_17886,N_16644,N_16655);
nand U17887 (N_17887,N_16695,N_16315);
and U17888 (N_17888,N_16523,N_16192);
nand U17889 (N_17889,N_16916,N_16595);
nor U17890 (N_17890,N_16668,N_16559);
or U17891 (N_17891,N_16031,N_16930);
xor U17892 (N_17892,N_16653,N_16821);
xor U17893 (N_17893,N_16990,N_16072);
nor U17894 (N_17894,N_16138,N_16497);
xor U17895 (N_17895,N_16640,N_16750);
xnor U17896 (N_17896,N_16367,N_16317);
nand U17897 (N_17897,N_16474,N_16111);
nand U17898 (N_17898,N_16895,N_16701);
or U17899 (N_17899,N_16946,N_16134);
nor U17900 (N_17900,N_16916,N_16002);
nor U17901 (N_17901,N_16977,N_16555);
xnor U17902 (N_17902,N_16556,N_16040);
xnor U17903 (N_17903,N_16216,N_16301);
xnor U17904 (N_17904,N_16829,N_16983);
or U17905 (N_17905,N_16960,N_16888);
or U17906 (N_17906,N_16516,N_16966);
nor U17907 (N_17907,N_16327,N_16026);
nand U17908 (N_17908,N_16872,N_16476);
xor U17909 (N_17909,N_16388,N_16782);
or U17910 (N_17910,N_16241,N_16420);
nand U17911 (N_17911,N_16266,N_16261);
and U17912 (N_17912,N_16237,N_16449);
nor U17913 (N_17913,N_16027,N_16783);
or U17914 (N_17914,N_16550,N_16736);
nor U17915 (N_17915,N_16318,N_16662);
xnor U17916 (N_17916,N_16762,N_16333);
xor U17917 (N_17917,N_16546,N_16438);
nor U17918 (N_17918,N_16718,N_16908);
or U17919 (N_17919,N_16213,N_16151);
nand U17920 (N_17920,N_16633,N_16051);
nor U17921 (N_17921,N_16266,N_16003);
xor U17922 (N_17922,N_16652,N_16576);
nand U17923 (N_17923,N_16293,N_16110);
nor U17924 (N_17924,N_16230,N_16314);
nand U17925 (N_17925,N_16174,N_16953);
xnor U17926 (N_17926,N_16363,N_16214);
and U17927 (N_17927,N_16644,N_16892);
xnor U17928 (N_17928,N_16905,N_16364);
and U17929 (N_17929,N_16369,N_16518);
nand U17930 (N_17930,N_16823,N_16069);
or U17931 (N_17931,N_16009,N_16971);
nor U17932 (N_17932,N_16142,N_16917);
nand U17933 (N_17933,N_16249,N_16896);
xor U17934 (N_17934,N_16067,N_16759);
or U17935 (N_17935,N_16337,N_16254);
nor U17936 (N_17936,N_16839,N_16638);
xor U17937 (N_17937,N_16224,N_16255);
or U17938 (N_17938,N_16702,N_16612);
and U17939 (N_17939,N_16043,N_16402);
xnor U17940 (N_17940,N_16221,N_16344);
and U17941 (N_17941,N_16899,N_16376);
xor U17942 (N_17942,N_16362,N_16614);
nor U17943 (N_17943,N_16244,N_16853);
nor U17944 (N_17944,N_16815,N_16257);
or U17945 (N_17945,N_16431,N_16593);
xor U17946 (N_17946,N_16750,N_16048);
and U17947 (N_17947,N_16621,N_16600);
nand U17948 (N_17948,N_16493,N_16089);
or U17949 (N_17949,N_16160,N_16288);
nor U17950 (N_17950,N_16180,N_16394);
and U17951 (N_17951,N_16992,N_16552);
and U17952 (N_17952,N_16716,N_16047);
nand U17953 (N_17953,N_16713,N_16323);
and U17954 (N_17954,N_16535,N_16123);
xor U17955 (N_17955,N_16857,N_16851);
xor U17956 (N_17956,N_16280,N_16642);
xnor U17957 (N_17957,N_16489,N_16364);
xnor U17958 (N_17958,N_16004,N_16010);
xnor U17959 (N_17959,N_16774,N_16358);
nor U17960 (N_17960,N_16501,N_16035);
nor U17961 (N_17961,N_16650,N_16179);
xnor U17962 (N_17962,N_16276,N_16091);
or U17963 (N_17963,N_16152,N_16166);
and U17964 (N_17964,N_16814,N_16427);
xnor U17965 (N_17965,N_16246,N_16135);
or U17966 (N_17966,N_16385,N_16187);
and U17967 (N_17967,N_16485,N_16713);
xnor U17968 (N_17968,N_16494,N_16650);
xor U17969 (N_17969,N_16540,N_16181);
xnor U17970 (N_17970,N_16808,N_16835);
xnor U17971 (N_17971,N_16951,N_16074);
and U17972 (N_17972,N_16382,N_16651);
nand U17973 (N_17973,N_16847,N_16766);
and U17974 (N_17974,N_16746,N_16235);
nor U17975 (N_17975,N_16693,N_16516);
nor U17976 (N_17976,N_16847,N_16898);
nand U17977 (N_17977,N_16557,N_16959);
nor U17978 (N_17978,N_16460,N_16826);
nand U17979 (N_17979,N_16663,N_16713);
and U17980 (N_17980,N_16340,N_16502);
or U17981 (N_17981,N_16100,N_16944);
xor U17982 (N_17982,N_16977,N_16723);
and U17983 (N_17983,N_16266,N_16921);
xnor U17984 (N_17984,N_16463,N_16202);
and U17985 (N_17985,N_16259,N_16879);
nand U17986 (N_17986,N_16166,N_16225);
and U17987 (N_17987,N_16782,N_16325);
or U17988 (N_17988,N_16402,N_16528);
nand U17989 (N_17989,N_16653,N_16332);
nor U17990 (N_17990,N_16510,N_16501);
and U17991 (N_17991,N_16998,N_16367);
xor U17992 (N_17992,N_16640,N_16848);
nand U17993 (N_17993,N_16872,N_16909);
nor U17994 (N_17994,N_16341,N_16460);
nand U17995 (N_17995,N_16710,N_16554);
nand U17996 (N_17996,N_16819,N_16279);
xnor U17997 (N_17997,N_16862,N_16358);
nand U17998 (N_17998,N_16770,N_16491);
xnor U17999 (N_17999,N_16784,N_16278);
nand U18000 (N_18000,N_17455,N_17287);
nand U18001 (N_18001,N_17331,N_17135);
xnor U18002 (N_18002,N_17677,N_17885);
xor U18003 (N_18003,N_17465,N_17581);
and U18004 (N_18004,N_17440,N_17250);
nand U18005 (N_18005,N_17973,N_17311);
and U18006 (N_18006,N_17411,N_17899);
and U18007 (N_18007,N_17922,N_17728);
nor U18008 (N_18008,N_17467,N_17236);
and U18009 (N_18009,N_17063,N_17735);
xor U18010 (N_18010,N_17818,N_17383);
or U18011 (N_18011,N_17351,N_17950);
or U18012 (N_18012,N_17346,N_17057);
nor U18013 (N_18013,N_17322,N_17141);
and U18014 (N_18014,N_17801,N_17679);
or U18015 (N_18015,N_17255,N_17772);
nor U18016 (N_18016,N_17364,N_17382);
xor U18017 (N_18017,N_17684,N_17290);
nor U18018 (N_18018,N_17976,N_17514);
or U18019 (N_18019,N_17261,N_17209);
nor U18020 (N_18020,N_17779,N_17075);
or U18021 (N_18021,N_17282,N_17632);
and U18022 (N_18022,N_17994,N_17725);
and U18023 (N_18023,N_17821,N_17252);
nand U18024 (N_18024,N_17017,N_17225);
and U18025 (N_18025,N_17855,N_17452);
or U18026 (N_18026,N_17985,N_17007);
nor U18027 (N_18027,N_17197,N_17582);
or U18028 (N_18028,N_17620,N_17592);
or U18029 (N_18029,N_17004,N_17165);
and U18030 (N_18030,N_17021,N_17228);
and U18031 (N_18031,N_17430,N_17029);
and U18032 (N_18032,N_17334,N_17519);
nor U18033 (N_18033,N_17489,N_17326);
nor U18034 (N_18034,N_17659,N_17476);
xor U18035 (N_18035,N_17655,N_17160);
and U18036 (N_18036,N_17940,N_17791);
and U18037 (N_18037,N_17518,N_17061);
nand U18038 (N_18038,N_17494,N_17926);
xnor U18039 (N_18039,N_17961,N_17258);
nand U18040 (N_18040,N_17148,N_17304);
xnor U18041 (N_18041,N_17826,N_17571);
xnor U18042 (N_18042,N_17115,N_17338);
nand U18043 (N_18043,N_17578,N_17937);
or U18044 (N_18044,N_17883,N_17403);
xnor U18045 (N_18045,N_17471,N_17915);
and U18046 (N_18046,N_17069,N_17595);
xnor U18047 (N_18047,N_17213,N_17834);
and U18048 (N_18048,N_17720,N_17907);
or U18049 (N_18049,N_17525,N_17897);
nand U18050 (N_18050,N_17757,N_17830);
nand U18051 (N_18051,N_17627,N_17876);
nand U18052 (N_18052,N_17675,N_17413);
xor U18053 (N_18053,N_17898,N_17929);
or U18054 (N_18054,N_17152,N_17234);
nor U18055 (N_18055,N_17888,N_17729);
nor U18056 (N_18056,N_17128,N_17805);
or U18057 (N_18057,N_17210,N_17773);
xor U18058 (N_18058,N_17886,N_17113);
xnor U18059 (N_18059,N_17536,N_17295);
or U18060 (N_18060,N_17217,N_17241);
and U18061 (N_18061,N_17512,N_17248);
and U18062 (N_18062,N_17739,N_17761);
nor U18063 (N_18063,N_17874,N_17185);
nor U18064 (N_18064,N_17917,N_17428);
or U18065 (N_18065,N_17035,N_17280);
nor U18066 (N_18066,N_17871,N_17590);
nand U18067 (N_18067,N_17373,N_17804);
nor U18068 (N_18068,N_17616,N_17624);
or U18069 (N_18069,N_17125,N_17506);
nor U18070 (N_18070,N_17169,N_17386);
and U18071 (N_18071,N_17817,N_17074);
nand U18072 (N_18072,N_17175,N_17780);
nor U18073 (N_18073,N_17755,N_17199);
nand U18074 (N_18074,N_17468,N_17363);
or U18075 (N_18075,N_17177,N_17221);
and U18076 (N_18076,N_17538,N_17544);
nor U18077 (N_18077,N_17835,N_17588);
nand U18078 (N_18078,N_17481,N_17243);
and U18079 (N_18079,N_17972,N_17150);
and U18080 (N_18080,N_17923,N_17060);
nand U18081 (N_18081,N_17587,N_17142);
and U18082 (N_18082,N_17919,N_17783);
xnor U18083 (N_18083,N_17018,N_17662);
nand U18084 (N_18084,N_17895,N_17957);
or U18085 (N_18085,N_17227,N_17577);
xor U18086 (N_18086,N_17505,N_17763);
and U18087 (N_18087,N_17466,N_17615);
xnor U18088 (N_18088,N_17104,N_17734);
nor U18089 (N_18089,N_17661,N_17054);
nand U18090 (N_18090,N_17349,N_17813);
xor U18091 (N_18091,N_17884,N_17245);
and U18092 (N_18092,N_17056,N_17597);
and U18093 (N_18093,N_17718,N_17703);
and U18094 (N_18094,N_17307,N_17510);
nand U18095 (N_18095,N_17106,N_17573);
nand U18096 (N_18096,N_17353,N_17443);
xnor U18097 (N_18097,N_17784,N_17977);
or U18098 (N_18098,N_17132,N_17006);
xor U18099 (N_18099,N_17020,N_17191);
and U18100 (N_18100,N_17508,N_17078);
nor U18101 (N_18101,N_17313,N_17031);
nand U18102 (N_18102,N_17497,N_17374);
nand U18103 (N_18103,N_17491,N_17921);
xor U18104 (N_18104,N_17194,N_17012);
or U18105 (N_18105,N_17291,N_17449);
xnor U18106 (N_18106,N_17186,N_17741);
xor U18107 (N_18107,N_17831,N_17118);
or U18108 (N_18108,N_17939,N_17523);
nand U18109 (N_18109,N_17712,N_17111);
xnor U18110 (N_18110,N_17669,N_17952);
xor U18111 (N_18111,N_17633,N_17664);
and U18112 (N_18112,N_17790,N_17266);
or U18113 (N_18113,N_17803,N_17429);
nand U18114 (N_18114,N_17814,N_17045);
nor U18115 (N_18115,N_17911,N_17833);
or U18116 (N_18116,N_17176,N_17325);
or U18117 (N_18117,N_17259,N_17656);
and U18118 (N_18118,N_17405,N_17279);
or U18119 (N_18119,N_17629,N_17609);
nand U18120 (N_18120,N_17232,N_17686);
nor U18121 (N_18121,N_17201,N_17963);
xor U18122 (N_18122,N_17960,N_17119);
or U18123 (N_18123,N_17242,N_17585);
xor U18124 (N_18124,N_17216,N_17460);
or U18125 (N_18125,N_17193,N_17740);
and U18126 (N_18126,N_17708,N_17516);
or U18127 (N_18127,N_17402,N_17726);
nand U18128 (N_18128,N_17869,N_17848);
xnor U18129 (N_18129,N_17947,N_17164);
nand U18130 (N_18130,N_17231,N_17626);
nand U18131 (N_18131,N_17161,N_17230);
and U18132 (N_18132,N_17011,N_17882);
or U18133 (N_18133,N_17001,N_17996);
or U18134 (N_18134,N_17704,N_17643);
xor U18135 (N_18135,N_17085,N_17859);
xor U18136 (N_18136,N_17215,N_17737);
or U18137 (N_18137,N_17842,N_17828);
xnor U18138 (N_18138,N_17219,N_17392);
nand U18139 (N_18139,N_17042,N_17114);
or U18140 (N_18140,N_17362,N_17569);
nand U18141 (N_18141,N_17076,N_17984);
nor U18142 (N_18142,N_17837,N_17660);
nor U18143 (N_18143,N_17877,N_17134);
nand U18144 (N_18144,N_17109,N_17495);
or U18145 (N_18145,N_17249,N_17576);
or U18146 (N_18146,N_17314,N_17167);
or U18147 (N_18147,N_17532,N_17556);
xor U18148 (N_18148,N_17274,N_17610);
or U18149 (N_18149,N_17044,N_17694);
nor U18150 (N_18150,N_17680,N_17158);
nor U18151 (N_18151,N_17438,N_17603);
xnor U18152 (N_18152,N_17381,N_17500);
or U18153 (N_18153,N_17435,N_17064);
and U18154 (N_18154,N_17327,N_17036);
nand U18155 (N_18155,N_17930,N_17000);
or U18156 (N_18156,N_17016,N_17564);
xnor U18157 (N_18157,N_17574,N_17296);
nor U18158 (N_18158,N_17579,N_17671);
nor U18159 (N_18159,N_17553,N_17836);
nand U18160 (N_18160,N_17529,N_17102);
nor U18161 (N_18161,N_17025,N_17964);
nor U18162 (N_18162,N_17336,N_17802);
xnor U18163 (N_18163,N_17567,N_17372);
or U18164 (N_18164,N_17945,N_17824);
nand U18165 (N_18165,N_17808,N_17370);
or U18166 (N_18166,N_17071,N_17395);
and U18167 (N_18167,N_17748,N_17070);
nand U18168 (N_18168,N_17584,N_17224);
nor U18169 (N_18169,N_17618,N_17909);
and U18170 (N_18170,N_17407,N_17146);
nand U18171 (N_18171,N_17463,N_17707);
or U18172 (N_18172,N_17752,N_17565);
xnor U18173 (N_18173,N_17867,N_17657);
xor U18174 (N_18174,N_17543,N_17724);
xor U18175 (N_18175,N_17744,N_17286);
nand U18176 (N_18176,N_17920,N_17200);
and U18177 (N_18177,N_17670,N_17348);
nor U18178 (N_18178,N_17124,N_17275);
or U18179 (N_18179,N_17753,N_17003);
nor U18180 (N_18180,N_17858,N_17086);
xor U18181 (N_18181,N_17781,N_17665);
nor U18182 (N_18182,N_17637,N_17103);
or U18183 (N_18183,N_17902,N_17663);
nand U18184 (N_18184,N_17490,N_17163);
xnor U18185 (N_18185,N_17580,N_17794);
or U18186 (N_18186,N_17184,N_17903);
or U18187 (N_18187,N_17051,N_17204);
and U18188 (N_18188,N_17196,N_17891);
nor U18189 (N_18189,N_17896,N_17501);
nor U18190 (N_18190,N_17059,N_17990);
nor U18191 (N_18191,N_17935,N_17092);
nand U18192 (N_18192,N_17782,N_17568);
and U18193 (N_18193,N_17598,N_17970);
xor U18194 (N_18194,N_17276,N_17980);
and U18195 (N_18195,N_17265,N_17082);
nor U18196 (N_18196,N_17116,N_17479);
nor U18197 (N_18197,N_17955,N_17853);
or U18198 (N_18198,N_17986,N_17890);
nand U18199 (N_18199,N_17562,N_17894);
or U18200 (N_18200,N_17554,N_17120);
nor U18201 (N_18201,N_17139,N_17202);
nor U18202 (N_18202,N_17932,N_17586);
nor U18203 (N_18203,N_17668,N_17376);
nand U18204 (N_18204,N_17218,N_17302);
nand U18205 (N_18205,N_17953,N_17371);
and U18206 (N_18206,N_17389,N_17840);
nand U18207 (N_18207,N_17785,N_17600);
nand U18208 (N_18208,N_17292,N_17845);
and U18209 (N_18209,N_17566,N_17974);
xor U18210 (N_18210,N_17238,N_17639);
nand U18211 (N_18211,N_17198,N_17531);
nor U18212 (N_18212,N_17206,N_17941);
or U18213 (N_18213,N_17760,N_17575);
and U18214 (N_18214,N_17699,N_17436);
nor U18215 (N_18215,N_17751,N_17749);
nand U18216 (N_18216,N_17502,N_17469);
nand U18217 (N_18217,N_17614,N_17727);
nor U18218 (N_18218,N_17642,N_17962);
and U18219 (N_18219,N_17880,N_17621);
nand U18220 (N_18220,N_17456,N_17179);
nand U18221 (N_18221,N_17667,N_17108);
or U18222 (N_18222,N_17687,N_17846);
nand U18223 (N_18223,N_17854,N_17852);
xor U18224 (N_18224,N_17251,N_17710);
xnor U18225 (N_18225,N_17358,N_17691);
or U18226 (N_18226,N_17969,N_17285);
nor U18227 (N_18227,N_17478,N_17795);
or U18228 (N_18228,N_17914,N_17422);
xor U18229 (N_18229,N_17560,N_17563);
nand U18230 (N_18230,N_17277,N_17454);
xor U18231 (N_18231,N_17247,N_17555);
xnor U18232 (N_18232,N_17938,N_17083);
or U18233 (N_18233,N_17404,N_17942);
and U18234 (N_18234,N_17384,N_17988);
nand U18235 (N_18235,N_17153,N_17442);
nor U18236 (N_18236,N_17240,N_17881);
xor U18237 (N_18237,N_17065,N_17205);
nor U18238 (N_18238,N_17284,N_17477);
and U18239 (N_18239,N_17320,N_17034);
or U18240 (N_18240,N_17480,N_17619);
or U18241 (N_18241,N_17617,N_17496);
xor U18242 (N_18242,N_17101,N_17352);
xor U18243 (N_18243,N_17446,N_17229);
nand U18244 (N_18244,N_17117,N_17589);
xor U18245 (N_18245,N_17674,N_17033);
and U18246 (N_18246,N_17298,N_17009);
and U18247 (N_18247,N_17388,N_17793);
and U18248 (N_18248,N_17546,N_17288);
and U18249 (N_18249,N_17166,N_17010);
xor U18250 (N_18250,N_17130,N_17638);
nor U18251 (N_18251,N_17379,N_17906);
or U18252 (N_18252,N_17154,N_17272);
nor U18253 (N_18253,N_17998,N_17812);
or U18254 (N_18254,N_17105,N_17263);
nor U18255 (N_18255,N_17385,N_17640);
or U18256 (N_18256,N_17474,N_17873);
nand U18257 (N_18257,N_17096,N_17702);
xnor U18258 (N_18258,N_17864,N_17698);
nor U18259 (N_18259,N_17432,N_17343);
and U18260 (N_18260,N_17337,N_17943);
nand U18261 (N_18261,N_17611,N_17099);
xnor U18262 (N_18262,N_17654,N_17345);
xor U18263 (N_18263,N_17123,N_17473);
and U18264 (N_18264,N_17851,N_17434);
or U18265 (N_18265,N_17122,N_17260);
nor U18266 (N_18266,N_17570,N_17742);
nand U18267 (N_18267,N_17989,N_17008);
or U18268 (N_18268,N_17424,N_17356);
nand U18269 (N_18269,N_17965,N_17912);
and U18270 (N_18270,N_17822,N_17246);
or U18271 (N_18271,N_17507,N_17765);
and U18272 (N_18272,N_17483,N_17539);
and U18273 (N_18273,N_17014,N_17268);
xnor U18274 (N_18274,N_17978,N_17625);
or U18275 (N_18275,N_17533,N_17530);
nand U18276 (N_18276,N_17015,N_17504);
xor U18277 (N_18277,N_17768,N_17809);
and U18278 (N_18278,N_17398,N_17548);
or U18279 (N_18279,N_17992,N_17860);
or U18280 (N_18280,N_17393,N_17079);
or U18281 (N_18281,N_17457,N_17333);
or U18282 (N_18282,N_17774,N_17341);
nor U18283 (N_18283,N_17652,N_17777);
or U18284 (N_18284,N_17606,N_17762);
and U18285 (N_18285,N_17170,N_17390);
or U18286 (N_18286,N_17181,N_17513);
or U18287 (N_18287,N_17237,N_17256);
xor U18288 (N_18288,N_17002,N_17900);
or U18289 (N_18289,N_17857,N_17613);
xnor U18290 (N_18290,N_17486,N_17281);
nor U18291 (N_18291,N_17872,N_17593);
nand U18292 (N_18292,N_17312,N_17315);
or U18293 (N_18293,N_17746,N_17844);
or U18294 (N_18294,N_17420,N_17596);
or U18295 (N_18295,N_17522,N_17073);
nor U18296 (N_18296,N_17391,N_17612);
and U18297 (N_18297,N_17366,N_17893);
and U18298 (N_18298,N_17622,N_17297);
and U18299 (N_18299,N_17717,N_17367);
and U18300 (N_18300,N_17511,N_17294);
nor U18301 (N_18301,N_17094,N_17815);
xnor U18302 (N_18302,N_17437,N_17820);
xor U18303 (N_18303,N_17925,N_17949);
nand U18304 (N_18304,N_17095,N_17887);
nor U18305 (N_18305,N_17147,N_17235);
or U18306 (N_18306,N_17701,N_17730);
nand U18307 (N_18307,N_17868,N_17770);
nand U18308 (N_18308,N_17360,N_17658);
or U18309 (N_18309,N_17975,N_17954);
nand U18310 (N_18310,N_17967,N_17958);
nand U18311 (N_18311,N_17174,N_17944);
and U18312 (N_18312,N_17155,N_17776);
or U18313 (N_18313,N_17630,N_17332);
nand U18314 (N_18314,N_17959,N_17318);
and U18315 (N_18315,N_17786,N_17487);
and U18316 (N_18316,N_17080,N_17892);
nor U18317 (N_18317,N_17695,N_17162);
or U18318 (N_18318,N_17041,N_17088);
nand U18319 (N_18319,N_17342,N_17453);
nand U18320 (N_18320,N_17715,N_17796);
and U18321 (N_18321,N_17207,N_17445);
nor U18322 (N_18322,N_17359,N_17396);
xnor U18323 (N_18323,N_17541,N_17168);
xor U18324 (N_18324,N_17875,N_17335);
and U18325 (N_18325,N_17019,N_17688);
and U18326 (N_18326,N_17330,N_17013);
xnor U18327 (N_18327,N_17788,N_17775);
or U18328 (N_18328,N_17458,N_17254);
or U18329 (N_18329,N_17636,N_17966);
xnor U18330 (N_18330,N_17324,N_17816);
and U18331 (N_18331,N_17527,N_17355);
and U18332 (N_18332,N_17306,N_17847);
nand U18333 (N_18333,N_17534,N_17097);
nor U18334 (N_18334,N_17350,N_17414);
and U18335 (N_18335,N_17451,N_17278);
and U18336 (N_18336,N_17934,N_17450);
nor U18337 (N_18337,N_17357,N_17133);
nand U18338 (N_18338,N_17412,N_17107);
and U18339 (N_18339,N_17754,N_17993);
xnor U18340 (N_18340,N_17321,N_17127);
nor U18341 (N_18341,N_17475,N_17825);
nand U18342 (N_18342,N_17055,N_17591);
nand U18343 (N_18343,N_17747,N_17220);
xnor U18344 (N_18344,N_17650,N_17439);
nand U18345 (N_18345,N_17849,N_17267);
or U18346 (N_18346,N_17889,N_17410);
or U18347 (N_18347,N_17126,N_17981);
nand U18348 (N_18348,N_17447,N_17623);
or U18349 (N_18349,N_17214,N_17273);
nor U18350 (N_18350,N_17005,N_17195);
or U18351 (N_18351,N_17540,N_17470);
or U18352 (N_18352,N_17838,N_17558);
nand U18353 (N_18353,N_17156,N_17602);
and U18354 (N_18354,N_17689,N_17696);
xnor U18355 (N_18355,N_17692,N_17293);
nor U18356 (N_18356,N_17448,N_17635);
xor U18357 (N_18357,N_17049,N_17946);
nor U18358 (N_18358,N_17211,N_17905);
nor U18359 (N_18359,N_17253,N_17736);
nand U18360 (N_18360,N_17983,N_17269);
nand U18361 (N_18361,N_17026,N_17528);
nand U18362 (N_18362,N_17672,N_17823);
or U18363 (N_18363,N_17991,N_17089);
nor U18364 (N_18364,N_17137,N_17948);
and U18365 (N_18365,N_17499,N_17819);
and U18366 (N_18366,N_17058,N_17862);
nand U18367 (N_18367,N_17310,N_17524);
nand U18368 (N_18368,N_17417,N_17608);
and U18369 (N_18369,N_17178,N_17607);
xnor U18370 (N_18370,N_17340,N_17931);
nor U18371 (N_18371,N_17423,N_17173);
or U18372 (N_18372,N_17918,N_17605);
xnor U18373 (N_18373,N_17087,N_17800);
and U18374 (N_18374,N_17394,N_17756);
or U18375 (N_18375,N_17188,N_17811);
or U18376 (N_18376,N_17262,N_17421);
nor U18377 (N_18377,N_17344,N_17492);
and U18378 (N_18378,N_17289,N_17572);
and U18379 (N_18379,N_17933,N_17767);
and U18380 (N_18380,N_17732,N_17425);
and U18381 (N_18381,N_17138,N_17361);
and U18382 (N_18382,N_17091,N_17713);
or U18383 (N_18383,N_17024,N_17271);
nand U18384 (N_18384,N_17419,N_17300);
nor U18385 (N_18385,N_17709,N_17913);
or U18386 (N_18386,N_17401,N_17787);
nand U18387 (N_18387,N_17317,N_17431);
and U18388 (N_18388,N_17515,N_17766);
nand U18389 (N_18389,N_17758,N_17182);
nand U18390 (N_18390,N_17239,N_17910);
nand U18391 (N_18391,N_17030,N_17745);
or U18392 (N_18392,N_17927,N_17062);
or U18393 (N_18393,N_17547,N_17829);
or U18394 (N_18394,N_17301,N_17807);
and U18395 (N_18395,N_17866,N_17244);
or U18396 (N_18396,N_17400,N_17144);
nor U18397 (N_18397,N_17676,N_17995);
xnor U18398 (N_18398,N_17878,N_17046);
nand U18399 (N_18399,N_17928,N_17208);
nor U18400 (N_18400,N_17649,N_17329);
xnor U18401 (N_18401,N_17264,N_17999);
nor U18402 (N_18402,N_17722,N_17861);
nand U18403 (N_18403,N_17233,N_17583);
nor U18404 (N_18404,N_17022,N_17043);
and U18405 (N_18405,N_17841,N_17979);
or U18406 (N_18406,N_17683,N_17693);
and U18407 (N_18407,N_17705,N_17759);
nor U18408 (N_18408,N_17968,N_17368);
nand U18409 (N_18409,N_17951,N_17549);
and U18410 (N_18410,N_17644,N_17171);
and U18411 (N_18411,N_17647,N_17427);
nor U18412 (N_18412,N_17850,N_17641);
or U18413 (N_18413,N_17462,N_17375);
nor U18414 (N_18414,N_17072,N_17032);
nand U18415 (N_18415,N_17347,N_17482);
xor U18416 (N_18416,N_17426,N_17149);
nor U18417 (N_18417,N_17924,N_17865);
nand U18418 (N_18418,N_17678,N_17040);
and U18419 (N_18419,N_17441,N_17810);
nor U18420 (N_18420,N_17697,N_17719);
or U18421 (N_18421,N_17319,N_17653);
nand U18422 (N_18422,N_17879,N_17493);
nor U18423 (N_18423,N_17339,N_17112);
or U18424 (N_18424,N_17711,N_17509);
nor U18425 (N_18425,N_17283,N_17673);
nand U18426 (N_18426,N_17223,N_17354);
or U18427 (N_18427,N_17646,N_17721);
and U18428 (N_18428,N_17444,N_17084);
and U18429 (N_18429,N_17081,N_17365);
and U18430 (N_18430,N_17634,N_17685);
or U18431 (N_18431,N_17778,N_17997);
and U18432 (N_18432,N_17485,N_17827);
nand U18433 (N_18433,N_17733,N_17901);
nor U18434 (N_18434,N_17526,N_17121);
nor U18435 (N_18435,N_17159,N_17459);
and U18436 (N_18436,N_17700,N_17464);
or U18437 (N_18437,N_17628,N_17789);
xor U18438 (N_18438,N_17050,N_17535);
nor U18439 (N_18439,N_17908,N_17380);
and U18440 (N_18440,N_17047,N_17328);
or U18441 (N_18441,N_17408,N_17461);
or U18442 (N_18442,N_17090,N_17257);
xor U18443 (N_18443,N_17764,N_17806);
xnor U18444 (N_18444,N_17187,N_17077);
nor U18445 (N_18445,N_17645,N_17798);
or U18446 (N_18446,N_17771,N_17066);
nor U18447 (N_18447,N_17309,N_17503);
and U18448 (N_18448,N_17378,N_17068);
nor U18449 (N_18449,N_17189,N_17706);
xnor U18450 (N_18450,N_17039,N_17738);
xnor U18451 (N_18451,N_17151,N_17415);
and U18452 (N_18452,N_17323,N_17870);
nor U18453 (N_18453,N_17028,N_17666);
nand U18454 (N_18454,N_17143,N_17100);
xnor U18455 (N_18455,N_17521,N_17140);
nor U18456 (N_18456,N_17690,N_17716);
or U18457 (N_18457,N_17832,N_17648);
and U18458 (N_18458,N_17517,N_17743);
and U18459 (N_18459,N_17416,N_17769);
nand U18460 (N_18460,N_17145,N_17936);
and U18461 (N_18461,N_17987,N_17797);
nor U18462 (N_18462,N_17537,N_17545);
xnor U18463 (N_18463,N_17203,N_17750);
or U18464 (N_18464,N_17601,N_17136);
and U18465 (N_18465,N_17406,N_17052);
or U18466 (N_18466,N_17863,N_17552);
nor U18467 (N_18467,N_17369,N_17542);
and U18468 (N_18468,N_17387,N_17682);
xor U18469 (N_18469,N_17037,N_17067);
nor U18470 (N_18470,N_17270,N_17098);
nor U18471 (N_18471,N_17308,N_17053);
nor U18472 (N_18472,N_17027,N_17550);
or U18473 (N_18473,N_17222,N_17714);
nand U18474 (N_18474,N_17520,N_17551);
and U18475 (N_18475,N_17484,N_17110);
nand U18476 (N_18476,N_17982,N_17916);
xnor U18477 (N_18477,N_17723,N_17183);
and U18478 (N_18478,N_17180,N_17731);
xnor U18479 (N_18479,N_17038,N_17472);
nand U18480 (N_18480,N_17904,N_17488);
nand U18481 (N_18481,N_17856,N_17157);
and U18482 (N_18482,N_17192,N_17226);
xor U18483 (N_18483,N_17409,N_17093);
nor U18484 (N_18484,N_17799,N_17190);
and U18485 (N_18485,N_17971,N_17129);
nand U18486 (N_18486,N_17559,N_17399);
nand U18487 (N_18487,N_17843,N_17316);
or U18488 (N_18488,N_17604,N_17631);
nor U18489 (N_18489,N_17557,N_17303);
nor U18490 (N_18490,N_17172,N_17498);
or U18491 (N_18491,N_17839,N_17212);
nor U18492 (N_18492,N_17023,N_17131);
xor U18493 (N_18493,N_17792,N_17305);
nor U18494 (N_18494,N_17377,N_17048);
nand U18495 (N_18495,N_17599,N_17956);
and U18496 (N_18496,N_17561,N_17594);
nand U18497 (N_18497,N_17681,N_17433);
nand U18498 (N_18498,N_17397,N_17299);
xnor U18499 (N_18499,N_17651,N_17418);
nor U18500 (N_18500,N_17711,N_17490);
and U18501 (N_18501,N_17539,N_17576);
or U18502 (N_18502,N_17486,N_17598);
nand U18503 (N_18503,N_17199,N_17736);
xnor U18504 (N_18504,N_17535,N_17743);
or U18505 (N_18505,N_17038,N_17172);
nand U18506 (N_18506,N_17384,N_17353);
or U18507 (N_18507,N_17110,N_17535);
nor U18508 (N_18508,N_17007,N_17437);
or U18509 (N_18509,N_17183,N_17589);
xor U18510 (N_18510,N_17124,N_17890);
nand U18511 (N_18511,N_17752,N_17715);
or U18512 (N_18512,N_17373,N_17939);
nor U18513 (N_18513,N_17783,N_17937);
xnor U18514 (N_18514,N_17318,N_17121);
xnor U18515 (N_18515,N_17421,N_17036);
nand U18516 (N_18516,N_17845,N_17400);
and U18517 (N_18517,N_17508,N_17469);
or U18518 (N_18518,N_17603,N_17411);
and U18519 (N_18519,N_17864,N_17788);
xor U18520 (N_18520,N_17278,N_17973);
xor U18521 (N_18521,N_17328,N_17399);
or U18522 (N_18522,N_17459,N_17298);
nor U18523 (N_18523,N_17602,N_17770);
nor U18524 (N_18524,N_17554,N_17574);
xnor U18525 (N_18525,N_17395,N_17996);
nor U18526 (N_18526,N_17461,N_17556);
and U18527 (N_18527,N_17211,N_17205);
or U18528 (N_18528,N_17151,N_17234);
nand U18529 (N_18529,N_17362,N_17325);
and U18530 (N_18530,N_17573,N_17892);
or U18531 (N_18531,N_17562,N_17871);
nor U18532 (N_18532,N_17104,N_17536);
xor U18533 (N_18533,N_17893,N_17902);
xnor U18534 (N_18534,N_17540,N_17093);
or U18535 (N_18535,N_17501,N_17109);
or U18536 (N_18536,N_17195,N_17505);
or U18537 (N_18537,N_17280,N_17209);
xnor U18538 (N_18538,N_17100,N_17528);
or U18539 (N_18539,N_17535,N_17012);
nand U18540 (N_18540,N_17017,N_17342);
or U18541 (N_18541,N_17852,N_17308);
nand U18542 (N_18542,N_17854,N_17693);
or U18543 (N_18543,N_17288,N_17671);
or U18544 (N_18544,N_17171,N_17134);
nor U18545 (N_18545,N_17102,N_17942);
xnor U18546 (N_18546,N_17920,N_17599);
or U18547 (N_18547,N_17271,N_17951);
nor U18548 (N_18548,N_17567,N_17020);
and U18549 (N_18549,N_17845,N_17044);
or U18550 (N_18550,N_17744,N_17686);
xor U18551 (N_18551,N_17611,N_17745);
xor U18552 (N_18552,N_17616,N_17537);
and U18553 (N_18553,N_17334,N_17338);
xor U18554 (N_18554,N_17574,N_17837);
xnor U18555 (N_18555,N_17861,N_17657);
and U18556 (N_18556,N_17920,N_17270);
and U18557 (N_18557,N_17514,N_17750);
and U18558 (N_18558,N_17257,N_17093);
or U18559 (N_18559,N_17115,N_17791);
nand U18560 (N_18560,N_17114,N_17082);
nand U18561 (N_18561,N_17877,N_17946);
nor U18562 (N_18562,N_17541,N_17830);
or U18563 (N_18563,N_17918,N_17781);
and U18564 (N_18564,N_17986,N_17446);
xor U18565 (N_18565,N_17872,N_17877);
or U18566 (N_18566,N_17472,N_17524);
and U18567 (N_18567,N_17797,N_17304);
nand U18568 (N_18568,N_17031,N_17198);
nand U18569 (N_18569,N_17069,N_17038);
nor U18570 (N_18570,N_17803,N_17738);
or U18571 (N_18571,N_17234,N_17318);
nor U18572 (N_18572,N_17229,N_17483);
xnor U18573 (N_18573,N_17131,N_17144);
and U18574 (N_18574,N_17870,N_17869);
nand U18575 (N_18575,N_17012,N_17848);
and U18576 (N_18576,N_17259,N_17941);
and U18577 (N_18577,N_17622,N_17386);
and U18578 (N_18578,N_17743,N_17601);
and U18579 (N_18579,N_17063,N_17734);
nand U18580 (N_18580,N_17332,N_17038);
xor U18581 (N_18581,N_17588,N_17510);
xnor U18582 (N_18582,N_17138,N_17286);
nor U18583 (N_18583,N_17937,N_17405);
or U18584 (N_18584,N_17479,N_17935);
and U18585 (N_18585,N_17837,N_17260);
and U18586 (N_18586,N_17580,N_17256);
nand U18587 (N_18587,N_17837,N_17486);
or U18588 (N_18588,N_17180,N_17965);
and U18589 (N_18589,N_17733,N_17333);
nand U18590 (N_18590,N_17633,N_17851);
and U18591 (N_18591,N_17511,N_17099);
and U18592 (N_18592,N_17157,N_17896);
and U18593 (N_18593,N_17132,N_17143);
xnor U18594 (N_18594,N_17806,N_17646);
nand U18595 (N_18595,N_17606,N_17313);
nor U18596 (N_18596,N_17275,N_17325);
nand U18597 (N_18597,N_17695,N_17522);
or U18598 (N_18598,N_17992,N_17956);
and U18599 (N_18599,N_17551,N_17068);
or U18600 (N_18600,N_17990,N_17289);
xor U18601 (N_18601,N_17770,N_17108);
and U18602 (N_18602,N_17088,N_17686);
and U18603 (N_18603,N_17334,N_17295);
nor U18604 (N_18604,N_17889,N_17147);
and U18605 (N_18605,N_17291,N_17376);
nor U18606 (N_18606,N_17452,N_17847);
xor U18607 (N_18607,N_17527,N_17722);
and U18608 (N_18608,N_17432,N_17421);
nor U18609 (N_18609,N_17628,N_17525);
xor U18610 (N_18610,N_17023,N_17472);
nand U18611 (N_18611,N_17640,N_17344);
nand U18612 (N_18612,N_17288,N_17280);
nand U18613 (N_18613,N_17452,N_17694);
xnor U18614 (N_18614,N_17538,N_17648);
xnor U18615 (N_18615,N_17039,N_17155);
nand U18616 (N_18616,N_17549,N_17939);
or U18617 (N_18617,N_17061,N_17004);
and U18618 (N_18618,N_17792,N_17518);
nor U18619 (N_18619,N_17112,N_17782);
or U18620 (N_18620,N_17790,N_17970);
or U18621 (N_18621,N_17516,N_17593);
or U18622 (N_18622,N_17292,N_17238);
xnor U18623 (N_18623,N_17299,N_17482);
nand U18624 (N_18624,N_17838,N_17429);
or U18625 (N_18625,N_17777,N_17638);
xor U18626 (N_18626,N_17189,N_17509);
xor U18627 (N_18627,N_17091,N_17240);
xor U18628 (N_18628,N_17747,N_17671);
nand U18629 (N_18629,N_17090,N_17662);
or U18630 (N_18630,N_17469,N_17517);
nor U18631 (N_18631,N_17975,N_17349);
xor U18632 (N_18632,N_17921,N_17256);
and U18633 (N_18633,N_17451,N_17816);
nand U18634 (N_18634,N_17093,N_17405);
or U18635 (N_18635,N_17700,N_17382);
nor U18636 (N_18636,N_17287,N_17108);
nor U18637 (N_18637,N_17471,N_17353);
and U18638 (N_18638,N_17814,N_17970);
xnor U18639 (N_18639,N_17589,N_17704);
xor U18640 (N_18640,N_17409,N_17926);
or U18641 (N_18641,N_17998,N_17272);
and U18642 (N_18642,N_17361,N_17534);
nor U18643 (N_18643,N_17524,N_17096);
xnor U18644 (N_18644,N_17687,N_17212);
or U18645 (N_18645,N_17269,N_17489);
xnor U18646 (N_18646,N_17448,N_17835);
xor U18647 (N_18647,N_17806,N_17943);
nor U18648 (N_18648,N_17797,N_17278);
nor U18649 (N_18649,N_17095,N_17837);
nand U18650 (N_18650,N_17224,N_17964);
or U18651 (N_18651,N_17674,N_17585);
and U18652 (N_18652,N_17952,N_17932);
nor U18653 (N_18653,N_17140,N_17820);
nor U18654 (N_18654,N_17993,N_17257);
and U18655 (N_18655,N_17724,N_17036);
or U18656 (N_18656,N_17801,N_17671);
and U18657 (N_18657,N_17825,N_17562);
nor U18658 (N_18658,N_17747,N_17748);
nor U18659 (N_18659,N_17163,N_17814);
nor U18660 (N_18660,N_17358,N_17408);
nand U18661 (N_18661,N_17465,N_17457);
and U18662 (N_18662,N_17218,N_17032);
or U18663 (N_18663,N_17773,N_17649);
xor U18664 (N_18664,N_17555,N_17753);
and U18665 (N_18665,N_17759,N_17933);
and U18666 (N_18666,N_17463,N_17081);
and U18667 (N_18667,N_17082,N_17360);
or U18668 (N_18668,N_17848,N_17827);
xnor U18669 (N_18669,N_17478,N_17830);
or U18670 (N_18670,N_17289,N_17564);
nor U18671 (N_18671,N_17253,N_17196);
and U18672 (N_18672,N_17476,N_17612);
or U18673 (N_18673,N_17303,N_17697);
xor U18674 (N_18674,N_17592,N_17299);
nand U18675 (N_18675,N_17167,N_17064);
or U18676 (N_18676,N_17092,N_17091);
or U18677 (N_18677,N_17808,N_17586);
xor U18678 (N_18678,N_17226,N_17983);
nand U18679 (N_18679,N_17413,N_17000);
nor U18680 (N_18680,N_17012,N_17341);
or U18681 (N_18681,N_17125,N_17760);
or U18682 (N_18682,N_17245,N_17085);
and U18683 (N_18683,N_17128,N_17537);
or U18684 (N_18684,N_17384,N_17840);
or U18685 (N_18685,N_17866,N_17879);
xnor U18686 (N_18686,N_17279,N_17477);
nand U18687 (N_18687,N_17796,N_17286);
xor U18688 (N_18688,N_17608,N_17089);
nand U18689 (N_18689,N_17869,N_17952);
nor U18690 (N_18690,N_17974,N_17464);
and U18691 (N_18691,N_17014,N_17481);
xor U18692 (N_18692,N_17509,N_17064);
and U18693 (N_18693,N_17429,N_17140);
or U18694 (N_18694,N_17857,N_17636);
and U18695 (N_18695,N_17363,N_17108);
nor U18696 (N_18696,N_17638,N_17169);
nand U18697 (N_18697,N_17737,N_17821);
nand U18698 (N_18698,N_17163,N_17347);
or U18699 (N_18699,N_17031,N_17813);
xnor U18700 (N_18700,N_17103,N_17959);
nor U18701 (N_18701,N_17907,N_17609);
nand U18702 (N_18702,N_17341,N_17475);
or U18703 (N_18703,N_17023,N_17994);
or U18704 (N_18704,N_17865,N_17191);
and U18705 (N_18705,N_17726,N_17925);
xnor U18706 (N_18706,N_17623,N_17047);
nand U18707 (N_18707,N_17483,N_17498);
nand U18708 (N_18708,N_17997,N_17328);
or U18709 (N_18709,N_17593,N_17008);
nand U18710 (N_18710,N_17123,N_17267);
nor U18711 (N_18711,N_17575,N_17278);
nor U18712 (N_18712,N_17907,N_17505);
nor U18713 (N_18713,N_17600,N_17738);
or U18714 (N_18714,N_17454,N_17596);
xor U18715 (N_18715,N_17001,N_17396);
or U18716 (N_18716,N_17554,N_17648);
and U18717 (N_18717,N_17016,N_17061);
or U18718 (N_18718,N_17468,N_17802);
nand U18719 (N_18719,N_17915,N_17853);
or U18720 (N_18720,N_17378,N_17896);
xor U18721 (N_18721,N_17286,N_17820);
and U18722 (N_18722,N_17055,N_17795);
nor U18723 (N_18723,N_17884,N_17951);
xnor U18724 (N_18724,N_17363,N_17054);
nand U18725 (N_18725,N_17048,N_17089);
and U18726 (N_18726,N_17855,N_17994);
and U18727 (N_18727,N_17150,N_17623);
nor U18728 (N_18728,N_17631,N_17579);
or U18729 (N_18729,N_17176,N_17657);
or U18730 (N_18730,N_17347,N_17599);
nand U18731 (N_18731,N_17677,N_17363);
or U18732 (N_18732,N_17780,N_17011);
or U18733 (N_18733,N_17067,N_17908);
or U18734 (N_18734,N_17239,N_17981);
or U18735 (N_18735,N_17654,N_17295);
nor U18736 (N_18736,N_17228,N_17861);
and U18737 (N_18737,N_17036,N_17081);
or U18738 (N_18738,N_17457,N_17581);
nand U18739 (N_18739,N_17935,N_17860);
xnor U18740 (N_18740,N_17472,N_17104);
and U18741 (N_18741,N_17359,N_17268);
xnor U18742 (N_18742,N_17059,N_17256);
xnor U18743 (N_18743,N_17378,N_17089);
nand U18744 (N_18744,N_17765,N_17031);
nor U18745 (N_18745,N_17447,N_17082);
and U18746 (N_18746,N_17555,N_17346);
nor U18747 (N_18747,N_17993,N_17240);
nand U18748 (N_18748,N_17202,N_17557);
xor U18749 (N_18749,N_17608,N_17781);
xor U18750 (N_18750,N_17041,N_17162);
or U18751 (N_18751,N_17016,N_17818);
nor U18752 (N_18752,N_17669,N_17310);
nor U18753 (N_18753,N_17240,N_17389);
or U18754 (N_18754,N_17253,N_17492);
nand U18755 (N_18755,N_17031,N_17144);
xnor U18756 (N_18756,N_17257,N_17458);
nor U18757 (N_18757,N_17447,N_17302);
nand U18758 (N_18758,N_17621,N_17116);
nand U18759 (N_18759,N_17914,N_17737);
nor U18760 (N_18760,N_17477,N_17095);
and U18761 (N_18761,N_17538,N_17470);
and U18762 (N_18762,N_17299,N_17110);
nand U18763 (N_18763,N_17576,N_17614);
or U18764 (N_18764,N_17207,N_17826);
nand U18765 (N_18765,N_17998,N_17398);
and U18766 (N_18766,N_17629,N_17825);
nor U18767 (N_18767,N_17659,N_17264);
and U18768 (N_18768,N_17880,N_17168);
or U18769 (N_18769,N_17900,N_17418);
and U18770 (N_18770,N_17430,N_17586);
nand U18771 (N_18771,N_17552,N_17230);
nand U18772 (N_18772,N_17089,N_17741);
or U18773 (N_18773,N_17897,N_17440);
and U18774 (N_18774,N_17293,N_17824);
nand U18775 (N_18775,N_17827,N_17336);
nor U18776 (N_18776,N_17710,N_17732);
and U18777 (N_18777,N_17092,N_17814);
xnor U18778 (N_18778,N_17023,N_17774);
and U18779 (N_18779,N_17534,N_17156);
nor U18780 (N_18780,N_17695,N_17291);
xor U18781 (N_18781,N_17524,N_17262);
nor U18782 (N_18782,N_17361,N_17765);
and U18783 (N_18783,N_17923,N_17606);
nand U18784 (N_18784,N_17386,N_17310);
nand U18785 (N_18785,N_17993,N_17071);
nor U18786 (N_18786,N_17557,N_17675);
nor U18787 (N_18787,N_17492,N_17628);
and U18788 (N_18788,N_17325,N_17157);
or U18789 (N_18789,N_17589,N_17511);
nor U18790 (N_18790,N_17635,N_17586);
xnor U18791 (N_18791,N_17381,N_17819);
xnor U18792 (N_18792,N_17007,N_17691);
and U18793 (N_18793,N_17544,N_17575);
nand U18794 (N_18794,N_17229,N_17544);
nand U18795 (N_18795,N_17962,N_17402);
xnor U18796 (N_18796,N_17210,N_17389);
nor U18797 (N_18797,N_17897,N_17898);
and U18798 (N_18798,N_17791,N_17633);
or U18799 (N_18799,N_17716,N_17602);
and U18800 (N_18800,N_17141,N_17154);
and U18801 (N_18801,N_17705,N_17639);
nor U18802 (N_18802,N_17239,N_17209);
nor U18803 (N_18803,N_17164,N_17432);
nand U18804 (N_18804,N_17382,N_17056);
nand U18805 (N_18805,N_17291,N_17756);
xor U18806 (N_18806,N_17245,N_17623);
nor U18807 (N_18807,N_17803,N_17925);
nand U18808 (N_18808,N_17963,N_17545);
xor U18809 (N_18809,N_17876,N_17555);
and U18810 (N_18810,N_17157,N_17824);
and U18811 (N_18811,N_17259,N_17809);
nor U18812 (N_18812,N_17757,N_17201);
and U18813 (N_18813,N_17647,N_17039);
xnor U18814 (N_18814,N_17885,N_17178);
or U18815 (N_18815,N_17472,N_17326);
nor U18816 (N_18816,N_17857,N_17264);
xor U18817 (N_18817,N_17107,N_17269);
or U18818 (N_18818,N_17238,N_17958);
xnor U18819 (N_18819,N_17092,N_17488);
nor U18820 (N_18820,N_17777,N_17129);
xnor U18821 (N_18821,N_17410,N_17933);
and U18822 (N_18822,N_17531,N_17573);
and U18823 (N_18823,N_17275,N_17822);
nor U18824 (N_18824,N_17355,N_17894);
and U18825 (N_18825,N_17855,N_17993);
nand U18826 (N_18826,N_17614,N_17144);
or U18827 (N_18827,N_17724,N_17883);
nand U18828 (N_18828,N_17635,N_17752);
or U18829 (N_18829,N_17438,N_17777);
nor U18830 (N_18830,N_17166,N_17639);
or U18831 (N_18831,N_17828,N_17839);
nor U18832 (N_18832,N_17722,N_17076);
nand U18833 (N_18833,N_17769,N_17581);
nor U18834 (N_18834,N_17336,N_17711);
nand U18835 (N_18835,N_17772,N_17194);
nor U18836 (N_18836,N_17768,N_17467);
nand U18837 (N_18837,N_17359,N_17591);
nand U18838 (N_18838,N_17399,N_17324);
nand U18839 (N_18839,N_17198,N_17714);
xor U18840 (N_18840,N_17781,N_17744);
or U18841 (N_18841,N_17140,N_17237);
nand U18842 (N_18842,N_17302,N_17493);
and U18843 (N_18843,N_17712,N_17087);
nor U18844 (N_18844,N_17462,N_17618);
nor U18845 (N_18845,N_17389,N_17334);
nor U18846 (N_18846,N_17063,N_17287);
or U18847 (N_18847,N_17866,N_17168);
and U18848 (N_18848,N_17048,N_17491);
nand U18849 (N_18849,N_17475,N_17353);
and U18850 (N_18850,N_17090,N_17645);
xor U18851 (N_18851,N_17307,N_17627);
xnor U18852 (N_18852,N_17023,N_17353);
nor U18853 (N_18853,N_17064,N_17421);
and U18854 (N_18854,N_17407,N_17058);
nor U18855 (N_18855,N_17227,N_17168);
xnor U18856 (N_18856,N_17183,N_17515);
nand U18857 (N_18857,N_17567,N_17945);
nor U18858 (N_18858,N_17587,N_17102);
nand U18859 (N_18859,N_17272,N_17624);
or U18860 (N_18860,N_17461,N_17972);
nor U18861 (N_18861,N_17795,N_17430);
and U18862 (N_18862,N_17325,N_17349);
and U18863 (N_18863,N_17708,N_17855);
nand U18864 (N_18864,N_17456,N_17529);
and U18865 (N_18865,N_17518,N_17659);
or U18866 (N_18866,N_17994,N_17496);
or U18867 (N_18867,N_17856,N_17301);
xnor U18868 (N_18868,N_17154,N_17891);
nor U18869 (N_18869,N_17551,N_17903);
xor U18870 (N_18870,N_17690,N_17356);
or U18871 (N_18871,N_17076,N_17226);
nand U18872 (N_18872,N_17976,N_17344);
xnor U18873 (N_18873,N_17268,N_17775);
or U18874 (N_18874,N_17364,N_17137);
or U18875 (N_18875,N_17114,N_17066);
xor U18876 (N_18876,N_17328,N_17756);
nor U18877 (N_18877,N_17558,N_17751);
and U18878 (N_18878,N_17853,N_17462);
nand U18879 (N_18879,N_17098,N_17011);
nor U18880 (N_18880,N_17256,N_17879);
and U18881 (N_18881,N_17338,N_17829);
nand U18882 (N_18882,N_17857,N_17685);
xnor U18883 (N_18883,N_17528,N_17821);
xnor U18884 (N_18884,N_17205,N_17395);
or U18885 (N_18885,N_17693,N_17528);
or U18886 (N_18886,N_17450,N_17763);
xnor U18887 (N_18887,N_17269,N_17639);
and U18888 (N_18888,N_17444,N_17850);
or U18889 (N_18889,N_17545,N_17610);
xor U18890 (N_18890,N_17072,N_17127);
and U18891 (N_18891,N_17923,N_17846);
nor U18892 (N_18892,N_17362,N_17934);
nor U18893 (N_18893,N_17464,N_17635);
xnor U18894 (N_18894,N_17015,N_17212);
xnor U18895 (N_18895,N_17638,N_17324);
nor U18896 (N_18896,N_17466,N_17831);
nand U18897 (N_18897,N_17799,N_17218);
xor U18898 (N_18898,N_17261,N_17461);
nor U18899 (N_18899,N_17192,N_17138);
or U18900 (N_18900,N_17154,N_17217);
nand U18901 (N_18901,N_17121,N_17520);
nand U18902 (N_18902,N_17427,N_17544);
and U18903 (N_18903,N_17236,N_17622);
nor U18904 (N_18904,N_17818,N_17919);
or U18905 (N_18905,N_17060,N_17979);
and U18906 (N_18906,N_17287,N_17075);
xor U18907 (N_18907,N_17779,N_17971);
xnor U18908 (N_18908,N_17592,N_17590);
nor U18909 (N_18909,N_17317,N_17680);
or U18910 (N_18910,N_17771,N_17922);
nor U18911 (N_18911,N_17640,N_17653);
nand U18912 (N_18912,N_17036,N_17037);
nand U18913 (N_18913,N_17362,N_17482);
nor U18914 (N_18914,N_17701,N_17646);
or U18915 (N_18915,N_17496,N_17420);
nand U18916 (N_18916,N_17662,N_17947);
or U18917 (N_18917,N_17074,N_17995);
nand U18918 (N_18918,N_17587,N_17265);
and U18919 (N_18919,N_17860,N_17293);
and U18920 (N_18920,N_17175,N_17988);
nor U18921 (N_18921,N_17010,N_17196);
and U18922 (N_18922,N_17150,N_17185);
or U18923 (N_18923,N_17901,N_17664);
nor U18924 (N_18924,N_17219,N_17012);
and U18925 (N_18925,N_17544,N_17560);
and U18926 (N_18926,N_17743,N_17754);
and U18927 (N_18927,N_17241,N_17627);
nor U18928 (N_18928,N_17939,N_17505);
nor U18929 (N_18929,N_17365,N_17797);
xor U18930 (N_18930,N_17427,N_17113);
nand U18931 (N_18931,N_17013,N_17976);
or U18932 (N_18932,N_17526,N_17314);
nand U18933 (N_18933,N_17278,N_17182);
nand U18934 (N_18934,N_17588,N_17107);
xnor U18935 (N_18935,N_17339,N_17453);
and U18936 (N_18936,N_17470,N_17202);
nand U18937 (N_18937,N_17728,N_17603);
or U18938 (N_18938,N_17401,N_17855);
and U18939 (N_18939,N_17892,N_17507);
nor U18940 (N_18940,N_17487,N_17535);
or U18941 (N_18941,N_17244,N_17932);
or U18942 (N_18942,N_17449,N_17641);
nand U18943 (N_18943,N_17445,N_17706);
and U18944 (N_18944,N_17883,N_17182);
or U18945 (N_18945,N_17354,N_17553);
or U18946 (N_18946,N_17219,N_17305);
nor U18947 (N_18947,N_17162,N_17692);
or U18948 (N_18948,N_17305,N_17569);
nor U18949 (N_18949,N_17374,N_17680);
and U18950 (N_18950,N_17036,N_17093);
or U18951 (N_18951,N_17669,N_17439);
xor U18952 (N_18952,N_17608,N_17487);
or U18953 (N_18953,N_17018,N_17330);
xnor U18954 (N_18954,N_17515,N_17322);
nand U18955 (N_18955,N_17696,N_17984);
or U18956 (N_18956,N_17775,N_17562);
nor U18957 (N_18957,N_17768,N_17000);
nand U18958 (N_18958,N_17756,N_17187);
nor U18959 (N_18959,N_17657,N_17927);
or U18960 (N_18960,N_17811,N_17717);
nand U18961 (N_18961,N_17192,N_17610);
nor U18962 (N_18962,N_17399,N_17491);
nand U18963 (N_18963,N_17452,N_17391);
and U18964 (N_18964,N_17246,N_17307);
nor U18965 (N_18965,N_17153,N_17709);
and U18966 (N_18966,N_17087,N_17040);
nor U18967 (N_18967,N_17130,N_17315);
nand U18968 (N_18968,N_17907,N_17801);
xor U18969 (N_18969,N_17147,N_17799);
xor U18970 (N_18970,N_17087,N_17415);
and U18971 (N_18971,N_17212,N_17311);
or U18972 (N_18972,N_17448,N_17524);
nand U18973 (N_18973,N_17658,N_17624);
xor U18974 (N_18974,N_17869,N_17797);
or U18975 (N_18975,N_17102,N_17484);
nand U18976 (N_18976,N_17502,N_17831);
and U18977 (N_18977,N_17902,N_17720);
and U18978 (N_18978,N_17096,N_17046);
xor U18979 (N_18979,N_17933,N_17008);
and U18980 (N_18980,N_17036,N_17291);
nand U18981 (N_18981,N_17742,N_17712);
and U18982 (N_18982,N_17368,N_17914);
or U18983 (N_18983,N_17937,N_17114);
and U18984 (N_18984,N_17222,N_17102);
and U18985 (N_18985,N_17295,N_17689);
xor U18986 (N_18986,N_17935,N_17574);
xnor U18987 (N_18987,N_17223,N_17838);
xor U18988 (N_18988,N_17681,N_17583);
nand U18989 (N_18989,N_17273,N_17080);
nor U18990 (N_18990,N_17511,N_17448);
nor U18991 (N_18991,N_17469,N_17588);
xor U18992 (N_18992,N_17004,N_17926);
nand U18993 (N_18993,N_17725,N_17631);
and U18994 (N_18994,N_17713,N_17992);
nand U18995 (N_18995,N_17044,N_17119);
xnor U18996 (N_18996,N_17844,N_17449);
or U18997 (N_18997,N_17746,N_17223);
and U18998 (N_18998,N_17435,N_17736);
xnor U18999 (N_18999,N_17619,N_17914);
xor U19000 (N_19000,N_18460,N_18229);
or U19001 (N_19001,N_18785,N_18479);
nor U19002 (N_19002,N_18354,N_18159);
and U19003 (N_19003,N_18459,N_18465);
xnor U19004 (N_19004,N_18601,N_18660);
nor U19005 (N_19005,N_18527,N_18834);
xor U19006 (N_19006,N_18184,N_18273);
nand U19007 (N_19007,N_18338,N_18244);
nor U19008 (N_19008,N_18900,N_18176);
nor U19009 (N_19009,N_18086,N_18635);
and U19010 (N_19010,N_18418,N_18431);
and U19011 (N_19011,N_18061,N_18873);
and U19012 (N_19012,N_18199,N_18435);
nand U19013 (N_19013,N_18943,N_18501);
or U19014 (N_19014,N_18809,N_18571);
nor U19015 (N_19015,N_18742,N_18801);
and U19016 (N_19016,N_18198,N_18220);
nand U19017 (N_19017,N_18657,N_18039);
nand U19018 (N_19018,N_18031,N_18941);
xnor U19019 (N_19019,N_18591,N_18085);
nor U19020 (N_19020,N_18561,N_18679);
and U19021 (N_19021,N_18186,N_18984);
and U19022 (N_19022,N_18293,N_18979);
xnor U19023 (N_19023,N_18971,N_18193);
xnor U19024 (N_19024,N_18934,N_18882);
nor U19025 (N_19025,N_18332,N_18304);
nand U19026 (N_19026,N_18776,N_18544);
nor U19027 (N_19027,N_18973,N_18262);
nor U19028 (N_19028,N_18877,N_18673);
nor U19029 (N_19029,N_18171,N_18274);
xor U19030 (N_19030,N_18416,N_18836);
nand U19031 (N_19031,N_18161,N_18843);
nor U19032 (N_19032,N_18598,N_18030);
nand U19033 (N_19033,N_18556,N_18287);
xnor U19034 (N_19034,N_18384,N_18335);
nand U19035 (N_19035,N_18940,N_18491);
or U19036 (N_19036,N_18683,N_18515);
and U19037 (N_19037,N_18604,N_18275);
xor U19038 (N_19038,N_18207,N_18883);
nor U19039 (N_19039,N_18234,N_18297);
nor U19040 (N_19040,N_18447,N_18745);
xnor U19041 (N_19041,N_18195,N_18254);
xnor U19042 (N_19042,N_18490,N_18853);
nand U19043 (N_19043,N_18811,N_18885);
nand U19044 (N_19044,N_18744,N_18863);
or U19045 (N_19045,N_18210,N_18830);
or U19046 (N_19046,N_18356,N_18305);
xnor U19047 (N_19047,N_18111,N_18956);
nor U19048 (N_19048,N_18955,N_18759);
nor U19049 (N_19049,N_18367,N_18027);
xor U19050 (N_19050,N_18552,N_18125);
or U19051 (N_19051,N_18179,N_18154);
xor U19052 (N_19052,N_18445,N_18052);
nor U19053 (N_19053,N_18730,N_18555);
or U19054 (N_19054,N_18063,N_18768);
and U19055 (N_19055,N_18020,N_18666);
or U19056 (N_19056,N_18642,N_18911);
and U19057 (N_19057,N_18622,N_18688);
xnor U19058 (N_19058,N_18716,N_18046);
nor U19059 (N_19059,N_18923,N_18392);
nand U19060 (N_19060,N_18303,N_18200);
or U19061 (N_19061,N_18441,N_18355);
xor U19062 (N_19062,N_18896,N_18675);
or U19063 (N_19063,N_18053,N_18495);
or U19064 (N_19064,N_18838,N_18764);
xnor U19065 (N_19065,N_18509,N_18954);
or U19066 (N_19066,N_18203,N_18858);
and U19067 (N_19067,N_18467,N_18283);
nand U19068 (N_19068,N_18607,N_18339);
nor U19069 (N_19069,N_18856,N_18708);
xnor U19070 (N_19070,N_18023,N_18074);
or U19071 (N_19071,N_18103,N_18301);
nor U19072 (N_19072,N_18786,N_18081);
xor U19073 (N_19073,N_18728,N_18779);
nand U19074 (N_19074,N_18763,N_18645);
xnor U19075 (N_19075,N_18357,N_18565);
and U19076 (N_19076,N_18288,N_18078);
and U19077 (N_19077,N_18976,N_18379);
nor U19078 (N_19078,N_18420,N_18757);
nor U19079 (N_19079,N_18543,N_18073);
nor U19080 (N_19080,N_18758,N_18483);
xor U19081 (N_19081,N_18450,N_18043);
or U19082 (N_19082,N_18414,N_18985);
or U19083 (N_19083,N_18328,N_18695);
or U19084 (N_19084,N_18071,N_18077);
and U19085 (N_19085,N_18542,N_18098);
or U19086 (N_19086,N_18331,N_18114);
nor U19087 (N_19087,N_18531,N_18204);
xnor U19088 (N_19088,N_18406,N_18549);
or U19089 (N_19089,N_18377,N_18580);
and U19090 (N_19090,N_18336,N_18806);
or U19091 (N_19091,N_18651,N_18163);
and U19092 (N_19092,N_18630,N_18430);
nand U19093 (N_19093,N_18101,N_18022);
nor U19094 (N_19094,N_18484,N_18533);
and U19095 (N_19095,N_18922,N_18284);
or U19096 (N_19096,N_18983,N_18676);
nand U19097 (N_19097,N_18162,N_18686);
or U19098 (N_19098,N_18534,N_18421);
nand U19099 (N_19099,N_18698,N_18032);
and U19100 (N_19100,N_18130,N_18812);
xnor U19101 (N_19101,N_18138,N_18342);
or U19102 (N_19102,N_18831,N_18899);
or U19103 (N_19103,N_18551,N_18021);
xor U19104 (N_19104,N_18146,N_18717);
and U19105 (N_19105,N_18135,N_18385);
and U19106 (N_19106,N_18295,N_18731);
and U19107 (N_19107,N_18257,N_18540);
nor U19108 (N_19108,N_18152,N_18627);
nor U19109 (N_19109,N_18616,N_18564);
and U19110 (N_19110,N_18149,N_18006);
xnor U19111 (N_19111,N_18058,N_18024);
or U19112 (N_19112,N_18326,N_18090);
or U19113 (N_19113,N_18999,N_18783);
nor U19114 (N_19114,N_18548,N_18916);
nor U19115 (N_19115,N_18319,N_18488);
xor U19116 (N_19116,N_18341,N_18833);
xor U19117 (N_19117,N_18394,N_18277);
nand U19118 (N_19118,N_18978,N_18276);
nor U19119 (N_19119,N_18312,N_18183);
nand U19120 (N_19120,N_18076,N_18122);
nand U19121 (N_19121,N_18034,N_18337);
or U19122 (N_19122,N_18787,N_18129);
nor U19123 (N_19123,N_18070,N_18166);
nand U19124 (N_19124,N_18474,N_18844);
nand U19125 (N_19125,N_18360,N_18599);
or U19126 (N_19126,N_18588,N_18835);
nand U19127 (N_19127,N_18422,N_18629);
nor U19128 (N_19128,N_18893,N_18603);
xor U19129 (N_19129,N_18788,N_18123);
xnor U19130 (N_19130,N_18496,N_18790);
or U19131 (N_19131,N_18712,N_18296);
and U19132 (N_19132,N_18938,N_18727);
and U19133 (N_19133,N_18109,N_18753);
nor U19134 (N_19134,N_18401,N_18452);
xor U19135 (N_19135,N_18944,N_18879);
nand U19136 (N_19136,N_18766,N_18316);
xor U19137 (N_19137,N_18674,N_18734);
and U19138 (N_19138,N_18269,N_18765);
and U19139 (N_19139,N_18760,N_18258);
nand U19140 (N_19140,N_18286,N_18915);
or U19141 (N_19141,N_18218,N_18793);
or U19142 (N_19142,N_18263,N_18921);
or U19143 (N_19143,N_18692,N_18614);
or U19144 (N_19144,N_18700,N_18212);
nor U19145 (N_19145,N_18772,N_18167);
nand U19146 (N_19146,N_18443,N_18750);
and U19147 (N_19147,N_18848,N_18550);
nand U19148 (N_19148,N_18347,N_18314);
or U19149 (N_19149,N_18298,N_18409);
xnor U19150 (N_19150,N_18609,N_18088);
or U19151 (N_19151,N_18028,N_18523);
nor U19152 (N_19152,N_18807,N_18637);
and U19153 (N_19153,N_18089,N_18762);
nand U19154 (N_19154,N_18980,N_18127);
nor U19155 (N_19155,N_18775,N_18749);
nor U19156 (N_19156,N_18148,N_18715);
nor U19157 (N_19157,N_18839,N_18823);
nor U19158 (N_19158,N_18315,N_18857);
and U19159 (N_19159,N_18568,N_18155);
and U19160 (N_19160,N_18214,N_18702);
xor U19161 (N_19161,N_18019,N_18663);
and U19162 (N_19162,N_18151,N_18623);
and U19163 (N_19163,N_18850,N_18656);
nor U19164 (N_19164,N_18388,N_18640);
nand U19165 (N_19165,N_18239,N_18577);
nor U19166 (N_19166,N_18570,N_18991);
nor U19167 (N_19167,N_18736,N_18156);
and U19168 (N_19168,N_18875,N_18461);
nor U19169 (N_19169,N_18164,N_18165);
xor U19170 (N_19170,N_18854,N_18080);
or U19171 (N_19171,N_18597,N_18795);
nor U19172 (N_19172,N_18932,N_18141);
nor U19173 (N_19173,N_18815,N_18767);
nand U19174 (N_19174,N_18035,N_18953);
or U19175 (N_19175,N_18366,N_18230);
xnor U19176 (N_19176,N_18824,N_18611);
nor U19177 (N_19177,N_18497,N_18411);
and U19178 (N_19178,N_18661,N_18669);
xnor U19179 (N_19179,N_18721,N_18405);
or U19180 (N_19180,N_18189,N_18937);
or U19181 (N_19181,N_18605,N_18247);
nor U19182 (N_19182,N_18935,N_18398);
or U19183 (N_19183,N_18904,N_18628);
xnor U19184 (N_19184,N_18792,N_18819);
and U19185 (N_19185,N_18102,N_18018);
xor U19186 (N_19186,N_18803,N_18389);
xnor U19187 (N_19187,N_18236,N_18814);
nand U19188 (N_19188,N_18691,N_18572);
nand U19189 (N_19189,N_18351,N_18837);
xnor U19190 (N_19190,N_18248,N_18290);
xnor U19191 (N_19191,N_18905,N_18222);
nand U19192 (N_19192,N_18323,N_18794);
nor U19193 (N_19193,N_18437,N_18910);
nor U19194 (N_19194,N_18476,N_18701);
and U19195 (N_19195,N_18802,N_18124);
xor U19196 (N_19196,N_18927,N_18902);
nor U19197 (N_19197,N_18646,N_18644);
and U19198 (N_19198,N_18499,N_18181);
xor U19199 (N_19199,N_18456,N_18267);
nand U19200 (N_19200,N_18096,N_18260);
nand U19201 (N_19201,N_18782,N_18880);
or U19202 (N_19202,N_18808,N_18002);
nor U19203 (N_19203,N_18348,N_18970);
or U19204 (N_19204,N_18928,N_18116);
and U19205 (N_19205,N_18192,N_18828);
and U19206 (N_19206,N_18737,N_18383);
or U19207 (N_19207,N_18404,N_18864);
nand U19208 (N_19208,N_18751,N_18489);
nor U19209 (N_19209,N_18574,N_18547);
or U19210 (N_19210,N_18374,N_18693);
xor U19211 (N_19211,N_18680,N_18826);
xnor U19212 (N_19212,N_18908,N_18706);
nor U19213 (N_19213,N_18557,N_18829);
xor U19214 (N_19214,N_18209,N_18719);
xor U19215 (N_19215,N_18126,N_18608);
xnor U19216 (N_19216,N_18796,N_18455);
xnor U19217 (N_19217,N_18412,N_18062);
xor U19218 (N_19218,N_18696,N_18237);
nor U19219 (N_19219,N_18517,N_18017);
xor U19220 (N_19220,N_18045,N_18318);
or U19221 (N_19221,N_18579,N_18147);
xnor U19222 (N_19222,N_18739,N_18906);
xnor U19223 (N_19223,N_18486,N_18079);
nand U19224 (N_19224,N_18399,N_18528);
or U19225 (N_19225,N_18137,N_18083);
xnor U19226 (N_19226,N_18475,N_18482);
xnor U19227 (N_19227,N_18641,N_18378);
or U19228 (N_19228,N_18056,N_18989);
and U19229 (N_19229,N_18936,N_18519);
nand U19230 (N_19230,N_18514,N_18748);
and U19231 (N_19231,N_18582,N_18066);
xor U19232 (N_19232,N_18865,N_18894);
and U19233 (N_19233,N_18967,N_18217);
xnor U19234 (N_19234,N_18321,N_18033);
and U19235 (N_19235,N_18402,N_18400);
nand U19236 (N_19236,N_18370,N_18308);
nand U19237 (N_19237,N_18180,N_18330);
or U19238 (N_19238,N_18912,N_18259);
nand U19239 (N_19239,N_18797,N_18117);
nand U19240 (N_19240,N_18131,N_18228);
xnor U19241 (N_19241,N_18747,N_18440);
or U19242 (N_19242,N_18092,N_18363);
and U19243 (N_19243,N_18699,N_18221);
or U19244 (N_19244,N_18995,N_18434);
or U19245 (N_19245,N_18016,N_18325);
nor U19246 (N_19246,N_18202,N_18051);
and U19247 (N_19247,N_18997,N_18177);
nand U19248 (N_19248,N_18920,N_18725);
or U19249 (N_19249,N_18756,N_18648);
xor U19250 (N_19250,N_18242,N_18684);
and U19251 (N_19251,N_18393,N_18966);
and U19252 (N_19252,N_18294,N_18403);
nor U19253 (N_19253,N_18265,N_18919);
or U19254 (N_19254,N_18996,N_18170);
or U19255 (N_19255,N_18633,N_18707);
or U19256 (N_19256,N_18243,N_18852);
nand U19257 (N_19257,N_18008,N_18506);
and U19258 (N_19258,N_18449,N_18726);
nor U19259 (N_19259,N_18494,N_18050);
or U19260 (N_19260,N_18365,N_18187);
nor U19261 (N_19261,N_18235,N_18216);
and U19262 (N_19262,N_18962,N_18458);
and U19263 (N_19263,N_18638,N_18709);
nor U19264 (N_19264,N_18150,N_18867);
and U19265 (N_19265,N_18649,N_18233);
or U19266 (N_19266,N_18282,N_18145);
nor U19267 (N_19267,N_18871,N_18559);
nor U19268 (N_19268,N_18291,N_18545);
xnor U19269 (N_19269,N_18659,N_18593);
nor U19270 (N_19270,N_18329,N_18773);
nand U19271 (N_19271,N_18798,N_18804);
and U19272 (N_19272,N_18949,N_18362);
and U19273 (N_19273,N_18268,N_18653);
nand U19274 (N_19274,N_18225,N_18047);
nand U19275 (N_19275,N_18974,N_18566);
and U19276 (N_19276,N_18194,N_18132);
and U19277 (N_19277,N_18832,N_18947);
nor U19278 (N_19278,N_18897,N_18252);
nand U19279 (N_19279,N_18253,N_18710);
xor U19280 (N_19280,N_18219,N_18480);
xnor U19281 (N_19281,N_18924,N_18818);
nand U19282 (N_19282,N_18168,N_18091);
nand U19283 (N_19283,N_18847,N_18396);
or U19284 (N_19284,N_18780,N_18816);
nand U19285 (N_19285,N_18595,N_18602);
xor U19286 (N_19286,N_18429,N_18413);
or U19287 (N_19287,N_18211,N_18589);
nor U19288 (N_19288,N_18586,N_18986);
and U19289 (N_19289,N_18560,N_18541);
and U19290 (N_19290,N_18391,N_18468);
and U19291 (N_19291,N_18678,N_18596);
nor U19292 (N_19292,N_18261,N_18878);
xnor U19293 (N_19293,N_18600,N_18038);
or U19294 (N_19294,N_18107,N_18432);
nand U19295 (N_19295,N_18278,N_18718);
nand U19296 (N_19296,N_18306,N_18946);
nand U19297 (N_19297,N_18191,N_18245);
xnor U19298 (N_19298,N_18099,N_18606);
and U19299 (N_19299,N_18160,N_18299);
xnor U19300 (N_19300,N_18142,N_18567);
and U19301 (N_19301,N_18036,N_18634);
xnor U19302 (N_19302,N_18082,N_18206);
nand U19303 (N_19303,N_18658,N_18057);
or U19304 (N_19304,N_18505,N_18358);
and U19305 (N_19305,N_18361,N_18397);
or U19306 (N_19306,N_18672,N_18881);
and U19307 (N_19307,N_18761,N_18272);
nor U19308 (N_19308,N_18256,N_18741);
or U19309 (N_19309,N_18842,N_18618);
and U19310 (N_19310,N_18525,N_18959);
xnor U19311 (N_19311,N_18558,N_18375);
nor U19312 (N_19312,N_18419,N_18025);
nor U19313 (N_19313,N_18487,N_18485);
nand U19314 (N_19314,N_18317,N_18553);
nand U19315 (N_19315,N_18887,N_18327);
and U19316 (N_19316,N_18791,N_18872);
and U19317 (N_19317,N_18714,N_18820);
nand U19318 (N_19318,N_18249,N_18895);
and U19319 (N_19319,N_18415,N_18015);
xnor U19320 (N_19320,N_18049,N_18250);
or U19321 (N_19321,N_18914,N_18428);
nor U19322 (N_19322,N_18913,N_18510);
or U19323 (N_19323,N_18581,N_18121);
or U19324 (N_19324,N_18344,N_18011);
nand U19325 (N_19325,N_18255,N_18470);
and U19326 (N_19326,N_18855,N_18067);
nor U19327 (N_19327,N_18992,N_18454);
nand U19328 (N_19328,N_18994,N_18975);
xor U19329 (N_19329,N_18457,N_18583);
or U19330 (N_19330,N_18529,N_18918);
nor U19331 (N_19331,N_18197,N_18439);
xor U19332 (N_19332,N_18563,N_18201);
nand U19333 (N_19333,N_18733,N_18427);
xor U19334 (N_19334,N_18827,N_18113);
and U19335 (N_19335,N_18013,N_18313);
or U19336 (N_19336,N_18650,N_18738);
nor U19337 (N_19337,N_18231,N_18119);
or U19338 (N_19338,N_18903,N_18898);
or U19339 (N_19339,N_18241,N_18746);
or U19340 (N_19340,N_18026,N_18590);
xor U19341 (N_19341,N_18185,N_18068);
nor U19342 (N_19342,N_18516,N_18226);
or U19343 (N_19343,N_18105,N_18215);
nand U19344 (N_19344,N_18526,N_18333);
or U19345 (N_19345,N_18931,N_18869);
xor U19346 (N_19346,N_18442,N_18382);
or U19347 (N_19347,N_18960,N_18535);
xnor U19348 (N_19348,N_18128,N_18810);
nand U19349 (N_19349,N_18538,N_18029);
nand U19350 (N_19350,N_18813,N_18264);
or U19351 (N_19351,N_18613,N_18524);
nor U19352 (N_19352,N_18668,N_18512);
nor U19353 (N_19353,N_18508,N_18961);
and U19354 (N_19354,N_18037,N_18270);
xor U19355 (N_19355,N_18386,N_18311);
nor U19356 (N_19356,N_18532,N_18682);
xnor U19357 (N_19357,N_18310,N_18481);
nand U19358 (N_19358,N_18740,N_18048);
and U19359 (N_19359,N_18448,N_18866);
nand U19360 (N_19360,N_18907,N_18477);
nor U19361 (N_19361,N_18578,N_18845);
nor U19362 (N_19362,N_18720,N_18890);
xnor U19363 (N_19363,N_18575,N_18951);
xnor U19364 (N_19364,N_18968,N_18000);
or U19365 (N_19365,N_18909,N_18594);
and U19366 (N_19366,N_18784,N_18643);
nand U19367 (N_19367,N_18300,N_18350);
and U19368 (N_19368,N_18075,N_18072);
xor U19369 (N_19369,N_18948,N_18988);
xor U19370 (N_19370,N_18945,N_18800);
xor U19371 (N_19371,N_18172,N_18743);
nand U19372 (N_19372,N_18112,N_18500);
nor U19373 (N_19373,N_18340,N_18901);
nor U19374 (N_19374,N_18208,N_18610);
nor U19375 (N_19375,N_18573,N_18530);
xor U19376 (N_19376,N_18417,N_18498);
xor U19377 (N_19377,N_18371,N_18926);
nand U19378 (N_19378,N_18585,N_18592);
or U19379 (N_19379,N_18965,N_18376);
nor U19380 (N_19380,N_18369,N_18054);
or U19381 (N_19381,N_18998,N_18139);
nor U19382 (N_19382,N_18182,N_18095);
or U19383 (N_19383,N_18424,N_18892);
nor U19384 (N_19384,N_18711,N_18677);
nor U19385 (N_19385,N_18463,N_18345);
and U19386 (N_19386,N_18694,N_18817);
nand U19387 (N_19387,N_18636,N_18868);
nand U19388 (N_19388,N_18713,N_18652);
or U19389 (N_19389,N_18120,N_18009);
nand U19390 (N_19390,N_18473,N_18562);
or U19391 (N_19391,N_18118,N_18410);
or U19392 (N_19392,N_18860,N_18140);
nand U19393 (N_19393,N_18735,N_18723);
and U19394 (N_19394,N_18175,N_18925);
or U19395 (N_19395,N_18939,N_18849);
nor U19396 (N_19396,N_18064,N_18466);
nand U19397 (N_19397,N_18755,N_18841);
nor U19398 (N_19398,N_18874,N_18408);
or U19399 (N_19399,N_18732,N_18930);
or U19400 (N_19400,N_18681,N_18617);
nor U19401 (N_19401,N_18624,N_18670);
nand U19402 (N_19402,N_18972,N_18087);
and U19403 (N_19403,N_18292,N_18188);
nand U19404 (N_19404,N_18825,N_18359);
and U19405 (N_19405,N_18352,N_18232);
nand U19406 (N_19406,N_18324,N_18639);
and U19407 (N_19407,N_18513,N_18504);
and U19408 (N_19408,N_18722,N_18704);
xor U19409 (N_19409,N_18134,N_18042);
xor U19410 (N_19410,N_18001,N_18821);
and U19411 (N_19411,N_18917,N_18060);
nor U19412 (N_19412,N_18368,N_18280);
or U19413 (N_19413,N_18343,N_18289);
or U19414 (N_19414,N_18334,N_18407);
nor U19415 (N_19415,N_18446,N_18133);
or U19416 (N_19416,N_18227,N_18539);
nor U19417 (N_19417,N_18472,N_18781);
xor U19418 (N_19418,N_18390,N_18667);
nand U19419 (N_19419,N_18840,N_18004);
or U19420 (N_19420,N_18507,N_18144);
nor U19421 (N_19421,N_18576,N_18870);
or U19422 (N_19422,N_18536,N_18502);
nor U19423 (N_19423,N_18822,N_18662);
xor U19424 (N_19424,N_18223,N_18805);
xor U19425 (N_19425,N_18381,N_18626);
nor U19426 (N_19426,N_18521,N_18655);
and U19427 (N_19427,N_18353,N_18309);
nor U19428 (N_19428,N_18373,N_18625);
nand U19429 (N_19429,N_18520,N_18349);
xnor U19430 (N_19430,N_18569,N_18307);
xor U19431 (N_19431,N_18007,N_18647);
and U19432 (N_19432,N_18136,N_18040);
nand U19433 (N_19433,N_18778,N_18157);
or U19434 (N_19434,N_18685,N_18158);
xor U19435 (N_19435,N_18729,N_18689);
xor U19436 (N_19436,N_18665,N_18703);
nor U19437 (N_19437,N_18453,N_18859);
and U19438 (N_19438,N_18436,N_18364);
and U19439 (N_19439,N_18451,N_18774);
nor U19440 (N_19440,N_18093,N_18205);
xnor U19441 (N_19441,N_18478,N_18469);
or U19442 (N_19442,N_18884,N_18503);
or U19443 (N_19443,N_18889,N_18380);
or U19444 (N_19444,N_18993,N_18433);
nor U19445 (N_19445,N_18554,N_18438);
nand U19446 (N_19446,N_18097,N_18612);
nor U19447 (N_19447,N_18084,N_18464);
nand U19448 (N_19448,N_18546,N_18518);
nor U19449 (N_19449,N_18003,N_18279);
nor U19450 (N_19450,N_18423,N_18108);
nor U19451 (N_19451,N_18963,N_18977);
nand U19452 (N_19452,N_18982,N_18104);
and U19453 (N_19453,N_18621,N_18705);
and U19454 (N_19454,N_18876,N_18322);
and U19455 (N_19455,N_18846,N_18511);
nand U19456 (N_19456,N_18690,N_18471);
nor U19457 (N_19457,N_18537,N_18789);
nand U19458 (N_19458,N_18632,N_18224);
xnor U19459 (N_19459,N_18271,N_18266);
xnor U19460 (N_19460,N_18664,N_18957);
or U19461 (N_19461,N_18929,N_18990);
nand U19462 (N_19462,N_18886,N_18861);
nor U19463 (N_19463,N_18115,N_18770);
nor U19464 (N_19464,N_18654,N_18281);
nor U19465 (N_19465,N_18987,N_18587);
nor U19466 (N_19466,N_18615,N_18754);
nor U19467 (N_19467,N_18981,N_18320);
nand U19468 (N_19468,N_18395,N_18799);
nor U19469 (N_19469,N_18190,N_18425);
xnor U19470 (N_19470,N_18933,N_18769);
and U19471 (N_19471,N_18251,N_18462);
or U19472 (N_19472,N_18238,N_18196);
or U19473 (N_19473,N_18041,N_18619);
nand U19474 (N_19474,N_18620,N_18246);
xnor U19475 (N_19475,N_18952,N_18106);
xor U19476 (N_19476,N_18143,N_18426);
xnor U19477 (N_19477,N_18942,N_18169);
nor U19478 (N_19478,N_18891,N_18958);
and U19479 (N_19479,N_18372,N_18173);
and U19480 (N_19480,N_18014,N_18724);
nor U19481 (N_19481,N_18010,N_18100);
xnor U19482 (N_19482,N_18777,N_18752);
nor U19483 (N_19483,N_18012,N_18285);
and U19484 (N_19484,N_18005,N_18044);
nand U19485 (N_19485,N_18697,N_18178);
and U19486 (N_19486,N_18771,N_18240);
nand U19487 (N_19487,N_18444,N_18069);
or U19488 (N_19488,N_18492,N_18174);
nand U19489 (N_19489,N_18631,N_18964);
nor U19490 (N_19490,N_18851,N_18059);
nor U19491 (N_19491,N_18055,N_18493);
or U19492 (N_19492,N_18687,N_18213);
and U19493 (N_19493,N_18969,N_18110);
nor U19494 (N_19494,N_18522,N_18153);
nand U19495 (N_19495,N_18950,N_18065);
nor U19496 (N_19496,N_18346,N_18584);
and U19497 (N_19497,N_18387,N_18888);
xor U19498 (N_19498,N_18671,N_18302);
or U19499 (N_19499,N_18862,N_18094);
xnor U19500 (N_19500,N_18681,N_18161);
nor U19501 (N_19501,N_18793,N_18252);
xnor U19502 (N_19502,N_18995,N_18832);
nand U19503 (N_19503,N_18825,N_18735);
nor U19504 (N_19504,N_18053,N_18241);
nand U19505 (N_19505,N_18084,N_18334);
nand U19506 (N_19506,N_18304,N_18701);
and U19507 (N_19507,N_18765,N_18166);
nor U19508 (N_19508,N_18791,N_18617);
nand U19509 (N_19509,N_18131,N_18360);
nor U19510 (N_19510,N_18138,N_18587);
or U19511 (N_19511,N_18676,N_18866);
xor U19512 (N_19512,N_18343,N_18439);
nand U19513 (N_19513,N_18999,N_18591);
or U19514 (N_19514,N_18706,N_18645);
and U19515 (N_19515,N_18879,N_18431);
or U19516 (N_19516,N_18723,N_18778);
xnor U19517 (N_19517,N_18060,N_18314);
and U19518 (N_19518,N_18754,N_18044);
or U19519 (N_19519,N_18141,N_18568);
or U19520 (N_19520,N_18176,N_18595);
xor U19521 (N_19521,N_18771,N_18302);
or U19522 (N_19522,N_18461,N_18090);
nor U19523 (N_19523,N_18362,N_18819);
or U19524 (N_19524,N_18665,N_18976);
nor U19525 (N_19525,N_18277,N_18862);
nor U19526 (N_19526,N_18952,N_18810);
and U19527 (N_19527,N_18735,N_18626);
nand U19528 (N_19528,N_18025,N_18438);
and U19529 (N_19529,N_18551,N_18171);
nor U19530 (N_19530,N_18998,N_18167);
nor U19531 (N_19531,N_18574,N_18463);
xnor U19532 (N_19532,N_18609,N_18141);
and U19533 (N_19533,N_18643,N_18105);
nand U19534 (N_19534,N_18456,N_18507);
xor U19535 (N_19535,N_18334,N_18758);
or U19536 (N_19536,N_18568,N_18618);
xor U19537 (N_19537,N_18198,N_18371);
nor U19538 (N_19538,N_18990,N_18810);
or U19539 (N_19539,N_18499,N_18482);
and U19540 (N_19540,N_18489,N_18247);
xnor U19541 (N_19541,N_18940,N_18885);
nand U19542 (N_19542,N_18008,N_18949);
or U19543 (N_19543,N_18406,N_18453);
xnor U19544 (N_19544,N_18997,N_18819);
or U19545 (N_19545,N_18228,N_18071);
xor U19546 (N_19546,N_18624,N_18040);
nand U19547 (N_19547,N_18966,N_18037);
or U19548 (N_19548,N_18101,N_18340);
or U19549 (N_19549,N_18460,N_18580);
or U19550 (N_19550,N_18115,N_18254);
or U19551 (N_19551,N_18964,N_18537);
and U19552 (N_19552,N_18746,N_18228);
nor U19553 (N_19553,N_18606,N_18550);
and U19554 (N_19554,N_18224,N_18516);
or U19555 (N_19555,N_18846,N_18460);
or U19556 (N_19556,N_18568,N_18457);
nand U19557 (N_19557,N_18471,N_18561);
nor U19558 (N_19558,N_18454,N_18779);
xnor U19559 (N_19559,N_18671,N_18076);
xor U19560 (N_19560,N_18193,N_18423);
and U19561 (N_19561,N_18802,N_18761);
nor U19562 (N_19562,N_18446,N_18481);
nor U19563 (N_19563,N_18594,N_18053);
or U19564 (N_19564,N_18536,N_18273);
and U19565 (N_19565,N_18961,N_18375);
and U19566 (N_19566,N_18304,N_18559);
xnor U19567 (N_19567,N_18396,N_18733);
nor U19568 (N_19568,N_18636,N_18218);
and U19569 (N_19569,N_18607,N_18560);
or U19570 (N_19570,N_18463,N_18610);
and U19571 (N_19571,N_18255,N_18827);
nor U19572 (N_19572,N_18358,N_18089);
nand U19573 (N_19573,N_18459,N_18533);
and U19574 (N_19574,N_18011,N_18832);
and U19575 (N_19575,N_18449,N_18344);
xor U19576 (N_19576,N_18807,N_18411);
nand U19577 (N_19577,N_18419,N_18213);
and U19578 (N_19578,N_18106,N_18353);
and U19579 (N_19579,N_18144,N_18655);
nand U19580 (N_19580,N_18568,N_18145);
and U19581 (N_19581,N_18431,N_18616);
nand U19582 (N_19582,N_18867,N_18197);
and U19583 (N_19583,N_18800,N_18397);
nor U19584 (N_19584,N_18360,N_18272);
or U19585 (N_19585,N_18869,N_18143);
nand U19586 (N_19586,N_18044,N_18758);
xor U19587 (N_19587,N_18187,N_18313);
and U19588 (N_19588,N_18011,N_18340);
or U19589 (N_19589,N_18137,N_18273);
or U19590 (N_19590,N_18463,N_18416);
nor U19591 (N_19591,N_18974,N_18885);
nand U19592 (N_19592,N_18601,N_18158);
and U19593 (N_19593,N_18693,N_18446);
or U19594 (N_19594,N_18452,N_18942);
nor U19595 (N_19595,N_18096,N_18259);
nor U19596 (N_19596,N_18333,N_18495);
nand U19597 (N_19597,N_18640,N_18455);
and U19598 (N_19598,N_18451,N_18174);
and U19599 (N_19599,N_18718,N_18437);
nand U19600 (N_19600,N_18178,N_18143);
xor U19601 (N_19601,N_18440,N_18960);
and U19602 (N_19602,N_18891,N_18822);
nor U19603 (N_19603,N_18726,N_18265);
xor U19604 (N_19604,N_18656,N_18922);
and U19605 (N_19605,N_18580,N_18122);
or U19606 (N_19606,N_18930,N_18459);
or U19607 (N_19607,N_18850,N_18728);
and U19608 (N_19608,N_18952,N_18752);
nor U19609 (N_19609,N_18486,N_18668);
or U19610 (N_19610,N_18079,N_18994);
nor U19611 (N_19611,N_18936,N_18794);
nand U19612 (N_19612,N_18235,N_18103);
and U19613 (N_19613,N_18557,N_18841);
and U19614 (N_19614,N_18947,N_18572);
or U19615 (N_19615,N_18073,N_18917);
nor U19616 (N_19616,N_18036,N_18737);
or U19617 (N_19617,N_18785,N_18444);
nand U19618 (N_19618,N_18302,N_18712);
nand U19619 (N_19619,N_18110,N_18529);
xnor U19620 (N_19620,N_18418,N_18482);
or U19621 (N_19621,N_18455,N_18328);
xor U19622 (N_19622,N_18963,N_18086);
nand U19623 (N_19623,N_18848,N_18062);
nor U19624 (N_19624,N_18569,N_18970);
nor U19625 (N_19625,N_18739,N_18684);
nor U19626 (N_19626,N_18286,N_18716);
xor U19627 (N_19627,N_18656,N_18967);
nand U19628 (N_19628,N_18648,N_18043);
and U19629 (N_19629,N_18723,N_18155);
and U19630 (N_19630,N_18817,N_18401);
nand U19631 (N_19631,N_18934,N_18916);
or U19632 (N_19632,N_18245,N_18141);
nand U19633 (N_19633,N_18918,N_18798);
nand U19634 (N_19634,N_18241,N_18041);
nor U19635 (N_19635,N_18718,N_18482);
xnor U19636 (N_19636,N_18934,N_18586);
nor U19637 (N_19637,N_18482,N_18094);
and U19638 (N_19638,N_18091,N_18361);
and U19639 (N_19639,N_18349,N_18950);
nand U19640 (N_19640,N_18130,N_18841);
and U19641 (N_19641,N_18846,N_18196);
nor U19642 (N_19642,N_18585,N_18213);
nor U19643 (N_19643,N_18511,N_18290);
or U19644 (N_19644,N_18512,N_18034);
nor U19645 (N_19645,N_18520,N_18371);
and U19646 (N_19646,N_18135,N_18803);
xor U19647 (N_19647,N_18466,N_18384);
or U19648 (N_19648,N_18657,N_18511);
and U19649 (N_19649,N_18441,N_18246);
nand U19650 (N_19650,N_18650,N_18856);
or U19651 (N_19651,N_18535,N_18688);
and U19652 (N_19652,N_18218,N_18916);
nand U19653 (N_19653,N_18028,N_18824);
xnor U19654 (N_19654,N_18757,N_18696);
or U19655 (N_19655,N_18987,N_18390);
and U19656 (N_19656,N_18859,N_18204);
nand U19657 (N_19657,N_18307,N_18853);
nand U19658 (N_19658,N_18991,N_18174);
nand U19659 (N_19659,N_18771,N_18376);
nand U19660 (N_19660,N_18774,N_18819);
nand U19661 (N_19661,N_18483,N_18313);
or U19662 (N_19662,N_18619,N_18154);
nand U19663 (N_19663,N_18061,N_18066);
nand U19664 (N_19664,N_18542,N_18589);
or U19665 (N_19665,N_18934,N_18764);
and U19666 (N_19666,N_18844,N_18851);
xor U19667 (N_19667,N_18842,N_18753);
nor U19668 (N_19668,N_18081,N_18218);
and U19669 (N_19669,N_18152,N_18909);
or U19670 (N_19670,N_18163,N_18938);
and U19671 (N_19671,N_18867,N_18225);
nor U19672 (N_19672,N_18759,N_18143);
or U19673 (N_19673,N_18086,N_18074);
xor U19674 (N_19674,N_18035,N_18177);
xor U19675 (N_19675,N_18904,N_18102);
nand U19676 (N_19676,N_18520,N_18820);
and U19677 (N_19677,N_18970,N_18989);
xor U19678 (N_19678,N_18212,N_18156);
xor U19679 (N_19679,N_18661,N_18087);
xnor U19680 (N_19680,N_18489,N_18253);
xnor U19681 (N_19681,N_18657,N_18710);
and U19682 (N_19682,N_18661,N_18362);
and U19683 (N_19683,N_18896,N_18023);
or U19684 (N_19684,N_18840,N_18005);
nand U19685 (N_19685,N_18159,N_18654);
or U19686 (N_19686,N_18012,N_18847);
or U19687 (N_19687,N_18134,N_18141);
nor U19688 (N_19688,N_18680,N_18799);
xor U19689 (N_19689,N_18374,N_18230);
or U19690 (N_19690,N_18520,N_18348);
or U19691 (N_19691,N_18347,N_18289);
or U19692 (N_19692,N_18984,N_18866);
xnor U19693 (N_19693,N_18665,N_18133);
and U19694 (N_19694,N_18415,N_18515);
xor U19695 (N_19695,N_18973,N_18607);
nor U19696 (N_19696,N_18103,N_18487);
or U19697 (N_19697,N_18667,N_18436);
nor U19698 (N_19698,N_18020,N_18171);
nor U19699 (N_19699,N_18426,N_18338);
or U19700 (N_19700,N_18447,N_18444);
or U19701 (N_19701,N_18982,N_18517);
or U19702 (N_19702,N_18589,N_18919);
nand U19703 (N_19703,N_18863,N_18469);
and U19704 (N_19704,N_18747,N_18258);
and U19705 (N_19705,N_18169,N_18569);
nand U19706 (N_19706,N_18041,N_18548);
nor U19707 (N_19707,N_18118,N_18658);
nand U19708 (N_19708,N_18309,N_18514);
and U19709 (N_19709,N_18201,N_18151);
xor U19710 (N_19710,N_18045,N_18766);
nor U19711 (N_19711,N_18375,N_18960);
nor U19712 (N_19712,N_18365,N_18916);
nand U19713 (N_19713,N_18556,N_18183);
xor U19714 (N_19714,N_18085,N_18326);
nand U19715 (N_19715,N_18401,N_18664);
and U19716 (N_19716,N_18997,N_18868);
nand U19717 (N_19717,N_18863,N_18038);
xnor U19718 (N_19718,N_18391,N_18547);
and U19719 (N_19719,N_18140,N_18961);
or U19720 (N_19720,N_18838,N_18664);
xor U19721 (N_19721,N_18425,N_18474);
nor U19722 (N_19722,N_18037,N_18482);
xnor U19723 (N_19723,N_18550,N_18815);
and U19724 (N_19724,N_18288,N_18307);
and U19725 (N_19725,N_18224,N_18939);
or U19726 (N_19726,N_18642,N_18393);
nand U19727 (N_19727,N_18374,N_18673);
nor U19728 (N_19728,N_18682,N_18024);
nor U19729 (N_19729,N_18702,N_18357);
xor U19730 (N_19730,N_18266,N_18999);
nor U19731 (N_19731,N_18713,N_18269);
or U19732 (N_19732,N_18210,N_18325);
nand U19733 (N_19733,N_18780,N_18257);
xor U19734 (N_19734,N_18028,N_18235);
or U19735 (N_19735,N_18734,N_18271);
or U19736 (N_19736,N_18530,N_18202);
and U19737 (N_19737,N_18352,N_18733);
nor U19738 (N_19738,N_18481,N_18724);
or U19739 (N_19739,N_18207,N_18073);
nand U19740 (N_19740,N_18813,N_18781);
nor U19741 (N_19741,N_18406,N_18515);
and U19742 (N_19742,N_18109,N_18682);
or U19743 (N_19743,N_18377,N_18803);
nand U19744 (N_19744,N_18472,N_18140);
xnor U19745 (N_19745,N_18993,N_18629);
or U19746 (N_19746,N_18665,N_18405);
and U19747 (N_19747,N_18664,N_18931);
xnor U19748 (N_19748,N_18051,N_18675);
nor U19749 (N_19749,N_18359,N_18007);
nand U19750 (N_19750,N_18117,N_18602);
or U19751 (N_19751,N_18256,N_18586);
nand U19752 (N_19752,N_18256,N_18045);
and U19753 (N_19753,N_18735,N_18694);
xnor U19754 (N_19754,N_18211,N_18462);
nor U19755 (N_19755,N_18037,N_18457);
nor U19756 (N_19756,N_18804,N_18103);
xor U19757 (N_19757,N_18904,N_18014);
nor U19758 (N_19758,N_18896,N_18222);
nor U19759 (N_19759,N_18427,N_18451);
or U19760 (N_19760,N_18322,N_18199);
and U19761 (N_19761,N_18887,N_18908);
and U19762 (N_19762,N_18189,N_18053);
or U19763 (N_19763,N_18932,N_18616);
or U19764 (N_19764,N_18705,N_18168);
and U19765 (N_19765,N_18554,N_18848);
nand U19766 (N_19766,N_18180,N_18952);
or U19767 (N_19767,N_18620,N_18685);
nand U19768 (N_19768,N_18727,N_18950);
xor U19769 (N_19769,N_18721,N_18540);
and U19770 (N_19770,N_18828,N_18284);
nand U19771 (N_19771,N_18869,N_18669);
xor U19772 (N_19772,N_18162,N_18727);
and U19773 (N_19773,N_18453,N_18315);
or U19774 (N_19774,N_18509,N_18337);
nor U19775 (N_19775,N_18421,N_18007);
or U19776 (N_19776,N_18589,N_18558);
nor U19777 (N_19777,N_18953,N_18268);
and U19778 (N_19778,N_18328,N_18236);
nand U19779 (N_19779,N_18101,N_18748);
and U19780 (N_19780,N_18123,N_18236);
and U19781 (N_19781,N_18473,N_18731);
and U19782 (N_19782,N_18928,N_18958);
xor U19783 (N_19783,N_18902,N_18418);
nand U19784 (N_19784,N_18669,N_18082);
or U19785 (N_19785,N_18373,N_18828);
xnor U19786 (N_19786,N_18836,N_18855);
nand U19787 (N_19787,N_18266,N_18524);
nand U19788 (N_19788,N_18507,N_18527);
nor U19789 (N_19789,N_18285,N_18552);
and U19790 (N_19790,N_18123,N_18599);
xnor U19791 (N_19791,N_18601,N_18874);
xor U19792 (N_19792,N_18004,N_18082);
nand U19793 (N_19793,N_18506,N_18890);
xnor U19794 (N_19794,N_18457,N_18720);
nor U19795 (N_19795,N_18500,N_18910);
or U19796 (N_19796,N_18015,N_18371);
or U19797 (N_19797,N_18264,N_18864);
and U19798 (N_19798,N_18057,N_18617);
xor U19799 (N_19799,N_18122,N_18435);
nor U19800 (N_19800,N_18750,N_18853);
or U19801 (N_19801,N_18588,N_18489);
or U19802 (N_19802,N_18721,N_18593);
nor U19803 (N_19803,N_18115,N_18079);
xor U19804 (N_19804,N_18628,N_18341);
or U19805 (N_19805,N_18323,N_18718);
or U19806 (N_19806,N_18831,N_18112);
and U19807 (N_19807,N_18050,N_18914);
and U19808 (N_19808,N_18025,N_18145);
nor U19809 (N_19809,N_18836,N_18334);
or U19810 (N_19810,N_18599,N_18092);
and U19811 (N_19811,N_18933,N_18175);
nor U19812 (N_19812,N_18790,N_18015);
nand U19813 (N_19813,N_18170,N_18760);
xnor U19814 (N_19814,N_18502,N_18266);
or U19815 (N_19815,N_18769,N_18790);
and U19816 (N_19816,N_18032,N_18557);
or U19817 (N_19817,N_18637,N_18857);
xnor U19818 (N_19818,N_18322,N_18908);
nand U19819 (N_19819,N_18658,N_18957);
nand U19820 (N_19820,N_18775,N_18535);
nand U19821 (N_19821,N_18963,N_18690);
or U19822 (N_19822,N_18404,N_18793);
and U19823 (N_19823,N_18683,N_18437);
or U19824 (N_19824,N_18527,N_18739);
xor U19825 (N_19825,N_18962,N_18149);
and U19826 (N_19826,N_18592,N_18104);
or U19827 (N_19827,N_18604,N_18028);
nor U19828 (N_19828,N_18723,N_18724);
nor U19829 (N_19829,N_18136,N_18534);
or U19830 (N_19830,N_18933,N_18068);
xor U19831 (N_19831,N_18930,N_18221);
and U19832 (N_19832,N_18680,N_18779);
and U19833 (N_19833,N_18896,N_18184);
nand U19834 (N_19834,N_18305,N_18809);
nor U19835 (N_19835,N_18531,N_18515);
nand U19836 (N_19836,N_18362,N_18262);
nand U19837 (N_19837,N_18432,N_18080);
nand U19838 (N_19838,N_18340,N_18774);
nand U19839 (N_19839,N_18582,N_18967);
and U19840 (N_19840,N_18175,N_18758);
or U19841 (N_19841,N_18895,N_18220);
xor U19842 (N_19842,N_18299,N_18055);
xor U19843 (N_19843,N_18252,N_18554);
xnor U19844 (N_19844,N_18468,N_18455);
and U19845 (N_19845,N_18102,N_18444);
nor U19846 (N_19846,N_18152,N_18771);
nand U19847 (N_19847,N_18033,N_18115);
or U19848 (N_19848,N_18736,N_18781);
and U19849 (N_19849,N_18473,N_18732);
and U19850 (N_19850,N_18356,N_18339);
xnor U19851 (N_19851,N_18395,N_18538);
nor U19852 (N_19852,N_18169,N_18026);
and U19853 (N_19853,N_18859,N_18443);
nor U19854 (N_19854,N_18613,N_18772);
nor U19855 (N_19855,N_18614,N_18541);
nand U19856 (N_19856,N_18836,N_18345);
and U19857 (N_19857,N_18102,N_18997);
or U19858 (N_19858,N_18172,N_18109);
and U19859 (N_19859,N_18721,N_18272);
xor U19860 (N_19860,N_18955,N_18561);
or U19861 (N_19861,N_18252,N_18487);
xor U19862 (N_19862,N_18472,N_18778);
xor U19863 (N_19863,N_18024,N_18916);
xnor U19864 (N_19864,N_18079,N_18310);
or U19865 (N_19865,N_18437,N_18207);
and U19866 (N_19866,N_18524,N_18516);
nor U19867 (N_19867,N_18657,N_18897);
nand U19868 (N_19868,N_18528,N_18836);
xor U19869 (N_19869,N_18044,N_18267);
nor U19870 (N_19870,N_18948,N_18503);
and U19871 (N_19871,N_18807,N_18562);
and U19872 (N_19872,N_18639,N_18284);
nand U19873 (N_19873,N_18138,N_18762);
nand U19874 (N_19874,N_18213,N_18111);
nand U19875 (N_19875,N_18861,N_18609);
nand U19876 (N_19876,N_18247,N_18892);
nor U19877 (N_19877,N_18421,N_18676);
or U19878 (N_19878,N_18902,N_18750);
or U19879 (N_19879,N_18775,N_18395);
nand U19880 (N_19880,N_18590,N_18725);
and U19881 (N_19881,N_18495,N_18849);
nand U19882 (N_19882,N_18852,N_18948);
xor U19883 (N_19883,N_18102,N_18558);
nand U19884 (N_19884,N_18714,N_18413);
xor U19885 (N_19885,N_18138,N_18581);
xnor U19886 (N_19886,N_18185,N_18648);
or U19887 (N_19887,N_18562,N_18202);
or U19888 (N_19888,N_18226,N_18348);
xnor U19889 (N_19889,N_18811,N_18054);
xnor U19890 (N_19890,N_18010,N_18418);
and U19891 (N_19891,N_18206,N_18500);
nand U19892 (N_19892,N_18849,N_18385);
nand U19893 (N_19893,N_18528,N_18987);
xor U19894 (N_19894,N_18439,N_18703);
xor U19895 (N_19895,N_18584,N_18873);
or U19896 (N_19896,N_18745,N_18744);
and U19897 (N_19897,N_18239,N_18889);
nand U19898 (N_19898,N_18868,N_18947);
nand U19899 (N_19899,N_18810,N_18711);
and U19900 (N_19900,N_18831,N_18677);
and U19901 (N_19901,N_18114,N_18207);
or U19902 (N_19902,N_18788,N_18264);
and U19903 (N_19903,N_18584,N_18792);
nor U19904 (N_19904,N_18620,N_18416);
nand U19905 (N_19905,N_18858,N_18144);
xor U19906 (N_19906,N_18161,N_18781);
nand U19907 (N_19907,N_18979,N_18143);
xor U19908 (N_19908,N_18841,N_18493);
or U19909 (N_19909,N_18033,N_18822);
nor U19910 (N_19910,N_18673,N_18019);
and U19911 (N_19911,N_18239,N_18232);
or U19912 (N_19912,N_18710,N_18079);
and U19913 (N_19913,N_18581,N_18528);
or U19914 (N_19914,N_18870,N_18193);
nor U19915 (N_19915,N_18674,N_18829);
nand U19916 (N_19916,N_18908,N_18408);
nand U19917 (N_19917,N_18476,N_18270);
nor U19918 (N_19918,N_18753,N_18826);
or U19919 (N_19919,N_18911,N_18216);
and U19920 (N_19920,N_18089,N_18330);
xnor U19921 (N_19921,N_18844,N_18166);
nand U19922 (N_19922,N_18242,N_18889);
and U19923 (N_19923,N_18673,N_18982);
nand U19924 (N_19924,N_18768,N_18848);
xnor U19925 (N_19925,N_18769,N_18878);
and U19926 (N_19926,N_18513,N_18526);
xnor U19927 (N_19927,N_18426,N_18899);
nand U19928 (N_19928,N_18683,N_18480);
and U19929 (N_19929,N_18000,N_18272);
and U19930 (N_19930,N_18825,N_18349);
nor U19931 (N_19931,N_18012,N_18004);
nor U19932 (N_19932,N_18986,N_18226);
nand U19933 (N_19933,N_18575,N_18876);
nor U19934 (N_19934,N_18749,N_18870);
xor U19935 (N_19935,N_18576,N_18264);
nor U19936 (N_19936,N_18737,N_18750);
and U19937 (N_19937,N_18988,N_18652);
xor U19938 (N_19938,N_18478,N_18561);
xor U19939 (N_19939,N_18857,N_18691);
and U19940 (N_19940,N_18677,N_18678);
or U19941 (N_19941,N_18945,N_18184);
nor U19942 (N_19942,N_18339,N_18166);
or U19943 (N_19943,N_18263,N_18420);
nand U19944 (N_19944,N_18883,N_18090);
nor U19945 (N_19945,N_18281,N_18711);
and U19946 (N_19946,N_18038,N_18727);
and U19947 (N_19947,N_18303,N_18245);
nor U19948 (N_19948,N_18217,N_18604);
nor U19949 (N_19949,N_18192,N_18229);
and U19950 (N_19950,N_18681,N_18844);
nand U19951 (N_19951,N_18707,N_18407);
nand U19952 (N_19952,N_18324,N_18934);
nand U19953 (N_19953,N_18148,N_18146);
nor U19954 (N_19954,N_18702,N_18688);
xnor U19955 (N_19955,N_18096,N_18407);
and U19956 (N_19956,N_18546,N_18527);
xnor U19957 (N_19957,N_18925,N_18271);
nand U19958 (N_19958,N_18980,N_18599);
xor U19959 (N_19959,N_18275,N_18484);
nand U19960 (N_19960,N_18017,N_18983);
xnor U19961 (N_19961,N_18306,N_18454);
nand U19962 (N_19962,N_18243,N_18422);
and U19963 (N_19963,N_18926,N_18997);
and U19964 (N_19964,N_18246,N_18081);
or U19965 (N_19965,N_18163,N_18782);
nor U19966 (N_19966,N_18185,N_18716);
nor U19967 (N_19967,N_18124,N_18100);
nand U19968 (N_19968,N_18950,N_18501);
nor U19969 (N_19969,N_18416,N_18102);
or U19970 (N_19970,N_18927,N_18505);
or U19971 (N_19971,N_18910,N_18983);
nand U19972 (N_19972,N_18802,N_18780);
or U19973 (N_19973,N_18481,N_18518);
xnor U19974 (N_19974,N_18726,N_18970);
xnor U19975 (N_19975,N_18100,N_18305);
nand U19976 (N_19976,N_18752,N_18723);
nor U19977 (N_19977,N_18024,N_18663);
or U19978 (N_19978,N_18090,N_18361);
nand U19979 (N_19979,N_18005,N_18761);
xor U19980 (N_19980,N_18379,N_18162);
or U19981 (N_19981,N_18045,N_18222);
nor U19982 (N_19982,N_18079,N_18381);
xor U19983 (N_19983,N_18941,N_18289);
and U19984 (N_19984,N_18902,N_18439);
or U19985 (N_19985,N_18834,N_18500);
xnor U19986 (N_19986,N_18093,N_18144);
xnor U19987 (N_19987,N_18812,N_18029);
nand U19988 (N_19988,N_18088,N_18316);
and U19989 (N_19989,N_18104,N_18707);
nor U19990 (N_19990,N_18427,N_18011);
xnor U19991 (N_19991,N_18523,N_18294);
nand U19992 (N_19992,N_18341,N_18183);
xnor U19993 (N_19993,N_18808,N_18148);
or U19994 (N_19994,N_18275,N_18661);
xnor U19995 (N_19995,N_18508,N_18375);
or U19996 (N_19996,N_18986,N_18807);
xnor U19997 (N_19997,N_18997,N_18766);
nor U19998 (N_19998,N_18195,N_18176);
or U19999 (N_19999,N_18016,N_18142);
and U20000 (N_20000,N_19906,N_19865);
nand U20001 (N_20001,N_19282,N_19530);
and U20002 (N_20002,N_19043,N_19246);
or U20003 (N_20003,N_19391,N_19356);
and U20004 (N_20004,N_19872,N_19135);
nand U20005 (N_20005,N_19484,N_19066);
xor U20006 (N_20006,N_19065,N_19307);
nor U20007 (N_20007,N_19201,N_19141);
nor U20008 (N_20008,N_19581,N_19310);
and U20009 (N_20009,N_19113,N_19738);
or U20010 (N_20010,N_19035,N_19231);
and U20011 (N_20011,N_19704,N_19215);
nor U20012 (N_20012,N_19680,N_19277);
xor U20013 (N_20013,N_19434,N_19538);
nor U20014 (N_20014,N_19705,N_19811);
or U20015 (N_20015,N_19303,N_19427);
or U20016 (N_20016,N_19436,N_19009);
and U20017 (N_20017,N_19404,N_19984);
or U20018 (N_20018,N_19195,N_19922);
nand U20019 (N_20019,N_19742,N_19622);
nor U20020 (N_20020,N_19809,N_19908);
nand U20021 (N_20021,N_19639,N_19881);
and U20022 (N_20022,N_19503,N_19118);
and U20023 (N_20023,N_19154,N_19358);
nor U20024 (N_20024,N_19591,N_19561);
or U20025 (N_20025,N_19890,N_19763);
or U20026 (N_20026,N_19407,N_19312);
or U20027 (N_20027,N_19776,N_19977);
nor U20028 (N_20028,N_19229,N_19518);
and U20029 (N_20029,N_19543,N_19996);
nand U20030 (N_20030,N_19083,N_19399);
and U20031 (N_20031,N_19167,N_19220);
nor U20032 (N_20032,N_19950,N_19219);
nor U20033 (N_20033,N_19058,N_19825);
nand U20034 (N_20034,N_19779,N_19678);
nor U20035 (N_20035,N_19819,N_19621);
and U20036 (N_20036,N_19535,N_19665);
and U20037 (N_20037,N_19021,N_19435);
or U20038 (N_20038,N_19304,N_19433);
nor U20039 (N_20039,N_19945,N_19280);
nor U20040 (N_20040,N_19800,N_19894);
nand U20041 (N_20041,N_19869,N_19656);
or U20042 (N_20042,N_19545,N_19744);
xor U20043 (N_20043,N_19699,N_19153);
xnor U20044 (N_20044,N_19971,N_19626);
nor U20045 (N_20045,N_19091,N_19550);
or U20046 (N_20046,N_19239,N_19953);
xnor U20047 (N_20047,N_19175,N_19264);
xnor U20048 (N_20048,N_19589,N_19863);
or U20049 (N_20049,N_19149,N_19462);
xor U20050 (N_20050,N_19921,N_19162);
nor U20051 (N_20051,N_19641,N_19857);
or U20052 (N_20052,N_19947,N_19269);
xnor U20053 (N_20053,N_19780,N_19853);
and U20054 (N_20054,N_19278,N_19488);
or U20055 (N_20055,N_19722,N_19520);
and U20056 (N_20056,N_19592,N_19198);
and U20057 (N_20057,N_19797,N_19406);
or U20058 (N_20058,N_19480,N_19748);
xor U20059 (N_20059,N_19601,N_19521);
nand U20060 (N_20060,N_19445,N_19335);
nor U20061 (N_20061,N_19205,N_19466);
xnor U20062 (N_20062,N_19218,N_19353);
nor U20063 (N_20063,N_19918,N_19425);
and U20064 (N_20064,N_19424,N_19207);
xnor U20065 (N_20065,N_19046,N_19346);
nor U20066 (N_20066,N_19327,N_19268);
xor U20067 (N_20067,N_19534,N_19919);
and U20068 (N_20068,N_19454,N_19831);
or U20069 (N_20069,N_19410,N_19861);
or U20070 (N_20070,N_19827,N_19372);
and U20071 (N_20071,N_19826,N_19573);
nor U20072 (N_20072,N_19528,N_19572);
and U20073 (N_20073,N_19288,N_19844);
or U20074 (N_20074,N_19851,N_19845);
xor U20075 (N_20075,N_19233,N_19176);
and U20076 (N_20076,N_19806,N_19962);
and U20077 (N_20077,N_19097,N_19004);
nand U20078 (N_20078,N_19839,N_19693);
nor U20079 (N_20079,N_19597,N_19690);
nand U20080 (N_20080,N_19557,N_19171);
and U20081 (N_20081,N_19392,N_19276);
and U20082 (N_20082,N_19813,N_19102);
nor U20083 (N_20083,N_19414,N_19739);
or U20084 (N_20084,N_19613,N_19368);
nand U20085 (N_20085,N_19757,N_19464);
and U20086 (N_20086,N_19493,N_19023);
nor U20087 (N_20087,N_19026,N_19605);
or U20088 (N_20088,N_19075,N_19234);
or U20089 (N_20089,N_19864,N_19305);
or U20090 (N_20090,N_19495,N_19266);
nand U20091 (N_20091,N_19405,N_19850);
nor U20092 (N_20092,N_19903,N_19973);
nor U20093 (N_20093,N_19609,N_19554);
nand U20094 (N_20094,N_19037,N_19259);
nand U20095 (N_20095,N_19700,N_19032);
nor U20096 (N_20096,N_19147,N_19519);
and U20097 (N_20097,N_19822,N_19526);
nor U20098 (N_20098,N_19416,N_19284);
xnor U20099 (N_20099,N_19096,N_19796);
nand U20100 (N_20100,N_19909,N_19238);
nand U20101 (N_20101,N_19753,N_19044);
and U20102 (N_20102,N_19453,N_19868);
or U20103 (N_20103,N_19442,N_19847);
and U20104 (N_20104,N_19062,N_19482);
nand U20105 (N_20105,N_19345,N_19884);
nor U20106 (N_20106,N_19401,N_19784);
and U20107 (N_20107,N_19669,N_19481);
and U20108 (N_20108,N_19529,N_19749);
or U20109 (N_20109,N_19511,N_19571);
xnor U20110 (N_20110,N_19450,N_19910);
or U20111 (N_20111,N_19247,N_19701);
or U20112 (N_20112,N_19017,N_19734);
nand U20113 (N_20113,N_19262,N_19712);
nand U20114 (N_20114,N_19575,N_19691);
and U20115 (N_20115,N_19173,N_19200);
nand U20116 (N_20116,N_19360,N_19491);
or U20117 (N_20117,N_19747,N_19988);
or U20118 (N_20118,N_19446,N_19761);
nand U20119 (N_20119,N_19951,N_19841);
xor U20120 (N_20120,N_19272,N_19965);
nor U20121 (N_20121,N_19187,N_19930);
and U20122 (N_20122,N_19460,N_19192);
nand U20123 (N_20123,N_19208,N_19283);
nand U20124 (N_20124,N_19513,N_19093);
nand U20125 (N_20125,N_19676,N_19620);
nor U20126 (N_20126,N_19323,N_19582);
nand U20127 (N_20127,N_19039,N_19981);
or U20128 (N_20128,N_19408,N_19946);
and U20129 (N_20129,N_19580,N_19386);
or U20130 (N_20130,N_19934,N_19459);
nand U20131 (N_20131,N_19928,N_19477);
or U20132 (N_20132,N_19158,N_19273);
nand U20133 (N_20133,N_19899,N_19190);
nor U20134 (N_20134,N_19512,N_19687);
or U20135 (N_20135,N_19880,N_19221);
nor U20136 (N_20136,N_19652,N_19810);
or U20137 (N_20137,N_19756,N_19030);
xnor U20138 (N_20138,N_19898,N_19183);
or U20139 (N_20139,N_19798,N_19937);
xor U20140 (N_20140,N_19476,N_19764);
xor U20141 (N_20141,N_19456,N_19465);
and U20142 (N_20142,N_19126,N_19213);
nand U20143 (N_20143,N_19105,N_19063);
and U20144 (N_20144,N_19235,N_19382);
or U20145 (N_20145,N_19119,N_19718);
xnor U20146 (N_20146,N_19578,N_19396);
and U20147 (N_20147,N_19522,N_19311);
or U20148 (N_20148,N_19536,N_19726);
xnor U20149 (N_20149,N_19210,N_19555);
or U20150 (N_20150,N_19943,N_19567);
and U20151 (N_20151,N_19352,N_19077);
or U20152 (N_20152,N_19684,N_19479);
nor U20153 (N_20153,N_19619,N_19330);
nand U20154 (N_20154,N_19289,N_19343);
or U20155 (N_20155,N_19308,N_19695);
or U20156 (N_20156,N_19650,N_19878);
nand U20157 (N_20157,N_19677,N_19562);
and U20158 (N_20158,N_19944,N_19969);
xnor U20159 (N_20159,N_19324,N_19270);
xnor U20160 (N_20160,N_19053,N_19031);
nand U20161 (N_20161,N_19257,N_19920);
nand U20162 (N_20162,N_19714,N_19008);
nor U20163 (N_20163,N_19789,N_19122);
xnor U20164 (N_20164,N_19166,N_19729);
xnor U20165 (N_20165,N_19750,N_19799);
nor U20166 (N_20166,N_19760,N_19549);
or U20167 (N_20167,N_19332,N_19936);
nand U20168 (N_20168,N_19683,N_19361);
or U20169 (N_20169,N_19426,N_19240);
xnor U20170 (N_20170,N_19820,N_19960);
and U20171 (N_20171,N_19751,N_19155);
nand U20172 (N_20172,N_19294,N_19672);
xor U20173 (N_20173,N_19527,N_19012);
nor U20174 (N_20174,N_19092,N_19873);
and U20175 (N_20175,N_19261,N_19029);
nor U20176 (N_20176,N_19523,N_19904);
nor U20177 (N_20177,N_19879,N_19888);
or U20178 (N_20178,N_19805,N_19431);
or U20179 (N_20179,N_19647,N_19774);
xnor U20180 (N_20180,N_19357,N_19929);
and U20181 (N_20181,N_19314,N_19161);
nor U20182 (N_20182,N_19508,N_19184);
nand U20183 (N_20183,N_19400,N_19979);
or U20184 (N_20184,N_19309,N_19733);
nand U20185 (N_20185,N_19098,N_19646);
xor U20186 (N_20186,N_19616,N_19380);
nand U20187 (N_20187,N_19611,N_19069);
nand U20188 (N_20188,N_19463,N_19139);
nand U20189 (N_20189,N_19721,N_19193);
nor U20190 (N_20190,N_19994,N_19395);
and U20191 (N_20191,N_19279,N_19300);
or U20192 (N_20192,N_19250,N_19338);
and U20193 (N_20193,N_19532,N_19711);
nor U20194 (N_20194,N_19603,N_19584);
and U20195 (N_20195,N_19131,N_19730);
and U20196 (N_20196,N_19001,N_19895);
xor U20197 (N_20197,N_19110,N_19381);
xnor U20198 (N_20198,N_19574,N_19777);
or U20199 (N_20199,N_19668,N_19255);
or U20200 (N_20200,N_19189,N_19507);
or U20201 (N_20201,N_19291,N_19398);
and U20202 (N_20202,N_19152,N_19054);
and U20203 (N_20203,N_19245,N_19350);
and U20204 (N_20204,N_19049,N_19686);
xnor U20205 (N_20205,N_19443,N_19048);
nor U20206 (N_20206,N_19143,N_19287);
nand U20207 (N_20207,N_19871,N_19657);
or U20208 (N_20208,N_19740,N_19814);
nor U20209 (N_20209,N_19963,N_19724);
xnor U20210 (N_20210,N_19074,N_19271);
nor U20211 (N_20211,N_19961,N_19710);
and U20212 (N_20212,N_19203,N_19145);
and U20213 (N_20213,N_19064,N_19995);
nor U20214 (N_20214,N_19662,N_19635);
nor U20215 (N_20215,N_19275,N_19293);
nor U20216 (N_20216,N_19829,N_19290);
or U20217 (N_20217,N_19320,N_19084);
and U20218 (N_20218,N_19397,N_19180);
xnor U20219 (N_20219,N_19886,N_19586);
nor U20220 (N_20220,N_19754,N_19915);
xnor U20221 (N_20221,N_19583,N_19882);
or U20222 (N_20222,N_19412,N_19376);
and U20223 (N_20223,N_19767,N_19254);
nand U20224 (N_20224,N_19373,N_19177);
and U20225 (N_20225,N_19912,N_19328);
nand U20226 (N_20226,N_19661,N_19978);
or U20227 (N_20227,N_19794,N_19674);
and U20228 (N_20228,N_19604,N_19204);
and U20229 (N_20229,N_19018,N_19423);
and U20230 (N_20230,N_19980,N_19025);
or U20231 (N_20231,N_19743,N_19109);
nor U20232 (N_20232,N_19660,N_19877);
and U20233 (N_20233,N_19354,N_19104);
and U20234 (N_20234,N_19552,N_19413);
nor U20235 (N_20235,N_19499,N_19889);
nor U20236 (N_20236,N_19157,N_19134);
and U20237 (N_20237,N_19485,N_19478);
nor U20238 (N_20238,N_19897,N_19014);
nor U20239 (N_20239,N_19607,N_19546);
or U20240 (N_20240,N_19033,N_19659);
or U20241 (N_20241,N_19371,N_19509);
or U20242 (N_20242,N_19461,N_19059);
nand U20243 (N_20243,N_19081,N_19876);
xor U20244 (N_20244,N_19388,N_19997);
xor U20245 (N_20245,N_19050,N_19156);
nand U20246 (N_20246,N_19663,N_19045);
and U20247 (N_20247,N_19627,N_19618);
nor U20248 (N_20248,N_19088,N_19011);
and U20249 (N_20249,N_19801,N_19441);
nand U20250 (N_20250,N_19206,N_19812);
and U20251 (N_20251,N_19212,N_19447);
and U20252 (N_20252,N_19094,N_19498);
xnor U20253 (N_20253,N_19384,N_19067);
nand U20254 (N_20254,N_19265,N_19028);
and U20255 (N_20255,N_19347,N_19887);
nand U20256 (N_20256,N_19020,N_19987);
nor U20257 (N_20257,N_19974,N_19121);
or U20258 (N_20258,N_19792,N_19103);
and U20259 (N_20259,N_19999,N_19417);
xnor U20260 (N_20260,N_19430,N_19344);
xnor U20261 (N_20261,N_19383,N_19612);
and U20262 (N_20262,N_19244,N_19927);
nor U20263 (N_20263,N_19688,N_19468);
nor U20264 (N_20264,N_19931,N_19642);
nor U20265 (N_20265,N_19992,N_19114);
nor U20266 (N_20266,N_19348,N_19164);
or U20267 (N_20267,N_19163,N_19697);
nor U20268 (N_20268,N_19653,N_19467);
nor U20269 (N_20269,N_19875,N_19632);
or U20270 (N_20270,N_19539,N_19892);
nand U20271 (N_20271,N_19140,N_19883);
nand U20272 (N_20272,N_19544,N_19630);
or U20273 (N_20273,N_19727,N_19804);
xor U20274 (N_20274,N_19148,N_19179);
and U20275 (N_20275,N_19939,N_19787);
or U20276 (N_20276,N_19651,N_19692);
nor U20277 (N_20277,N_19194,N_19696);
and U20278 (N_20278,N_19599,N_19896);
xor U20279 (N_20279,N_19551,N_19533);
xnor U20280 (N_20280,N_19086,N_19336);
or U20281 (N_20281,N_19949,N_19076);
or U20282 (N_20282,N_19941,N_19858);
xnor U20283 (N_20283,N_19752,N_19515);
nand U20284 (N_20284,N_19199,N_19321);
nor U20285 (N_20285,N_19333,N_19319);
and U20286 (N_20286,N_19082,N_19640);
nor U20287 (N_20287,N_19051,N_19379);
or U20288 (N_20288,N_19237,N_19267);
and U20289 (N_20289,N_19146,N_19795);
nor U20290 (N_20290,N_19563,N_19745);
nand U20291 (N_20291,N_19566,N_19629);
or U20292 (N_20292,N_19355,N_19577);
nor U20293 (N_20293,N_19003,N_19842);
nor U20294 (N_20294,N_19998,N_19337);
xor U20295 (N_20295,N_19833,N_19124);
nand U20296 (N_20296,N_19986,N_19227);
nand U20297 (N_20297,N_19060,N_19438);
nand U20298 (N_20298,N_19496,N_19341);
and U20299 (N_20299,N_19365,N_19393);
and U20300 (N_20300,N_19057,N_19191);
nor U20301 (N_20301,N_19732,N_19449);
nand U20302 (N_20302,N_19252,N_19602);
nor U20303 (N_20303,N_19223,N_19295);
nand U20304 (N_20304,N_19068,N_19976);
or U20305 (N_20305,N_19517,N_19633);
xnor U20306 (N_20306,N_19715,N_19224);
nor U20307 (N_20307,N_19556,N_19564);
or U20308 (N_20308,N_19185,N_19429);
or U20309 (N_20309,N_19600,N_19168);
nor U20310 (N_20310,N_19785,N_19548);
and U20311 (N_20311,N_19637,N_19838);
and U20312 (N_20312,N_19169,N_19428);
or U20313 (N_20313,N_19793,N_19905);
xnor U20314 (N_20314,N_19643,N_19862);
nor U20315 (N_20315,N_19542,N_19855);
xor U20316 (N_20316,N_19924,N_19115);
nor U20317 (N_20317,N_19367,N_19615);
and U20318 (N_20318,N_19666,N_19492);
xnor U20319 (N_20319,N_19772,N_19728);
and U20320 (N_20320,N_19242,N_19648);
nor U20321 (N_20321,N_19101,N_19547);
and U20322 (N_20322,N_19832,N_19133);
or U20323 (N_20323,N_19385,N_19689);
nand U20324 (N_20324,N_19170,N_19497);
and U20325 (N_20325,N_19759,N_19364);
and U20326 (N_20326,N_19595,N_19174);
nand U20327 (N_20327,N_19013,N_19671);
xor U20328 (N_20328,N_19860,N_19249);
or U20329 (N_20329,N_19420,N_19596);
and U20330 (N_20330,N_19954,N_19933);
or U20331 (N_20331,N_19389,N_19253);
nand U20332 (N_20332,N_19403,N_19849);
or U20333 (N_20333,N_19111,N_19716);
nor U20334 (N_20334,N_19725,N_19501);
nor U20335 (N_20335,N_19955,N_19658);
nor U20336 (N_20336,N_19196,N_19274);
nand U20337 (N_20337,N_19306,N_19486);
and U20338 (N_20338,N_19243,N_19706);
and U20339 (N_20339,N_19072,N_19673);
and U20340 (N_20340,N_19803,N_19409);
nand U20341 (N_20341,N_19993,N_19840);
nand U20342 (N_20342,N_19956,N_19494);
nand U20343 (N_20343,N_19452,N_19823);
nand U20344 (N_20344,N_19052,N_19322);
nor U20345 (N_20345,N_19137,N_19634);
nor U20346 (N_20346,N_19590,N_19870);
nor U20347 (N_20347,N_19448,N_19006);
xnor U20348 (N_20348,N_19808,N_19349);
xnor U20349 (N_20349,N_19316,N_19078);
nand U20350 (N_20350,N_19225,N_19585);
and U20351 (N_20351,N_19975,N_19329);
xnor U20352 (N_20352,N_19339,N_19024);
nand U20353 (N_20353,N_19297,N_19859);
nand U20354 (N_20354,N_19432,N_19655);
and U20355 (N_20355,N_19893,N_19649);
or U20356 (N_20356,N_19325,N_19375);
xor U20357 (N_20357,N_19359,N_19902);
xnor U20358 (N_20358,N_19598,N_19594);
nor U20359 (N_20359,N_19186,N_19606);
nand U20360 (N_20360,N_19151,N_19932);
nand U20361 (N_20361,N_19768,N_19970);
nand U20362 (N_20362,N_19457,N_19834);
and U20363 (N_20363,N_19991,N_19900);
xnor U20364 (N_20364,N_19298,N_19781);
or U20365 (N_20365,N_19854,N_19913);
nand U20366 (N_20366,N_19846,N_19470);
nand U20367 (N_20367,N_19516,N_19016);
or U20368 (N_20368,N_19762,N_19856);
xnor U20369 (N_20369,N_19340,N_19318);
nand U20370 (N_20370,N_19758,N_19818);
nor U20371 (N_20371,N_19369,N_19125);
and U20372 (N_20372,N_19773,N_19681);
nand U20373 (N_20373,N_19036,N_19654);
and U20374 (N_20374,N_19766,N_19989);
or U20375 (N_20375,N_19469,N_19982);
or U20376 (N_20376,N_19807,N_19061);
and U20377 (N_20377,N_19150,N_19326);
xor U20378 (N_20378,N_19130,N_19073);
or U20379 (N_20379,N_19473,N_19458);
nor U20380 (N_20380,N_19685,N_19852);
xor U20381 (N_20381,N_19007,N_19707);
or U20382 (N_20382,N_19116,N_19541);
nor U20383 (N_20383,N_19022,N_19990);
xor U20384 (N_20384,N_19315,N_19444);
nand U20385 (N_20385,N_19940,N_19588);
and U20386 (N_20386,N_19471,N_19958);
nor U20387 (N_20387,N_19019,N_19182);
and U20388 (N_20388,N_19292,N_19002);
nand U20389 (N_20389,N_19117,N_19694);
nor U20390 (N_20390,N_19217,N_19769);
and U20391 (N_20391,N_19967,N_19972);
and U20392 (N_20392,N_19474,N_19165);
nor U20393 (N_20393,N_19682,N_19709);
and U20394 (N_20394,N_19631,N_19313);
xnor U20395 (N_20395,N_19948,N_19874);
nand U20396 (N_20396,N_19506,N_19080);
nor U20397 (N_20397,N_19926,N_19891);
xnor U20398 (N_20398,N_19828,N_19351);
or U20399 (N_20399,N_19765,N_19723);
and U20400 (N_20400,N_19128,N_19702);
xor U20401 (N_20401,N_19000,N_19957);
or U20402 (N_20402,N_19679,N_19746);
nand U20403 (N_20403,N_19815,N_19472);
nor U20404 (N_20404,N_19228,N_19377);
nand U20405 (N_20405,N_19144,N_19487);
nor U20406 (N_20406,N_19079,N_19342);
and U20407 (N_20407,N_19136,N_19568);
nand U20408 (N_20408,N_19959,N_19628);
nand U20409 (N_20409,N_19771,N_19451);
or U20410 (N_20410,N_19241,N_19782);
xnor U20411 (N_20411,N_19363,N_19087);
or U20412 (N_20412,N_19085,N_19214);
or U20413 (N_20413,N_19222,N_19100);
and U20414 (N_20414,N_19731,N_19755);
nor U20415 (N_20415,N_19917,N_19178);
nor U20416 (N_20416,N_19071,N_19636);
nand U20417 (N_20417,N_19402,N_19056);
nor U20418 (N_20418,N_19387,N_19778);
xnor U20419 (N_20419,N_19617,N_19505);
and U20420 (N_20420,N_19034,N_19565);
or U20421 (N_20421,N_19670,N_19202);
xor U20422 (N_20422,N_19188,N_19708);
and U20423 (N_20423,N_19741,N_19537);
and U20424 (N_20424,N_19286,N_19587);
or U20425 (N_20425,N_19835,N_19703);
nor U20426 (N_20426,N_19302,N_19090);
and U20427 (N_20427,N_19964,N_19843);
and U20428 (N_20428,N_19258,N_19041);
or U20429 (N_20429,N_19916,N_19524);
nand U20430 (N_20430,N_19230,N_19579);
or U20431 (N_20431,N_19260,N_19719);
or U20432 (N_20432,N_19817,N_19667);
or U20433 (N_20433,N_19129,N_19500);
nand U20434 (N_20434,N_19558,N_19514);
or U20435 (N_20435,N_19263,N_19938);
nor U20436 (N_20436,N_19394,N_19209);
nand U20437 (N_20437,N_19942,N_19027);
nor U20438 (N_20438,N_19127,N_19421);
nor U20439 (N_20439,N_19783,N_19770);
nand U20440 (N_20440,N_19455,N_19107);
or U20441 (N_20441,N_19923,N_19985);
nand U20442 (N_20442,N_19390,N_19256);
nor U20443 (N_20443,N_19483,N_19138);
nor U20444 (N_20444,N_19285,N_19281);
and U20445 (N_20445,N_19197,N_19251);
or U20446 (N_20446,N_19422,N_19510);
and U20447 (N_20447,N_19362,N_19106);
nor U20448 (N_20448,N_19331,N_19914);
or U20449 (N_20449,N_19120,N_19296);
nand U20450 (N_20450,N_19015,N_19415);
or U20451 (N_20451,N_19816,N_19614);
nor U20452 (N_20452,N_19216,N_19952);
and U20453 (N_20453,N_19983,N_19005);
nand U20454 (N_20454,N_19720,N_19791);
and U20455 (N_20455,N_19042,N_19698);
or U20456 (N_20456,N_19560,N_19236);
or U20457 (N_20457,N_19624,N_19625);
xnor U20458 (N_20458,N_19525,N_19644);
nor U20459 (N_20459,N_19786,N_19374);
and U20460 (N_20460,N_19966,N_19047);
or U20461 (N_20461,N_19038,N_19502);
nor U20462 (N_20462,N_19735,N_19248);
and U20463 (N_20463,N_19569,N_19717);
xor U20464 (N_20464,N_19301,N_19490);
and U20465 (N_20465,N_19867,N_19317);
nand U20466 (N_20466,N_19675,N_19010);
or U20467 (N_20467,N_19848,N_19925);
nor U20468 (N_20468,N_19089,N_19713);
or U20469 (N_20469,N_19645,N_19070);
and U20470 (N_20470,N_19638,N_19437);
or U20471 (N_20471,N_19559,N_19211);
or U20472 (N_20472,N_19378,N_19531);
xor U20473 (N_20473,N_19099,N_19370);
nor U20474 (N_20474,N_19334,N_19837);
nand U20475 (N_20475,N_19593,N_19775);
nor U20476 (N_20476,N_19830,N_19181);
nor U20477 (N_20477,N_19159,N_19576);
nand U20478 (N_20478,N_19299,N_19132);
and U20479 (N_20479,N_19440,N_19112);
xnor U20480 (N_20480,N_19911,N_19736);
nor U20481 (N_20481,N_19836,N_19142);
xnor U20482 (N_20482,N_19737,N_19411);
xor U20483 (N_20483,N_19824,N_19821);
nor U20484 (N_20484,N_19540,N_19623);
or U20485 (N_20485,N_19172,N_19968);
nor U20486 (N_20486,N_19108,N_19504);
nor U20487 (N_20487,N_19553,N_19885);
nor U20488 (N_20488,N_19907,N_19040);
or U20489 (N_20489,N_19788,N_19160);
nor U20490 (N_20490,N_19935,N_19610);
nand U20491 (N_20491,N_19608,N_19055);
xor U20492 (N_20492,N_19790,N_19419);
nand U20493 (N_20493,N_19366,N_19802);
nor U20494 (N_20494,N_19489,N_19866);
and U20495 (N_20495,N_19475,N_19418);
xnor U20496 (N_20496,N_19226,N_19570);
nor U20497 (N_20497,N_19232,N_19095);
or U20498 (N_20498,N_19439,N_19123);
or U20499 (N_20499,N_19901,N_19664);
xor U20500 (N_20500,N_19858,N_19863);
or U20501 (N_20501,N_19787,N_19862);
nor U20502 (N_20502,N_19918,N_19491);
nand U20503 (N_20503,N_19419,N_19355);
nand U20504 (N_20504,N_19954,N_19634);
nor U20505 (N_20505,N_19615,N_19510);
nand U20506 (N_20506,N_19423,N_19389);
or U20507 (N_20507,N_19286,N_19691);
xor U20508 (N_20508,N_19973,N_19333);
nand U20509 (N_20509,N_19251,N_19990);
nand U20510 (N_20510,N_19781,N_19297);
nor U20511 (N_20511,N_19240,N_19119);
nand U20512 (N_20512,N_19035,N_19629);
nand U20513 (N_20513,N_19860,N_19980);
xnor U20514 (N_20514,N_19643,N_19359);
or U20515 (N_20515,N_19655,N_19881);
xor U20516 (N_20516,N_19050,N_19011);
and U20517 (N_20517,N_19001,N_19957);
and U20518 (N_20518,N_19039,N_19375);
nor U20519 (N_20519,N_19530,N_19129);
xor U20520 (N_20520,N_19426,N_19845);
nor U20521 (N_20521,N_19637,N_19599);
xnor U20522 (N_20522,N_19860,N_19332);
and U20523 (N_20523,N_19598,N_19637);
nor U20524 (N_20524,N_19224,N_19166);
xnor U20525 (N_20525,N_19048,N_19870);
xor U20526 (N_20526,N_19537,N_19730);
xnor U20527 (N_20527,N_19934,N_19467);
and U20528 (N_20528,N_19582,N_19781);
xor U20529 (N_20529,N_19896,N_19457);
nand U20530 (N_20530,N_19203,N_19033);
xnor U20531 (N_20531,N_19801,N_19141);
nor U20532 (N_20532,N_19482,N_19280);
xnor U20533 (N_20533,N_19885,N_19131);
and U20534 (N_20534,N_19329,N_19706);
nor U20535 (N_20535,N_19526,N_19899);
xor U20536 (N_20536,N_19472,N_19731);
and U20537 (N_20537,N_19630,N_19579);
or U20538 (N_20538,N_19032,N_19957);
nand U20539 (N_20539,N_19892,N_19096);
or U20540 (N_20540,N_19377,N_19381);
and U20541 (N_20541,N_19771,N_19521);
xor U20542 (N_20542,N_19025,N_19300);
xor U20543 (N_20543,N_19932,N_19238);
nor U20544 (N_20544,N_19411,N_19072);
and U20545 (N_20545,N_19104,N_19934);
xnor U20546 (N_20546,N_19222,N_19741);
or U20547 (N_20547,N_19406,N_19248);
nand U20548 (N_20548,N_19696,N_19577);
nor U20549 (N_20549,N_19265,N_19536);
and U20550 (N_20550,N_19854,N_19384);
xor U20551 (N_20551,N_19474,N_19156);
or U20552 (N_20552,N_19296,N_19285);
nor U20553 (N_20553,N_19467,N_19366);
xor U20554 (N_20554,N_19528,N_19922);
nand U20555 (N_20555,N_19414,N_19601);
or U20556 (N_20556,N_19159,N_19329);
and U20557 (N_20557,N_19879,N_19329);
and U20558 (N_20558,N_19583,N_19217);
or U20559 (N_20559,N_19812,N_19511);
or U20560 (N_20560,N_19410,N_19560);
and U20561 (N_20561,N_19402,N_19681);
xnor U20562 (N_20562,N_19895,N_19679);
xor U20563 (N_20563,N_19548,N_19799);
or U20564 (N_20564,N_19930,N_19026);
nand U20565 (N_20565,N_19579,N_19756);
nor U20566 (N_20566,N_19470,N_19353);
or U20567 (N_20567,N_19920,N_19250);
nor U20568 (N_20568,N_19238,N_19302);
or U20569 (N_20569,N_19452,N_19953);
nor U20570 (N_20570,N_19171,N_19505);
and U20571 (N_20571,N_19094,N_19646);
nand U20572 (N_20572,N_19115,N_19821);
nand U20573 (N_20573,N_19367,N_19420);
and U20574 (N_20574,N_19328,N_19955);
xor U20575 (N_20575,N_19773,N_19700);
and U20576 (N_20576,N_19362,N_19076);
xnor U20577 (N_20577,N_19540,N_19886);
nand U20578 (N_20578,N_19565,N_19428);
nand U20579 (N_20579,N_19086,N_19433);
nor U20580 (N_20580,N_19449,N_19935);
nand U20581 (N_20581,N_19078,N_19292);
nand U20582 (N_20582,N_19979,N_19309);
nor U20583 (N_20583,N_19699,N_19227);
nor U20584 (N_20584,N_19066,N_19752);
and U20585 (N_20585,N_19955,N_19323);
nor U20586 (N_20586,N_19055,N_19227);
and U20587 (N_20587,N_19760,N_19636);
nor U20588 (N_20588,N_19501,N_19408);
nand U20589 (N_20589,N_19125,N_19212);
nor U20590 (N_20590,N_19237,N_19280);
xnor U20591 (N_20591,N_19344,N_19461);
xor U20592 (N_20592,N_19681,N_19107);
nand U20593 (N_20593,N_19306,N_19271);
nand U20594 (N_20594,N_19913,N_19874);
xnor U20595 (N_20595,N_19233,N_19000);
nand U20596 (N_20596,N_19649,N_19785);
nor U20597 (N_20597,N_19288,N_19547);
and U20598 (N_20598,N_19138,N_19615);
nor U20599 (N_20599,N_19857,N_19853);
and U20600 (N_20600,N_19430,N_19597);
nand U20601 (N_20601,N_19060,N_19433);
and U20602 (N_20602,N_19131,N_19726);
or U20603 (N_20603,N_19602,N_19982);
xor U20604 (N_20604,N_19770,N_19275);
and U20605 (N_20605,N_19405,N_19968);
nor U20606 (N_20606,N_19581,N_19287);
nand U20607 (N_20607,N_19549,N_19260);
nand U20608 (N_20608,N_19201,N_19910);
xnor U20609 (N_20609,N_19066,N_19386);
nor U20610 (N_20610,N_19649,N_19501);
nand U20611 (N_20611,N_19347,N_19882);
nand U20612 (N_20612,N_19919,N_19432);
nor U20613 (N_20613,N_19945,N_19938);
or U20614 (N_20614,N_19115,N_19414);
xor U20615 (N_20615,N_19962,N_19440);
nand U20616 (N_20616,N_19649,N_19913);
nor U20617 (N_20617,N_19693,N_19589);
and U20618 (N_20618,N_19261,N_19553);
and U20619 (N_20619,N_19650,N_19902);
nor U20620 (N_20620,N_19500,N_19171);
and U20621 (N_20621,N_19230,N_19380);
nor U20622 (N_20622,N_19814,N_19775);
nor U20623 (N_20623,N_19117,N_19492);
or U20624 (N_20624,N_19948,N_19439);
nor U20625 (N_20625,N_19938,N_19488);
or U20626 (N_20626,N_19177,N_19215);
xor U20627 (N_20627,N_19706,N_19893);
nor U20628 (N_20628,N_19484,N_19140);
nand U20629 (N_20629,N_19385,N_19803);
or U20630 (N_20630,N_19573,N_19128);
xnor U20631 (N_20631,N_19433,N_19674);
nor U20632 (N_20632,N_19888,N_19748);
nand U20633 (N_20633,N_19001,N_19023);
nor U20634 (N_20634,N_19971,N_19037);
nor U20635 (N_20635,N_19951,N_19344);
and U20636 (N_20636,N_19866,N_19878);
xnor U20637 (N_20637,N_19385,N_19663);
and U20638 (N_20638,N_19683,N_19723);
nand U20639 (N_20639,N_19177,N_19788);
nor U20640 (N_20640,N_19656,N_19768);
xnor U20641 (N_20641,N_19994,N_19300);
nor U20642 (N_20642,N_19788,N_19825);
nand U20643 (N_20643,N_19423,N_19865);
xnor U20644 (N_20644,N_19016,N_19411);
or U20645 (N_20645,N_19155,N_19941);
and U20646 (N_20646,N_19100,N_19677);
and U20647 (N_20647,N_19152,N_19580);
nand U20648 (N_20648,N_19611,N_19441);
or U20649 (N_20649,N_19359,N_19313);
and U20650 (N_20650,N_19604,N_19971);
nand U20651 (N_20651,N_19910,N_19672);
or U20652 (N_20652,N_19645,N_19591);
xnor U20653 (N_20653,N_19725,N_19635);
or U20654 (N_20654,N_19437,N_19355);
and U20655 (N_20655,N_19323,N_19992);
or U20656 (N_20656,N_19473,N_19475);
nand U20657 (N_20657,N_19071,N_19005);
nor U20658 (N_20658,N_19044,N_19740);
or U20659 (N_20659,N_19299,N_19660);
xnor U20660 (N_20660,N_19724,N_19048);
and U20661 (N_20661,N_19748,N_19695);
xnor U20662 (N_20662,N_19598,N_19347);
or U20663 (N_20663,N_19309,N_19661);
and U20664 (N_20664,N_19946,N_19414);
and U20665 (N_20665,N_19643,N_19410);
nor U20666 (N_20666,N_19456,N_19518);
nor U20667 (N_20667,N_19502,N_19332);
xor U20668 (N_20668,N_19499,N_19756);
and U20669 (N_20669,N_19860,N_19247);
and U20670 (N_20670,N_19072,N_19611);
nor U20671 (N_20671,N_19765,N_19945);
nand U20672 (N_20672,N_19002,N_19782);
nor U20673 (N_20673,N_19689,N_19220);
and U20674 (N_20674,N_19873,N_19790);
and U20675 (N_20675,N_19645,N_19370);
nand U20676 (N_20676,N_19272,N_19990);
or U20677 (N_20677,N_19991,N_19764);
nor U20678 (N_20678,N_19055,N_19694);
and U20679 (N_20679,N_19000,N_19075);
nor U20680 (N_20680,N_19301,N_19195);
xnor U20681 (N_20681,N_19594,N_19041);
or U20682 (N_20682,N_19161,N_19083);
nand U20683 (N_20683,N_19174,N_19296);
nor U20684 (N_20684,N_19705,N_19703);
and U20685 (N_20685,N_19914,N_19366);
or U20686 (N_20686,N_19720,N_19251);
xnor U20687 (N_20687,N_19302,N_19461);
nand U20688 (N_20688,N_19398,N_19046);
or U20689 (N_20689,N_19346,N_19188);
and U20690 (N_20690,N_19315,N_19636);
and U20691 (N_20691,N_19719,N_19969);
nor U20692 (N_20692,N_19598,N_19491);
xnor U20693 (N_20693,N_19239,N_19183);
and U20694 (N_20694,N_19843,N_19555);
and U20695 (N_20695,N_19965,N_19389);
or U20696 (N_20696,N_19511,N_19397);
nor U20697 (N_20697,N_19063,N_19422);
or U20698 (N_20698,N_19223,N_19428);
xor U20699 (N_20699,N_19282,N_19031);
or U20700 (N_20700,N_19963,N_19966);
nand U20701 (N_20701,N_19605,N_19840);
and U20702 (N_20702,N_19258,N_19119);
nor U20703 (N_20703,N_19735,N_19294);
nand U20704 (N_20704,N_19762,N_19646);
nor U20705 (N_20705,N_19798,N_19975);
and U20706 (N_20706,N_19849,N_19963);
nor U20707 (N_20707,N_19493,N_19120);
or U20708 (N_20708,N_19202,N_19083);
xnor U20709 (N_20709,N_19131,N_19810);
or U20710 (N_20710,N_19001,N_19930);
or U20711 (N_20711,N_19651,N_19299);
xnor U20712 (N_20712,N_19597,N_19936);
and U20713 (N_20713,N_19982,N_19517);
or U20714 (N_20714,N_19004,N_19770);
and U20715 (N_20715,N_19012,N_19482);
or U20716 (N_20716,N_19603,N_19263);
xnor U20717 (N_20717,N_19817,N_19039);
nand U20718 (N_20718,N_19721,N_19219);
xor U20719 (N_20719,N_19173,N_19325);
and U20720 (N_20720,N_19493,N_19944);
or U20721 (N_20721,N_19509,N_19682);
xor U20722 (N_20722,N_19609,N_19689);
nor U20723 (N_20723,N_19227,N_19279);
xor U20724 (N_20724,N_19642,N_19772);
and U20725 (N_20725,N_19959,N_19658);
nor U20726 (N_20726,N_19443,N_19211);
nor U20727 (N_20727,N_19437,N_19446);
nor U20728 (N_20728,N_19211,N_19174);
and U20729 (N_20729,N_19283,N_19108);
nand U20730 (N_20730,N_19486,N_19344);
nor U20731 (N_20731,N_19677,N_19245);
xnor U20732 (N_20732,N_19014,N_19895);
nand U20733 (N_20733,N_19545,N_19390);
and U20734 (N_20734,N_19840,N_19220);
xor U20735 (N_20735,N_19641,N_19736);
or U20736 (N_20736,N_19842,N_19443);
nor U20737 (N_20737,N_19149,N_19591);
or U20738 (N_20738,N_19620,N_19362);
nand U20739 (N_20739,N_19524,N_19213);
nor U20740 (N_20740,N_19425,N_19197);
xnor U20741 (N_20741,N_19915,N_19363);
and U20742 (N_20742,N_19738,N_19220);
or U20743 (N_20743,N_19505,N_19813);
and U20744 (N_20744,N_19478,N_19492);
nor U20745 (N_20745,N_19469,N_19894);
nor U20746 (N_20746,N_19993,N_19881);
xor U20747 (N_20747,N_19824,N_19271);
nand U20748 (N_20748,N_19903,N_19353);
nand U20749 (N_20749,N_19878,N_19142);
nand U20750 (N_20750,N_19778,N_19455);
and U20751 (N_20751,N_19266,N_19199);
xor U20752 (N_20752,N_19362,N_19118);
xor U20753 (N_20753,N_19937,N_19894);
or U20754 (N_20754,N_19095,N_19384);
nand U20755 (N_20755,N_19796,N_19966);
xnor U20756 (N_20756,N_19261,N_19789);
xnor U20757 (N_20757,N_19390,N_19992);
and U20758 (N_20758,N_19311,N_19744);
xor U20759 (N_20759,N_19535,N_19541);
nor U20760 (N_20760,N_19140,N_19071);
xor U20761 (N_20761,N_19102,N_19782);
or U20762 (N_20762,N_19905,N_19960);
xnor U20763 (N_20763,N_19591,N_19255);
nand U20764 (N_20764,N_19841,N_19729);
and U20765 (N_20765,N_19371,N_19802);
xnor U20766 (N_20766,N_19869,N_19453);
nor U20767 (N_20767,N_19926,N_19537);
nand U20768 (N_20768,N_19922,N_19483);
xor U20769 (N_20769,N_19359,N_19050);
nor U20770 (N_20770,N_19218,N_19442);
xnor U20771 (N_20771,N_19483,N_19531);
or U20772 (N_20772,N_19525,N_19940);
and U20773 (N_20773,N_19014,N_19369);
nand U20774 (N_20774,N_19508,N_19379);
and U20775 (N_20775,N_19153,N_19546);
nor U20776 (N_20776,N_19053,N_19631);
or U20777 (N_20777,N_19215,N_19790);
nand U20778 (N_20778,N_19408,N_19230);
and U20779 (N_20779,N_19421,N_19380);
nor U20780 (N_20780,N_19931,N_19961);
or U20781 (N_20781,N_19303,N_19138);
and U20782 (N_20782,N_19730,N_19660);
nor U20783 (N_20783,N_19807,N_19991);
nand U20784 (N_20784,N_19153,N_19128);
xor U20785 (N_20785,N_19491,N_19172);
nor U20786 (N_20786,N_19114,N_19306);
nor U20787 (N_20787,N_19993,N_19096);
xor U20788 (N_20788,N_19958,N_19577);
nand U20789 (N_20789,N_19217,N_19552);
or U20790 (N_20790,N_19948,N_19613);
nand U20791 (N_20791,N_19671,N_19977);
nand U20792 (N_20792,N_19423,N_19477);
xor U20793 (N_20793,N_19668,N_19314);
xor U20794 (N_20794,N_19170,N_19723);
and U20795 (N_20795,N_19540,N_19897);
nor U20796 (N_20796,N_19409,N_19298);
or U20797 (N_20797,N_19617,N_19124);
or U20798 (N_20798,N_19360,N_19359);
nand U20799 (N_20799,N_19201,N_19447);
and U20800 (N_20800,N_19906,N_19568);
xnor U20801 (N_20801,N_19217,N_19655);
and U20802 (N_20802,N_19955,N_19461);
and U20803 (N_20803,N_19003,N_19930);
and U20804 (N_20804,N_19488,N_19942);
or U20805 (N_20805,N_19170,N_19218);
or U20806 (N_20806,N_19250,N_19117);
nor U20807 (N_20807,N_19601,N_19441);
nand U20808 (N_20808,N_19752,N_19084);
xnor U20809 (N_20809,N_19061,N_19128);
xnor U20810 (N_20810,N_19011,N_19345);
nor U20811 (N_20811,N_19689,N_19087);
and U20812 (N_20812,N_19255,N_19004);
and U20813 (N_20813,N_19532,N_19151);
nand U20814 (N_20814,N_19346,N_19246);
and U20815 (N_20815,N_19234,N_19444);
nand U20816 (N_20816,N_19229,N_19228);
or U20817 (N_20817,N_19305,N_19339);
xnor U20818 (N_20818,N_19188,N_19621);
nor U20819 (N_20819,N_19038,N_19590);
nand U20820 (N_20820,N_19412,N_19599);
xnor U20821 (N_20821,N_19973,N_19984);
xor U20822 (N_20822,N_19431,N_19038);
nor U20823 (N_20823,N_19372,N_19574);
nor U20824 (N_20824,N_19358,N_19809);
and U20825 (N_20825,N_19247,N_19012);
xnor U20826 (N_20826,N_19233,N_19619);
nand U20827 (N_20827,N_19735,N_19884);
xnor U20828 (N_20828,N_19970,N_19622);
and U20829 (N_20829,N_19267,N_19812);
nand U20830 (N_20830,N_19844,N_19388);
nor U20831 (N_20831,N_19100,N_19631);
nor U20832 (N_20832,N_19273,N_19614);
xor U20833 (N_20833,N_19818,N_19587);
xor U20834 (N_20834,N_19488,N_19307);
xnor U20835 (N_20835,N_19181,N_19735);
and U20836 (N_20836,N_19712,N_19177);
nand U20837 (N_20837,N_19654,N_19843);
and U20838 (N_20838,N_19067,N_19219);
and U20839 (N_20839,N_19140,N_19450);
or U20840 (N_20840,N_19730,N_19293);
xnor U20841 (N_20841,N_19455,N_19893);
nand U20842 (N_20842,N_19214,N_19847);
nor U20843 (N_20843,N_19899,N_19053);
nor U20844 (N_20844,N_19812,N_19516);
nor U20845 (N_20845,N_19064,N_19825);
nand U20846 (N_20846,N_19628,N_19853);
xnor U20847 (N_20847,N_19790,N_19366);
or U20848 (N_20848,N_19642,N_19877);
or U20849 (N_20849,N_19870,N_19730);
xnor U20850 (N_20850,N_19082,N_19217);
nor U20851 (N_20851,N_19047,N_19289);
xnor U20852 (N_20852,N_19929,N_19530);
nor U20853 (N_20853,N_19307,N_19755);
nor U20854 (N_20854,N_19620,N_19280);
or U20855 (N_20855,N_19124,N_19140);
nand U20856 (N_20856,N_19184,N_19463);
nand U20857 (N_20857,N_19202,N_19421);
or U20858 (N_20858,N_19557,N_19524);
xor U20859 (N_20859,N_19634,N_19978);
and U20860 (N_20860,N_19376,N_19393);
nor U20861 (N_20861,N_19852,N_19407);
or U20862 (N_20862,N_19725,N_19375);
and U20863 (N_20863,N_19881,N_19415);
nand U20864 (N_20864,N_19188,N_19160);
xor U20865 (N_20865,N_19142,N_19016);
xnor U20866 (N_20866,N_19415,N_19061);
xor U20867 (N_20867,N_19788,N_19197);
nor U20868 (N_20868,N_19147,N_19467);
xor U20869 (N_20869,N_19373,N_19868);
nand U20870 (N_20870,N_19439,N_19452);
or U20871 (N_20871,N_19233,N_19381);
or U20872 (N_20872,N_19086,N_19256);
and U20873 (N_20873,N_19895,N_19043);
or U20874 (N_20874,N_19123,N_19374);
nor U20875 (N_20875,N_19158,N_19341);
or U20876 (N_20876,N_19154,N_19962);
nor U20877 (N_20877,N_19341,N_19525);
xor U20878 (N_20878,N_19965,N_19406);
xnor U20879 (N_20879,N_19097,N_19841);
and U20880 (N_20880,N_19148,N_19201);
xnor U20881 (N_20881,N_19648,N_19512);
nand U20882 (N_20882,N_19681,N_19645);
xnor U20883 (N_20883,N_19035,N_19738);
nand U20884 (N_20884,N_19316,N_19229);
and U20885 (N_20885,N_19096,N_19889);
or U20886 (N_20886,N_19100,N_19730);
nor U20887 (N_20887,N_19039,N_19077);
xnor U20888 (N_20888,N_19144,N_19424);
nor U20889 (N_20889,N_19215,N_19614);
and U20890 (N_20890,N_19339,N_19522);
or U20891 (N_20891,N_19867,N_19108);
nor U20892 (N_20892,N_19349,N_19451);
nor U20893 (N_20893,N_19012,N_19996);
xor U20894 (N_20894,N_19952,N_19392);
and U20895 (N_20895,N_19158,N_19128);
and U20896 (N_20896,N_19543,N_19085);
nor U20897 (N_20897,N_19895,N_19734);
or U20898 (N_20898,N_19465,N_19847);
and U20899 (N_20899,N_19500,N_19874);
and U20900 (N_20900,N_19789,N_19290);
xor U20901 (N_20901,N_19309,N_19706);
nand U20902 (N_20902,N_19591,N_19114);
nor U20903 (N_20903,N_19121,N_19029);
xnor U20904 (N_20904,N_19548,N_19173);
nand U20905 (N_20905,N_19874,N_19460);
and U20906 (N_20906,N_19460,N_19392);
nand U20907 (N_20907,N_19782,N_19354);
nor U20908 (N_20908,N_19941,N_19029);
or U20909 (N_20909,N_19481,N_19393);
and U20910 (N_20910,N_19637,N_19158);
and U20911 (N_20911,N_19074,N_19031);
nand U20912 (N_20912,N_19796,N_19220);
nand U20913 (N_20913,N_19896,N_19959);
nor U20914 (N_20914,N_19207,N_19169);
xor U20915 (N_20915,N_19680,N_19102);
xor U20916 (N_20916,N_19431,N_19534);
xor U20917 (N_20917,N_19430,N_19787);
and U20918 (N_20918,N_19452,N_19230);
and U20919 (N_20919,N_19148,N_19936);
xor U20920 (N_20920,N_19962,N_19254);
and U20921 (N_20921,N_19390,N_19527);
and U20922 (N_20922,N_19726,N_19018);
or U20923 (N_20923,N_19417,N_19653);
and U20924 (N_20924,N_19348,N_19975);
or U20925 (N_20925,N_19132,N_19171);
nor U20926 (N_20926,N_19103,N_19871);
or U20927 (N_20927,N_19169,N_19718);
nand U20928 (N_20928,N_19426,N_19269);
and U20929 (N_20929,N_19196,N_19399);
or U20930 (N_20930,N_19946,N_19224);
xnor U20931 (N_20931,N_19803,N_19843);
or U20932 (N_20932,N_19235,N_19173);
nand U20933 (N_20933,N_19224,N_19495);
and U20934 (N_20934,N_19747,N_19091);
xnor U20935 (N_20935,N_19288,N_19099);
xnor U20936 (N_20936,N_19935,N_19918);
nor U20937 (N_20937,N_19878,N_19883);
and U20938 (N_20938,N_19668,N_19818);
or U20939 (N_20939,N_19308,N_19254);
xnor U20940 (N_20940,N_19625,N_19924);
and U20941 (N_20941,N_19297,N_19330);
or U20942 (N_20942,N_19662,N_19873);
or U20943 (N_20943,N_19144,N_19460);
nor U20944 (N_20944,N_19050,N_19647);
nor U20945 (N_20945,N_19866,N_19278);
and U20946 (N_20946,N_19385,N_19497);
nor U20947 (N_20947,N_19913,N_19904);
and U20948 (N_20948,N_19264,N_19971);
nor U20949 (N_20949,N_19876,N_19690);
nor U20950 (N_20950,N_19505,N_19714);
nor U20951 (N_20951,N_19268,N_19881);
nand U20952 (N_20952,N_19641,N_19467);
nand U20953 (N_20953,N_19376,N_19162);
nand U20954 (N_20954,N_19517,N_19907);
or U20955 (N_20955,N_19994,N_19762);
and U20956 (N_20956,N_19000,N_19087);
or U20957 (N_20957,N_19557,N_19110);
or U20958 (N_20958,N_19088,N_19961);
xnor U20959 (N_20959,N_19026,N_19303);
xor U20960 (N_20960,N_19053,N_19617);
or U20961 (N_20961,N_19578,N_19896);
nor U20962 (N_20962,N_19744,N_19258);
xnor U20963 (N_20963,N_19855,N_19408);
nor U20964 (N_20964,N_19836,N_19988);
xnor U20965 (N_20965,N_19912,N_19420);
or U20966 (N_20966,N_19559,N_19118);
nand U20967 (N_20967,N_19853,N_19906);
or U20968 (N_20968,N_19332,N_19381);
or U20969 (N_20969,N_19429,N_19418);
nor U20970 (N_20970,N_19947,N_19384);
or U20971 (N_20971,N_19185,N_19957);
or U20972 (N_20972,N_19244,N_19251);
nand U20973 (N_20973,N_19543,N_19485);
nor U20974 (N_20974,N_19758,N_19972);
nand U20975 (N_20975,N_19814,N_19405);
or U20976 (N_20976,N_19167,N_19393);
nand U20977 (N_20977,N_19766,N_19628);
and U20978 (N_20978,N_19781,N_19760);
and U20979 (N_20979,N_19562,N_19971);
nor U20980 (N_20980,N_19910,N_19353);
or U20981 (N_20981,N_19666,N_19455);
or U20982 (N_20982,N_19445,N_19777);
xor U20983 (N_20983,N_19282,N_19723);
nand U20984 (N_20984,N_19164,N_19450);
nor U20985 (N_20985,N_19024,N_19330);
nand U20986 (N_20986,N_19271,N_19494);
or U20987 (N_20987,N_19738,N_19588);
nor U20988 (N_20988,N_19143,N_19750);
nand U20989 (N_20989,N_19397,N_19579);
nor U20990 (N_20990,N_19080,N_19010);
or U20991 (N_20991,N_19346,N_19087);
xor U20992 (N_20992,N_19782,N_19316);
and U20993 (N_20993,N_19774,N_19694);
or U20994 (N_20994,N_19953,N_19767);
and U20995 (N_20995,N_19811,N_19160);
or U20996 (N_20996,N_19545,N_19228);
nand U20997 (N_20997,N_19586,N_19591);
nand U20998 (N_20998,N_19222,N_19977);
nor U20999 (N_20999,N_19488,N_19748);
or U21000 (N_21000,N_20019,N_20945);
xor U21001 (N_21001,N_20709,N_20968);
and U21002 (N_21002,N_20859,N_20041);
nor U21003 (N_21003,N_20869,N_20635);
or U21004 (N_21004,N_20867,N_20233);
and U21005 (N_21005,N_20681,N_20285);
xor U21006 (N_21006,N_20797,N_20081);
and U21007 (N_21007,N_20316,N_20781);
xnor U21008 (N_21008,N_20282,N_20250);
nor U21009 (N_21009,N_20683,N_20536);
or U21010 (N_21010,N_20795,N_20470);
xnor U21011 (N_21011,N_20412,N_20409);
or U21012 (N_21012,N_20106,N_20070);
xor U21013 (N_21013,N_20909,N_20407);
or U21014 (N_21014,N_20135,N_20394);
or U21015 (N_21015,N_20473,N_20025);
and U21016 (N_21016,N_20446,N_20943);
nand U21017 (N_21017,N_20461,N_20191);
nand U21018 (N_21018,N_20879,N_20865);
and U21019 (N_21019,N_20200,N_20954);
nor U21020 (N_21020,N_20667,N_20239);
or U21021 (N_21021,N_20017,N_20918);
or U21022 (N_21022,N_20792,N_20207);
and U21023 (N_21023,N_20843,N_20028);
nor U21024 (N_21024,N_20161,N_20529);
nand U21025 (N_21025,N_20122,N_20910);
nand U21026 (N_21026,N_20054,N_20834);
and U21027 (N_21027,N_20671,N_20167);
nand U21028 (N_21028,N_20607,N_20690);
nand U21029 (N_21029,N_20352,N_20895);
xor U21030 (N_21030,N_20655,N_20182);
or U21031 (N_21031,N_20697,N_20720);
or U21032 (N_21032,N_20248,N_20705);
xnor U21033 (N_21033,N_20382,N_20469);
and U21034 (N_21034,N_20622,N_20351);
and U21035 (N_21035,N_20547,N_20863);
or U21036 (N_21036,N_20586,N_20058);
and U21037 (N_21037,N_20814,N_20732);
nand U21038 (N_21038,N_20179,N_20397);
and U21039 (N_21039,N_20296,N_20321);
xnor U21040 (N_21040,N_20903,N_20988);
xnor U21041 (N_21041,N_20114,N_20046);
nand U21042 (N_21042,N_20064,N_20127);
nor U21043 (N_21043,N_20454,N_20789);
nand U21044 (N_21044,N_20381,N_20308);
xnor U21045 (N_21045,N_20142,N_20436);
and U21046 (N_21046,N_20265,N_20383);
and U21047 (N_21047,N_20221,N_20953);
or U21048 (N_21048,N_20237,N_20348);
or U21049 (N_21049,N_20992,N_20568);
or U21050 (N_21050,N_20557,N_20659);
nand U21051 (N_21051,N_20688,N_20669);
and U21052 (N_21052,N_20026,N_20293);
nand U21053 (N_21053,N_20991,N_20978);
and U21054 (N_21054,N_20993,N_20141);
nor U21055 (N_21055,N_20483,N_20323);
and U21056 (N_21056,N_20481,N_20877);
nand U21057 (N_21057,N_20596,N_20636);
xor U21058 (N_21058,N_20353,N_20494);
or U21059 (N_21059,N_20180,N_20121);
and U21060 (N_21060,N_20914,N_20400);
nor U21061 (N_21061,N_20820,N_20042);
or U21062 (N_21062,N_20299,N_20260);
and U21063 (N_21063,N_20885,N_20662);
nor U21064 (N_21064,N_20768,N_20939);
and U21065 (N_21065,N_20804,N_20380);
nor U21066 (N_21066,N_20595,N_20949);
nand U21067 (N_21067,N_20350,N_20994);
xnor U21068 (N_21068,N_20816,N_20444);
or U21069 (N_21069,N_20823,N_20787);
nand U21070 (N_21070,N_20783,N_20424);
and U21071 (N_21071,N_20192,N_20388);
or U21072 (N_21072,N_20138,N_20246);
nand U21073 (N_21073,N_20916,N_20226);
and U21074 (N_21074,N_20827,N_20936);
or U21075 (N_21075,N_20396,N_20116);
nand U21076 (N_21076,N_20302,N_20230);
nand U21077 (N_21077,N_20585,N_20724);
and U21078 (N_21078,N_20187,N_20015);
nand U21079 (N_21079,N_20366,N_20673);
or U21080 (N_21080,N_20432,N_20218);
and U21081 (N_21081,N_20440,N_20000);
and U21082 (N_21082,N_20128,N_20984);
and U21083 (N_21083,N_20882,N_20220);
or U21084 (N_21084,N_20641,N_20008);
nor U21085 (N_21085,N_20088,N_20699);
xnor U21086 (N_21086,N_20848,N_20840);
nand U21087 (N_21087,N_20602,N_20307);
nand U21088 (N_21088,N_20811,N_20368);
xnor U21089 (N_21089,N_20420,N_20534);
nand U21090 (N_21090,N_20485,N_20457);
nor U21091 (N_21091,N_20247,N_20103);
nand U21092 (N_21092,N_20204,N_20793);
xor U21093 (N_21093,N_20467,N_20549);
nor U21094 (N_21094,N_20810,N_20267);
nor U21095 (N_21095,N_20005,N_20484);
nor U21096 (N_21096,N_20580,N_20670);
nor U21097 (N_21097,N_20309,N_20698);
nor U21098 (N_21098,N_20271,N_20137);
nand U21099 (N_21099,N_20259,N_20036);
xor U21100 (N_21100,N_20718,N_20480);
nand U21101 (N_21101,N_20740,N_20983);
and U21102 (N_21102,N_20962,N_20278);
nor U21103 (N_21103,N_20035,N_20047);
nor U21104 (N_21104,N_20244,N_20117);
nand U21105 (N_21105,N_20490,N_20208);
nor U21106 (N_21106,N_20492,N_20775);
or U21107 (N_21107,N_20704,N_20503);
nor U21108 (N_21108,N_20177,N_20249);
or U21109 (N_21109,N_20504,N_20707);
nand U21110 (N_21110,N_20361,N_20068);
or U21111 (N_21111,N_20158,N_20442);
nand U21112 (N_21112,N_20099,N_20798);
nor U21113 (N_21113,N_20448,N_20858);
or U21114 (N_21114,N_20710,N_20006);
nand U21115 (N_21115,N_20884,N_20313);
nand U21116 (N_21116,N_20059,N_20845);
xor U21117 (N_21117,N_20268,N_20819);
and U21118 (N_21118,N_20164,N_20876);
and U21119 (N_21119,N_20300,N_20971);
xnor U21120 (N_21120,N_20856,N_20927);
and U21121 (N_21121,N_20439,N_20986);
and U21122 (N_21122,N_20615,N_20033);
and U21123 (N_21123,N_20173,N_20152);
nand U21124 (N_21124,N_20011,N_20094);
nand U21125 (N_21125,N_20087,N_20241);
nand U21126 (N_21126,N_20433,N_20332);
and U21127 (N_21127,N_20889,N_20955);
or U21128 (N_21128,N_20371,N_20280);
nand U21129 (N_21129,N_20010,N_20051);
or U21130 (N_21130,N_20465,N_20419);
nor U21131 (N_21131,N_20112,N_20330);
or U21132 (N_21132,N_20832,N_20190);
nand U21133 (N_21133,N_20501,N_20611);
nand U21134 (N_21134,N_20500,N_20921);
xor U21135 (N_21135,N_20310,N_20703);
nor U21136 (N_21136,N_20555,N_20691);
and U21137 (N_21137,N_20211,N_20014);
or U21138 (N_21138,N_20657,N_20275);
and U21139 (N_21139,N_20303,N_20561);
nor U21140 (N_21140,N_20496,N_20893);
xnor U21141 (N_21141,N_20728,N_20423);
xor U21142 (N_21142,N_20734,N_20217);
nand U21143 (N_21143,N_20159,N_20739);
nor U21144 (N_21144,N_20023,N_20540);
xnor U21145 (N_21145,N_20813,N_20318);
xnor U21146 (N_21146,N_20196,N_20593);
and U21147 (N_21147,N_20076,N_20195);
xnor U21148 (N_21148,N_20377,N_20109);
nor U21149 (N_21149,N_20189,N_20385);
nor U21150 (N_21150,N_20078,N_20689);
nor U21151 (N_21151,N_20693,N_20007);
xor U21152 (N_21152,N_20924,N_20450);
or U21153 (N_21153,N_20564,N_20315);
nand U21154 (N_21154,N_20735,N_20842);
nand U21155 (N_21155,N_20578,N_20629);
xnor U21156 (N_21156,N_20966,N_20755);
nor U21157 (N_21157,N_20232,N_20590);
xor U21158 (N_21158,N_20676,N_20144);
and U21159 (N_21159,N_20526,N_20603);
xor U21160 (N_21160,N_20626,N_20995);
nand U21161 (N_21161,N_20651,N_20998);
nor U21162 (N_21162,N_20290,N_20235);
or U21163 (N_21163,N_20686,N_20123);
nand U21164 (N_21164,N_20741,N_20101);
xnor U21165 (N_21165,N_20415,N_20165);
or U21166 (N_21166,N_20880,N_20402);
or U21167 (N_21167,N_20086,N_20589);
and U21168 (N_21168,N_20980,N_20654);
and U21169 (N_21169,N_20289,N_20841);
and U21170 (N_21170,N_20941,N_20608);
or U21171 (N_21171,N_20069,N_20982);
xnor U21172 (N_21172,N_20610,N_20169);
nand U21173 (N_21173,N_20520,N_20521);
nor U21174 (N_21174,N_20393,N_20538);
nand U21175 (N_21175,N_20258,N_20126);
nor U21176 (N_21176,N_20493,N_20408);
or U21177 (N_21177,N_20134,N_20588);
or U21178 (N_21178,N_20652,N_20796);
xnor U21179 (N_21179,N_20738,N_20261);
xnor U21180 (N_21180,N_20899,N_20510);
xor U21181 (N_21181,N_20364,N_20614);
nor U21182 (N_21182,N_20294,N_20306);
nor U21183 (N_21183,N_20030,N_20786);
xor U21184 (N_21184,N_20194,N_20723);
and U21185 (N_21185,N_20482,N_20012);
nand U21186 (N_21186,N_20852,N_20486);
xor U21187 (N_21187,N_20210,N_20276);
xor U21188 (N_21188,N_20744,N_20021);
or U21189 (N_21189,N_20176,N_20150);
or U21190 (N_21190,N_20868,N_20048);
and U21191 (N_21191,N_20600,N_20097);
xnor U21192 (N_21192,N_20038,N_20253);
nor U21193 (N_21193,N_20245,N_20319);
or U21194 (N_21194,N_20024,N_20228);
nor U21195 (N_21195,N_20696,N_20763);
nor U21196 (N_21196,N_20251,N_20748);
or U21197 (N_21197,N_20767,N_20760);
xor U21198 (N_21198,N_20085,N_20912);
or U21199 (N_21199,N_20314,N_20851);
and U21200 (N_21200,N_20073,N_20799);
and U21201 (N_21201,N_20757,N_20824);
and U21202 (N_21202,N_20238,N_20131);
or U21203 (N_21203,N_20902,N_20900);
nand U21204 (N_21204,N_20964,N_20630);
or U21205 (N_21205,N_20650,N_20782);
or U21206 (N_21206,N_20612,N_20206);
or U21207 (N_21207,N_20032,N_20989);
or U21208 (N_21208,N_20414,N_20441);
or U21209 (N_21209,N_20581,N_20618);
xor U21210 (N_21210,N_20277,N_20960);
and U21211 (N_21211,N_20874,N_20777);
nor U21212 (N_21212,N_20171,N_20297);
or U21213 (N_21213,N_20411,N_20427);
nand U21214 (N_21214,N_20067,N_20742);
nand U21215 (N_21215,N_20359,N_20556);
nor U21216 (N_21216,N_20052,N_20236);
nand U21217 (N_21217,N_20719,N_20129);
xor U21218 (N_21218,N_20766,N_20716);
or U21219 (N_21219,N_20507,N_20160);
xnor U21220 (N_21220,N_20802,N_20771);
or U21221 (N_21221,N_20202,N_20756);
and U21222 (N_21222,N_20682,N_20996);
and U21223 (N_21223,N_20497,N_20357);
nor U21224 (N_21224,N_20562,N_20864);
nor U21225 (N_21225,N_20554,N_20034);
or U21226 (N_21226,N_20475,N_20234);
nor U21227 (N_21227,N_20198,N_20892);
xor U21228 (N_21228,N_20107,N_20649);
nand U21229 (N_21229,N_20931,N_20706);
nor U21230 (N_21230,N_20929,N_20515);
and U21231 (N_21231,N_20794,N_20273);
nand U21232 (N_21232,N_20074,N_20336);
or U21233 (N_21233,N_20460,N_20754);
and U21234 (N_21234,N_20431,N_20045);
or U21235 (N_21235,N_20745,N_20115);
nor U21236 (N_21236,N_20222,N_20360);
xnor U21237 (N_21237,N_20214,N_20404);
xor U21238 (N_21238,N_20301,N_20124);
and U21239 (N_21239,N_20132,N_20624);
nor U21240 (N_21240,N_20712,N_20977);
or U21241 (N_21241,N_20317,N_20219);
or U21242 (N_21242,N_20295,N_20434);
nand U21243 (N_21243,N_20209,N_20039);
or U21244 (N_21244,N_20616,N_20896);
nor U21245 (N_21245,N_20040,N_20018);
or U21246 (N_21246,N_20257,N_20660);
nor U21247 (N_21247,N_20417,N_20826);
and U21248 (N_21248,N_20619,N_20764);
nor U21249 (N_21249,N_20333,N_20174);
or U21250 (N_21250,N_20110,N_20471);
xnor U21251 (N_21251,N_20778,N_20283);
nand U21252 (N_21252,N_20188,N_20027);
or U21253 (N_21253,N_20558,N_20288);
and U21254 (N_21254,N_20438,N_20565);
and U21255 (N_21255,N_20425,N_20606);
nand U21256 (N_21256,N_20592,N_20508);
nor U21257 (N_21257,N_20653,N_20057);
or U21258 (N_21258,N_20906,N_20911);
and U21259 (N_21259,N_20937,N_20981);
or U21260 (N_21260,N_20518,N_20747);
xnor U21261 (N_21261,N_20472,N_20844);
or U21262 (N_21262,N_20965,N_20729);
and U21263 (N_21263,N_20274,N_20574);
nand U21264 (N_21264,N_20113,N_20525);
xnor U21265 (N_21265,N_20118,N_20016);
nand U21266 (N_21266,N_20416,N_20464);
or U21267 (N_21267,N_20715,N_20779);
nand U21268 (N_21268,N_20551,N_20263);
or U21269 (N_21269,N_20356,N_20083);
nand U21270 (N_21270,N_20104,N_20587);
and U21271 (N_21271,N_20505,N_20020);
xor U21272 (N_21272,N_20506,N_20095);
xor U21273 (N_21273,N_20146,N_20346);
nand U21274 (N_21274,N_20969,N_20362);
xnor U21275 (N_21275,N_20695,N_20495);
or U21276 (N_21276,N_20203,N_20722);
or U21277 (N_21277,N_20976,N_20455);
or U21278 (N_21278,N_20835,N_20163);
and U21279 (N_21279,N_20421,N_20759);
and U21280 (N_21280,N_20942,N_20817);
nand U21281 (N_21281,N_20511,N_20328);
nor U21282 (N_21282,N_20063,N_20435);
xnor U21283 (N_21283,N_20426,N_20084);
or U21284 (N_21284,N_20546,N_20270);
nor U21285 (N_21285,N_20363,N_20948);
or U21286 (N_21286,N_20527,N_20430);
and U21287 (N_21287,N_20451,N_20956);
and U21288 (N_21288,N_20347,N_20001);
and U21289 (N_21289,N_20139,N_20774);
and U21290 (N_21290,N_20224,N_20919);
nor U21291 (N_21291,N_20279,N_20231);
or U21292 (N_21292,N_20866,N_20502);
and U21293 (N_21293,N_20913,N_20523);
and U21294 (N_21294,N_20331,N_20049);
and U21295 (N_21295,N_20367,N_20684);
xnor U21296 (N_21296,N_20120,N_20379);
or U21297 (N_21297,N_20456,N_20157);
xnor U21298 (N_21298,N_20569,N_20952);
nand U21299 (N_21299,N_20644,N_20447);
nor U21300 (N_21300,N_20901,N_20638);
nand U21301 (N_21301,N_20335,N_20055);
xnor U21302 (N_21302,N_20805,N_20609);
or U21303 (N_21303,N_20422,N_20656);
or U21304 (N_21304,N_20583,N_20401);
or U21305 (N_21305,N_20898,N_20077);
xnor U21306 (N_21306,N_20050,N_20098);
nor U21307 (N_21307,N_20997,N_20979);
nor U21308 (N_21308,N_20240,N_20631);
and U21309 (N_21309,N_20013,N_20700);
and U21310 (N_21310,N_20272,N_20543);
and U21311 (N_21311,N_20329,N_20664);
or U21312 (N_21312,N_20658,N_20100);
nor U21313 (N_21313,N_20545,N_20837);
xnor U21314 (N_21314,N_20762,N_20907);
nand U21315 (N_21315,N_20476,N_20009);
and U21316 (N_21316,N_20354,N_20256);
nand U21317 (N_21317,N_20509,N_20125);
and U21318 (N_21318,N_20524,N_20037);
nor U21319 (N_21319,N_20111,N_20389);
nand U21320 (N_21320,N_20711,N_20855);
or U21321 (N_21321,N_20839,N_20205);
nor U21322 (N_21322,N_20946,N_20881);
and U21323 (N_21323,N_20730,N_20854);
or U21324 (N_21324,N_20452,N_20458);
nand U21325 (N_21325,N_20242,N_20891);
or U21326 (N_21326,N_20053,N_20384);
nand U21327 (N_21327,N_20186,N_20633);
nand U21328 (N_21328,N_20090,N_20254);
nor U21329 (N_21329,N_20340,N_20533);
nand U21330 (N_21330,N_20604,N_20692);
or U21331 (N_21331,N_20894,N_20575);
xnor U21332 (N_21332,N_20872,N_20570);
nand U21333 (N_21333,N_20072,N_20229);
nand U21334 (N_21334,N_20080,N_20553);
and U21335 (N_21335,N_20957,N_20365);
nand U21336 (N_21336,N_20803,N_20445);
and U21337 (N_21337,N_20031,N_20769);
or U21338 (N_21338,N_20950,N_20579);
xnor U21339 (N_21339,N_20043,N_20643);
nor U21340 (N_21340,N_20065,N_20305);
xor U21341 (N_21341,N_20974,N_20522);
xor U21342 (N_21342,N_20512,N_20871);
nor U21343 (N_21343,N_20286,N_20888);
nand U21344 (N_21344,N_20550,N_20628);
nor U21345 (N_21345,N_20930,N_20905);
or U21346 (N_21346,N_20646,N_20625);
nand U21347 (N_21347,N_20772,N_20062);
and U21348 (N_21348,N_20990,N_20639);
and U21349 (N_21349,N_20358,N_20985);
or U21350 (N_21350,N_20560,N_20532);
or U21351 (N_21351,N_20822,N_20721);
nand U21352 (N_21352,N_20599,N_20082);
and U21353 (N_21353,N_20645,N_20665);
or U21354 (N_21354,N_20694,N_20491);
nor U21355 (N_21355,N_20369,N_20535);
and U21356 (N_21356,N_20002,N_20634);
or U21357 (N_21357,N_20264,N_20743);
and U21358 (N_21358,N_20847,N_20136);
nand U21359 (N_21359,N_20725,N_20003);
xor U21360 (N_21360,N_20806,N_20726);
nand U21361 (N_21361,N_20373,N_20934);
or U21362 (N_21362,N_20405,N_20374);
or U21363 (N_21363,N_20514,N_20620);
and U21364 (N_21364,N_20197,N_20920);
nand U21365 (N_21365,N_20531,N_20119);
and U21366 (N_21366,N_20341,N_20075);
or U21367 (N_21367,N_20917,N_20386);
nor U21368 (N_21368,N_20212,N_20582);
xnor U21369 (N_21369,N_20459,N_20621);
xnor U21370 (N_21370,N_20466,N_20923);
or U21371 (N_21371,N_20761,N_20327);
xnor U21372 (N_21372,N_20216,N_20701);
nor U21373 (N_21373,N_20833,N_20828);
nor U21374 (N_21374,N_20963,N_20105);
xor U21375 (N_21375,N_20972,N_20821);
nor U21376 (N_21376,N_20029,N_20398);
or U21377 (N_21377,N_20825,N_20155);
and U21378 (N_21378,N_20453,N_20344);
nor U21379 (N_21379,N_20838,N_20750);
or U21380 (N_21380,N_20784,N_20181);
and U21381 (N_21381,N_20944,N_20970);
xor U21382 (N_21382,N_20809,N_20175);
xor U21383 (N_21383,N_20737,N_20668);
xor U21384 (N_21384,N_20935,N_20544);
and U21385 (N_21385,N_20370,N_20566);
or U21386 (N_21386,N_20498,N_20056);
nand U21387 (N_21387,N_20479,N_20375);
or U21388 (N_21388,N_20349,N_20951);
and U21389 (N_21389,N_20145,N_20800);
or U21390 (N_21390,N_20790,N_20717);
nand U21391 (N_21391,N_20940,N_20975);
nor U21392 (N_21392,N_20890,N_20227);
nand U21393 (N_21393,N_20573,N_20462);
or U21394 (N_21394,N_20168,N_20713);
nor U21395 (N_21395,N_20322,N_20185);
and U21396 (N_21396,N_20861,N_20584);
and U21397 (N_21397,N_20973,N_20287);
or U21398 (N_21398,N_20304,N_20147);
nor U21399 (N_21399,N_20831,N_20675);
or U21400 (N_21400,N_20887,N_20102);
nand U21401 (N_21401,N_20926,N_20812);
and U21402 (N_21402,N_20378,N_20829);
nor U21403 (N_21403,N_20666,N_20291);
xnor U21404 (N_21404,N_20623,N_20266);
nand U21405 (N_21405,N_20904,N_20915);
or U21406 (N_21406,N_20345,N_20878);
or U21407 (N_21407,N_20680,N_20079);
nor U21408 (N_21408,N_20199,N_20488);
and U21409 (N_21409,N_20776,N_20066);
nand U21410 (N_21410,N_20463,N_20958);
and U21411 (N_21411,N_20849,N_20243);
nand U21412 (N_21412,N_20674,N_20752);
nor U21413 (N_21413,N_20537,N_20807);
nand U21414 (N_21414,N_20961,N_20836);
or U21415 (N_21415,N_20642,N_20292);
nor U21416 (N_21416,N_20516,N_20947);
and U21417 (N_21417,N_20133,N_20928);
xor U21418 (N_21418,N_20753,N_20539);
and U21419 (N_21419,N_20572,N_20938);
or U21420 (N_21420,N_20418,N_20376);
xor U21421 (N_21421,N_20959,N_20342);
nor U21422 (N_21422,N_20967,N_20213);
xnor U21423 (N_21423,N_20474,N_20791);
or U21424 (N_21424,N_20758,N_20428);
nor U21425 (N_21425,N_20044,N_20178);
and U21426 (N_21426,N_20410,N_20403);
nor U21427 (N_21427,N_20343,N_20677);
nor U21428 (N_21428,N_20326,N_20765);
and U21429 (N_21429,N_20387,N_20223);
xnor U21430 (N_21430,N_20391,N_20801);
xor U21431 (N_21431,N_20563,N_20339);
and U21432 (N_21432,N_20089,N_20148);
xor U21433 (N_21433,N_20437,N_20468);
nand U21434 (N_21434,N_20255,N_20156);
and U21435 (N_21435,N_20685,N_20818);
xnor U21436 (N_21436,N_20215,N_20727);
and U21437 (N_21437,N_20857,N_20672);
nor U21438 (N_21438,N_20092,N_20311);
nand U21439 (N_21439,N_20225,N_20637);
nor U21440 (N_21440,N_20172,N_20022);
and U21441 (N_21441,N_20542,N_20337);
nand U21442 (N_21442,N_20846,N_20751);
xor U21443 (N_21443,N_20183,N_20749);
nand U21444 (N_21444,N_20334,N_20541);
and U21445 (N_21445,N_20489,N_20567);
and U21446 (N_21446,N_20091,N_20449);
nor U21447 (N_21447,N_20850,N_20162);
and U21448 (N_21448,N_20594,N_20519);
or U21449 (N_21449,N_20853,N_20605);
nand U21450 (N_21450,N_20269,N_20298);
and U21451 (N_21451,N_20613,N_20576);
nand U21452 (N_21452,N_20154,N_20151);
xnor U21453 (N_21453,N_20780,N_20886);
and U21454 (N_21454,N_20143,N_20193);
nand U21455 (N_21455,N_20736,N_20478);
xnor U21456 (N_21456,N_20108,N_20617);
xor U21457 (N_21457,N_20548,N_20678);
nor U21458 (N_21458,N_20788,N_20601);
or U21459 (N_21459,N_20252,N_20281);
xor U21460 (N_21460,N_20773,N_20663);
or U21461 (N_21461,N_20443,N_20679);
nand U21462 (N_21462,N_20140,N_20399);
nand U21463 (N_21463,N_20395,N_20325);
nor U21464 (N_21464,N_20731,N_20770);
xnor U21465 (N_21465,N_20627,N_20096);
nand U21466 (N_21466,N_20922,N_20093);
and U21467 (N_21467,N_20648,N_20413);
nand U21468 (N_21468,N_20390,N_20830);
or U21469 (N_21469,N_20597,N_20513);
and U21470 (N_21470,N_20355,N_20708);
and U21471 (N_21471,N_20591,N_20487);
and U21472 (N_21472,N_20687,N_20528);
and U21473 (N_21473,N_20184,N_20130);
nand U21474 (N_21474,N_20999,N_20647);
or U21475 (N_21475,N_20987,N_20873);
xor U21476 (N_21476,N_20429,N_20632);
and U21477 (N_21477,N_20571,N_20559);
xnor U21478 (N_21478,N_20517,N_20933);
nor U21479 (N_21479,N_20808,N_20061);
nor U21480 (N_21480,N_20733,N_20925);
xor U21481 (N_21481,N_20153,N_20284);
xnor U21482 (N_21482,N_20702,N_20714);
xnor U21483 (N_21483,N_20883,N_20166);
and U21484 (N_21484,N_20661,N_20870);
nand U21485 (N_21485,N_20785,N_20060);
xor U21486 (N_21486,N_20149,N_20477);
xnor U21487 (N_21487,N_20577,N_20372);
nor U21488 (N_21488,N_20499,N_20406);
nor U21489 (N_21489,N_20530,N_20815);
nand U21490 (N_21490,N_20071,N_20170);
xor U21491 (N_21491,N_20875,N_20908);
and U21492 (N_21492,N_20552,N_20860);
nand U21493 (N_21493,N_20201,N_20862);
and U21494 (N_21494,N_20338,N_20640);
xnor U21495 (N_21495,N_20004,N_20324);
or U21496 (N_21496,N_20312,N_20932);
and U21497 (N_21497,N_20746,N_20897);
nand U21498 (N_21498,N_20392,N_20598);
xor U21499 (N_21499,N_20262,N_20320);
nor U21500 (N_21500,N_20200,N_20937);
nand U21501 (N_21501,N_20184,N_20332);
xnor U21502 (N_21502,N_20222,N_20382);
nor U21503 (N_21503,N_20171,N_20107);
or U21504 (N_21504,N_20286,N_20360);
or U21505 (N_21505,N_20951,N_20647);
nor U21506 (N_21506,N_20317,N_20214);
and U21507 (N_21507,N_20968,N_20523);
nor U21508 (N_21508,N_20944,N_20409);
and U21509 (N_21509,N_20345,N_20996);
nor U21510 (N_21510,N_20545,N_20740);
nor U21511 (N_21511,N_20633,N_20513);
nor U21512 (N_21512,N_20328,N_20745);
and U21513 (N_21513,N_20798,N_20735);
or U21514 (N_21514,N_20084,N_20363);
and U21515 (N_21515,N_20949,N_20537);
and U21516 (N_21516,N_20503,N_20302);
xnor U21517 (N_21517,N_20700,N_20582);
xnor U21518 (N_21518,N_20441,N_20206);
or U21519 (N_21519,N_20612,N_20199);
nor U21520 (N_21520,N_20207,N_20147);
nor U21521 (N_21521,N_20209,N_20555);
and U21522 (N_21522,N_20148,N_20623);
xnor U21523 (N_21523,N_20849,N_20815);
xnor U21524 (N_21524,N_20666,N_20247);
and U21525 (N_21525,N_20639,N_20598);
nand U21526 (N_21526,N_20237,N_20166);
nor U21527 (N_21527,N_20862,N_20311);
nand U21528 (N_21528,N_20383,N_20456);
or U21529 (N_21529,N_20142,N_20017);
nand U21530 (N_21530,N_20035,N_20633);
or U21531 (N_21531,N_20070,N_20827);
and U21532 (N_21532,N_20113,N_20475);
and U21533 (N_21533,N_20990,N_20562);
and U21534 (N_21534,N_20577,N_20419);
nand U21535 (N_21535,N_20797,N_20548);
nor U21536 (N_21536,N_20999,N_20060);
and U21537 (N_21537,N_20280,N_20387);
and U21538 (N_21538,N_20367,N_20531);
or U21539 (N_21539,N_20400,N_20728);
nand U21540 (N_21540,N_20332,N_20283);
and U21541 (N_21541,N_20705,N_20807);
nand U21542 (N_21542,N_20373,N_20733);
nor U21543 (N_21543,N_20376,N_20427);
nand U21544 (N_21544,N_20451,N_20928);
nand U21545 (N_21545,N_20976,N_20985);
or U21546 (N_21546,N_20930,N_20618);
nand U21547 (N_21547,N_20437,N_20952);
xnor U21548 (N_21548,N_20565,N_20031);
nand U21549 (N_21549,N_20058,N_20399);
or U21550 (N_21550,N_20180,N_20054);
nor U21551 (N_21551,N_20262,N_20182);
nand U21552 (N_21552,N_20673,N_20112);
and U21553 (N_21553,N_20296,N_20037);
nor U21554 (N_21554,N_20487,N_20474);
or U21555 (N_21555,N_20884,N_20335);
nand U21556 (N_21556,N_20820,N_20364);
or U21557 (N_21557,N_20621,N_20920);
or U21558 (N_21558,N_20437,N_20593);
or U21559 (N_21559,N_20148,N_20171);
nor U21560 (N_21560,N_20419,N_20018);
xor U21561 (N_21561,N_20029,N_20748);
nor U21562 (N_21562,N_20618,N_20892);
nand U21563 (N_21563,N_20761,N_20426);
and U21564 (N_21564,N_20040,N_20074);
and U21565 (N_21565,N_20382,N_20687);
nand U21566 (N_21566,N_20736,N_20752);
or U21567 (N_21567,N_20360,N_20292);
nand U21568 (N_21568,N_20774,N_20429);
nor U21569 (N_21569,N_20026,N_20294);
nor U21570 (N_21570,N_20388,N_20311);
nor U21571 (N_21571,N_20699,N_20840);
nor U21572 (N_21572,N_20181,N_20244);
nor U21573 (N_21573,N_20075,N_20029);
or U21574 (N_21574,N_20982,N_20705);
and U21575 (N_21575,N_20551,N_20983);
nand U21576 (N_21576,N_20211,N_20738);
or U21577 (N_21577,N_20718,N_20038);
or U21578 (N_21578,N_20756,N_20310);
xor U21579 (N_21579,N_20032,N_20307);
nor U21580 (N_21580,N_20151,N_20569);
nand U21581 (N_21581,N_20478,N_20283);
and U21582 (N_21582,N_20309,N_20630);
xnor U21583 (N_21583,N_20600,N_20477);
and U21584 (N_21584,N_20087,N_20834);
xnor U21585 (N_21585,N_20963,N_20013);
xor U21586 (N_21586,N_20527,N_20602);
xor U21587 (N_21587,N_20611,N_20475);
and U21588 (N_21588,N_20373,N_20421);
xor U21589 (N_21589,N_20077,N_20808);
or U21590 (N_21590,N_20706,N_20522);
and U21591 (N_21591,N_20888,N_20490);
xor U21592 (N_21592,N_20939,N_20960);
xnor U21593 (N_21593,N_20257,N_20935);
or U21594 (N_21594,N_20267,N_20549);
xnor U21595 (N_21595,N_20421,N_20883);
and U21596 (N_21596,N_20817,N_20807);
nor U21597 (N_21597,N_20844,N_20628);
and U21598 (N_21598,N_20277,N_20095);
or U21599 (N_21599,N_20454,N_20844);
xnor U21600 (N_21600,N_20564,N_20189);
nor U21601 (N_21601,N_20406,N_20724);
nor U21602 (N_21602,N_20405,N_20991);
and U21603 (N_21603,N_20941,N_20903);
xnor U21604 (N_21604,N_20082,N_20990);
and U21605 (N_21605,N_20676,N_20508);
and U21606 (N_21606,N_20473,N_20798);
and U21607 (N_21607,N_20523,N_20601);
or U21608 (N_21608,N_20767,N_20915);
nand U21609 (N_21609,N_20593,N_20478);
or U21610 (N_21610,N_20119,N_20634);
nor U21611 (N_21611,N_20931,N_20563);
nor U21612 (N_21612,N_20731,N_20925);
xnor U21613 (N_21613,N_20647,N_20166);
or U21614 (N_21614,N_20256,N_20190);
and U21615 (N_21615,N_20661,N_20492);
or U21616 (N_21616,N_20615,N_20193);
xor U21617 (N_21617,N_20416,N_20128);
nor U21618 (N_21618,N_20058,N_20779);
nand U21619 (N_21619,N_20349,N_20539);
or U21620 (N_21620,N_20247,N_20144);
nor U21621 (N_21621,N_20352,N_20639);
nor U21622 (N_21622,N_20347,N_20751);
or U21623 (N_21623,N_20610,N_20248);
xor U21624 (N_21624,N_20143,N_20579);
nor U21625 (N_21625,N_20927,N_20582);
or U21626 (N_21626,N_20368,N_20033);
xnor U21627 (N_21627,N_20557,N_20773);
nand U21628 (N_21628,N_20563,N_20552);
nor U21629 (N_21629,N_20893,N_20925);
nor U21630 (N_21630,N_20574,N_20428);
and U21631 (N_21631,N_20488,N_20621);
and U21632 (N_21632,N_20745,N_20428);
nand U21633 (N_21633,N_20711,N_20376);
xnor U21634 (N_21634,N_20200,N_20782);
and U21635 (N_21635,N_20267,N_20092);
or U21636 (N_21636,N_20282,N_20956);
xor U21637 (N_21637,N_20610,N_20069);
and U21638 (N_21638,N_20156,N_20458);
nor U21639 (N_21639,N_20605,N_20023);
and U21640 (N_21640,N_20103,N_20797);
and U21641 (N_21641,N_20899,N_20427);
xor U21642 (N_21642,N_20254,N_20800);
xnor U21643 (N_21643,N_20847,N_20315);
nor U21644 (N_21644,N_20389,N_20254);
nor U21645 (N_21645,N_20427,N_20109);
nor U21646 (N_21646,N_20728,N_20116);
nand U21647 (N_21647,N_20722,N_20531);
or U21648 (N_21648,N_20775,N_20807);
nand U21649 (N_21649,N_20154,N_20410);
nand U21650 (N_21650,N_20234,N_20440);
and U21651 (N_21651,N_20283,N_20246);
nand U21652 (N_21652,N_20579,N_20479);
and U21653 (N_21653,N_20771,N_20380);
xnor U21654 (N_21654,N_20921,N_20528);
nand U21655 (N_21655,N_20990,N_20314);
and U21656 (N_21656,N_20553,N_20393);
nand U21657 (N_21657,N_20153,N_20125);
and U21658 (N_21658,N_20945,N_20159);
and U21659 (N_21659,N_20968,N_20849);
nor U21660 (N_21660,N_20107,N_20038);
xnor U21661 (N_21661,N_20222,N_20088);
nor U21662 (N_21662,N_20637,N_20149);
and U21663 (N_21663,N_20355,N_20312);
and U21664 (N_21664,N_20225,N_20439);
or U21665 (N_21665,N_20772,N_20900);
or U21666 (N_21666,N_20143,N_20073);
or U21667 (N_21667,N_20044,N_20621);
nor U21668 (N_21668,N_20442,N_20564);
xor U21669 (N_21669,N_20550,N_20723);
or U21670 (N_21670,N_20727,N_20904);
and U21671 (N_21671,N_20814,N_20780);
and U21672 (N_21672,N_20016,N_20444);
or U21673 (N_21673,N_20127,N_20659);
or U21674 (N_21674,N_20131,N_20445);
or U21675 (N_21675,N_20554,N_20051);
and U21676 (N_21676,N_20457,N_20096);
and U21677 (N_21677,N_20505,N_20144);
and U21678 (N_21678,N_20724,N_20926);
nor U21679 (N_21679,N_20573,N_20324);
nor U21680 (N_21680,N_20164,N_20685);
nor U21681 (N_21681,N_20623,N_20075);
xor U21682 (N_21682,N_20451,N_20979);
nand U21683 (N_21683,N_20115,N_20928);
and U21684 (N_21684,N_20351,N_20833);
and U21685 (N_21685,N_20167,N_20772);
xor U21686 (N_21686,N_20622,N_20499);
xor U21687 (N_21687,N_20085,N_20521);
and U21688 (N_21688,N_20624,N_20262);
nand U21689 (N_21689,N_20014,N_20520);
nor U21690 (N_21690,N_20197,N_20975);
nor U21691 (N_21691,N_20918,N_20528);
nand U21692 (N_21692,N_20827,N_20454);
nor U21693 (N_21693,N_20684,N_20604);
or U21694 (N_21694,N_20615,N_20175);
and U21695 (N_21695,N_20675,N_20670);
and U21696 (N_21696,N_20555,N_20925);
xnor U21697 (N_21697,N_20672,N_20943);
nand U21698 (N_21698,N_20260,N_20582);
nand U21699 (N_21699,N_20321,N_20668);
or U21700 (N_21700,N_20463,N_20735);
and U21701 (N_21701,N_20750,N_20211);
nor U21702 (N_21702,N_20878,N_20847);
xnor U21703 (N_21703,N_20689,N_20301);
xor U21704 (N_21704,N_20627,N_20433);
xor U21705 (N_21705,N_20584,N_20317);
xor U21706 (N_21706,N_20686,N_20515);
or U21707 (N_21707,N_20563,N_20864);
and U21708 (N_21708,N_20721,N_20573);
xor U21709 (N_21709,N_20631,N_20065);
and U21710 (N_21710,N_20773,N_20673);
or U21711 (N_21711,N_20697,N_20925);
or U21712 (N_21712,N_20473,N_20403);
and U21713 (N_21713,N_20372,N_20488);
nand U21714 (N_21714,N_20492,N_20806);
nor U21715 (N_21715,N_20847,N_20816);
or U21716 (N_21716,N_20853,N_20259);
or U21717 (N_21717,N_20920,N_20993);
or U21718 (N_21718,N_20232,N_20422);
xnor U21719 (N_21719,N_20448,N_20746);
xor U21720 (N_21720,N_20463,N_20323);
nor U21721 (N_21721,N_20989,N_20717);
or U21722 (N_21722,N_20036,N_20049);
nor U21723 (N_21723,N_20670,N_20860);
nor U21724 (N_21724,N_20958,N_20007);
and U21725 (N_21725,N_20310,N_20373);
xnor U21726 (N_21726,N_20213,N_20898);
nand U21727 (N_21727,N_20139,N_20445);
or U21728 (N_21728,N_20433,N_20884);
xnor U21729 (N_21729,N_20624,N_20270);
xnor U21730 (N_21730,N_20771,N_20892);
and U21731 (N_21731,N_20013,N_20948);
or U21732 (N_21732,N_20775,N_20593);
and U21733 (N_21733,N_20665,N_20921);
and U21734 (N_21734,N_20667,N_20716);
and U21735 (N_21735,N_20464,N_20713);
or U21736 (N_21736,N_20276,N_20773);
nor U21737 (N_21737,N_20237,N_20803);
or U21738 (N_21738,N_20672,N_20263);
xor U21739 (N_21739,N_20157,N_20161);
and U21740 (N_21740,N_20703,N_20602);
and U21741 (N_21741,N_20771,N_20390);
or U21742 (N_21742,N_20608,N_20931);
or U21743 (N_21743,N_20157,N_20272);
and U21744 (N_21744,N_20408,N_20124);
xnor U21745 (N_21745,N_20311,N_20161);
and U21746 (N_21746,N_20253,N_20707);
nor U21747 (N_21747,N_20737,N_20574);
xor U21748 (N_21748,N_20559,N_20761);
or U21749 (N_21749,N_20904,N_20043);
and U21750 (N_21750,N_20230,N_20014);
nor U21751 (N_21751,N_20075,N_20248);
and U21752 (N_21752,N_20287,N_20391);
and U21753 (N_21753,N_20824,N_20745);
and U21754 (N_21754,N_20937,N_20285);
nand U21755 (N_21755,N_20950,N_20947);
nor U21756 (N_21756,N_20371,N_20059);
nand U21757 (N_21757,N_20941,N_20565);
and U21758 (N_21758,N_20512,N_20554);
nor U21759 (N_21759,N_20898,N_20441);
or U21760 (N_21760,N_20987,N_20051);
and U21761 (N_21761,N_20292,N_20834);
and U21762 (N_21762,N_20028,N_20329);
nand U21763 (N_21763,N_20173,N_20196);
xor U21764 (N_21764,N_20099,N_20174);
or U21765 (N_21765,N_20858,N_20889);
xnor U21766 (N_21766,N_20165,N_20953);
or U21767 (N_21767,N_20036,N_20102);
nand U21768 (N_21768,N_20684,N_20735);
or U21769 (N_21769,N_20731,N_20057);
xnor U21770 (N_21770,N_20034,N_20246);
or U21771 (N_21771,N_20780,N_20204);
nor U21772 (N_21772,N_20286,N_20134);
and U21773 (N_21773,N_20744,N_20135);
nor U21774 (N_21774,N_20627,N_20761);
nand U21775 (N_21775,N_20077,N_20703);
xnor U21776 (N_21776,N_20753,N_20923);
nand U21777 (N_21777,N_20789,N_20318);
nor U21778 (N_21778,N_20544,N_20419);
or U21779 (N_21779,N_20254,N_20211);
xnor U21780 (N_21780,N_20051,N_20773);
xnor U21781 (N_21781,N_20827,N_20588);
xnor U21782 (N_21782,N_20133,N_20888);
nor U21783 (N_21783,N_20383,N_20155);
or U21784 (N_21784,N_20404,N_20513);
nor U21785 (N_21785,N_20350,N_20477);
and U21786 (N_21786,N_20462,N_20753);
and U21787 (N_21787,N_20024,N_20171);
nor U21788 (N_21788,N_20577,N_20491);
and U21789 (N_21789,N_20366,N_20168);
xor U21790 (N_21790,N_20131,N_20637);
nand U21791 (N_21791,N_20626,N_20811);
xnor U21792 (N_21792,N_20631,N_20392);
nand U21793 (N_21793,N_20624,N_20220);
nand U21794 (N_21794,N_20523,N_20887);
and U21795 (N_21795,N_20906,N_20087);
and U21796 (N_21796,N_20232,N_20352);
nand U21797 (N_21797,N_20101,N_20325);
xnor U21798 (N_21798,N_20115,N_20483);
nor U21799 (N_21799,N_20345,N_20769);
nor U21800 (N_21800,N_20122,N_20967);
or U21801 (N_21801,N_20148,N_20404);
nand U21802 (N_21802,N_20276,N_20751);
nand U21803 (N_21803,N_20833,N_20887);
or U21804 (N_21804,N_20270,N_20072);
nand U21805 (N_21805,N_20457,N_20370);
and U21806 (N_21806,N_20702,N_20292);
or U21807 (N_21807,N_20640,N_20957);
or U21808 (N_21808,N_20295,N_20696);
nand U21809 (N_21809,N_20680,N_20343);
nand U21810 (N_21810,N_20209,N_20394);
and U21811 (N_21811,N_20267,N_20400);
or U21812 (N_21812,N_20904,N_20817);
nor U21813 (N_21813,N_20720,N_20583);
nor U21814 (N_21814,N_20759,N_20603);
nor U21815 (N_21815,N_20808,N_20884);
nand U21816 (N_21816,N_20996,N_20184);
and U21817 (N_21817,N_20926,N_20351);
and U21818 (N_21818,N_20755,N_20426);
nand U21819 (N_21819,N_20318,N_20013);
and U21820 (N_21820,N_20065,N_20517);
or U21821 (N_21821,N_20906,N_20226);
nor U21822 (N_21822,N_20201,N_20141);
or U21823 (N_21823,N_20449,N_20381);
nor U21824 (N_21824,N_20608,N_20437);
or U21825 (N_21825,N_20582,N_20141);
xnor U21826 (N_21826,N_20527,N_20693);
nand U21827 (N_21827,N_20260,N_20911);
and U21828 (N_21828,N_20799,N_20749);
nor U21829 (N_21829,N_20668,N_20858);
nor U21830 (N_21830,N_20812,N_20776);
nand U21831 (N_21831,N_20702,N_20574);
and U21832 (N_21832,N_20400,N_20554);
nor U21833 (N_21833,N_20577,N_20000);
or U21834 (N_21834,N_20742,N_20029);
and U21835 (N_21835,N_20088,N_20883);
xor U21836 (N_21836,N_20578,N_20636);
xor U21837 (N_21837,N_20521,N_20956);
and U21838 (N_21838,N_20490,N_20946);
nand U21839 (N_21839,N_20444,N_20126);
and U21840 (N_21840,N_20141,N_20226);
nor U21841 (N_21841,N_20394,N_20576);
xnor U21842 (N_21842,N_20323,N_20661);
xnor U21843 (N_21843,N_20829,N_20270);
and U21844 (N_21844,N_20862,N_20272);
or U21845 (N_21845,N_20315,N_20415);
nand U21846 (N_21846,N_20397,N_20382);
xor U21847 (N_21847,N_20791,N_20994);
nor U21848 (N_21848,N_20119,N_20472);
and U21849 (N_21849,N_20540,N_20854);
or U21850 (N_21850,N_20523,N_20155);
nor U21851 (N_21851,N_20770,N_20638);
xor U21852 (N_21852,N_20588,N_20913);
nor U21853 (N_21853,N_20654,N_20820);
or U21854 (N_21854,N_20858,N_20455);
nand U21855 (N_21855,N_20817,N_20556);
and U21856 (N_21856,N_20998,N_20155);
or U21857 (N_21857,N_20179,N_20552);
nor U21858 (N_21858,N_20600,N_20023);
and U21859 (N_21859,N_20906,N_20808);
nor U21860 (N_21860,N_20907,N_20560);
nand U21861 (N_21861,N_20740,N_20714);
nor U21862 (N_21862,N_20994,N_20288);
or U21863 (N_21863,N_20875,N_20752);
and U21864 (N_21864,N_20201,N_20033);
xor U21865 (N_21865,N_20413,N_20480);
and U21866 (N_21866,N_20086,N_20513);
xnor U21867 (N_21867,N_20135,N_20208);
and U21868 (N_21868,N_20812,N_20958);
and U21869 (N_21869,N_20433,N_20208);
xnor U21870 (N_21870,N_20094,N_20386);
or U21871 (N_21871,N_20968,N_20407);
and U21872 (N_21872,N_20661,N_20697);
nor U21873 (N_21873,N_20740,N_20722);
and U21874 (N_21874,N_20191,N_20938);
or U21875 (N_21875,N_20374,N_20249);
and U21876 (N_21876,N_20161,N_20213);
nand U21877 (N_21877,N_20621,N_20557);
xnor U21878 (N_21878,N_20879,N_20502);
xnor U21879 (N_21879,N_20709,N_20474);
or U21880 (N_21880,N_20235,N_20255);
nor U21881 (N_21881,N_20585,N_20731);
nand U21882 (N_21882,N_20390,N_20337);
xnor U21883 (N_21883,N_20580,N_20961);
nor U21884 (N_21884,N_20764,N_20285);
xnor U21885 (N_21885,N_20544,N_20018);
nand U21886 (N_21886,N_20009,N_20013);
nor U21887 (N_21887,N_20408,N_20635);
and U21888 (N_21888,N_20305,N_20030);
and U21889 (N_21889,N_20665,N_20187);
xnor U21890 (N_21890,N_20875,N_20463);
nand U21891 (N_21891,N_20823,N_20431);
nor U21892 (N_21892,N_20483,N_20971);
nand U21893 (N_21893,N_20293,N_20134);
and U21894 (N_21894,N_20934,N_20785);
or U21895 (N_21895,N_20501,N_20632);
xor U21896 (N_21896,N_20757,N_20790);
or U21897 (N_21897,N_20025,N_20657);
xnor U21898 (N_21898,N_20573,N_20691);
and U21899 (N_21899,N_20574,N_20437);
xnor U21900 (N_21900,N_20456,N_20187);
nor U21901 (N_21901,N_20923,N_20963);
and U21902 (N_21902,N_20656,N_20355);
or U21903 (N_21903,N_20699,N_20131);
and U21904 (N_21904,N_20264,N_20318);
nor U21905 (N_21905,N_20073,N_20617);
nand U21906 (N_21906,N_20657,N_20818);
xor U21907 (N_21907,N_20588,N_20586);
nand U21908 (N_21908,N_20112,N_20087);
or U21909 (N_21909,N_20793,N_20293);
or U21910 (N_21910,N_20570,N_20734);
and U21911 (N_21911,N_20622,N_20739);
nand U21912 (N_21912,N_20071,N_20548);
and U21913 (N_21913,N_20510,N_20616);
and U21914 (N_21914,N_20958,N_20015);
nor U21915 (N_21915,N_20955,N_20863);
or U21916 (N_21916,N_20278,N_20403);
nor U21917 (N_21917,N_20777,N_20320);
and U21918 (N_21918,N_20801,N_20010);
xnor U21919 (N_21919,N_20892,N_20349);
nand U21920 (N_21920,N_20838,N_20027);
xor U21921 (N_21921,N_20421,N_20409);
nand U21922 (N_21922,N_20888,N_20021);
xor U21923 (N_21923,N_20715,N_20767);
nor U21924 (N_21924,N_20830,N_20860);
and U21925 (N_21925,N_20352,N_20875);
nand U21926 (N_21926,N_20890,N_20394);
or U21927 (N_21927,N_20614,N_20374);
or U21928 (N_21928,N_20636,N_20980);
and U21929 (N_21929,N_20881,N_20867);
nand U21930 (N_21930,N_20230,N_20999);
nor U21931 (N_21931,N_20201,N_20447);
and U21932 (N_21932,N_20467,N_20918);
nor U21933 (N_21933,N_20236,N_20578);
nor U21934 (N_21934,N_20519,N_20550);
nand U21935 (N_21935,N_20296,N_20541);
and U21936 (N_21936,N_20064,N_20861);
xnor U21937 (N_21937,N_20144,N_20176);
and U21938 (N_21938,N_20434,N_20949);
nand U21939 (N_21939,N_20373,N_20469);
nor U21940 (N_21940,N_20312,N_20105);
nor U21941 (N_21941,N_20235,N_20419);
nand U21942 (N_21942,N_20406,N_20853);
nand U21943 (N_21943,N_20707,N_20678);
and U21944 (N_21944,N_20042,N_20689);
xor U21945 (N_21945,N_20528,N_20870);
or U21946 (N_21946,N_20296,N_20152);
or U21947 (N_21947,N_20460,N_20702);
nand U21948 (N_21948,N_20241,N_20848);
or U21949 (N_21949,N_20939,N_20773);
and U21950 (N_21950,N_20795,N_20805);
xnor U21951 (N_21951,N_20286,N_20146);
xnor U21952 (N_21952,N_20685,N_20557);
nor U21953 (N_21953,N_20425,N_20625);
nor U21954 (N_21954,N_20808,N_20545);
nor U21955 (N_21955,N_20849,N_20734);
nand U21956 (N_21956,N_20562,N_20929);
or U21957 (N_21957,N_20097,N_20896);
nor U21958 (N_21958,N_20368,N_20743);
or U21959 (N_21959,N_20967,N_20406);
or U21960 (N_21960,N_20096,N_20941);
xnor U21961 (N_21961,N_20852,N_20646);
and U21962 (N_21962,N_20363,N_20092);
and U21963 (N_21963,N_20326,N_20949);
nand U21964 (N_21964,N_20784,N_20034);
and U21965 (N_21965,N_20859,N_20511);
xnor U21966 (N_21966,N_20230,N_20272);
or U21967 (N_21967,N_20261,N_20410);
nor U21968 (N_21968,N_20680,N_20361);
xnor U21969 (N_21969,N_20017,N_20865);
xor U21970 (N_21970,N_20808,N_20987);
nand U21971 (N_21971,N_20849,N_20806);
nor U21972 (N_21972,N_20768,N_20547);
nor U21973 (N_21973,N_20654,N_20094);
and U21974 (N_21974,N_20915,N_20328);
or U21975 (N_21975,N_20724,N_20658);
nand U21976 (N_21976,N_20740,N_20348);
xnor U21977 (N_21977,N_20155,N_20234);
xor U21978 (N_21978,N_20281,N_20224);
nand U21979 (N_21979,N_20033,N_20839);
nor U21980 (N_21980,N_20690,N_20019);
or U21981 (N_21981,N_20648,N_20775);
xnor U21982 (N_21982,N_20586,N_20548);
nand U21983 (N_21983,N_20765,N_20532);
nor U21984 (N_21984,N_20909,N_20100);
or U21985 (N_21985,N_20234,N_20889);
nand U21986 (N_21986,N_20301,N_20965);
xnor U21987 (N_21987,N_20229,N_20029);
nor U21988 (N_21988,N_20318,N_20511);
xor U21989 (N_21989,N_20634,N_20742);
xor U21990 (N_21990,N_20314,N_20305);
or U21991 (N_21991,N_20839,N_20070);
xor U21992 (N_21992,N_20128,N_20282);
nor U21993 (N_21993,N_20793,N_20604);
nand U21994 (N_21994,N_20230,N_20195);
nand U21995 (N_21995,N_20643,N_20875);
or U21996 (N_21996,N_20243,N_20278);
xnor U21997 (N_21997,N_20382,N_20757);
or U21998 (N_21998,N_20944,N_20256);
nand U21999 (N_21999,N_20955,N_20658);
nor U22000 (N_22000,N_21316,N_21463);
and U22001 (N_22001,N_21657,N_21485);
xnor U22002 (N_22002,N_21214,N_21336);
or U22003 (N_22003,N_21756,N_21548);
and U22004 (N_22004,N_21389,N_21585);
nor U22005 (N_22005,N_21113,N_21326);
nor U22006 (N_22006,N_21294,N_21965);
nand U22007 (N_22007,N_21377,N_21735);
and U22008 (N_22008,N_21971,N_21388);
nand U22009 (N_22009,N_21524,N_21659);
nor U22010 (N_22010,N_21872,N_21790);
nand U22011 (N_22011,N_21644,N_21533);
or U22012 (N_22012,N_21291,N_21748);
nand U22013 (N_22013,N_21117,N_21525);
or U22014 (N_22014,N_21369,N_21039);
nor U22015 (N_22015,N_21399,N_21241);
xnor U22016 (N_22016,N_21408,N_21407);
or U22017 (N_22017,N_21036,N_21430);
and U22018 (N_22018,N_21034,N_21398);
xor U22019 (N_22019,N_21444,N_21484);
or U22020 (N_22020,N_21172,N_21370);
and U22021 (N_22021,N_21378,N_21826);
and U22022 (N_22022,N_21562,N_21539);
nand U22023 (N_22023,N_21312,N_21390);
and U22024 (N_22024,N_21675,N_21783);
or U22025 (N_22025,N_21052,N_21637);
or U22026 (N_22026,N_21220,N_21365);
xnor U22027 (N_22027,N_21605,N_21740);
or U22028 (N_22028,N_21357,N_21116);
and U22029 (N_22029,N_21344,N_21033);
and U22030 (N_22030,N_21082,N_21178);
nor U22031 (N_22031,N_21645,N_21292);
or U22032 (N_22032,N_21635,N_21986);
xor U22033 (N_22033,N_21202,N_21342);
and U22034 (N_22034,N_21274,N_21838);
or U22035 (N_22035,N_21909,N_21624);
and U22036 (N_22036,N_21273,N_21654);
or U22037 (N_22037,N_21295,N_21417);
xnor U22038 (N_22038,N_21574,N_21331);
nor U22039 (N_22039,N_21797,N_21360);
and U22040 (N_22040,N_21834,N_21696);
nor U22041 (N_22041,N_21560,N_21705);
and U22042 (N_22042,N_21785,N_21545);
xor U22043 (N_22043,N_21043,N_21306);
xor U22044 (N_22044,N_21961,N_21795);
or U22045 (N_22045,N_21698,N_21508);
or U22046 (N_22046,N_21411,N_21054);
or U22047 (N_22047,N_21459,N_21721);
or U22048 (N_22048,N_21104,N_21750);
nor U22049 (N_22049,N_21908,N_21249);
xnor U22050 (N_22050,N_21400,N_21019);
xnor U22051 (N_22051,N_21450,N_21824);
and U22052 (N_22052,N_21185,N_21121);
or U22053 (N_22053,N_21046,N_21325);
or U22054 (N_22054,N_21367,N_21672);
xnor U22055 (N_22055,N_21636,N_21324);
nand U22056 (N_22056,N_21849,N_21240);
nand U22057 (N_22057,N_21936,N_21772);
nor U22058 (N_22058,N_21296,N_21126);
or U22059 (N_22059,N_21979,N_21706);
nand U22060 (N_22060,N_21288,N_21681);
and U22061 (N_22061,N_21262,N_21171);
and U22062 (N_22062,N_21693,N_21014);
nand U22063 (N_22063,N_21017,N_21943);
nor U22064 (N_22064,N_21267,N_21075);
nand U22065 (N_22065,N_21487,N_21608);
xnor U22066 (N_22066,N_21649,N_21521);
nor U22067 (N_22067,N_21879,N_21155);
nor U22068 (N_22068,N_21841,N_21412);
nor U22069 (N_22069,N_21072,N_21372);
xor U22070 (N_22070,N_21232,N_21168);
nand U22071 (N_22071,N_21974,N_21467);
or U22072 (N_22072,N_21310,N_21596);
nor U22073 (N_22073,N_21527,N_21753);
nor U22074 (N_22074,N_21153,N_21800);
and U22075 (N_22075,N_21192,N_21875);
and U22076 (N_22076,N_21685,N_21130);
nand U22077 (N_22077,N_21090,N_21056);
xor U22078 (N_22078,N_21897,N_21106);
nand U22079 (N_22079,N_21453,N_21237);
and U22080 (N_22080,N_21458,N_21105);
nand U22081 (N_22081,N_21819,N_21405);
or U22082 (N_22082,N_21402,N_21499);
and U22083 (N_22083,N_21384,N_21958);
nand U22084 (N_22084,N_21020,N_21754);
and U22085 (N_22085,N_21991,N_21821);
xnor U22086 (N_22086,N_21855,N_21639);
xor U22087 (N_22087,N_21710,N_21012);
xnor U22088 (N_22088,N_21018,N_21536);
nand U22089 (N_22089,N_21253,N_21630);
xnor U22090 (N_22090,N_21766,N_21895);
nor U22091 (N_22091,N_21788,N_21469);
xor U22092 (N_22092,N_21422,N_21009);
nor U22093 (N_22093,N_21179,N_21787);
nor U22094 (N_22094,N_21601,N_21147);
nand U22095 (N_22095,N_21223,N_21462);
xor U22096 (N_22096,N_21751,N_21689);
and U22097 (N_22097,N_21794,N_21193);
nor U22098 (N_22098,N_21423,N_21994);
nor U22099 (N_22099,N_21940,N_21079);
nand U22100 (N_22100,N_21504,N_21057);
or U22101 (N_22101,N_21478,N_21626);
nor U22102 (N_22102,N_21953,N_21929);
or U22103 (N_22103,N_21629,N_21470);
nand U22104 (N_22104,N_21066,N_21268);
nand U22105 (N_22105,N_21133,N_21150);
or U22106 (N_22106,N_21815,N_21221);
or U22107 (N_22107,N_21436,N_21386);
and U22108 (N_22108,N_21161,N_21146);
xor U22109 (N_22109,N_21726,N_21903);
or U22110 (N_22110,N_21503,N_21498);
nor U22111 (N_22111,N_21523,N_21374);
or U22112 (N_22112,N_21990,N_21714);
nand U22113 (N_22113,N_21472,N_21317);
nor U22114 (N_22114,N_21617,N_21570);
or U22115 (N_22115,N_21233,N_21439);
and U22116 (N_22116,N_21140,N_21535);
nor U22117 (N_22117,N_21625,N_21230);
xor U22118 (N_22118,N_21989,N_21874);
xnor U22119 (N_22119,N_21746,N_21114);
nand U22120 (N_22120,N_21846,N_21736);
or U22121 (N_22121,N_21259,N_21102);
xnor U22122 (N_22122,N_21432,N_21631);
and U22123 (N_22123,N_21290,N_21087);
or U22124 (N_22124,N_21803,N_21951);
nand U22125 (N_22125,N_21277,N_21301);
and U22126 (N_22126,N_21900,N_21906);
and U22127 (N_22127,N_21712,N_21802);
xnor U22128 (N_22128,N_21600,N_21582);
nand U22129 (N_22129,N_21859,N_21798);
xor U22130 (N_22130,N_21435,N_21777);
and U22131 (N_22131,N_21424,N_21073);
nor U22132 (N_22132,N_21686,N_21473);
xor U22133 (N_22133,N_21238,N_21759);
nand U22134 (N_22134,N_21843,N_21078);
nor U22135 (N_22135,N_21169,N_21068);
xor U22136 (N_22136,N_21881,N_21889);
nand U22137 (N_22137,N_21392,N_21069);
nor U22138 (N_22138,N_21466,N_21032);
nand U22139 (N_22139,N_21722,N_21383);
nor U22140 (N_22140,N_21419,N_21611);
or U22141 (N_22141,N_21885,N_21825);
nand U22142 (N_22142,N_21853,N_21065);
xor U22143 (N_22143,N_21454,N_21373);
xnor U22144 (N_22144,N_21627,N_21856);
and U22145 (N_22145,N_21510,N_21250);
nor U22146 (N_22146,N_21127,N_21850);
nand U22147 (N_22147,N_21148,N_21460);
xnor U22148 (N_22148,N_21718,N_21599);
nand U22149 (N_22149,N_21186,N_21760);
or U22150 (N_22150,N_21304,N_21282);
xnor U22151 (N_22151,N_21298,N_21120);
nor U22152 (N_22152,N_21547,N_21932);
nand U22153 (N_22153,N_21406,N_21719);
nor U22154 (N_22154,N_21609,N_21684);
or U22155 (N_22155,N_21658,N_21898);
xor U22156 (N_22156,N_21835,N_21362);
or U22157 (N_22157,N_21403,N_21567);
xnor U22158 (N_22158,N_21299,N_21752);
nand U22159 (N_22159,N_21100,N_21715);
nor U22160 (N_22160,N_21334,N_21845);
nand U22161 (N_22161,N_21941,N_21784);
nand U22162 (N_22162,N_21865,N_21808);
nor U22163 (N_22163,N_21123,N_21468);
and U22164 (N_22164,N_21348,N_21028);
xnor U22165 (N_22165,N_21429,N_21180);
xor U22166 (N_22166,N_21176,N_21410);
nor U22167 (N_22167,N_21812,N_21966);
and U22168 (N_22168,N_21836,N_21345);
or U22169 (N_22169,N_21329,N_21190);
and U22170 (N_22170,N_21285,N_21578);
or U22171 (N_22171,N_21269,N_21888);
and U22172 (N_22172,N_21321,N_21199);
and U22173 (N_22173,N_21053,N_21287);
nor U22174 (N_22174,N_21051,N_21441);
nor U22175 (N_22175,N_21647,N_21911);
xor U22176 (N_22176,N_21242,N_21813);
and U22177 (N_22177,N_21944,N_21284);
or U22178 (N_22178,N_21025,N_21341);
and U22179 (N_22179,N_21902,N_21040);
xor U22180 (N_22180,N_21883,N_21666);
or U22181 (N_22181,N_21164,N_21747);
and U22182 (N_22182,N_21416,N_21828);
nand U22183 (N_22183,N_21045,N_21391);
or U22184 (N_22184,N_21692,N_21058);
or U22185 (N_22185,N_21505,N_21952);
xor U22186 (N_22186,N_21376,N_21912);
nor U22187 (N_22187,N_21584,N_21962);
xor U22188 (N_22188,N_21877,N_21077);
nor U22189 (N_22189,N_21985,N_21976);
or U22190 (N_22190,N_21244,N_21758);
nand U22191 (N_22191,N_21517,N_21091);
and U22192 (N_22192,N_21229,N_21713);
nand U22193 (N_22193,N_21049,N_21670);
or U22194 (N_22194,N_21420,N_21189);
nor U22195 (N_22195,N_21216,N_21160);
or U22196 (N_22196,N_21021,N_21923);
xor U22197 (N_22197,N_21425,N_21254);
nor U22198 (N_22198,N_21447,N_21081);
xnor U22199 (N_22199,N_21501,N_21543);
xnor U22200 (N_22200,N_21925,N_21776);
xor U22201 (N_22201,N_21955,N_21279);
or U22202 (N_22202,N_21101,N_21676);
or U22203 (N_22203,N_21683,N_21768);
and U22204 (N_22204,N_21699,N_21822);
nor U22205 (N_22205,N_21210,N_21837);
nor U22206 (N_22206,N_21327,N_21571);
xnor U22207 (N_22207,N_21007,N_21455);
xnor U22208 (N_22208,N_21380,N_21805);
and U22209 (N_22209,N_21694,N_21509);
nand U22210 (N_22210,N_21188,N_21948);
nand U22211 (N_22211,N_21476,N_21661);
xnor U22212 (N_22212,N_21048,N_21479);
or U22213 (N_22213,N_21482,N_21993);
or U22214 (N_22214,N_21174,N_21709);
nor U22215 (N_22215,N_21055,N_21745);
nand U22216 (N_22216,N_21302,N_21083);
and U22217 (N_22217,N_21443,N_21983);
nor U22218 (N_22218,N_21332,N_21440);
or U22219 (N_22219,N_21208,N_21303);
or U22220 (N_22220,N_21395,N_21265);
nor U22221 (N_22221,N_21764,N_21024);
nor U22222 (N_22222,N_21842,N_21434);
or U22223 (N_22223,N_21810,N_21518);
and U22224 (N_22224,N_21433,N_21177);
nand U22225 (N_22225,N_21729,N_21089);
nand U22226 (N_22226,N_21592,N_21531);
nand U22227 (N_22227,N_21149,N_21212);
and U22228 (N_22228,N_21500,N_21491);
or U22229 (N_22229,N_21309,N_21001);
and U22230 (N_22230,N_21204,N_21774);
xor U22231 (N_22231,N_21278,N_21763);
and U22232 (N_22232,N_21137,N_21931);
nor U22233 (N_22233,N_21643,N_21583);
xnor U22234 (N_22234,N_21196,N_21623);
or U22235 (N_22235,N_21339,N_21158);
nand U22236 (N_22236,N_21218,N_21839);
nor U22237 (N_22237,N_21280,N_21243);
nand U22238 (N_22238,N_21998,N_21157);
nand U22239 (N_22239,N_21896,N_21311);
nand U22240 (N_22240,N_21234,N_21445);
and U22241 (N_22241,N_21136,N_21431);
nor U22242 (N_22242,N_21641,N_21067);
and U22243 (N_22243,N_21970,N_21323);
nand U22244 (N_22244,N_21401,N_21580);
and U22245 (N_22245,N_21222,N_21559);
nor U22246 (N_22246,N_21938,N_21110);
or U22247 (N_22247,N_21610,N_21115);
or U22248 (N_22248,N_21356,N_21663);
xnor U22249 (N_22249,N_21621,N_21328);
nand U22250 (N_22250,N_21118,N_21595);
nor U22251 (N_22251,N_21270,N_21546);
or U22252 (N_22252,N_21465,N_21381);
xor U22253 (N_22253,N_21063,N_21135);
nand U22254 (N_22254,N_21042,N_21236);
nor U22255 (N_22255,N_21086,N_21483);
and U22256 (N_22256,N_21716,N_21907);
or U22257 (N_22257,N_21071,N_21702);
or U22258 (N_22258,N_21198,N_21502);
or U22259 (N_22259,N_21779,N_21248);
and U22260 (N_22260,N_21044,N_21612);
xnor U22261 (N_22261,N_21870,N_21530);
nand U22262 (N_22262,N_21963,N_21191);
xnor U22263 (N_22263,N_21343,N_21004);
and U22264 (N_22264,N_21495,N_21840);
nor U22265 (N_22265,N_21552,N_21996);
nor U22266 (N_22266,N_21194,N_21833);
or U22267 (N_22267,N_21697,N_21029);
nand U22268 (N_22268,N_21142,N_21568);
or U22269 (N_22269,N_21939,N_21588);
nor U22270 (N_22270,N_21921,N_21603);
nor U22271 (N_22271,N_21041,N_21480);
or U22272 (N_22272,N_21008,N_21184);
nand U22273 (N_22273,N_21464,N_21335);
nor U22274 (N_22274,N_21563,N_21512);
or U22275 (N_22275,N_21969,N_21717);
nand U22276 (N_22276,N_21662,N_21516);
nor U22277 (N_22277,N_21978,N_21181);
or U22278 (N_22278,N_21919,N_21217);
and U22279 (N_22279,N_21477,N_21964);
xor U22280 (N_22280,N_21030,N_21809);
and U22281 (N_22281,N_21848,N_21129);
nand U22282 (N_22282,N_21108,N_21806);
and U22283 (N_22283,N_21461,N_21572);
or U22284 (N_22284,N_21260,N_21844);
nand U22285 (N_22285,N_21475,N_21213);
xnor U22286 (N_22286,N_21337,N_21154);
nand U22287 (N_22287,N_21182,N_21308);
nor U22288 (N_22288,N_21554,N_21598);
xor U22289 (N_22289,N_21700,N_21725);
nand U22290 (N_22290,N_21526,N_21375);
and U22291 (N_22291,N_21438,N_21225);
and U22292 (N_22292,N_21830,N_21928);
or U22293 (N_22293,N_21566,N_21781);
nand U22294 (N_22294,N_21674,N_21305);
xnor U22295 (N_22295,N_21607,N_21946);
xnor U22296 (N_22296,N_21255,N_21338);
xor U22297 (N_22297,N_21997,N_21935);
or U22298 (N_22298,N_21999,N_21371);
nand U22299 (N_22299,N_21442,N_21141);
or U22300 (N_22300,N_21786,N_21387);
nor U22301 (N_22301,N_21728,N_21910);
or U22302 (N_22302,N_21869,N_21289);
nor U22303 (N_22303,N_21061,N_21924);
xor U22304 (N_22304,N_21251,N_21557);
xor U22305 (N_22305,N_21780,N_21980);
xnor U22306 (N_22306,N_21358,N_21680);
or U22307 (N_22307,N_21823,N_21755);
xor U22308 (N_22308,N_21871,N_21576);
xnor U22309 (N_22309,N_21891,N_21593);
xnor U22310 (N_22310,N_21734,N_21037);
and U22311 (N_22311,N_21205,N_21333);
xor U22312 (N_22312,N_21981,N_21927);
nor U22313 (N_22313,N_21085,N_21209);
nand U22314 (N_22314,N_21606,N_21655);
xnor U22315 (N_22315,N_21227,N_21651);
or U22316 (N_22316,N_21937,N_21144);
nand U22317 (N_22317,N_21861,N_21586);
or U22318 (N_22318,N_21541,N_21668);
or U22319 (N_22319,N_21047,N_21741);
xor U22320 (N_22320,N_21984,N_21271);
and U22321 (N_22321,N_21064,N_21514);
nand U22322 (N_22322,N_21421,N_21995);
nor U22323 (N_22323,N_21264,N_21669);
nor U22324 (N_22324,N_21540,N_21132);
nand U22325 (N_22325,N_21281,N_21261);
nand U22326 (N_22326,N_21368,N_21197);
nor U22327 (N_22327,N_21544,N_21350);
nor U22328 (N_22328,N_21211,N_21972);
and U22329 (N_22329,N_21860,N_21930);
nor U22330 (N_22330,N_21070,N_21183);
nor U22331 (N_22331,N_21415,N_21307);
xor U22332 (N_22332,N_21364,N_21553);
nor U22333 (N_22333,N_21515,N_21899);
or U22334 (N_22334,N_21796,N_21537);
nor U22335 (N_22335,N_21762,N_21076);
xnor U22336 (N_22336,N_21330,N_21143);
nand U22337 (N_22337,N_21867,N_21616);
nor U22338 (N_22338,N_21773,N_21492);
and U22339 (N_22339,N_21200,N_21497);
or U22340 (N_22340,N_21131,N_21414);
or U22341 (N_22341,N_21743,N_21322);
and U22342 (N_22342,N_21538,N_21876);
nand U22343 (N_22343,N_21708,N_21002);
xnor U22344 (N_22344,N_21170,N_21506);
and U22345 (N_22345,N_21992,N_21128);
nor U22346 (N_22346,N_21084,N_21088);
and U22347 (N_22347,N_21707,N_21000);
and U22348 (N_22348,N_21765,N_21818);
or U22349 (N_22349,N_21577,N_21949);
nor U22350 (N_22350,N_21532,N_21166);
and U22351 (N_22351,N_21319,N_21013);
or U22352 (N_22352,N_21950,N_21581);
or U22353 (N_22353,N_21203,N_21226);
xor U22354 (N_22354,N_21093,N_21062);
nand U22355 (N_22355,N_21245,N_21152);
nor U22356 (N_22356,N_21878,N_21379);
and U22357 (N_22357,N_21125,N_21832);
xnor U22358 (N_22358,N_21614,N_21456);
and U22359 (N_22359,N_21915,N_21315);
nor U22360 (N_22360,N_21493,N_21711);
and U22361 (N_22361,N_21022,N_21829);
nor U22362 (N_22362,N_21382,N_21235);
nor U22363 (N_22363,N_21446,N_21122);
nor U22364 (N_22364,N_21761,N_21393);
and U22365 (N_22365,N_21224,N_21988);
or U22366 (N_22366,N_21096,N_21397);
or U22367 (N_22367,N_21723,N_21792);
and U22368 (N_22368,N_21917,N_21778);
xnor U22369 (N_22369,N_21945,N_21258);
nand U22370 (N_22370,N_21320,N_21664);
or U22371 (N_22371,N_21507,N_21489);
xor U22372 (N_22372,N_21868,N_21542);
nand U22373 (N_22373,N_21366,N_21124);
or U22374 (N_22374,N_21886,N_21451);
or U22375 (N_22375,N_21276,N_21769);
xnor U22376 (N_22376,N_21488,N_21050);
nor U22377 (N_22377,N_21145,N_21591);
nor U22378 (N_22378,N_21256,N_21638);
and U22379 (N_22379,N_21863,N_21318);
nor U22380 (N_22380,N_21968,N_21272);
and U22381 (N_22381,N_21413,N_21920);
and U22382 (N_22382,N_21092,N_21820);
nor U22383 (N_22383,N_21804,N_21257);
nor U22384 (N_22384,N_21660,N_21977);
nor U22385 (N_22385,N_21854,N_21165);
nand U22386 (N_22386,N_21656,N_21799);
nor U22387 (N_22387,N_21916,N_21426);
and U22388 (N_22388,N_21252,N_21791);
nor U22389 (N_22389,N_21471,N_21494);
xor U22390 (N_22390,N_21982,N_21687);
xor U22391 (N_22391,N_21733,N_21112);
or U22392 (N_22392,N_21757,N_21703);
nand U22393 (N_22393,N_21195,N_21026);
nor U22394 (N_22394,N_21187,N_21887);
nor U22395 (N_22395,N_21107,N_21967);
and U22396 (N_22396,N_21678,N_21619);
nor U22397 (N_22397,N_21520,N_21807);
nand U22398 (N_22398,N_21904,N_21486);
and U22399 (N_22399,N_21219,N_21695);
xnor U22400 (N_22400,N_21138,N_21015);
and U22401 (N_22401,N_21060,N_21633);
nor U22402 (N_22402,N_21720,N_21094);
or U22403 (N_22403,N_21097,N_21167);
nor U22404 (N_22404,N_21119,N_21427);
and U22405 (N_22405,N_21103,N_21847);
nand U22406 (N_22406,N_21628,N_21960);
nor U22407 (N_22407,N_21266,N_21111);
nor U22408 (N_22408,N_21139,N_21038);
xnor U22409 (N_22409,N_21355,N_21031);
nor U22410 (N_22410,N_21852,N_21749);
or U22411 (N_22411,N_21549,N_21851);
nor U22412 (N_22412,N_21648,N_21173);
nor U22413 (N_22413,N_21347,N_21573);
and U22414 (N_22414,N_21359,N_21589);
nand U22415 (N_22415,N_21396,N_21739);
nor U22416 (N_22416,N_21613,N_21690);
xor U22417 (N_22417,N_21490,N_21016);
nand U22418 (N_22418,N_21363,N_21206);
or U22419 (N_22419,N_21511,N_21594);
or U22420 (N_22420,N_21522,N_21297);
nor U22421 (N_22421,N_21575,N_21394);
nand U22422 (N_22422,N_21679,N_21474);
and U22423 (N_22423,N_21098,N_21449);
nand U22424 (N_22424,N_21620,N_21457);
nand U22425 (N_22425,N_21286,N_21528);
nor U22426 (N_22426,N_21163,N_21957);
nand U22427 (N_22427,N_21864,N_21564);
or U22428 (N_22428,N_21561,N_21095);
nand U22429 (N_22429,N_21003,N_21565);
and U22430 (N_22430,N_21361,N_21215);
xor U22431 (N_22431,N_21727,N_21622);
nor U22432 (N_22432,N_21775,N_21156);
nor U22433 (N_22433,N_21738,N_21558);
or U22434 (N_22434,N_21602,N_21691);
xnor U22435 (N_22435,N_21956,N_21882);
and U22436 (N_22436,N_21134,N_21035);
nor U22437 (N_22437,N_21933,N_21671);
nor U22438 (N_22438,N_21201,N_21080);
or U22439 (N_22439,N_21247,N_21811);
xnor U22440 (N_22440,N_21448,N_21529);
and U22441 (N_22441,N_21918,N_21099);
nor U22442 (N_22442,N_21634,N_21892);
or U22443 (N_22443,N_21346,N_21615);
xor U22444 (N_22444,N_21858,N_21894);
and U22445 (N_22445,N_21428,N_21831);
nor U22446 (N_22446,N_21228,N_21349);
nand U22447 (N_22447,N_21263,N_21246);
xor U22448 (N_22448,N_21737,N_21437);
nand U22449 (N_22449,N_21677,N_21814);
nand U22450 (N_22450,N_21481,N_21640);
nor U22451 (N_22451,N_21513,N_21519);
nand U22452 (N_22452,N_21947,N_21731);
and U22453 (N_22453,N_21959,N_21642);
nor U22454 (N_22454,N_21352,N_21159);
nand U22455 (N_22455,N_21632,N_21275);
nand U22456 (N_22456,N_21353,N_21880);
xor U22457 (N_22457,N_21385,N_21354);
nor U22458 (N_22458,N_21742,N_21816);
or U22459 (N_22459,N_21732,N_21618);
nand U22460 (N_22460,N_21801,N_21300);
or U22461 (N_22461,N_21109,N_21162);
and U22462 (N_22462,N_21688,N_21597);
nand U22463 (N_22463,N_21817,N_21730);
xor U22464 (N_22464,N_21239,N_21027);
nor U22465 (N_22465,N_21665,N_21351);
or U22466 (N_22466,N_21496,N_21231);
or U22467 (N_22467,N_21418,N_21023);
and U22468 (N_22468,N_21866,N_21975);
xnor U22469 (N_22469,N_21207,N_21770);
and U22470 (N_22470,N_21793,N_21059);
and U22471 (N_22471,N_21452,N_21650);
and U22472 (N_22472,N_21827,N_21873);
nor U22473 (N_22473,N_21652,N_21011);
nor U22474 (N_22474,N_21901,N_21550);
nand U22475 (N_22475,N_21005,N_21724);
or U22476 (N_22476,N_21175,N_21587);
and U22477 (N_22477,N_21914,N_21590);
and U22478 (N_22478,N_21074,N_21922);
and U22479 (N_22479,N_21667,N_21926);
or U22480 (N_22480,N_21555,N_21704);
nand U22481 (N_22481,N_21556,N_21942);
nor U22482 (N_22482,N_21404,N_21913);
nand U22483 (N_22483,N_21782,N_21789);
and U22484 (N_22484,N_21771,N_21744);
nand U22485 (N_22485,N_21151,N_21569);
xor U22486 (N_22486,N_21283,N_21973);
nor U22487 (N_22487,N_21767,N_21884);
nand U22488 (N_22488,N_21890,N_21987);
xnor U22489 (N_22489,N_21409,N_21314);
and U22490 (N_22490,N_21673,N_21905);
and U22491 (N_22491,N_21340,N_21646);
or U22492 (N_22492,N_21313,N_21293);
and U22493 (N_22493,N_21701,N_21862);
and U22494 (N_22494,N_21579,N_21682);
xor U22495 (N_22495,N_21653,N_21006);
nor U22496 (N_22496,N_21934,N_21010);
nor U22497 (N_22497,N_21551,N_21604);
xor U22498 (N_22498,N_21534,N_21857);
nand U22499 (N_22499,N_21893,N_21954);
nor U22500 (N_22500,N_21249,N_21738);
xor U22501 (N_22501,N_21072,N_21181);
and U22502 (N_22502,N_21247,N_21482);
or U22503 (N_22503,N_21090,N_21208);
nor U22504 (N_22504,N_21441,N_21285);
nor U22505 (N_22505,N_21180,N_21465);
xor U22506 (N_22506,N_21069,N_21432);
or U22507 (N_22507,N_21948,N_21434);
nand U22508 (N_22508,N_21032,N_21146);
or U22509 (N_22509,N_21837,N_21198);
xor U22510 (N_22510,N_21453,N_21545);
xor U22511 (N_22511,N_21664,N_21771);
nor U22512 (N_22512,N_21184,N_21404);
nand U22513 (N_22513,N_21235,N_21987);
nor U22514 (N_22514,N_21115,N_21320);
nor U22515 (N_22515,N_21504,N_21054);
xnor U22516 (N_22516,N_21899,N_21838);
nand U22517 (N_22517,N_21507,N_21404);
xor U22518 (N_22518,N_21045,N_21971);
nand U22519 (N_22519,N_21636,N_21551);
nand U22520 (N_22520,N_21222,N_21280);
and U22521 (N_22521,N_21175,N_21929);
and U22522 (N_22522,N_21162,N_21834);
xnor U22523 (N_22523,N_21328,N_21616);
and U22524 (N_22524,N_21669,N_21307);
or U22525 (N_22525,N_21250,N_21641);
nor U22526 (N_22526,N_21614,N_21732);
nor U22527 (N_22527,N_21593,N_21197);
xor U22528 (N_22528,N_21245,N_21623);
and U22529 (N_22529,N_21029,N_21284);
nor U22530 (N_22530,N_21960,N_21063);
and U22531 (N_22531,N_21315,N_21295);
nand U22532 (N_22532,N_21474,N_21693);
nor U22533 (N_22533,N_21609,N_21871);
nor U22534 (N_22534,N_21907,N_21689);
or U22535 (N_22535,N_21557,N_21551);
or U22536 (N_22536,N_21986,N_21630);
or U22537 (N_22537,N_21998,N_21230);
nor U22538 (N_22538,N_21305,N_21306);
nor U22539 (N_22539,N_21444,N_21297);
nor U22540 (N_22540,N_21541,N_21255);
and U22541 (N_22541,N_21123,N_21219);
or U22542 (N_22542,N_21687,N_21729);
xor U22543 (N_22543,N_21039,N_21488);
nand U22544 (N_22544,N_21038,N_21551);
nand U22545 (N_22545,N_21771,N_21750);
or U22546 (N_22546,N_21021,N_21942);
and U22547 (N_22547,N_21984,N_21942);
and U22548 (N_22548,N_21648,N_21646);
nand U22549 (N_22549,N_21944,N_21723);
xor U22550 (N_22550,N_21403,N_21673);
nand U22551 (N_22551,N_21528,N_21479);
nand U22552 (N_22552,N_21657,N_21574);
and U22553 (N_22553,N_21115,N_21290);
xor U22554 (N_22554,N_21128,N_21036);
nor U22555 (N_22555,N_21722,N_21275);
and U22556 (N_22556,N_21481,N_21120);
and U22557 (N_22557,N_21011,N_21259);
and U22558 (N_22558,N_21990,N_21962);
xnor U22559 (N_22559,N_21331,N_21611);
nand U22560 (N_22560,N_21973,N_21964);
nor U22561 (N_22561,N_21529,N_21344);
nand U22562 (N_22562,N_21633,N_21294);
nor U22563 (N_22563,N_21822,N_21926);
xor U22564 (N_22564,N_21620,N_21847);
or U22565 (N_22565,N_21035,N_21211);
or U22566 (N_22566,N_21265,N_21282);
nand U22567 (N_22567,N_21449,N_21110);
or U22568 (N_22568,N_21857,N_21353);
nand U22569 (N_22569,N_21689,N_21587);
nor U22570 (N_22570,N_21976,N_21021);
nand U22571 (N_22571,N_21614,N_21985);
nor U22572 (N_22572,N_21798,N_21074);
or U22573 (N_22573,N_21133,N_21812);
or U22574 (N_22574,N_21096,N_21004);
nand U22575 (N_22575,N_21750,N_21274);
nor U22576 (N_22576,N_21877,N_21725);
nand U22577 (N_22577,N_21084,N_21066);
or U22578 (N_22578,N_21762,N_21459);
xnor U22579 (N_22579,N_21572,N_21600);
or U22580 (N_22580,N_21469,N_21246);
or U22581 (N_22581,N_21492,N_21899);
nor U22582 (N_22582,N_21813,N_21051);
or U22583 (N_22583,N_21287,N_21979);
or U22584 (N_22584,N_21325,N_21850);
nand U22585 (N_22585,N_21289,N_21058);
and U22586 (N_22586,N_21350,N_21343);
nand U22587 (N_22587,N_21194,N_21758);
and U22588 (N_22588,N_21141,N_21560);
and U22589 (N_22589,N_21965,N_21178);
nand U22590 (N_22590,N_21621,N_21313);
and U22591 (N_22591,N_21864,N_21593);
or U22592 (N_22592,N_21504,N_21038);
nand U22593 (N_22593,N_21285,N_21922);
and U22594 (N_22594,N_21976,N_21811);
nor U22595 (N_22595,N_21984,N_21669);
nor U22596 (N_22596,N_21112,N_21006);
or U22597 (N_22597,N_21888,N_21610);
nand U22598 (N_22598,N_21748,N_21716);
xnor U22599 (N_22599,N_21085,N_21718);
or U22600 (N_22600,N_21005,N_21460);
nand U22601 (N_22601,N_21108,N_21218);
nand U22602 (N_22602,N_21868,N_21855);
xor U22603 (N_22603,N_21700,N_21996);
xor U22604 (N_22604,N_21924,N_21600);
and U22605 (N_22605,N_21204,N_21437);
xnor U22606 (N_22606,N_21514,N_21319);
xnor U22607 (N_22607,N_21642,N_21975);
xnor U22608 (N_22608,N_21187,N_21808);
nand U22609 (N_22609,N_21408,N_21888);
nand U22610 (N_22610,N_21760,N_21722);
or U22611 (N_22611,N_21978,N_21440);
nand U22612 (N_22612,N_21599,N_21963);
and U22613 (N_22613,N_21772,N_21579);
nor U22614 (N_22614,N_21756,N_21456);
nor U22615 (N_22615,N_21992,N_21687);
xor U22616 (N_22616,N_21425,N_21307);
and U22617 (N_22617,N_21026,N_21778);
and U22618 (N_22618,N_21570,N_21620);
or U22619 (N_22619,N_21296,N_21270);
xor U22620 (N_22620,N_21142,N_21124);
nor U22621 (N_22621,N_21726,N_21378);
nor U22622 (N_22622,N_21224,N_21426);
nor U22623 (N_22623,N_21153,N_21240);
or U22624 (N_22624,N_21129,N_21698);
and U22625 (N_22625,N_21040,N_21165);
xnor U22626 (N_22626,N_21164,N_21099);
or U22627 (N_22627,N_21247,N_21916);
nor U22628 (N_22628,N_21307,N_21846);
xor U22629 (N_22629,N_21128,N_21202);
nor U22630 (N_22630,N_21649,N_21946);
or U22631 (N_22631,N_21444,N_21146);
or U22632 (N_22632,N_21785,N_21542);
nor U22633 (N_22633,N_21270,N_21688);
and U22634 (N_22634,N_21392,N_21481);
xnor U22635 (N_22635,N_21567,N_21952);
nand U22636 (N_22636,N_21929,N_21669);
nor U22637 (N_22637,N_21151,N_21717);
nand U22638 (N_22638,N_21929,N_21654);
and U22639 (N_22639,N_21760,N_21288);
or U22640 (N_22640,N_21984,N_21030);
nor U22641 (N_22641,N_21893,N_21913);
nand U22642 (N_22642,N_21258,N_21829);
nor U22643 (N_22643,N_21895,N_21984);
nor U22644 (N_22644,N_21823,N_21948);
and U22645 (N_22645,N_21947,N_21369);
nor U22646 (N_22646,N_21176,N_21773);
xnor U22647 (N_22647,N_21478,N_21471);
xnor U22648 (N_22648,N_21580,N_21747);
xnor U22649 (N_22649,N_21563,N_21660);
or U22650 (N_22650,N_21840,N_21505);
nor U22651 (N_22651,N_21083,N_21783);
xor U22652 (N_22652,N_21947,N_21280);
xnor U22653 (N_22653,N_21215,N_21466);
and U22654 (N_22654,N_21140,N_21564);
nand U22655 (N_22655,N_21536,N_21027);
or U22656 (N_22656,N_21283,N_21072);
nor U22657 (N_22657,N_21771,N_21898);
nor U22658 (N_22658,N_21176,N_21156);
or U22659 (N_22659,N_21293,N_21307);
or U22660 (N_22660,N_21461,N_21318);
or U22661 (N_22661,N_21952,N_21346);
nand U22662 (N_22662,N_21210,N_21694);
and U22663 (N_22663,N_21917,N_21452);
or U22664 (N_22664,N_21566,N_21759);
nor U22665 (N_22665,N_21938,N_21678);
nand U22666 (N_22666,N_21175,N_21297);
or U22667 (N_22667,N_21603,N_21650);
xnor U22668 (N_22668,N_21082,N_21138);
nor U22669 (N_22669,N_21182,N_21546);
nand U22670 (N_22670,N_21437,N_21863);
xnor U22671 (N_22671,N_21756,N_21741);
xor U22672 (N_22672,N_21138,N_21915);
nor U22673 (N_22673,N_21464,N_21835);
and U22674 (N_22674,N_21133,N_21126);
or U22675 (N_22675,N_21789,N_21921);
nand U22676 (N_22676,N_21547,N_21702);
xnor U22677 (N_22677,N_21988,N_21586);
nor U22678 (N_22678,N_21179,N_21644);
xnor U22679 (N_22679,N_21885,N_21732);
nor U22680 (N_22680,N_21064,N_21508);
nand U22681 (N_22681,N_21303,N_21943);
or U22682 (N_22682,N_21280,N_21905);
nor U22683 (N_22683,N_21015,N_21228);
or U22684 (N_22684,N_21736,N_21901);
nand U22685 (N_22685,N_21309,N_21189);
nor U22686 (N_22686,N_21126,N_21861);
nand U22687 (N_22687,N_21559,N_21626);
and U22688 (N_22688,N_21014,N_21732);
nand U22689 (N_22689,N_21000,N_21369);
and U22690 (N_22690,N_21480,N_21003);
nor U22691 (N_22691,N_21030,N_21104);
or U22692 (N_22692,N_21159,N_21388);
and U22693 (N_22693,N_21870,N_21188);
nand U22694 (N_22694,N_21501,N_21549);
nand U22695 (N_22695,N_21767,N_21582);
xnor U22696 (N_22696,N_21912,N_21438);
xor U22697 (N_22697,N_21080,N_21301);
and U22698 (N_22698,N_21470,N_21023);
and U22699 (N_22699,N_21442,N_21764);
and U22700 (N_22700,N_21843,N_21233);
nor U22701 (N_22701,N_21211,N_21721);
or U22702 (N_22702,N_21957,N_21785);
nor U22703 (N_22703,N_21082,N_21539);
nand U22704 (N_22704,N_21724,N_21900);
nand U22705 (N_22705,N_21892,N_21331);
xnor U22706 (N_22706,N_21906,N_21625);
nand U22707 (N_22707,N_21510,N_21829);
and U22708 (N_22708,N_21093,N_21022);
nor U22709 (N_22709,N_21509,N_21695);
nand U22710 (N_22710,N_21029,N_21592);
nor U22711 (N_22711,N_21746,N_21686);
nor U22712 (N_22712,N_21570,N_21186);
and U22713 (N_22713,N_21924,N_21381);
or U22714 (N_22714,N_21222,N_21453);
nand U22715 (N_22715,N_21969,N_21744);
and U22716 (N_22716,N_21806,N_21606);
nor U22717 (N_22717,N_21318,N_21449);
or U22718 (N_22718,N_21403,N_21078);
nor U22719 (N_22719,N_21270,N_21710);
nor U22720 (N_22720,N_21447,N_21411);
nand U22721 (N_22721,N_21368,N_21628);
or U22722 (N_22722,N_21772,N_21658);
and U22723 (N_22723,N_21245,N_21827);
nand U22724 (N_22724,N_21982,N_21761);
xor U22725 (N_22725,N_21491,N_21928);
and U22726 (N_22726,N_21610,N_21742);
nand U22727 (N_22727,N_21702,N_21208);
and U22728 (N_22728,N_21021,N_21316);
nand U22729 (N_22729,N_21489,N_21733);
or U22730 (N_22730,N_21095,N_21357);
or U22731 (N_22731,N_21001,N_21418);
nor U22732 (N_22732,N_21680,N_21246);
or U22733 (N_22733,N_21611,N_21297);
xnor U22734 (N_22734,N_21345,N_21539);
nand U22735 (N_22735,N_21656,N_21300);
or U22736 (N_22736,N_21249,N_21286);
xor U22737 (N_22737,N_21529,N_21943);
or U22738 (N_22738,N_21977,N_21142);
xnor U22739 (N_22739,N_21064,N_21125);
xor U22740 (N_22740,N_21085,N_21997);
nand U22741 (N_22741,N_21333,N_21381);
xor U22742 (N_22742,N_21936,N_21078);
nand U22743 (N_22743,N_21472,N_21345);
or U22744 (N_22744,N_21114,N_21509);
xnor U22745 (N_22745,N_21146,N_21838);
and U22746 (N_22746,N_21152,N_21128);
and U22747 (N_22747,N_21976,N_21897);
or U22748 (N_22748,N_21931,N_21645);
and U22749 (N_22749,N_21518,N_21755);
and U22750 (N_22750,N_21894,N_21049);
nor U22751 (N_22751,N_21381,N_21115);
nor U22752 (N_22752,N_21078,N_21074);
nor U22753 (N_22753,N_21063,N_21446);
nand U22754 (N_22754,N_21498,N_21829);
or U22755 (N_22755,N_21186,N_21823);
or U22756 (N_22756,N_21516,N_21349);
or U22757 (N_22757,N_21322,N_21633);
nand U22758 (N_22758,N_21229,N_21775);
xnor U22759 (N_22759,N_21610,N_21205);
nor U22760 (N_22760,N_21699,N_21266);
and U22761 (N_22761,N_21848,N_21280);
nand U22762 (N_22762,N_21236,N_21963);
xnor U22763 (N_22763,N_21997,N_21516);
nor U22764 (N_22764,N_21009,N_21703);
nand U22765 (N_22765,N_21329,N_21467);
xnor U22766 (N_22766,N_21815,N_21235);
or U22767 (N_22767,N_21506,N_21754);
or U22768 (N_22768,N_21853,N_21546);
xor U22769 (N_22769,N_21284,N_21700);
nand U22770 (N_22770,N_21664,N_21869);
or U22771 (N_22771,N_21235,N_21206);
nor U22772 (N_22772,N_21456,N_21398);
xnor U22773 (N_22773,N_21097,N_21627);
xnor U22774 (N_22774,N_21673,N_21379);
and U22775 (N_22775,N_21990,N_21694);
nor U22776 (N_22776,N_21336,N_21911);
and U22777 (N_22777,N_21550,N_21545);
or U22778 (N_22778,N_21649,N_21296);
xnor U22779 (N_22779,N_21930,N_21471);
or U22780 (N_22780,N_21217,N_21834);
nand U22781 (N_22781,N_21561,N_21748);
or U22782 (N_22782,N_21997,N_21431);
or U22783 (N_22783,N_21812,N_21266);
nand U22784 (N_22784,N_21645,N_21755);
or U22785 (N_22785,N_21262,N_21911);
or U22786 (N_22786,N_21466,N_21864);
or U22787 (N_22787,N_21819,N_21121);
or U22788 (N_22788,N_21865,N_21791);
xnor U22789 (N_22789,N_21287,N_21921);
nor U22790 (N_22790,N_21563,N_21189);
or U22791 (N_22791,N_21857,N_21784);
nor U22792 (N_22792,N_21401,N_21002);
nand U22793 (N_22793,N_21263,N_21645);
and U22794 (N_22794,N_21503,N_21795);
and U22795 (N_22795,N_21267,N_21534);
or U22796 (N_22796,N_21276,N_21059);
or U22797 (N_22797,N_21562,N_21510);
nand U22798 (N_22798,N_21130,N_21675);
or U22799 (N_22799,N_21646,N_21914);
and U22800 (N_22800,N_21374,N_21133);
xor U22801 (N_22801,N_21033,N_21592);
xnor U22802 (N_22802,N_21937,N_21129);
or U22803 (N_22803,N_21039,N_21071);
nand U22804 (N_22804,N_21185,N_21753);
or U22805 (N_22805,N_21582,N_21652);
or U22806 (N_22806,N_21864,N_21356);
nand U22807 (N_22807,N_21678,N_21816);
and U22808 (N_22808,N_21047,N_21842);
nor U22809 (N_22809,N_21230,N_21402);
or U22810 (N_22810,N_21869,N_21754);
xnor U22811 (N_22811,N_21766,N_21564);
nor U22812 (N_22812,N_21384,N_21754);
and U22813 (N_22813,N_21891,N_21637);
and U22814 (N_22814,N_21810,N_21450);
and U22815 (N_22815,N_21087,N_21644);
xnor U22816 (N_22816,N_21671,N_21382);
xor U22817 (N_22817,N_21611,N_21566);
and U22818 (N_22818,N_21701,N_21585);
xor U22819 (N_22819,N_21365,N_21670);
xor U22820 (N_22820,N_21332,N_21486);
nand U22821 (N_22821,N_21857,N_21333);
or U22822 (N_22822,N_21378,N_21419);
nand U22823 (N_22823,N_21860,N_21079);
nor U22824 (N_22824,N_21740,N_21492);
and U22825 (N_22825,N_21451,N_21782);
nand U22826 (N_22826,N_21730,N_21560);
and U22827 (N_22827,N_21170,N_21519);
xnor U22828 (N_22828,N_21246,N_21772);
xnor U22829 (N_22829,N_21966,N_21865);
xor U22830 (N_22830,N_21774,N_21341);
nand U22831 (N_22831,N_21988,N_21928);
xor U22832 (N_22832,N_21403,N_21117);
xnor U22833 (N_22833,N_21418,N_21102);
nand U22834 (N_22834,N_21474,N_21460);
and U22835 (N_22835,N_21089,N_21808);
nand U22836 (N_22836,N_21422,N_21559);
nand U22837 (N_22837,N_21142,N_21129);
and U22838 (N_22838,N_21390,N_21622);
or U22839 (N_22839,N_21321,N_21049);
nor U22840 (N_22840,N_21404,N_21104);
nor U22841 (N_22841,N_21192,N_21122);
and U22842 (N_22842,N_21939,N_21411);
nor U22843 (N_22843,N_21507,N_21137);
or U22844 (N_22844,N_21711,N_21011);
nor U22845 (N_22845,N_21966,N_21891);
nor U22846 (N_22846,N_21148,N_21589);
nor U22847 (N_22847,N_21415,N_21269);
nor U22848 (N_22848,N_21908,N_21670);
or U22849 (N_22849,N_21283,N_21315);
nor U22850 (N_22850,N_21850,N_21207);
xnor U22851 (N_22851,N_21668,N_21652);
nor U22852 (N_22852,N_21915,N_21317);
nand U22853 (N_22853,N_21770,N_21343);
nand U22854 (N_22854,N_21615,N_21843);
and U22855 (N_22855,N_21444,N_21112);
xor U22856 (N_22856,N_21315,N_21304);
and U22857 (N_22857,N_21079,N_21194);
and U22858 (N_22858,N_21164,N_21825);
nor U22859 (N_22859,N_21853,N_21481);
xnor U22860 (N_22860,N_21815,N_21993);
nand U22861 (N_22861,N_21485,N_21807);
xor U22862 (N_22862,N_21774,N_21919);
xor U22863 (N_22863,N_21537,N_21523);
nand U22864 (N_22864,N_21074,N_21949);
nor U22865 (N_22865,N_21157,N_21163);
xor U22866 (N_22866,N_21850,N_21731);
or U22867 (N_22867,N_21346,N_21306);
or U22868 (N_22868,N_21826,N_21930);
or U22869 (N_22869,N_21215,N_21390);
or U22870 (N_22870,N_21339,N_21143);
and U22871 (N_22871,N_21053,N_21184);
or U22872 (N_22872,N_21927,N_21040);
nand U22873 (N_22873,N_21322,N_21896);
xor U22874 (N_22874,N_21096,N_21683);
nor U22875 (N_22875,N_21510,N_21420);
xor U22876 (N_22876,N_21939,N_21153);
and U22877 (N_22877,N_21285,N_21319);
and U22878 (N_22878,N_21056,N_21228);
nand U22879 (N_22879,N_21824,N_21210);
or U22880 (N_22880,N_21122,N_21463);
and U22881 (N_22881,N_21188,N_21077);
nor U22882 (N_22882,N_21910,N_21822);
or U22883 (N_22883,N_21291,N_21851);
or U22884 (N_22884,N_21061,N_21103);
nand U22885 (N_22885,N_21195,N_21091);
and U22886 (N_22886,N_21628,N_21609);
or U22887 (N_22887,N_21884,N_21995);
nand U22888 (N_22888,N_21340,N_21861);
nand U22889 (N_22889,N_21425,N_21576);
or U22890 (N_22890,N_21081,N_21893);
nor U22891 (N_22891,N_21388,N_21679);
xnor U22892 (N_22892,N_21874,N_21322);
and U22893 (N_22893,N_21386,N_21337);
nand U22894 (N_22894,N_21178,N_21923);
nor U22895 (N_22895,N_21138,N_21591);
and U22896 (N_22896,N_21097,N_21111);
nand U22897 (N_22897,N_21144,N_21707);
or U22898 (N_22898,N_21680,N_21436);
nor U22899 (N_22899,N_21886,N_21308);
and U22900 (N_22900,N_21278,N_21729);
or U22901 (N_22901,N_21965,N_21281);
and U22902 (N_22902,N_21229,N_21924);
or U22903 (N_22903,N_21978,N_21337);
and U22904 (N_22904,N_21802,N_21144);
and U22905 (N_22905,N_21176,N_21172);
or U22906 (N_22906,N_21930,N_21069);
nor U22907 (N_22907,N_21185,N_21619);
or U22908 (N_22908,N_21517,N_21594);
nand U22909 (N_22909,N_21753,N_21994);
and U22910 (N_22910,N_21557,N_21921);
nor U22911 (N_22911,N_21165,N_21011);
and U22912 (N_22912,N_21249,N_21853);
nor U22913 (N_22913,N_21713,N_21107);
and U22914 (N_22914,N_21062,N_21472);
nand U22915 (N_22915,N_21870,N_21647);
nand U22916 (N_22916,N_21300,N_21843);
nand U22917 (N_22917,N_21914,N_21689);
nor U22918 (N_22918,N_21238,N_21697);
nand U22919 (N_22919,N_21481,N_21905);
xor U22920 (N_22920,N_21537,N_21675);
nand U22921 (N_22921,N_21683,N_21645);
nand U22922 (N_22922,N_21507,N_21899);
or U22923 (N_22923,N_21752,N_21078);
and U22924 (N_22924,N_21299,N_21884);
nor U22925 (N_22925,N_21981,N_21173);
or U22926 (N_22926,N_21347,N_21076);
and U22927 (N_22927,N_21271,N_21974);
and U22928 (N_22928,N_21161,N_21889);
nand U22929 (N_22929,N_21518,N_21376);
and U22930 (N_22930,N_21596,N_21042);
or U22931 (N_22931,N_21553,N_21298);
or U22932 (N_22932,N_21285,N_21613);
xor U22933 (N_22933,N_21967,N_21067);
xnor U22934 (N_22934,N_21132,N_21467);
nand U22935 (N_22935,N_21340,N_21234);
nor U22936 (N_22936,N_21543,N_21355);
xnor U22937 (N_22937,N_21782,N_21541);
nand U22938 (N_22938,N_21970,N_21238);
xnor U22939 (N_22939,N_21699,N_21767);
xnor U22940 (N_22940,N_21933,N_21403);
xor U22941 (N_22941,N_21660,N_21914);
nor U22942 (N_22942,N_21803,N_21955);
and U22943 (N_22943,N_21270,N_21503);
xnor U22944 (N_22944,N_21100,N_21896);
and U22945 (N_22945,N_21930,N_21399);
xor U22946 (N_22946,N_21142,N_21058);
xnor U22947 (N_22947,N_21472,N_21244);
or U22948 (N_22948,N_21962,N_21501);
and U22949 (N_22949,N_21603,N_21297);
or U22950 (N_22950,N_21816,N_21378);
nand U22951 (N_22951,N_21388,N_21576);
nor U22952 (N_22952,N_21242,N_21407);
nor U22953 (N_22953,N_21769,N_21641);
nor U22954 (N_22954,N_21378,N_21097);
and U22955 (N_22955,N_21577,N_21184);
and U22956 (N_22956,N_21291,N_21147);
or U22957 (N_22957,N_21353,N_21711);
nor U22958 (N_22958,N_21646,N_21094);
xnor U22959 (N_22959,N_21644,N_21601);
nor U22960 (N_22960,N_21416,N_21296);
xor U22961 (N_22961,N_21606,N_21571);
nand U22962 (N_22962,N_21966,N_21490);
nor U22963 (N_22963,N_21320,N_21782);
or U22964 (N_22964,N_21340,N_21352);
nand U22965 (N_22965,N_21195,N_21547);
xnor U22966 (N_22966,N_21111,N_21661);
nor U22967 (N_22967,N_21571,N_21607);
xnor U22968 (N_22968,N_21771,N_21636);
or U22969 (N_22969,N_21722,N_21551);
or U22970 (N_22970,N_21792,N_21322);
nand U22971 (N_22971,N_21573,N_21403);
or U22972 (N_22972,N_21227,N_21726);
nor U22973 (N_22973,N_21310,N_21365);
nor U22974 (N_22974,N_21429,N_21548);
nor U22975 (N_22975,N_21418,N_21414);
nand U22976 (N_22976,N_21653,N_21300);
nand U22977 (N_22977,N_21605,N_21213);
or U22978 (N_22978,N_21191,N_21143);
xor U22979 (N_22979,N_21956,N_21585);
xor U22980 (N_22980,N_21601,N_21828);
nor U22981 (N_22981,N_21700,N_21912);
or U22982 (N_22982,N_21835,N_21209);
or U22983 (N_22983,N_21403,N_21780);
nand U22984 (N_22984,N_21977,N_21638);
xor U22985 (N_22985,N_21263,N_21833);
or U22986 (N_22986,N_21387,N_21768);
and U22987 (N_22987,N_21041,N_21536);
xnor U22988 (N_22988,N_21043,N_21299);
xnor U22989 (N_22989,N_21247,N_21724);
xnor U22990 (N_22990,N_21581,N_21506);
and U22991 (N_22991,N_21937,N_21171);
or U22992 (N_22992,N_21332,N_21529);
nor U22993 (N_22993,N_21767,N_21252);
xnor U22994 (N_22994,N_21313,N_21049);
or U22995 (N_22995,N_21133,N_21162);
and U22996 (N_22996,N_21508,N_21252);
or U22997 (N_22997,N_21268,N_21182);
xor U22998 (N_22998,N_21792,N_21003);
nor U22999 (N_22999,N_21100,N_21441);
xor U23000 (N_23000,N_22278,N_22985);
xnor U23001 (N_23001,N_22010,N_22740);
and U23002 (N_23002,N_22576,N_22963);
nand U23003 (N_23003,N_22606,N_22760);
or U23004 (N_23004,N_22149,N_22035);
or U23005 (N_23005,N_22747,N_22689);
xor U23006 (N_23006,N_22499,N_22437);
xnor U23007 (N_23007,N_22845,N_22702);
xnor U23008 (N_23008,N_22434,N_22113);
xor U23009 (N_23009,N_22106,N_22508);
or U23010 (N_23010,N_22743,N_22513);
nand U23011 (N_23011,N_22838,N_22954);
or U23012 (N_23012,N_22156,N_22700);
and U23013 (N_23013,N_22286,N_22738);
nor U23014 (N_23014,N_22175,N_22770);
and U23015 (N_23015,N_22983,N_22996);
xnor U23016 (N_23016,N_22557,N_22116);
nand U23017 (N_23017,N_22020,N_22707);
xnor U23018 (N_23018,N_22716,N_22455);
nor U23019 (N_23019,N_22739,N_22960);
nor U23020 (N_23020,N_22181,N_22772);
xor U23021 (N_23021,N_22890,N_22706);
nor U23022 (N_23022,N_22443,N_22241);
nor U23023 (N_23023,N_22386,N_22814);
and U23024 (N_23024,N_22379,N_22038);
and U23025 (N_23025,N_22327,N_22541);
xor U23026 (N_23026,N_22840,N_22193);
xor U23027 (N_23027,N_22503,N_22001);
nand U23028 (N_23028,N_22063,N_22006);
or U23029 (N_23029,N_22041,N_22151);
nor U23030 (N_23030,N_22782,N_22101);
xor U23031 (N_23031,N_22756,N_22600);
xor U23032 (N_23032,N_22886,N_22989);
nand U23033 (N_23033,N_22209,N_22311);
nand U23034 (N_23034,N_22257,N_22627);
xnor U23035 (N_23035,N_22710,N_22573);
nand U23036 (N_23036,N_22245,N_22687);
and U23037 (N_23037,N_22642,N_22092);
xor U23038 (N_23038,N_22381,N_22711);
and U23039 (N_23039,N_22862,N_22216);
and U23040 (N_23040,N_22164,N_22514);
xor U23041 (N_23041,N_22787,N_22359);
and U23042 (N_23042,N_22352,N_22653);
or U23043 (N_23043,N_22833,N_22993);
or U23044 (N_23044,N_22728,N_22540);
and U23045 (N_23045,N_22918,N_22030);
nand U23046 (N_23046,N_22506,N_22342);
nand U23047 (N_23047,N_22696,N_22808);
nor U23048 (N_23048,N_22575,N_22086);
and U23049 (N_23049,N_22774,N_22496);
xor U23050 (N_23050,N_22162,N_22959);
and U23051 (N_23051,N_22910,N_22318);
nand U23052 (N_23052,N_22465,N_22248);
xor U23053 (N_23053,N_22072,N_22394);
nor U23054 (N_23054,N_22812,N_22762);
or U23055 (N_23055,N_22228,N_22238);
and U23056 (N_23056,N_22049,N_22779);
xnor U23057 (N_23057,N_22045,N_22708);
and U23058 (N_23058,N_22801,N_22222);
or U23059 (N_23059,N_22119,N_22961);
xnor U23060 (N_23060,N_22877,N_22403);
nand U23061 (N_23061,N_22153,N_22486);
xnor U23062 (N_23062,N_22863,N_22387);
nor U23063 (N_23063,N_22721,N_22899);
or U23064 (N_23064,N_22681,N_22893);
nand U23065 (N_23065,N_22665,N_22539);
or U23066 (N_23066,N_22628,N_22614);
xor U23067 (N_23067,N_22570,N_22538);
nand U23068 (N_23068,N_22651,N_22444);
nor U23069 (N_23069,N_22326,N_22192);
xor U23070 (N_23070,N_22531,N_22805);
nor U23071 (N_23071,N_22075,N_22726);
xnor U23072 (N_23072,N_22841,N_22777);
or U23073 (N_23073,N_22406,N_22210);
or U23074 (N_23074,N_22139,N_22367);
nor U23075 (N_23075,N_22360,N_22942);
or U23076 (N_23076,N_22565,N_22727);
and U23077 (N_23077,N_22357,N_22013);
nor U23078 (N_23078,N_22264,N_22130);
nand U23079 (N_23079,N_22981,N_22551);
nor U23080 (N_23080,N_22811,N_22517);
xnor U23081 (N_23081,N_22867,N_22261);
nor U23082 (N_23082,N_22888,N_22876);
nand U23083 (N_23083,N_22043,N_22464);
or U23084 (N_23084,N_22339,N_22157);
or U23085 (N_23085,N_22929,N_22645);
or U23086 (N_23086,N_22980,N_22510);
and U23087 (N_23087,N_22401,N_22578);
and U23088 (N_23088,N_22125,N_22376);
nand U23089 (N_23089,N_22127,N_22921);
and U23090 (N_23090,N_22112,N_22477);
nor U23091 (N_23091,N_22036,N_22287);
nand U23092 (N_23092,N_22108,N_22236);
nand U23093 (N_23093,N_22999,N_22003);
nor U23094 (N_23094,N_22646,N_22518);
and U23095 (N_23095,N_22660,N_22306);
xnor U23096 (N_23096,N_22221,N_22136);
nor U23097 (N_23097,N_22611,N_22201);
xor U23098 (N_23098,N_22263,N_22804);
or U23099 (N_23099,N_22100,N_22958);
and U23100 (N_23100,N_22412,N_22884);
nor U23101 (N_23101,N_22023,N_22429);
xnor U23102 (N_23102,N_22355,N_22493);
nor U23103 (N_23103,N_22008,N_22577);
nand U23104 (N_23104,N_22559,N_22823);
or U23105 (N_23105,N_22522,N_22976);
or U23106 (N_23106,N_22968,N_22067);
nand U23107 (N_23107,N_22198,N_22189);
nor U23108 (N_23108,N_22898,N_22633);
xnor U23109 (N_23109,N_22419,N_22077);
or U23110 (N_23110,N_22583,N_22374);
nor U23111 (N_23111,N_22511,N_22074);
xor U23112 (N_23112,N_22759,N_22864);
xor U23113 (N_23113,N_22347,N_22810);
nand U23114 (N_23114,N_22613,N_22025);
and U23115 (N_23115,N_22421,N_22068);
or U23116 (N_23116,N_22620,N_22832);
xor U23117 (N_23117,N_22949,N_22753);
nand U23118 (N_23118,N_22322,N_22334);
nand U23119 (N_23119,N_22822,N_22213);
nand U23120 (N_23120,N_22219,N_22816);
nor U23121 (N_23121,N_22338,N_22553);
or U23122 (N_23122,N_22887,N_22644);
and U23123 (N_23123,N_22361,N_22117);
xor U23124 (N_23124,N_22647,N_22495);
xnor U23125 (N_23125,N_22071,N_22973);
or U23126 (N_23126,N_22861,N_22695);
or U23127 (N_23127,N_22826,N_22214);
xor U23128 (N_23128,N_22567,N_22280);
or U23129 (N_23129,N_22525,N_22215);
and U23130 (N_23130,N_22017,N_22672);
nor U23131 (N_23131,N_22792,N_22796);
and U23132 (N_23132,N_22470,N_22185);
and U23133 (N_23133,N_22791,N_22285);
nor U23134 (N_23134,N_22969,N_22643);
or U23135 (N_23135,N_22605,N_22485);
nor U23136 (N_23136,N_22093,N_22384);
and U23137 (N_23137,N_22232,N_22200);
nor U23138 (N_23138,N_22667,N_22988);
nor U23139 (N_23139,N_22450,N_22661);
nand U23140 (N_23140,N_22820,N_22415);
and U23141 (N_23141,N_22199,N_22436);
xor U23142 (N_23142,N_22408,N_22598);
xnor U23143 (N_23143,N_22732,N_22947);
and U23144 (N_23144,N_22195,N_22521);
nand U23145 (N_23145,N_22764,N_22941);
and U23146 (N_23146,N_22719,N_22244);
or U23147 (N_23147,N_22362,N_22031);
or U23148 (N_23148,N_22693,N_22196);
nor U23149 (N_23149,N_22677,N_22170);
or U23150 (N_23150,N_22602,N_22720);
xnor U23151 (N_23151,N_22622,N_22967);
nor U23152 (N_23152,N_22590,N_22396);
and U23153 (N_23153,N_22836,N_22656);
or U23154 (N_23154,N_22848,N_22502);
and U23155 (N_23155,N_22766,N_22407);
xnor U23156 (N_23156,N_22229,N_22048);
xor U23157 (N_23157,N_22410,N_22372);
nand U23158 (N_23158,N_22472,N_22892);
nand U23159 (N_23159,N_22579,N_22448);
and U23160 (N_23160,N_22858,N_22416);
xnor U23161 (N_23161,N_22270,N_22731);
nor U23162 (N_23162,N_22891,N_22223);
xor U23163 (N_23163,N_22377,N_22011);
and U23164 (N_23164,N_22128,N_22191);
nor U23165 (N_23165,N_22019,N_22735);
or U23166 (N_23166,N_22122,N_22922);
nand U23167 (N_23167,N_22267,N_22262);
nor U23168 (N_23168,N_22755,N_22424);
xnor U23169 (N_23169,N_22723,N_22088);
xor U23170 (N_23170,N_22725,N_22050);
nor U23171 (N_23171,N_22737,N_22505);
nand U23172 (N_23172,N_22780,N_22998);
nand U23173 (N_23173,N_22869,N_22631);
and U23174 (N_23174,N_22524,N_22055);
xor U23175 (N_23175,N_22282,N_22784);
xnor U23176 (N_23176,N_22303,N_22369);
and U23177 (N_23177,N_22205,N_22639);
nor U23178 (N_23178,N_22736,N_22005);
nand U23179 (N_23179,N_22875,N_22435);
and U23180 (N_23180,N_22178,N_22310);
nor U23181 (N_23181,N_22987,N_22333);
and U23182 (N_23182,N_22479,N_22305);
and U23183 (N_23183,N_22830,N_22155);
xnor U23184 (N_23184,N_22393,N_22586);
xnor U23185 (N_23185,N_22857,N_22649);
or U23186 (N_23186,N_22794,N_22924);
and U23187 (N_23187,N_22596,N_22659);
xnor U23188 (N_23188,N_22227,N_22217);
nor U23189 (N_23189,N_22474,N_22203);
and U23190 (N_23190,N_22276,N_22516);
nor U23191 (N_23191,N_22914,N_22817);
xnor U23192 (N_23192,N_22272,N_22373);
or U23193 (N_23193,N_22546,N_22397);
and U23194 (N_23194,N_22500,N_22060);
and U23195 (N_23195,N_22501,N_22348);
and U23196 (N_23196,N_22288,N_22901);
or U23197 (N_23197,N_22617,N_22463);
xnor U23198 (N_23198,N_22466,N_22004);
nand U23199 (N_23199,N_22957,N_22691);
xnor U23200 (N_23200,N_22658,N_22626);
nor U23201 (N_23201,N_22392,N_22591);
or U23202 (N_23202,N_22775,N_22344);
and U23203 (N_23203,N_22484,N_22945);
and U23204 (N_23204,N_22593,N_22849);
and U23205 (N_23205,N_22131,N_22635);
nand U23206 (N_23206,N_22654,N_22032);
nor U23207 (N_23207,N_22793,N_22800);
nor U23208 (N_23208,N_22595,N_22618);
nand U23209 (N_23209,N_22313,N_22225);
or U23210 (N_23210,N_22684,N_22330);
nand U23211 (N_23211,N_22529,N_22097);
xnor U23212 (N_23212,N_22574,N_22169);
nor U23213 (N_23213,N_22123,N_22970);
nand U23214 (N_23214,N_22928,N_22194);
nand U23215 (N_23215,N_22445,N_22323);
nand U23216 (N_23216,N_22294,N_22519);
nor U23217 (N_23217,N_22425,N_22184);
nand U23218 (N_23218,N_22490,N_22230);
or U23219 (N_23219,N_22834,N_22426);
nor U23220 (N_23220,N_22588,N_22964);
nor U23221 (N_23221,N_22204,N_22829);
nor U23222 (N_23222,N_22905,N_22129);
nor U23223 (N_23223,N_22678,N_22274);
xor U23224 (N_23224,N_22388,N_22478);
or U23225 (N_23225,N_22972,N_22370);
nand U23226 (N_23226,N_22281,N_22815);
nand U23227 (N_23227,N_22457,N_22473);
nand U23228 (N_23228,N_22992,N_22778);
nor U23229 (N_23229,N_22632,N_22343);
nand U23230 (N_23230,N_22309,N_22580);
or U23231 (N_23231,N_22955,N_22065);
nor U23232 (N_23232,N_22398,N_22034);
or U23233 (N_23233,N_22081,N_22509);
nand U23234 (N_23234,N_22956,N_22391);
nand U23235 (N_23235,N_22558,N_22094);
or U23236 (N_23236,N_22676,N_22975);
and U23237 (N_23237,N_22612,N_22172);
nor U23238 (N_23238,N_22610,N_22028);
nor U23239 (N_23239,N_22110,N_22908);
and U23240 (N_23240,N_22758,N_22137);
or U23241 (N_23241,N_22289,N_22087);
or U23242 (N_23242,N_22752,N_22483);
nand U23243 (N_23243,N_22233,N_22096);
xor U23244 (N_23244,N_22231,N_22866);
nand U23245 (N_23245,N_22159,N_22919);
nand U23246 (N_23246,N_22648,N_22940);
xor U23247 (N_23247,N_22247,N_22083);
and U23248 (N_23248,N_22991,N_22277);
nor U23249 (N_23249,N_22675,N_22293);
xnor U23250 (N_23250,N_22084,N_22349);
xnor U23251 (N_23251,N_22895,N_22066);
nand U23252 (N_23252,N_22183,N_22115);
nor U23253 (N_23253,N_22748,N_22329);
and U23254 (N_23254,N_22440,N_22847);
nand U23255 (N_23255,N_22694,N_22021);
xnor U23256 (N_23256,N_22053,N_22202);
nand U23257 (N_23257,N_22138,N_22033);
or U23258 (N_23258,N_22813,N_22368);
xor U23259 (N_23259,N_22843,N_22979);
nor U23260 (N_23260,N_22641,N_22315);
nor U23261 (N_23261,N_22176,N_22534);
xnor U23262 (N_23262,N_22930,N_22913);
nand U23263 (N_23263,N_22581,N_22317);
nor U23264 (N_23264,N_22383,N_22044);
xnor U23265 (N_23265,N_22916,N_22745);
and U23266 (N_23266,N_22560,N_22168);
or U23267 (N_23267,N_22603,N_22173);
nand U23268 (N_23268,N_22056,N_22301);
xnor U23269 (N_23269,N_22615,N_22144);
or U23270 (N_23270,N_22442,N_22366);
or U23271 (N_23271,N_22734,N_22167);
nor U23272 (N_23272,N_22265,N_22365);
nor U23273 (N_23273,N_22091,N_22134);
and U23274 (N_23274,N_22844,N_22704);
nor U23275 (N_23275,N_22533,N_22389);
or U23276 (N_23276,N_22337,N_22104);
xor U23277 (N_23277,N_22548,N_22331);
nand U23278 (N_23278,N_22554,N_22917);
or U23279 (N_23279,N_22385,N_22809);
nand U23280 (N_23280,N_22163,N_22312);
nand U23281 (N_23281,N_22015,N_22798);
nor U23282 (N_23282,N_22607,N_22564);
nor U23283 (N_23283,N_22432,N_22399);
xor U23284 (N_23284,N_22042,N_22934);
xor U23285 (N_23285,N_22405,N_22126);
or U23286 (N_23286,N_22824,N_22089);
nor U23287 (N_23287,N_22664,N_22180);
xnor U23288 (N_23288,N_22255,N_22630);
nand U23289 (N_23289,N_22480,N_22915);
or U23290 (N_23290,N_22860,N_22971);
nand U23291 (N_23291,N_22962,N_22489);
xor U23292 (N_23292,N_22275,N_22135);
nor U23293 (N_23293,N_22253,N_22240);
or U23294 (N_23294,N_22118,N_22498);
or U23295 (N_23295,N_22492,N_22059);
or U23296 (N_23296,N_22121,N_22190);
and U23297 (N_23297,N_22951,N_22268);
nor U23298 (N_23298,N_22346,N_22585);
or U23299 (N_23299,N_22304,N_22781);
xnor U23300 (N_23300,N_22939,N_22460);
xor U23301 (N_23301,N_22571,N_22828);
and U23302 (N_23302,N_22773,N_22390);
and U23303 (N_23303,N_22754,N_22601);
nand U23304 (N_23304,N_22446,N_22894);
or U23305 (N_23305,N_22336,N_22179);
xor U23306 (N_23306,N_22783,N_22024);
nor U23307 (N_23307,N_22459,N_22938);
or U23308 (N_23308,N_22324,N_22458);
nand U23309 (N_23309,N_22160,N_22948);
nand U23310 (N_23310,N_22378,N_22690);
or U23311 (N_23311,N_22920,N_22872);
or U23312 (N_23312,N_22873,N_22523);
xnor U23313 (N_23313,N_22143,N_22604);
or U23314 (N_23314,N_22047,N_22952);
nor U23315 (N_23315,N_22371,N_22284);
xnor U23316 (N_23316,N_22109,N_22133);
nor U23317 (N_23317,N_22683,N_22657);
nand U23318 (N_23318,N_22904,N_22402);
nor U23319 (N_23319,N_22880,N_22467);
xor U23320 (N_23320,N_22741,N_22882);
xnor U23321 (N_23321,N_22532,N_22789);
xnor U23322 (N_23322,N_22332,N_22543);
xnor U23323 (N_23323,N_22197,N_22174);
nand U23324 (N_23324,N_22099,N_22846);
xor U23325 (N_23325,N_22224,N_22943);
and U23326 (N_23326,N_22290,N_22986);
xor U23327 (N_23327,N_22624,N_22431);
or U23328 (N_23328,N_22569,N_22208);
nand U23329 (N_23329,N_22680,N_22249);
and U23330 (N_23330,N_22854,N_22350);
or U23331 (N_23331,N_22400,N_22562);
nor U23332 (N_23332,N_22650,N_22563);
nor U23333 (N_23333,N_22026,N_22572);
xor U23334 (N_23334,N_22380,N_22902);
and U23335 (N_23335,N_22556,N_22655);
and U23336 (N_23336,N_22321,N_22243);
nand U23337 (N_23337,N_22364,N_22923);
and U23338 (N_23338,N_22291,N_22561);
nand U23339 (N_23339,N_22619,N_22530);
nand U23340 (N_23340,N_22307,N_22266);
nand U23341 (N_23341,N_22358,N_22427);
nand U23342 (N_23342,N_22166,N_22422);
nor U23343 (N_23343,N_22395,N_22636);
or U23344 (N_23344,N_22051,N_22932);
nor U23345 (N_23345,N_22767,N_22080);
nor U23346 (N_23346,N_22242,N_22714);
xnor U23347 (N_23347,N_22608,N_22666);
nor U23348 (N_23348,N_22273,N_22152);
xnor U23349 (N_23349,N_22878,N_22621);
nor U23350 (N_23350,N_22933,N_22682);
or U23351 (N_23351,N_22016,N_22982);
or U23352 (N_23352,N_22146,N_22868);
nor U23353 (N_23353,N_22404,N_22881);
or U23354 (N_23354,N_22430,N_22413);
or U23355 (N_23355,N_22111,N_22461);
nor U23356 (N_23356,N_22452,N_22990);
xnor U23357 (N_23357,N_22308,N_22507);
and U23358 (N_23358,N_22438,N_22148);
and U23359 (N_23359,N_22686,N_22865);
nand U23360 (N_23360,N_22742,N_22252);
or U23361 (N_23361,N_22504,N_22925);
xnor U23362 (N_23362,N_22977,N_22078);
or U23363 (N_23363,N_22314,N_22763);
or U23364 (N_23364,N_22000,N_22802);
nand U23365 (N_23365,N_22512,N_22488);
xnor U23366 (N_23366,N_22037,N_22211);
nand U23367 (N_23367,N_22147,N_22002);
nor U23368 (N_23368,N_22296,N_22014);
xor U23369 (N_23369,N_22462,N_22629);
xor U23370 (N_23370,N_22729,N_22837);
xor U23371 (N_23371,N_22965,N_22145);
or U23372 (N_23372,N_22871,N_22827);
nand U23373 (N_23373,N_22382,N_22698);
and U23374 (N_23374,N_22715,N_22730);
xor U23375 (N_23375,N_22420,N_22995);
xnor U23376 (N_23376,N_22453,N_22414);
nor U23377 (N_23377,N_22544,N_22879);
xnor U23378 (N_23378,N_22946,N_22454);
xor U23379 (N_23379,N_22733,N_22476);
nand U23380 (N_23380,N_22375,N_22098);
and U23381 (N_23381,N_22771,N_22102);
or U23382 (N_23382,N_22839,N_22718);
or U23383 (N_23383,N_22701,N_22212);
or U23384 (N_23384,N_22254,N_22353);
and U23385 (N_23385,N_22335,N_22447);
xnor U23386 (N_23386,N_22937,N_22746);
and U23387 (N_23387,N_22825,N_22589);
and U23388 (N_23388,N_22269,N_22883);
nor U23389 (N_23389,N_22070,N_22885);
or U23390 (N_23390,N_22107,N_22064);
and U23391 (N_23391,N_22206,N_22161);
or U23392 (N_23392,N_22757,N_22668);
nand U23393 (N_23393,N_22132,N_22251);
xor U23394 (N_23394,N_22842,N_22114);
xor U23395 (N_23395,N_22906,N_22054);
or U23396 (N_23396,N_22316,N_22853);
nand U23397 (N_23397,N_22340,N_22697);
nand U23398 (N_23398,N_22363,N_22090);
or U23399 (N_23399,N_22487,N_22870);
and U23400 (N_23400,N_22984,N_22768);
nor U23401 (N_23401,N_22471,N_22069);
nor U23402 (N_23402,N_22302,N_22936);
nand U23403 (N_23403,N_22256,N_22012);
and U23404 (N_23404,N_22526,N_22061);
nor U23405 (N_23405,N_22803,N_22897);
and U23406 (N_23406,N_22931,N_22186);
nor U23407 (N_23407,N_22491,N_22859);
nand U23408 (N_23408,N_22515,N_22165);
or U23409 (N_23409,N_22142,N_22835);
nor U23410 (N_23410,N_22785,N_22950);
nor U23411 (N_23411,N_22409,N_22351);
nand U23412 (N_23412,N_22703,N_22027);
and U23413 (N_23413,N_22679,N_22537);
nor U23414 (N_23414,N_22239,N_22062);
or U23415 (N_23415,N_22007,N_22547);
xnor U23416 (N_23416,N_22926,N_22260);
xor U23417 (N_23417,N_22482,N_22765);
and U23418 (N_23418,N_22594,N_22788);
nand U23419 (N_23419,N_22283,N_22769);
xor U23420 (N_23420,N_22029,N_22587);
xor U23421 (N_23421,N_22456,N_22799);
or U23422 (N_23422,N_22207,N_22354);
nand U23423 (N_23423,N_22712,N_22699);
or U23424 (N_23424,N_22433,N_22124);
and U23425 (N_23425,N_22625,N_22623);
nor U23426 (N_23426,N_22751,N_22927);
and U23427 (N_23427,N_22057,N_22674);
nor U23428 (N_23428,N_22896,N_22806);
nand U23429 (N_23429,N_22085,N_22549);
and U23430 (N_23430,N_22441,N_22079);
nand U23431 (N_23431,N_22966,N_22009);
or U23432 (N_23432,N_22235,N_22497);
xnor U23433 (N_23433,N_22912,N_22692);
or U23434 (N_23434,N_22807,N_22411);
xnor U23435 (N_23435,N_22328,N_22671);
or U23436 (N_23436,N_22582,N_22713);
and U23437 (N_23437,N_22609,N_22226);
nand U23438 (N_23438,N_22439,N_22974);
nor U23439 (N_23439,N_22909,N_22761);
nand U23440 (N_23440,N_22994,N_22978);
and U23441 (N_23441,N_22592,N_22237);
xnor U23442 (N_23442,N_22542,N_22907);
or U23443 (N_23443,N_22105,N_22299);
and U23444 (N_23444,N_22856,N_22250);
and U23445 (N_23445,N_22776,N_22652);
nor U23446 (N_23446,N_22259,N_22295);
nand U23447 (N_23447,N_22150,N_22140);
or U23448 (N_23448,N_22082,N_22046);
nor U23449 (N_23449,N_22550,N_22171);
or U23450 (N_23450,N_22935,N_22744);
nand U23451 (N_23451,N_22058,N_22022);
nand U23452 (N_23452,N_22889,N_22188);
and U23453 (N_23453,N_22218,N_22786);
nor U23454 (N_23454,N_22634,N_22423);
nand U23455 (N_23455,N_22120,N_22177);
nor U23456 (N_23456,N_22527,N_22790);
nand U23457 (N_23457,N_22795,N_22319);
and U23458 (N_23458,N_22182,N_22076);
or U23459 (N_23459,N_22852,N_22717);
nand U23460 (N_23460,N_22039,N_22356);
nand U23461 (N_23461,N_22494,N_22481);
xor U23462 (N_23462,N_22345,N_22536);
and U23463 (N_23463,N_22095,N_22320);
or U23464 (N_23464,N_22688,N_22292);
or U23465 (N_23465,N_22750,N_22451);
nor U23466 (N_23466,N_22475,N_22428);
xnor U23467 (N_23467,N_22797,N_22662);
nand U23468 (N_23468,N_22831,N_22663);
xnor U23469 (N_23469,N_22040,N_22749);
nor U23470 (N_23470,N_22325,N_22903);
or U23471 (N_23471,N_22545,N_22997);
nor U23472 (N_23472,N_22555,N_22246);
nor U23473 (N_23473,N_22449,N_22552);
xnor U23474 (N_23474,N_22418,N_22818);
xor U23475 (N_23475,N_22584,N_22535);
nand U23476 (N_23476,N_22911,N_22468);
nor U23477 (N_23477,N_22052,N_22851);
and U23478 (N_23478,N_22724,N_22821);
nand U23479 (N_23479,N_22953,N_22566);
xor U23480 (N_23480,N_22669,N_22234);
and U23481 (N_23481,N_22722,N_22637);
or U23482 (N_23482,N_22685,N_22220);
or U23483 (N_23483,N_22819,N_22597);
and U23484 (N_23484,N_22673,N_22855);
and U23485 (N_23485,N_22297,N_22638);
or U23486 (N_23486,N_22158,N_22417);
and U23487 (N_23487,N_22141,N_22279);
and U23488 (N_23488,N_22874,N_22709);
and U23489 (N_23489,N_22599,N_22154);
xor U23490 (N_23490,N_22944,N_22018);
or U23491 (N_23491,N_22271,N_22298);
and U23492 (N_23492,N_22469,N_22073);
nand U23493 (N_23493,N_22187,N_22705);
nor U23494 (N_23494,N_22616,N_22850);
and U23495 (N_23495,N_22670,N_22900);
or U23496 (N_23496,N_22520,N_22341);
nor U23497 (N_23497,N_22258,N_22568);
xnor U23498 (N_23498,N_22300,N_22103);
xnor U23499 (N_23499,N_22528,N_22640);
nor U23500 (N_23500,N_22053,N_22466);
nor U23501 (N_23501,N_22520,N_22008);
nand U23502 (N_23502,N_22125,N_22404);
and U23503 (N_23503,N_22233,N_22329);
xnor U23504 (N_23504,N_22775,N_22735);
nor U23505 (N_23505,N_22439,N_22409);
nand U23506 (N_23506,N_22541,N_22002);
xnor U23507 (N_23507,N_22292,N_22739);
or U23508 (N_23508,N_22307,N_22867);
xor U23509 (N_23509,N_22455,N_22440);
nor U23510 (N_23510,N_22983,N_22372);
nor U23511 (N_23511,N_22120,N_22374);
or U23512 (N_23512,N_22754,N_22694);
nand U23513 (N_23513,N_22530,N_22873);
xor U23514 (N_23514,N_22639,N_22530);
nand U23515 (N_23515,N_22391,N_22406);
nor U23516 (N_23516,N_22089,N_22401);
nor U23517 (N_23517,N_22906,N_22259);
and U23518 (N_23518,N_22373,N_22828);
nand U23519 (N_23519,N_22975,N_22091);
nand U23520 (N_23520,N_22140,N_22823);
and U23521 (N_23521,N_22565,N_22820);
xor U23522 (N_23522,N_22523,N_22026);
or U23523 (N_23523,N_22588,N_22503);
xnor U23524 (N_23524,N_22174,N_22406);
or U23525 (N_23525,N_22818,N_22478);
xnor U23526 (N_23526,N_22155,N_22092);
xnor U23527 (N_23527,N_22147,N_22695);
and U23528 (N_23528,N_22569,N_22532);
nor U23529 (N_23529,N_22408,N_22187);
nand U23530 (N_23530,N_22765,N_22466);
or U23531 (N_23531,N_22564,N_22471);
nor U23532 (N_23532,N_22039,N_22436);
nand U23533 (N_23533,N_22037,N_22403);
xor U23534 (N_23534,N_22807,N_22742);
and U23535 (N_23535,N_22128,N_22149);
or U23536 (N_23536,N_22466,N_22556);
nor U23537 (N_23537,N_22936,N_22982);
xor U23538 (N_23538,N_22430,N_22954);
and U23539 (N_23539,N_22585,N_22111);
and U23540 (N_23540,N_22332,N_22325);
and U23541 (N_23541,N_22282,N_22558);
and U23542 (N_23542,N_22485,N_22325);
nand U23543 (N_23543,N_22816,N_22842);
and U23544 (N_23544,N_22294,N_22177);
or U23545 (N_23545,N_22303,N_22895);
nor U23546 (N_23546,N_22205,N_22911);
and U23547 (N_23547,N_22098,N_22184);
nand U23548 (N_23548,N_22013,N_22870);
and U23549 (N_23549,N_22922,N_22297);
xor U23550 (N_23550,N_22493,N_22453);
and U23551 (N_23551,N_22955,N_22843);
nand U23552 (N_23552,N_22579,N_22190);
xnor U23553 (N_23553,N_22281,N_22353);
xnor U23554 (N_23554,N_22808,N_22420);
or U23555 (N_23555,N_22758,N_22470);
and U23556 (N_23556,N_22959,N_22477);
nand U23557 (N_23557,N_22284,N_22579);
nand U23558 (N_23558,N_22623,N_22759);
or U23559 (N_23559,N_22028,N_22939);
nor U23560 (N_23560,N_22112,N_22249);
and U23561 (N_23561,N_22611,N_22659);
and U23562 (N_23562,N_22562,N_22336);
and U23563 (N_23563,N_22900,N_22321);
and U23564 (N_23564,N_22388,N_22397);
or U23565 (N_23565,N_22851,N_22106);
nor U23566 (N_23566,N_22985,N_22623);
nor U23567 (N_23567,N_22614,N_22811);
or U23568 (N_23568,N_22419,N_22393);
nand U23569 (N_23569,N_22643,N_22586);
or U23570 (N_23570,N_22151,N_22894);
nor U23571 (N_23571,N_22125,N_22424);
nand U23572 (N_23572,N_22013,N_22391);
and U23573 (N_23573,N_22178,N_22837);
and U23574 (N_23574,N_22729,N_22727);
xnor U23575 (N_23575,N_22994,N_22876);
and U23576 (N_23576,N_22102,N_22902);
nand U23577 (N_23577,N_22692,N_22331);
and U23578 (N_23578,N_22091,N_22682);
nand U23579 (N_23579,N_22742,N_22703);
xnor U23580 (N_23580,N_22095,N_22663);
nand U23581 (N_23581,N_22570,N_22661);
or U23582 (N_23582,N_22973,N_22272);
and U23583 (N_23583,N_22942,N_22862);
xnor U23584 (N_23584,N_22036,N_22009);
or U23585 (N_23585,N_22850,N_22878);
or U23586 (N_23586,N_22509,N_22163);
xnor U23587 (N_23587,N_22827,N_22329);
or U23588 (N_23588,N_22774,N_22358);
or U23589 (N_23589,N_22015,N_22073);
nand U23590 (N_23590,N_22891,N_22478);
nor U23591 (N_23591,N_22419,N_22465);
nand U23592 (N_23592,N_22298,N_22294);
and U23593 (N_23593,N_22488,N_22229);
xnor U23594 (N_23594,N_22762,N_22300);
and U23595 (N_23595,N_22556,N_22571);
nor U23596 (N_23596,N_22133,N_22111);
xnor U23597 (N_23597,N_22359,N_22732);
or U23598 (N_23598,N_22632,N_22947);
xor U23599 (N_23599,N_22122,N_22197);
and U23600 (N_23600,N_22005,N_22184);
nor U23601 (N_23601,N_22815,N_22552);
nor U23602 (N_23602,N_22616,N_22704);
and U23603 (N_23603,N_22341,N_22933);
xnor U23604 (N_23604,N_22368,N_22004);
nand U23605 (N_23605,N_22791,N_22626);
nor U23606 (N_23606,N_22698,N_22880);
xor U23607 (N_23607,N_22379,N_22566);
and U23608 (N_23608,N_22632,N_22066);
nand U23609 (N_23609,N_22765,N_22699);
xnor U23610 (N_23610,N_22047,N_22324);
xnor U23611 (N_23611,N_22149,N_22752);
nor U23612 (N_23612,N_22778,N_22601);
or U23613 (N_23613,N_22965,N_22383);
or U23614 (N_23614,N_22614,N_22145);
nor U23615 (N_23615,N_22126,N_22288);
nand U23616 (N_23616,N_22207,N_22451);
nand U23617 (N_23617,N_22922,N_22154);
or U23618 (N_23618,N_22525,N_22954);
nand U23619 (N_23619,N_22965,N_22776);
or U23620 (N_23620,N_22704,N_22663);
nand U23621 (N_23621,N_22096,N_22013);
or U23622 (N_23622,N_22622,N_22187);
nand U23623 (N_23623,N_22862,N_22543);
or U23624 (N_23624,N_22554,N_22958);
nor U23625 (N_23625,N_22933,N_22213);
or U23626 (N_23626,N_22023,N_22359);
and U23627 (N_23627,N_22338,N_22030);
and U23628 (N_23628,N_22721,N_22378);
nand U23629 (N_23629,N_22211,N_22047);
and U23630 (N_23630,N_22971,N_22277);
or U23631 (N_23631,N_22738,N_22727);
nand U23632 (N_23632,N_22860,N_22471);
and U23633 (N_23633,N_22466,N_22050);
and U23634 (N_23634,N_22724,N_22451);
nand U23635 (N_23635,N_22704,N_22501);
xor U23636 (N_23636,N_22019,N_22914);
and U23637 (N_23637,N_22259,N_22063);
xor U23638 (N_23638,N_22544,N_22582);
nor U23639 (N_23639,N_22634,N_22900);
nand U23640 (N_23640,N_22732,N_22723);
xor U23641 (N_23641,N_22364,N_22902);
and U23642 (N_23642,N_22950,N_22116);
nor U23643 (N_23643,N_22178,N_22256);
xnor U23644 (N_23644,N_22524,N_22522);
and U23645 (N_23645,N_22916,N_22929);
nand U23646 (N_23646,N_22616,N_22183);
and U23647 (N_23647,N_22333,N_22473);
xnor U23648 (N_23648,N_22445,N_22606);
nand U23649 (N_23649,N_22055,N_22406);
or U23650 (N_23650,N_22240,N_22306);
and U23651 (N_23651,N_22815,N_22921);
xor U23652 (N_23652,N_22035,N_22454);
or U23653 (N_23653,N_22270,N_22611);
xor U23654 (N_23654,N_22478,N_22176);
xnor U23655 (N_23655,N_22574,N_22017);
nand U23656 (N_23656,N_22803,N_22163);
or U23657 (N_23657,N_22525,N_22651);
nand U23658 (N_23658,N_22892,N_22750);
nand U23659 (N_23659,N_22823,N_22199);
nor U23660 (N_23660,N_22918,N_22750);
nand U23661 (N_23661,N_22274,N_22138);
xnor U23662 (N_23662,N_22575,N_22497);
nand U23663 (N_23663,N_22248,N_22626);
xnor U23664 (N_23664,N_22969,N_22604);
nor U23665 (N_23665,N_22769,N_22230);
xnor U23666 (N_23666,N_22859,N_22363);
nor U23667 (N_23667,N_22160,N_22231);
or U23668 (N_23668,N_22539,N_22083);
or U23669 (N_23669,N_22680,N_22142);
nor U23670 (N_23670,N_22320,N_22288);
nand U23671 (N_23671,N_22850,N_22908);
xnor U23672 (N_23672,N_22157,N_22282);
nor U23673 (N_23673,N_22346,N_22711);
xnor U23674 (N_23674,N_22171,N_22595);
nor U23675 (N_23675,N_22324,N_22537);
and U23676 (N_23676,N_22822,N_22251);
xor U23677 (N_23677,N_22956,N_22596);
xor U23678 (N_23678,N_22697,N_22876);
xnor U23679 (N_23679,N_22123,N_22112);
nand U23680 (N_23680,N_22023,N_22203);
nand U23681 (N_23681,N_22159,N_22625);
nor U23682 (N_23682,N_22347,N_22334);
or U23683 (N_23683,N_22198,N_22337);
and U23684 (N_23684,N_22774,N_22990);
xor U23685 (N_23685,N_22717,N_22700);
nor U23686 (N_23686,N_22382,N_22526);
and U23687 (N_23687,N_22682,N_22344);
xor U23688 (N_23688,N_22477,N_22715);
nand U23689 (N_23689,N_22108,N_22468);
or U23690 (N_23690,N_22998,N_22188);
nor U23691 (N_23691,N_22023,N_22823);
xnor U23692 (N_23692,N_22133,N_22090);
xnor U23693 (N_23693,N_22626,N_22397);
nor U23694 (N_23694,N_22666,N_22391);
nor U23695 (N_23695,N_22200,N_22796);
or U23696 (N_23696,N_22186,N_22237);
and U23697 (N_23697,N_22527,N_22738);
nor U23698 (N_23698,N_22938,N_22206);
and U23699 (N_23699,N_22720,N_22229);
and U23700 (N_23700,N_22717,N_22285);
nor U23701 (N_23701,N_22445,N_22415);
and U23702 (N_23702,N_22326,N_22362);
nor U23703 (N_23703,N_22581,N_22874);
or U23704 (N_23704,N_22697,N_22398);
nor U23705 (N_23705,N_22942,N_22783);
or U23706 (N_23706,N_22933,N_22052);
and U23707 (N_23707,N_22537,N_22598);
or U23708 (N_23708,N_22923,N_22019);
nand U23709 (N_23709,N_22901,N_22193);
xnor U23710 (N_23710,N_22323,N_22754);
xnor U23711 (N_23711,N_22976,N_22022);
or U23712 (N_23712,N_22343,N_22777);
and U23713 (N_23713,N_22932,N_22184);
xnor U23714 (N_23714,N_22137,N_22872);
nand U23715 (N_23715,N_22718,N_22667);
xor U23716 (N_23716,N_22863,N_22080);
nor U23717 (N_23717,N_22681,N_22412);
nor U23718 (N_23718,N_22210,N_22361);
or U23719 (N_23719,N_22642,N_22774);
and U23720 (N_23720,N_22937,N_22154);
nand U23721 (N_23721,N_22487,N_22232);
xnor U23722 (N_23722,N_22595,N_22665);
xnor U23723 (N_23723,N_22679,N_22160);
or U23724 (N_23724,N_22037,N_22428);
or U23725 (N_23725,N_22004,N_22853);
nor U23726 (N_23726,N_22255,N_22544);
nor U23727 (N_23727,N_22425,N_22334);
nand U23728 (N_23728,N_22993,N_22096);
and U23729 (N_23729,N_22350,N_22912);
nand U23730 (N_23730,N_22989,N_22239);
nand U23731 (N_23731,N_22850,N_22253);
nor U23732 (N_23732,N_22897,N_22354);
and U23733 (N_23733,N_22589,N_22099);
or U23734 (N_23734,N_22608,N_22330);
nand U23735 (N_23735,N_22829,N_22084);
nor U23736 (N_23736,N_22315,N_22406);
or U23737 (N_23737,N_22181,N_22724);
nor U23738 (N_23738,N_22688,N_22019);
or U23739 (N_23739,N_22271,N_22095);
nor U23740 (N_23740,N_22345,N_22371);
nand U23741 (N_23741,N_22424,N_22641);
nand U23742 (N_23742,N_22529,N_22496);
nor U23743 (N_23743,N_22715,N_22850);
nand U23744 (N_23744,N_22031,N_22378);
nor U23745 (N_23745,N_22853,N_22900);
nor U23746 (N_23746,N_22870,N_22369);
and U23747 (N_23747,N_22003,N_22275);
or U23748 (N_23748,N_22579,N_22526);
nand U23749 (N_23749,N_22829,N_22566);
xnor U23750 (N_23750,N_22827,N_22696);
or U23751 (N_23751,N_22191,N_22352);
and U23752 (N_23752,N_22403,N_22456);
nor U23753 (N_23753,N_22127,N_22808);
nand U23754 (N_23754,N_22719,N_22627);
xor U23755 (N_23755,N_22545,N_22301);
and U23756 (N_23756,N_22820,N_22725);
and U23757 (N_23757,N_22616,N_22233);
or U23758 (N_23758,N_22438,N_22411);
nand U23759 (N_23759,N_22158,N_22080);
nor U23760 (N_23760,N_22681,N_22954);
and U23761 (N_23761,N_22063,N_22699);
or U23762 (N_23762,N_22352,N_22018);
or U23763 (N_23763,N_22281,N_22311);
nand U23764 (N_23764,N_22366,N_22203);
or U23765 (N_23765,N_22141,N_22880);
and U23766 (N_23766,N_22516,N_22631);
nor U23767 (N_23767,N_22503,N_22396);
and U23768 (N_23768,N_22594,N_22805);
xor U23769 (N_23769,N_22391,N_22490);
xnor U23770 (N_23770,N_22283,N_22705);
nor U23771 (N_23771,N_22185,N_22072);
nor U23772 (N_23772,N_22491,N_22492);
xor U23773 (N_23773,N_22363,N_22238);
xor U23774 (N_23774,N_22573,N_22518);
xor U23775 (N_23775,N_22661,N_22598);
or U23776 (N_23776,N_22259,N_22147);
nor U23777 (N_23777,N_22201,N_22185);
and U23778 (N_23778,N_22183,N_22399);
and U23779 (N_23779,N_22762,N_22489);
nand U23780 (N_23780,N_22464,N_22081);
xnor U23781 (N_23781,N_22089,N_22100);
and U23782 (N_23782,N_22448,N_22768);
and U23783 (N_23783,N_22034,N_22193);
nand U23784 (N_23784,N_22796,N_22210);
nand U23785 (N_23785,N_22268,N_22674);
or U23786 (N_23786,N_22457,N_22210);
or U23787 (N_23787,N_22886,N_22855);
nand U23788 (N_23788,N_22258,N_22909);
nor U23789 (N_23789,N_22946,N_22834);
nor U23790 (N_23790,N_22239,N_22669);
and U23791 (N_23791,N_22231,N_22157);
and U23792 (N_23792,N_22437,N_22579);
nor U23793 (N_23793,N_22796,N_22919);
or U23794 (N_23794,N_22446,N_22657);
nor U23795 (N_23795,N_22131,N_22555);
nor U23796 (N_23796,N_22907,N_22968);
or U23797 (N_23797,N_22125,N_22374);
nor U23798 (N_23798,N_22036,N_22588);
nand U23799 (N_23799,N_22287,N_22672);
and U23800 (N_23800,N_22591,N_22051);
nand U23801 (N_23801,N_22257,N_22120);
and U23802 (N_23802,N_22529,N_22212);
xor U23803 (N_23803,N_22711,N_22369);
and U23804 (N_23804,N_22175,N_22313);
nor U23805 (N_23805,N_22309,N_22296);
nand U23806 (N_23806,N_22153,N_22272);
nand U23807 (N_23807,N_22764,N_22307);
nand U23808 (N_23808,N_22646,N_22307);
or U23809 (N_23809,N_22649,N_22006);
or U23810 (N_23810,N_22055,N_22418);
nor U23811 (N_23811,N_22325,N_22870);
or U23812 (N_23812,N_22984,N_22460);
xnor U23813 (N_23813,N_22267,N_22277);
or U23814 (N_23814,N_22001,N_22016);
nor U23815 (N_23815,N_22074,N_22177);
and U23816 (N_23816,N_22043,N_22628);
and U23817 (N_23817,N_22848,N_22789);
and U23818 (N_23818,N_22075,N_22084);
or U23819 (N_23819,N_22365,N_22942);
xor U23820 (N_23820,N_22696,N_22490);
nand U23821 (N_23821,N_22900,N_22315);
nand U23822 (N_23822,N_22974,N_22876);
xor U23823 (N_23823,N_22055,N_22829);
nor U23824 (N_23824,N_22617,N_22984);
and U23825 (N_23825,N_22522,N_22640);
or U23826 (N_23826,N_22218,N_22644);
or U23827 (N_23827,N_22130,N_22619);
and U23828 (N_23828,N_22516,N_22792);
nand U23829 (N_23829,N_22399,N_22209);
and U23830 (N_23830,N_22386,N_22099);
nor U23831 (N_23831,N_22521,N_22481);
and U23832 (N_23832,N_22005,N_22447);
xor U23833 (N_23833,N_22058,N_22651);
xnor U23834 (N_23834,N_22573,N_22543);
nor U23835 (N_23835,N_22836,N_22563);
and U23836 (N_23836,N_22655,N_22457);
xor U23837 (N_23837,N_22392,N_22134);
xor U23838 (N_23838,N_22052,N_22376);
nor U23839 (N_23839,N_22119,N_22223);
and U23840 (N_23840,N_22029,N_22918);
and U23841 (N_23841,N_22813,N_22506);
or U23842 (N_23842,N_22486,N_22865);
nand U23843 (N_23843,N_22137,N_22135);
nand U23844 (N_23844,N_22567,N_22792);
nor U23845 (N_23845,N_22448,N_22488);
or U23846 (N_23846,N_22389,N_22013);
or U23847 (N_23847,N_22005,N_22563);
or U23848 (N_23848,N_22321,N_22669);
and U23849 (N_23849,N_22438,N_22986);
or U23850 (N_23850,N_22189,N_22079);
xor U23851 (N_23851,N_22626,N_22245);
or U23852 (N_23852,N_22770,N_22282);
xor U23853 (N_23853,N_22332,N_22927);
nand U23854 (N_23854,N_22843,N_22861);
nand U23855 (N_23855,N_22485,N_22449);
nand U23856 (N_23856,N_22017,N_22768);
nor U23857 (N_23857,N_22699,N_22998);
nand U23858 (N_23858,N_22023,N_22873);
xnor U23859 (N_23859,N_22451,N_22592);
xnor U23860 (N_23860,N_22275,N_22454);
nand U23861 (N_23861,N_22068,N_22453);
nand U23862 (N_23862,N_22921,N_22508);
or U23863 (N_23863,N_22989,N_22332);
nand U23864 (N_23864,N_22243,N_22049);
or U23865 (N_23865,N_22446,N_22145);
and U23866 (N_23866,N_22212,N_22788);
nor U23867 (N_23867,N_22707,N_22855);
and U23868 (N_23868,N_22634,N_22517);
nor U23869 (N_23869,N_22819,N_22647);
and U23870 (N_23870,N_22798,N_22921);
nand U23871 (N_23871,N_22497,N_22351);
nor U23872 (N_23872,N_22984,N_22485);
or U23873 (N_23873,N_22680,N_22447);
nor U23874 (N_23874,N_22036,N_22181);
nand U23875 (N_23875,N_22212,N_22232);
and U23876 (N_23876,N_22820,N_22717);
xor U23877 (N_23877,N_22596,N_22399);
and U23878 (N_23878,N_22819,N_22555);
nor U23879 (N_23879,N_22585,N_22219);
nand U23880 (N_23880,N_22570,N_22799);
and U23881 (N_23881,N_22154,N_22475);
and U23882 (N_23882,N_22545,N_22253);
xor U23883 (N_23883,N_22230,N_22531);
nand U23884 (N_23884,N_22193,N_22891);
nor U23885 (N_23885,N_22590,N_22926);
nor U23886 (N_23886,N_22425,N_22215);
or U23887 (N_23887,N_22557,N_22277);
nor U23888 (N_23888,N_22397,N_22328);
xnor U23889 (N_23889,N_22899,N_22931);
or U23890 (N_23890,N_22580,N_22924);
and U23891 (N_23891,N_22651,N_22325);
nor U23892 (N_23892,N_22947,N_22060);
nand U23893 (N_23893,N_22172,N_22814);
xor U23894 (N_23894,N_22228,N_22999);
and U23895 (N_23895,N_22932,N_22908);
nor U23896 (N_23896,N_22985,N_22015);
nor U23897 (N_23897,N_22099,N_22137);
nor U23898 (N_23898,N_22963,N_22349);
nor U23899 (N_23899,N_22436,N_22202);
or U23900 (N_23900,N_22735,N_22031);
nor U23901 (N_23901,N_22761,N_22808);
or U23902 (N_23902,N_22197,N_22458);
xor U23903 (N_23903,N_22366,N_22969);
or U23904 (N_23904,N_22148,N_22055);
nand U23905 (N_23905,N_22387,N_22767);
and U23906 (N_23906,N_22200,N_22868);
xor U23907 (N_23907,N_22442,N_22992);
or U23908 (N_23908,N_22579,N_22907);
or U23909 (N_23909,N_22144,N_22674);
and U23910 (N_23910,N_22397,N_22208);
or U23911 (N_23911,N_22515,N_22001);
xor U23912 (N_23912,N_22789,N_22282);
and U23913 (N_23913,N_22279,N_22203);
or U23914 (N_23914,N_22447,N_22050);
and U23915 (N_23915,N_22060,N_22963);
or U23916 (N_23916,N_22505,N_22008);
nor U23917 (N_23917,N_22894,N_22451);
and U23918 (N_23918,N_22828,N_22527);
or U23919 (N_23919,N_22602,N_22893);
and U23920 (N_23920,N_22537,N_22703);
nor U23921 (N_23921,N_22966,N_22173);
and U23922 (N_23922,N_22219,N_22580);
nor U23923 (N_23923,N_22049,N_22134);
or U23924 (N_23924,N_22490,N_22842);
nor U23925 (N_23925,N_22398,N_22687);
and U23926 (N_23926,N_22054,N_22013);
or U23927 (N_23927,N_22355,N_22621);
xor U23928 (N_23928,N_22395,N_22129);
and U23929 (N_23929,N_22627,N_22791);
or U23930 (N_23930,N_22441,N_22551);
nand U23931 (N_23931,N_22708,N_22380);
or U23932 (N_23932,N_22981,N_22488);
or U23933 (N_23933,N_22779,N_22012);
xor U23934 (N_23934,N_22311,N_22750);
xor U23935 (N_23935,N_22634,N_22513);
and U23936 (N_23936,N_22790,N_22759);
nand U23937 (N_23937,N_22564,N_22642);
or U23938 (N_23938,N_22559,N_22011);
and U23939 (N_23939,N_22185,N_22375);
and U23940 (N_23940,N_22277,N_22849);
or U23941 (N_23941,N_22309,N_22011);
and U23942 (N_23942,N_22537,N_22410);
xnor U23943 (N_23943,N_22663,N_22638);
nor U23944 (N_23944,N_22071,N_22308);
or U23945 (N_23945,N_22398,N_22842);
or U23946 (N_23946,N_22766,N_22437);
and U23947 (N_23947,N_22709,N_22297);
or U23948 (N_23948,N_22236,N_22977);
xnor U23949 (N_23949,N_22767,N_22108);
nor U23950 (N_23950,N_22946,N_22605);
and U23951 (N_23951,N_22503,N_22447);
xnor U23952 (N_23952,N_22676,N_22165);
or U23953 (N_23953,N_22229,N_22515);
nor U23954 (N_23954,N_22227,N_22004);
and U23955 (N_23955,N_22725,N_22926);
and U23956 (N_23956,N_22880,N_22637);
xnor U23957 (N_23957,N_22901,N_22057);
or U23958 (N_23958,N_22105,N_22408);
nor U23959 (N_23959,N_22874,N_22880);
or U23960 (N_23960,N_22769,N_22458);
and U23961 (N_23961,N_22850,N_22367);
nor U23962 (N_23962,N_22582,N_22149);
and U23963 (N_23963,N_22251,N_22451);
xor U23964 (N_23964,N_22603,N_22397);
nand U23965 (N_23965,N_22308,N_22494);
nor U23966 (N_23966,N_22318,N_22565);
and U23967 (N_23967,N_22609,N_22336);
and U23968 (N_23968,N_22586,N_22605);
xnor U23969 (N_23969,N_22568,N_22068);
nor U23970 (N_23970,N_22967,N_22496);
nand U23971 (N_23971,N_22648,N_22682);
nor U23972 (N_23972,N_22240,N_22075);
and U23973 (N_23973,N_22267,N_22387);
or U23974 (N_23974,N_22489,N_22741);
and U23975 (N_23975,N_22863,N_22065);
or U23976 (N_23976,N_22987,N_22771);
or U23977 (N_23977,N_22139,N_22514);
nand U23978 (N_23978,N_22463,N_22744);
nor U23979 (N_23979,N_22647,N_22710);
nor U23980 (N_23980,N_22964,N_22633);
or U23981 (N_23981,N_22703,N_22991);
nand U23982 (N_23982,N_22422,N_22580);
nand U23983 (N_23983,N_22819,N_22145);
or U23984 (N_23984,N_22838,N_22270);
or U23985 (N_23985,N_22894,N_22201);
nand U23986 (N_23986,N_22956,N_22677);
nor U23987 (N_23987,N_22239,N_22004);
and U23988 (N_23988,N_22761,N_22664);
nor U23989 (N_23989,N_22144,N_22581);
and U23990 (N_23990,N_22542,N_22460);
nand U23991 (N_23991,N_22440,N_22607);
xnor U23992 (N_23992,N_22109,N_22490);
nor U23993 (N_23993,N_22977,N_22468);
nand U23994 (N_23994,N_22746,N_22930);
xnor U23995 (N_23995,N_22718,N_22517);
and U23996 (N_23996,N_22651,N_22723);
xor U23997 (N_23997,N_22936,N_22690);
xor U23998 (N_23998,N_22955,N_22407);
or U23999 (N_23999,N_22368,N_22224);
or U24000 (N_24000,N_23389,N_23862);
nand U24001 (N_24001,N_23962,N_23296);
or U24002 (N_24002,N_23416,N_23275);
xor U24003 (N_24003,N_23395,N_23852);
nor U24004 (N_24004,N_23387,N_23298);
or U24005 (N_24005,N_23950,N_23163);
or U24006 (N_24006,N_23767,N_23727);
or U24007 (N_24007,N_23044,N_23219);
xor U24008 (N_24008,N_23685,N_23015);
or U24009 (N_24009,N_23051,N_23064);
and U24010 (N_24010,N_23789,N_23142);
nor U24011 (N_24011,N_23835,N_23990);
and U24012 (N_24012,N_23761,N_23354);
nand U24013 (N_24013,N_23877,N_23840);
xor U24014 (N_24014,N_23363,N_23755);
xnor U24015 (N_24015,N_23763,N_23650);
nor U24016 (N_24016,N_23826,N_23057);
nand U24017 (N_24017,N_23979,N_23252);
nand U24018 (N_24018,N_23831,N_23579);
or U24019 (N_24019,N_23312,N_23381);
or U24020 (N_24020,N_23746,N_23666);
nand U24021 (N_24021,N_23527,N_23739);
or U24022 (N_24022,N_23589,N_23616);
xnor U24023 (N_24023,N_23654,N_23683);
and U24024 (N_24024,N_23211,N_23350);
or U24025 (N_24025,N_23580,N_23166);
and U24026 (N_24026,N_23251,N_23138);
nor U24027 (N_24027,N_23472,N_23720);
nor U24028 (N_24028,N_23817,N_23897);
or U24029 (N_24029,N_23823,N_23022);
or U24030 (N_24030,N_23906,N_23581);
nor U24031 (N_24031,N_23006,N_23253);
nand U24032 (N_24032,N_23286,N_23262);
nand U24033 (N_24033,N_23490,N_23200);
nand U24034 (N_24034,N_23038,N_23427);
nor U24035 (N_24035,N_23300,N_23629);
and U24036 (N_24036,N_23222,N_23775);
nor U24037 (N_24037,N_23773,N_23317);
xor U24038 (N_24038,N_23738,N_23446);
nor U24039 (N_24039,N_23807,N_23541);
nand U24040 (N_24040,N_23788,N_23287);
or U24041 (N_24041,N_23443,N_23011);
nand U24042 (N_24042,N_23643,N_23682);
nand U24043 (N_24043,N_23938,N_23343);
or U24044 (N_24044,N_23434,N_23543);
and U24045 (N_24045,N_23456,N_23503);
xor U24046 (N_24046,N_23876,N_23139);
xnor U24047 (N_24047,N_23491,N_23315);
or U24048 (N_24048,N_23153,N_23610);
nand U24049 (N_24049,N_23230,N_23644);
or U24050 (N_24050,N_23124,N_23680);
xnor U24051 (N_24051,N_23658,N_23393);
and U24052 (N_24052,N_23694,N_23929);
or U24053 (N_24053,N_23321,N_23220);
or U24054 (N_24054,N_23168,N_23570);
or U24055 (N_24055,N_23645,N_23417);
and U24056 (N_24056,N_23040,N_23511);
or U24057 (N_24057,N_23132,N_23041);
nor U24058 (N_24058,N_23633,N_23954);
or U24059 (N_24059,N_23690,N_23035);
or U24060 (N_24060,N_23802,N_23554);
xor U24061 (N_24061,N_23029,N_23195);
or U24062 (N_24062,N_23236,N_23249);
nand U24063 (N_24063,N_23401,N_23391);
xor U24064 (N_24064,N_23159,N_23608);
nand U24065 (N_24065,N_23677,N_23901);
xor U24066 (N_24066,N_23282,N_23707);
and U24067 (N_24067,N_23146,N_23357);
xnor U24068 (N_24068,N_23538,N_23463);
or U24069 (N_24069,N_23425,N_23593);
and U24070 (N_24070,N_23127,N_23697);
and U24071 (N_24071,N_23001,N_23246);
xor U24072 (N_24072,N_23973,N_23803);
and U24073 (N_24073,N_23323,N_23989);
nand U24074 (N_24074,N_23367,N_23301);
xor U24075 (N_24075,N_23382,N_23325);
nor U24076 (N_24076,N_23705,N_23488);
xnor U24077 (N_24077,N_23829,N_23477);
and U24078 (N_24078,N_23194,N_23234);
xor U24079 (N_24079,N_23742,N_23936);
xor U24080 (N_24080,N_23276,N_23261);
and U24081 (N_24081,N_23945,N_23341);
nand U24082 (N_24082,N_23749,N_23157);
nand U24083 (N_24083,N_23713,N_23948);
xor U24084 (N_24084,N_23576,N_23624);
nor U24085 (N_24085,N_23991,N_23602);
xor U24086 (N_24086,N_23806,N_23167);
nor U24087 (N_24087,N_23328,N_23724);
xor U24088 (N_24088,N_23759,N_23953);
xnor U24089 (N_24089,N_23704,N_23860);
or U24090 (N_24090,N_23519,N_23055);
or U24091 (N_24091,N_23218,N_23320);
nand U24092 (N_24092,N_23059,N_23052);
nor U24093 (N_24093,N_23304,N_23465);
nand U24094 (N_24094,N_23113,N_23451);
and U24095 (N_24095,N_23760,N_23797);
and U24096 (N_24096,N_23182,N_23088);
or U24097 (N_24097,N_23319,N_23747);
nor U24098 (N_24098,N_23787,N_23856);
nand U24099 (N_24099,N_23444,N_23932);
nand U24100 (N_24100,N_23708,N_23410);
and U24101 (N_24101,N_23104,N_23118);
or U24102 (N_24102,N_23732,N_23611);
nor U24103 (N_24103,N_23668,N_23617);
and U24104 (N_24104,N_23965,N_23696);
nor U24105 (N_24105,N_23635,N_23984);
nand U24106 (N_24106,N_23597,N_23330);
xnor U24107 (N_24107,N_23303,N_23657);
nor U24108 (N_24108,N_23116,N_23332);
nor U24109 (N_24109,N_23480,N_23891);
nand U24110 (N_24110,N_23148,N_23756);
xnor U24111 (N_24111,N_23333,N_23196);
and U24112 (N_24112,N_23865,N_23562);
and U24113 (N_24113,N_23499,N_23368);
and U24114 (N_24114,N_23385,N_23125);
xnor U24115 (N_24115,N_23339,N_23086);
nor U24116 (N_24116,N_23032,N_23620);
nand U24117 (N_24117,N_23069,N_23378);
nand U24118 (N_24118,N_23075,N_23178);
nor U24119 (N_24119,N_23447,N_23590);
nand U24120 (N_24120,N_23625,N_23497);
or U24121 (N_24121,N_23937,N_23008);
xnor U24122 (N_24122,N_23873,N_23245);
nor U24123 (N_24123,N_23437,N_23049);
or U24124 (N_24124,N_23294,N_23054);
or U24125 (N_24125,N_23946,N_23264);
xnor U24126 (N_24126,N_23248,N_23729);
nor U24127 (N_24127,N_23288,N_23476);
and U24128 (N_24128,N_23693,N_23914);
xnor U24129 (N_24129,N_23295,N_23846);
or U24130 (N_24130,N_23943,N_23553);
xnor U24131 (N_24131,N_23013,N_23719);
xor U24132 (N_24132,N_23436,N_23723);
nor U24133 (N_24133,N_23801,N_23675);
nor U24134 (N_24134,N_23237,N_23297);
nand U24135 (N_24135,N_23386,N_23688);
xor U24136 (N_24136,N_23710,N_23165);
nor U24137 (N_24137,N_23601,N_23868);
nor U24138 (N_24138,N_23795,N_23867);
nand U24139 (N_24139,N_23047,N_23291);
nor U24140 (N_24140,N_23569,N_23875);
nand U24141 (N_24141,N_23213,N_23784);
nand U24142 (N_24142,N_23671,N_23808);
nor U24143 (N_24143,N_23709,N_23575);
or U24144 (N_24144,N_23703,N_23306);
nor U24145 (N_24145,N_23772,N_23383);
xor U24146 (N_24146,N_23985,N_23435);
and U24147 (N_24147,N_23641,N_23560);
nor U24148 (N_24148,N_23370,N_23796);
and U24149 (N_24149,N_23198,N_23440);
nor U24150 (N_24150,N_23799,N_23878);
nor U24151 (N_24151,N_23670,N_23818);
nor U24152 (N_24152,N_23966,N_23266);
nand U24153 (N_24153,N_23004,N_23563);
or U24154 (N_24154,N_23986,N_23618);
xnor U24155 (N_24155,N_23505,N_23882);
and U24156 (N_24156,N_23971,N_23056);
nand U24157 (N_24157,N_23764,N_23250);
nor U24158 (N_24158,N_23176,N_23058);
nor U24159 (N_24159,N_23769,N_23949);
or U24160 (N_24160,N_23905,N_23825);
and U24161 (N_24161,N_23552,N_23702);
or U24162 (N_24162,N_23335,N_23407);
nor U24163 (N_24163,N_23183,N_23881);
nor U24164 (N_24164,N_23130,N_23374);
nand U24165 (N_24165,N_23507,N_23631);
or U24166 (N_24166,N_23115,N_23811);
nor U24167 (N_24167,N_23351,N_23915);
and U24168 (N_24168,N_23596,N_23980);
xor U24169 (N_24169,N_23197,N_23030);
nor U24170 (N_24170,N_23981,N_23924);
and U24171 (N_24171,N_23455,N_23508);
xor U24172 (N_24172,N_23923,N_23396);
xor U24173 (N_24173,N_23655,N_23963);
nand U24174 (N_24174,N_23174,N_23672);
nor U24175 (N_24175,N_23947,N_23571);
xnor U24176 (N_24176,N_23336,N_23184);
xor U24177 (N_24177,N_23564,N_23212);
xnor U24178 (N_24178,N_23762,N_23091);
xnor U24179 (N_24179,N_23819,N_23096);
or U24180 (N_24180,N_23090,N_23585);
nand U24181 (N_24181,N_23186,N_23513);
or U24182 (N_24182,N_23942,N_23689);
nand U24183 (N_24183,N_23718,N_23352);
xnor U24184 (N_24184,N_23952,N_23827);
nand U24185 (N_24185,N_23170,N_23050);
nor U24186 (N_24186,N_23957,N_23861);
nor U24187 (N_24187,N_23036,N_23140);
nand U24188 (N_24188,N_23793,N_23510);
xnor U24189 (N_24189,N_23630,N_23667);
and U24190 (N_24190,N_23814,N_23886);
nand U24191 (N_24191,N_23838,N_23893);
nor U24192 (N_24192,N_23310,N_23398);
xor U24193 (N_24193,N_23229,N_23975);
nor U24194 (N_24194,N_23175,N_23782);
or U24195 (N_24195,N_23226,N_23375);
nand U24196 (N_24196,N_23518,N_23792);
and U24197 (N_24197,N_23372,N_23686);
or U24198 (N_24198,N_23565,N_23016);
and U24199 (N_24199,N_23334,N_23376);
and U24200 (N_24200,N_23123,N_23384);
nor U24201 (N_24201,N_23223,N_23752);
nand U24202 (N_24202,N_23969,N_23337);
nand U24203 (N_24203,N_23774,N_23870);
or U24204 (N_24204,N_23780,N_23885);
or U24205 (N_24205,N_23895,N_23520);
or U24206 (N_24206,N_23639,N_23421);
or U24207 (N_24207,N_23545,N_23445);
xor U24208 (N_24208,N_23257,N_23344);
xnor U24209 (N_24209,N_23745,N_23740);
nand U24210 (N_24210,N_23208,N_23765);
or U24211 (N_24211,N_23149,N_23781);
nand U24212 (N_24212,N_23516,N_23135);
xor U24213 (N_24213,N_23299,N_23105);
or U24214 (N_24214,N_23485,N_23327);
nor U24215 (N_24215,N_23626,N_23144);
nand U24216 (N_24216,N_23449,N_23786);
nand U24217 (N_24217,N_23837,N_23632);
xor U24218 (N_24218,N_23857,N_23768);
nor U24219 (N_24219,N_23623,N_23804);
or U24220 (N_24220,N_23272,N_23646);
nand U24221 (N_24221,N_23188,N_23173);
xor U24222 (N_24222,N_23240,N_23152);
nand U24223 (N_24223,N_23479,N_23995);
xor U24224 (N_24224,N_23441,N_23627);
and U24225 (N_24225,N_23892,N_23241);
and U24226 (N_24226,N_23400,N_23959);
and U24227 (N_24227,N_23664,N_23235);
nor U24228 (N_24228,N_23730,N_23528);
xnor U24229 (N_24229,N_23190,N_23369);
or U24230 (N_24230,N_23031,N_23869);
xnor U24231 (N_24231,N_23504,N_23353);
or U24232 (N_24232,N_23100,N_23120);
and U24233 (N_24233,N_23087,N_23277);
xnor U24234 (N_24234,N_23033,N_23854);
and U24235 (N_24235,N_23753,N_23813);
and U24236 (N_24236,N_23556,N_23996);
or U24237 (N_24237,N_23907,N_23547);
or U24238 (N_24238,N_23551,N_23733);
and U24239 (N_24239,N_23018,N_23207);
nor U24240 (N_24240,N_23592,N_23815);
xnor U24241 (N_24241,N_23656,N_23955);
nor U24242 (N_24242,N_23874,N_23619);
and U24243 (N_24243,N_23659,N_23107);
nor U24244 (N_24244,N_23637,N_23439);
nor U24245 (N_24245,N_23524,N_23177);
or U24246 (N_24246,N_23478,N_23648);
xor U24247 (N_24247,N_23487,N_23598);
and U24248 (N_24248,N_23758,N_23077);
xor U24249 (N_24249,N_23506,N_23082);
xor U24250 (N_24250,N_23968,N_23380);
or U24251 (N_24251,N_23314,N_23572);
or U24252 (N_24252,N_23063,N_23422);
nand U24253 (N_24253,N_23512,N_23413);
xnor U24254 (N_24254,N_23308,N_23322);
or U24255 (N_24255,N_23366,N_23928);
nand U24256 (N_24256,N_23475,N_23536);
nor U24257 (N_24257,N_23271,N_23855);
nor U24258 (N_24258,N_23360,N_23238);
and U24259 (N_24259,N_23070,N_23992);
xor U24260 (N_24260,N_23509,N_23150);
or U24261 (N_24261,N_23399,N_23482);
and U24262 (N_24262,N_23028,N_23112);
nor U24263 (N_24263,N_23956,N_23205);
nand U24264 (N_24264,N_23215,N_23798);
xor U24265 (N_24265,N_23607,N_23158);
and U24266 (N_24266,N_23883,N_23530);
nor U24267 (N_24267,N_23859,N_23525);
nand U24268 (N_24268,N_23599,N_23734);
nand U24269 (N_24269,N_23181,N_23092);
xor U24270 (N_24270,N_23279,N_23824);
nand U24271 (N_24271,N_23089,N_23448);
and U24272 (N_24272,N_23588,N_23459);
nor U24273 (N_24273,N_23858,N_23866);
and U24274 (N_24274,N_23024,N_23548);
nor U24275 (N_24275,N_23757,N_23160);
nand U24276 (N_24276,N_23532,N_23843);
nor U24277 (N_24277,N_23392,N_23609);
and U24278 (N_24278,N_23900,N_23429);
and U24279 (N_24279,N_23539,N_23326);
nor U24280 (N_24280,N_23199,N_23841);
nand U24281 (N_24281,N_23910,N_23430);
nand U24282 (N_24282,N_23162,N_23974);
and U24283 (N_24283,N_23231,N_23483);
or U24284 (N_24284,N_23404,N_23978);
or U24285 (N_24285,N_23243,N_23192);
and U24286 (N_24286,N_23566,N_23102);
xnor U24287 (N_24287,N_23678,N_23676);
nand U24288 (N_24288,N_23529,N_23591);
or U24289 (N_24289,N_23023,N_23958);
or U24290 (N_24290,N_23342,N_23106);
xnor U24291 (N_24291,N_23373,N_23716);
and U24292 (N_24292,N_23982,N_23048);
nor U24293 (N_24293,N_23292,N_23085);
nor U24294 (N_24294,N_23486,N_23239);
nor U24295 (N_24295,N_23642,N_23154);
and U24296 (N_24296,N_23256,N_23636);
and U24297 (N_24297,N_23406,N_23894);
and U24298 (N_24298,N_23833,N_23573);
nand U24299 (N_24299,N_23390,N_23555);
and U24300 (N_24300,N_23331,N_23695);
xnor U24301 (N_24301,N_23791,N_23535);
or U24302 (N_24302,N_23805,N_23358);
nand U24303 (N_24303,N_23426,N_23584);
nor U24304 (N_24304,N_23533,N_23045);
xnor U24305 (N_24305,N_23103,N_23832);
nor U24306 (N_24306,N_23133,N_23498);
xor U24307 (N_24307,N_23462,N_23501);
or U24308 (N_24308,N_23293,N_23042);
and U24309 (N_24309,N_23233,N_23081);
and U24310 (N_24310,N_23839,N_23109);
nand U24311 (N_24311,N_23419,N_23290);
xnor U24312 (N_24312,N_23021,N_23779);
or U24313 (N_24313,N_23468,N_23951);
or U24314 (N_24314,N_23364,N_23020);
nor U24315 (N_24315,N_23987,N_23647);
and U24316 (N_24316,N_23534,N_23771);
or U24317 (N_24317,N_23717,N_23141);
nand U24318 (N_24318,N_23776,N_23442);
or U24319 (N_24319,N_23423,N_23848);
or U24320 (N_24320,N_23638,N_23681);
and U24321 (N_24321,N_23076,N_23691);
xnor U24322 (N_24322,N_23122,N_23496);
xnor U24323 (N_24323,N_23994,N_23930);
or U24324 (N_24324,N_23414,N_23522);
nor U24325 (N_24325,N_23000,N_23884);
and U24326 (N_24326,N_23349,N_23114);
or U24327 (N_24327,N_23921,N_23466);
xnor U24328 (N_24328,N_23108,N_23202);
nor U24329 (N_24329,N_23454,N_23822);
or U24330 (N_24330,N_23471,N_23898);
xnor U24331 (N_24331,N_23844,N_23889);
or U24332 (N_24332,N_23777,N_23922);
nor U24333 (N_24333,N_23722,N_23228);
nor U24334 (N_24334,N_23067,N_23415);
or U24335 (N_24335,N_23544,N_23428);
xor U24336 (N_24336,N_23568,N_23830);
and U24337 (N_24337,N_23467,N_23613);
nand U24338 (N_24338,N_23934,N_23692);
and U24339 (N_24339,N_23080,N_23281);
nand U24340 (N_24340,N_23143,N_23359);
nor U24341 (N_24341,N_23595,N_23706);
and U24342 (N_24342,N_23071,N_23003);
xnor U24343 (N_24343,N_23715,N_23880);
nand U24344 (N_24344,N_23347,N_23227);
or U24345 (N_24345,N_23871,N_23816);
and U24346 (N_24346,N_23721,N_23098);
xnor U24347 (N_24347,N_23621,N_23517);
or U24348 (N_24348,N_23210,N_23812);
and U24349 (N_24349,N_23604,N_23450);
and U24350 (N_24350,N_23136,N_23944);
or U24351 (N_24351,N_23268,N_23134);
nor U24352 (N_24352,N_23318,N_23411);
nand U24353 (N_24353,N_23362,N_23699);
xor U24354 (N_24354,N_23302,N_23976);
xor U24355 (N_24355,N_23917,N_23131);
and U24356 (N_24356,N_23743,N_23927);
nor U24357 (N_24357,N_23244,N_23864);
nor U24358 (N_24358,N_23156,N_23043);
and U24359 (N_24359,N_23918,N_23999);
xnor U24360 (N_24360,N_23770,N_23684);
xor U24361 (N_24361,N_23561,N_23495);
or U24362 (N_24362,N_23255,N_23967);
xnor U24363 (N_24363,N_23307,N_23014);
nand U24364 (N_24364,N_23171,N_23484);
nand U24365 (N_24365,N_23649,N_23099);
and U24366 (N_24366,N_23735,N_23094);
nor U24367 (N_24367,N_23204,N_23515);
and U24368 (N_24368,N_23260,N_23540);
and U24369 (N_24369,N_23217,N_23305);
nand U24370 (N_24370,N_23010,N_23101);
nor U24371 (N_24371,N_23567,N_23800);
and U24372 (N_24372,N_23725,N_23652);
nand U24373 (N_24373,N_23007,N_23850);
xnor U24374 (N_24374,N_23845,N_23500);
nor U24375 (N_24375,N_23203,N_23606);
xor U24376 (N_24376,N_23377,N_23418);
xor U24377 (N_24377,N_23474,N_23265);
or U24378 (N_24378,N_23053,N_23909);
or U24379 (N_24379,N_23469,N_23842);
nor U24380 (N_24380,N_23698,N_23438);
nor U24381 (N_24381,N_23062,N_23066);
nor U24382 (N_24382,N_23324,N_23461);
nand U24383 (N_24383,N_23521,N_23887);
nand U24384 (N_24384,N_23285,N_23037);
nand U24385 (N_24385,N_23674,N_23065);
xnor U24386 (N_24386,N_23026,N_23494);
xor U24387 (N_24387,N_23258,N_23712);
or U24388 (N_24388,N_23577,N_23514);
nand U24389 (N_24389,N_23888,N_23221);
and U24390 (N_24390,N_23179,N_23458);
or U24391 (N_24391,N_23612,N_23005);
or U24392 (N_24392,N_23111,N_23214);
nand U24393 (N_24393,N_23432,N_23269);
xnor U24394 (N_24394,N_23820,N_23559);
nand U24395 (N_24395,N_23397,N_23361);
and U24396 (N_24396,N_23473,N_23919);
or U24397 (N_24397,N_23460,N_23232);
or U24398 (N_24398,N_23651,N_23964);
xnor U24399 (N_24399,N_23983,N_23126);
nor U24400 (N_24400,N_23110,N_23206);
xnor U24401 (N_24401,N_23941,N_23673);
nand U24402 (N_24402,N_23828,N_23169);
nand U24403 (N_24403,N_23481,N_23821);
nor U24404 (N_24404,N_23492,N_23464);
or U24405 (N_24405,N_23750,N_23201);
nor U24406 (N_24406,N_23316,N_23574);
xor U24407 (N_24407,N_23270,N_23714);
nor U24408 (N_24408,N_23961,N_23355);
and U24409 (N_24409,N_23640,N_23039);
nor U24410 (N_24410,N_23977,N_23209);
nor U24411 (N_24411,N_23879,N_23736);
or U24412 (N_24412,N_23453,N_23216);
xor U24413 (N_24413,N_23557,N_23379);
nor U24414 (N_24414,N_23172,N_23603);
and U24415 (N_24415,N_23913,N_23371);
and U24416 (N_24416,N_23145,N_23412);
nor U24417 (N_24417,N_23084,N_23147);
and U24418 (N_24418,N_23117,N_23726);
or U24419 (N_24419,N_23810,N_23161);
xnor U24420 (N_24420,N_23155,N_23939);
nand U24421 (N_24421,N_23970,N_23072);
xnor U24422 (N_24422,N_23558,N_23653);
xor U24423 (N_24423,N_23017,N_23549);
or U24424 (N_24424,N_23283,N_23034);
xor U24425 (N_24425,N_23263,N_23701);
and U24426 (N_24426,N_23002,N_23537);
and U24427 (N_24427,N_23502,N_23079);
xnor U24428 (N_24428,N_23687,N_23225);
xor U24429 (N_24429,N_23960,N_23600);
xor U24430 (N_24430,N_23899,N_23311);
nand U24431 (N_24431,N_23766,N_23546);
and U24432 (N_24432,N_23409,N_23849);
and U24433 (N_24433,N_23137,N_23912);
nand U24434 (N_24434,N_23151,N_23457);
nand U24435 (N_24435,N_23242,N_23911);
or U24436 (N_24436,N_23920,N_23452);
nor U24437 (N_24437,N_23073,N_23634);
nor U24438 (N_24438,N_23908,N_23700);
and U24439 (N_24439,N_23289,N_23836);
nand U24440 (N_24440,N_23345,N_23313);
or U24441 (N_24441,N_23904,N_23489);
or U24442 (N_24442,N_23129,N_23737);
and U24443 (N_24443,N_23189,N_23185);
nor U24444 (N_24444,N_23273,N_23594);
nand U24445 (N_24445,N_23046,N_23744);
xnor U24446 (N_24446,N_23025,N_23420);
nor U24447 (N_24447,N_23346,N_23550);
nand U24448 (N_24448,N_23662,N_23931);
nor U24449 (N_24449,N_23794,N_23403);
nor U24450 (N_24450,N_23863,N_23180);
and U24451 (N_24451,N_23078,N_23587);
xnor U24452 (N_24452,N_23061,N_23348);
nor U24453 (N_24453,N_23128,N_23164);
or U24454 (N_24454,N_23402,N_23972);
xor U24455 (N_24455,N_23997,N_23661);
or U24456 (N_24456,N_23728,N_23224);
and U24457 (N_24457,N_23405,N_23582);
and U24458 (N_24458,N_23778,N_23068);
or U24459 (N_24459,N_23365,N_23338);
xor U24460 (N_24460,N_23083,N_23935);
nand U24461 (N_24461,N_23526,N_23916);
and U24462 (N_24462,N_23431,N_23748);
or U24463 (N_24463,N_23902,N_23191);
nand U24464 (N_24464,N_23284,N_23340);
nor U24465 (N_24465,N_23896,N_23267);
nand U24466 (N_24466,N_23940,N_23586);
nor U24467 (N_24467,N_23847,N_23993);
and U24468 (N_24468,N_23009,N_23388);
nor U24469 (N_24469,N_23097,N_23998);
and U24470 (N_24470,N_23711,N_23925);
and U24471 (N_24471,N_23628,N_23027);
nand U24472 (N_24472,N_23060,N_23663);
xor U24473 (N_24473,N_23622,N_23278);
nand U24474 (N_24474,N_23309,N_23988);
xnor U24475 (N_24475,N_23751,N_23853);
xnor U24476 (N_24476,N_23121,N_23119);
nor U24477 (N_24477,N_23274,N_23809);
or U24478 (N_24478,N_23433,N_23731);
and U24479 (N_24479,N_23424,N_23523);
or U24480 (N_24480,N_23679,N_23741);
nor U24481 (N_24481,N_23254,N_23259);
and U24482 (N_24482,N_23890,N_23903);
nand U24483 (N_24483,N_23093,N_23785);
nor U24484 (N_24484,N_23790,N_23665);
nand U24485 (N_24485,N_23531,N_23280);
xor U24486 (N_24486,N_23019,N_23394);
xor U24487 (N_24487,N_23660,N_23933);
nor U24488 (N_24488,N_23605,N_23408);
nor U24489 (N_24489,N_23851,N_23834);
nand U24490 (N_24490,N_23095,N_23356);
nand U24491 (N_24491,N_23872,N_23754);
and U24492 (N_24492,N_23187,N_23470);
or U24493 (N_24493,N_23614,N_23783);
xnor U24494 (N_24494,N_23583,N_23193);
and U24495 (N_24495,N_23926,N_23247);
xor U24496 (N_24496,N_23615,N_23493);
and U24497 (N_24497,N_23542,N_23578);
and U24498 (N_24498,N_23669,N_23074);
or U24499 (N_24499,N_23329,N_23012);
nor U24500 (N_24500,N_23092,N_23682);
nor U24501 (N_24501,N_23172,N_23538);
or U24502 (N_24502,N_23201,N_23223);
xnor U24503 (N_24503,N_23980,N_23999);
or U24504 (N_24504,N_23071,N_23465);
xnor U24505 (N_24505,N_23134,N_23506);
and U24506 (N_24506,N_23641,N_23084);
xor U24507 (N_24507,N_23860,N_23745);
or U24508 (N_24508,N_23236,N_23375);
and U24509 (N_24509,N_23151,N_23987);
and U24510 (N_24510,N_23015,N_23069);
xnor U24511 (N_24511,N_23827,N_23846);
and U24512 (N_24512,N_23139,N_23526);
xor U24513 (N_24513,N_23169,N_23359);
and U24514 (N_24514,N_23039,N_23985);
nor U24515 (N_24515,N_23159,N_23665);
xnor U24516 (N_24516,N_23634,N_23704);
and U24517 (N_24517,N_23449,N_23881);
and U24518 (N_24518,N_23057,N_23005);
and U24519 (N_24519,N_23951,N_23117);
nor U24520 (N_24520,N_23757,N_23025);
and U24521 (N_24521,N_23718,N_23675);
or U24522 (N_24522,N_23535,N_23454);
and U24523 (N_24523,N_23622,N_23356);
or U24524 (N_24524,N_23660,N_23212);
and U24525 (N_24525,N_23155,N_23334);
or U24526 (N_24526,N_23640,N_23502);
nand U24527 (N_24527,N_23638,N_23348);
and U24528 (N_24528,N_23052,N_23817);
xor U24529 (N_24529,N_23405,N_23409);
and U24530 (N_24530,N_23444,N_23963);
nand U24531 (N_24531,N_23804,N_23930);
and U24532 (N_24532,N_23903,N_23158);
nor U24533 (N_24533,N_23810,N_23656);
xor U24534 (N_24534,N_23759,N_23849);
xnor U24535 (N_24535,N_23445,N_23656);
or U24536 (N_24536,N_23902,N_23772);
and U24537 (N_24537,N_23989,N_23058);
xnor U24538 (N_24538,N_23697,N_23669);
nand U24539 (N_24539,N_23418,N_23280);
nand U24540 (N_24540,N_23746,N_23010);
nor U24541 (N_24541,N_23875,N_23472);
and U24542 (N_24542,N_23641,N_23337);
nand U24543 (N_24543,N_23251,N_23749);
and U24544 (N_24544,N_23442,N_23809);
nor U24545 (N_24545,N_23799,N_23700);
nor U24546 (N_24546,N_23813,N_23088);
xnor U24547 (N_24547,N_23778,N_23368);
nor U24548 (N_24548,N_23274,N_23679);
nand U24549 (N_24549,N_23534,N_23317);
nand U24550 (N_24550,N_23571,N_23979);
or U24551 (N_24551,N_23502,N_23174);
xnor U24552 (N_24552,N_23561,N_23537);
nor U24553 (N_24553,N_23220,N_23807);
nand U24554 (N_24554,N_23000,N_23565);
nor U24555 (N_24555,N_23891,N_23622);
nand U24556 (N_24556,N_23820,N_23836);
nor U24557 (N_24557,N_23478,N_23249);
and U24558 (N_24558,N_23899,N_23904);
xnor U24559 (N_24559,N_23208,N_23917);
xor U24560 (N_24560,N_23716,N_23287);
nor U24561 (N_24561,N_23718,N_23392);
nand U24562 (N_24562,N_23008,N_23615);
nor U24563 (N_24563,N_23185,N_23758);
nand U24564 (N_24564,N_23654,N_23168);
and U24565 (N_24565,N_23503,N_23090);
and U24566 (N_24566,N_23518,N_23617);
or U24567 (N_24567,N_23573,N_23670);
or U24568 (N_24568,N_23485,N_23280);
or U24569 (N_24569,N_23948,N_23581);
or U24570 (N_24570,N_23013,N_23607);
xor U24571 (N_24571,N_23948,N_23174);
xnor U24572 (N_24572,N_23477,N_23095);
nand U24573 (N_24573,N_23082,N_23174);
nand U24574 (N_24574,N_23011,N_23904);
and U24575 (N_24575,N_23085,N_23274);
nor U24576 (N_24576,N_23096,N_23516);
and U24577 (N_24577,N_23141,N_23796);
nand U24578 (N_24578,N_23660,N_23032);
nor U24579 (N_24579,N_23733,N_23713);
nand U24580 (N_24580,N_23263,N_23936);
xnor U24581 (N_24581,N_23748,N_23900);
or U24582 (N_24582,N_23339,N_23858);
nand U24583 (N_24583,N_23273,N_23123);
nor U24584 (N_24584,N_23611,N_23089);
or U24585 (N_24585,N_23902,N_23560);
nor U24586 (N_24586,N_23740,N_23322);
and U24587 (N_24587,N_23469,N_23336);
xnor U24588 (N_24588,N_23148,N_23940);
or U24589 (N_24589,N_23754,N_23091);
nor U24590 (N_24590,N_23219,N_23199);
xor U24591 (N_24591,N_23811,N_23867);
nand U24592 (N_24592,N_23491,N_23159);
nor U24593 (N_24593,N_23340,N_23120);
and U24594 (N_24594,N_23428,N_23293);
nand U24595 (N_24595,N_23714,N_23782);
nor U24596 (N_24596,N_23014,N_23827);
nor U24597 (N_24597,N_23071,N_23661);
or U24598 (N_24598,N_23732,N_23469);
nand U24599 (N_24599,N_23811,N_23107);
or U24600 (N_24600,N_23589,N_23244);
or U24601 (N_24601,N_23245,N_23616);
and U24602 (N_24602,N_23459,N_23335);
nand U24603 (N_24603,N_23474,N_23968);
nor U24604 (N_24604,N_23784,N_23950);
and U24605 (N_24605,N_23525,N_23926);
nor U24606 (N_24606,N_23299,N_23887);
nor U24607 (N_24607,N_23920,N_23386);
and U24608 (N_24608,N_23147,N_23236);
nand U24609 (N_24609,N_23321,N_23999);
nand U24610 (N_24610,N_23780,N_23131);
and U24611 (N_24611,N_23689,N_23181);
nand U24612 (N_24612,N_23027,N_23572);
or U24613 (N_24613,N_23107,N_23407);
or U24614 (N_24614,N_23434,N_23372);
nor U24615 (N_24615,N_23702,N_23322);
and U24616 (N_24616,N_23222,N_23687);
and U24617 (N_24617,N_23540,N_23996);
and U24618 (N_24618,N_23622,N_23917);
xor U24619 (N_24619,N_23940,N_23971);
and U24620 (N_24620,N_23389,N_23145);
nor U24621 (N_24621,N_23037,N_23655);
xnor U24622 (N_24622,N_23968,N_23522);
nor U24623 (N_24623,N_23224,N_23543);
and U24624 (N_24624,N_23590,N_23010);
or U24625 (N_24625,N_23099,N_23140);
nor U24626 (N_24626,N_23713,N_23901);
or U24627 (N_24627,N_23102,N_23663);
and U24628 (N_24628,N_23125,N_23483);
and U24629 (N_24629,N_23627,N_23347);
xor U24630 (N_24630,N_23384,N_23521);
and U24631 (N_24631,N_23743,N_23040);
nand U24632 (N_24632,N_23786,N_23800);
nand U24633 (N_24633,N_23398,N_23508);
nand U24634 (N_24634,N_23522,N_23206);
xnor U24635 (N_24635,N_23662,N_23082);
or U24636 (N_24636,N_23362,N_23840);
nor U24637 (N_24637,N_23915,N_23640);
or U24638 (N_24638,N_23022,N_23854);
nand U24639 (N_24639,N_23079,N_23663);
nor U24640 (N_24640,N_23240,N_23898);
xnor U24641 (N_24641,N_23992,N_23788);
xor U24642 (N_24642,N_23379,N_23740);
nand U24643 (N_24643,N_23900,N_23825);
or U24644 (N_24644,N_23332,N_23597);
nand U24645 (N_24645,N_23489,N_23105);
and U24646 (N_24646,N_23064,N_23703);
and U24647 (N_24647,N_23672,N_23749);
nand U24648 (N_24648,N_23913,N_23696);
xnor U24649 (N_24649,N_23302,N_23943);
and U24650 (N_24650,N_23334,N_23682);
and U24651 (N_24651,N_23797,N_23877);
or U24652 (N_24652,N_23507,N_23874);
nor U24653 (N_24653,N_23075,N_23662);
and U24654 (N_24654,N_23079,N_23829);
nand U24655 (N_24655,N_23443,N_23719);
xnor U24656 (N_24656,N_23070,N_23248);
nor U24657 (N_24657,N_23201,N_23517);
or U24658 (N_24658,N_23033,N_23163);
and U24659 (N_24659,N_23225,N_23193);
or U24660 (N_24660,N_23723,N_23777);
nor U24661 (N_24661,N_23885,N_23698);
or U24662 (N_24662,N_23806,N_23539);
xor U24663 (N_24663,N_23351,N_23568);
xnor U24664 (N_24664,N_23058,N_23089);
nand U24665 (N_24665,N_23803,N_23529);
nand U24666 (N_24666,N_23026,N_23773);
or U24667 (N_24667,N_23879,N_23443);
and U24668 (N_24668,N_23303,N_23885);
or U24669 (N_24669,N_23877,N_23423);
or U24670 (N_24670,N_23302,N_23646);
and U24671 (N_24671,N_23627,N_23747);
or U24672 (N_24672,N_23529,N_23094);
nand U24673 (N_24673,N_23138,N_23510);
and U24674 (N_24674,N_23145,N_23179);
xor U24675 (N_24675,N_23301,N_23873);
nor U24676 (N_24676,N_23616,N_23119);
nor U24677 (N_24677,N_23322,N_23840);
nor U24678 (N_24678,N_23849,N_23503);
xor U24679 (N_24679,N_23684,N_23816);
nor U24680 (N_24680,N_23941,N_23344);
nor U24681 (N_24681,N_23959,N_23058);
nor U24682 (N_24682,N_23523,N_23673);
or U24683 (N_24683,N_23871,N_23000);
nand U24684 (N_24684,N_23653,N_23298);
and U24685 (N_24685,N_23145,N_23963);
and U24686 (N_24686,N_23403,N_23326);
nand U24687 (N_24687,N_23729,N_23214);
and U24688 (N_24688,N_23643,N_23755);
or U24689 (N_24689,N_23213,N_23997);
nor U24690 (N_24690,N_23216,N_23010);
nor U24691 (N_24691,N_23660,N_23823);
xor U24692 (N_24692,N_23167,N_23420);
xnor U24693 (N_24693,N_23024,N_23161);
nand U24694 (N_24694,N_23584,N_23118);
xor U24695 (N_24695,N_23294,N_23061);
or U24696 (N_24696,N_23250,N_23920);
xor U24697 (N_24697,N_23069,N_23499);
xnor U24698 (N_24698,N_23098,N_23374);
xor U24699 (N_24699,N_23802,N_23918);
xnor U24700 (N_24700,N_23763,N_23224);
or U24701 (N_24701,N_23961,N_23111);
and U24702 (N_24702,N_23415,N_23885);
nor U24703 (N_24703,N_23913,N_23218);
nand U24704 (N_24704,N_23229,N_23364);
xnor U24705 (N_24705,N_23260,N_23218);
and U24706 (N_24706,N_23708,N_23080);
or U24707 (N_24707,N_23821,N_23951);
nand U24708 (N_24708,N_23535,N_23711);
nor U24709 (N_24709,N_23743,N_23903);
and U24710 (N_24710,N_23000,N_23698);
nor U24711 (N_24711,N_23059,N_23133);
nand U24712 (N_24712,N_23634,N_23772);
xnor U24713 (N_24713,N_23410,N_23984);
and U24714 (N_24714,N_23897,N_23732);
nor U24715 (N_24715,N_23845,N_23714);
xor U24716 (N_24716,N_23790,N_23238);
nor U24717 (N_24717,N_23087,N_23315);
xnor U24718 (N_24718,N_23110,N_23272);
nor U24719 (N_24719,N_23569,N_23351);
xnor U24720 (N_24720,N_23737,N_23320);
and U24721 (N_24721,N_23471,N_23197);
nand U24722 (N_24722,N_23405,N_23551);
and U24723 (N_24723,N_23884,N_23396);
nand U24724 (N_24724,N_23457,N_23697);
and U24725 (N_24725,N_23557,N_23399);
nand U24726 (N_24726,N_23397,N_23344);
or U24727 (N_24727,N_23064,N_23749);
nor U24728 (N_24728,N_23916,N_23986);
nor U24729 (N_24729,N_23089,N_23731);
nor U24730 (N_24730,N_23520,N_23692);
nor U24731 (N_24731,N_23179,N_23586);
or U24732 (N_24732,N_23895,N_23552);
nor U24733 (N_24733,N_23184,N_23578);
or U24734 (N_24734,N_23969,N_23297);
or U24735 (N_24735,N_23112,N_23030);
xnor U24736 (N_24736,N_23031,N_23333);
and U24737 (N_24737,N_23664,N_23180);
nand U24738 (N_24738,N_23039,N_23507);
nor U24739 (N_24739,N_23251,N_23891);
nor U24740 (N_24740,N_23281,N_23962);
and U24741 (N_24741,N_23242,N_23124);
nand U24742 (N_24742,N_23232,N_23126);
nand U24743 (N_24743,N_23075,N_23566);
and U24744 (N_24744,N_23602,N_23907);
xor U24745 (N_24745,N_23270,N_23977);
and U24746 (N_24746,N_23919,N_23173);
and U24747 (N_24747,N_23382,N_23346);
nand U24748 (N_24748,N_23872,N_23756);
xnor U24749 (N_24749,N_23540,N_23654);
and U24750 (N_24750,N_23093,N_23454);
nor U24751 (N_24751,N_23713,N_23180);
nor U24752 (N_24752,N_23957,N_23376);
xnor U24753 (N_24753,N_23063,N_23260);
nor U24754 (N_24754,N_23613,N_23630);
nor U24755 (N_24755,N_23348,N_23739);
nor U24756 (N_24756,N_23038,N_23856);
xnor U24757 (N_24757,N_23573,N_23769);
or U24758 (N_24758,N_23495,N_23206);
nor U24759 (N_24759,N_23223,N_23901);
nand U24760 (N_24760,N_23012,N_23127);
nand U24761 (N_24761,N_23163,N_23376);
nor U24762 (N_24762,N_23880,N_23464);
and U24763 (N_24763,N_23112,N_23520);
nor U24764 (N_24764,N_23873,N_23797);
and U24765 (N_24765,N_23145,N_23312);
and U24766 (N_24766,N_23704,N_23471);
and U24767 (N_24767,N_23521,N_23180);
or U24768 (N_24768,N_23423,N_23899);
and U24769 (N_24769,N_23556,N_23821);
nand U24770 (N_24770,N_23595,N_23412);
and U24771 (N_24771,N_23668,N_23341);
or U24772 (N_24772,N_23012,N_23194);
xor U24773 (N_24773,N_23525,N_23369);
and U24774 (N_24774,N_23697,N_23586);
or U24775 (N_24775,N_23496,N_23115);
and U24776 (N_24776,N_23273,N_23742);
nor U24777 (N_24777,N_23351,N_23400);
nor U24778 (N_24778,N_23043,N_23830);
or U24779 (N_24779,N_23510,N_23377);
and U24780 (N_24780,N_23984,N_23650);
xor U24781 (N_24781,N_23730,N_23445);
or U24782 (N_24782,N_23480,N_23472);
or U24783 (N_24783,N_23785,N_23124);
nor U24784 (N_24784,N_23334,N_23453);
nor U24785 (N_24785,N_23089,N_23215);
or U24786 (N_24786,N_23191,N_23751);
nand U24787 (N_24787,N_23414,N_23026);
and U24788 (N_24788,N_23341,N_23600);
nand U24789 (N_24789,N_23997,N_23012);
and U24790 (N_24790,N_23406,N_23517);
nor U24791 (N_24791,N_23662,N_23900);
or U24792 (N_24792,N_23772,N_23502);
or U24793 (N_24793,N_23113,N_23798);
or U24794 (N_24794,N_23012,N_23287);
nand U24795 (N_24795,N_23961,N_23630);
nand U24796 (N_24796,N_23228,N_23129);
and U24797 (N_24797,N_23667,N_23954);
or U24798 (N_24798,N_23393,N_23914);
and U24799 (N_24799,N_23180,N_23652);
or U24800 (N_24800,N_23228,N_23276);
nor U24801 (N_24801,N_23424,N_23873);
nand U24802 (N_24802,N_23944,N_23219);
and U24803 (N_24803,N_23901,N_23152);
nor U24804 (N_24804,N_23516,N_23918);
and U24805 (N_24805,N_23487,N_23199);
and U24806 (N_24806,N_23383,N_23421);
xor U24807 (N_24807,N_23077,N_23846);
xor U24808 (N_24808,N_23180,N_23906);
or U24809 (N_24809,N_23518,N_23650);
xnor U24810 (N_24810,N_23327,N_23297);
or U24811 (N_24811,N_23701,N_23790);
xor U24812 (N_24812,N_23266,N_23302);
and U24813 (N_24813,N_23414,N_23383);
nand U24814 (N_24814,N_23724,N_23703);
nor U24815 (N_24815,N_23816,N_23762);
and U24816 (N_24816,N_23875,N_23231);
nand U24817 (N_24817,N_23300,N_23455);
and U24818 (N_24818,N_23228,N_23918);
nand U24819 (N_24819,N_23040,N_23609);
or U24820 (N_24820,N_23526,N_23404);
nor U24821 (N_24821,N_23576,N_23661);
and U24822 (N_24822,N_23790,N_23783);
nand U24823 (N_24823,N_23501,N_23668);
and U24824 (N_24824,N_23050,N_23031);
xnor U24825 (N_24825,N_23165,N_23914);
or U24826 (N_24826,N_23547,N_23431);
or U24827 (N_24827,N_23218,N_23224);
and U24828 (N_24828,N_23519,N_23211);
or U24829 (N_24829,N_23992,N_23505);
nor U24830 (N_24830,N_23667,N_23127);
xnor U24831 (N_24831,N_23854,N_23182);
xor U24832 (N_24832,N_23218,N_23696);
nand U24833 (N_24833,N_23472,N_23370);
or U24834 (N_24834,N_23688,N_23880);
nand U24835 (N_24835,N_23324,N_23187);
nand U24836 (N_24836,N_23833,N_23053);
nor U24837 (N_24837,N_23940,N_23235);
and U24838 (N_24838,N_23424,N_23673);
nand U24839 (N_24839,N_23836,N_23149);
nor U24840 (N_24840,N_23756,N_23847);
and U24841 (N_24841,N_23472,N_23077);
nand U24842 (N_24842,N_23916,N_23527);
and U24843 (N_24843,N_23194,N_23656);
nor U24844 (N_24844,N_23217,N_23142);
nand U24845 (N_24845,N_23363,N_23676);
xnor U24846 (N_24846,N_23518,N_23321);
nand U24847 (N_24847,N_23145,N_23440);
or U24848 (N_24848,N_23511,N_23129);
nor U24849 (N_24849,N_23096,N_23699);
and U24850 (N_24850,N_23893,N_23652);
and U24851 (N_24851,N_23794,N_23528);
nand U24852 (N_24852,N_23538,N_23017);
xor U24853 (N_24853,N_23421,N_23170);
nand U24854 (N_24854,N_23604,N_23124);
or U24855 (N_24855,N_23415,N_23108);
or U24856 (N_24856,N_23387,N_23221);
nand U24857 (N_24857,N_23904,N_23942);
and U24858 (N_24858,N_23486,N_23041);
nand U24859 (N_24859,N_23768,N_23566);
or U24860 (N_24860,N_23972,N_23139);
nor U24861 (N_24861,N_23988,N_23788);
nand U24862 (N_24862,N_23909,N_23864);
and U24863 (N_24863,N_23816,N_23022);
nor U24864 (N_24864,N_23244,N_23930);
nand U24865 (N_24865,N_23587,N_23757);
nand U24866 (N_24866,N_23549,N_23736);
or U24867 (N_24867,N_23400,N_23728);
nor U24868 (N_24868,N_23131,N_23781);
nand U24869 (N_24869,N_23592,N_23046);
xor U24870 (N_24870,N_23443,N_23185);
and U24871 (N_24871,N_23093,N_23064);
nor U24872 (N_24872,N_23240,N_23661);
nor U24873 (N_24873,N_23798,N_23229);
nor U24874 (N_24874,N_23970,N_23792);
or U24875 (N_24875,N_23763,N_23860);
nor U24876 (N_24876,N_23488,N_23501);
or U24877 (N_24877,N_23629,N_23471);
nand U24878 (N_24878,N_23521,N_23525);
and U24879 (N_24879,N_23727,N_23596);
and U24880 (N_24880,N_23043,N_23860);
nand U24881 (N_24881,N_23856,N_23383);
or U24882 (N_24882,N_23883,N_23519);
nand U24883 (N_24883,N_23701,N_23767);
nand U24884 (N_24884,N_23639,N_23755);
and U24885 (N_24885,N_23242,N_23704);
or U24886 (N_24886,N_23050,N_23897);
or U24887 (N_24887,N_23430,N_23906);
xor U24888 (N_24888,N_23961,N_23618);
or U24889 (N_24889,N_23592,N_23060);
xnor U24890 (N_24890,N_23877,N_23121);
or U24891 (N_24891,N_23520,N_23482);
or U24892 (N_24892,N_23669,N_23753);
nor U24893 (N_24893,N_23983,N_23789);
nand U24894 (N_24894,N_23487,N_23187);
and U24895 (N_24895,N_23943,N_23466);
or U24896 (N_24896,N_23163,N_23016);
and U24897 (N_24897,N_23409,N_23609);
nand U24898 (N_24898,N_23565,N_23489);
nor U24899 (N_24899,N_23234,N_23277);
and U24900 (N_24900,N_23408,N_23101);
nand U24901 (N_24901,N_23584,N_23770);
or U24902 (N_24902,N_23362,N_23477);
nand U24903 (N_24903,N_23855,N_23107);
and U24904 (N_24904,N_23377,N_23588);
nand U24905 (N_24905,N_23199,N_23721);
or U24906 (N_24906,N_23105,N_23776);
nor U24907 (N_24907,N_23016,N_23816);
nand U24908 (N_24908,N_23018,N_23618);
and U24909 (N_24909,N_23773,N_23068);
nand U24910 (N_24910,N_23303,N_23672);
or U24911 (N_24911,N_23555,N_23128);
nand U24912 (N_24912,N_23025,N_23247);
or U24913 (N_24913,N_23799,N_23314);
xor U24914 (N_24914,N_23347,N_23561);
and U24915 (N_24915,N_23171,N_23532);
and U24916 (N_24916,N_23119,N_23886);
nand U24917 (N_24917,N_23812,N_23777);
and U24918 (N_24918,N_23926,N_23517);
and U24919 (N_24919,N_23835,N_23880);
and U24920 (N_24920,N_23931,N_23331);
nor U24921 (N_24921,N_23484,N_23222);
nor U24922 (N_24922,N_23761,N_23280);
xor U24923 (N_24923,N_23837,N_23154);
and U24924 (N_24924,N_23355,N_23016);
xnor U24925 (N_24925,N_23465,N_23365);
xor U24926 (N_24926,N_23497,N_23707);
and U24927 (N_24927,N_23525,N_23849);
and U24928 (N_24928,N_23820,N_23694);
or U24929 (N_24929,N_23396,N_23390);
and U24930 (N_24930,N_23437,N_23955);
or U24931 (N_24931,N_23598,N_23112);
and U24932 (N_24932,N_23300,N_23229);
nand U24933 (N_24933,N_23879,N_23754);
nor U24934 (N_24934,N_23742,N_23848);
and U24935 (N_24935,N_23597,N_23265);
or U24936 (N_24936,N_23556,N_23118);
or U24937 (N_24937,N_23047,N_23845);
and U24938 (N_24938,N_23579,N_23957);
xnor U24939 (N_24939,N_23292,N_23067);
xnor U24940 (N_24940,N_23734,N_23450);
xnor U24941 (N_24941,N_23455,N_23661);
nor U24942 (N_24942,N_23204,N_23718);
xor U24943 (N_24943,N_23205,N_23860);
and U24944 (N_24944,N_23255,N_23772);
nor U24945 (N_24945,N_23307,N_23819);
and U24946 (N_24946,N_23740,N_23749);
nor U24947 (N_24947,N_23112,N_23220);
or U24948 (N_24948,N_23163,N_23492);
and U24949 (N_24949,N_23877,N_23313);
nor U24950 (N_24950,N_23671,N_23494);
or U24951 (N_24951,N_23008,N_23001);
xnor U24952 (N_24952,N_23576,N_23668);
and U24953 (N_24953,N_23608,N_23579);
nor U24954 (N_24954,N_23220,N_23446);
and U24955 (N_24955,N_23652,N_23758);
xor U24956 (N_24956,N_23939,N_23932);
and U24957 (N_24957,N_23611,N_23515);
nand U24958 (N_24958,N_23107,N_23678);
nand U24959 (N_24959,N_23990,N_23305);
nor U24960 (N_24960,N_23844,N_23778);
and U24961 (N_24961,N_23184,N_23136);
nor U24962 (N_24962,N_23239,N_23269);
nor U24963 (N_24963,N_23621,N_23576);
nor U24964 (N_24964,N_23246,N_23580);
nand U24965 (N_24965,N_23570,N_23477);
nand U24966 (N_24966,N_23037,N_23390);
nor U24967 (N_24967,N_23587,N_23657);
xnor U24968 (N_24968,N_23866,N_23288);
xor U24969 (N_24969,N_23656,N_23784);
or U24970 (N_24970,N_23988,N_23686);
or U24971 (N_24971,N_23466,N_23415);
nor U24972 (N_24972,N_23963,N_23660);
or U24973 (N_24973,N_23773,N_23861);
or U24974 (N_24974,N_23363,N_23968);
and U24975 (N_24975,N_23966,N_23414);
nand U24976 (N_24976,N_23978,N_23762);
or U24977 (N_24977,N_23259,N_23734);
or U24978 (N_24978,N_23501,N_23785);
or U24979 (N_24979,N_23098,N_23459);
xnor U24980 (N_24980,N_23912,N_23974);
nor U24981 (N_24981,N_23764,N_23366);
nand U24982 (N_24982,N_23106,N_23273);
nand U24983 (N_24983,N_23044,N_23587);
nand U24984 (N_24984,N_23019,N_23838);
nor U24985 (N_24985,N_23074,N_23480);
or U24986 (N_24986,N_23426,N_23240);
or U24987 (N_24987,N_23143,N_23571);
xor U24988 (N_24988,N_23341,N_23941);
nor U24989 (N_24989,N_23030,N_23670);
nor U24990 (N_24990,N_23162,N_23043);
nor U24991 (N_24991,N_23267,N_23439);
and U24992 (N_24992,N_23509,N_23216);
xnor U24993 (N_24993,N_23430,N_23696);
nand U24994 (N_24994,N_23488,N_23054);
nor U24995 (N_24995,N_23882,N_23227);
nand U24996 (N_24996,N_23365,N_23110);
xor U24997 (N_24997,N_23075,N_23308);
nand U24998 (N_24998,N_23416,N_23064);
xor U24999 (N_24999,N_23885,N_23306);
xnor UO_0 (O_0,N_24160,N_24025);
nor UO_1 (O_1,N_24432,N_24594);
xor UO_2 (O_2,N_24762,N_24219);
xor UO_3 (O_3,N_24171,N_24189);
nor UO_4 (O_4,N_24424,N_24497);
or UO_5 (O_5,N_24835,N_24356);
xnor UO_6 (O_6,N_24578,N_24047);
and UO_7 (O_7,N_24111,N_24276);
xnor UO_8 (O_8,N_24183,N_24469);
nor UO_9 (O_9,N_24508,N_24096);
nand UO_10 (O_10,N_24650,N_24030);
and UO_11 (O_11,N_24077,N_24263);
and UO_12 (O_12,N_24336,N_24655);
xnor UO_13 (O_13,N_24476,N_24954);
or UO_14 (O_14,N_24233,N_24141);
xnor UO_15 (O_15,N_24317,N_24454);
nor UO_16 (O_16,N_24584,N_24274);
nand UO_17 (O_17,N_24975,N_24653);
xnor UO_18 (O_18,N_24491,N_24394);
xnor UO_19 (O_19,N_24235,N_24044);
nand UO_20 (O_20,N_24884,N_24215);
nor UO_21 (O_21,N_24677,N_24011);
nor UO_22 (O_22,N_24679,N_24240);
nor UO_23 (O_23,N_24278,N_24797);
nand UO_24 (O_24,N_24376,N_24669);
nor UO_25 (O_25,N_24720,N_24614);
xnor UO_26 (O_26,N_24507,N_24831);
xor UO_27 (O_27,N_24362,N_24123);
nand UO_28 (O_28,N_24637,N_24404);
nand UO_29 (O_29,N_24664,N_24602);
or UO_30 (O_30,N_24072,N_24449);
or UO_31 (O_31,N_24087,N_24898);
nand UO_32 (O_32,N_24868,N_24562);
xnor UO_33 (O_33,N_24100,N_24828);
nor UO_34 (O_34,N_24147,N_24808);
and UO_35 (O_35,N_24528,N_24838);
nor UO_36 (O_36,N_24731,N_24176);
and UO_37 (O_37,N_24146,N_24866);
nand UO_38 (O_38,N_24569,N_24040);
nand UO_39 (O_39,N_24220,N_24857);
nand UO_40 (O_40,N_24284,N_24861);
nand UO_41 (O_41,N_24204,N_24987);
nand UO_42 (O_42,N_24525,N_24092);
or UO_43 (O_43,N_24000,N_24870);
xnor UO_44 (O_44,N_24696,N_24994);
or UO_45 (O_45,N_24611,N_24557);
nand UO_46 (O_46,N_24254,N_24805);
or UO_47 (O_47,N_24417,N_24211);
and UO_48 (O_48,N_24206,N_24523);
or UO_49 (O_49,N_24467,N_24144);
xnor UO_50 (O_50,N_24398,N_24676);
xor UO_51 (O_51,N_24588,N_24707);
nand UO_52 (O_52,N_24896,N_24161);
nand UO_53 (O_53,N_24648,N_24208);
nor UO_54 (O_54,N_24132,N_24667);
xnor UO_55 (O_55,N_24344,N_24200);
and UO_56 (O_56,N_24524,N_24290);
or UO_57 (O_57,N_24463,N_24458);
and UO_58 (O_58,N_24652,N_24783);
and UO_59 (O_59,N_24081,N_24957);
or UO_60 (O_60,N_24370,N_24542);
and UO_61 (O_61,N_24430,N_24076);
nand UO_62 (O_62,N_24479,N_24829);
nor UO_63 (O_63,N_24156,N_24409);
or UO_64 (O_64,N_24801,N_24715);
xnor UO_65 (O_65,N_24251,N_24443);
nor UO_66 (O_66,N_24164,N_24891);
xor UO_67 (O_67,N_24711,N_24505);
and UO_68 (O_68,N_24833,N_24811);
and UO_69 (O_69,N_24924,N_24547);
nor UO_70 (O_70,N_24486,N_24559);
xnor UO_71 (O_71,N_24597,N_24026);
xnor UO_72 (O_72,N_24418,N_24522);
nand UO_73 (O_73,N_24060,N_24333);
and UO_74 (O_74,N_24166,N_24107);
nand UO_75 (O_75,N_24089,N_24633);
nand UO_76 (O_76,N_24198,N_24751);
or UO_77 (O_77,N_24538,N_24612);
and UO_78 (O_78,N_24120,N_24540);
xnor UO_79 (O_79,N_24130,N_24860);
nand UO_80 (O_80,N_24464,N_24150);
nor UO_81 (O_81,N_24721,N_24606);
nor UO_82 (O_82,N_24798,N_24493);
and UO_83 (O_83,N_24482,N_24440);
nand UO_84 (O_84,N_24425,N_24776);
and UO_85 (O_85,N_24143,N_24043);
nor UO_86 (O_86,N_24188,N_24148);
and UO_87 (O_87,N_24314,N_24999);
or UO_88 (O_88,N_24134,N_24061);
or UO_89 (O_89,N_24307,N_24590);
nand UO_90 (O_90,N_24136,N_24907);
and UO_91 (O_91,N_24444,N_24615);
xnor UO_92 (O_92,N_24018,N_24295);
xnor UO_93 (O_93,N_24347,N_24197);
xnor UO_94 (O_94,N_24520,N_24638);
or UO_95 (O_95,N_24790,N_24227);
and UO_96 (O_96,N_24007,N_24078);
and UO_97 (O_97,N_24623,N_24970);
nand UO_98 (O_98,N_24519,N_24242);
nor UO_99 (O_99,N_24475,N_24576);
nor UO_100 (O_100,N_24747,N_24599);
or UO_101 (O_101,N_24665,N_24930);
or UO_102 (O_102,N_24313,N_24434);
nand UO_103 (O_103,N_24743,N_24330);
and UO_104 (O_104,N_24905,N_24315);
or UO_105 (O_105,N_24341,N_24929);
nand UO_106 (O_106,N_24323,N_24617);
nand UO_107 (O_107,N_24022,N_24695);
nand UO_108 (O_108,N_24155,N_24733);
nand UO_109 (O_109,N_24858,N_24014);
or UO_110 (O_110,N_24224,N_24827);
nand UO_111 (O_111,N_24897,N_24471);
and UO_112 (O_112,N_24735,N_24563);
or UO_113 (O_113,N_24958,N_24572);
or UO_114 (O_114,N_24543,N_24549);
xor UO_115 (O_115,N_24748,N_24772);
nand UO_116 (O_116,N_24277,N_24480);
nand UO_117 (O_117,N_24710,N_24327);
xnor UO_118 (O_118,N_24969,N_24191);
or UO_119 (O_119,N_24324,N_24862);
xor UO_120 (O_120,N_24103,N_24113);
nand UO_121 (O_121,N_24369,N_24951);
xnor UO_122 (O_122,N_24066,N_24008);
nand UO_123 (O_123,N_24792,N_24610);
or UO_124 (O_124,N_24158,N_24825);
nor UO_125 (O_125,N_24624,N_24561);
and UO_126 (O_126,N_24462,N_24109);
and UO_127 (O_127,N_24770,N_24996);
and UO_128 (O_128,N_24820,N_24573);
nand UO_129 (O_129,N_24049,N_24989);
nor UO_130 (O_130,N_24744,N_24775);
and UO_131 (O_131,N_24169,N_24498);
nor UO_132 (O_132,N_24429,N_24332);
or UO_133 (O_133,N_24074,N_24746);
nand UO_134 (O_134,N_24977,N_24680);
xor UO_135 (O_135,N_24338,N_24700);
nor UO_136 (O_136,N_24364,N_24387);
nand UO_137 (O_137,N_24869,N_24035);
xnor UO_138 (O_138,N_24237,N_24504);
xor UO_139 (O_139,N_24302,N_24319);
and UO_140 (O_140,N_24657,N_24340);
xor UO_141 (O_141,N_24998,N_24938);
nor UO_142 (O_142,N_24410,N_24816);
nor UO_143 (O_143,N_24806,N_24532);
xor UO_144 (O_144,N_24021,N_24085);
nand UO_145 (O_145,N_24565,N_24567);
and UO_146 (O_146,N_24289,N_24736);
nor UO_147 (O_147,N_24548,N_24872);
nand UO_148 (O_148,N_24162,N_24834);
nand UO_149 (O_149,N_24228,N_24768);
xor UO_150 (O_150,N_24239,N_24604);
xor UO_151 (O_151,N_24603,N_24084);
xnor UO_152 (O_152,N_24714,N_24687);
nor UO_153 (O_153,N_24069,N_24613);
nor UO_154 (O_154,N_24979,N_24017);
and UO_155 (O_155,N_24071,N_24737);
and UO_156 (O_156,N_24546,N_24598);
xnor UO_157 (O_157,N_24264,N_24029);
xor UO_158 (O_158,N_24659,N_24564);
xor UO_159 (O_159,N_24075,N_24972);
or UO_160 (O_160,N_24133,N_24620);
and UO_161 (O_161,N_24342,N_24439);
nand UO_162 (O_162,N_24566,N_24729);
nor UO_163 (O_163,N_24119,N_24037);
or UO_164 (O_164,N_24823,N_24019);
xor UO_165 (O_165,N_24756,N_24851);
nand UO_166 (O_166,N_24789,N_24309);
xnor UO_167 (O_167,N_24045,N_24042);
and UO_168 (O_168,N_24099,N_24261);
and UO_169 (O_169,N_24916,N_24438);
nor UO_170 (O_170,N_24182,N_24587);
nand UO_171 (O_171,N_24764,N_24329);
xnor UO_172 (O_172,N_24609,N_24755);
xnor UO_173 (O_173,N_24765,N_24153);
nor UO_174 (O_174,N_24163,N_24506);
or UO_175 (O_175,N_24780,N_24436);
nor UO_176 (O_176,N_24173,N_24388);
nor UO_177 (O_177,N_24052,N_24016);
or UO_178 (O_178,N_24408,N_24810);
xnor UO_179 (O_179,N_24948,N_24003);
or UO_180 (O_180,N_24852,N_24126);
xnor UO_181 (O_181,N_24205,N_24413);
xnor UO_182 (O_182,N_24510,N_24990);
and UO_183 (O_183,N_24168,N_24817);
nor UO_184 (O_184,N_24112,N_24670);
nand UO_185 (O_185,N_24488,N_24796);
or UO_186 (O_186,N_24651,N_24672);
or UO_187 (O_187,N_24225,N_24766);
or UO_188 (O_188,N_24331,N_24943);
nor UO_189 (O_189,N_24115,N_24353);
and UO_190 (O_190,N_24684,N_24967);
nand UO_191 (O_191,N_24175,N_24708);
nor UO_192 (O_192,N_24232,N_24064);
nand UO_193 (O_193,N_24051,N_24361);
nand UO_194 (O_194,N_24279,N_24947);
or UO_195 (O_195,N_24705,N_24785);
or UO_196 (O_196,N_24842,N_24526);
or UO_197 (O_197,N_24568,N_24988);
or UO_198 (O_198,N_24591,N_24793);
and UO_199 (O_199,N_24596,N_24763);
nand UO_200 (O_200,N_24268,N_24297);
xnor UO_201 (O_201,N_24854,N_24402);
xor UO_202 (O_202,N_24445,N_24478);
xor UO_203 (O_203,N_24640,N_24723);
or UO_204 (O_204,N_24586,N_24005);
or UO_205 (O_205,N_24675,N_24724);
or UO_206 (O_206,N_24180,N_24583);
nand UO_207 (O_207,N_24393,N_24236);
nor UO_208 (O_208,N_24804,N_24460);
and UO_209 (O_209,N_24028,N_24855);
nor UO_210 (O_210,N_24814,N_24374);
xnor UO_211 (O_211,N_24271,N_24216);
nor UO_212 (O_212,N_24683,N_24065);
and UO_213 (O_213,N_24642,N_24784);
xor UO_214 (O_214,N_24844,N_24091);
xor UO_215 (O_215,N_24346,N_24135);
or UO_216 (O_216,N_24259,N_24571);
xnor UO_217 (O_217,N_24618,N_24978);
xnor UO_218 (O_218,N_24560,N_24058);
nand UO_219 (O_219,N_24968,N_24285);
nor UO_220 (O_220,N_24272,N_24223);
nand UO_221 (O_221,N_24213,N_24848);
and UO_222 (O_222,N_24974,N_24971);
and UO_223 (O_223,N_24310,N_24252);
nand UO_224 (O_224,N_24366,N_24073);
nor UO_225 (O_225,N_24773,N_24453);
and UO_226 (O_226,N_24411,N_24145);
and UO_227 (O_227,N_24193,N_24114);
nor UO_228 (O_228,N_24982,N_24316);
and UO_229 (O_229,N_24928,N_24986);
xor UO_230 (O_230,N_24845,N_24400);
or UO_231 (O_231,N_24448,N_24673);
or UO_232 (O_232,N_24405,N_24836);
nor UO_233 (O_233,N_24949,N_24824);
nand UO_234 (O_234,N_24849,N_24688);
xnor UO_235 (O_235,N_24709,N_24671);
and UO_236 (O_236,N_24937,N_24122);
xnor UO_237 (O_237,N_24095,N_24094);
and UO_238 (O_238,N_24229,N_24426);
or UO_239 (O_239,N_24457,N_24984);
nand UO_240 (O_240,N_24830,N_24935);
xnor UO_241 (O_241,N_24416,N_24865);
nor UO_242 (O_242,N_24367,N_24450);
or UO_243 (O_243,N_24082,N_24345);
nand UO_244 (O_244,N_24382,N_24280);
or UO_245 (O_245,N_24786,N_24983);
and UO_246 (O_246,N_24513,N_24779);
or UO_247 (O_247,N_24527,N_24068);
or UO_248 (O_248,N_24257,N_24373);
nand UO_249 (O_249,N_24759,N_24435);
or UO_250 (O_250,N_24901,N_24555);
nand UO_251 (O_251,N_24847,N_24992);
nand UO_252 (O_252,N_24149,N_24819);
nand UO_253 (O_253,N_24887,N_24803);
xor UO_254 (O_254,N_24976,N_24377);
nor UO_255 (O_255,N_24015,N_24249);
xnor UO_256 (O_256,N_24492,N_24911);
nor UO_257 (O_257,N_24697,N_24012);
xor UO_258 (O_258,N_24900,N_24931);
or UO_259 (O_259,N_24774,N_24904);
nor UO_260 (O_260,N_24207,N_24010);
nor UO_261 (O_261,N_24230,N_24485);
nor UO_262 (O_262,N_24646,N_24875);
nor UO_263 (O_263,N_24881,N_24939);
or UO_264 (O_264,N_24080,N_24262);
xnor UO_265 (O_265,N_24922,N_24758);
nand UO_266 (O_266,N_24945,N_24856);
nand UO_267 (O_267,N_24266,N_24481);
nor UO_268 (O_268,N_24529,N_24500);
nor UO_269 (O_269,N_24964,N_24873);
xor UO_270 (O_270,N_24632,N_24248);
and UO_271 (O_271,N_24247,N_24956);
and UO_272 (O_272,N_24809,N_24628);
nand UO_273 (O_273,N_24477,N_24864);
or UO_274 (O_274,N_24291,N_24116);
xor UO_275 (O_275,N_24258,N_24306);
xnor UO_276 (O_276,N_24575,N_24407);
or UO_277 (O_277,N_24118,N_24159);
nand UO_278 (O_278,N_24494,N_24605);
and UO_279 (O_279,N_24360,N_24455);
xor UO_280 (O_280,N_24267,N_24020);
xnor UO_281 (O_281,N_24589,N_24032);
xnor UO_282 (O_282,N_24574,N_24517);
and UO_283 (O_283,N_24050,N_24055);
or UO_284 (O_284,N_24698,N_24694);
or UO_285 (O_285,N_24321,N_24304);
xnor UO_286 (O_286,N_24878,N_24788);
or UO_287 (O_287,N_24178,N_24348);
and UO_288 (O_288,N_24371,N_24666);
or UO_289 (O_289,N_24401,N_24151);
nand UO_290 (O_290,N_24013,N_24212);
nand UO_291 (O_291,N_24414,N_24433);
or UO_292 (O_292,N_24093,N_24877);
and UO_293 (O_293,N_24850,N_24663);
and UO_294 (O_294,N_24647,N_24961);
xnor UO_295 (O_295,N_24892,N_24837);
nand UO_296 (O_296,N_24919,N_24383);
nand UO_297 (O_297,N_24940,N_24921);
and UO_298 (O_298,N_24337,N_24446);
nor UO_299 (O_299,N_24728,N_24600);
and UO_300 (O_300,N_24318,N_24518);
or UO_301 (O_301,N_24357,N_24509);
xnor UO_302 (O_302,N_24658,N_24138);
nor UO_303 (O_303,N_24722,N_24214);
nand UO_304 (O_304,N_24305,N_24385);
xor UO_305 (O_305,N_24350,N_24131);
and UO_306 (O_306,N_24893,N_24375);
nor UO_307 (O_307,N_24771,N_24502);
or UO_308 (O_308,N_24853,N_24201);
xor UO_309 (O_309,N_24355,N_24955);
or UO_310 (O_310,N_24157,N_24795);
and UO_311 (O_311,N_24920,N_24128);
and UO_312 (O_312,N_24472,N_24706);
xor UO_313 (O_313,N_24098,N_24351);
nand UO_314 (O_314,N_24883,N_24942);
nor UO_315 (O_315,N_24534,N_24154);
or UO_316 (O_316,N_24807,N_24459);
nand UO_317 (O_317,N_24265,N_24322);
nand UO_318 (O_318,N_24752,N_24281);
nand UO_319 (O_319,N_24033,N_24750);
or UO_320 (O_320,N_24124,N_24950);
nor UO_321 (O_321,N_24447,N_24354);
or UO_322 (O_322,N_24885,N_24913);
xnor UO_323 (O_323,N_24769,N_24902);
or UO_324 (O_324,N_24428,N_24726);
and UO_325 (O_325,N_24358,N_24048);
nor UO_326 (O_326,N_24363,N_24412);
nor UO_327 (O_327,N_24129,N_24293);
nand UO_328 (O_328,N_24923,N_24953);
and UO_329 (O_329,N_24456,N_24420);
nand UO_330 (O_330,N_24577,N_24915);
or UO_331 (O_331,N_24719,N_24580);
nand UO_332 (O_332,N_24914,N_24741);
and UO_333 (O_333,N_24004,N_24874);
or UO_334 (O_334,N_24406,N_24470);
xor UO_335 (O_335,N_24973,N_24501);
nand UO_336 (O_336,N_24423,N_24691);
xnor UO_337 (O_337,N_24952,N_24503);
xnor UO_338 (O_338,N_24941,N_24841);
or UO_339 (O_339,N_24644,N_24760);
and UO_340 (O_340,N_24717,N_24621);
and UO_341 (O_341,N_24067,N_24303);
nand UO_342 (O_342,N_24300,N_24545);
and UO_343 (O_343,N_24859,N_24101);
or UO_344 (O_344,N_24791,N_24023);
and UO_345 (O_345,N_24876,N_24312);
and UO_346 (O_346,N_24582,N_24894);
or UO_347 (O_347,N_24718,N_24946);
and UO_348 (O_348,N_24185,N_24753);
and UO_349 (O_349,N_24702,N_24889);
and UO_350 (O_350,N_24685,N_24932);
or UO_351 (O_351,N_24392,N_24121);
nor UO_352 (O_352,N_24630,N_24140);
and UO_353 (O_353,N_24372,N_24541);
nor UO_354 (O_354,N_24343,N_24738);
or UO_355 (O_355,N_24815,N_24437);
nand UO_356 (O_356,N_24622,N_24761);
or UO_357 (O_357,N_24745,N_24104);
and UO_358 (O_358,N_24287,N_24083);
xor UO_359 (O_359,N_24311,N_24794);
or UO_360 (O_360,N_24662,N_24693);
and UO_361 (O_361,N_24593,N_24002);
and UO_362 (O_362,N_24034,N_24521);
nand UO_363 (O_363,N_24734,N_24253);
or UO_364 (O_364,N_24725,N_24511);
or UO_365 (O_365,N_24699,N_24553);
and UO_366 (O_366,N_24390,N_24867);
nand UO_367 (O_367,N_24704,N_24294);
and UO_368 (O_368,N_24403,N_24550);
xnor UO_369 (O_369,N_24056,N_24800);
or UO_370 (O_370,N_24256,N_24754);
xnor UO_371 (O_371,N_24627,N_24378);
xnor UO_372 (O_372,N_24452,N_24778);
nand UO_373 (O_373,N_24328,N_24419);
nand UO_374 (O_374,N_24202,N_24282);
or UO_375 (O_375,N_24209,N_24079);
or UO_376 (O_376,N_24442,N_24165);
or UO_377 (O_377,N_24490,N_24234);
nand UO_378 (O_378,N_24535,N_24682);
xor UO_379 (O_379,N_24906,N_24912);
nand UO_380 (O_380,N_24152,N_24554);
nor UO_381 (O_381,N_24740,N_24537);
nor UO_382 (O_382,N_24465,N_24641);
nand UO_383 (O_383,N_24441,N_24057);
nand UO_384 (O_384,N_24246,N_24395);
or UO_385 (O_385,N_24006,N_24993);
and UO_386 (O_386,N_24713,N_24585);
or UO_387 (O_387,N_24298,N_24245);
or UO_388 (O_388,N_24187,N_24626);
nor UO_389 (O_389,N_24551,N_24552);
nor UO_390 (O_390,N_24712,N_24960);
nand UO_391 (O_391,N_24690,N_24487);
and UO_392 (O_392,N_24097,N_24727);
nor UO_393 (O_393,N_24217,N_24062);
nor UO_394 (O_394,N_24832,N_24918);
and UO_395 (O_395,N_24879,N_24299);
nand UO_396 (O_396,N_24255,N_24701);
nor UO_397 (O_397,N_24739,N_24269);
and UO_398 (O_398,N_24515,N_24530);
nor UO_399 (O_399,N_24339,N_24359);
xnor UO_400 (O_400,N_24415,N_24558);
or UO_401 (O_401,N_24601,N_24787);
nor UO_402 (O_402,N_24241,N_24273);
xor UO_403 (O_403,N_24936,N_24927);
and UO_404 (O_404,N_24222,N_24451);
or UO_405 (O_405,N_24296,N_24461);
nand UO_406 (O_406,N_24196,N_24473);
or UO_407 (O_407,N_24668,N_24431);
nand UO_408 (O_408,N_24105,N_24818);
nand UO_409 (O_409,N_24981,N_24592);
or UO_410 (O_410,N_24926,N_24368);
or UO_411 (O_411,N_24194,N_24777);
nor UO_412 (O_412,N_24260,N_24656);
xor UO_413 (O_413,N_24167,N_24767);
nor UO_414 (O_414,N_24802,N_24396);
nor UO_415 (O_415,N_24039,N_24352);
or UO_416 (O_416,N_24674,N_24581);
or UO_417 (O_417,N_24041,N_24086);
nand UO_418 (O_418,N_24474,N_24326);
nand UO_419 (O_419,N_24839,N_24365);
nand UO_420 (O_420,N_24110,N_24962);
xor UO_421 (O_421,N_24749,N_24221);
or UO_422 (O_422,N_24716,N_24944);
nor UO_423 (O_423,N_24181,N_24489);
nor UO_424 (O_424,N_24880,N_24177);
or UO_425 (O_425,N_24031,N_24172);
or UO_426 (O_426,N_24635,N_24995);
nor UO_427 (O_427,N_24389,N_24334);
or UO_428 (O_428,N_24625,N_24125);
and UO_429 (O_429,N_24629,N_24822);
and UO_430 (O_430,N_24886,N_24619);
xor UO_431 (O_431,N_24533,N_24966);
or UO_432 (O_432,N_24639,N_24985);
nand UO_433 (O_433,N_24757,N_24512);
xnor UO_434 (O_434,N_24910,N_24001);
nand UO_435 (O_435,N_24495,N_24218);
and UO_436 (O_436,N_24899,N_24643);
and UO_437 (O_437,N_24391,N_24102);
xnor UO_438 (O_438,N_24963,N_24270);
nand UO_439 (O_439,N_24381,N_24649);
and UO_440 (O_440,N_24631,N_24732);
or UO_441 (O_441,N_24514,N_24275);
or UO_442 (O_442,N_24933,N_24195);
nand UO_443 (O_443,N_24636,N_24840);
or UO_444 (O_444,N_24654,N_24127);
nand UO_445 (O_445,N_24024,N_24616);
and UO_446 (O_446,N_24250,N_24380);
nand UO_447 (O_447,N_24179,N_24226);
nor UO_448 (O_448,N_24421,N_24009);
xnor UO_449 (O_449,N_24645,N_24579);
nor UO_450 (O_450,N_24903,N_24308);
nand UO_451 (O_451,N_24496,N_24634);
xor UO_452 (O_452,N_24106,N_24117);
or UO_453 (O_453,N_24386,N_24283);
xnor UO_454 (O_454,N_24399,N_24203);
nand UO_455 (O_455,N_24142,N_24925);
nor UO_456 (O_456,N_24484,N_24499);
and UO_457 (O_457,N_24781,N_24063);
xnor UO_458 (O_458,N_24539,N_24595);
or UO_459 (O_459,N_24826,N_24190);
nand UO_460 (O_460,N_24917,N_24384);
xor UO_461 (O_461,N_24909,N_24607);
nor UO_462 (O_462,N_24730,N_24556);
and UO_463 (O_463,N_24813,N_24070);
nand UO_464 (O_464,N_24544,N_24821);
nand UO_465 (O_465,N_24799,N_24054);
or UO_466 (O_466,N_24038,N_24689);
and UO_467 (O_467,N_24882,N_24139);
nor UO_468 (O_468,N_24516,N_24703);
or UO_469 (O_469,N_24335,N_24301);
xnor UO_470 (O_470,N_24934,N_24046);
and UO_471 (O_471,N_24320,N_24243);
nor UO_472 (O_472,N_24325,N_24843);
xor UO_473 (O_473,N_24036,N_24686);
nand UO_474 (O_474,N_24184,N_24186);
and UO_475 (O_475,N_24108,N_24090);
xor UO_476 (O_476,N_24483,N_24570);
nand UO_477 (O_477,N_24660,N_24863);
or UO_478 (O_478,N_24980,N_24397);
nand UO_479 (O_479,N_24661,N_24888);
and UO_480 (O_480,N_24174,N_24536);
or UO_481 (O_481,N_24292,N_24238);
or UO_482 (O_482,N_24210,N_24059);
or UO_483 (O_483,N_24890,N_24053);
nor UO_484 (O_484,N_24379,N_24681);
nand UO_485 (O_485,N_24027,N_24782);
and UO_486 (O_486,N_24199,N_24427);
xnor UO_487 (O_487,N_24349,N_24231);
and UO_488 (O_488,N_24192,N_24959);
xnor UO_489 (O_489,N_24895,N_24244);
and UO_490 (O_490,N_24871,N_24088);
or UO_491 (O_491,N_24846,N_24137);
nand UO_492 (O_492,N_24170,N_24997);
or UO_493 (O_493,N_24908,N_24812);
or UO_494 (O_494,N_24466,N_24288);
nor UO_495 (O_495,N_24965,N_24692);
nand UO_496 (O_496,N_24468,N_24422);
xor UO_497 (O_497,N_24742,N_24286);
xnor UO_498 (O_498,N_24991,N_24678);
or UO_499 (O_499,N_24531,N_24608);
xnor UO_500 (O_500,N_24092,N_24804);
or UO_501 (O_501,N_24626,N_24733);
and UO_502 (O_502,N_24510,N_24377);
nor UO_503 (O_503,N_24613,N_24308);
or UO_504 (O_504,N_24046,N_24915);
xnor UO_505 (O_505,N_24241,N_24699);
and UO_506 (O_506,N_24294,N_24124);
nand UO_507 (O_507,N_24522,N_24554);
and UO_508 (O_508,N_24796,N_24823);
nor UO_509 (O_509,N_24213,N_24430);
xor UO_510 (O_510,N_24456,N_24635);
or UO_511 (O_511,N_24136,N_24723);
or UO_512 (O_512,N_24235,N_24742);
or UO_513 (O_513,N_24523,N_24522);
xnor UO_514 (O_514,N_24569,N_24261);
xnor UO_515 (O_515,N_24113,N_24636);
nand UO_516 (O_516,N_24363,N_24875);
and UO_517 (O_517,N_24981,N_24165);
or UO_518 (O_518,N_24118,N_24200);
and UO_519 (O_519,N_24615,N_24652);
or UO_520 (O_520,N_24592,N_24656);
nor UO_521 (O_521,N_24787,N_24582);
or UO_522 (O_522,N_24429,N_24527);
nor UO_523 (O_523,N_24985,N_24345);
nor UO_524 (O_524,N_24715,N_24536);
nand UO_525 (O_525,N_24340,N_24237);
nor UO_526 (O_526,N_24784,N_24820);
and UO_527 (O_527,N_24043,N_24210);
nand UO_528 (O_528,N_24362,N_24053);
nand UO_529 (O_529,N_24502,N_24730);
and UO_530 (O_530,N_24798,N_24601);
xor UO_531 (O_531,N_24513,N_24061);
and UO_532 (O_532,N_24471,N_24148);
nand UO_533 (O_533,N_24099,N_24479);
and UO_534 (O_534,N_24132,N_24509);
and UO_535 (O_535,N_24154,N_24375);
xor UO_536 (O_536,N_24889,N_24503);
xnor UO_537 (O_537,N_24587,N_24459);
xnor UO_538 (O_538,N_24258,N_24151);
and UO_539 (O_539,N_24405,N_24991);
nor UO_540 (O_540,N_24921,N_24050);
or UO_541 (O_541,N_24670,N_24279);
nor UO_542 (O_542,N_24168,N_24064);
nor UO_543 (O_543,N_24421,N_24194);
and UO_544 (O_544,N_24068,N_24481);
nor UO_545 (O_545,N_24688,N_24600);
and UO_546 (O_546,N_24401,N_24127);
nor UO_547 (O_547,N_24176,N_24710);
nor UO_548 (O_548,N_24458,N_24069);
or UO_549 (O_549,N_24697,N_24451);
xnor UO_550 (O_550,N_24902,N_24444);
nand UO_551 (O_551,N_24291,N_24702);
or UO_552 (O_552,N_24459,N_24250);
xnor UO_553 (O_553,N_24835,N_24636);
or UO_554 (O_554,N_24402,N_24400);
and UO_555 (O_555,N_24198,N_24375);
and UO_556 (O_556,N_24366,N_24984);
and UO_557 (O_557,N_24760,N_24519);
nor UO_558 (O_558,N_24338,N_24616);
xnor UO_559 (O_559,N_24880,N_24164);
and UO_560 (O_560,N_24700,N_24001);
xnor UO_561 (O_561,N_24452,N_24811);
or UO_562 (O_562,N_24893,N_24972);
and UO_563 (O_563,N_24624,N_24762);
xor UO_564 (O_564,N_24588,N_24135);
nand UO_565 (O_565,N_24315,N_24389);
nand UO_566 (O_566,N_24308,N_24379);
nand UO_567 (O_567,N_24355,N_24574);
or UO_568 (O_568,N_24563,N_24162);
and UO_569 (O_569,N_24472,N_24059);
nor UO_570 (O_570,N_24144,N_24436);
nor UO_571 (O_571,N_24061,N_24295);
nor UO_572 (O_572,N_24420,N_24599);
and UO_573 (O_573,N_24461,N_24711);
xor UO_574 (O_574,N_24207,N_24622);
xor UO_575 (O_575,N_24072,N_24528);
xnor UO_576 (O_576,N_24339,N_24720);
nand UO_577 (O_577,N_24180,N_24278);
or UO_578 (O_578,N_24023,N_24256);
xnor UO_579 (O_579,N_24248,N_24650);
or UO_580 (O_580,N_24765,N_24554);
nor UO_581 (O_581,N_24633,N_24634);
nor UO_582 (O_582,N_24105,N_24621);
nor UO_583 (O_583,N_24424,N_24734);
nor UO_584 (O_584,N_24307,N_24339);
and UO_585 (O_585,N_24847,N_24506);
nor UO_586 (O_586,N_24274,N_24394);
nor UO_587 (O_587,N_24289,N_24739);
and UO_588 (O_588,N_24494,N_24871);
or UO_589 (O_589,N_24958,N_24100);
and UO_590 (O_590,N_24240,N_24551);
nor UO_591 (O_591,N_24323,N_24167);
xor UO_592 (O_592,N_24132,N_24540);
nand UO_593 (O_593,N_24164,N_24444);
xor UO_594 (O_594,N_24457,N_24391);
nor UO_595 (O_595,N_24179,N_24379);
or UO_596 (O_596,N_24271,N_24840);
xnor UO_597 (O_597,N_24548,N_24147);
xor UO_598 (O_598,N_24541,N_24299);
nand UO_599 (O_599,N_24646,N_24199);
nand UO_600 (O_600,N_24084,N_24698);
or UO_601 (O_601,N_24158,N_24482);
nand UO_602 (O_602,N_24590,N_24555);
and UO_603 (O_603,N_24282,N_24885);
and UO_604 (O_604,N_24498,N_24776);
nand UO_605 (O_605,N_24015,N_24534);
nand UO_606 (O_606,N_24603,N_24125);
or UO_607 (O_607,N_24331,N_24350);
nor UO_608 (O_608,N_24067,N_24010);
nor UO_609 (O_609,N_24231,N_24979);
or UO_610 (O_610,N_24541,N_24368);
or UO_611 (O_611,N_24477,N_24087);
nand UO_612 (O_612,N_24826,N_24617);
xor UO_613 (O_613,N_24933,N_24644);
xor UO_614 (O_614,N_24219,N_24721);
and UO_615 (O_615,N_24968,N_24233);
and UO_616 (O_616,N_24891,N_24642);
or UO_617 (O_617,N_24595,N_24426);
nand UO_618 (O_618,N_24978,N_24998);
nor UO_619 (O_619,N_24997,N_24179);
nor UO_620 (O_620,N_24937,N_24853);
nand UO_621 (O_621,N_24087,N_24824);
or UO_622 (O_622,N_24345,N_24149);
and UO_623 (O_623,N_24972,N_24001);
xor UO_624 (O_624,N_24453,N_24076);
nand UO_625 (O_625,N_24204,N_24290);
or UO_626 (O_626,N_24000,N_24717);
or UO_627 (O_627,N_24036,N_24476);
xor UO_628 (O_628,N_24939,N_24043);
nand UO_629 (O_629,N_24814,N_24575);
xor UO_630 (O_630,N_24268,N_24023);
or UO_631 (O_631,N_24506,N_24840);
or UO_632 (O_632,N_24810,N_24138);
or UO_633 (O_633,N_24007,N_24142);
and UO_634 (O_634,N_24617,N_24927);
or UO_635 (O_635,N_24279,N_24706);
and UO_636 (O_636,N_24163,N_24394);
and UO_637 (O_637,N_24701,N_24325);
nand UO_638 (O_638,N_24104,N_24557);
nor UO_639 (O_639,N_24961,N_24358);
xnor UO_640 (O_640,N_24029,N_24470);
nand UO_641 (O_641,N_24642,N_24617);
and UO_642 (O_642,N_24747,N_24409);
nand UO_643 (O_643,N_24975,N_24287);
xnor UO_644 (O_644,N_24869,N_24536);
or UO_645 (O_645,N_24561,N_24790);
and UO_646 (O_646,N_24241,N_24775);
nor UO_647 (O_647,N_24114,N_24282);
and UO_648 (O_648,N_24549,N_24177);
or UO_649 (O_649,N_24807,N_24245);
nand UO_650 (O_650,N_24283,N_24883);
xor UO_651 (O_651,N_24124,N_24303);
and UO_652 (O_652,N_24523,N_24131);
nand UO_653 (O_653,N_24741,N_24708);
nor UO_654 (O_654,N_24858,N_24264);
xnor UO_655 (O_655,N_24578,N_24643);
nand UO_656 (O_656,N_24994,N_24928);
nor UO_657 (O_657,N_24267,N_24543);
nor UO_658 (O_658,N_24994,N_24676);
nand UO_659 (O_659,N_24202,N_24875);
nor UO_660 (O_660,N_24673,N_24287);
nand UO_661 (O_661,N_24203,N_24660);
or UO_662 (O_662,N_24730,N_24346);
nor UO_663 (O_663,N_24312,N_24323);
nand UO_664 (O_664,N_24411,N_24029);
nand UO_665 (O_665,N_24928,N_24940);
nor UO_666 (O_666,N_24479,N_24003);
nand UO_667 (O_667,N_24237,N_24525);
nor UO_668 (O_668,N_24100,N_24110);
and UO_669 (O_669,N_24787,N_24345);
nand UO_670 (O_670,N_24923,N_24074);
nand UO_671 (O_671,N_24245,N_24134);
or UO_672 (O_672,N_24181,N_24484);
nor UO_673 (O_673,N_24421,N_24732);
or UO_674 (O_674,N_24950,N_24103);
or UO_675 (O_675,N_24397,N_24400);
xnor UO_676 (O_676,N_24206,N_24590);
xnor UO_677 (O_677,N_24004,N_24921);
or UO_678 (O_678,N_24423,N_24904);
xor UO_679 (O_679,N_24143,N_24489);
and UO_680 (O_680,N_24251,N_24989);
and UO_681 (O_681,N_24881,N_24173);
xnor UO_682 (O_682,N_24367,N_24162);
or UO_683 (O_683,N_24963,N_24161);
nand UO_684 (O_684,N_24207,N_24469);
nand UO_685 (O_685,N_24290,N_24515);
nor UO_686 (O_686,N_24207,N_24160);
and UO_687 (O_687,N_24875,N_24186);
nor UO_688 (O_688,N_24299,N_24747);
nand UO_689 (O_689,N_24502,N_24397);
or UO_690 (O_690,N_24708,N_24900);
nand UO_691 (O_691,N_24097,N_24141);
nor UO_692 (O_692,N_24496,N_24275);
nor UO_693 (O_693,N_24138,N_24228);
nand UO_694 (O_694,N_24803,N_24789);
nor UO_695 (O_695,N_24155,N_24358);
or UO_696 (O_696,N_24914,N_24556);
xnor UO_697 (O_697,N_24326,N_24588);
nand UO_698 (O_698,N_24950,N_24909);
or UO_699 (O_699,N_24256,N_24363);
nand UO_700 (O_700,N_24179,N_24716);
xor UO_701 (O_701,N_24658,N_24401);
or UO_702 (O_702,N_24714,N_24319);
nand UO_703 (O_703,N_24192,N_24889);
nand UO_704 (O_704,N_24186,N_24809);
or UO_705 (O_705,N_24069,N_24587);
xnor UO_706 (O_706,N_24998,N_24139);
or UO_707 (O_707,N_24533,N_24335);
nor UO_708 (O_708,N_24083,N_24371);
or UO_709 (O_709,N_24303,N_24883);
nand UO_710 (O_710,N_24842,N_24437);
nor UO_711 (O_711,N_24099,N_24550);
nor UO_712 (O_712,N_24695,N_24813);
or UO_713 (O_713,N_24779,N_24207);
nand UO_714 (O_714,N_24940,N_24833);
nor UO_715 (O_715,N_24573,N_24766);
xnor UO_716 (O_716,N_24812,N_24742);
nor UO_717 (O_717,N_24801,N_24988);
nand UO_718 (O_718,N_24153,N_24043);
and UO_719 (O_719,N_24219,N_24958);
nor UO_720 (O_720,N_24583,N_24968);
nand UO_721 (O_721,N_24322,N_24034);
nor UO_722 (O_722,N_24473,N_24390);
nor UO_723 (O_723,N_24007,N_24527);
and UO_724 (O_724,N_24004,N_24897);
xnor UO_725 (O_725,N_24871,N_24408);
or UO_726 (O_726,N_24692,N_24661);
nor UO_727 (O_727,N_24687,N_24999);
nor UO_728 (O_728,N_24215,N_24293);
nand UO_729 (O_729,N_24629,N_24777);
and UO_730 (O_730,N_24624,N_24018);
nor UO_731 (O_731,N_24681,N_24237);
nand UO_732 (O_732,N_24578,N_24375);
nand UO_733 (O_733,N_24659,N_24416);
nor UO_734 (O_734,N_24544,N_24313);
xor UO_735 (O_735,N_24151,N_24165);
and UO_736 (O_736,N_24245,N_24481);
or UO_737 (O_737,N_24974,N_24509);
xnor UO_738 (O_738,N_24196,N_24532);
or UO_739 (O_739,N_24016,N_24523);
or UO_740 (O_740,N_24550,N_24823);
nor UO_741 (O_741,N_24145,N_24122);
or UO_742 (O_742,N_24267,N_24753);
and UO_743 (O_743,N_24202,N_24616);
or UO_744 (O_744,N_24071,N_24250);
nand UO_745 (O_745,N_24649,N_24729);
and UO_746 (O_746,N_24888,N_24555);
nand UO_747 (O_747,N_24522,N_24074);
xnor UO_748 (O_748,N_24992,N_24361);
nor UO_749 (O_749,N_24097,N_24484);
nand UO_750 (O_750,N_24126,N_24499);
and UO_751 (O_751,N_24682,N_24868);
and UO_752 (O_752,N_24358,N_24460);
nor UO_753 (O_753,N_24388,N_24502);
and UO_754 (O_754,N_24735,N_24254);
or UO_755 (O_755,N_24213,N_24075);
nor UO_756 (O_756,N_24282,N_24247);
xnor UO_757 (O_757,N_24040,N_24321);
nand UO_758 (O_758,N_24384,N_24224);
or UO_759 (O_759,N_24372,N_24178);
xnor UO_760 (O_760,N_24062,N_24536);
and UO_761 (O_761,N_24448,N_24586);
nor UO_762 (O_762,N_24057,N_24547);
nor UO_763 (O_763,N_24546,N_24570);
and UO_764 (O_764,N_24970,N_24814);
or UO_765 (O_765,N_24788,N_24659);
nand UO_766 (O_766,N_24174,N_24461);
nand UO_767 (O_767,N_24300,N_24268);
xor UO_768 (O_768,N_24007,N_24316);
xnor UO_769 (O_769,N_24161,N_24456);
xor UO_770 (O_770,N_24790,N_24140);
nor UO_771 (O_771,N_24163,N_24724);
nor UO_772 (O_772,N_24121,N_24105);
nor UO_773 (O_773,N_24881,N_24383);
nor UO_774 (O_774,N_24608,N_24410);
nand UO_775 (O_775,N_24460,N_24058);
or UO_776 (O_776,N_24913,N_24508);
or UO_777 (O_777,N_24061,N_24287);
nor UO_778 (O_778,N_24818,N_24025);
xor UO_779 (O_779,N_24886,N_24585);
and UO_780 (O_780,N_24654,N_24785);
xnor UO_781 (O_781,N_24410,N_24558);
or UO_782 (O_782,N_24558,N_24389);
or UO_783 (O_783,N_24957,N_24311);
nand UO_784 (O_784,N_24725,N_24937);
and UO_785 (O_785,N_24320,N_24683);
nand UO_786 (O_786,N_24496,N_24250);
and UO_787 (O_787,N_24962,N_24662);
nand UO_788 (O_788,N_24574,N_24121);
or UO_789 (O_789,N_24648,N_24122);
nor UO_790 (O_790,N_24401,N_24778);
and UO_791 (O_791,N_24087,N_24520);
or UO_792 (O_792,N_24074,N_24680);
and UO_793 (O_793,N_24369,N_24483);
and UO_794 (O_794,N_24777,N_24229);
xor UO_795 (O_795,N_24213,N_24486);
or UO_796 (O_796,N_24979,N_24412);
xnor UO_797 (O_797,N_24267,N_24946);
nand UO_798 (O_798,N_24142,N_24668);
nor UO_799 (O_799,N_24428,N_24696);
xor UO_800 (O_800,N_24363,N_24247);
and UO_801 (O_801,N_24777,N_24848);
or UO_802 (O_802,N_24640,N_24336);
nand UO_803 (O_803,N_24434,N_24288);
xor UO_804 (O_804,N_24009,N_24483);
xnor UO_805 (O_805,N_24265,N_24531);
or UO_806 (O_806,N_24749,N_24178);
or UO_807 (O_807,N_24502,N_24061);
or UO_808 (O_808,N_24003,N_24285);
nor UO_809 (O_809,N_24029,N_24311);
xor UO_810 (O_810,N_24870,N_24912);
nor UO_811 (O_811,N_24607,N_24005);
xor UO_812 (O_812,N_24725,N_24463);
nor UO_813 (O_813,N_24506,N_24721);
nand UO_814 (O_814,N_24518,N_24616);
and UO_815 (O_815,N_24701,N_24211);
or UO_816 (O_816,N_24793,N_24114);
or UO_817 (O_817,N_24460,N_24783);
nand UO_818 (O_818,N_24580,N_24257);
and UO_819 (O_819,N_24813,N_24850);
nand UO_820 (O_820,N_24446,N_24712);
nor UO_821 (O_821,N_24204,N_24129);
nand UO_822 (O_822,N_24573,N_24154);
or UO_823 (O_823,N_24830,N_24416);
or UO_824 (O_824,N_24995,N_24376);
nor UO_825 (O_825,N_24323,N_24431);
nor UO_826 (O_826,N_24642,N_24414);
xor UO_827 (O_827,N_24769,N_24117);
nor UO_828 (O_828,N_24282,N_24273);
or UO_829 (O_829,N_24448,N_24390);
or UO_830 (O_830,N_24568,N_24199);
or UO_831 (O_831,N_24894,N_24764);
or UO_832 (O_832,N_24020,N_24906);
nor UO_833 (O_833,N_24547,N_24046);
and UO_834 (O_834,N_24196,N_24533);
xor UO_835 (O_835,N_24236,N_24302);
nand UO_836 (O_836,N_24986,N_24097);
or UO_837 (O_837,N_24758,N_24415);
nand UO_838 (O_838,N_24371,N_24949);
xnor UO_839 (O_839,N_24972,N_24865);
xnor UO_840 (O_840,N_24119,N_24090);
nor UO_841 (O_841,N_24647,N_24025);
and UO_842 (O_842,N_24764,N_24866);
or UO_843 (O_843,N_24546,N_24312);
or UO_844 (O_844,N_24304,N_24824);
nand UO_845 (O_845,N_24572,N_24795);
and UO_846 (O_846,N_24688,N_24446);
or UO_847 (O_847,N_24604,N_24078);
nor UO_848 (O_848,N_24291,N_24376);
or UO_849 (O_849,N_24013,N_24424);
nand UO_850 (O_850,N_24372,N_24890);
and UO_851 (O_851,N_24792,N_24363);
xnor UO_852 (O_852,N_24975,N_24091);
nand UO_853 (O_853,N_24389,N_24240);
nor UO_854 (O_854,N_24696,N_24905);
nor UO_855 (O_855,N_24083,N_24569);
or UO_856 (O_856,N_24878,N_24070);
and UO_857 (O_857,N_24459,N_24423);
nor UO_858 (O_858,N_24882,N_24612);
nand UO_859 (O_859,N_24813,N_24721);
nand UO_860 (O_860,N_24581,N_24282);
nor UO_861 (O_861,N_24505,N_24694);
nand UO_862 (O_862,N_24663,N_24705);
and UO_863 (O_863,N_24755,N_24359);
nand UO_864 (O_864,N_24750,N_24252);
nand UO_865 (O_865,N_24959,N_24898);
nand UO_866 (O_866,N_24583,N_24588);
nor UO_867 (O_867,N_24935,N_24387);
nand UO_868 (O_868,N_24057,N_24601);
and UO_869 (O_869,N_24038,N_24096);
nor UO_870 (O_870,N_24059,N_24915);
or UO_871 (O_871,N_24967,N_24364);
or UO_872 (O_872,N_24317,N_24826);
nor UO_873 (O_873,N_24873,N_24607);
nor UO_874 (O_874,N_24420,N_24879);
and UO_875 (O_875,N_24362,N_24413);
nor UO_876 (O_876,N_24431,N_24222);
nor UO_877 (O_877,N_24304,N_24772);
and UO_878 (O_878,N_24923,N_24900);
xor UO_879 (O_879,N_24614,N_24112);
or UO_880 (O_880,N_24906,N_24402);
nor UO_881 (O_881,N_24997,N_24834);
or UO_882 (O_882,N_24851,N_24314);
nor UO_883 (O_883,N_24230,N_24904);
or UO_884 (O_884,N_24727,N_24667);
xnor UO_885 (O_885,N_24091,N_24010);
or UO_886 (O_886,N_24817,N_24365);
and UO_887 (O_887,N_24156,N_24467);
nand UO_888 (O_888,N_24909,N_24541);
or UO_889 (O_889,N_24321,N_24630);
or UO_890 (O_890,N_24860,N_24561);
and UO_891 (O_891,N_24491,N_24217);
or UO_892 (O_892,N_24343,N_24438);
nand UO_893 (O_893,N_24131,N_24633);
or UO_894 (O_894,N_24432,N_24398);
or UO_895 (O_895,N_24339,N_24800);
nor UO_896 (O_896,N_24835,N_24447);
xor UO_897 (O_897,N_24139,N_24379);
and UO_898 (O_898,N_24518,N_24055);
or UO_899 (O_899,N_24997,N_24073);
and UO_900 (O_900,N_24657,N_24318);
xnor UO_901 (O_901,N_24963,N_24042);
nand UO_902 (O_902,N_24984,N_24970);
and UO_903 (O_903,N_24757,N_24615);
or UO_904 (O_904,N_24870,N_24479);
xnor UO_905 (O_905,N_24417,N_24146);
and UO_906 (O_906,N_24956,N_24187);
and UO_907 (O_907,N_24191,N_24501);
or UO_908 (O_908,N_24534,N_24786);
nand UO_909 (O_909,N_24213,N_24743);
nand UO_910 (O_910,N_24434,N_24059);
nor UO_911 (O_911,N_24746,N_24430);
xor UO_912 (O_912,N_24132,N_24771);
nand UO_913 (O_913,N_24670,N_24628);
nor UO_914 (O_914,N_24006,N_24086);
and UO_915 (O_915,N_24719,N_24539);
xnor UO_916 (O_916,N_24399,N_24904);
nor UO_917 (O_917,N_24109,N_24182);
xnor UO_918 (O_918,N_24495,N_24236);
nand UO_919 (O_919,N_24677,N_24445);
or UO_920 (O_920,N_24088,N_24634);
and UO_921 (O_921,N_24403,N_24624);
xor UO_922 (O_922,N_24402,N_24211);
or UO_923 (O_923,N_24936,N_24129);
nand UO_924 (O_924,N_24420,N_24940);
and UO_925 (O_925,N_24510,N_24715);
and UO_926 (O_926,N_24522,N_24596);
or UO_927 (O_927,N_24930,N_24545);
nand UO_928 (O_928,N_24745,N_24827);
or UO_929 (O_929,N_24009,N_24132);
nor UO_930 (O_930,N_24196,N_24444);
or UO_931 (O_931,N_24966,N_24173);
nand UO_932 (O_932,N_24196,N_24657);
nor UO_933 (O_933,N_24390,N_24346);
and UO_934 (O_934,N_24359,N_24550);
xor UO_935 (O_935,N_24161,N_24140);
nand UO_936 (O_936,N_24014,N_24132);
nand UO_937 (O_937,N_24527,N_24550);
and UO_938 (O_938,N_24667,N_24503);
nor UO_939 (O_939,N_24817,N_24513);
nand UO_940 (O_940,N_24763,N_24479);
nand UO_941 (O_941,N_24843,N_24665);
and UO_942 (O_942,N_24601,N_24084);
and UO_943 (O_943,N_24448,N_24925);
and UO_944 (O_944,N_24093,N_24776);
xor UO_945 (O_945,N_24690,N_24219);
xnor UO_946 (O_946,N_24491,N_24642);
or UO_947 (O_947,N_24810,N_24861);
nand UO_948 (O_948,N_24675,N_24131);
and UO_949 (O_949,N_24670,N_24249);
xor UO_950 (O_950,N_24151,N_24055);
nand UO_951 (O_951,N_24605,N_24236);
nor UO_952 (O_952,N_24585,N_24795);
xnor UO_953 (O_953,N_24912,N_24748);
or UO_954 (O_954,N_24313,N_24716);
nand UO_955 (O_955,N_24459,N_24179);
nand UO_956 (O_956,N_24167,N_24046);
nor UO_957 (O_957,N_24822,N_24593);
nand UO_958 (O_958,N_24361,N_24479);
nor UO_959 (O_959,N_24446,N_24295);
nor UO_960 (O_960,N_24649,N_24499);
and UO_961 (O_961,N_24658,N_24677);
nand UO_962 (O_962,N_24800,N_24061);
xnor UO_963 (O_963,N_24277,N_24702);
xnor UO_964 (O_964,N_24268,N_24184);
nand UO_965 (O_965,N_24659,N_24213);
and UO_966 (O_966,N_24137,N_24710);
and UO_967 (O_967,N_24077,N_24634);
xor UO_968 (O_968,N_24768,N_24648);
or UO_969 (O_969,N_24800,N_24205);
and UO_970 (O_970,N_24566,N_24973);
nand UO_971 (O_971,N_24834,N_24082);
xnor UO_972 (O_972,N_24683,N_24297);
or UO_973 (O_973,N_24678,N_24564);
xnor UO_974 (O_974,N_24568,N_24610);
nand UO_975 (O_975,N_24897,N_24479);
or UO_976 (O_976,N_24686,N_24291);
or UO_977 (O_977,N_24474,N_24850);
and UO_978 (O_978,N_24650,N_24203);
nand UO_979 (O_979,N_24095,N_24226);
or UO_980 (O_980,N_24854,N_24065);
or UO_981 (O_981,N_24449,N_24933);
and UO_982 (O_982,N_24086,N_24860);
xor UO_983 (O_983,N_24402,N_24837);
nand UO_984 (O_984,N_24551,N_24502);
and UO_985 (O_985,N_24451,N_24804);
xor UO_986 (O_986,N_24031,N_24772);
or UO_987 (O_987,N_24890,N_24369);
xor UO_988 (O_988,N_24368,N_24367);
xnor UO_989 (O_989,N_24166,N_24809);
nand UO_990 (O_990,N_24221,N_24378);
and UO_991 (O_991,N_24048,N_24273);
xor UO_992 (O_992,N_24055,N_24411);
and UO_993 (O_993,N_24578,N_24398);
nand UO_994 (O_994,N_24027,N_24223);
or UO_995 (O_995,N_24849,N_24162);
nand UO_996 (O_996,N_24432,N_24826);
and UO_997 (O_997,N_24162,N_24981);
or UO_998 (O_998,N_24506,N_24768);
or UO_999 (O_999,N_24044,N_24215);
or UO_1000 (O_1000,N_24174,N_24194);
nand UO_1001 (O_1001,N_24632,N_24359);
nand UO_1002 (O_1002,N_24699,N_24748);
and UO_1003 (O_1003,N_24730,N_24718);
nor UO_1004 (O_1004,N_24438,N_24845);
nor UO_1005 (O_1005,N_24314,N_24712);
nor UO_1006 (O_1006,N_24608,N_24877);
nor UO_1007 (O_1007,N_24167,N_24654);
or UO_1008 (O_1008,N_24598,N_24356);
nand UO_1009 (O_1009,N_24340,N_24772);
xor UO_1010 (O_1010,N_24362,N_24164);
and UO_1011 (O_1011,N_24227,N_24165);
and UO_1012 (O_1012,N_24758,N_24299);
xnor UO_1013 (O_1013,N_24731,N_24739);
xnor UO_1014 (O_1014,N_24060,N_24752);
xnor UO_1015 (O_1015,N_24014,N_24239);
nor UO_1016 (O_1016,N_24608,N_24406);
xnor UO_1017 (O_1017,N_24334,N_24642);
nand UO_1018 (O_1018,N_24817,N_24085);
or UO_1019 (O_1019,N_24043,N_24370);
nor UO_1020 (O_1020,N_24591,N_24563);
nor UO_1021 (O_1021,N_24309,N_24821);
nor UO_1022 (O_1022,N_24152,N_24068);
xnor UO_1023 (O_1023,N_24496,N_24283);
or UO_1024 (O_1024,N_24469,N_24532);
xor UO_1025 (O_1025,N_24336,N_24439);
xor UO_1026 (O_1026,N_24215,N_24147);
nor UO_1027 (O_1027,N_24664,N_24431);
xor UO_1028 (O_1028,N_24093,N_24667);
nor UO_1029 (O_1029,N_24408,N_24853);
nand UO_1030 (O_1030,N_24866,N_24055);
nor UO_1031 (O_1031,N_24944,N_24533);
or UO_1032 (O_1032,N_24079,N_24382);
and UO_1033 (O_1033,N_24525,N_24582);
nand UO_1034 (O_1034,N_24977,N_24813);
xnor UO_1035 (O_1035,N_24443,N_24369);
xor UO_1036 (O_1036,N_24741,N_24307);
and UO_1037 (O_1037,N_24847,N_24855);
or UO_1038 (O_1038,N_24041,N_24153);
nor UO_1039 (O_1039,N_24739,N_24569);
xor UO_1040 (O_1040,N_24387,N_24978);
or UO_1041 (O_1041,N_24197,N_24050);
nor UO_1042 (O_1042,N_24241,N_24455);
nand UO_1043 (O_1043,N_24338,N_24484);
and UO_1044 (O_1044,N_24437,N_24713);
nor UO_1045 (O_1045,N_24745,N_24533);
nor UO_1046 (O_1046,N_24192,N_24613);
and UO_1047 (O_1047,N_24322,N_24271);
nor UO_1048 (O_1048,N_24953,N_24251);
xnor UO_1049 (O_1049,N_24065,N_24702);
and UO_1050 (O_1050,N_24690,N_24525);
nand UO_1051 (O_1051,N_24867,N_24547);
nor UO_1052 (O_1052,N_24752,N_24206);
nor UO_1053 (O_1053,N_24997,N_24061);
nand UO_1054 (O_1054,N_24892,N_24776);
nand UO_1055 (O_1055,N_24723,N_24357);
nor UO_1056 (O_1056,N_24391,N_24756);
nor UO_1057 (O_1057,N_24067,N_24285);
nor UO_1058 (O_1058,N_24613,N_24874);
nand UO_1059 (O_1059,N_24043,N_24353);
nand UO_1060 (O_1060,N_24198,N_24961);
or UO_1061 (O_1061,N_24036,N_24594);
xor UO_1062 (O_1062,N_24847,N_24449);
nor UO_1063 (O_1063,N_24056,N_24657);
xnor UO_1064 (O_1064,N_24583,N_24485);
nor UO_1065 (O_1065,N_24109,N_24952);
xor UO_1066 (O_1066,N_24925,N_24516);
xnor UO_1067 (O_1067,N_24476,N_24086);
and UO_1068 (O_1068,N_24495,N_24526);
nor UO_1069 (O_1069,N_24246,N_24264);
and UO_1070 (O_1070,N_24925,N_24520);
nor UO_1071 (O_1071,N_24410,N_24381);
xnor UO_1072 (O_1072,N_24766,N_24996);
or UO_1073 (O_1073,N_24209,N_24842);
or UO_1074 (O_1074,N_24863,N_24594);
or UO_1075 (O_1075,N_24722,N_24847);
xor UO_1076 (O_1076,N_24311,N_24475);
nand UO_1077 (O_1077,N_24338,N_24762);
nor UO_1078 (O_1078,N_24397,N_24945);
xnor UO_1079 (O_1079,N_24680,N_24330);
nor UO_1080 (O_1080,N_24872,N_24004);
xor UO_1081 (O_1081,N_24291,N_24771);
and UO_1082 (O_1082,N_24968,N_24341);
xnor UO_1083 (O_1083,N_24533,N_24804);
nor UO_1084 (O_1084,N_24671,N_24977);
nand UO_1085 (O_1085,N_24283,N_24347);
and UO_1086 (O_1086,N_24978,N_24601);
and UO_1087 (O_1087,N_24253,N_24913);
nand UO_1088 (O_1088,N_24415,N_24306);
xor UO_1089 (O_1089,N_24273,N_24999);
nand UO_1090 (O_1090,N_24965,N_24608);
or UO_1091 (O_1091,N_24338,N_24467);
xnor UO_1092 (O_1092,N_24749,N_24996);
or UO_1093 (O_1093,N_24164,N_24781);
xnor UO_1094 (O_1094,N_24402,N_24020);
and UO_1095 (O_1095,N_24608,N_24861);
nor UO_1096 (O_1096,N_24631,N_24597);
and UO_1097 (O_1097,N_24176,N_24447);
or UO_1098 (O_1098,N_24459,N_24766);
xor UO_1099 (O_1099,N_24474,N_24023);
or UO_1100 (O_1100,N_24426,N_24621);
nor UO_1101 (O_1101,N_24630,N_24222);
or UO_1102 (O_1102,N_24658,N_24163);
or UO_1103 (O_1103,N_24831,N_24307);
nand UO_1104 (O_1104,N_24517,N_24737);
xor UO_1105 (O_1105,N_24872,N_24108);
nor UO_1106 (O_1106,N_24685,N_24235);
nor UO_1107 (O_1107,N_24024,N_24152);
or UO_1108 (O_1108,N_24467,N_24844);
and UO_1109 (O_1109,N_24097,N_24644);
nand UO_1110 (O_1110,N_24998,N_24683);
or UO_1111 (O_1111,N_24115,N_24398);
nand UO_1112 (O_1112,N_24472,N_24148);
xnor UO_1113 (O_1113,N_24561,N_24890);
nor UO_1114 (O_1114,N_24121,N_24094);
xnor UO_1115 (O_1115,N_24853,N_24682);
nor UO_1116 (O_1116,N_24384,N_24760);
nand UO_1117 (O_1117,N_24755,N_24464);
xnor UO_1118 (O_1118,N_24229,N_24215);
nand UO_1119 (O_1119,N_24653,N_24046);
nand UO_1120 (O_1120,N_24137,N_24325);
xor UO_1121 (O_1121,N_24546,N_24437);
and UO_1122 (O_1122,N_24557,N_24604);
nor UO_1123 (O_1123,N_24056,N_24341);
xnor UO_1124 (O_1124,N_24569,N_24337);
xnor UO_1125 (O_1125,N_24583,N_24234);
nand UO_1126 (O_1126,N_24676,N_24375);
and UO_1127 (O_1127,N_24343,N_24188);
and UO_1128 (O_1128,N_24041,N_24766);
nor UO_1129 (O_1129,N_24487,N_24717);
xor UO_1130 (O_1130,N_24023,N_24633);
or UO_1131 (O_1131,N_24039,N_24386);
nor UO_1132 (O_1132,N_24972,N_24316);
nand UO_1133 (O_1133,N_24317,N_24120);
and UO_1134 (O_1134,N_24743,N_24299);
xnor UO_1135 (O_1135,N_24212,N_24010);
nor UO_1136 (O_1136,N_24243,N_24238);
nand UO_1137 (O_1137,N_24456,N_24198);
nor UO_1138 (O_1138,N_24905,N_24431);
nor UO_1139 (O_1139,N_24739,N_24951);
or UO_1140 (O_1140,N_24614,N_24028);
and UO_1141 (O_1141,N_24903,N_24405);
xor UO_1142 (O_1142,N_24053,N_24691);
nand UO_1143 (O_1143,N_24934,N_24570);
and UO_1144 (O_1144,N_24489,N_24516);
or UO_1145 (O_1145,N_24197,N_24070);
or UO_1146 (O_1146,N_24617,N_24498);
xor UO_1147 (O_1147,N_24245,N_24882);
or UO_1148 (O_1148,N_24560,N_24595);
nor UO_1149 (O_1149,N_24311,N_24574);
nor UO_1150 (O_1150,N_24154,N_24122);
xor UO_1151 (O_1151,N_24049,N_24876);
and UO_1152 (O_1152,N_24922,N_24387);
or UO_1153 (O_1153,N_24176,N_24668);
and UO_1154 (O_1154,N_24039,N_24802);
or UO_1155 (O_1155,N_24943,N_24713);
xnor UO_1156 (O_1156,N_24694,N_24803);
nor UO_1157 (O_1157,N_24000,N_24705);
nand UO_1158 (O_1158,N_24147,N_24720);
xnor UO_1159 (O_1159,N_24387,N_24781);
nor UO_1160 (O_1160,N_24964,N_24645);
nor UO_1161 (O_1161,N_24521,N_24849);
xnor UO_1162 (O_1162,N_24439,N_24632);
nand UO_1163 (O_1163,N_24100,N_24637);
nor UO_1164 (O_1164,N_24344,N_24654);
and UO_1165 (O_1165,N_24492,N_24740);
xnor UO_1166 (O_1166,N_24107,N_24401);
and UO_1167 (O_1167,N_24857,N_24363);
xor UO_1168 (O_1168,N_24103,N_24828);
xor UO_1169 (O_1169,N_24728,N_24547);
nand UO_1170 (O_1170,N_24265,N_24586);
nand UO_1171 (O_1171,N_24745,N_24281);
xnor UO_1172 (O_1172,N_24483,N_24937);
and UO_1173 (O_1173,N_24885,N_24950);
or UO_1174 (O_1174,N_24855,N_24625);
or UO_1175 (O_1175,N_24418,N_24708);
xnor UO_1176 (O_1176,N_24925,N_24808);
or UO_1177 (O_1177,N_24983,N_24930);
nor UO_1178 (O_1178,N_24610,N_24425);
nand UO_1179 (O_1179,N_24518,N_24724);
or UO_1180 (O_1180,N_24317,N_24426);
and UO_1181 (O_1181,N_24667,N_24150);
xnor UO_1182 (O_1182,N_24215,N_24927);
nand UO_1183 (O_1183,N_24465,N_24699);
and UO_1184 (O_1184,N_24319,N_24999);
and UO_1185 (O_1185,N_24544,N_24778);
nor UO_1186 (O_1186,N_24624,N_24545);
nor UO_1187 (O_1187,N_24061,N_24198);
xnor UO_1188 (O_1188,N_24280,N_24059);
or UO_1189 (O_1189,N_24957,N_24568);
or UO_1190 (O_1190,N_24910,N_24847);
or UO_1191 (O_1191,N_24145,N_24975);
xnor UO_1192 (O_1192,N_24349,N_24466);
xor UO_1193 (O_1193,N_24022,N_24974);
or UO_1194 (O_1194,N_24314,N_24213);
xnor UO_1195 (O_1195,N_24846,N_24351);
xor UO_1196 (O_1196,N_24512,N_24264);
and UO_1197 (O_1197,N_24638,N_24474);
or UO_1198 (O_1198,N_24187,N_24372);
or UO_1199 (O_1199,N_24860,N_24617);
nor UO_1200 (O_1200,N_24964,N_24431);
nand UO_1201 (O_1201,N_24405,N_24819);
or UO_1202 (O_1202,N_24393,N_24720);
and UO_1203 (O_1203,N_24907,N_24651);
and UO_1204 (O_1204,N_24073,N_24454);
nor UO_1205 (O_1205,N_24394,N_24732);
and UO_1206 (O_1206,N_24411,N_24313);
and UO_1207 (O_1207,N_24357,N_24936);
and UO_1208 (O_1208,N_24012,N_24207);
nor UO_1209 (O_1209,N_24632,N_24426);
xnor UO_1210 (O_1210,N_24500,N_24513);
xor UO_1211 (O_1211,N_24281,N_24357);
and UO_1212 (O_1212,N_24958,N_24130);
or UO_1213 (O_1213,N_24266,N_24910);
or UO_1214 (O_1214,N_24505,N_24246);
or UO_1215 (O_1215,N_24766,N_24084);
and UO_1216 (O_1216,N_24050,N_24394);
or UO_1217 (O_1217,N_24928,N_24373);
nor UO_1218 (O_1218,N_24781,N_24370);
nand UO_1219 (O_1219,N_24239,N_24162);
and UO_1220 (O_1220,N_24705,N_24807);
and UO_1221 (O_1221,N_24719,N_24476);
and UO_1222 (O_1222,N_24344,N_24509);
nand UO_1223 (O_1223,N_24022,N_24485);
or UO_1224 (O_1224,N_24406,N_24089);
nor UO_1225 (O_1225,N_24215,N_24352);
nand UO_1226 (O_1226,N_24943,N_24152);
nor UO_1227 (O_1227,N_24375,N_24704);
nand UO_1228 (O_1228,N_24810,N_24668);
nand UO_1229 (O_1229,N_24593,N_24971);
or UO_1230 (O_1230,N_24213,N_24463);
nand UO_1231 (O_1231,N_24111,N_24154);
nor UO_1232 (O_1232,N_24349,N_24859);
xnor UO_1233 (O_1233,N_24358,N_24493);
nand UO_1234 (O_1234,N_24487,N_24939);
or UO_1235 (O_1235,N_24690,N_24097);
and UO_1236 (O_1236,N_24079,N_24733);
and UO_1237 (O_1237,N_24071,N_24878);
xnor UO_1238 (O_1238,N_24883,N_24265);
or UO_1239 (O_1239,N_24283,N_24448);
nand UO_1240 (O_1240,N_24137,N_24196);
nand UO_1241 (O_1241,N_24416,N_24198);
nand UO_1242 (O_1242,N_24631,N_24912);
nand UO_1243 (O_1243,N_24372,N_24962);
nor UO_1244 (O_1244,N_24567,N_24649);
nor UO_1245 (O_1245,N_24835,N_24696);
nand UO_1246 (O_1246,N_24054,N_24017);
or UO_1247 (O_1247,N_24009,N_24989);
or UO_1248 (O_1248,N_24890,N_24671);
or UO_1249 (O_1249,N_24952,N_24679);
and UO_1250 (O_1250,N_24999,N_24341);
nand UO_1251 (O_1251,N_24493,N_24166);
xor UO_1252 (O_1252,N_24549,N_24547);
xnor UO_1253 (O_1253,N_24317,N_24570);
and UO_1254 (O_1254,N_24174,N_24381);
nand UO_1255 (O_1255,N_24788,N_24276);
and UO_1256 (O_1256,N_24087,N_24670);
nor UO_1257 (O_1257,N_24744,N_24373);
nor UO_1258 (O_1258,N_24118,N_24999);
nand UO_1259 (O_1259,N_24960,N_24420);
or UO_1260 (O_1260,N_24537,N_24997);
or UO_1261 (O_1261,N_24223,N_24584);
or UO_1262 (O_1262,N_24586,N_24875);
or UO_1263 (O_1263,N_24522,N_24770);
nand UO_1264 (O_1264,N_24128,N_24020);
or UO_1265 (O_1265,N_24983,N_24615);
or UO_1266 (O_1266,N_24351,N_24211);
nand UO_1267 (O_1267,N_24612,N_24628);
nor UO_1268 (O_1268,N_24456,N_24523);
or UO_1269 (O_1269,N_24314,N_24956);
nand UO_1270 (O_1270,N_24091,N_24725);
xor UO_1271 (O_1271,N_24055,N_24512);
nand UO_1272 (O_1272,N_24765,N_24928);
nand UO_1273 (O_1273,N_24410,N_24096);
xor UO_1274 (O_1274,N_24060,N_24365);
xor UO_1275 (O_1275,N_24734,N_24942);
xnor UO_1276 (O_1276,N_24484,N_24730);
nand UO_1277 (O_1277,N_24263,N_24649);
or UO_1278 (O_1278,N_24444,N_24097);
nand UO_1279 (O_1279,N_24800,N_24228);
and UO_1280 (O_1280,N_24126,N_24982);
nand UO_1281 (O_1281,N_24317,N_24632);
nand UO_1282 (O_1282,N_24498,N_24077);
nand UO_1283 (O_1283,N_24267,N_24135);
or UO_1284 (O_1284,N_24144,N_24819);
xor UO_1285 (O_1285,N_24800,N_24201);
and UO_1286 (O_1286,N_24412,N_24066);
or UO_1287 (O_1287,N_24507,N_24876);
or UO_1288 (O_1288,N_24013,N_24022);
nor UO_1289 (O_1289,N_24513,N_24316);
xor UO_1290 (O_1290,N_24294,N_24720);
xnor UO_1291 (O_1291,N_24727,N_24067);
nand UO_1292 (O_1292,N_24057,N_24283);
and UO_1293 (O_1293,N_24127,N_24898);
nor UO_1294 (O_1294,N_24349,N_24599);
and UO_1295 (O_1295,N_24581,N_24661);
or UO_1296 (O_1296,N_24635,N_24188);
and UO_1297 (O_1297,N_24534,N_24807);
xor UO_1298 (O_1298,N_24738,N_24206);
nand UO_1299 (O_1299,N_24999,N_24107);
nor UO_1300 (O_1300,N_24451,N_24919);
nand UO_1301 (O_1301,N_24553,N_24083);
xor UO_1302 (O_1302,N_24173,N_24509);
nand UO_1303 (O_1303,N_24224,N_24200);
nand UO_1304 (O_1304,N_24664,N_24756);
and UO_1305 (O_1305,N_24199,N_24783);
or UO_1306 (O_1306,N_24397,N_24622);
nand UO_1307 (O_1307,N_24511,N_24662);
or UO_1308 (O_1308,N_24694,N_24262);
or UO_1309 (O_1309,N_24003,N_24107);
and UO_1310 (O_1310,N_24065,N_24444);
nor UO_1311 (O_1311,N_24448,N_24442);
nand UO_1312 (O_1312,N_24901,N_24805);
nand UO_1313 (O_1313,N_24305,N_24912);
xnor UO_1314 (O_1314,N_24283,N_24425);
or UO_1315 (O_1315,N_24381,N_24618);
nand UO_1316 (O_1316,N_24107,N_24020);
or UO_1317 (O_1317,N_24259,N_24168);
or UO_1318 (O_1318,N_24621,N_24454);
nand UO_1319 (O_1319,N_24673,N_24986);
and UO_1320 (O_1320,N_24553,N_24414);
and UO_1321 (O_1321,N_24462,N_24027);
or UO_1322 (O_1322,N_24151,N_24913);
nand UO_1323 (O_1323,N_24723,N_24867);
or UO_1324 (O_1324,N_24922,N_24579);
or UO_1325 (O_1325,N_24927,N_24561);
or UO_1326 (O_1326,N_24618,N_24338);
and UO_1327 (O_1327,N_24679,N_24444);
nand UO_1328 (O_1328,N_24461,N_24227);
or UO_1329 (O_1329,N_24230,N_24050);
nor UO_1330 (O_1330,N_24304,N_24509);
xnor UO_1331 (O_1331,N_24223,N_24621);
xor UO_1332 (O_1332,N_24249,N_24734);
or UO_1333 (O_1333,N_24545,N_24220);
xnor UO_1334 (O_1334,N_24758,N_24523);
or UO_1335 (O_1335,N_24442,N_24724);
nor UO_1336 (O_1336,N_24011,N_24075);
nor UO_1337 (O_1337,N_24162,N_24487);
or UO_1338 (O_1338,N_24038,N_24353);
and UO_1339 (O_1339,N_24329,N_24111);
or UO_1340 (O_1340,N_24357,N_24969);
or UO_1341 (O_1341,N_24709,N_24183);
nand UO_1342 (O_1342,N_24964,N_24534);
nand UO_1343 (O_1343,N_24367,N_24906);
or UO_1344 (O_1344,N_24550,N_24224);
xnor UO_1345 (O_1345,N_24514,N_24507);
nand UO_1346 (O_1346,N_24927,N_24465);
nand UO_1347 (O_1347,N_24015,N_24679);
nand UO_1348 (O_1348,N_24217,N_24747);
or UO_1349 (O_1349,N_24100,N_24304);
or UO_1350 (O_1350,N_24517,N_24116);
and UO_1351 (O_1351,N_24423,N_24506);
xor UO_1352 (O_1352,N_24589,N_24605);
xor UO_1353 (O_1353,N_24103,N_24281);
nand UO_1354 (O_1354,N_24867,N_24034);
nor UO_1355 (O_1355,N_24853,N_24747);
xnor UO_1356 (O_1356,N_24610,N_24977);
nor UO_1357 (O_1357,N_24212,N_24811);
nor UO_1358 (O_1358,N_24310,N_24160);
xor UO_1359 (O_1359,N_24228,N_24090);
xnor UO_1360 (O_1360,N_24325,N_24602);
and UO_1361 (O_1361,N_24707,N_24424);
and UO_1362 (O_1362,N_24841,N_24339);
nand UO_1363 (O_1363,N_24081,N_24996);
nand UO_1364 (O_1364,N_24380,N_24042);
nand UO_1365 (O_1365,N_24611,N_24379);
xor UO_1366 (O_1366,N_24908,N_24557);
nor UO_1367 (O_1367,N_24784,N_24921);
nor UO_1368 (O_1368,N_24813,N_24020);
or UO_1369 (O_1369,N_24996,N_24800);
nor UO_1370 (O_1370,N_24845,N_24562);
nor UO_1371 (O_1371,N_24886,N_24376);
xnor UO_1372 (O_1372,N_24728,N_24686);
xor UO_1373 (O_1373,N_24182,N_24689);
xnor UO_1374 (O_1374,N_24709,N_24130);
or UO_1375 (O_1375,N_24780,N_24843);
and UO_1376 (O_1376,N_24316,N_24634);
nand UO_1377 (O_1377,N_24133,N_24446);
and UO_1378 (O_1378,N_24462,N_24630);
nand UO_1379 (O_1379,N_24956,N_24563);
or UO_1380 (O_1380,N_24875,N_24530);
and UO_1381 (O_1381,N_24675,N_24514);
xnor UO_1382 (O_1382,N_24276,N_24495);
nor UO_1383 (O_1383,N_24177,N_24677);
xnor UO_1384 (O_1384,N_24037,N_24766);
xor UO_1385 (O_1385,N_24614,N_24085);
nand UO_1386 (O_1386,N_24044,N_24312);
and UO_1387 (O_1387,N_24700,N_24646);
nand UO_1388 (O_1388,N_24987,N_24048);
nor UO_1389 (O_1389,N_24801,N_24647);
nand UO_1390 (O_1390,N_24192,N_24395);
nor UO_1391 (O_1391,N_24864,N_24026);
and UO_1392 (O_1392,N_24039,N_24470);
xor UO_1393 (O_1393,N_24117,N_24129);
nand UO_1394 (O_1394,N_24097,N_24550);
or UO_1395 (O_1395,N_24850,N_24950);
nor UO_1396 (O_1396,N_24593,N_24024);
nand UO_1397 (O_1397,N_24688,N_24095);
or UO_1398 (O_1398,N_24143,N_24682);
xnor UO_1399 (O_1399,N_24691,N_24325);
nand UO_1400 (O_1400,N_24565,N_24430);
or UO_1401 (O_1401,N_24661,N_24834);
or UO_1402 (O_1402,N_24555,N_24540);
nor UO_1403 (O_1403,N_24101,N_24046);
or UO_1404 (O_1404,N_24849,N_24718);
nor UO_1405 (O_1405,N_24876,N_24599);
and UO_1406 (O_1406,N_24563,N_24725);
or UO_1407 (O_1407,N_24228,N_24549);
or UO_1408 (O_1408,N_24541,N_24193);
xnor UO_1409 (O_1409,N_24856,N_24622);
nor UO_1410 (O_1410,N_24508,N_24178);
or UO_1411 (O_1411,N_24806,N_24281);
nand UO_1412 (O_1412,N_24403,N_24569);
and UO_1413 (O_1413,N_24558,N_24447);
or UO_1414 (O_1414,N_24851,N_24650);
nor UO_1415 (O_1415,N_24749,N_24711);
or UO_1416 (O_1416,N_24440,N_24870);
xnor UO_1417 (O_1417,N_24815,N_24961);
and UO_1418 (O_1418,N_24873,N_24029);
or UO_1419 (O_1419,N_24257,N_24870);
and UO_1420 (O_1420,N_24864,N_24900);
xor UO_1421 (O_1421,N_24535,N_24413);
nor UO_1422 (O_1422,N_24611,N_24102);
nor UO_1423 (O_1423,N_24999,N_24973);
and UO_1424 (O_1424,N_24417,N_24834);
or UO_1425 (O_1425,N_24385,N_24021);
or UO_1426 (O_1426,N_24653,N_24628);
nand UO_1427 (O_1427,N_24875,N_24776);
and UO_1428 (O_1428,N_24256,N_24667);
and UO_1429 (O_1429,N_24580,N_24870);
nor UO_1430 (O_1430,N_24665,N_24364);
nor UO_1431 (O_1431,N_24412,N_24502);
or UO_1432 (O_1432,N_24723,N_24620);
nand UO_1433 (O_1433,N_24691,N_24402);
nand UO_1434 (O_1434,N_24796,N_24983);
xnor UO_1435 (O_1435,N_24872,N_24994);
xnor UO_1436 (O_1436,N_24090,N_24879);
and UO_1437 (O_1437,N_24060,N_24825);
nand UO_1438 (O_1438,N_24311,N_24162);
nand UO_1439 (O_1439,N_24219,N_24792);
xnor UO_1440 (O_1440,N_24493,N_24124);
nand UO_1441 (O_1441,N_24939,N_24807);
and UO_1442 (O_1442,N_24869,N_24045);
xnor UO_1443 (O_1443,N_24573,N_24295);
or UO_1444 (O_1444,N_24942,N_24522);
nor UO_1445 (O_1445,N_24382,N_24964);
nand UO_1446 (O_1446,N_24933,N_24503);
or UO_1447 (O_1447,N_24473,N_24134);
and UO_1448 (O_1448,N_24852,N_24574);
xor UO_1449 (O_1449,N_24539,N_24138);
and UO_1450 (O_1450,N_24724,N_24813);
or UO_1451 (O_1451,N_24953,N_24846);
or UO_1452 (O_1452,N_24343,N_24437);
xnor UO_1453 (O_1453,N_24017,N_24157);
nor UO_1454 (O_1454,N_24003,N_24919);
xor UO_1455 (O_1455,N_24503,N_24768);
nand UO_1456 (O_1456,N_24676,N_24897);
nor UO_1457 (O_1457,N_24794,N_24901);
and UO_1458 (O_1458,N_24852,N_24954);
or UO_1459 (O_1459,N_24546,N_24734);
and UO_1460 (O_1460,N_24768,N_24477);
or UO_1461 (O_1461,N_24833,N_24707);
nor UO_1462 (O_1462,N_24297,N_24696);
nor UO_1463 (O_1463,N_24243,N_24065);
xor UO_1464 (O_1464,N_24461,N_24957);
nor UO_1465 (O_1465,N_24404,N_24955);
and UO_1466 (O_1466,N_24791,N_24799);
and UO_1467 (O_1467,N_24560,N_24248);
or UO_1468 (O_1468,N_24369,N_24179);
nor UO_1469 (O_1469,N_24201,N_24982);
nor UO_1470 (O_1470,N_24678,N_24881);
and UO_1471 (O_1471,N_24908,N_24890);
nor UO_1472 (O_1472,N_24485,N_24027);
or UO_1473 (O_1473,N_24338,N_24854);
and UO_1474 (O_1474,N_24453,N_24820);
and UO_1475 (O_1475,N_24098,N_24163);
nor UO_1476 (O_1476,N_24039,N_24081);
nand UO_1477 (O_1477,N_24398,N_24849);
or UO_1478 (O_1478,N_24245,N_24754);
xor UO_1479 (O_1479,N_24815,N_24449);
or UO_1480 (O_1480,N_24813,N_24429);
nand UO_1481 (O_1481,N_24090,N_24626);
or UO_1482 (O_1482,N_24886,N_24090);
nand UO_1483 (O_1483,N_24742,N_24302);
nand UO_1484 (O_1484,N_24277,N_24350);
and UO_1485 (O_1485,N_24005,N_24734);
and UO_1486 (O_1486,N_24117,N_24552);
and UO_1487 (O_1487,N_24092,N_24489);
and UO_1488 (O_1488,N_24795,N_24333);
nand UO_1489 (O_1489,N_24029,N_24060);
nor UO_1490 (O_1490,N_24477,N_24983);
xnor UO_1491 (O_1491,N_24220,N_24150);
and UO_1492 (O_1492,N_24593,N_24931);
xnor UO_1493 (O_1493,N_24009,N_24234);
nand UO_1494 (O_1494,N_24201,N_24971);
nor UO_1495 (O_1495,N_24432,N_24372);
xnor UO_1496 (O_1496,N_24607,N_24378);
nor UO_1497 (O_1497,N_24602,N_24796);
xnor UO_1498 (O_1498,N_24930,N_24157);
xnor UO_1499 (O_1499,N_24665,N_24401);
or UO_1500 (O_1500,N_24529,N_24569);
and UO_1501 (O_1501,N_24208,N_24643);
or UO_1502 (O_1502,N_24468,N_24675);
and UO_1503 (O_1503,N_24811,N_24344);
or UO_1504 (O_1504,N_24137,N_24005);
nor UO_1505 (O_1505,N_24572,N_24275);
and UO_1506 (O_1506,N_24160,N_24390);
nor UO_1507 (O_1507,N_24857,N_24904);
xor UO_1508 (O_1508,N_24152,N_24520);
nor UO_1509 (O_1509,N_24044,N_24077);
or UO_1510 (O_1510,N_24840,N_24296);
and UO_1511 (O_1511,N_24532,N_24406);
xor UO_1512 (O_1512,N_24548,N_24862);
and UO_1513 (O_1513,N_24088,N_24861);
nand UO_1514 (O_1514,N_24552,N_24499);
nor UO_1515 (O_1515,N_24119,N_24293);
nand UO_1516 (O_1516,N_24020,N_24465);
and UO_1517 (O_1517,N_24918,N_24898);
nand UO_1518 (O_1518,N_24405,N_24219);
nor UO_1519 (O_1519,N_24942,N_24995);
and UO_1520 (O_1520,N_24344,N_24596);
and UO_1521 (O_1521,N_24491,N_24111);
nand UO_1522 (O_1522,N_24594,N_24262);
xor UO_1523 (O_1523,N_24557,N_24294);
nand UO_1524 (O_1524,N_24478,N_24725);
nand UO_1525 (O_1525,N_24052,N_24961);
xor UO_1526 (O_1526,N_24693,N_24759);
or UO_1527 (O_1527,N_24149,N_24251);
or UO_1528 (O_1528,N_24381,N_24495);
nor UO_1529 (O_1529,N_24972,N_24035);
nand UO_1530 (O_1530,N_24161,N_24172);
or UO_1531 (O_1531,N_24721,N_24532);
nand UO_1532 (O_1532,N_24876,N_24877);
nor UO_1533 (O_1533,N_24979,N_24105);
or UO_1534 (O_1534,N_24901,N_24880);
nand UO_1535 (O_1535,N_24497,N_24153);
nor UO_1536 (O_1536,N_24856,N_24892);
nor UO_1537 (O_1537,N_24637,N_24390);
and UO_1538 (O_1538,N_24313,N_24898);
xor UO_1539 (O_1539,N_24386,N_24005);
or UO_1540 (O_1540,N_24048,N_24649);
and UO_1541 (O_1541,N_24136,N_24607);
or UO_1542 (O_1542,N_24589,N_24484);
and UO_1543 (O_1543,N_24887,N_24555);
xnor UO_1544 (O_1544,N_24724,N_24871);
nor UO_1545 (O_1545,N_24166,N_24585);
and UO_1546 (O_1546,N_24339,N_24558);
nor UO_1547 (O_1547,N_24533,N_24502);
nor UO_1548 (O_1548,N_24094,N_24628);
xnor UO_1549 (O_1549,N_24167,N_24550);
xor UO_1550 (O_1550,N_24377,N_24781);
and UO_1551 (O_1551,N_24038,N_24661);
xnor UO_1552 (O_1552,N_24161,N_24875);
xnor UO_1553 (O_1553,N_24502,N_24229);
nor UO_1554 (O_1554,N_24700,N_24618);
and UO_1555 (O_1555,N_24170,N_24418);
and UO_1556 (O_1556,N_24510,N_24553);
xnor UO_1557 (O_1557,N_24068,N_24409);
and UO_1558 (O_1558,N_24629,N_24548);
xnor UO_1559 (O_1559,N_24949,N_24715);
xor UO_1560 (O_1560,N_24223,N_24582);
xor UO_1561 (O_1561,N_24315,N_24290);
nand UO_1562 (O_1562,N_24181,N_24130);
or UO_1563 (O_1563,N_24717,N_24200);
xnor UO_1564 (O_1564,N_24193,N_24951);
nand UO_1565 (O_1565,N_24335,N_24298);
and UO_1566 (O_1566,N_24816,N_24874);
nor UO_1567 (O_1567,N_24269,N_24836);
nor UO_1568 (O_1568,N_24522,N_24376);
nor UO_1569 (O_1569,N_24533,N_24286);
nor UO_1570 (O_1570,N_24414,N_24238);
xor UO_1571 (O_1571,N_24001,N_24973);
nand UO_1572 (O_1572,N_24750,N_24248);
nand UO_1573 (O_1573,N_24083,N_24416);
nor UO_1574 (O_1574,N_24227,N_24488);
nand UO_1575 (O_1575,N_24690,N_24025);
or UO_1576 (O_1576,N_24685,N_24561);
xnor UO_1577 (O_1577,N_24528,N_24147);
and UO_1578 (O_1578,N_24883,N_24801);
xor UO_1579 (O_1579,N_24080,N_24817);
or UO_1580 (O_1580,N_24829,N_24237);
nand UO_1581 (O_1581,N_24564,N_24849);
nand UO_1582 (O_1582,N_24251,N_24147);
and UO_1583 (O_1583,N_24579,N_24788);
nor UO_1584 (O_1584,N_24939,N_24109);
nand UO_1585 (O_1585,N_24696,N_24977);
or UO_1586 (O_1586,N_24412,N_24536);
xnor UO_1587 (O_1587,N_24939,N_24748);
nand UO_1588 (O_1588,N_24803,N_24984);
xnor UO_1589 (O_1589,N_24321,N_24891);
or UO_1590 (O_1590,N_24543,N_24695);
nor UO_1591 (O_1591,N_24298,N_24421);
nand UO_1592 (O_1592,N_24099,N_24354);
nor UO_1593 (O_1593,N_24249,N_24952);
or UO_1594 (O_1594,N_24890,N_24155);
and UO_1595 (O_1595,N_24916,N_24855);
xnor UO_1596 (O_1596,N_24535,N_24343);
nor UO_1597 (O_1597,N_24035,N_24872);
xor UO_1598 (O_1598,N_24936,N_24246);
xor UO_1599 (O_1599,N_24960,N_24713);
or UO_1600 (O_1600,N_24996,N_24997);
and UO_1601 (O_1601,N_24382,N_24640);
and UO_1602 (O_1602,N_24771,N_24060);
nor UO_1603 (O_1603,N_24969,N_24108);
nand UO_1604 (O_1604,N_24615,N_24396);
and UO_1605 (O_1605,N_24632,N_24508);
nand UO_1606 (O_1606,N_24538,N_24473);
nand UO_1607 (O_1607,N_24557,N_24094);
xnor UO_1608 (O_1608,N_24220,N_24909);
nand UO_1609 (O_1609,N_24171,N_24628);
xnor UO_1610 (O_1610,N_24553,N_24400);
nor UO_1611 (O_1611,N_24622,N_24111);
nand UO_1612 (O_1612,N_24469,N_24193);
nor UO_1613 (O_1613,N_24101,N_24907);
and UO_1614 (O_1614,N_24661,N_24863);
xor UO_1615 (O_1615,N_24904,N_24111);
and UO_1616 (O_1616,N_24143,N_24778);
nor UO_1617 (O_1617,N_24093,N_24719);
nand UO_1618 (O_1618,N_24032,N_24041);
nor UO_1619 (O_1619,N_24937,N_24680);
nand UO_1620 (O_1620,N_24751,N_24092);
and UO_1621 (O_1621,N_24152,N_24478);
or UO_1622 (O_1622,N_24373,N_24839);
nand UO_1623 (O_1623,N_24673,N_24905);
and UO_1624 (O_1624,N_24070,N_24784);
xnor UO_1625 (O_1625,N_24750,N_24533);
and UO_1626 (O_1626,N_24780,N_24501);
nor UO_1627 (O_1627,N_24887,N_24772);
xnor UO_1628 (O_1628,N_24786,N_24934);
or UO_1629 (O_1629,N_24580,N_24684);
xor UO_1630 (O_1630,N_24850,N_24074);
or UO_1631 (O_1631,N_24373,N_24248);
xor UO_1632 (O_1632,N_24085,N_24742);
and UO_1633 (O_1633,N_24731,N_24581);
xor UO_1634 (O_1634,N_24458,N_24050);
nand UO_1635 (O_1635,N_24948,N_24586);
nor UO_1636 (O_1636,N_24196,N_24333);
nand UO_1637 (O_1637,N_24524,N_24873);
and UO_1638 (O_1638,N_24497,N_24127);
and UO_1639 (O_1639,N_24333,N_24530);
nand UO_1640 (O_1640,N_24084,N_24103);
xnor UO_1641 (O_1641,N_24596,N_24822);
or UO_1642 (O_1642,N_24970,N_24000);
xor UO_1643 (O_1643,N_24592,N_24485);
nor UO_1644 (O_1644,N_24103,N_24352);
or UO_1645 (O_1645,N_24402,N_24137);
and UO_1646 (O_1646,N_24155,N_24400);
nor UO_1647 (O_1647,N_24045,N_24956);
nor UO_1648 (O_1648,N_24132,N_24029);
and UO_1649 (O_1649,N_24783,N_24145);
and UO_1650 (O_1650,N_24188,N_24305);
or UO_1651 (O_1651,N_24974,N_24087);
and UO_1652 (O_1652,N_24647,N_24281);
or UO_1653 (O_1653,N_24972,N_24788);
xnor UO_1654 (O_1654,N_24754,N_24261);
xor UO_1655 (O_1655,N_24542,N_24393);
and UO_1656 (O_1656,N_24258,N_24270);
nand UO_1657 (O_1657,N_24276,N_24033);
nor UO_1658 (O_1658,N_24773,N_24319);
and UO_1659 (O_1659,N_24973,N_24044);
and UO_1660 (O_1660,N_24054,N_24309);
xnor UO_1661 (O_1661,N_24674,N_24039);
xnor UO_1662 (O_1662,N_24829,N_24551);
nand UO_1663 (O_1663,N_24387,N_24153);
or UO_1664 (O_1664,N_24977,N_24452);
and UO_1665 (O_1665,N_24005,N_24717);
xnor UO_1666 (O_1666,N_24622,N_24525);
or UO_1667 (O_1667,N_24997,N_24902);
nand UO_1668 (O_1668,N_24614,N_24499);
nor UO_1669 (O_1669,N_24668,N_24422);
or UO_1670 (O_1670,N_24782,N_24021);
nor UO_1671 (O_1671,N_24000,N_24421);
nor UO_1672 (O_1672,N_24456,N_24143);
xnor UO_1673 (O_1673,N_24340,N_24001);
nor UO_1674 (O_1674,N_24221,N_24344);
xor UO_1675 (O_1675,N_24257,N_24073);
and UO_1676 (O_1676,N_24389,N_24602);
nor UO_1677 (O_1677,N_24780,N_24623);
nor UO_1678 (O_1678,N_24029,N_24890);
nand UO_1679 (O_1679,N_24938,N_24641);
or UO_1680 (O_1680,N_24254,N_24689);
or UO_1681 (O_1681,N_24542,N_24680);
nor UO_1682 (O_1682,N_24579,N_24954);
nand UO_1683 (O_1683,N_24827,N_24642);
xor UO_1684 (O_1684,N_24029,N_24040);
nor UO_1685 (O_1685,N_24846,N_24848);
xor UO_1686 (O_1686,N_24064,N_24540);
and UO_1687 (O_1687,N_24254,N_24241);
nand UO_1688 (O_1688,N_24572,N_24618);
or UO_1689 (O_1689,N_24342,N_24159);
and UO_1690 (O_1690,N_24290,N_24573);
or UO_1691 (O_1691,N_24684,N_24739);
and UO_1692 (O_1692,N_24819,N_24512);
xnor UO_1693 (O_1693,N_24597,N_24395);
xnor UO_1694 (O_1694,N_24467,N_24082);
nand UO_1695 (O_1695,N_24338,N_24942);
or UO_1696 (O_1696,N_24694,N_24925);
xor UO_1697 (O_1697,N_24307,N_24847);
nor UO_1698 (O_1698,N_24125,N_24210);
nor UO_1699 (O_1699,N_24821,N_24767);
xnor UO_1700 (O_1700,N_24915,N_24916);
or UO_1701 (O_1701,N_24558,N_24987);
nand UO_1702 (O_1702,N_24062,N_24490);
or UO_1703 (O_1703,N_24370,N_24653);
nor UO_1704 (O_1704,N_24371,N_24274);
nand UO_1705 (O_1705,N_24876,N_24741);
nor UO_1706 (O_1706,N_24508,N_24496);
xnor UO_1707 (O_1707,N_24609,N_24410);
nand UO_1708 (O_1708,N_24332,N_24817);
nand UO_1709 (O_1709,N_24838,N_24713);
nand UO_1710 (O_1710,N_24051,N_24036);
or UO_1711 (O_1711,N_24831,N_24736);
or UO_1712 (O_1712,N_24894,N_24593);
and UO_1713 (O_1713,N_24665,N_24880);
xor UO_1714 (O_1714,N_24418,N_24906);
and UO_1715 (O_1715,N_24703,N_24606);
xor UO_1716 (O_1716,N_24140,N_24310);
and UO_1717 (O_1717,N_24113,N_24229);
xnor UO_1718 (O_1718,N_24589,N_24351);
nor UO_1719 (O_1719,N_24164,N_24229);
nor UO_1720 (O_1720,N_24222,N_24580);
or UO_1721 (O_1721,N_24544,N_24185);
or UO_1722 (O_1722,N_24365,N_24377);
xor UO_1723 (O_1723,N_24428,N_24420);
xnor UO_1724 (O_1724,N_24440,N_24558);
or UO_1725 (O_1725,N_24670,N_24994);
and UO_1726 (O_1726,N_24196,N_24017);
and UO_1727 (O_1727,N_24364,N_24547);
and UO_1728 (O_1728,N_24782,N_24325);
nand UO_1729 (O_1729,N_24643,N_24509);
nor UO_1730 (O_1730,N_24405,N_24065);
nand UO_1731 (O_1731,N_24827,N_24629);
nor UO_1732 (O_1732,N_24947,N_24426);
xor UO_1733 (O_1733,N_24729,N_24063);
or UO_1734 (O_1734,N_24058,N_24095);
nand UO_1735 (O_1735,N_24972,N_24682);
and UO_1736 (O_1736,N_24899,N_24995);
and UO_1737 (O_1737,N_24657,N_24741);
nor UO_1738 (O_1738,N_24582,N_24255);
nand UO_1739 (O_1739,N_24342,N_24216);
or UO_1740 (O_1740,N_24570,N_24896);
and UO_1741 (O_1741,N_24763,N_24408);
or UO_1742 (O_1742,N_24408,N_24130);
nor UO_1743 (O_1743,N_24926,N_24696);
nor UO_1744 (O_1744,N_24254,N_24084);
and UO_1745 (O_1745,N_24200,N_24255);
and UO_1746 (O_1746,N_24490,N_24257);
xnor UO_1747 (O_1747,N_24173,N_24338);
xnor UO_1748 (O_1748,N_24669,N_24325);
and UO_1749 (O_1749,N_24581,N_24703);
nor UO_1750 (O_1750,N_24212,N_24523);
xnor UO_1751 (O_1751,N_24245,N_24732);
nor UO_1752 (O_1752,N_24986,N_24655);
or UO_1753 (O_1753,N_24739,N_24308);
nand UO_1754 (O_1754,N_24858,N_24254);
nor UO_1755 (O_1755,N_24714,N_24219);
and UO_1756 (O_1756,N_24343,N_24037);
nand UO_1757 (O_1757,N_24573,N_24373);
nor UO_1758 (O_1758,N_24085,N_24247);
nand UO_1759 (O_1759,N_24470,N_24248);
or UO_1760 (O_1760,N_24189,N_24014);
xor UO_1761 (O_1761,N_24964,N_24603);
xnor UO_1762 (O_1762,N_24329,N_24484);
nand UO_1763 (O_1763,N_24251,N_24273);
or UO_1764 (O_1764,N_24773,N_24618);
or UO_1765 (O_1765,N_24797,N_24422);
nand UO_1766 (O_1766,N_24698,N_24615);
nand UO_1767 (O_1767,N_24635,N_24852);
nand UO_1768 (O_1768,N_24412,N_24372);
nand UO_1769 (O_1769,N_24158,N_24436);
xnor UO_1770 (O_1770,N_24902,N_24343);
nor UO_1771 (O_1771,N_24557,N_24234);
or UO_1772 (O_1772,N_24096,N_24431);
nand UO_1773 (O_1773,N_24385,N_24722);
nand UO_1774 (O_1774,N_24270,N_24890);
and UO_1775 (O_1775,N_24766,N_24357);
nor UO_1776 (O_1776,N_24021,N_24176);
or UO_1777 (O_1777,N_24494,N_24920);
and UO_1778 (O_1778,N_24117,N_24464);
xnor UO_1779 (O_1779,N_24740,N_24221);
xnor UO_1780 (O_1780,N_24314,N_24260);
and UO_1781 (O_1781,N_24947,N_24364);
or UO_1782 (O_1782,N_24555,N_24266);
and UO_1783 (O_1783,N_24341,N_24575);
nand UO_1784 (O_1784,N_24072,N_24249);
xor UO_1785 (O_1785,N_24133,N_24636);
nor UO_1786 (O_1786,N_24625,N_24349);
and UO_1787 (O_1787,N_24267,N_24866);
and UO_1788 (O_1788,N_24106,N_24612);
nand UO_1789 (O_1789,N_24088,N_24629);
and UO_1790 (O_1790,N_24681,N_24784);
nand UO_1791 (O_1791,N_24217,N_24937);
nor UO_1792 (O_1792,N_24051,N_24118);
xnor UO_1793 (O_1793,N_24785,N_24280);
or UO_1794 (O_1794,N_24896,N_24546);
nor UO_1795 (O_1795,N_24603,N_24045);
and UO_1796 (O_1796,N_24727,N_24673);
xnor UO_1797 (O_1797,N_24423,N_24041);
or UO_1798 (O_1798,N_24606,N_24969);
nand UO_1799 (O_1799,N_24356,N_24627);
xnor UO_1800 (O_1800,N_24459,N_24879);
nor UO_1801 (O_1801,N_24893,N_24529);
xor UO_1802 (O_1802,N_24566,N_24875);
nand UO_1803 (O_1803,N_24019,N_24967);
nand UO_1804 (O_1804,N_24214,N_24610);
xnor UO_1805 (O_1805,N_24928,N_24171);
or UO_1806 (O_1806,N_24183,N_24772);
nand UO_1807 (O_1807,N_24399,N_24044);
and UO_1808 (O_1808,N_24847,N_24516);
nor UO_1809 (O_1809,N_24487,N_24636);
nor UO_1810 (O_1810,N_24711,N_24356);
or UO_1811 (O_1811,N_24265,N_24097);
and UO_1812 (O_1812,N_24242,N_24654);
nand UO_1813 (O_1813,N_24516,N_24088);
and UO_1814 (O_1814,N_24215,N_24534);
nand UO_1815 (O_1815,N_24579,N_24798);
nor UO_1816 (O_1816,N_24841,N_24906);
or UO_1817 (O_1817,N_24896,N_24927);
and UO_1818 (O_1818,N_24599,N_24532);
nor UO_1819 (O_1819,N_24535,N_24344);
nor UO_1820 (O_1820,N_24837,N_24343);
or UO_1821 (O_1821,N_24970,N_24255);
nor UO_1822 (O_1822,N_24078,N_24635);
or UO_1823 (O_1823,N_24775,N_24526);
nor UO_1824 (O_1824,N_24609,N_24778);
and UO_1825 (O_1825,N_24831,N_24673);
and UO_1826 (O_1826,N_24157,N_24998);
nand UO_1827 (O_1827,N_24575,N_24398);
and UO_1828 (O_1828,N_24601,N_24116);
nor UO_1829 (O_1829,N_24224,N_24127);
and UO_1830 (O_1830,N_24002,N_24372);
and UO_1831 (O_1831,N_24605,N_24956);
nand UO_1832 (O_1832,N_24883,N_24310);
nor UO_1833 (O_1833,N_24077,N_24166);
or UO_1834 (O_1834,N_24017,N_24927);
nor UO_1835 (O_1835,N_24355,N_24630);
or UO_1836 (O_1836,N_24158,N_24676);
or UO_1837 (O_1837,N_24496,N_24996);
nand UO_1838 (O_1838,N_24867,N_24659);
nor UO_1839 (O_1839,N_24319,N_24075);
or UO_1840 (O_1840,N_24265,N_24572);
nand UO_1841 (O_1841,N_24409,N_24997);
or UO_1842 (O_1842,N_24322,N_24018);
nand UO_1843 (O_1843,N_24273,N_24657);
or UO_1844 (O_1844,N_24928,N_24247);
nand UO_1845 (O_1845,N_24619,N_24928);
nand UO_1846 (O_1846,N_24103,N_24730);
nor UO_1847 (O_1847,N_24056,N_24002);
and UO_1848 (O_1848,N_24163,N_24195);
nor UO_1849 (O_1849,N_24325,N_24838);
or UO_1850 (O_1850,N_24052,N_24531);
or UO_1851 (O_1851,N_24232,N_24726);
or UO_1852 (O_1852,N_24553,N_24600);
nand UO_1853 (O_1853,N_24700,N_24884);
nand UO_1854 (O_1854,N_24108,N_24239);
nand UO_1855 (O_1855,N_24105,N_24589);
and UO_1856 (O_1856,N_24867,N_24324);
nand UO_1857 (O_1857,N_24979,N_24779);
and UO_1858 (O_1858,N_24233,N_24594);
or UO_1859 (O_1859,N_24033,N_24034);
nand UO_1860 (O_1860,N_24101,N_24311);
xnor UO_1861 (O_1861,N_24945,N_24054);
nor UO_1862 (O_1862,N_24713,N_24346);
and UO_1863 (O_1863,N_24318,N_24524);
nor UO_1864 (O_1864,N_24909,N_24433);
nand UO_1865 (O_1865,N_24906,N_24005);
nand UO_1866 (O_1866,N_24293,N_24852);
or UO_1867 (O_1867,N_24094,N_24648);
xnor UO_1868 (O_1868,N_24155,N_24876);
and UO_1869 (O_1869,N_24579,N_24468);
or UO_1870 (O_1870,N_24926,N_24198);
and UO_1871 (O_1871,N_24742,N_24464);
nand UO_1872 (O_1872,N_24131,N_24637);
xnor UO_1873 (O_1873,N_24779,N_24008);
nor UO_1874 (O_1874,N_24236,N_24908);
or UO_1875 (O_1875,N_24531,N_24330);
xor UO_1876 (O_1876,N_24879,N_24761);
xor UO_1877 (O_1877,N_24299,N_24881);
xnor UO_1878 (O_1878,N_24661,N_24928);
and UO_1879 (O_1879,N_24815,N_24090);
nor UO_1880 (O_1880,N_24862,N_24432);
nor UO_1881 (O_1881,N_24359,N_24795);
or UO_1882 (O_1882,N_24641,N_24772);
or UO_1883 (O_1883,N_24864,N_24975);
nand UO_1884 (O_1884,N_24484,N_24934);
nor UO_1885 (O_1885,N_24430,N_24082);
nor UO_1886 (O_1886,N_24422,N_24826);
and UO_1887 (O_1887,N_24375,N_24518);
nor UO_1888 (O_1888,N_24372,N_24332);
and UO_1889 (O_1889,N_24905,N_24189);
nand UO_1890 (O_1890,N_24985,N_24861);
or UO_1891 (O_1891,N_24749,N_24320);
and UO_1892 (O_1892,N_24746,N_24524);
or UO_1893 (O_1893,N_24744,N_24205);
or UO_1894 (O_1894,N_24803,N_24118);
and UO_1895 (O_1895,N_24157,N_24043);
xnor UO_1896 (O_1896,N_24962,N_24738);
or UO_1897 (O_1897,N_24023,N_24682);
and UO_1898 (O_1898,N_24553,N_24611);
xor UO_1899 (O_1899,N_24938,N_24716);
or UO_1900 (O_1900,N_24308,N_24836);
nor UO_1901 (O_1901,N_24830,N_24592);
or UO_1902 (O_1902,N_24120,N_24543);
nor UO_1903 (O_1903,N_24901,N_24124);
or UO_1904 (O_1904,N_24493,N_24400);
or UO_1905 (O_1905,N_24084,N_24710);
or UO_1906 (O_1906,N_24146,N_24622);
nand UO_1907 (O_1907,N_24705,N_24743);
or UO_1908 (O_1908,N_24860,N_24290);
and UO_1909 (O_1909,N_24397,N_24361);
and UO_1910 (O_1910,N_24883,N_24331);
nor UO_1911 (O_1911,N_24395,N_24614);
nor UO_1912 (O_1912,N_24851,N_24249);
xnor UO_1913 (O_1913,N_24984,N_24112);
nor UO_1914 (O_1914,N_24014,N_24653);
xnor UO_1915 (O_1915,N_24580,N_24038);
or UO_1916 (O_1916,N_24837,N_24269);
nor UO_1917 (O_1917,N_24928,N_24796);
nand UO_1918 (O_1918,N_24415,N_24819);
xnor UO_1919 (O_1919,N_24581,N_24839);
nor UO_1920 (O_1920,N_24326,N_24044);
nor UO_1921 (O_1921,N_24906,N_24069);
nand UO_1922 (O_1922,N_24507,N_24607);
nor UO_1923 (O_1923,N_24584,N_24776);
or UO_1924 (O_1924,N_24431,N_24483);
xnor UO_1925 (O_1925,N_24563,N_24666);
or UO_1926 (O_1926,N_24538,N_24253);
nand UO_1927 (O_1927,N_24615,N_24538);
nor UO_1928 (O_1928,N_24341,N_24717);
nor UO_1929 (O_1929,N_24613,N_24290);
xnor UO_1930 (O_1930,N_24989,N_24890);
nand UO_1931 (O_1931,N_24869,N_24647);
nand UO_1932 (O_1932,N_24337,N_24285);
and UO_1933 (O_1933,N_24117,N_24666);
xor UO_1934 (O_1934,N_24719,N_24401);
nor UO_1935 (O_1935,N_24860,N_24244);
xnor UO_1936 (O_1936,N_24561,N_24585);
xor UO_1937 (O_1937,N_24239,N_24389);
or UO_1938 (O_1938,N_24026,N_24029);
or UO_1939 (O_1939,N_24354,N_24195);
or UO_1940 (O_1940,N_24663,N_24210);
nor UO_1941 (O_1941,N_24901,N_24321);
and UO_1942 (O_1942,N_24915,N_24564);
and UO_1943 (O_1943,N_24311,N_24862);
nand UO_1944 (O_1944,N_24093,N_24790);
xnor UO_1945 (O_1945,N_24316,N_24225);
nor UO_1946 (O_1946,N_24261,N_24439);
or UO_1947 (O_1947,N_24668,N_24904);
and UO_1948 (O_1948,N_24233,N_24798);
nor UO_1949 (O_1949,N_24099,N_24397);
nand UO_1950 (O_1950,N_24978,N_24339);
nor UO_1951 (O_1951,N_24547,N_24457);
or UO_1952 (O_1952,N_24325,N_24104);
xor UO_1953 (O_1953,N_24917,N_24486);
nor UO_1954 (O_1954,N_24096,N_24999);
or UO_1955 (O_1955,N_24103,N_24189);
or UO_1956 (O_1956,N_24133,N_24058);
nand UO_1957 (O_1957,N_24931,N_24462);
or UO_1958 (O_1958,N_24538,N_24983);
and UO_1959 (O_1959,N_24596,N_24342);
xnor UO_1960 (O_1960,N_24866,N_24538);
nand UO_1961 (O_1961,N_24291,N_24380);
nand UO_1962 (O_1962,N_24051,N_24239);
xnor UO_1963 (O_1963,N_24035,N_24440);
and UO_1964 (O_1964,N_24628,N_24003);
nand UO_1965 (O_1965,N_24915,N_24574);
nand UO_1966 (O_1966,N_24571,N_24545);
or UO_1967 (O_1967,N_24683,N_24780);
and UO_1968 (O_1968,N_24260,N_24706);
xnor UO_1969 (O_1969,N_24228,N_24834);
and UO_1970 (O_1970,N_24182,N_24835);
nand UO_1971 (O_1971,N_24176,N_24117);
and UO_1972 (O_1972,N_24706,N_24661);
xnor UO_1973 (O_1973,N_24121,N_24088);
nand UO_1974 (O_1974,N_24680,N_24517);
xor UO_1975 (O_1975,N_24487,N_24499);
xor UO_1976 (O_1976,N_24887,N_24084);
xnor UO_1977 (O_1977,N_24652,N_24772);
or UO_1978 (O_1978,N_24283,N_24565);
or UO_1979 (O_1979,N_24875,N_24909);
nand UO_1980 (O_1980,N_24700,N_24742);
nand UO_1981 (O_1981,N_24619,N_24316);
nor UO_1982 (O_1982,N_24987,N_24499);
and UO_1983 (O_1983,N_24556,N_24561);
and UO_1984 (O_1984,N_24486,N_24195);
nor UO_1985 (O_1985,N_24245,N_24597);
xor UO_1986 (O_1986,N_24970,N_24589);
nand UO_1987 (O_1987,N_24667,N_24656);
and UO_1988 (O_1988,N_24619,N_24779);
nand UO_1989 (O_1989,N_24555,N_24267);
or UO_1990 (O_1990,N_24340,N_24156);
xnor UO_1991 (O_1991,N_24620,N_24350);
nand UO_1992 (O_1992,N_24714,N_24958);
or UO_1993 (O_1993,N_24900,N_24345);
nand UO_1994 (O_1994,N_24419,N_24488);
xnor UO_1995 (O_1995,N_24077,N_24898);
and UO_1996 (O_1996,N_24220,N_24984);
nor UO_1997 (O_1997,N_24267,N_24271);
nor UO_1998 (O_1998,N_24832,N_24852);
xor UO_1999 (O_1999,N_24397,N_24448);
nor UO_2000 (O_2000,N_24647,N_24035);
nand UO_2001 (O_2001,N_24476,N_24803);
or UO_2002 (O_2002,N_24395,N_24997);
nor UO_2003 (O_2003,N_24253,N_24090);
nand UO_2004 (O_2004,N_24329,N_24371);
and UO_2005 (O_2005,N_24824,N_24622);
xnor UO_2006 (O_2006,N_24291,N_24951);
or UO_2007 (O_2007,N_24692,N_24764);
and UO_2008 (O_2008,N_24664,N_24810);
nor UO_2009 (O_2009,N_24982,N_24964);
and UO_2010 (O_2010,N_24232,N_24335);
or UO_2011 (O_2011,N_24088,N_24917);
or UO_2012 (O_2012,N_24561,N_24718);
and UO_2013 (O_2013,N_24274,N_24919);
or UO_2014 (O_2014,N_24499,N_24512);
nor UO_2015 (O_2015,N_24796,N_24642);
or UO_2016 (O_2016,N_24477,N_24924);
and UO_2017 (O_2017,N_24490,N_24362);
xnor UO_2018 (O_2018,N_24447,N_24201);
and UO_2019 (O_2019,N_24266,N_24762);
nand UO_2020 (O_2020,N_24245,N_24259);
and UO_2021 (O_2021,N_24205,N_24038);
xor UO_2022 (O_2022,N_24992,N_24207);
and UO_2023 (O_2023,N_24921,N_24415);
nor UO_2024 (O_2024,N_24504,N_24285);
and UO_2025 (O_2025,N_24892,N_24100);
nand UO_2026 (O_2026,N_24667,N_24738);
nand UO_2027 (O_2027,N_24404,N_24621);
or UO_2028 (O_2028,N_24369,N_24789);
xnor UO_2029 (O_2029,N_24175,N_24431);
xnor UO_2030 (O_2030,N_24774,N_24405);
or UO_2031 (O_2031,N_24829,N_24345);
and UO_2032 (O_2032,N_24863,N_24999);
xor UO_2033 (O_2033,N_24262,N_24012);
or UO_2034 (O_2034,N_24109,N_24634);
and UO_2035 (O_2035,N_24331,N_24373);
nand UO_2036 (O_2036,N_24473,N_24092);
xnor UO_2037 (O_2037,N_24410,N_24117);
xnor UO_2038 (O_2038,N_24996,N_24392);
nor UO_2039 (O_2039,N_24064,N_24664);
nor UO_2040 (O_2040,N_24169,N_24521);
and UO_2041 (O_2041,N_24646,N_24197);
or UO_2042 (O_2042,N_24588,N_24802);
and UO_2043 (O_2043,N_24305,N_24936);
nor UO_2044 (O_2044,N_24928,N_24462);
and UO_2045 (O_2045,N_24234,N_24540);
nor UO_2046 (O_2046,N_24686,N_24875);
xnor UO_2047 (O_2047,N_24349,N_24099);
and UO_2048 (O_2048,N_24394,N_24925);
and UO_2049 (O_2049,N_24413,N_24717);
nand UO_2050 (O_2050,N_24874,N_24262);
nand UO_2051 (O_2051,N_24896,N_24483);
and UO_2052 (O_2052,N_24877,N_24167);
nor UO_2053 (O_2053,N_24975,N_24924);
nand UO_2054 (O_2054,N_24106,N_24109);
or UO_2055 (O_2055,N_24573,N_24806);
nand UO_2056 (O_2056,N_24868,N_24870);
and UO_2057 (O_2057,N_24153,N_24812);
and UO_2058 (O_2058,N_24138,N_24323);
and UO_2059 (O_2059,N_24215,N_24412);
nand UO_2060 (O_2060,N_24881,N_24557);
or UO_2061 (O_2061,N_24223,N_24300);
nor UO_2062 (O_2062,N_24852,N_24219);
nor UO_2063 (O_2063,N_24937,N_24812);
nand UO_2064 (O_2064,N_24535,N_24448);
and UO_2065 (O_2065,N_24564,N_24598);
nor UO_2066 (O_2066,N_24672,N_24349);
nor UO_2067 (O_2067,N_24276,N_24623);
nand UO_2068 (O_2068,N_24913,N_24122);
xnor UO_2069 (O_2069,N_24791,N_24955);
and UO_2070 (O_2070,N_24595,N_24530);
and UO_2071 (O_2071,N_24683,N_24236);
and UO_2072 (O_2072,N_24125,N_24533);
nand UO_2073 (O_2073,N_24099,N_24252);
nor UO_2074 (O_2074,N_24232,N_24607);
or UO_2075 (O_2075,N_24015,N_24798);
or UO_2076 (O_2076,N_24566,N_24655);
nand UO_2077 (O_2077,N_24414,N_24146);
xnor UO_2078 (O_2078,N_24094,N_24096);
xor UO_2079 (O_2079,N_24278,N_24673);
nand UO_2080 (O_2080,N_24774,N_24286);
xnor UO_2081 (O_2081,N_24710,N_24599);
nor UO_2082 (O_2082,N_24942,N_24343);
nor UO_2083 (O_2083,N_24904,N_24359);
nor UO_2084 (O_2084,N_24934,N_24204);
and UO_2085 (O_2085,N_24970,N_24656);
and UO_2086 (O_2086,N_24439,N_24000);
nand UO_2087 (O_2087,N_24663,N_24615);
nor UO_2088 (O_2088,N_24774,N_24914);
nand UO_2089 (O_2089,N_24239,N_24280);
xor UO_2090 (O_2090,N_24714,N_24872);
xor UO_2091 (O_2091,N_24634,N_24982);
xnor UO_2092 (O_2092,N_24870,N_24704);
and UO_2093 (O_2093,N_24997,N_24526);
nor UO_2094 (O_2094,N_24100,N_24882);
xnor UO_2095 (O_2095,N_24191,N_24400);
and UO_2096 (O_2096,N_24367,N_24105);
xor UO_2097 (O_2097,N_24222,N_24872);
or UO_2098 (O_2098,N_24430,N_24196);
nand UO_2099 (O_2099,N_24037,N_24877);
xnor UO_2100 (O_2100,N_24966,N_24423);
and UO_2101 (O_2101,N_24029,N_24282);
nor UO_2102 (O_2102,N_24586,N_24216);
nand UO_2103 (O_2103,N_24821,N_24807);
or UO_2104 (O_2104,N_24953,N_24836);
nand UO_2105 (O_2105,N_24962,N_24676);
nor UO_2106 (O_2106,N_24368,N_24483);
nor UO_2107 (O_2107,N_24839,N_24023);
xnor UO_2108 (O_2108,N_24200,N_24662);
and UO_2109 (O_2109,N_24032,N_24703);
nor UO_2110 (O_2110,N_24269,N_24895);
and UO_2111 (O_2111,N_24863,N_24299);
nand UO_2112 (O_2112,N_24857,N_24792);
xnor UO_2113 (O_2113,N_24300,N_24038);
nand UO_2114 (O_2114,N_24830,N_24220);
and UO_2115 (O_2115,N_24059,N_24104);
or UO_2116 (O_2116,N_24526,N_24742);
xnor UO_2117 (O_2117,N_24218,N_24239);
or UO_2118 (O_2118,N_24836,N_24321);
xor UO_2119 (O_2119,N_24418,N_24121);
xnor UO_2120 (O_2120,N_24382,N_24454);
nor UO_2121 (O_2121,N_24340,N_24637);
nand UO_2122 (O_2122,N_24961,N_24050);
or UO_2123 (O_2123,N_24883,N_24621);
nand UO_2124 (O_2124,N_24956,N_24229);
xnor UO_2125 (O_2125,N_24069,N_24897);
and UO_2126 (O_2126,N_24890,N_24092);
nor UO_2127 (O_2127,N_24706,N_24715);
xor UO_2128 (O_2128,N_24341,N_24674);
nand UO_2129 (O_2129,N_24214,N_24158);
xnor UO_2130 (O_2130,N_24197,N_24909);
nand UO_2131 (O_2131,N_24744,N_24997);
xor UO_2132 (O_2132,N_24071,N_24331);
or UO_2133 (O_2133,N_24306,N_24368);
nand UO_2134 (O_2134,N_24569,N_24915);
and UO_2135 (O_2135,N_24935,N_24897);
or UO_2136 (O_2136,N_24928,N_24238);
or UO_2137 (O_2137,N_24957,N_24198);
and UO_2138 (O_2138,N_24940,N_24004);
nor UO_2139 (O_2139,N_24636,N_24194);
and UO_2140 (O_2140,N_24492,N_24037);
xor UO_2141 (O_2141,N_24159,N_24223);
xor UO_2142 (O_2142,N_24851,N_24965);
or UO_2143 (O_2143,N_24830,N_24872);
and UO_2144 (O_2144,N_24510,N_24036);
nand UO_2145 (O_2145,N_24356,N_24614);
or UO_2146 (O_2146,N_24854,N_24525);
nor UO_2147 (O_2147,N_24061,N_24117);
or UO_2148 (O_2148,N_24978,N_24837);
and UO_2149 (O_2149,N_24857,N_24108);
or UO_2150 (O_2150,N_24944,N_24053);
nor UO_2151 (O_2151,N_24067,N_24465);
or UO_2152 (O_2152,N_24448,N_24906);
and UO_2153 (O_2153,N_24192,N_24770);
nor UO_2154 (O_2154,N_24124,N_24229);
nand UO_2155 (O_2155,N_24341,N_24197);
nor UO_2156 (O_2156,N_24229,N_24964);
nand UO_2157 (O_2157,N_24492,N_24746);
nor UO_2158 (O_2158,N_24893,N_24289);
and UO_2159 (O_2159,N_24303,N_24210);
nand UO_2160 (O_2160,N_24636,N_24042);
xor UO_2161 (O_2161,N_24117,N_24233);
nor UO_2162 (O_2162,N_24037,N_24838);
nor UO_2163 (O_2163,N_24915,N_24135);
or UO_2164 (O_2164,N_24208,N_24406);
nand UO_2165 (O_2165,N_24971,N_24121);
and UO_2166 (O_2166,N_24957,N_24363);
or UO_2167 (O_2167,N_24135,N_24219);
xnor UO_2168 (O_2168,N_24007,N_24587);
xor UO_2169 (O_2169,N_24783,N_24021);
xor UO_2170 (O_2170,N_24564,N_24702);
xnor UO_2171 (O_2171,N_24320,N_24149);
nand UO_2172 (O_2172,N_24021,N_24198);
nor UO_2173 (O_2173,N_24413,N_24335);
xnor UO_2174 (O_2174,N_24836,N_24375);
xor UO_2175 (O_2175,N_24108,N_24569);
nand UO_2176 (O_2176,N_24859,N_24368);
xor UO_2177 (O_2177,N_24440,N_24234);
xnor UO_2178 (O_2178,N_24340,N_24788);
xor UO_2179 (O_2179,N_24222,N_24001);
xnor UO_2180 (O_2180,N_24005,N_24368);
nand UO_2181 (O_2181,N_24263,N_24286);
nor UO_2182 (O_2182,N_24399,N_24773);
xnor UO_2183 (O_2183,N_24210,N_24327);
or UO_2184 (O_2184,N_24615,N_24452);
xor UO_2185 (O_2185,N_24059,N_24798);
xnor UO_2186 (O_2186,N_24233,N_24659);
and UO_2187 (O_2187,N_24758,N_24533);
xnor UO_2188 (O_2188,N_24310,N_24791);
xor UO_2189 (O_2189,N_24470,N_24088);
or UO_2190 (O_2190,N_24170,N_24589);
nor UO_2191 (O_2191,N_24188,N_24963);
nor UO_2192 (O_2192,N_24286,N_24930);
nand UO_2193 (O_2193,N_24168,N_24719);
or UO_2194 (O_2194,N_24434,N_24545);
nor UO_2195 (O_2195,N_24863,N_24883);
xor UO_2196 (O_2196,N_24180,N_24132);
nor UO_2197 (O_2197,N_24547,N_24356);
xor UO_2198 (O_2198,N_24921,N_24998);
nand UO_2199 (O_2199,N_24185,N_24312);
and UO_2200 (O_2200,N_24155,N_24344);
and UO_2201 (O_2201,N_24077,N_24928);
xor UO_2202 (O_2202,N_24095,N_24001);
or UO_2203 (O_2203,N_24241,N_24618);
nand UO_2204 (O_2204,N_24878,N_24627);
nor UO_2205 (O_2205,N_24759,N_24228);
xor UO_2206 (O_2206,N_24994,N_24552);
or UO_2207 (O_2207,N_24524,N_24901);
or UO_2208 (O_2208,N_24618,N_24841);
nor UO_2209 (O_2209,N_24294,N_24583);
nor UO_2210 (O_2210,N_24250,N_24577);
nand UO_2211 (O_2211,N_24226,N_24325);
and UO_2212 (O_2212,N_24704,N_24031);
or UO_2213 (O_2213,N_24637,N_24908);
and UO_2214 (O_2214,N_24639,N_24636);
or UO_2215 (O_2215,N_24824,N_24956);
nor UO_2216 (O_2216,N_24410,N_24009);
nand UO_2217 (O_2217,N_24000,N_24551);
or UO_2218 (O_2218,N_24087,N_24403);
nor UO_2219 (O_2219,N_24022,N_24901);
and UO_2220 (O_2220,N_24536,N_24947);
nand UO_2221 (O_2221,N_24751,N_24335);
xnor UO_2222 (O_2222,N_24591,N_24839);
nand UO_2223 (O_2223,N_24890,N_24897);
nand UO_2224 (O_2224,N_24261,N_24454);
xor UO_2225 (O_2225,N_24951,N_24933);
or UO_2226 (O_2226,N_24040,N_24664);
nor UO_2227 (O_2227,N_24322,N_24399);
and UO_2228 (O_2228,N_24533,N_24535);
nand UO_2229 (O_2229,N_24621,N_24098);
nand UO_2230 (O_2230,N_24765,N_24560);
xor UO_2231 (O_2231,N_24412,N_24638);
xor UO_2232 (O_2232,N_24634,N_24189);
and UO_2233 (O_2233,N_24698,N_24169);
and UO_2234 (O_2234,N_24169,N_24723);
xnor UO_2235 (O_2235,N_24551,N_24875);
nand UO_2236 (O_2236,N_24368,N_24717);
nor UO_2237 (O_2237,N_24936,N_24948);
nor UO_2238 (O_2238,N_24600,N_24780);
and UO_2239 (O_2239,N_24207,N_24867);
nor UO_2240 (O_2240,N_24195,N_24176);
and UO_2241 (O_2241,N_24044,N_24851);
nand UO_2242 (O_2242,N_24446,N_24616);
or UO_2243 (O_2243,N_24676,N_24847);
nor UO_2244 (O_2244,N_24688,N_24813);
xor UO_2245 (O_2245,N_24833,N_24495);
or UO_2246 (O_2246,N_24154,N_24599);
nor UO_2247 (O_2247,N_24448,N_24707);
xor UO_2248 (O_2248,N_24527,N_24468);
or UO_2249 (O_2249,N_24499,N_24677);
nor UO_2250 (O_2250,N_24785,N_24497);
and UO_2251 (O_2251,N_24298,N_24984);
and UO_2252 (O_2252,N_24070,N_24696);
nand UO_2253 (O_2253,N_24179,N_24344);
nand UO_2254 (O_2254,N_24317,N_24820);
or UO_2255 (O_2255,N_24864,N_24101);
nand UO_2256 (O_2256,N_24915,N_24197);
or UO_2257 (O_2257,N_24504,N_24433);
and UO_2258 (O_2258,N_24158,N_24911);
nor UO_2259 (O_2259,N_24934,N_24328);
nor UO_2260 (O_2260,N_24948,N_24227);
and UO_2261 (O_2261,N_24650,N_24919);
or UO_2262 (O_2262,N_24023,N_24601);
nand UO_2263 (O_2263,N_24843,N_24295);
and UO_2264 (O_2264,N_24874,N_24122);
xor UO_2265 (O_2265,N_24638,N_24429);
or UO_2266 (O_2266,N_24455,N_24642);
xnor UO_2267 (O_2267,N_24054,N_24299);
nor UO_2268 (O_2268,N_24204,N_24461);
and UO_2269 (O_2269,N_24475,N_24076);
nand UO_2270 (O_2270,N_24695,N_24236);
and UO_2271 (O_2271,N_24016,N_24721);
nor UO_2272 (O_2272,N_24884,N_24366);
or UO_2273 (O_2273,N_24836,N_24495);
or UO_2274 (O_2274,N_24321,N_24973);
nor UO_2275 (O_2275,N_24137,N_24152);
nor UO_2276 (O_2276,N_24701,N_24361);
nor UO_2277 (O_2277,N_24948,N_24687);
nand UO_2278 (O_2278,N_24616,N_24104);
or UO_2279 (O_2279,N_24752,N_24729);
nand UO_2280 (O_2280,N_24050,N_24008);
and UO_2281 (O_2281,N_24768,N_24777);
nand UO_2282 (O_2282,N_24729,N_24004);
or UO_2283 (O_2283,N_24115,N_24300);
or UO_2284 (O_2284,N_24133,N_24894);
and UO_2285 (O_2285,N_24630,N_24522);
nor UO_2286 (O_2286,N_24017,N_24329);
xnor UO_2287 (O_2287,N_24296,N_24272);
and UO_2288 (O_2288,N_24505,N_24957);
or UO_2289 (O_2289,N_24057,N_24454);
and UO_2290 (O_2290,N_24037,N_24204);
or UO_2291 (O_2291,N_24433,N_24351);
or UO_2292 (O_2292,N_24779,N_24654);
or UO_2293 (O_2293,N_24172,N_24024);
or UO_2294 (O_2294,N_24385,N_24808);
and UO_2295 (O_2295,N_24011,N_24669);
or UO_2296 (O_2296,N_24412,N_24806);
nor UO_2297 (O_2297,N_24193,N_24984);
nor UO_2298 (O_2298,N_24575,N_24616);
or UO_2299 (O_2299,N_24674,N_24573);
xor UO_2300 (O_2300,N_24766,N_24407);
xnor UO_2301 (O_2301,N_24131,N_24930);
or UO_2302 (O_2302,N_24980,N_24391);
nor UO_2303 (O_2303,N_24249,N_24916);
xnor UO_2304 (O_2304,N_24816,N_24026);
nor UO_2305 (O_2305,N_24371,N_24023);
and UO_2306 (O_2306,N_24915,N_24885);
nand UO_2307 (O_2307,N_24441,N_24949);
xnor UO_2308 (O_2308,N_24121,N_24522);
nor UO_2309 (O_2309,N_24263,N_24454);
xnor UO_2310 (O_2310,N_24223,N_24821);
and UO_2311 (O_2311,N_24843,N_24099);
xnor UO_2312 (O_2312,N_24266,N_24027);
nand UO_2313 (O_2313,N_24097,N_24579);
or UO_2314 (O_2314,N_24852,N_24802);
nor UO_2315 (O_2315,N_24515,N_24010);
and UO_2316 (O_2316,N_24789,N_24332);
nor UO_2317 (O_2317,N_24206,N_24041);
nor UO_2318 (O_2318,N_24622,N_24247);
xnor UO_2319 (O_2319,N_24602,N_24699);
xor UO_2320 (O_2320,N_24146,N_24562);
or UO_2321 (O_2321,N_24295,N_24929);
xnor UO_2322 (O_2322,N_24148,N_24043);
nor UO_2323 (O_2323,N_24681,N_24170);
nor UO_2324 (O_2324,N_24410,N_24652);
xor UO_2325 (O_2325,N_24690,N_24463);
nand UO_2326 (O_2326,N_24684,N_24896);
xor UO_2327 (O_2327,N_24628,N_24760);
and UO_2328 (O_2328,N_24265,N_24601);
and UO_2329 (O_2329,N_24559,N_24789);
and UO_2330 (O_2330,N_24691,N_24938);
and UO_2331 (O_2331,N_24300,N_24274);
xor UO_2332 (O_2332,N_24771,N_24478);
and UO_2333 (O_2333,N_24909,N_24494);
nand UO_2334 (O_2334,N_24856,N_24826);
nand UO_2335 (O_2335,N_24831,N_24951);
or UO_2336 (O_2336,N_24592,N_24540);
or UO_2337 (O_2337,N_24290,N_24133);
xor UO_2338 (O_2338,N_24125,N_24232);
nand UO_2339 (O_2339,N_24257,N_24484);
nand UO_2340 (O_2340,N_24661,N_24032);
nor UO_2341 (O_2341,N_24935,N_24967);
or UO_2342 (O_2342,N_24934,N_24442);
nor UO_2343 (O_2343,N_24225,N_24090);
or UO_2344 (O_2344,N_24437,N_24930);
xnor UO_2345 (O_2345,N_24463,N_24803);
or UO_2346 (O_2346,N_24714,N_24201);
xor UO_2347 (O_2347,N_24052,N_24410);
xor UO_2348 (O_2348,N_24941,N_24020);
nor UO_2349 (O_2349,N_24183,N_24609);
xnor UO_2350 (O_2350,N_24038,N_24296);
nor UO_2351 (O_2351,N_24520,N_24432);
and UO_2352 (O_2352,N_24164,N_24172);
nor UO_2353 (O_2353,N_24098,N_24540);
nor UO_2354 (O_2354,N_24021,N_24348);
nor UO_2355 (O_2355,N_24373,N_24513);
nor UO_2356 (O_2356,N_24008,N_24961);
xor UO_2357 (O_2357,N_24712,N_24337);
and UO_2358 (O_2358,N_24601,N_24014);
xnor UO_2359 (O_2359,N_24993,N_24803);
and UO_2360 (O_2360,N_24845,N_24370);
nand UO_2361 (O_2361,N_24940,N_24083);
xnor UO_2362 (O_2362,N_24534,N_24535);
xor UO_2363 (O_2363,N_24265,N_24819);
xor UO_2364 (O_2364,N_24054,N_24679);
or UO_2365 (O_2365,N_24727,N_24485);
nor UO_2366 (O_2366,N_24436,N_24364);
nand UO_2367 (O_2367,N_24277,N_24252);
nor UO_2368 (O_2368,N_24384,N_24137);
or UO_2369 (O_2369,N_24661,N_24770);
xor UO_2370 (O_2370,N_24791,N_24197);
xnor UO_2371 (O_2371,N_24038,N_24500);
and UO_2372 (O_2372,N_24588,N_24713);
xnor UO_2373 (O_2373,N_24832,N_24907);
nor UO_2374 (O_2374,N_24523,N_24335);
and UO_2375 (O_2375,N_24485,N_24498);
nand UO_2376 (O_2376,N_24430,N_24889);
and UO_2377 (O_2377,N_24514,N_24797);
nor UO_2378 (O_2378,N_24341,N_24842);
nor UO_2379 (O_2379,N_24129,N_24861);
nor UO_2380 (O_2380,N_24794,N_24856);
and UO_2381 (O_2381,N_24666,N_24321);
and UO_2382 (O_2382,N_24331,N_24884);
nor UO_2383 (O_2383,N_24863,N_24316);
nand UO_2384 (O_2384,N_24847,N_24162);
xnor UO_2385 (O_2385,N_24108,N_24088);
and UO_2386 (O_2386,N_24876,N_24208);
and UO_2387 (O_2387,N_24860,N_24681);
nand UO_2388 (O_2388,N_24226,N_24103);
or UO_2389 (O_2389,N_24007,N_24633);
nor UO_2390 (O_2390,N_24180,N_24104);
nor UO_2391 (O_2391,N_24760,N_24224);
and UO_2392 (O_2392,N_24546,N_24104);
and UO_2393 (O_2393,N_24872,N_24067);
or UO_2394 (O_2394,N_24858,N_24779);
nor UO_2395 (O_2395,N_24802,N_24895);
and UO_2396 (O_2396,N_24589,N_24764);
xor UO_2397 (O_2397,N_24350,N_24467);
nor UO_2398 (O_2398,N_24337,N_24719);
nor UO_2399 (O_2399,N_24055,N_24473);
and UO_2400 (O_2400,N_24845,N_24225);
and UO_2401 (O_2401,N_24820,N_24121);
xnor UO_2402 (O_2402,N_24213,N_24612);
and UO_2403 (O_2403,N_24972,N_24355);
xnor UO_2404 (O_2404,N_24229,N_24154);
nor UO_2405 (O_2405,N_24959,N_24081);
xnor UO_2406 (O_2406,N_24827,N_24321);
nor UO_2407 (O_2407,N_24249,N_24311);
and UO_2408 (O_2408,N_24562,N_24895);
nand UO_2409 (O_2409,N_24981,N_24598);
nor UO_2410 (O_2410,N_24267,N_24226);
xnor UO_2411 (O_2411,N_24539,N_24793);
nand UO_2412 (O_2412,N_24969,N_24138);
nor UO_2413 (O_2413,N_24000,N_24833);
xnor UO_2414 (O_2414,N_24355,N_24885);
or UO_2415 (O_2415,N_24633,N_24856);
and UO_2416 (O_2416,N_24103,N_24596);
xor UO_2417 (O_2417,N_24621,N_24126);
xor UO_2418 (O_2418,N_24599,N_24618);
nand UO_2419 (O_2419,N_24638,N_24293);
or UO_2420 (O_2420,N_24897,N_24898);
xnor UO_2421 (O_2421,N_24448,N_24591);
xnor UO_2422 (O_2422,N_24064,N_24083);
and UO_2423 (O_2423,N_24655,N_24654);
or UO_2424 (O_2424,N_24679,N_24785);
nand UO_2425 (O_2425,N_24785,N_24882);
or UO_2426 (O_2426,N_24967,N_24718);
or UO_2427 (O_2427,N_24996,N_24228);
nor UO_2428 (O_2428,N_24285,N_24595);
or UO_2429 (O_2429,N_24590,N_24535);
nor UO_2430 (O_2430,N_24166,N_24777);
and UO_2431 (O_2431,N_24718,N_24366);
nand UO_2432 (O_2432,N_24943,N_24047);
xnor UO_2433 (O_2433,N_24701,N_24420);
nor UO_2434 (O_2434,N_24719,N_24501);
nor UO_2435 (O_2435,N_24301,N_24073);
and UO_2436 (O_2436,N_24111,N_24476);
nor UO_2437 (O_2437,N_24168,N_24261);
nor UO_2438 (O_2438,N_24825,N_24930);
or UO_2439 (O_2439,N_24549,N_24901);
and UO_2440 (O_2440,N_24411,N_24478);
nor UO_2441 (O_2441,N_24662,N_24544);
xor UO_2442 (O_2442,N_24748,N_24991);
nand UO_2443 (O_2443,N_24138,N_24026);
nor UO_2444 (O_2444,N_24695,N_24146);
nand UO_2445 (O_2445,N_24296,N_24013);
nor UO_2446 (O_2446,N_24517,N_24607);
nand UO_2447 (O_2447,N_24459,N_24115);
or UO_2448 (O_2448,N_24667,N_24510);
or UO_2449 (O_2449,N_24184,N_24484);
and UO_2450 (O_2450,N_24343,N_24479);
nand UO_2451 (O_2451,N_24702,N_24295);
or UO_2452 (O_2452,N_24398,N_24148);
xor UO_2453 (O_2453,N_24286,N_24828);
and UO_2454 (O_2454,N_24370,N_24291);
nor UO_2455 (O_2455,N_24231,N_24463);
xor UO_2456 (O_2456,N_24918,N_24257);
nor UO_2457 (O_2457,N_24846,N_24812);
nand UO_2458 (O_2458,N_24244,N_24618);
or UO_2459 (O_2459,N_24345,N_24827);
and UO_2460 (O_2460,N_24798,N_24608);
nand UO_2461 (O_2461,N_24012,N_24985);
nor UO_2462 (O_2462,N_24906,N_24038);
or UO_2463 (O_2463,N_24383,N_24752);
or UO_2464 (O_2464,N_24176,N_24236);
or UO_2465 (O_2465,N_24411,N_24259);
nor UO_2466 (O_2466,N_24547,N_24338);
or UO_2467 (O_2467,N_24796,N_24010);
nand UO_2468 (O_2468,N_24682,N_24889);
and UO_2469 (O_2469,N_24542,N_24384);
and UO_2470 (O_2470,N_24861,N_24933);
nor UO_2471 (O_2471,N_24365,N_24332);
nor UO_2472 (O_2472,N_24460,N_24635);
xnor UO_2473 (O_2473,N_24401,N_24580);
nor UO_2474 (O_2474,N_24710,N_24965);
xnor UO_2475 (O_2475,N_24515,N_24226);
nor UO_2476 (O_2476,N_24623,N_24415);
nand UO_2477 (O_2477,N_24932,N_24250);
xnor UO_2478 (O_2478,N_24538,N_24161);
xor UO_2479 (O_2479,N_24989,N_24614);
and UO_2480 (O_2480,N_24250,N_24519);
and UO_2481 (O_2481,N_24363,N_24558);
or UO_2482 (O_2482,N_24027,N_24471);
nand UO_2483 (O_2483,N_24847,N_24687);
or UO_2484 (O_2484,N_24339,N_24036);
nor UO_2485 (O_2485,N_24419,N_24538);
xor UO_2486 (O_2486,N_24980,N_24990);
and UO_2487 (O_2487,N_24940,N_24200);
xnor UO_2488 (O_2488,N_24189,N_24558);
or UO_2489 (O_2489,N_24684,N_24631);
or UO_2490 (O_2490,N_24107,N_24773);
and UO_2491 (O_2491,N_24038,N_24674);
xnor UO_2492 (O_2492,N_24292,N_24109);
nand UO_2493 (O_2493,N_24760,N_24262);
and UO_2494 (O_2494,N_24205,N_24672);
nand UO_2495 (O_2495,N_24904,N_24889);
nor UO_2496 (O_2496,N_24054,N_24490);
xor UO_2497 (O_2497,N_24033,N_24917);
xnor UO_2498 (O_2498,N_24435,N_24601);
nand UO_2499 (O_2499,N_24489,N_24411);
xnor UO_2500 (O_2500,N_24862,N_24660);
or UO_2501 (O_2501,N_24548,N_24199);
and UO_2502 (O_2502,N_24126,N_24096);
xor UO_2503 (O_2503,N_24938,N_24792);
xor UO_2504 (O_2504,N_24037,N_24933);
nor UO_2505 (O_2505,N_24050,N_24207);
xor UO_2506 (O_2506,N_24523,N_24937);
nand UO_2507 (O_2507,N_24403,N_24299);
nor UO_2508 (O_2508,N_24037,N_24995);
and UO_2509 (O_2509,N_24430,N_24154);
and UO_2510 (O_2510,N_24358,N_24162);
or UO_2511 (O_2511,N_24599,N_24453);
and UO_2512 (O_2512,N_24630,N_24484);
or UO_2513 (O_2513,N_24018,N_24331);
xor UO_2514 (O_2514,N_24337,N_24682);
nor UO_2515 (O_2515,N_24262,N_24585);
or UO_2516 (O_2516,N_24596,N_24042);
or UO_2517 (O_2517,N_24240,N_24165);
nor UO_2518 (O_2518,N_24109,N_24295);
or UO_2519 (O_2519,N_24210,N_24902);
xnor UO_2520 (O_2520,N_24001,N_24925);
and UO_2521 (O_2521,N_24329,N_24063);
or UO_2522 (O_2522,N_24321,N_24912);
nor UO_2523 (O_2523,N_24171,N_24224);
xnor UO_2524 (O_2524,N_24391,N_24866);
and UO_2525 (O_2525,N_24950,N_24636);
and UO_2526 (O_2526,N_24870,N_24874);
and UO_2527 (O_2527,N_24252,N_24513);
nand UO_2528 (O_2528,N_24648,N_24364);
and UO_2529 (O_2529,N_24839,N_24465);
nor UO_2530 (O_2530,N_24102,N_24281);
nor UO_2531 (O_2531,N_24080,N_24054);
xnor UO_2532 (O_2532,N_24036,N_24264);
nor UO_2533 (O_2533,N_24274,N_24094);
xnor UO_2534 (O_2534,N_24727,N_24467);
nand UO_2535 (O_2535,N_24118,N_24105);
nand UO_2536 (O_2536,N_24914,N_24545);
nand UO_2537 (O_2537,N_24452,N_24648);
nand UO_2538 (O_2538,N_24797,N_24382);
or UO_2539 (O_2539,N_24345,N_24327);
or UO_2540 (O_2540,N_24336,N_24397);
or UO_2541 (O_2541,N_24307,N_24392);
xnor UO_2542 (O_2542,N_24116,N_24659);
xor UO_2543 (O_2543,N_24131,N_24102);
xnor UO_2544 (O_2544,N_24692,N_24673);
and UO_2545 (O_2545,N_24951,N_24185);
xor UO_2546 (O_2546,N_24581,N_24521);
and UO_2547 (O_2547,N_24491,N_24275);
and UO_2548 (O_2548,N_24778,N_24392);
xor UO_2549 (O_2549,N_24622,N_24356);
xnor UO_2550 (O_2550,N_24185,N_24585);
nand UO_2551 (O_2551,N_24979,N_24777);
and UO_2552 (O_2552,N_24356,N_24710);
nor UO_2553 (O_2553,N_24300,N_24176);
and UO_2554 (O_2554,N_24262,N_24209);
and UO_2555 (O_2555,N_24809,N_24050);
or UO_2556 (O_2556,N_24877,N_24718);
nor UO_2557 (O_2557,N_24663,N_24465);
xnor UO_2558 (O_2558,N_24645,N_24585);
or UO_2559 (O_2559,N_24798,N_24451);
and UO_2560 (O_2560,N_24396,N_24315);
xnor UO_2561 (O_2561,N_24861,N_24682);
and UO_2562 (O_2562,N_24347,N_24232);
or UO_2563 (O_2563,N_24168,N_24490);
nand UO_2564 (O_2564,N_24553,N_24549);
xor UO_2565 (O_2565,N_24109,N_24480);
xor UO_2566 (O_2566,N_24101,N_24545);
or UO_2567 (O_2567,N_24702,N_24476);
nand UO_2568 (O_2568,N_24133,N_24235);
nand UO_2569 (O_2569,N_24010,N_24265);
and UO_2570 (O_2570,N_24321,N_24385);
xor UO_2571 (O_2571,N_24008,N_24085);
or UO_2572 (O_2572,N_24509,N_24415);
nor UO_2573 (O_2573,N_24102,N_24862);
and UO_2574 (O_2574,N_24827,N_24571);
or UO_2575 (O_2575,N_24222,N_24546);
nand UO_2576 (O_2576,N_24306,N_24366);
and UO_2577 (O_2577,N_24917,N_24265);
or UO_2578 (O_2578,N_24016,N_24322);
and UO_2579 (O_2579,N_24629,N_24440);
xor UO_2580 (O_2580,N_24989,N_24656);
and UO_2581 (O_2581,N_24391,N_24928);
or UO_2582 (O_2582,N_24451,N_24960);
and UO_2583 (O_2583,N_24388,N_24688);
and UO_2584 (O_2584,N_24910,N_24379);
or UO_2585 (O_2585,N_24916,N_24049);
xnor UO_2586 (O_2586,N_24911,N_24298);
xor UO_2587 (O_2587,N_24587,N_24537);
and UO_2588 (O_2588,N_24569,N_24126);
and UO_2589 (O_2589,N_24980,N_24958);
nor UO_2590 (O_2590,N_24678,N_24372);
nand UO_2591 (O_2591,N_24102,N_24267);
and UO_2592 (O_2592,N_24312,N_24386);
nor UO_2593 (O_2593,N_24289,N_24578);
or UO_2594 (O_2594,N_24425,N_24512);
nand UO_2595 (O_2595,N_24576,N_24539);
nor UO_2596 (O_2596,N_24839,N_24037);
nand UO_2597 (O_2597,N_24246,N_24393);
nand UO_2598 (O_2598,N_24278,N_24121);
nor UO_2599 (O_2599,N_24811,N_24601);
nor UO_2600 (O_2600,N_24077,N_24558);
xor UO_2601 (O_2601,N_24553,N_24131);
or UO_2602 (O_2602,N_24179,N_24070);
or UO_2603 (O_2603,N_24761,N_24695);
and UO_2604 (O_2604,N_24310,N_24766);
and UO_2605 (O_2605,N_24723,N_24831);
nand UO_2606 (O_2606,N_24703,N_24308);
or UO_2607 (O_2607,N_24286,N_24013);
xnor UO_2608 (O_2608,N_24624,N_24939);
xor UO_2609 (O_2609,N_24310,N_24184);
and UO_2610 (O_2610,N_24180,N_24730);
and UO_2611 (O_2611,N_24765,N_24349);
and UO_2612 (O_2612,N_24916,N_24212);
xor UO_2613 (O_2613,N_24759,N_24050);
and UO_2614 (O_2614,N_24267,N_24481);
nand UO_2615 (O_2615,N_24658,N_24190);
xnor UO_2616 (O_2616,N_24563,N_24947);
and UO_2617 (O_2617,N_24724,N_24008);
xor UO_2618 (O_2618,N_24315,N_24164);
and UO_2619 (O_2619,N_24979,N_24392);
xor UO_2620 (O_2620,N_24840,N_24588);
or UO_2621 (O_2621,N_24043,N_24394);
or UO_2622 (O_2622,N_24180,N_24255);
nor UO_2623 (O_2623,N_24971,N_24759);
or UO_2624 (O_2624,N_24599,N_24088);
xor UO_2625 (O_2625,N_24058,N_24728);
or UO_2626 (O_2626,N_24988,N_24212);
xor UO_2627 (O_2627,N_24247,N_24818);
nor UO_2628 (O_2628,N_24476,N_24590);
and UO_2629 (O_2629,N_24043,N_24633);
nor UO_2630 (O_2630,N_24915,N_24752);
xnor UO_2631 (O_2631,N_24097,N_24181);
xor UO_2632 (O_2632,N_24283,N_24640);
nand UO_2633 (O_2633,N_24186,N_24801);
nand UO_2634 (O_2634,N_24210,N_24877);
nand UO_2635 (O_2635,N_24284,N_24652);
nor UO_2636 (O_2636,N_24075,N_24154);
nand UO_2637 (O_2637,N_24432,N_24717);
nor UO_2638 (O_2638,N_24070,N_24512);
nor UO_2639 (O_2639,N_24066,N_24919);
nand UO_2640 (O_2640,N_24951,N_24900);
or UO_2641 (O_2641,N_24045,N_24400);
nand UO_2642 (O_2642,N_24170,N_24349);
nor UO_2643 (O_2643,N_24150,N_24637);
xnor UO_2644 (O_2644,N_24224,N_24587);
nand UO_2645 (O_2645,N_24523,N_24386);
or UO_2646 (O_2646,N_24705,N_24762);
nor UO_2647 (O_2647,N_24351,N_24042);
and UO_2648 (O_2648,N_24100,N_24039);
xor UO_2649 (O_2649,N_24106,N_24912);
and UO_2650 (O_2650,N_24929,N_24731);
nor UO_2651 (O_2651,N_24119,N_24245);
nor UO_2652 (O_2652,N_24757,N_24080);
nand UO_2653 (O_2653,N_24619,N_24615);
or UO_2654 (O_2654,N_24215,N_24559);
nor UO_2655 (O_2655,N_24304,N_24694);
or UO_2656 (O_2656,N_24118,N_24225);
nor UO_2657 (O_2657,N_24208,N_24022);
nor UO_2658 (O_2658,N_24366,N_24470);
nor UO_2659 (O_2659,N_24786,N_24635);
nand UO_2660 (O_2660,N_24788,N_24940);
nor UO_2661 (O_2661,N_24393,N_24226);
nand UO_2662 (O_2662,N_24680,N_24882);
xnor UO_2663 (O_2663,N_24638,N_24320);
nand UO_2664 (O_2664,N_24725,N_24402);
nor UO_2665 (O_2665,N_24431,N_24763);
nand UO_2666 (O_2666,N_24060,N_24287);
nor UO_2667 (O_2667,N_24879,N_24401);
nor UO_2668 (O_2668,N_24331,N_24563);
nand UO_2669 (O_2669,N_24197,N_24058);
nand UO_2670 (O_2670,N_24324,N_24718);
nor UO_2671 (O_2671,N_24476,N_24915);
and UO_2672 (O_2672,N_24209,N_24633);
xnor UO_2673 (O_2673,N_24384,N_24590);
nand UO_2674 (O_2674,N_24959,N_24219);
xor UO_2675 (O_2675,N_24774,N_24562);
nor UO_2676 (O_2676,N_24395,N_24392);
nor UO_2677 (O_2677,N_24940,N_24970);
and UO_2678 (O_2678,N_24199,N_24922);
or UO_2679 (O_2679,N_24957,N_24254);
nor UO_2680 (O_2680,N_24829,N_24048);
nand UO_2681 (O_2681,N_24754,N_24672);
xnor UO_2682 (O_2682,N_24331,N_24739);
or UO_2683 (O_2683,N_24938,N_24386);
or UO_2684 (O_2684,N_24007,N_24974);
and UO_2685 (O_2685,N_24642,N_24917);
or UO_2686 (O_2686,N_24394,N_24034);
and UO_2687 (O_2687,N_24080,N_24322);
and UO_2688 (O_2688,N_24644,N_24355);
and UO_2689 (O_2689,N_24875,N_24015);
nand UO_2690 (O_2690,N_24562,N_24712);
and UO_2691 (O_2691,N_24710,N_24038);
xnor UO_2692 (O_2692,N_24481,N_24136);
xnor UO_2693 (O_2693,N_24367,N_24165);
nor UO_2694 (O_2694,N_24279,N_24824);
and UO_2695 (O_2695,N_24286,N_24035);
nand UO_2696 (O_2696,N_24614,N_24780);
and UO_2697 (O_2697,N_24840,N_24784);
nand UO_2698 (O_2698,N_24704,N_24326);
nor UO_2699 (O_2699,N_24738,N_24917);
xnor UO_2700 (O_2700,N_24107,N_24463);
and UO_2701 (O_2701,N_24734,N_24777);
and UO_2702 (O_2702,N_24838,N_24772);
xnor UO_2703 (O_2703,N_24877,N_24875);
nand UO_2704 (O_2704,N_24748,N_24979);
and UO_2705 (O_2705,N_24454,N_24321);
nand UO_2706 (O_2706,N_24780,N_24115);
or UO_2707 (O_2707,N_24557,N_24126);
nand UO_2708 (O_2708,N_24119,N_24054);
nand UO_2709 (O_2709,N_24386,N_24623);
and UO_2710 (O_2710,N_24261,N_24472);
nand UO_2711 (O_2711,N_24618,N_24823);
nand UO_2712 (O_2712,N_24805,N_24784);
and UO_2713 (O_2713,N_24315,N_24157);
and UO_2714 (O_2714,N_24993,N_24162);
or UO_2715 (O_2715,N_24227,N_24260);
and UO_2716 (O_2716,N_24898,N_24299);
nand UO_2717 (O_2717,N_24867,N_24631);
nand UO_2718 (O_2718,N_24262,N_24296);
xnor UO_2719 (O_2719,N_24666,N_24998);
nand UO_2720 (O_2720,N_24411,N_24346);
and UO_2721 (O_2721,N_24797,N_24314);
nor UO_2722 (O_2722,N_24782,N_24966);
and UO_2723 (O_2723,N_24662,N_24540);
nor UO_2724 (O_2724,N_24464,N_24267);
nand UO_2725 (O_2725,N_24498,N_24872);
nand UO_2726 (O_2726,N_24943,N_24883);
nor UO_2727 (O_2727,N_24658,N_24337);
and UO_2728 (O_2728,N_24640,N_24903);
and UO_2729 (O_2729,N_24644,N_24657);
or UO_2730 (O_2730,N_24741,N_24627);
or UO_2731 (O_2731,N_24469,N_24905);
nand UO_2732 (O_2732,N_24121,N_24011);
and UO_2733 (O_2733,N_24409,N_24268);
and UO_2734 (O_2734,N_24327,N_24469);
nor UO_2735 (O_2735,N_24279,N_24104);
nand UO_2736 (O_2736,N_24406,N_24554);
xor UO_2737 (O_2737,N_24955,N_24667);
nor UO_2738 (O_2738,N_24205,N_24017);
xnor UO_2739 (O_2739,N_24029,N_24512);
xnor UO_2740 (O_2740,N_24172,N_24039);
nand UO_2741 (O_2741,N_24424,N_24117);
nor UO_2742 (O_2742,N_24879,N_24433);
or UO_2743 (O_2743,N_24336,N_24681);
or UO_2744 (O_2744,N_24389,N_24581);
and UO_2745 (O_2745,N_24080,N_24352);
or UO_2746 (O_2746,N_24190,N_24587);
or UO_2747 (O_2747,N_24518,N_24124);
nor UO_2748 (O_2748,N_24212,N_24188);
and UO_2749 (O_2749,N_24014,N_24815);
and UO_2750 (O_2750,N_24930,N_24883);
nor UO_2751 (O_2751,N_24039,N_24772);
or UO_2752 (O_2752,N_24569,N_24360);
nand UO_2753 (O_2753,N_24163,N_24302);
nor UO_2754 (O_2754,N_24367,N_24213);
xnor UO_2755 (O_2755,N_24369,N_24958);
xnor UO_2756 (O_2756,N_24521,N_24094);
or UO_2757 (O_2757,N_24706,N_24804);
xor UO_2758 (O_2758,N_24941,N_24821);
and UO_2759 (O_2759,N_24488,N_24309);
nor UO_2760 (O_2760,N_24284,N_24033);
nor UO_2761 (O_2761,N_24125,N_24651);
and UO_2762 (O_2762,N_24544,N_24598);
or UO_2763 (O_2763,N_24444,N_24371);
and UO_2764 (O_2764,N_24999,N_24680);
and UO_2765 (O_2765,N_24858,N_24600);
or UO_2766 (O_2766,N_24933,N_24251);
nand UO_2767 (O_2767,N_24318,N_24145);
xor UO_2768 (O_2768,N_24439,N_24938);
and UO_2769 (O_2769,N_24289,N_24947);
nor UO_2770 (O_2770,N_24750,N_24988);
xnor UO_2771 (O_2771,N_24905,N_24894);
or UO_2772 (O_2772,N_24754,N_24930);
or UO_2773 (O_2773,N_24431,N_24662);
nand UO_2774 (O_2774,N_24870,N_24325);
and UO_2775 (O_2775,N_24983,N_24534);
nor UO_2776 (O_2776,N_24288,N_24788);
xor UO_2777 (O_2777,N_24556,N_24954);
xor UO_2778 (O_2778,N_24096,N_24412);
nor UO_2779 (O_2779,N_24329,N_24642);
and UO_2780 (O_2780,N_24184,N_24289);
nor UO_2781 (O_2781,N_24070,N_24909);
nor UO_2782 (O_2782,N_24794,N_24668);
xor UO_2783 (O_2783,N_24585,N_24934);
or UO_2784 (O_2784,N_24580,N_24578);
or UO_2785 (O_2785,N_24900,N_24571);
xnor UO_2786 (O_2786,N_24979,N_24822);
xor UO_2787 (O_2787,N_24875,N_24506);
nand UO_2788 (O_2788,N_24162,N_24015);
and UO_2789 (O_2789,N_24767,N_24777);
or UO_2790 (O_2790,N_24651,N_24661);
or UO_2791 (O_2791,N_24575,N_24373);
nand UO_2792 (O_2792,N_24853,N_24113);
xnor UO_2793 (O_2793,N_24385,N_24217);
nor UO_2794 (O_2794,N_24072,N_24802);
or UO_2795 (O_2795,N_24794,N_24882);
nor UO_2796 (O_2796,N_24469,N_24191);
or UO_2797 (O_2797,N_24384,N_24517);
nor UO_2798 (O_2798,N_24085,N_24350);
nor UO_2799 (O_2799,N_24323,N_24533);
nand UO_2800 (O_2800,N_24068,N_24069);
nand UO_2801 (O_2801,N_24352,N_24686);
xnor UO_2802 (O_2802,N_24176,N_24210);
nand UO_2803 (O_2803,N_24052,N_24810);
nand UO_2804 (O_2804,N_24196,N_24465);
nor UO_2805 (O_2805,N_24477,N_24869);
and UO_2806 (O_2806,N_24358,N_24912);
xor UO_2807 (O_2807,N_24178,N_24156);
and UO_2808 (O_2808,N_24134,N_24088);
or UO_2809 (O_2809,N_24620,N_24704);
nor UO_2810 (O_2810,N_24297,N_24655);
nand UO_2811 (O_2811,N_24926,N_24907);
nand UO_2812 (O_2812,N_24122,N_24223);
and UO_2813 (O_2813,N_24942,N_24198);
nand UO_2814 (O_2814,N_24590,N_24975);
xnor UO_2815 (O_2815,N_24528,N_24833);
xnor UO_2816 (O_2816,N_24903,N_24262);
nor UO_2817 (O_2817,N_24562,N_24748);
nand UO_2818 (O_2818,N_24247,N_24235);
nand UO_2819 (O_2819,N_24535,N_24157);
nor UO_2820 (O_2820,N_24998,N_24214);
and UO_2821 (O_2821,N_24262,N_24095);
xnor UO_2822 (O_2822,N_24413,N_24494);
nor UO_2823 (O_2823,N_24657,N_24098);
xor UO_2824 (O_2824,N_24026,N_24000);
xnor UO_2825 (O_2825,N_24524,N_24215);
nor UO_2826 (O_2826,N_24980,N_24205);
xor UO_2827 (O_2827,N_24245,N_24869);
and UO_2828 (O_2828,N_24481,N_24744);
and UO_2829 (O_2829,N_24296,N_24999);
xor UO_2830 (O_2830,N_24849,N_24101);
nand UO_2831 (O_2831,N_24074,N_24682);
and UO_2832 (O_2832,N_24446,N_24705);
nand UO_2833 (O_2833,N_24091,N_24451);
or UO_2834 (O_2834,N_24405,N_24369);
nor UO_2835 (O_2835,N_24913,N_24531);
xor UO_2836 (O_2836,N_24275,N_24064);
nor UO_2837 (O_2837,N_24741,N_24797);
or UO_2838 (O_2838,N_24648,N_24451);
nor UO_2839 (O_2839,N_24286,N_24992);
nor UO_2840 (O_2840,N_24884,N_24892);
and UO_2841 (O_2841,N_24708,N_24098);
nor UO_2842 (O_2842,N_24992,N_24745);
nand UO_2843 (O_2843,N_24571,N_24284);
or UO_2844 (O_2844,N_24150,N_24696);
xor UO_2845 (O_2845,N_24308,N_24505);
xor UO_2846 (O_2846,N_24668,N_24229);
and UO_2847 (O_2847,N_24303,N_24954);
and UO_2848 (O_2848,N_24019,N_24081);
and UO_2849 (O_2849,N_24252,N_24283);
nand UO_2850 (O_2850,N_24669,N_24000);
and UO_2851 (O_2851,N_24929,N_24485);
or UO_2852 (O_2852,N_24881,N_24764);
or UO_2853 (O_2853,N_24145,N_24495);
or UO_2854 (O_2854,N_24115,N_24747);
or UO_2855 (O_2855,N_24792,N_24946);
or UO_2856 (O_2856,N_24840,N_24679);
nor UO_2857 (O_2857,N_24802,N_24579);
nand UO_2858 (O_2858,N_24630,N_24141);
or UO_2859 (O_2859,N_24075,N_24332);
nand UO_2860 (O_2860,N_24007,N_24840);
xor UO_2861 (O_2861,N_24218,N_24560);
nand UO_2862 (O_2862,N_24782,N_24710);
nor UO_2863 (O_2863,N_24790,N_24711);
nor UO_2864 (O_2864,N_24502,N_24965);
and UO_2865 (O_2865,N_24678,N_24491);
and UO_2866 (O_2866,N_24159,N_24695);
nand UO_2867 (O_2867,N_24299,N_24979);
and UO_2868 (O_2868,N_24305,N_24715);
or UO_2869 (O_2869,N_24430,N_24885);
nand UO_2870 (O_2870,N_24552,N_24431);
or UO_2871 (O_2871,N_24683,N_24515);
or UO_2872 (O_2872,N_24851,N_24896);
xor UO_2873 (O_2873,N_24271,N_24737);
or UO_2874 (O_2874,N_24440,N_24458);
or UO_2875 (O_2875,N_24116,N_24461);
nand UO_2876 (O_2876,N_24169,N_24535);
nand UO_2877 (O_2877,N_24062,N_24534);
nor UO_2878 (O_2878,N_24884,N_24829);
xnor UO_2879 (O_2879,N_24719,N_24704);
xnor UO_2880 (O_2880,N_24412,N_24267);
nand UO_2881 (O_2881,N_24897,N_24966);
and UO_2882 (O_2882,N_24275,N_24405);
or UO_2883 (O_2883,N_24337,N_24362);
nand UO_2884 (O_2884,N_24212,N_24710);
xor UO_2885 (O_2885,N_24700,N_24432);
nor UO_2886 (O_2886,N_24855,N_24084);
xor UO_2887 (O_2887,N_24672,N_24327);
nand UO_2888 (O_2888,N_24186,N_24471);
nor UO_2889 (O_2889,N_24828,N_24581);
xnor UO_2890 (O_2890,N_24087,N_24596);
or UO_2891 (O_2891,N_24243,N_24467);
nor UO_2892 (O_2892,N_24983,N_24587);
nand UO_2893 (O_2893,N_24552,N_24033);
nand UO_2894 (O_2894,N_24033,N_24607);
xor UO_2895 (O_2895,N_24812,N_24698);
and UO_2896 (O_2896,N_24049,N_24021);
nand UO_2897 (O_2897,N_24361,N_24568);
nor UO_2898 (O_2898,N_24109,N_24912);
nand UO_2899 (O_2899,N_24154,N_24541);
or UO_2900 (O_2900,N_24307,N_24134);
nor UO_2901 (O_2901,N_24418,N_24386);
and UO_2902 (O_2902,N_24704,N_24063);
nor UO_2903 (O_2903,N_24769,N_24467);
or UO_2904 (O_2904,N_24236,N_24352);
or UO_2905 (O_2905,N_24629,N_24745);
nor UO_2906 (O_2906,N_24797,N_24670);
xor UO_2907 (O_2907,N_24029,N_24868);
nand UO_2908 (O_2908,N_24636,N_24273);
or UO_2909 (O_2909,N_24319,N_24083);
nand UO_2910 (O_2910,N_24737,N_24695);
nand UO_2911 (O_2911,N_24799,N_24452);
and UO_2912 (O_2912,N_24746,N_24386);
or UO_2913 (O_2913,N_24002,N_24665);
or UO_2914 (O_2914,N_24783,N_24163);
xnor UO_2915 (O_2915,N_24118,N_24095);
or UO_2916 (O_2916,N_24615,N_24506);
nand UO_2917 (O_2917,N_24321,N_24971);
nand UO_2918 (O_2918,N_24949,N_24173);
and UO_2919 (O_2919,N_24028,N_24456);
nand UO_2920 (O_2920,N_24152,N_24055);
nor UO_2921 (O_2921,N_24124,N_24999);
xnor UO_2922 (O_2922,N_24113,N_24253);
nand UO_2923 (O_2923,N_24572,N_24827);
nand UO_2924 (O_2924,N_24685,N_24942);
and UO_2925 (O_2925,N_24600,N_24258);
xnor UO_2926 (O_2926,N_24905,N_24599);
xor UO_2927 (O_2927,N_24612,N_24277);
and UO_2928 (O_2928,N_24757,N_24632);
xnor UO_2929 (O_2929,N_24286,N_24621);
nor UO_2930 (O_2930,N_24861,N_24904);
or UO_2931 (O_2931,N_24683,N_24041);
nand UO_2932 (O_2932,N_24588,N_24152);
nand UO_2933 (O_2933,N_24753,N_24381);
and UO_2934 (O_2934,N_24907,N_24968);
or UO_2935 (O_2935,N_24485,N_24153);
nor UO_2936 (O_2936,N_24053,N_24287);
nor UO_2937 (O_2937,N_24475,N_24589);
nand UO_2938 (O_2938,N_24100,N_24308);
nor UO_2939 (O_2939,N_24546,N_24490);
and UO_2940 (O_2940,N_24694,N_24000);
nor UO_2941 (O_2941,N_24517,N_24113);
nor UO_2942 (O_2942,N_24813,N_24819);
nor UO_2943 (O_2943,N_24040,N_24426);
nor UO_2944 (O_2944,N_24096,N_24233);
or UO_2945 (O_2945,N_24788,N_24508);
nor UO_2946 (O_2946,N_24651,N_24276);
nor UO_2947 (O_2947,N_24888,N_24046);
xnor UO_2948 (O_2948,N_24581,N_24158);
and UO_2949 (O_2949,N_24185,N_24114);
nand UO_2950 (O_2950,N_24774,N_24099);
xor UO_2951 (O_2951,N_24172,N_24401);
and UO_2952 (O_2952,N_24390,N_24541);
or UO_2953 (O_2953,N_24492,N_24227);
and UO_2954 (O_2954,N_24186,N_24948);
xor UO_2955 (O_2955,N_24556,N_24749);
or UO_2956 (O_2956,N_24223,N_24843);
nor UO_2957 (O_2957,N_24161,N_24987);
xor UO_2958 (O_2958,N_24846,N_24133);
xor UO_2959 (O_2959,N_24109,N_24048);
or UO_2960 (O_2960,N_24760,N_24569);
xnor UO_2961 (O_2961,N_24882,N_24975);
xor UO_2962 (O_2962,N_24279,N_24775);
nand UO_2963 (O_2963,N_24326,N_24924);
nand UO_2964 (O_2964,N_24985,N_24541);
xor UO_2965 (O_2965,N_24177,N_24420);
nand UO_2966 (O_2966,N_24329,N_24944);
nor UO_2967 (O_2967,N_24578,N_24677);
or UO_2968 (O_2968,N_24048,N_24969);
nor UO_2969 (O_2969,N_24162,N_24031);
xnor UO_2970 (O_2970,N_24433,N_24919);
or UO_2971 (O_2971,N_24702,N_24066);
xor UO_2972 (O_2972,N_24452,N_24217);
and UO_2973 (O_2973,N_24197,N_24556);
and UO_2974 (O_2974,N_24295,N_24655);
xnor UO_2975 (O_2975,N_24390,N_24018);
xor UO_2976 (O_2976,N_24885,N_24424);
and UO_2977 (O_2977,N_24702,N_24535);
or UO_2978 (O_2978,N_24094,N_24589);
and UO_2979 (O_2979,N_24178,N_24848);
or UO_2980 (O_2980,N_24602,N_24118);
and UO_2981 (O_2981,N_24166,N_24434);
and UO_2982 (O_2982,N_24686,N_24032);
and UO_2983 (O_2983,N_24975,N_24679);
or UO_2984 (O_2984,N_24243,N_24123);
nand UO_2985 (O_2985,N_24887,N_24116);
xnor UO_2986 (O_2986,N_24102,N_24731);
nor UO_2987 (O_2987,N_24856,N_24418);
or UO_2988 (O_2988,N_24490,N_24617);
nor UO_2989 (O_2989,N_24306,N_24132);
nor UO_2990 (O_2990,N_24347,N_24358);
nor UO_2991 (O_2991,N_24829,N_24176);
nor UO_2992 (O_2992,N_24133,N_24587);
xnor UO_2993 (O_2993,N_24558,N_24655);
or UO_2994 (O_2994,N_24599,N_24564);
and UO_2995 (O_2995,N_24442,N_24102);
nor UO_2996 (O_2996,N_24188,N_24662);
or UO_2997 (O_2997,N_24198,N_24381);
or UO_2998 (O_2998,N_24736,N_24890);
nor UO_2999 (O_2999,N_24471,N_24753);
endmodule