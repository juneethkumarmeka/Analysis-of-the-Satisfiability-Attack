module basic_2500_25000_3000_5_levels_5xor_4(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999;
nor U0 (N_0,In_821,In_2367);
and U1 (N_1,In_2353,In_1705);
or U2 (N_2,In_725,In_69);
nor U3 (N_3,In_132,In_833);
nor U4 (N_4,In_1713,In_949);
nand U5 (N_5,In_2309,In_1220);
nand U6 (N_6,In_2371,In_1081);
xor U7 (N_7,In_883,In_1632);
or U8 (N_8,In_535,In_727);
nor U9 (N_9,In_1960,In_1766);
or U10 (N_10,In_1091,In_360);
nor U11 (N_11,In_506,In_2108);
nor U12 (N_12,In_434,In_967);
and U13 (N_13,In_2124,In_410);
xnor U14 (N_14,In_60,In_548);
or U15 (N_15,In_1250,In_287);
or U16 (N_16,In_3,In_2094);
or U17 (N_17,In_311,In_910);
nor U18 (N_18,In_464,In_2217);
nor U19 (N_19,In_1127,In_773);
nor U20 (N_20,In_1404,In_553);
or U21 (N_21,In_67,In_2191);
nor U22 (N_22,In_622,In_640);
and U23 (N_23,In_2223,In_1102);
or U24 (N_24,In_1697,In_73);
nand U25 (N_25,In_181,In_1674);
nor U26 (N_26,In_2262,In_1225);
nor U27 (N_27,In_1295,In_1280);
or U28 (N_28,In_816,In_194);
nor U29 (N_29,In_1971,In_306);
or U30 (N_30,In_2358,In_1039);
nand U31 (N_31,In_1712,In_2376);
nand U32 (N_32,In_184,In_1930);
or U33 (N_33,In_2374,In_722);
nand U34 (N_34,In_1851,In_2026);
and U35 (N_35,In_30,In_644);
and U36 (N_36,In_323,In_361);
xnor U37 (N_37,In_766,In_1980);
or U38 (N_38,In_403,In_242);
or U39 (N_39,In_927,In_1588);
nand U40 (N_40,In_2206,In_1579);
nand U41 (N_41,In_2444,In_1140);
nand U42 (N_42,In_704,In_587);
nand U43 (N_43,In_2265,In_1950);
and U44 (N_44,In_1887,In_782);
or U45 (N_45,In_1551,In_613);
nand U46 (N_46,In_1163,In_2413);
nor U47 (N_47,In_527,In_583);
nand U48 (N_48,In_1360,In_2000);
xnor U49 (N_49,In_335,In_2137);
and U50 (N_50,In_2150,In_2487);
or U51 (N_51,In_1745,In_1424);
and U52 (N_52,In_2233,In_2245);
and U53 (N_53,In_532,In_777);
nand U54 (N_54,In_1032,In_2404);
nor U55 (N_55,In_1235,In_1903);
or U56 (N_56,In_59,In_747);
or U57 (N_57,In_1353,In_693);
or U58 (N_58,In_1033,In_1813);
nor U59 (N_59,In_1179,In_1724);
xnor U60 (N_60,In_51,In_761);
nor U61 (N_61,In_2337,In_1227);
and U62 (N_62,In_947,In_2461);
nor U63 (N_63,In_516,In_1336);
or U64 (N_64,In_2342,In_364);
nand U65 (N_65,In_1349,In_1202);
or U66 (N_66,In_2095,In_2441);
nand U67 (N_67,In_2381,In_2133);
nand U68 (N_68,In_2119,In_913);
nor U69 (N_69,In_2323,In_402);
nor U70 (N_70,In_1271,In_1583);
or U71 (N_71,In_1332,In_1325);
nor U72 (N_72,In_2406,In_749);
and U73 (N_73,In_246,In_209);
nand U74 (N_74,In_1307,In_1512);
or U75 (N_75,In_860,In_524);
and U76 (N_76,In_1728,In_2230);
nand U77 (N_77,In_1617,In_938);
or U78 (N_78,In_353,In_685);
nand U79 (N_79,In_1226,In_2134);
nand U80 (N_80,In_1460,In_1900);
or U81 (N_81,In_750,In_2391);
or U82 (N_82,In_2295,In_2074);
or U83 (N_83,In_2473,In_1982);
nand U84 (N_84,In_1340,In_1078);
xnor U85 (N_85,In_1389,In_479);
nand U86 (N_86,In_2048,In_661);
or U87 (N_87,In_2215,In_1128);
xor U88 (N_88,In_591,In_1186);
nand U89 (N_89,In_957,In_1578);
nand U90 (N_90,In_2282,In_2332);
nor U91 (N_91,In_128,In_1470);
or U92 (N_92,In_44,In_2116);
nand U93 (N_93,In_656,In_2361);
or U94 (N_94,In_814,In_2152);
nor U95 (N_95,In_1774,In_2315);
nand U96 (N_96,In_2314,In_2477);
nor U97 (N_97,In_373,In_966);
or U98 (N_98,In_1620,In_953);
nand U99 (N_99,In_902,In_1953);
xor U100 (N_100,In_1158,In_376);
or U101 (N_101,In_1937,In_309);
nand U102 (N_102,In_564,In_372);
or U103 (N_103,In_1863,In_114);
nand U104 (N_104,In_1939,In_2159);
or U105 (N_105,In_998,In_1204);
or U106 (N_106,In_793,In_1594);
xor U107 (N_107,In_174,In_11);
nor U108 (N_108,In_1639,In_743);
or U109 (N_109,In_1875,In_2260);
or U110 (N_110,In_1795,In_1597);
and U111 (N_111,In_1616,In_24);
and U112 (N_112,In_476,In_419);
nor U113 (N_113,In_256,In_1439);
nor U114 (N_114,In_248,In_1309);
nand U115 (N_115,In_1839,In_1775);
or U116 (N_116,In_1811,In_1831);
nor U117 (N_117,In_960,In_121);
nor U118 (N_118,In_2242,In_2446);
nand U119 (N_119,In_2231,In_1941);
nor U120 (N_120,In_58,In_1880);
or U121 (N_121,In_1466,In_2436);
nand U122 (N_122,In_342,In_838);
nand U123 (N_123,In_1672,In_2033);
and U124 (N_124,In_1195,In_1363);
nand U125 (N_125,In_278,In_507);
and U126 (N_126,In_2083,In_956);
nor U127 (N_127,In_1454,In_284);
nor U128 (N_128,In_299,In_1281);
or U129 (N_129,In_1592,In_2059);
nor U130 (N_130,In_258,In_76);
and U131 (N_131,In_490,In_64);
nor U132 (N_132,In_254,In_33);
and U133 (N_133,In_842,In_2345);
nor U134 (N_134,In_16,In_120);
nand U135 (N_135,In_1114,In_2478);
nor U136 (N_136,In_1737,In_540);
nor U137 (N_137,In_2271,In_433);
xor U138 (N_138,In_1997,In_2);
nand U139 (N_139,In_2110,In_1191);
xor U140 (N_140,In_1729,In_815);
xnor U141 (N_141,In_1254,In_1432);
or U142 (N_142,In_1571,In_1874);
nand U143 (N_143,In_2330,In_1515);
and U144 (N_144,In_559,In_1096);
nor U145 (N_145,In_374,In_878);
and U146 (N_146,In_1927,In_1733);
nand U147 (N_147,In_362,In_710);
nand U148 (N_148,In_1399,In_1804);
and U149 (N_149,In_634,In_269);
nor U150 (N_150,In_897,In_2034);
nand U151 (N_151,In_1929,In_1159);
nand U152 (N_152,In_2320,In_2160);
nor U153 (N_153,In_615,In_1170);
and U154 (N_154,In_1287,In_1582);
nand U155 (N_155,In_454,In_53);
nand U156 (N_156,In_713,In_443);
xnor U157 (N_157,In_500,In_1074);
nand U158 (N_158,In_684,In_1099);
nand U159 (N_159,In_2174,In_1650);
and U160 (N_160,In_1896,In_2482);
nor U161 (N_161,In_46,In_397);
nor U162 (N_162,In_2486,In_2300);
nor U163 (N_163,In_980,In_983);
nand U164 (N_164,In_590,In_2302);
xor U165 (N_165,In_682,In_347);
xor U166 (N_166,In_890,In_936);
xor U167 (N_167,In_230,In_1507);
xor U168 (N_168,In_2331,In_2355);
nand U169 (N_169,In_762,In_1272);
nand U170 (N_170,In_260,In_455);
nor U171 (N_171,In_146,In_2415);
or U172 (N_172,In_292,In_2283);
or U173 (N_173,In_1805,In_700);
or U174 (N_174,In_432,In_934);
or U175 (N_175,In_848,In_151);
xnor U176 (N_176,In_2209,In_1637);
or U177 (N_177,In_442,In_2165);
nor U178 (N_178,In_1,In_914);
nor U179 (N_179,In_2204,In_1669);
nor U180 (N_180,In_2025,In_2259);
nor U181 (N_181,In_1700,In_937);
nor U182 (N_182,In_1401,In_1249);
or U183 (N_183,In_2229,In_745);
and U184 (N_184,In_972,In_1122);
and U185 (N_185,In_2328,In_1567);
nor U186 (N_186,In_1921,In_1867);
xor U187 (N_187,In_889,In_1564);
nor U188 (N_188,In_529,In_893);
nor U189 (N_189,In_1498,In_203);
or U190 (N_190,In_90,In_2449);
and U191 (N_191,In_1345,In_961);
or U192 (N_192,In_2481,In_2219);
xnor U193 (N_193,In_257,In_1502);
nor U194 (N_194,In_1691,In_1403);
or U195 (N_195,In_794,In_1386);
or U196 (N_196,In_1025,In_1801);
and U197 (N_197,In_1414,In_1964);
nand U198 (N_198,In_2032,In_1892);
xnor U199 (N_199,In_593,In_2263);
and U200 (N_200,In_2009,In_1850);
nor U201 (N_201,In_2424,In_2344);
or U202 (N_202,In_267,In_769);
xnor U203 (N_203,In_1459,In_1208);
or U204 (N_204,In_1685,In_1837);
nor U205 (N_205,In_1082,In_941);
nand U206 (N_206,In_1180,In_1968);
and U207 (N_207,In_1715,In_1017);
nand U208 (N_208,In_539,In_1488);
nand U209 (N_209,In_499,In_222);
or U210 (N_210,In_1977,In_1716);
nand U211 (N_211,In_1561,In_1311);
nor U212 (N_212,In_15,In_2427);
or U213 (N_213,In_711,In_185);
or U214 (N_214,In_1653,In_1086);
xor U215 (N_215,In_217,In_1651);
and U216 (N_216,In_896,In_1750);
or U217 (N_217,In_720,In_1652);
nor U218 (N_218,In_2196,In_71);
and U219 (N_219,In_2352,In_1031);
or U220 (N_220,In_1269,In_669);
or U221 (N_221,In_1814,In_2128);
or U222 (N_222,In_1238,In_996);
nand U223 (N_223,In_1731,In_510);
xor U224 (N_224,In_1215,In_224);
and U225 (N_225,In_1398,In_449);
xor U226 (N_226,In_2222,In_1264);
or U227 (N_227,In_850,In_1011);
nand U228 (N_228,In_1261,In_1445);
nand U229 (N_229,In_965,In_1560);
nor U230 (N_230,In_776,In_118);
and U231 (N_231,In_265,In_32);
or U232 (N_232,In_1618,In_1566);
nor U233 (N_233,In_2170,In_52);
nor U234 (N_234,In_2101,In_66);
nand U235 (N_235,In_2483,In_1640);
nor U236 (N_236,In_45,In_2372);
nand U237 (N_237,In_1768,In_2365);
or U238 (N_238,In_467,In_1647);
nand U239 (N_239,In_199,In_2258);
nor U240 (N_240,In_509,In_2416);
and U241 (N_241,In_1144,In_135);
and U242 (N_242,In_1408,In_551);
nand U243 (N_243,In_1040,In_1510);
nand U244 (N_244,In_456,In_85);
nor U245 (N_245,In_923,In_1948);
nor U246 (N_246,In_1256,In_742);
and U247 (N_247,In_512,In_1243);
nand U248 (N_248,In_1660,In_2202);
nor U249 (N_249,In_993,In_918);
nor U250 (N_250,In_1166,In_2243);
nand U251 (N_251,In_1075,In_1423);
and U252 (N_252,In_2126,In_220);
nor U253 (N_253,In_475,In_2154);
or U254 (N_254,In_1026,In_674);
nand U255 (N_255,In_473,In_1662);
nand U256 (N_256,In_1276,In_1781);
and U257 (N_257,In_1574,In_1956);
nand U258 (N_258,In_1558,In_2179);
and U259 (N_259,In_1629,In_2253);
and U260 (N_260,In_378,In_2019);
nor U261 (N_261,In_1743,In_1120);
and U262 (N_262,In_886,In_1211);
or U263 (N_263,In_2426,In_1077);
and U264 (N_264,In_2285,In_317);
nor U265 (N_265,In_137,In_2383);
or U266 (N_266,In_515,In_2364);
or U267 (N_267,In_631,In_1701);
nor U268 (N_268,In_1151,In_420);
or U269 (N_269,In_581,In_1036);
nor U270 (N_270,In_2192,In_2220);
nor U271 (N_271,In_903,In_817);
nand U272 (N_272,In_2425,In_554);
nand U273 (N_273,In_1904,In_321);
nor U274 (N_274,In_1698,In_493);
nor U275 (N_275,In_1736,In_1044);
nand U276 (N_276,In_2004,In_1293);
and U277 (N_277,In_2490,In_251);
or U278 (N_278,In_1193,In_399);
nor U279 (N_279,In_1954,In_329);
nor U280 (N_280,In_2351,In_1499);
or U281 (N_281,In_1570,In_416);
nand U282 (N_282,In_2306,In_2072);
nand U283 (N_283,In_2378,In_1614);
nor U284 (N_284,In_54,In_1456);
and U285 (N_285,In_1236,In_1174);
nor U286 (N_286,In_1189,In_840);
or U287 (N_287,In_1504,In_1885);
nand U288 (N_288,In_1059,In_2363);
xor U289 (N_289,In_1819,In_1992);
or U290 (N_290,In_423,In_2054);
nor U291 (N_291,In_2311,In_1374);
or U292 (N_292,In_1975,In_1920);
and U293 (N_293,In_4,In_2275);
and U294 (N_294,In_1428,In_1710);
or U295 (N_295,In_1440,In_351);
and U296 (N_296,In_2147,In_310);
and U297 (N_297,In_1371,In_2168);
or U298 (N_298,In_228,In_169);
nand U299 (N_299,In_1562,In_1200);
nand U300 (N_300,In_979,In_407);
xor U301 (N_301,In_1829,In_1649);
or U302 (N_302,In_20,In_2050);
or U303 (N_303,In_1780,In_1330);
nand U304 (N_304,In_1142,In_2341);
nor U305 (N_305,In_2014,In_2234);
nand U306 (N_306,In_812,In_330);
nor U307 (N_307,In_1988,In_789);
nand U308 (N_308,In_1344,In_1239);
or U309 (N_309,In_1268,In_1708);
and U310 (N_310,In_1480,In_1922);
nand U311 (N_311,In_1334,In_806);
and U312 (N_312,In_2312,In_89);
or U313 (N_313,In_1857,In_731);
or U314 (N_314,In_678,In_2431);
nor U315 (N_315,In_2296,In_1914);
nor U316 (N_316,In_874,In_1773);
or U317 (N_317,In_431,In_1931);
or U318 (N_318,In_1265,In_546);
and U319 (N_319,In_569,In_763);
and U320 (N_320,In_675,In_1905);
or U321 (N_321,In_1240,In_1732);
and U322 (N_322,In_1491,In_668);
and U323 (N_323,In_1843,In_2278);
and U324 (N_324,In_2380,In_1019);
xnor U325 (N_325,In_2041,In_86);
nand U326 (N_326,In_568,In_1071);
xor U327 (N_327,In_945,In_715);
or U328 (N_328,In_1520,In_1110);
or U329 (N_329,In_161,In_2304);
nor U330 (N_330,In_2244,In_809);
xnor U331 (N_331,In_2452,In_1744);
and U332 (N_332,In_383,In_1521);
xnor U333 (N_333,In_2286,In_2075);
or U334 (N_334,In_468,In_608);
and U335 (N_335,In_1377,In_709);
nand U336 (N_336,In_1161,In_1767);
and U337 (N_337,In_435,In_2102);
xor U338 (N_338,In_1052,In_892);
nand U339 (N_339,In_1476,In_925);
nand U340 (N_340,In_1757,In_1915);
and U341 (N_341,In_1546,In_714);
and U342 (N_342,In_628,In_599);
nand U343 (N_343,In_110,In_692);
and U344 (N_344,In_1109,In_1884);
and U345 (N_345,In_982,In_1633);
or U346 (N_346,In_1497,In_1323);
xor U347 (N_347,In_2162,In_2011);
or U348 (N_348,In_2013,In_1846);
xnor U349 (N_349,In_577,In_1918);
or U350 (N_350,In_2002,In_999);
nor U351 (N_351,In_1262,In_1746);
xor U352 (N_352,In_1636,In_2068);
or U353 (N_353,In_40,In_2113);
or U354 (N_354,In_1910,In_1119);
nor U355 (N_355,In_345,In_2027);
nor U356 (N_356,In_116,In_803);
or U357 (N_357,In_650,In_2280);
and U358 (N_358,In_1835,In_630);
and U359 (N_359,In_677,In_520);
xnor U360 (N_360,In_2333,In_603);
and U361 (N_361,In_839,In_1783);
nor U362 (N_362,In_514,In_202);
nor U363 (N_363,In_325,In_272);
and U364 (N_364,In_2012,In_1419);
and U365 (N_365,In_2135,In_1027);
or U366 (N_366,In_2293,In_1245);
nor U367 (N_367,In_1694,In_1348);
nor U368 (N_368,In_1912,In_2190);
nor U369 (N_369,In_853,In_1518);
nor U370 (N_370,In_2069,In_1290);
or U371 (N_371,In_1763,In_2484);
nor U372 (N_372,In_1641,In_7);
or U373 (N_373,In_1343,In_2003);
and U374 (N_374,In_415,In_666);
or U375 (N_375,In_2397,In_1544);
and U376 (N_376,In_1500,In_1381);
nand U377 (N_377,In_1508,In_88);
xor U378 (N_378,In_83,In_707);
nand U379 (N_379,In_1505,In_1690);
nand U380 (N_380,In_505,In_332);
or U381 (N_381,In_138,In_1065);
and U382 (N_382,In_1949,In_1598);
or U383 (N_383,In_845,In_75);
nand U384 (N_384,In_2479,In_1793);
nor U385 (N_385,In_328,In_648);
nor U386 (N_386,In_1187,In_275);
and U387 (N_387,In_1324,In_1387);
nor U388 (N_388,In_1755,In_2457);
and U389 (N_389,In_2281,In_2439);
nor U390 (N_390,In_606,In_1608);
or U391 (N_391,In_542,In_1972);
nand U392 (N_392,In_129,In_1447);
or U393 (N_393,In_969,In_1085);
or U394 (N_394,In_1625,In_1003);
nor U395 (N_395,In_741,In_991);
nand U396 (N_396,In_1361,In_1658);
or U397 (N_397,In_736,In_767);
nor U398 (N_398,In_98,In_296);
nand U399 (N_399,In_227,In_1932);
and U400 (N_400,In_905,In_43);
and U401 (N_401,In_37,In_189);
nor U402 (N_402,In_1292,In_2145);
nand U403 (N_403,In_754,In_786);
xor U404 (N_404,In_933,In_825);
and U405 (N_405,In_641,In_1329);
xor U406 (N_406,In_1199,In_438);
nor U407 (N_407,In_1366,In_1540);
nor U408 (N_408,In_2065,In_1494);
nor U409 (N_409,In_852,In_105);
xnor U410 (N_410,In_274,In_653);
or U411 (N_411,In_642,In_2335);
xnor U412 (N_412,In_450,In_1824);
nand U413 (N_413,In_2136,In_654);
nor U414 (N_414,In_91,In_2467);
nor U415 (N_415,In_1224,In_2084);
and U416 (N_416,In_1664,In_1635);
nand U417 (N_417,In_344,In_1911);
nor U418 (N_418,In_1942,In_1084);
and U419 (N_419,In_2496,In_1316);
nor U420 (N_420,In_101,In_2148);
nand U421 (N_421,In_1945,In_2232);
nand U422 (N_422,In_1565,In_1899);
or U423 (N_423,In_1661,In_1792);
and U424 (N_424,In_1034,In_1529);
nand U425 (N_425,In_1441,In_2182);
or U426 (N_426,In_521,In_322);
or U427 (N_427,In_2326,In_1858);
nor U428 (N_428,In_47,In_1986);
and U429 (N_429,In_1060,In_1994);
nor U430 (N_430,In_901,In_1021);
or U431 (N_431,In_1545,In_352);
and U432 (N_432,In_2151,In_1646);
nor U433 (N_433,In_2188,In_462);
nand U434 (N_434,In_2146,In_1559);
nand U435 (N_435,In_457,In_526);
nor U436 (N_436,In_2158,In_863);
nor U437 (N_437,In_2430,In_125);
nor U438 (N_438,In_82,In_1178);
or U439 (N_439,In_975,In_234);
nor U440 (N_440,In_1001,In_314);
nand U441 (N_441,In_728,In_2298);
or U442 (N_442,In_1897,In_1602);
and U443 (N_443,In_1798,In_2247);
or U444 (N_444,In_1258,In_688);
or U445 (N_445,In_180,In_1749);
nor U446 (N_446,In_846,In_319);
or U447 (N_447,In_2035,In_1943);
and U448 (N_448,In_2103,In_1513);
nor U449 (N_449,In_1908,In_193);
and U450 (N_450,In_1064,In_1524);
nor U451 (N_451,In_1042,In_2339);
nand U452 (N_452,In_734,In_103);
and U453 (N_453,In_210,In_977);
nand U454 (N_454,In_788,In_156);
and U455 (N_455,In_2143,In_1596);
and U456 (N_456,In_25,In_229);
nor U457 (N_457,In_1058,In_2305);
and U458 (N_458,In_1709,In_1072);
and U459 (N_459,In_876,In_1828);
nor U460 (N_460,In_1823,In_34);
xor U461 (N_461,In_2429,In_147);
or U462 (N_462,In_1877,In_84);
nor U463 (N_463,In_504,In_488);
nor U464 (N_464,In_1010,In_1587);
xor U465 (N_465,In_1740,In_1742);
nand U466 (N_466,In_2086,In_1963);
nand U467 (N_467,In_1359,In_1467);
or U468 (N_468,In_1643,In_213);
nand U469 (N_469,In_1300,In_1893);
nand U470 (N_470,In_2031,In_679);
xnor U471 (N_471,In_643,In_1981);
nor U472 (N_472,In_2419,In_276);
nor U473 (N_473,In_658,In_2052);
nand U474 (N_474,In_501,In_1868);
nor U475 (N_475,In_440,In_729);
xnor U476 (N_476,In_609,In_2277);
nand U477 (N_477,In_293,In_1004);
or U478 (N_478,In_1420,In_1248);
and U479 (N_479,In_1808,In_1156);
nor U480 (N_480,In_1628,In_1418);
nor U481 (N_481,In_149,In_2403);
and U482 (N_482,In_827,In_2212);
xor U483 (N_483,In_1063,In_1785);
or U484 (N_484,In_1770,In_584);
or U485 (N_485,In_1861,In_1146);
nor U486 (N_486,In_2017,In_396);
or U487 (N_487,In_404,In_177);
or U488 (N_488,In_1341,In_1397);
or U489 (N_489,In_1041,In_1591);
or U490 (N_490,In_358,In_139);
nor U491 (N_491,In_541,In_1400);
nand U492 (N_492,In_1849,In_1306);
nand U493 (N_493,In_141,In_1326);
nor U494 (N_494,In_952,In_2297);
xor U495 (N_495,In_1989,In_676);
and U496 (N_496,In_2303,In_408);
and U497 (N_497,In_563,In_142);
or U498 (N_498,In_703,In_2241);
xor U499 (N_499,In_2301,In_2294);
nand U500 (N_500,In_1362,In_2347);
xor U501 (N_501,In_572,In_544);
nor U502 (N_502,In_390,In_708);
nor U503 (N_503,In_849,In_1879);
or U504 (N_504,In_2433,In_779);
and U505 (N_505,In_600,In_958);
and U506 (N_506,In_1465,In_695);
nor U507 (N_507,In_381,In_757);
nand U508 (N_508,In_701,In_2197);
nand U509 (N_509,In_2238,In_122);
or U510 (N_510,In_2125,In_623);
nor U511 (N_511,In_2288,In_1531);
nor U512 (N_512,In_875,In_1229);
nand U513 (N_513,In_2428,In_1097);
nor U514 (N_514,In_205,In_1279);
nand U515 (N_515,In_1006,In_1369);
nand U516 (N_516,In_1047,In_318);
or U517 (N_517,In_931,In_2121);
nor U518 (N_518,In_2104,In_626);
nand U519 (N_519,In_206,In_2016);
and U520 (N_520,In_2099,In_1543);
nor U521 (N_521,In_2474,In_1575);
nand U522 (N_522,In_38,In_1748);
nand U523 (N_523,In_1055,In_2184);
nor U524 (N_524,In_724,In_22);
xor U525 (N_525,In_1503,In_2499);
nor U526 (N_526,In_525,In_1130);
or U527 (N_527,In_494,In_2491);
or U528 (N_528,In_2393,In_57);
nand U529 (N_529,In_18,In_2088);
nor U530 (N_530,In_1080,In_2357);
and U531 (N_531,In_607,In_215);
or U532 (N_532,In_637,In_1385);
and U533 (N_533,In_1217,In_212);
or U534 (N_534,In_1969,In_106);
nand U535 (N_535,In_1557,In_2161);
nand U536 (N_536,In_1511,In_1103);
nor U537 (N_537,In_739,In_1133);
or U538 (N_538,In_962,In_1985);
nor U539 (N_539,In_1528,In_486);
nor U540 (N_540,In_451,In_900);
or U541 (N_541,In_130,In_124);
and U542 (N_542,In_1426,In_697);
nand U543 (N_543,In_2468,In_1354);
nor U544 (N_544,In_2316,In_1286);
or U545 (N_545,In_772,In_1169);
nand U546 (N_546,In_262,In_774);
or U547 (N_547,In_1944,In_1143);
and U548 (N_548,In_1391,In_1378);
or U549 (N_549,In_1882,In_1132);
nand U550 (N_550,In_1294,In_158);
nor U551 (N_551,In_1194,In_1536);
nand U552 (N_552,In_19,In_197);
or U553 (N_553,In_1895,In_1422);
and U554 (N_554,In_289,In_2096);
nor U555 (N_555,In_411,In_1952);
nand U556 (N_556,In_1462,In_1112);
nor U557 (N_557,In_1541,In_756);
nand U558 (N_558,In_1802,In_986);
nand U559 (N_559,In_36,In_1607);
and U560 (N_560,In_102,In_557);
nor U561 (N_561,In_547,In_398);
or U562 (N_562,In_368,In_2465);
nand U563 (N_563,In_2193,In_469);
or U564 (N_564,In_1610,In_981);
nor U565 (N_565,In_698,In_1255);
or U566 (N_566,In_444,In_2251);
nand U567 (N_567,In_1150,In_1585);
nor U568 (N_568,In_1832,In_1527);
nor U569 (N_569,In_2062,In_1364);
nand U570 (N_570,In_1393,In_785);
nand U571 (N_571,In_2382,In_439);
and U572 (N_572,In_1417,In_99);
nor U573 (N_573,In_929,In_2249);
nor U574 (N_574,In_2422,In_2390);
and U575 (N_575,In_759,In_1367);
xor U576 (N_576,In_297,In_2049);
nand U577 (N_577,In_477,In_1394);
nand U578 (N_578,In_441,In_582);
nand U579 (N_579,In_81,In_2180);
or U580 (N_580,In_1656,In_190);
nand U581 (N_581,In_992,In_1600);
and U582 (N_582,In_1926,In_2144);
nor U583 (N_583,In_2153,In_195);
and U584 (N_584,In_1093,In_2284);
nor U585 (N_585,In_2476,In_1232);
xor U586 (N_586,In_2020,In_625);
xor U587 (N_587,In_882,In_471);
and U588 (N_588,In_1320,In_2336);
nor U589 (N_589,In_1589,In_166);
nand U590 (N_590,In_183,In_1259);
xnor U591 (N_591,In_1117,In_1492);
nand U592 (N_592,In_856,In_744);
or U593 (N_593,In_459,In_2213);
and U594 (N_594,In_884,In_2132);
xor U595 (N_595,In_1305,In_348);
nor U596 (N_596,In_263,In_2167);
or U597 (N_597,In_2093,In_1212);
nand U598 (N_598,In_990,In_820);
xor U599 (N_599,In_336,In_2292);
nor U600 (N_600,In_1384,In_77);
nor U601 (N_601,In_42,In_472);
and U602 (N_602,In_68,In_1807);
and U603 (N_603,In_2343,In_796);
xor U604 (N_604,In_2409,In_1427);
and U605 (N_605,In_1779,In_1197);
and U606 (N_606,In_808,In_270);
nor U607 (N_607,In_338,In_1335);
and U608 (N_608,In_1889,In_517);
xnor U609 (N_609,In_1153,In_1553);
xnor U610 (N_610,In_1535,In_823);
and U611 (N_611,In_119,In_175);
nor U612 (N_612,In_616,In_1175);
xor U613 (N_613,In_2256,In_2080);
and U614 (N_614,In_244,In_621);
xnor U615 (N_615,In_2402,In_1350);
xor U616 (N_616,In_1318,In_813);
or U617 (N_617,In_915,In_872);
nand U618 (N_618,In_1630,In_2495);
nor U619 (N_619,In_1452,In_1425);
nor U620 (N_620,In_2432,In_1727);
nand U621 (N_621,In_1090,In_596);
and U622 (N_622,In_312,In_926);
or U623 (N_623,In_690,In_409);
nor U624 (N_624,In_133,In_1296);
nand U625 (N_625,In_253,In_271);
nor U626 (N_626,In_1431,In_906);
or U627 (N_627,In_1782,In_895);
xor U628 (N_628,In_1444,In_1554);
nor U629 (N_629,In_1667,In_841);
nor U630 (N_630,In_1501,In_1834);
nor U631 (N_631,In_2440,In_375);
xnor U632 (N_632,In_1778,In_426);
or U633 (N_633,In_2420,In_851);
or U634 (N_634,In_1023,In_1627);
or U635 (N_635,In_1182,In_2200);
nor U636 (N_636,In_755,In_2463);
and U637 (N_637,In_2010,In_847);
and U638 (N_638,In_1680,In_924);
and U639 (N_639,In_810,In_732);
or U640 (N_640,In_1152,In_1984);
nand U641 (N_641,In_948,In_888);
nand U642 (N_642,In_1678,In_1888);
nor U643 (N_643,In_2157,In_2071);
or U644 (N_644,In_1449,In_1437);
nand U645 (N_645,In_1210,In_1057);
and U646 (N_646,In_595,In_921);
nand U647 (N_647,In_696,In_31);
and U648 (N_648,In_2462,In_1881);
and U649 (N_649,In_87,In_487);
and U650 (N_650,In_2254,In_2239);
and U651 (N_651,In_489,In_1263);
xnor U652 (N_652,In_160,In_370);
nand U653 (N_653,In_1747,In_1067);
or U654 (N_654,In_1853,In_1718);
nor U655 (N_655,In_2272,In_916);
and U656 (N_656,In_2362,In_49);
or U657 (N_657,In_1517,In_2115);
nor U658 (N_658,In_1869,In_341);
nor U659 (N_659,In_1372,In_1886);
nor U660 (N_660,In_1991,In_2356);
nand U661 (N_661,In_1176,In_1671);
nor U662 (N_662,In_2266,In_406);
or U663 (N_663,In_288,In_1720);
nor U664 (N_664,In_2181,In_346);
or U665 (N_665,In_1809,In_1907);
nand U666 (N_666,In_2079,In_718);
nor U667 (N_667,In_1689,In_2081);
nand U668 (N_668,In_1822,In_908);
and U669 (N_669,In_1406,In_327);
xnor U670 (N_670,In_706,In_112);
nand U671 (N_671,In_123,In_1840);
nor U672 (N_672,In_1430,In_2106);
nand U673 (N_673,In_143,In_1357);
or U674 (N_674,In_324,In_1909);
nand U675 (N_675,In_478,In_2221);
or U676 (N_676,In_1753,In_1358);
or U677 (N_677,In_482,In_150);
or U678 (N_678,In_1407,In_2276);
and U679 (N_679,In_824,In_1872);
or U680 (N_680,In_1160,In_864);
or U681 (N_681,In_1957,In_955);
or U682 (N_682,In_1810,In_1477);
nor U683 (N_683,In_178,In_1569);
nor U684 (N_684,In_522,In_805);
nand U685 (N_685,In_61,In_1730);
nand U686 (N_686,In_2471,In_392);
nor U687 (N_687,In_333,In_1523);
nand U688 (N_688,In_687,In_2090);
nand U689 (N_689,In_453,In_1018);
and U690 (N_690,In_1009,In_1157);
xor U691 (N_691,In_23,In_491);
nand U692 (N_692,In_1368,In_1221);
nor U693 (N_693,In_208,In_2291);
nand U694 (N_694,In_386,In_1319);
nor U695 (N_695,In_571,In_2493);
or U696 (N_696,In_617,In_1684);
or U697 (N_697,In_873,In_1866);
and U698 (N_698,In_534,In_1842);
xor U699 (N_699,In_313,In_1666);
nor U700 (N_700,In_508,In_80);
and U701 (N_701,In_2171,In_2317);
and U702 (N_702,In_1821,In_870);
xor U703 (N_703,In_1721,In_2227);
and U704 (N_704,In_1472,In_1676);
and U705 (N_705,In_401,In_295);
nand U706 (N_706,In_1891,In_1734);
nand U707 (N_707,In_2114,In_1273);
nand U708 (N_708,In_294,In_780);
or U709 (N_709,In_586,In_1219);
or U710 (N_710,In_738,In_950);
nand U711 (N_711,In_1833,In_252);
or U712 (N_712,In_588,In_1644);
xnor U713 (N_713,In_1266,In_1576);
nor U714 (N_714,In_2042,In_1754);
and U715 (N_715,In_2257,In_2111);
or U716 (N_716,In_1020,In_951);
or U717 (N_717,In_393,In_605);
and U718 (N_718,In_1190,In_2248);
or U719 (N_719,In_1234,In_1129);
and U720 (N_720,In_286,In_662);
nor U721 (N_721,In_1648,In_2001);
nand U722 (N_722,In_273,In_2109);
and U723 (N_723,In_250,In_1464);
nor U724 (N_724,In_349,In_597);
nor U725 (N_725,In_1482,In_1681);
nor U726 (N_726,In_1222,In_2489);
nand U727 (N_727,In_1495,In_954);
and U728 (N_728,In_1141,In_2058);
and U729 (N_729,In_1380,In_1446);
nand U730 (N_730,In_795,In_2226);
and U731 (N_731,In_1919,In_1762);
nor U732 (N_732,In_2379,In_837);
nand U733 (N_733,In_1390,In_2290);
xnor U734 (N_734,In_1841,In_1605);
or U735 (N_735,In_148,In_1304);
xor U736 (N_736,In_1759,In_2321);
or U737 (N_737,In_748,In_2028);
nand U738 (N_738,In_1966,In_320);
nor U739 (N_739,In_787,In_13);
xnor U740 (N_740,In_1463,In_2030);
or U741 (N_741,In_1458,In_1274);
and U742 (N_742,In_2060,In_369);
nand U743 (N_743,In_928,In_726);
nor U744 (N_744,In_277,In_1634);
and U745 (N_745,In_1183,In_359);
nor U746 (N_746,In_480,In_1167);
nand U747 (N_747,In_2046,In_186);
nand U748 (N_748,In_2454,In_618);
or U749 (N_749,In_1735,In_1601);
nand U750 (N_750,In_1365,In_1095);
nand U751 (N_751,In_2036,In_2389);
or U752 (N_752,In_533,In_2299);
nor U753 (N_753,In_1312,In_778);
nor U754 (N_754,In_939,In_1246);
and U755 (N_755,In_55,In_1015);
or U756 (N_756,In_1797,In_2497);
nand U757 (N_757,In_604,In_502);
and U758 (N_758,In_2319,In_2414);
nand U759 (N_759,In_418,In_2224);
and U760 (N_760,In_1088,In_1164);
xnor U761 (N_761,In_1356,In_232);
xor U762 (N_762,In_2423,In_1764);
nand U763 (N_763,In_1453,In_1302);
nand U764 (N_764,In_624,In_855);
nor U765 (N_765,In_1029,In_784);
nor U766 (N_766,In_496,In_1752);
and U767 (N_767,In_95,In_2194);
and U768 (N_768,In_41,In_1894);
or U769 (N_769,In_448,In_1707);
or U770 (N_770,In_619,In_460);
nor U771 (N_771,In_1089,In_2120);
and U772 (N_772,In_1990,In_1845);
xor U773 (N_773,In_1496,In_6);
or U774 (N_774,In_1121,In_1116);
nand U775 (N_775,In_1549,In_366);
nor U776 (N_776,In_2417,In_282);
and U777 (N_777,In_236,In_1469);
xor U778 (N_778,In_2172,In_1277);
or U779 (N_779,In_316,In_667);
nand U780 (N_780,In_2240,In_1642);
or U781 (N_781,In_307,In_1855);
xor U782 (N_782,In_247,In_340);
nand U783 (N_783,In_2396,In_1218);
nand U784 (N_784,In_1609,In_2123);
and U785 (N_785,In_943,In_93);
nor U786 (N_786,In_1534,In_1624);
and U787 (N_787,In_1012,In_549);
nand U788 (N_788,In_1124,In_164);
and U789 (N_789,In_1675,In_1902);
nor U790 (N_790,In_1976,In_1673);
nor U791 (N_791,In_1196,In_470);
nand U792 (N_792,In_1291,In_163);
and U793 (N_793,In_1233,In_2261);
and U794 (N_794,In_279,In_2398);
nor U795 (N_795,In_1475,In_1933);
or U796 (N_796,In_594,In_1228);
nor U797 (N_797,In_2408,In_1631);
nor U798 (N_798,In_1856,In_2040);
nor U799 (N_799,In_865,In_1703);
nand U800 (N_800,In_1339,In_1936);
or U801 (N_801,In_1765,In_1198);
nor U802 (N_802,In_2273,In_223);
and U803 (N_803,In_665,In_2360);
and U804 (N_804,In_1862,In_237);
nor U805 (N_805,In_758,In_1205);
or U806 (N_806,In_5,In_2329);
nor U807 (N_807,In_1315,In_1448);
nand U808 (N_808,In_1471,In_836);
and U809 (N_809,In_167,In_2472);
and U810 (N_810,In_1978,In_1136);
xnor U811 (N_811,In_1815,In_1370);
and U812 (N_812,In_1351,In_179);
xor U813 (N_813,In_377,In_1230);
and U814 (N_814,In_2434,In_1168);
nand U815 (N_815,In_238,In_154);
and U816 (N_816,In_134,In_1794);
nor U817 (N_817,In_1595,In_694);
nand U818 (N_818,In_1995,In_917);
xnor U819 (N_819,In_1485,In_391);
or U820 (N_820,In_1677,In_394);
or U821 (N_821,In_2097,In_854);
nand U822 (N_822,In_413,In_2395);
nor U823 (N_823,In_48,In_481);
and U824 (N_824,In_2061,In_2183);
or U825 (N_825,In_1016,In_791);
nand U826 (N_826,In_2375,In_1438);
nor U827 (N_827,In_2401,In_187);
or U828 (N_828,In_880,In_385);
nor U829 (N_829,In_513,In_2350);
nand U830 (N_830,In_2322,In_2359);
nor U831 (N_831,In_2055,In_2087);
or U832 (N_832,In_1657,In_894);
or U833 (N_833,In_2007,In_1532);
xnor U834 (N_834,In_2334,In_2201);
or U835 (N_835,In_1134,In_638);
and U836 (N_836,In_1688,In_1873);
xnor U837 (N_837,In_131,In_1126);
nand U838 (N_838,In_1474,In_1584);
or U839 (N_839,In_1951,In_680);
and U840 (N_840,In_2450,In_670);
nand U841 (N_841,In_200,In_2207);
nor U842 (N_842,In_241,In_2122);
nand U843 (N_843,In_2459,In_1812);
or U844 (N_844,In_610,In_866);
nor U845 (N_845,In_363,In_1244);
or U846 (N_846,In_1590,In_2447);
or U847 (N_847,In_660,In_611);
nor U848 (N_848,In_445,In_126);
xnor U849 (N_849,In_783,In_484);
or U850 (N_850,In_627,In_1201);
nor U851 (N_851,In_1615,In_405);
or U852 (N_852,In_912,In_932);
xnor U853 (N_853,In_2443,In_800);
or U854 (N_854,In_1852,In_1870);
nor U855 (N_855,In_1148,In_869);
and U856 (N_856,In_530,In_1702);
or U857 (N_857,In_1073,In_28);
nand U858 (N_858,In_1024,In_466);
xnor U859 (N_859,In_2129,In_1416);
and U860 (N_860,In_198,In_528);
nor U861 (N_861,In_689,In_170);
xor U862 (N_862,In_1940,In_1247);
or U863 (N_863,In_1686,In_2250);
nor U864 (N_864,In_337,In_165);
or U865 (N_865,In_664,In_2022);
or U866 (N_866,In_1938,In_1654);
nor U867 (N_867,In_483,In_831);
and U868 (N_868,In_1928,In_109);
nand U869 (N_869,In_940,In_968);
nand U870 (N_870,In_1137,In_1756);
nor U871 (N_871,In_1655,In_1530);
nor U872 (N_872,In_97,In_1037);
or U873 (N_873,In_2044,In_764);
and U874 (N_874,In_716,In_1790);
and U875 (N_875,In_2264,In_400);
nand U876 (N_876,In_585,In_1860);
and U877 (N_877,In_752,In_2073);
or U878 (N_878,In_2480,In_1412);
nor U879 (N_879,In_214,In_1796);
nor U880 (N_880,In_930,In_1288);
nor U881 (N_881,In_1383,In_1299);
nand U882 (N_882,In_162,In_2164);
nand U883 (N_883,In_2464,In_1337);
nor U884 (N_884,In_1695,In_2156);
nor U885 (N_885,In_2392,In_465);
nor U886 (N_886,In_2173,In_1599);
and U887 (N_887,In_1776,In_1946);
nor U888 (N_888,In_1723,In_2056);
xnor U889 (N_889,In_565,In_1489);
and U890 (N_890,In_1048,In_2274);
nand U891 (N_891,In_1739,In_580);
nand U892 (N_892,In_1301,In_1342);
nand U893 (N_893,In_1706,In_2252);
nand U894 (N_894,In_2057,In_29);
and U895 (N_895,In_1548,In_2270);
nand U896 (N_896,In_705,In_2469);
nand U897 (N_897,In_2394,In_2178);
and U898 (N_898,In_1847,In_2346);
nand U899 (N_899,In_1223,In_1604);
nor U900 (N_900,In_536,In_1313);
nand U901 (N_901,In_2373,In_1623);
nand U902 (N_902,In_1818,In_1395);
nand U903 (N_903,In_629,In_1049);
or U904 (N_904,In_2366,In_1786);
nand U905 (N_905,In_830,In_74);
and U906 (N_906,In_382,In_281);
nor U907 (N_907,In_683,In_291);
xnor U908 (N_908,In_1619,In_1050);
or U909 (N_909,In_790,In_1092);
xor U910 (N_910,In_2198,In_881);
or U911 (N_911,In_859,In_826);
xnor U912 (N_912,In_1069,In_207);
and U913 (N_913,In_2418,In_424);
nand U914 (N_914,In_1409,In_1461);
or U915 (N_915,In_2218,In_985);
or U916 (N_916,In_305,In_976);
nand U917 (N_917,In_573,In_1188);
nand U918 (N_918,In_1022,In_1045);
nand U919 (N_919,In_70,In_1967);
and U920 (N_920,In_2131,In_2199);
and U921 (N_921,In_2177,In_1149);
and U922 (N_922,In_0,In_1355);
nor U923 (N_923,In_1486,In_988);
nand U924 (N_924,In_843,In_552);
nor U925 (N_925,In_730,In_2466);
and U926 (N_926,In_574,In_231);
or U927 (N_927,In_384,In_2092);
or U928 (N_928,In_2051,In_1457);
nand U929 (N_929,In_699,In_1155);
nor U930 (N_930,In_1061,In_898);
and U931 (N_931,In_2118,In_1070);
nor U932 (N_932,In_1593,In_427);
nor U933 (N_933,In_639,In_218);
nor U934 (N_934,In_2163,In_1692);
nor U935 (N_935,In_1865,In_461);
nand U936 (N_936,In_1322,In_2130);
nor U937 (N_937,In_485,In_2187);
or U938 (N_938,In_601,In_1522);
or U939 (N_939,In_1722,In_100);
nor U940 (N_940,In_1278,In_1925);
or U941 (N_941,In_1468,In_63);
and U942 (N_942,In_891,In_2176);
nand U943 (N_943,In_1487,In_1484);
nor U944 (N_944,In_2387,In_2047);
and U945 (N_945,In_1935,In_2112);
and U946 (N_946,In_1154,In_2185);
or U947 (N_947,In_1621,In_2067);
nand U948 (N_948,In_1665,In_2141);
and U949 (N_949,In_531,In_1267);
and U950 (N_950,In_1005,In_1704);
xnor U951 (N_951,In_56,In_1572);
or U952 (N_952,In_1493,In_1115);
and U953 (N_953,In_655,In_380);
xor U954 (N_954,In_2149,In_2155);
or U955 (N_955,In_1934,In_1979);
nand U956 (N_956,In_204,In_173);
nor U957 (N_957,In_636,In_219);
nand U958 (N_958,In_2029,In_243);
nand U959 (N_959,In_1973,In_1526);
nand U960 (N_960,In_799,In_188);
nor U961 (N_961,In_1827,In_620);
nor U962 (N_962,In_2228,In_1777);
and U963 (N_963,In_111,In_1799);
nor U964 (N_964,In_1800,In_1816);
and U965 (N_965,In_561,In_646);
nor U966 (N_966,In_1213,In_935);
nand U967 (N_967,In_1580,In_598);
or U968 (N_968,In_1803,In_1725);
nand U969 (N_969,In_819,In_647);
nand U970 (N_970,In_1830,In_50);
nand U971 (N_971,In_1451,In_765);
or U972 (N_972,In_2327,In_944);
nor U973 (N_973,In_2492,In_1917);
or U974 (N_974,In_2005,In_1854);
nand U975 (N_975,In_1118,In_152);
and U976 (N_976,In_868,In_172);
or U977 (N_977,In_1581,In_1683);
and U978 (N_978,In_537,In_775);
nand U979 (N_979,In_1586,In_1123);
nor U980 (N_980,In_1376,In_2410);
nand U981 (N_981,In_1192,In_1923);
or U982 (N_982,In_107,In_1890);
nor U983 (N_983,In_1958,In_1687);
nor U984 (N_984,In_2340,In_1825);
xnor U985 (N_985,In_1696,In_1924);
nand U986 (N_986,In_92,In_523);
nor U987 (N_987,In_538,In_1242);
xor U988 (N_988,In_2142,In_1603);
xnor U989 (N_989,In_1413,In_1275);
nor U990 (N_990,In_1547,In_2399);
nor U991 (N_991,In_153,In_1516);
nor U992 (N_992,In_437,In_2117);
nor U993 (N_993,In_576,In_899);
and U994 (N_994,In_171,In_495);
and U995 (N_995,In_1145,In_2458);
and U996 (N_996,In_62,In_226);
nand U997 (N_997,In_919,In_1659);
and U998 (N_998,In_556,In_614);
and U999 (N_999,In_2189,In_1901);
and U1000 (N_1000,In_2078,In_350);
and U1001 (N_1001,In_2455,In_1788);
and U1002 (N_1002,In_717,In_1864);
nand U1003 (N_1003,In_2400,In_1612);
nand U1004 (N_1004,In_1308,In_1285);
and U1005 (N_1005,In_2203,In_602);
nand U1006 (N_1006,In_1231,In_1375);
xnor U1007 (N_1007,In_771,In_239);
nand U1008 (N_1008,In_1455,In_657);
and U1009 (N_1009,In_144,In_1577);
nor U1010 (N_1010,In_1382,In_1999);
nand U1011 (N_1011,In_2435,In_1333);
and U1012 (N_1012,In_2015,In_2310);
or U1013 (N_1013,In_2070,In_1836);
and U1014 (N_1014,In_2100,In_2039);
or U1015 (N_1015,In_1346,In_302);
nand U1016 (N_1016,In_1913,In_1450);
nor U1017 (N_1017,In_315,In_2370);
nand U1018 (N_1018,In_355,In_1314);
nor U1019 (N_1019,In_261,In_1388);
and U1020 (N_1020,In_356,In_1206);
and U1021 (N_1021,In_1100,In_343);
and U1022 (N_1022,In_567,In_1347);
nor U1023 (N_1023,In_1297,In_9);
nand U1024 (N_1024,In_12,In_1682);
nor U1025 (N_1025,In_2138,In_176);
nor U1026 (N_1026,In_2307,In_304);
or U1027 (N_1027,In_1043,In_963);
and U1028 (N_1028,In_1392,In_211);
and U1029 (N_1029,In_1556,In_719);
nor U1030 (N_1030,In_159,In_1373);
nand U1031 (N_1031,In_1791,In_264);
nand U1032 (N_1032,In_974,In_2236);
nand U1033 (N_1033,In_555,In_1436);
or U1034 (N_1034,In_1717,In_832);
and U1035 (N_1035,In_2066,In_1883);
nand U1036 (N_1036,In_1916,In_1046);
nand U1037 (N_1037,In_545,In_2175);
or U1038 (N_1038,In_10,In_1525);
or U1039 (N_1039,In_645,In_301);
nand U1040 (N_1040,In_2498,In_298);
nand U1041 (N_1041,In_429,In_942);
nand U1042 (N_1042,In_550,In_1481);
and U1043 (N_1043,In_1961,In_395);
and U1044 (N_1044,In_1751,In_1898);
or U1045 (N_1045,In_1959,In_196);
nor U1046 (N_1046,In_2208,In_1568);
nor U1047 (N_1047,In_425,In_1998);
or U1048 (N_1048,In_973,In_2267);
or U1049 (N_1049,In_2225,In_2437);
xnor U1050 (N_1050,In_922,In_1303);
nand U1051 (N_1051,In_1817,In_2438);
nand U1052 (N_1052,In_798,In_649);
nand U1053 (N_1053,In_671,In_1970);
or U1054 (N_1054,In_191,In_2023);
and U1055 (N_1055,In_822,In_861);
or U1056 (N_1056,In_1670,In_145);
nor U1057 (N_1057,In_511,In_365);
nand U1058 (N_1058,In_94,In_1411);
xor U1059 (N_1059,In_1162,In_1165);
xor U1060 (N_1060,In_818,In_2076);
or U1061 (N_1061,In_1135,In_570);
nand U1062 (N_1062,In_27,In_2038);
nor U1063 (N_1063,In_1008,In_235);
nand U1064 (N_1064,In_2494,In_1014);
nand U1065 (N_1065,In_17,In_417);
or U1066 (N_1066,In_2169,In_753);
and U1067 (N_1067,In_760,In_108);
nand U1068 (N_1068,In_2255,In_2246);
xnor U1069 (N_1069,In_1719,In_2354);
nand U1070 (N_1070,In_1251,In_474);
nor U1071 (N_1071,In_1611,In_2318);
nor U1072 (N_1072,In_1002,In_155);
nand U1073 (N_1073,In_1806,In_2313);
or U1074 (N_1074,In_2338,In_2485);
xnor U1075 (N_1075,In_1209,In_1878);
nand U1076 (N_1076,In_1327,In_339);
nand U1077 (N_1077,In_1083,In_1435);
nand U1078 (N_1078,In_558,In_2386);
and U1079 (N_1079,In_1859,In_1216);
nor U1080 (N_1080,In_300,In_1125);
nand U1081 (N_1081,In_2369,In_283);
or U1082 (N_1082,In_2384,In_388);
xor U1083 (N_1083,In_1035,In_1848);
nand U1084 (N_1084,In_1252,In_303);
nor U1085 (N_1085,In_2210,In_994);
nand U1086 (N_1086,In_104,In_1000);
nand U1087 (N_1087,In_26,In_1284);
nand U1088 (N_1088,In_518,In_1054);
or U1089 (N_1089,In_1537,In_1068);
or U1090 (N_1090,In_2140,In_2089);
nand U1091 (N_1091,In_240,In_259);
nor U1092 (N_1092,In_2289,In_1947);
nand U1093 (N_1093,In_811,In_1030);
nor U1094 (N_1094,In_1051,In_2421);
nor U1095 (N_1095,In_96,In_1563);
and U1096 (N_1096,In_2085,In_964);
and U1097 (N_1097,In_79,In_681);
and U1098 (N_1098,In_245,In_1514);
and U1099 (N_1099,In_1270,In_2445);
nor U1100 (N_1100,In_255,In_1613);
nand U1101 (N_1101,In_168,In_746);
and U1102 (N_1102,In_673,In_858);
xnor U1103 (N_1103,In_566,In_2385);
nand U1104 (N_1104,In_1761,In_1415);
nor U1105 (N_1105,In_1769,In_592);
and U1106 (N_1106,In_1410,In_2064);
nor U1107 (N_1107,In_1317,In_140);
and U1108 (N_1108,In_612,In_216);
and U1109 (N_1109,In_1555,In_225);
nand U1110 (N_1110,In_672,In_2098);
or U1111 (N_1111,In_984,In_1996);
or U1112 (N_1112,In_1352,In_2324);
and U1113 (N_1113,In_422,In_987);
nor U1114 (N_1114,In_446,In_686);
or U1115 (N_1115,In_1079,In_249);
nor U1116 (N_1116,In_1622,In_1289);
nand U1117 (N_1117,In_1062,In_192);
and U1118 (N_1118,In_357,In_1007);
nand U1119 (N_1119,In_997,In_280);
nor U1120 (N_1120,In_1038,In_35);
and U1121 (N_1121,In_1138,In_702);
nor U1122 (N_1122,In_1108,In_157);
or U1123 (N_1123,In_1679,In_1962);
nand U1124 (N_1124,In_578,In_844);
and U1125 (N_1125,In_2442,In_1538);
nand U1126 (N_1126,In_723,In_971);
or U1127 (N_1127,In_1106,In_862);
xnor U1128 (N_1128,In_1442,In_2043);
xor U1129 (N_1129,In_8,In_39);
and U1130 (N_1130,In_1519,In_1711);
nor U1131 (N_1131,In_354,In_887);
nand U1132 (N_1132,In_907,In_430);
nor U1133 (N_1133,In_562,In_1331);
or U1134 (N_1134,In_871,In_503);
and U1135 (N_1135,In_1338,In_2195);
or U1136 (N_1136,In_575,In_579);
or U1137 (N_1137,In_115,In_1974);
xnor U1138 (N_1138,In_2308,In_1771);
or U1139 (N_1139,In_885,In_2063);
nand U1140 (N_1140,In_1645,In_1506);
nand U1141 (N_1141,In_1490,In_1396);
and U1142 (N_1142,In_635,In_807);
nor U1143 (N_1143,In_1257,In_1107);
or U1144 (N_1144,In_2127,In_1076);
xor U1145 (N_1145,In_712,In_2139);
and U1146 (N_1146,In_1113,In_326);
nand U1147 (N_1147,In_978,In_266);
nand U1148 (N_1148,In_1328,In_543);
or U1149 (N_1149,In_2053,In_1434);
or U1150 (N_1150,In_1638,In_2448);
nand U1151 (N_1151,In_1429,In_920);
nor U1152 (N_1152,In_1871,In_452);
or U1153 (N_1153,In_2368,In_447);
and U1154 (N_1154,In_221,In_2211);
and U1155 (N_1155,In_2460,In_1173);
nand U1156 (N_1156,In_2456,In_1310);
or U1157 (N_1157,In_781,In_589);
or U1158 (N_1158,In_379,In_663);
and U1159 (N_1159,In_387,In_1478);
xor U1160 (N_1160,In_633,In_1087);
xnor U1161 (N_1161,In_1379,In_2451);
and U1162 (N_1162,In_2105,In_2453);
or U1163 (N_1163,In_2216,In_1402);
nand U1164 (N_1164,In_835,In_946);
or U1165 (N_1165,In_2214,In_1726);
or U1166 (N_1166,In_1056,In_421);
or U1167 (N_1167,In_2018,In_792);
nand U1168 (N_1168,In_233,In_651);
and U1169 (N_1169,In_389,In_1714);
or U1170 (N_1170,In_201,In_1663);
or U1171 (N_1171,In_1573,In_331);
nor U1172 (N_1172,In_2325,In_2006);
and U1173 (N_1173,In_1241,In_2021);
and U1174 (N_1174,In_1421,In_1101);
and U1175 (N_1175,In_1139,In_721);
nor U1176 (N_1176,In_458,In_2091);
or U1177 (N_1177,In_117,In_2205);
and U1178 (N_1178,In_1321,In_770);
nor U1179 (N_1179,In_2268,In_1013);
nor U1180 (N_1180,In_1131,In_804);
or U1181 (N_1181,In_1760,In_1838);
nand U1182 (N_1182,In_1104,In_1207);
nand U1183 (N_1183,In_519,In_857);
nand U1184 (N_1184,In_911,In_2008);
xnor U1185 (N_1185,In_2045,In_14);
or U1186 (N_1186,In_2269,In_1826);
or U1187 (N_1187,In_1172,In_127);
or U1188 (N_1188,In_1993,In_1260);
nand U1189 (N_1189,In_751,In_1772);
nor U1190 (N_1190,In_1542,In_308);
or U1191 (N_1191,In_1983,In_2235);
or U1192 (N_1192,In_1876,In_2186);
nand U1193 (N_1193,In_904,In_959);
nand U1194 (N_1194,In_1820,In_1214);
or U1195 (N_1195,In_2107,In_652);
and U1196 (N_1196,In_2470,In_1105);
or U1197 (N_1197,In_1147,In_1784);
nor U1198 (N_1198,In_285,In_1552);
nand U1199 (N_1199,In_2488,In_801);
nor U1200 (N_1200,In_2475,In_1283);
nor U1201 (N_1201,In_414,In_909);
and U1202 (N_1202,In_2279,In_428);
or U1203 (N_1203,In_367,In_828);
nand U1204 (N_1204,In_1787,In_1171);
nor U1205 (N_1205,In_1965,In_2082);
or U1206 (N_1206,In_2412,In_1509);
or U1207 (N_1207,In_1606,In_1028);
nor U1208 (N_1208,In_463,In_867);
and U1209 (N_1209,In_1181,In_1298);
or U1210 (N_1210,In_136,In_2411);
nor U1211 (N_1211,In_1539,In_1253);
or U1212 (N_1212,In_879,In_2024);
and U1213 (N_1213,In_2077,In_1433);
nand U1214 (N_1214,In_1483,In_1738);
and U1215 (N_1215,In_1203,In_1185);
nand U1216 (N_1216,In_691,In_740);
nand U1217 (N_1217,In_1668,In_659);
nand U1218 (N_1218,In_797,In_2037);
nor U1219 (N_1219,In_1789,In_1473);
or U1220 (N_1220,In_970,In_1094);
or U1221 (N_1221,In_1479,In_2388);
or U1222 (N_1222,In_2349,In_1066);
and U1223 (N_1223,In_492,In_436);
and U1224 (N_1224,In_1237,In_268);
and U1225 (N_1225,In_21,In_334);
nand U1226 (N_1226,In_2348,In_1987);
nor U1227 (N_1227,In_877,In_2237);
nand U1228 (N_1228,In_113,In_768);
nor U1229 (N_1229,In_2377,In_829);
and U1230 (N_1230,In_802,In_560);
nand U1231 (N_1231,In_632,In_1693);
and U1232 (N_1232,In_1184,In_72);
and U1233 (N_1233,In_65,In_2166);
or U1234 (N_1234,In_733,In_1550);
or U1235 (N_1235,In_1443,In_2405);
nand U1236 (N_1236,In_2287,In_1177);
or U1237 (N_1237,In_78,In_989);
and U1238 (N_1238,In_1405,In_1955);
nor U1239 (N_1239,In_1533,In_1906);
nor U1240 (N_1240,In_1111,In_737);
nor U1241 (N_1241,In_1741,In_2407);
and U1242 (N_1242,In_1758,In_182);
and U1243 (N_1243,In_1282,In_1699);
nor U1244 (N_1244,In_1053,In_834);
nand U1245 (N_1245,In_371,In_735);
or U1246 (N_1246,In_412,In_995);
nand U1247 (N_1247,In_498,In_1626);
nor U1248 (N_1248,In_497,In_290);
or U1249 (N_1249,In_1098,In_1844);
and U1250 (N_1250,In_1395,In_1166);
nand U1251 (N_1251,In_1169,In_109);
nor U1252 (N_1252,In_2479,In_63);
nor U1253 (N_1253,In_2079,In_1246);
and U1254 (N_1254,In_1181,In_861);
and U1255 (N_1255,In_740,In_1073);
and U1256 (N_1256,In_1571,In_2499);
nor U1257 (N_1257,In_2419,In_362);
or U1258 (N_1258,In_94,In_1591);
or U1259 (N_1259,In_360,In_1137);
xor U1260 (N_1260,In_1587,In_1211);
nand U1261 (N_1261,In_2115,In_1537);
nand U1262 (N_1262,In_2099,In_406);
xor U1263 (N_1263,In_1608,In_1345);
or U1264 (N_1264,In_1177,In_106);
nor U1265 (N_1265,In_2256,In_51);
nand U1266 (N_1266,In_2119,In_1701);
nand U1267 (N_1267,In_503,In_1556);
nand U1268 (N_1268,In_818,In_1230);
nand U1269 (N_1269,In_666,In_2115);
xor U1270 (N_1270,In_1889,In_2428);
nor U1271 (N_1271,In_739,In_1796);
xor U1272 (N_1272,In_1525,In_1190);
or U1273 (N_1273,In_489,In_1212);
nand U1274 (N_1274,In_1246,In_995);
nand U1275 (N_1275,In_2414,In_472);
nor U1276 (N_1276,In_921,In_527);
nor U1277 (N_1277,In_1739,In_2051);
and U1278 (N_1278,In_1643,In_1278);
and U1279 (N_1279,In_465,In_2131);
or U1280 (N_1280,In_2118,In_646);
and U1281 (N_1281,In_2464,In_2344);
or U1282 (N_1282,In_630,In_1662);
nand U1283 (N_1283,In_1358,In_1599);
and U1284 (N_1284,In_1286,In_1172);
nor U1285 (N_1285,In_425,In_1563);
or U1286 (N_1286,In_143,In_1836);
nand U1287 (N_1287,In_2152,In_1237);
nor U1288 (N_1288,In_1542,In_387);
or U1289 (N_1289,In_1746,In_840);
xor U1290 (N_1290,In_1350,In_653);
nand U1291 (N_1291,In_873,In_240);
nand U1292 (N_1292,In_1985,In_456);
nand U1293 (N_1293,In_837,In_1342);
and U1294 (N_1294,In_936,In_1177);
or U1295 (N_1295,In_2218,In_446);
or U1296 (N_1296,In_1518,In_592);
nor U1297 (N_1297,In_830,In_2099);
xor U1298 (N_1298,In_1533,In_2175);
nor U1299 (N_1299,In_1168,In_1740);
or U1300 (N_1300,In_1282,In_1755);
or U1301 (N_1301,In_58,In_340);
nor U1302 (N_1302,In_502,In_2484);
or U1303 (N_1303,In_445,In_888);
nand U1304 (N_1304,In_1402,In_2284);
or U1305 (N_1305,In_1702,In_701);
or U1306 (N_1306,In_1506,In_563);
nand U1307 (N_1307,In_427,In_2317);
and U1308 (N_1308,In_1125,In_1903);
nand U1309 (N_1309,In_505,In_1775);
or U1310 (N_1310,In_1631,In_701);
nor U1311 (N_1311,In_611,In_1695);
nand U1312 (N_1312,In_371,In_1249);
or U1313 (N_1313,In_133,In_2184);
nand U1314 (N_1314,In_2114,In_1086);
xor U1315 (N_1315,In_2164,In_1401);
and U1316 (N_1316,In_990,In_96);
nor U1317 (N_1317,In_1935,In_981);
or U1318 (N_1318,In_133,In_2422);
and U1319 (N_1319,In_1836,In_1627);
nor U1320 (N_1320,In_1635,In_2477);
nor U1321 (N_1321,In_1169,In_907);
xor U1322 (N_1322,In_457,In_885);
or U1323 (N_1323,In_652,In_1933);
or U1324 (N_1324,In_1846,In_2238);
and U1325 (N_1325,In_1844,In_1508);
nand U1326 (N_1326,In_1793,In_2496);
nand U1327 (N_1327,In_2420,In_2478);
nor U1328 (N_1328,In_169,In_1900);
nor U1329 (N_1329,In_1698,In_292);
or U1330 (N_1330,In_2025,In_343);
nand U1331 (N_1331,In_1776,In_262);
xnor U1332 (N_1332,In_311,In_1963);
xor U1333 (N_1333,In_2290,In_2164);
or U1334 (N_1334,In_1868,In_43);
and U1335 (N_1335,In_2218,In_1157);
and U1336 (N_1336,In_1378,In_36);
nand U1337 (N_1337,In_1334,In_1581);
and U1338 (N_1338,In_374,In_654);
nand U1339 (N_1339,In_245,In_2478);
nor U1340 (N_1340,In_736,In_1386);
and U1341 (N_1341,In_582,In_2312);
or U1342 (N_1342,In_1047,In_1130);
and U1343 (N_1343,In_2183,In_247);
nor U1344 (N_1344,In_1325,In_2022);
and U1345 (N_1345,In_1330,In_459);
nor U1346 (N_1346,In_840,In_1147);
xor U1347 (N_1347,In_2195,In_989);
or U1348 (N_1348,In_940,In_742);
nand U1349 (N_1349,In_2375,In_538);
or U1350 (N_1350,In_488,In_607);
or U1351 (N_1351,In_2121,In_414);
nand U1352 (N_1352,In_2016,In_1513);
or U1353 (N_1353,In_1114,In_1990);
or U1354 (N_1354,In_1244,In_2293);
nor U1355 (N_1355,In_1957,In_106);
and U1356 (N_1356,In_1132,In_997);
and U1357 (N_1357,In_1782,In_798);
and U1358 (N_1358,In_923,In_1036);
and U1359 (N_1359,In_150,In_175);
or U1360 (N_1360,In_437,In_895);
nand U1361 (N_1361,In_842,In_470);
and U1362 (N_1362,In_2232,In_1312);
nor U1363 (N_1363,In_476,In_1245);
xnor U1364 (N_1364,In_479,In_2019);
and U1365 (N_1365,In_982,In_913);
xor U1366 (N_1366,In_2438,In_2257);
xor U1367 (N_1367,In_831,In_101);
or U1368 (N_1368,In_1807,In_433);
nand U1369 (N_1369,In_27,In_952);
and U1370 (N_1370,In_1082,In_1632);
nand U1371 (N_1371,In_2494,In_68);
nor U1372 (N_1372,In_395,In_916);
nor U1373 (N_1373,In_941,In_2146);
or U1374 (N_1374,In_2204,In_882);
nor U1375 (N_1375,In_646,In_2023);
nor U1376 (N_1376,In_1416,In_604);
or U1377 (N_1377,In_433,In_1994);
xnor U1378 (N_1378,In_2320,In_2250);
and U1379 (N_1379,In_1159,In_441);
nand U1380 (N_1380,In_473,In_2043);
or U1381 (N_1381,In_1449,In_2443);
and U1382 (N_1382,In_470,In_600);
or U1383 (N_1383,In_1270,In_1571);
or U1384 (N_1384,In_2337,In_767);
nor U1385 (N_1385,In_1509,In_331);
or U1386 (N_1386,In_1647,In_477);
or U1387 (N_1387,In_22,In_2394);
or U1388 (N_1388,In_165,In_1979);
and U1389 (N_1389,In_2192,In_2066);
nand U1390 (N_1390,In_1932,In_661);
nor U1391 (N_1391,In_320,In_1678);
nor U1392 (N_1392,In_465,In_1802);
nand U1393 (N_1393,In_2053,In_1342);
xor U1394 (N_1394,In_506,In_1189);
nor U1395 (N_1395,In_1970,In_789);
and U1396 (N_1396,In_2078,In_2056);
nand U1397 (N_1397,In_2173,In_1792);
and U1398 (N_1398,In_1486,In_1740);
nor U1399 (N_1399,In_2144,In_414);
or U1400 (N_1400,In_1219,In_2161);
or U1401 (N_1401,In_193,In_618);
nand U1402 (N_1402,In_366,In_66);
nor U1403 (N_1403,In_1682,In_2304);
or U1404 (N_1404,In_1605,In_2000);
or U1405 (N_1405,In_2325,In_2033);
nor U1406 (N_1406,In_2418,In_1377);
or U1407 (N_1407,In_185,In_329);
or U1408 (N_1408,In_1151,In_1575);
nor U1409 (N_1409,In_1766,In_108);
and U1410 (N_1410,In_741,In_293);
and U1411 (N_1411,In_426,In_1491);
nand U1412 (N_1412,In_2174,In_1973);
nand U1413 (N_1413,In_2029,In_793);
and U1414 (N_1414,In_1543,In_831);
nand U1415 (N_1415,In_1247,In_1177);
nand U1416 (N_1416,In_1479,In_1512);
or U1417 (N_1417,In_2099,In_2104);
nand U1418 (N_1418,In_1188,In_2139);
or U1419 (N_1419,In_1552,In_1994);
nand U1420 (N_1420,In_1590,In_1476);
and U1421 (N_1421,In_450,In_1275);
and U1422 (N_1422,In_1228,In_336);
xor U1423 (N_1423,In_2149,In_988);
or U1424 (N_1424,In_559,In_1026);
nor U1425 (N_1425,In_214,In_295);
nand U1426 (N_1426,In_268,In_600);
and U1427 (N_1427,In_1342,In_156);
xor U1428 (N_1428,In_185,In_2226);
xnor U1429 (N_1429,In_787,In_1452);
xor U1430 (N_1430,In_789,In_744);
xnor U1431 (N_1431,In_218,In_1746);
nor U1432 (N_1432,In_1541,In_1046);
or U1433 (N_1433,In_1559,In_199);
nand U1434 (N_1434,In_1328,In_898);
nand U1435 (N_1435,In_67,In_187);
nand U1436 (N_1436,In_191,In_617);
nor U1437 (N_1437,In_744,In_142);
xor U1438 (N_1438,In_1776,In_165);
and U1439 (N_1439,In_1087,In_315);
nor U1440 (N_1440,In_1216,In_871);
nand U1441 (N_1441,In_1008,In_795);
or U1442 (N_1442,In_1996,In_175);
and U1443 (N_1443,In_2102,In_721);
and U1444 (N_1444,In_2337,In_27);
and U1445 (N_1445,In_618,In_2048);
nor U1446 (N_1446,In_2055,In_758);
nand U1447 (N_1447,In_1136,In_1894);
nor U1448 (N_1448,In_1765,In_2374);
or U1449 (N_1449,In_469,In_1184);
and U1450 (N_1450,In_267,In_1135);
or U1451 (N_1451,In_229,In_511);
nor U1452 (N_1452,In_1925,In_585);
and U1453 (N_1453,In_441,In_246);
nand U1454 (N_1454,In_1973,In_1036);
xor U1455 (N_1455,In_1038,In_364);
nand U1456 (N_1456,In_86,In_2110);
nand U1457 (N_1457,In_2163,In_1976);
nand U1458 (N_1458,In_1411,In_1372);
nand U1459 (N_1459,In_814,In_1039);
or U1460 (N_1460,In_1240,In_1481);
xnor U1461 (N_1461,In_1675,In_1563);
nor U1462 (N_1462,In_237,In_321);
nand U1463 (N_1463,In_356,In_1938);
xnor U1464 (N_1464,In_21,In_1407);
or U1465 (N_1465,In_1035,In_2140);
or U1466 (N_1466,In_1360,In_625);
and U1467 (N_1467,In_1195,In_1791);
or U1468 (N_1468,In_2019,In_1251);
xnor U1469 (N_1469,In_1403,In_1018);
or U1470 (N_1470,In_1155,In_1909);
xor U1471 (N_1471,In_87,In_405);
nand U1472 (N_1472,In_1751,In_1378);
nand U1473 (N_1473,In_1466,In_376);
nand U1474 (N_1474,In_2326,In_203);
and U1475 (N_1475,In_1041,In_2437);
nor U1476 (N_1476,In_604,In_2335);
or U1477 (N_1477,In_1135,In_2250);
or U1478 (N_1478,In_2442,In_1561);
xor U1479 (N_1479,In_91,In_665);
or U1480 (N_1480,In_438,In_1429);
nor U1481 (N_1481,In_2259,In_1556);
nor U1482 (N_1482,In_1282,In_1989);
and U1483 (N_1483,In_2419,In_196);
and U1484 (N_1484,In_2203,In_321);
or U1485 (N_1485,In_105,In_2491);
nor U1486 (N_1486,In_1209,In_2454);
or U1487 (N_1487,In_1066,In_1747);
nor U1488 (N_1488,In_2010,In_1473);
and U1489 (N_1489,In_2449,In_2137);
xor U1490 (N_1490,In_881,In_2245);
or U1491 (N_1491,In_1322,In_1806);
nor U1492 (N_1492,In_532,In_1372);
and U1493 (N_1493,In_1386,In_2387);
or U1494 (N_1494,In_1296,In_778);
xor U1495 (N_1495,In_2122,In_1212);
nor U1496 (N_1496,In_607,In_546);
xnor U1497 (N_1497,In_1832,In_1671);
nor U1498 (N_1498,In_2105,In_592);
xor U1499 (N_1499,In_1610,In_670);
and U1500 (N_1500,In_316,In_1078);
or U1501 (N_1501,In_786,In_712);
and U1502 (N_1502,In_1425,In_2289);
or U1503 (N_1503,In_432,In_761);
nand U1504 (N_1504,In_103,In_1475);
or U1505 (N_1505,In_1244,In_12);
nand U1506 (N_1506,In_200,In_1695);
nand U1507 (N_1507,In_514,In_957);
or U1508 (N_1508,In_449,In_17);
nor U1509 (N_1509,In_1402,In_774);
nor U1510 (N_1510,In_135,In_27);
or U1511 (N_1511,In_110,In_731);
nand U1512 (N_1512,In_868,In_1273);
nor U1513 (N_1513,In_2351,In_879);
and U1514 (N_1514,In_2295,In_2086);
and U1515 (N_1515,In_1810,In_1956);
or U1516 (N_1516,In_241,In_2109);
or U1517 (N_1517,In_1784,In_360);
nor U1518 (N_1518,In_201,In_1408);
nor U1519 (N_1519,In_1119,In_480);
nor U1520 (N_1520,In_198,In_409);
or U1521 (N_1521,In_519,In_1135);
nor U1522 (N_1522,In_180,In_749);
or U1523 (N_1523,In_646,In_2043);
xor U1524 (N_1524,In_1567,In_204);
nor U1525 (N_1525,In_505,In_676);
nand U1526 (N_1526,In_679,In_1837);
nand U1527 (N_1527,In_2050,In_331);
nor U1528 (N_1528,In_704,In_2095);
xor U1529 (N_1529,In_2392,In_1767);
and U1530 (N_1530,In_1542,In_482);
nor U1531 (N_1531,In_1899,In_121);
or U1532 (N_1532,In_60,In_2034);
nor U1533 (N_1533,In_1372,In_221);
and U1534 (N_1534,In_182,In_2212);
and U1535 (N_1535,In_1111,In_531);
and U1536 (N_1536,In_368,In_317);
nand U1537 (N_1537,In_2014,In_1056);
nor U1538 (N_1538,In_2400,In_2362);
or U1539 (N_1539,In_396,In_2140);
nor U1540 (N_1540,In_1063,In_374);
nand U1541 (N_1541,In_2398,In_1469);
xor U1542 (N_1542,In_2431,In_2333);
nand U1543 (N_1543,In_2139,In_2303);
nand U1544 (N_1544,In_2464,In_169);
and U1545 (N_1545,In_433,In_625);
xor U1546 (N_1546,In_2313,In_389);
or U1547 (N_1547,In_1818,In_694);
nor U1548 (N_1548,In_1893,In_2119);
and U1549 (N_1549,In_155,In_2046);
or U1550 (N_1550,In_447,In_2100);
nor U1551 (N_1551,In_1831,In_2091);
or U1552 (N_1552,In_427,In_585);
or U1553 (N_1553,In_721,In_68);
nand U1554 (N_1554,In_446,In_2334);
and U1555 (N_1555,In_2224,In_698);
or U1556 (N_1556,In_1863,In_857);
nor U1557 (N_1557,In_2395,In_1633);
and U1558 (N_1558,In_2341,In_2461);
or U1559 (N_1559,In_127,In_1272);
nand U1560 (N_1560,In_2182,In_1463);
nor U1561 (N_1561,In_1601,In_146);
or U1562 (N_1562,In_2121,In_1789);
or U1563 (N_1563,In_1377,In_2130);
or U1564 (N_1564,In_60,In_2208);
or U1565 (N_1565,In_2356,In_2472);
or U1566 (N_1566,In_355,In_305);
and U1567 (N_1567,In_165,In_595);
nor U1568 (N_1568,In_832,In_1246);
or U1569 (N_1569,In_2311,In_0);
and U1570 (N_1570,In_700,In_1290);
or U1571 (N_1571,In_142,In_1776);
nand U1572 (N_1572,In_776,In_2470);
or U1573 (N_1573,In_171,In_3);
nor U1574 (N_1574,In_1848,In_2143);
or U1575 (N_1575,In_2080,In_2184);
or U1576 (N_1576,In_1970,In_2470);
xor U1577 (N_1577,In_508,In_1118);
or U1578 (N_1578,In_131,In_1297);
xor U1579 (N_1579,In_543,In_836);
or U1580 (N_1580,In_1162,In_1497);
or U1581 (N_1581,In_2411,In_257);
or U1582 (N_1582,In_1289,In_1244);
nor U1583 (N_1583,In_1673,In_1431);
and U1584 (N_1584,In_1048,In_406);
or U1585 (N_1585,In_348,In_1797);
nand U1586 (N_1586,In_626,In_1445);
and U1587 (N_1587,In_110,In_275);
nand U1588 (N_1588,In_659,In_2420);
nor U1589 (N_1589,In_2209,In_103);
nand U1590 (N_1590,In_1328,In_2309);
and U1591 (N_1591,In_1854,In_706);
xnor U1592 (N_1592,In_2021,In_2225);
or U1593 (N_1593,In_29,In_2408);
nand U1594 (N_1594,In_1196,In_498);
and U1595 (N_1595,In_5,In_325);
xor U1596 (N_1596,In_1985,In_683);
nand U1597 (N_1597,In_530,In_2177);
nand U1598 (N_1598,In_1487,In_866);
and U1599 (N_1599,In_1949,In_205);
and U1600 (N_1600,In_922,In_1984);
and U1601 (N_1601,In_2010,In_541);
or U1602 (N_1602,In_803,In_95);
nand U1603 (N_1603,In_1553,In_2229);
xor U1604 (N_1604,In_1955,In_978);
and U1605 (N_1605,In_1700,In_390);
or U1606 (N_1606,In_974,In_422);
and U1607 (N_1607,In_196,In_2348);
and U1608 (N_1608,In_2229,In_1639);
nand U1609 (N_1609,In_1270,In_237);
or U1610 (N_1610,In_1372,In_1678);
or U1611 (N_1611,In_375,In_311);
or U1612 (N_1612,In_2490,In_775);
and U1613 (N_1613,In_2407,In_1218);
nor U1614 (N_1614,In_2259,In_155);
nand U1615 (N_1615,In_491,In_400);
nor U1616 (N_1616,In_86,In_81);
nor U1617 (N_1617,In_1058,In_2300);
and U1618 (N_1618,In_1397,In_553);
or U1619 (N_1619,In_1396,In_1406);
or U1620 (N_1620,In_218,In_1261);
nand U1621 (N_1621,In_489,In_1369);
xnor U1622 (N_1622,In_550,In_670);
or U1623 (N_1623,In_2046,In_2152);
or U1624 (N_1624,In_1390,In_1985);
or U1625 (N_1625,In_29,In_1154);
nand U1626 (N_1626,In_709,In_240);
nand U1627 (N_1627,In_1080,In_468);
nand U1628 (N_1628,In_1343,In_705);
and U1629 (N_1629,In_1359,In_86);
nand U1630 (N_1630,In_1313,In_1560);
nand U1631 (N_1631,In_1345,In_107);
xor U1632 (N_1632,In_1394,In_1299);
and U1633 (N_1633,In_1235,In_382);
nand U1634 (N_1634,In_2278,In_2219);
or U1635 (N_1635,In_2213,In_58);
and U1636 (N_1636,In_1409,In_2012);
nand U1637 (N_1637,In_1087,In_1030);
and U1638 (N_1638,In_1701,In_729);
nor U1639 (N_1639,In_998,In_1264);
and U1640 (N_1640,In_495,In_1144);
or U1641 (N_1641,In_2421,In_699);
nor U1642 (N_1642,In_1140,In_1291);
nand U1643 (N_1643,In_2304,In_4);
nor U1644 (N_1644,In_1968,In_2494);
or U1645 (N_1645,In_2187,In_1806);
nor U1646 (N_1646,In_1958,In_1162);
nor U1647 (N_1647,In_2097,In_2294);
nand U1648 (N_1648,In_1770,In_1907);
nand U1649 (N_1649,In_903,In_1038);
or U1650 (N_1650,In_616,In_519);
or U1651 (N_1651,In_292,In_1023);
nor U1652 (N_1652,In_482,In_539);
or U1653 (N_1653,In_332,In_371);
or U1654 (N_1654,In_944,In_2233);
or U1655 (N_1655,In_1049,In_1698);
or U1656 (N_1656,In_1004,In_2118);
nand U1657 (N_1657,In_823,In_1306);
xnor U1658 (N_1658,In_1282,In_29);
and U1659 (N_1659,In_2048,In_0);
nand U1660 (N_1660,In_1147,In_2461);
nor U1661 (N_1661,In_860,In_224);
and U1662 (N_1662,In_560,In_573);
nor U1663 (N_1663,In_2186,In_983);
nand U1664 (N_1664,In_1616,In_620);
and U1665 (N_1665,In_1063,In_820);
nor U1666 (N_1666,In_1350,In_1097);
nor U1667 (N_1667,In_2078,In_1142);
or U1668 (N_1668,In_1768,In_2137);
nand U1669 (N_1669,In_2430,In_1691);
nor U1670 (N_1670,In_2301,In_616);
nor U1671 (N_1671,In_628,In_1485);
nand U1672 (N_1672,In_619,In_1180);
xnor U1673 (N_1673,In_262,In_296);
and U1674 (N_1674,In_1108,In_1175);
nor U1675 (N_1675,In_273,In_2046);
and U1676 (N_1676,In_1880,In_885);
or U1677 (N_1677,In_937,In_1992);
or U1678 (N_1678,In_308,In_39);
and U1679 (N_1679,In_1177,In_1992);
nor U1680 (N_1680,In_176,In_181);
nor U1681 (N_1681,In_1031,In_728);
xnor U1682 (N_1682,In_2480,In_2283);
nor U1683 (N_1683,In_748,In_9);
nor U1684 (N_1684,In_1502,In_1801);
and U1685 (N_1685,In_237,In_1723);
nor U1686 (N_1686,In_1802,In_2473);
nand U1687 (N_1687,In_1465,In_98);
nand U1688 (N_1688,In_276,In_1041);
nand U1689 (N_1689,In_1837,In_516);
and U1690 (N_1690,In_321,In_1745);
nand U1691 (N_1691,In_863,In_910);
xnor U1692 (N_1692,In_1907,In_1935);
and U1693 (N_1693,In_705,In_1516);
nor U1694 (N_1694,In_667,In_633);
xnor U1695 (N_1695,In_1206,In_647);
and U1696 (N_1696,In_1801,In_258);
nor U1697 (N_1697,In_12,In_1710);
nand U1698 (N_1698,In_2123,In_1480);
nand U1699 (N_1699,In_490,In_1238);
and U1700 (N_1700,In_1704,In_803);
nor U1701 (N_1701,In_89,In_1915);
nand U1702 (N_1702,In_2415,In_348);
nor U1703 (N_1703,In_1333,In_1149);
or U1704 (N_1704,In_1789,In_2266);
xor U1705 (N_1705,In_2286,In_1392);
or U1706 (N_1706,In_213,In_1564);
nand U1707 (N_1707,In_638,In_1047);
xnor U1708 (N_1708,In_820,In_1006);
nor U1709 (N_1709,In_1259,In_1958);
and U1710 (N_1710,In_411,In_196);
and U1711 (N_1711,In_337,In_461);
xnor U1712 (N_1712,In_2457,In_2094);
xor U1713 (N_1713,In_1320,In_1954);
xor U1714 (N_1714,In_649,In_1293);
nand U1715 (N_1715,In_2311,In_2197);
nand U1716 (N_1716,In_1378,In_1277);
nand U1717 (N_1717,In_1390,In_566);
nand U1718 (N_1718,In_1502,In_1185);
or U1719 (N_1719,In_1732,In_997);
and U1720 (N_1720,In_1882,In_74);
nand U1721 (N_1721,In_496,In_747);
or U1722 (N_1722,In_1330,In_46);
nor U1723 (N_1723,In_490,In_873);
xnor U1724 (N_1724,In_218,In_380);
nor U1725 (N_1725,In_548,In_2404);
nand U1726 (N_1726,In_2271,In_1711);
nor U1727 (N_1727,In_1709,In_268);
nor U1728 (N_1728,In_2350,In_2111);
xor U1729 (N_1729,In_487,In_304);
nand U1730 (N_1730,In_986,In_2324);
and U1731 (N_1731,In_65,In_222);
nor U1732 (N_1732,In_150,In_363);
nand U1733 (N_1733,In_670,In_2259);
nor U1734 (N_1734,In_572,In_497);
xor U1735 (N_1735,In_809,In_1158);
nand U1736 (N_1736,In_1369,In_1126);
nand U1737 (N_1737,In_153,In_1327);
and U1738 (N_1738,In_1207,In_2007);
nor U1739 (N_1739,In_2280,In_1953);
nand U1740 (N_1740,In_1479,In_2353);
nand U1741 (N_1741,In_594,In_1651);
or U1742 (N_1742,In_2244,In_1557);
and U1743 (N_1743,In_1749,In_2099);
and U1744 (N_1744,In_1746,In_1411);
or U1745 (N_1745,In_1293,In_2165);
and U1746 (N_1746,In_1786,In_195);
nor U1747 (N_1747,In_1572,In_98);
or U1748 (N_1748,In_449,In_1838);
and U1749 (N_1749,In_2000,In_739);
nor U1750 (N_1750,In_2425,In_440);
nor U1751 (N_1751,In_1885,In_1971);
or U1752 (N_1752,In_948,In_1039);
and U1753 (N_1753,In_2141,In_886);
nor U1754 (N_1754,In_1317,In_1992);
nor U1755 (N_1755,In_2337,In_819);
nand U1756 (N_1756,In_2265,In_345);
or U1757 (N_1757,In_77,In_2100);
or U1758 (N_1758,In_472,In_244);
or U1759 (N_1759,In_339,In_2351);
and U1760 (N_1760,In_671,In_1485);
nand U1761 (N_1761,In_1784,In_1481);
nor U1762 (N_1762,In_1608,In_2432);
and U1763 (N_1763,In_68,In_1786);
and U1764 (N_1764,In_2218,In_1857);
nor U1765 (N_1765,In_1682,In_1931);
and U1766 (N_1766,In_2394,In_1621);
nand U1767 (N_1767,In_829,In_2407);
nor U1768 (N_1768,In_1435,In_369);
or U1769 (N_1769,In_1404,In_134);
nor U1770 (N_1770,In_1255,In_1717);
nor U1771 (N_1771,In_2160,In_1508);
nor U1772 (N_1772,In_229,In_1550);
and U1773 (N_1773,In_141,In_901);
or U1774 (N_1774,In_239,In_320);
and U1775 (N_1775,In_906,In_1157);
and U1776 (N_1776,In_1335,In_1804);
and U1777 (N_1777,In_454,In_2270);
or U1778 (N_1778,In_2376,In_2434);
and U1779 (N_1779,In_2061,In_735);
and U1780 (N_1780,In_136,In_888);
nor U1781 (N_1781,In_982,In_151);
or U1782 (N_1782,In_1883,In_1088);
nand U1783 (N_1783,In_2016,In_759);
nor U1784 (N_1784,In_1041,In_1514);
nand U1785 (N_1785,In_324,In_856);
nand U1786 (N_1786,In_665,In_1193);
nor U1787 (N_1787,In_588,In_966);
and U1788 (N_1788,In_1381,In_1704);
nor U1789 (N_1789,In_914,In_494);
or U1790 (N_1790,In_709,In_1094);
or U1791 (N_1791,In_1945,In_974);
nand U1792 (N_1792,In_552,In_779);
nor U1793 (N_1793,In_146,In_681);
xor U1794 (N_1794,In_163,In_1474);
nand U1795 (N_1795,In_484,In_1171);
nand U1796 (N_1796,In_2061,In_235);
and U1797 (N_1797,In_2062,In_937);
and U1798 (N_1798,In_1143,In_2387);
nor U1799 (N_1799,In_1736,In_1878);
nand U1800 (N_1800,In_2394,In_2076);
nor U1801 (N_1801,In_1875,In_781);
or U1802 (N_1802,In_2473,In_2221);
and U1803 (N_1803,In_2279,In_26);
and U1804 (N_1804,In_1518,In_1956);
xor U1805 (N_1805,In_150,In_1104);
and U1806 (N_1806,In_1353,In_1270);
xnor U1807 (N_1807,In_2314,In_185);
or U1808 (N_1808,In_1043,In_1003);
xor U1809 (N_1809,In_1968,In_1016);
nand U1810 (N_1810,In_800,In_218);
nand U1811 (N_1811,In_2249,In_1372);
or U1812 (N_1812,In_24,In_1642);
and U1813 (N_1813,In_1623,In_1021);
xor U1814 (N_1814,In_1466,In_1444);
nand U1815 (N_1815,In_1229,In_1165);
and U1816 (N_1816,In_2214,In_1516);
or U1817 (N_1817,In_2252,In_610);
xor U1818 (N_1818,In_1912,In_1293);
or U1819 (N_1819,In_1171,In_470);
nand U1820 (N_1820,In_231,In_723);
nor U1821 (N_1821,In_1985,In_337);
nand U1822 (N_1822,In_1745,In_557);
and U1823 (N_1823,In_1524,In_893);
or U1824 (N_1824,In_2031,In_2166);
and U1825 (N_1825,In_1151,In_1285);
xnor U1826 (N_1826,In_2230,In_2271);
nor U1827 (N_1827,In_1953,In_1205);
or U1828 (N_1828,In_606,In_1508);
xor U1829 (N_1829,In_2327,In_1258);
and U1830 (N_1830,In_2394,In_2212);
nor U1831 (N_1831,In_1627,In_629);
and U1832 (N_1832,In_721,In_325);
or U1833 (N_1833,In_2154,In_1705);
and U1834 (N_1834,In_312,In_155);
and U1835 (N_1835,In_2152,In_1101);
nor U1836 (N_1836,In_1491,In_1001);
nand U1837 (N_1837,In_1393,In_1413);
or U1838 (N_1838,In_824,In_2056);
nor U1839 (N_1839,In_1524,In_2134);
nor U1840 (N_1840,In_2259,In_279);
or U1841 (N_1841,In_2450,In_964);
or U1842 (N_1842,In_1937,In_444);
or U1843 (N_1843,In_293,In_2350);
nand U1844 (N_1844,In_1916,In_1058);
or U1845 (N_1845,In_395,In_389);
and U1846 (N_1846,In_1582,In_824);
and U1847 (N_1847,In_1449,In_1110);
or U1848 (N_1848,In_802,In_1285);
nand U1849 (N_1849,In_489,In_87);
nand U1850 (N_1850,In_1202,In_1521);
nand U1851 (N_1851,In_831,In_1488);
nand U1852 (N_1852,In_907,In_1256);
xnor U1853 (N_1853,In_732,In_422);
or U1854 (N_1854,In_1164,In_324);
nor U1855 (N_1855,In_2368,In_373);
nor U1856 (N_1856,In_1141,In_1242);
and U1857 (N_1857,In_1593,In_1680);
xnor U1858 (N_1858,In_111,In_1506);
nor U1859 (N_1859,In_2373,In_1163);
nand U1860 (N_1860,In_1536,In_899);
nand U1861 (N_1861,In_2104,In_1195);
xnor U1862 (N_1862,In_1950,In_1182);
nor U1863 (N_1863,In_1601,In_1455);
and U1864 (N_1864,In_1753,In_1429);
or U1865 (N_1865,In_977,In_340);
and U1866 (N_1866,In_1714,In_1226);
and U1867 (N_1867,In_682,In_2219);
nor U1868 (N_1868,In_1838,In_1831);
or U1869 (N_1869,In_2192,In_1779);
nand U1870 (N_1870,In_1408,In_390);
nand U1871 (N_1871,In_668,In_1429);
nor U1872 (N_1872,In_46,In_1441);
xnor U1873 (N_1873,In_722,In_1799);
or U1874 (N_1874,In_657,In_871);
nand U1875 (N_1875,In_1546,In_749);
nor U1876 (N_1876,In_2225,In_1832);
or U1877 (N_1877,In_1574,In_1990);
nand U1878 (N_1878,In_1810,In_401);
and U1879 (N_1879,In_729,In_2153);
nor U1880 (N_1880,In_1676,In_1108);
xnor U1881 (N_1881,In_1869,In_538);
nand U1882 (N_1882,In_2176,In_2310);
nand U1883 (N_1883,In_242,In_375);
and U1884 (N_1884,In_1729,In_2490);
or U1885 (N_1885,In_283,In_2389);
nand U1886 (N_1886,In_2435,In_74);
nor U1887 (N_1887,In_1867,In_471);
and U1888 (N_1888,In_556,In_771);
nand U1889 (N_1889,In_1871,In_2058);
and U1890 (N_1890,In_1551,In_246);
and U1891 (N_1891,In_2032,In_1113);
and U1892 (N_1892,In_2358,In_2239);
and U1893 (N_1893,In_2382,In_1897);
xnor U1894 (N_1894,In_1130,In_389);
nand U1895 (N_1895,In_417,In_534);
nand U1896 (N_1896,In_1447,In_1070);
nand U1897 (N_1897,In_429,In_1726);
and U1898 (N_1898,In_1,In_2393);
or U1899 (N_1899,In_2172,In_226);
and U1900 (N_1900,In_1325,In_1797);
nor U1901 (N_1901,In_2238,In_1956);
and U1902 (N_1902,In_623,In_725);
xor U1903 (N_1903,In_1390,In_370);
and U1904 (N_1904,In_1499,In_1405);
nor U1905 (N_1905,In_1404,In_2464);
or U1906 (N_1906,In_2121,In_2105);
or U1907 (N_1907,In_723,In_230);
and U1908 (N_1908,In_199,In_2261);
nor U1909 (N_1909,In_1414,In_391);
nand U1910 (N_1910,In_1846,In_1910);
nor U1911 (N_1911,In_506,In_2330);
nand U1912 (N_1912,In_382,In_1127);
nor U1913 (N_1913,In_1144,In_2377);
and U1914 (N_1914,In_2404,In_1662);
and U1915 (N_1915,In_976,In_338);
or U1916 (N_1916,In_1532,In_98);
nor U1917 (N_1917,In_12,In_291);
nand U1918 (N_1918,In_1677,In_990);
and U1919 (N_1919,In_1663,In_1312);
and U1920 (N_1920,In_1085,In_322);
xnor U1921 (N_1921,In_1383,In_919);
xnor U1922 (N_1922,In_1815,In_1950);
nand U1923 (N_1923,In_1450,In_43);
nand U1924 (N_1924,In_317,In_300);
or U1925 (N_1925,In_708,In_371);
nor U1926 (N_1926,In_477,In_865);
xor U1927 (N_1927,In_1141,In_1429);
nand U1928 (N_1928,In_1622,In_1523);
nand U1929 (N_1929,In_2192,In_94);
or U1930 (N_1930,In_277,In_1454);
nor U1931 (N_1931,In_404,In_1335);
nor U1932 (N_1932,In_2280,In_2007);
or U1933 (N_1933,In_2349,In_1328);
or U1934 (N_1934,In_2359,In_115);
and U1935 (N_1935,In_1718,In_2171);
nor U1936 (N_1936,In_252,In_1654);
and U1937 (N_1937,In_260,In_1440);
and U1938 (N_1938,In_1554,In_1962);
nor U1939 (N_1939,In_2108,In_1787);
nor U1940 (N_1940,In_845,In_1657);
nor U1941 (N_1941,In_2396,In_896);
and U1942 (N_1942,In_1587,In_1369);
and U1943 (N_1943,In_1162,In_767);
nand U1944 (N_1944,In_180,In_764);
nor U1945 (N_1945,In_2271,In_2483);
nand U1946 (N_1946,In_2256,In_948);
xor U1947 (N_1947,In_1580,In_61);
xor U1948 (N_1948,In_2368,In_787);
xnor U1949 (N_1949,In_596,In_2491);
nand U1950 (N_1950,In_612,In_2195);
nand U1951 (N_1951,In_82,In_264);
and U1952 (N_1952,In_1664,In_1299);
nand U1953 (N_1953,In_1695,In_1915);
nor U1954 (N_1954,In_648,In_230);
and U1955 (N_1955,In_1932,In_457);
and U1956 (N_1956,In_92,In_1954);
and U1957 (N_1957,In_575,In_312);
xnor U1958 (N_1958,In_1864,In_1954);
or U1959 (N_1959,In_2287,In_499);
or U1960 (N_1960,In_1972,In_817);
nor U1961 (N_1961,In_1911,In_1779);
or U1962 (N_1962,In_2189,In_616);
nand U1963 (N_1963,In_1311,In_968);
nand U1964 (N_1964,In_242,In_2238);
and U1965 (N_1965,In_672,In_1347);
and U1966 (N_1966,In_1921,In_89);
and U1967 (N_1967,In_521,In_1632);
xnor U1968 (N_1968,In_1781,In_958);
xor U1969 (N_1969,In_777,In_964);
nand U1970 (N_1970,In_1073,In_1001);
or U1971 (N_1971,In_151,In_2066);
and U1972 (N_1972,In_769,In_127);
and U1973 (N_1973,In_36,In_1206);
nand U1974 (N_1974,In_2427,In_97);
and U1975 (N_1975,In_281,In_1310);
nand U1976 (N_1976,In_2203,In_2063);
xor U1977 (N_1977,In_1537,In_242);
and U1978 (N_1978,In_2458,In_929);
nand U1979 (N_1979,In_115,In_2029);
and U1980 (N_1980,In_2470,In_860);
nor U1981 (N_1981,In_1232,In_457);
nor U1982 (N_1982,In_1268,In_1801);
nor U1983 (N_1983,In_1684,In_2141);
and U1984 (N_1984,In_2232,In_955);
xnor U1985 (N_1985,In_726,In_1613);
xor U1986 (N_1986,In_958,In_1630);
nand U1987 (N_1987,In_1979,In_81);
or U1988 (N_1988,In_326,In_2266);
or U1989 (N_1989,In_1394,In_1213);
or U1990 (N_1990,In_859,In_1026);
or U1991 (N_1991,In_623,In_1040);
xnor U1992 (N_1992,In_1785,In_649);
nor U1993 (N_1993,In_150,In_727);
nand U1994 (N_1994,In_1020,In_2096);
or U1995 (N_1995,In_2246,In_2482);
nand U1996 (N_1996,In_1318,In_2451);
nand U1997 (N_1997,In_2334,In_1194);
or U1998 (N_1998,In_189,In_1397);
nor U1999 (N_1999,In_1379,In_942);
and U2000 (N_2000,In_1029,In_1239);
xor U2001 (N_2001,In_72,In_1819);
nor U2002 (N_2002,In_2170,In_1567);
nand U2003 (N_2003,In_411,In_1639);
nand U2004 (N_2004,In_997,In_951);
nand U2005 (N_2005,In_705,In_787);
xnor U2006 (N_2006,In_69,In_2107);
xor U2007 (N_2007,In_437,In_1393);
xnor U2008 (N_2008,In_1638,In_1864);
xor U2009 (N_2009,In_477,In_39);
nand U2010 (N_2010,In_1480,In_2302);
nand U2011 (N_2011,In_890,In_2075);
and U2012 (N_2012,In_184,In_1583);
nand U2013 (N_2013,In_698,In_303);
and U2014 (N_2014,In_2326,In_93);
nor U2015 (N_2015,In_1538,In_2358);
and U2016 (N_2016,In_2181,In_1889);
nor U2017 (N_2017,In_1273,In_1348);
nand U2018 (N_2018,In_427,In_1263);
or U2019 (N_2019,In_1896,In_2287);
or U2020 (N_2020,In_1209,In_67);
nor U2021 (N_2021,In_540,In_884);
nand U2022 (N_2022,In_2410,In_1446);
nor U2023 (N_2023,In_1182,In_727);
xor U2024 (N_2024,In_1135,In_1192);
nand U2025 (N_2025,In_1408,In_750);
nand U2026 (N_2026,In_1605,In_1722);
nor U2027 (N_2027,In_858,In_2075);
nand U2028 (N_2028,In_580,In_1443);
or U2029 (N_2029,In_375,In_2344);
or U2030 (N_2030,In_2259,In_2335);
and U2031 (N_2031,In_1352,In_1215);
and U2032 (N_2032,In_2064,In_32);
or U2033 (N_2033,In_484,In_1594);
nor U2034 (N_2034,In_219,In_1199);
or U2035 (N_2035,In_1117,In_838);
or U2036 (N_2036,In_122,In_2228);
nor U2037 (N_2037,In_176,In_1593);
and U2038 (N_2038,In_2285,In_2245);
and U2039 (N_2039,In_172,In_888);
nand U2040 (N_2040,In_269,In_1530);
xnor U2041 (N_2041,In_542,In_1986);
nand U2042 (N_2042,In_981,In_2477);
and U2043 (N_2043,In_1329,In_1026);
or U2044 (N_2044,In_154,In_2260);
and U2045 (N_2045,In_62,In_434);
nor U2046 (N_2046,In_1568,In_935);
nor U2047 (N_2047,In_727,In_1220);
xor U2048 (N_2048,In_1968,In_1483);
nand U2049 (N_2049,In_758,In_499);
or U2050 (N_2050,In_2250,In_1544);
or U2051 (N_2051,In_205,In_1025);
xnor U2052 (N_2052,In_880,In_570);
nand U2053 (N_2053,In_1287,In_1531);
nor U2054 (N_2054,In_308,In_730);
and U2055 (N_2055,In_206,In_2146);
or U2056 (N_2056,In_1899,In_1529);
xnor U2057 (N_2057,In_527,In_1087);
nor U2058 (N_2058,In_171,In_945);
nor U2059 (N_2059,In_235,In_626);
nand U2060 (N_2060,In_2311,In_1402);
and U2061 (N_2061,In_2101,In_2205);
and U2062 (N_2062,In_1670,In_97);
nor U2063 (N_2063,In_1891,In_684);
xnor U2064 (N_2064,In_2233,In_2021);
nor U2065 (N_2065,In_1723,In_1929);
and U2066 (N_2066,In_167,In_475);
nor U2067 (N_2067,In_509,In_1172);
nand U2068 (N_2068,In_1195,In_2350);
or U2069 (N_2069,In_2417,In_2488);
or U2070 (N_2070,In_1115,In_2255);
xnor U2071 (N_2071,In_1220,In_2005);
nand U2072 (N_2072,In_2354,In_1527);
xnor U2073 (N_2073,In_670,In_2238);
nor U2074 (N_2074,In_2128,In_1695);
or U2075 (N_2075,In_2036,In_783);
xnor U2076 (N_2076,In_2442,In_1416);
and U2077 (N_2077,In_2436,In_1229);
and U2078 (N_2078,In_1190,In_752);
and U2079 (N_2079,In_139,In_966);
or U2080 (N_2080,In_841,In_488);
nand U2081 (N_2081,In_1097,In_54);
or U2082 (N_2082,In_2247,In_987);
nor U2083 (N_2083,In_1683,In_1924);
and U2084 (N_2084,In_192,In_1510);
and U2085 (N_2085,In_1023,In_393);
nand U2086 (N_2086,In_343,In_2116);
nand U2087 (N_2087,In_2122,In_1818);
or U2088 (N_2088,In_734,In_538);
or U2089 (N_2089,In_748,In_2440);
xor U2090 (N_2090,In_1752,In_2339);
nand U2091 (N_2091,In_1222,In_629);
and U2092 (N_2092,In_1312,In_1509);
nand U2093 (N_2093,In_2247,In_1186);
nor U2094 (N_2094,In_1159,In_2446);
or U2095 (N_2095,In_1684,In_1855);
or U2096 (N_2096,In_507,In_1089);
nor U2097 (N_2097,In_1347,In_450);
nor U2098 (N_2098,In_496,In_1542);
and U2099 (N_2099,In_286,In_2225);
or U2100 (N_2100,In_1869,In_1123);
nand U2101 (N_2101,In_2010,In_235);
nor U2102 (N_2102,In_54,In_147);
nand U2103 (N_2103,In_1094,In_1861);
or U2104 (N_2104,In_530,In_615);
or U2105 (N_2105,In_898,In_1091);
or U2106 (N_2106,In_127,In_1268);
and U2107 (N_2107,In_1730,In_1511);
nand U2108 (N_2108,In_1228,In_499);
and U2109 (N_2109,In_2476,In_2077);
nand U2110 (N_2110,In_1177,In_1611);
nand U2111 (N_2111,In_129,In_463);
and U2112 (N_2112,In_833,In_1169);
and U2113 (N_2113,In_998,In_836);
and U2114 (N_2114,In_1883,In_164);
or U2115 (N_2115,In_1596,In_1693);
and U2116 (N_2116,In_1489,In_240);
and U2117 (N_2117,In_987,In_2017);
or U2118 (N_2118,In_1840,In_1382);
nand U2119 (N_2119,In_428,In_190);
nand U2120 (N_2120,In_1040,In_633);
nand U2121 (N_2121,In_309,In_2252);
nand U2122 (N_2122,In_2410,In_1315);
and U2123 (N_2123,In_1960,In_1711);
nor U2124 (N_2124,In_1766,In_918);
nor U2125 (N_2125,In_11,In_1176);
nand U2126 (N_2126,In_953,In_2300);
nand U2127 (N_2127,In_1799,In_1013);
nand U2128 (N_2128,In_2020,In_378);
nand U2129 (N_2129,In_1009,In_2298);
or U2130 (N_2130,In_1347,In_2400);
nand U2131 (N_2131,In_596,In_1014);
nor U2132 (N_2132,In_376,In_1594);
and U2133 (N_2133,In_1030,In_1600);
or U2134 (N_2134,In_1620,In_2390);
and U2135 (N_2135,In_1924,In_958);
xor U2136 (N_2136,In_2469,In_1747);
or U2137 (N_2137,In_82,In_1711);
nor U2138 (N_2138,In_19,In_1121);
or U2139 (N_2139,In_1326,In_792);
and U2140 (N_2140,In_1175,In_280);
xnor U2141 (N_2141,In_352,In_1430);
and U2142 (N_2142,In_2065,In_1302);
nand U2143 (N_2143,In_1938,In_1860);
or U2144 (N_2144,In_460,In_2195);
or U2145 (N_2145,In_2086,In_1296);
and U2146 (N_2146,In_1796,In_950);
or U2147 (N_2147,In_2194,In_231);
and U2148 (N_2148,In_2441,In_2124);
nand U2149 (N_2149,In_1378,In_1013);
and U2150 (N_2150,In_979,In_1678);
nor U2151 (N_2151,In_550,In_381);
nand U2152 (N_2152,In_1575,In_2356);
nand U2153 (N_2153,In_1643,In_1609);
and U2154 (N_2154,In_2405,In_295);
xnor U2155 (N_2155,In_2143,In_57);
nor U2156 (N_2156,In_1121,In_961);
nor U2157 (N_2157,In_862,In_1343);
xnor U2158 (N_2158,In_180,In_1928);
nand U2159 (N_2159,In_1153,In_484);
nand U2160 (N_2160,In_1005,In_807);
nor U2161 (N_2161,In_2018,In_2138);
or U2162 (N_2162,In_2006,In_2493);
nor U2163 (N_2163,In_1744,In_477);
and U2164 (N_2164,In_505,In_1696);
nor U2165 (N_2165,In_337,In_571);
nand U2166 (N_2166,In_2306,In_1575);
nand U2167 (N_2167,In_593,In_724);
nor U2168 (N_2168,In_2362,In_1566);
nor U2169 (N_2169,In_1715,In_575);
nand U2170 (N_2170,In_1871,In_1615);
xor U2171 (N_2171,In_262,In_1304);
nand U2172 (N_2172,In_1943,In_1243);
xor U2173 (N_2173,In_1410,In_1944);
or U2174 (N_2174,In_1749,In_1637);
nor U2175 (N_2175,In_2058,In_1392);
nor U2176 (N_2176,In_2327,In_1572);
and U2177 (N_2177,In_474,In_499);
nor U2178 (N_2178,In_489,In_1636);
nand U2179 (N_2179,In_484,In_1870);
nor U2180 (N_2180,In_600,In_2212);
nand U2181 (N_2181,In_577,In_2095);
nand U2182 (N_2182,In_428,In_2326);
nor U2183 (N_2183,In_2116,In_2267);
nand U2184 (N_2184,In_191,In_1292);
nor U2185 (N_2185,In_1790,In_68);
or U2186 (N_2186,In_2232,In_2289);
nor U2187 (N_2187,In_1700,In_1948);
nand U2188 (N_2188,In_1832,In_2161);
nor U2189 (N_2189,In_2220,In_70);
and U2190 (N_2190,In_1992,In_1657);
and U2191 (N_2191,In_2179,In_2192);
xor U2192 (N_2192,In_2266,In_2480);
nand U2193 (N_2193,In_2300,In_1244);
and U2194 (N_2194,In_293,In_1119);
xnor U2195 (N_2195,In_544,In_1585);
or U2196 (N_2196,In_2383,In_2003);
and U2197 (N_2197,In_880,In_1648);
nand U2198 (N_2198,In_529,In_2414);
nand U2199 (N_2199,In_1504,In_2261);
nand U2200 (N_2200,In_90,In_876);
nor U2201 (N_2201,In_259,In_717);
or U2202 (N_2202,In_141,In_556);
nand U2203 (N_2203,In_2368,In_1507);
nand U2204 (N_2204,In_946,In_385);
xor U2205 (N_2205,In_849,In_1896);
or U2206 (N_2206,In_1332,In_1513);
nor U2207 (N_2207,In_2451,In_2394);
nor U2208 (N_2208,In_761,In_2230);
or U2209 (N_2209,In_615,In_529);
or U2210 (N_2210,In_388,In_2278);
or U2211 (N_2211,In_101,In_929);
nor U2212 (N_2212,In_760,In_448);
and U2213 (N_2213,In_828,In_930);
nor U2214 (N_2214,In_511,In_146);
or U2215 (N_2215,In_181,In_1125);
and U2216 (N_2216,In_2098,In_1929);
and U2217 (N_2217,In_832,In_1163);
or U2218 (N_2218,In_1446,In_542);
nor U2219 (N_2219,In_2179,In_2485);
or U2220 (N_2220,In_2329,In_495);
xor U2221 (N_2221,In_2325,In_2386);
nand U2222 (N_2222,In_1642,In_1509);
nand U2223 (N_2223,In_2281,In_788);
xnor U2224 (N_2224,In_817,In_939);
and U2225 (N_2225,In_2369,In_1128);
nor U2226 (N_2226,In_763,In_377);
nor U2227 (N_2227,In_859,In_1750);
nor U2228 (N_2228,In_1548,In_1899);
nor U2229 (N_2229,In_1779,In_1394);
nand U2230 (N_2230,In_1554,In_210);
and U2231 (N_2231,In_416,In_1037);
or U2232 (N_2232,In_426,In_1578);
nor U2233 (N_2233,In_1407,In_1261);
or U2234 (N_2234,In_1344,In_1330);
nand U2235 (N_2235,In_837,In_1509);
nand U2236 (N_2236,In_1692,In_105);
nand U2237 (N_2237,In_2285,In_2077);
nor U2238 (N_2238,In_487,In_1528);
nor U2239 (N_2239,In_1778,In_261);
and U2240 (N_2240,In_215,In_969);
or U2241 (N_2241,In_2455,In_715);
nor U2242 (N_2242,In_1542,In_2047);
nand U2243 (N_2243,In_271,In_2417);
and U2244 (N_2244,In_1630,In_1034);
and U2245 (N_2245,In_801,In_1044);
or U2246 (N_2246,In_567,In_1426);
xnor U2247 (N_2247,In_1380,In_2185);
nor U2248 (N_2248,In_847,In_1953);
nand U2249 (N_2249,In_1741,In_278);
nand U2250 (N_2250,In_2093,In_1832);
and U2251 (N_2251,In_1572,In_1126);
or U2252 (N_2252,In_275,In_1708);
nand U2253 (N_2253,In_1614,In_1005);
and U2254 (N_2254,In_1550,In_974);
nand U2255 (N_2255,In_2250,In_648);
nand U2256 (N_2256,In_1137,In_2041);
or U2257 (N_2257,In_593,In_2229);
nand U2258 (N_2258,In_2059,In_135);
nand U2259 (N_2259,In_47,In_226);
xnor U2260 (N_2260,In_1146,In_314);
nand U2261 (N_2261,In_1038,In_2323);
or U2262 (N_2262,In_229,In_1120);
nand U2263 (N_2263,In_622,In_1426);
xnor U2264 (N_2264,In_1197,In_173);
xnor U2265 (N_2265,In_172,In_2122);
and U2266 (N_2266,In_934,In_277);
nand U2267 (N_2267,In_1105,In_2109);
nor U2268 (N_2268,In_467,In_748);
and U2269 (N_2269,In_119,In_698);
nor U2270 (N_2270,In_580,In_924);
and U2271 (N_2271,In_2400,In_887);
nand U2272 (N_2272,In_853,In_2136);
or U2273 (N_2273,In_289,In_1409);
xor U2274 (N_2274,In_1223,In_2475);
nor U2275 (N_2275,In_1215,In_2378);
nor U2276 (N_2276,In_1627,In_805);
or U2277 (N_2277,In_1101,In_286);
or U2278 (N_2278,In_983,In_1958);
nand U2279 (N_2279,In_666,In_920);
and U2280 (N_2280,In_1655,In_1418);
nor U2281 (N_2281,In_1184,In_242);
xnor U2282 (N_2282,In_1792,In_1498);
nand U2283 (N_2283,In_1883,In_1391);
nor U2284 (N_2284,In_1748,In_840);
nor U2285 (N_2285,In_266,In_26);
and U2286 (N_2286,In_818,In_2137);
nand U2287 (N_2287,In_2487,In_1441);
or U2288 (N_2288,In_1994,In_2099);
nand U2289 (N_2289,In_898,In_1235);
or U2290 (N_2290,In_1687,In_2001);
nor U2291 (N_2291,In_433,In_1650);
or U2292 (N_2292,In_1741,In_794);
nand U2293 (N_2293,In_29,In_1198);
nor U2294 (N_2294,In_1827,In_2260);
or U2295 (N_2295,In_231,In_1597);
and U2296 (N_2296,In_2461,In_6);
and U2297 (N_2297,In_334,In_320);
xor U2298 (N_2298,In_893,In_2465);
nand U2299 (N_2299,In_2329,In_2157);
and U2300 (N_2300,In_37,In_1249);
nor U2301 (N_2301,In_1947,In_1306);
and U2302 (N_2302,In_625,In_602);
and U2303 (N_2303,In_1482,In_316);
nor U2304 (N_2304,In_265,In_662);
nor U2305 (N_2305,In_2340,In_416);
or U2306 (N_2306,In_514,In_1364);
and U2307 (N_2307,In_1015,In_924);
nand U2308 (N_2308,In_401,In_1921);
nand U2309 (N_2309,In_827,In_402);
and U2310 (N_2310,In_1769,In_2180);
and U2311 (N_2311,In_1544,In_507);
nand U2312 (N_2312,In_870,In_2114);
or U2313 (N_2313,In_1208,In_704);
nand U2314 (N_2314,In_1888,In_1771);
nand U2315 (N_2315,In_2260,In_2390);
nor U2316 (N_2316,In_138,In_274);
and U2317 (N_2317,In_1059,In_32);
or U2318 (N_2318,In_2277,In_908);
nor U2319 (N_2319,In_552,In_1242);
or U2320 (N_2320,In_1244,In_862);
and U2321 (N_2321,In_106,In_692);
or U2322 (N_2322,In_967,In_2430);
nand U2323 (N_2323,In_1654,In_2224);
and U2324 (N_2324,In_782,In_625);
nor U2325 (N_2325,In_972,In_1853);
xor U2326 (N_2326,In_2111,In_1957);
nand U2327 (N_2327,In_68,In_2386);
xor U2328 (N_2328,In_1503,In_523);
nor U2329 (N_2329,In_1867,In_106);
or U2330 (N_2330,In_845,In_2156);
nor U2331 (N_2331,In_826,In_214);
xnor U2332 (N_2332,In_1714,In_1644);
nor U2333 (N_2333,In_87,In_1301);
nand U2334 (N_2334,In_508,In_1812);
and U2335 (N_2335,In_360,In_1698);
nor U2336 (N_2336,In_288,In_1700);
nand U2337 (N_2337,In_462,In_2207);
nor U2338 (N_2338,In_938,In_1663);
or U2339 (N_2339,In_1508,In_780);
nor U2340 (N_2340,In_511,In_1829);
nand U2341 (N_2341,In_218,In_1299);
nor U2342 (N_2342,In_571,In_915);
or U2343 (N_2343,In_1957,In_2283);
nand U2344 (N_2344,In_986,In_785);
and U2345 (N_2345,In_207,In_1586);
nor U2346 (N_2346,In_378,In_1518);
xnor U2347 (N_2347,In_791,In_181);
nor U2348 (N_2348,In_1213,In_1046);
and U2349 (N_2349,In_826,In_1980);
or U2350 (N_2350,In_15,In_806);
xnor U2351 (N_2351,In_195,In_1341);
nand U2352 (N_2352,In_780,In_845);
and U2353 (N_2353,In_2089,In_1884);
or U2354 (N_2354,In_447,In_1253);
or U2355 (N_2355,In_857,In_1811);
nand U2356 (N_2356,In_572,In_1689);
or U2357 (N_2357,In_48,In_142);
nand U2358 (N_2358,In_2244,In_1880);
nor U2359 (N_2359,In_315,In_619);
or U2360 (N_2360,In_1810,In_1150);
nor U2361 (N_2361,In_1443,In_2092);
nor U2362 (N_2362,In_788,In_1628);
nor U2363 (N_2363,In_1263,In_708);
and U2364 (N_2364,In_1036,In_1381);
nor U2365 (N_2365,In_257,In_1137);
nor U2366 (N_2366,In_1735,In_141);
xor U2367 (N_2367,In_37,In_1222);
or U2368 (N_2368,In_1837,In_788);
and U2369 (N_2369,In_2476,In_458);
nand U2370 (N_2370,In_2245,In_916);
nand U2371 (N_2371,In_1700,In_295);
or U2372 (N_2372,In_179,In_452);
nor U2373 (N_2373,In_1834,In_887);
or U2374 (N_2374,In_34,In_1651);
nor U2375 (N_2375,In_1615,In_506);
nand U2376 (N_2376,In_1511,In_1366);
and U2377 (N_2377,In_2125,In_1666);
and U2378 (N_2378,In_146,In_910);
or U2379 (N_2379,In_715,In_2413);
or U2380 (N_2380,In_1670,In_2071);
nand U2381 (N_2381,In_1218,In_541);
or U2382 (N_2382,In_2440,In_330);
nand U2383 (N_2383,In_2350,In_638);
or U2384 (N_2384,In_1843,In_543);
and U2385 (N_2385,In_2250,In_2216);
xnor U2386 (N_2386,In_1580,In_7);
nand U2387 (N_2387,In_124,In_2252);
or U2388 (N_2388,In_1050,In_624);
nand U2389 (N_2389,In_449,In_1932);
nor U2390 (N_2390,In_652,In_1439);
or U2391 (N_2391,In_2427,In_1617);
and U2392 (N_2392,In_1476,In_960);
or U2393 (N_2393,In_456,In_708);
nor U2394 (N_2394,In_1137,In_1521);
or U2395 (N_2395,In_68,In_865);
or U2396 (N_2396,In_17,In_1874);
nand U2397 (N_2397,In_1964,In_905);
and U2398 (N_2398,In_6,In_1130);
and U2399 (N_2399,In_691,In_2310);
xnor U2400 (N_2400,In_1085,In_401);
nand U2401 (N_2401,In_2202,In_1043);
nand U2402 (N_2402,In_241,In_110);
or U2403 (N_2403,In_1145,In_371);
nor U2404 (N_2404,In_925,In_2452);
or U2405 (N_2405,In_1775,In_1770);
or U2406 (N_2406,In_1149,In_2263);
nand U2407 (N_2407,In_1964,In_1435);
or U2408 (N_2408,In_231,In_879);
nor U2409 (N_2409,In_1798,In_1348);
or U2410 (N_2410,In_2049,In_2335);
and U2411 (N_2411,In_2399,In_661);
nand U2412 (N_2412,In_737,In_1508);
and U2413 (N_2413,In_674,In_510);
or U2414 (N_2414,In_1000,In_1160);
nor U2415 (N_2415,In_892,In_2030);
xor U2416 (N_2416,In_1631,In_332);
or U2417 (N_2417,In_84,In_1424);
nor U2418 (N_2418,In_96,In_544);
nand U2419 (N_2419,In_1638,In_1980);
and U2420 (N_2420,In_339,In_2099);
or U2421 (N_2421,In_1105,In_742);
nand U2422 (N_2422,In_2267,In_992);
nand U2423 (N_2423,In_2322,In_833);
nand U2424 (N_2424,In_1415,In_1813);
nand U2425 (N_2425,In_934,In_946);
nand U2426 (N_2426,In_2488,In_1223);
xnor U2427 (N_2427,In_1263,In_1024);
xor U2428 (N_2428,In_493,In_1977);
nor U2429 (N_2429,In_315,In_1390);
or U2430 (N_2430,In_2260,In_614);
and U2431 (N_2431,In_1837,In_1957);
or U2432 (N_2432,In_2460,In_1924);
or U2433 (N_2433,In_1796,In_930);
and U2434 (N_2434,In_2,In_486);
nor U2435 (N_2435,In_1330,In_1228);
and U2436 (N_2436,In_2081,In_321);
nand U2437 (N_2437,In_476,In_249);
or U2438 (N_2438,In_1444,In_420);
nor U2439 (N_2439,In_1851,In_1433);
nor U2440 (N_2440,In_1042,In_87);
and U2441 (N_2441,In_1030,In_2080);
nor U2442 (N_2442,In_1747,In_293);
or U2443 (N_2443,In_1924,In_2219);
and U2444 (N_2444,In_988,In_82);
nand U2445 (N_2445,In_1257,In_138);
nor U2446 (N_2446,In_2344,In_1864);
or U2447 (N_2447,In_1431,In_598);
nor U2448 (N_2448,In_2273,In_85);
nand U2449 (N_2449,In_928,In_1437);
nor U2450 (N_2450,In_1972,In_311);
nor U2451 (N_2451,In_2191,In_1205);
and U2452 (N_2452,In_80,In_1936);
and U2453 (N_2453,In_619,In_1914);
xor U2454 (N_2454,In_1995,In_588);
xnor U2455 (N_2455,In_949,In_2209);
nand U2456 (N_2456,In_474,In_1632);
nor U2457 (N_2457,In_1089,In_1970);
nand U2458 (N_2458,In_2401,In_555);
nand U2459 (N_2459,In_2216,In_1395);
and U2460 (N_2460,In_58,In_1584);
nand U2461 (N_2461,In_714,In_324);
nor U2462 (N_2462,In_1718,In_1366);
or U2463 (N_2463,In_492,In_717);
nor U2464 (N_2464,In_753,In_1428);
nor U2465 (N_2465,In_1224,In_34);
nor U2466 (N_2466,In_807,In_1121);
or U2467 (N_2467,In_485,In_953);
nand U2468 (N_2468,In_29,In_1148);
nor U2469 (N_2469,In_2098,In_2088);
nand U2470 (N_2470,In_1162,In_316);
nor U2471 (N_2471,In_2007,In_1717);
nor U2472 (N_2472,In_543,In_105);
or U2473 (N_2473,In_721,In_1227);
xor U2474 (N_2474,In_771,In_750);
nor U2475 (N_2475,In_203,In_1150);
and U2476 (N_2476,In_2413,In_942);
xnor U2477 (N_2477,In_1926,In_1076);
and U2478 (N_2478,In_908,In_1593);
and U2479 (N_2479,In_585,In_2480);
or U2480 (N_2480,In_493,In_959);
and U2481 (N_2481,In_190,In_1985);
xnor U2482 (N_2482,In_1996,In_704);
and U2483 (N_2483,In_1458,In_1539);
xor U2484 (N_2484,In_1302,In_2195);
or U2485 (N_2485,In_936,In_120);
and U2486 (N_2486,In_652,In_1711);
or U2487 (N_2487,In_82,In_1975);
and U2488 (N_2488,In_1717,In_1380);
or U2489 (N_2489,In_1742,In_2258);
xor U2490 (N_2490,In_2380,In_1326);
and U2491 (N_2491,In_1197,In_2181);
nor U2492 (N_2492,In_1403,In_215);
nor U2493 (N_2493,In_2122,In_148);
or U2494 (N_2494,In_2244,In_1748);
and U2495 (N_2495,In_888,In_179);
or U2496 (N_2496,In_1632,In_1595);
xnor U2497 (N_2497,In_723,In_1145);
nor U2498 (N_2498,In_676,In_954);
xnor U2499 (N_2499,In_2197,In_2080);
nor U2500 (N_2500,In_1966,In_1828);
or U2501 (N_2501,In_1695,In_1333);
xor U2502 (N_2502,In_184,In_2152);
nand U2503 (N_2503,In_2173,In_2374);
nand U2504 (N_2504,In_1388,In_2158);
nor U2505 (N_2505,In_2384,In_1816);
nand U2506 (N_2506,In_1085,In_734);
nor U2507 (N_2507,In_179,In_1211);
nor U2508 (N_2508,In_1591,In_1139);
or U2509 (N_2509,In_1463,In_2451);
nand U2510 (N_2510,In_1561,In_1026);
nor U2511 (N_2511,In_2398,In_2273);
and U2512 (N_2512,In_428,In_338);
xor U2513 (N_2513,In_650,In_1534);
and U2514 (N_2514,In_1408,In_620);
or U2515 (N_2515,In_1917,In_823);
xor U2516 (N_2516,In_210,In_2385);
nand U2517 (N_2517,In_849,In_938);
and U2518 (N_2518,In_845,In_742);
nand U2519 (N_2519,In_2098,In_2238);
nor U2520 (N_2520,In_2197,In_877);
nand U2521 (N_2521,In_911,In_1186);
or U2522 (N_2522,In_1046,In_916);
and U2523 (N_2523,In_2042,In_1392);
xor U2524 (N_2524,In_384,In_2034);
nor U2525 (N_2525,In_840,In_1020);
and U2526 (N_2526,In_146,In_1164);
or U2527 (N_2527,In_2301,In_2090);
or U2528 (N_2528,In_1767,In_1939);
and U2529 (N_2529,In_975,In_1255);
nor U2530 (N_2530,In_972,In_2068);
and U2531 (N_2531,In_563,In_1232);
nand U2532 (N_2532,In_567,In_2334);
or U2533 (N_2533,In_758,In_1113);
and U2534 (N_2534,In_657,In_2401);
nand U2535 (N_2535,In_1918,In_200);
or U2536 (N_2536,In_1620,In_1276);
nand U2537 (N_2537,In_2173,In_390);
or U2538 (N_2538,In_993,In_1687);
xnor U2539 (N_2539,In_1867,In_2262);
xor U2540 (N_2540,In_1011,In_800);
and U2541 (N_2541,In_1145,In_1766);
nor U2542 (N_2542,In_1602,In_2469);
nor U2543 (N_2543,In_801,In_69);
xnor U2544 (N_2544,In_250,In_881);
or U2545 (N_2545,In_1674,In_301);
nor U2546 (N_2546,In_1295,In_2428);
or U2547 (N_2547,In_33,In_1930);
nor U2548 (N_2548,In_1887,In_1244);
nor U2549 (N_2549,In_360,In_630);
or U2550 (N_2550,In_1126,In_185);
or U2551 (N_2551,In_2002,In_44);
or U2552 (N_2552,In_1601,In_2439);
nand U2553 (N_2553,In_922,In_795);
xnor U2554 (N_2554,In_643,In_904);
or U2555 (N_2555,In_1857,In_1085);
nand U2556 (N_2556,In_2272,In_687);
nand U2557 (N_2557,In_1756,In_413);
and U2558 (N_2558,In_579,In_2190);
or U2559 (N_2559,In_1386,In_264);
nor U2560 (N_2560,In_937,In_1646);
nor U2561 (N_2561,In_1853,In_635);
or U2562 (N_2562,In_1400,In_154);
or U2563 (N_2563,In_681,In_2151);
xnor U2564 (N_2564,In_2037,In_1368);
nand U2565 (N_2565,In_1417,In_1329);
and U2566 (N_2566,In_60,In_66);
xnor U2567 (N_2567,In_733,In_726);
and U2568 (N_2568,In_2447,In_1203);
or U2569 (N_2569,In_1143,In_1603);
and U2570 (N_2570,In_136,In_2267);
nand U2571 (N_2571,In_1352,In_1952);
xor U2572 (N_2572,In_271,In_549);
nand U2573 (N_2573,In_2332,In_2094);
and U2574 (N_2574,In_2135,In_1835);
nand U2575 (N_2575,In_1998,In_1614);
and U2576 (N_2576,In_747,In_1416);
nor U2577 (N_2577,In_2056,In_1408);
and U2578 (N_2578,In_42,In_2454);
and U2579 (N_2579,In_2261,In_2069);
and U2580 (N_2580,In_1244,In_1291);
nor U2581 (N_2581,In_912,In_1990);
xor U2582 (N_2582,In_1506,In_1545);
nor U2583 (N_2583,In_2214,In_2473);
nor U2584 (N_2584,In_1017,In_490);
and U2585 (N_2585,In_1822,In_2160);
nand U2586 (N_2586,In_1496,In_2327);
or U2587 (N_2587,In_669,In_60);
or U2588 (N_2588,In_2439,In_1454);
nor U2589 (N_2589,In_713,In_982);
and U2590 (N_2590,In_1748,In_823);
xor U2591 (N_2591,In_157,In_454);
and U2592 (N_2592,In_2147,In_531);
xnor U2593 (N_2593,In_2284,In_2224);
and U2594 (N_2594,In_445,In_1574);
nand U2595 (N_2595,In_2140,In_779);
nand U2596 (N_2596,In_284,In_2448);
nor U2597 (N_2597,In_1750,In_887);
nor U2598 (N_2598,In_1248,In_2253);
or U2599 (N_2599,In_2095,In_1879);
or U2600 (N_2600,In_649,In_1254);
nor U2601 (N_2601,In_1489,In_105);
nor U2602 (N_2602,In_491,In_1051);
and U2603 (N_2603,In_1912,In_492);
xor U2604 (N_2604,In_211,In_291);
nand U2605 (N_2605,In_1540,In_1259);
nand U2606 (N_2606,In_2007,In_1557);
or U2607 (N_2607,In_356,In_1461);
nor U2608 (N_2608,In_294,In_1239);
nand U2609 (N_2609,In_2015,In_2128);
and U2610 (N_2610,In_1054,In_1605);
xor U2611 (N_2611,In_832,In_1956);
and U2612 (N_2612,In_1868,In_1479);
or U2613 (N_2613,In_2471,In_1512);
nand U2614 (N_2614,In_2095,In_1624);
nor U2615 (N_2615,In_684,In_2195);
or U2616 (N_2616,In_663,In_281);
and U2617 (N_2617,In_2302,In_1813);
nor U2618 (N_2618,In_97,In_1793);
nor U2619 (N_2619,In_227,In_2206);
nand U2620 (N_2620,In_1239,In_1568);
and U2621 (N_2621,In_2186,In_247);
nand U2622 (N_2622,In_902,In_562);
nor U2623 (N_2623,In_174,In_1968);
nand U2624 (N_2624,In_1029,In_2069);
nor U2625 (N_2625,In_1373,In_1797);
and U2626 (N_2626,In_325,In_764);
and U2627 (N_2627,In_1132,In_469);
xor U2628 (N_2628,In_1770,In_2464);
or U2629 (N_2629,In_148,In_1078);
or U2630 (N_2630,In_1110,In_2392);
xor U2631 (N_2631,In_2326,In_1904);
nor U2632 (N_2632,In_928,In_2252);
nand U2633 (N_2633,In_891,In_1746);
or U2634 (N_2634,In_575,In_751);
or U2635 (N_2635,In_1034,In_608);
nand U2636 (N_2636,In_1896,In_2231);
or U2637 (N_2637,In_225,In_1590);
nor U2638 (N_2638,In_1474,In_2297);
and U2639 (N_2639,In_677,In_1134);
and U2640 (N_2640,In_86,In_1796);
and U2641 (N_2641,In_2162,In_1311);
and U2642 (N_2642,In_2308,In_1937);
and U2643 (N_2643,In_517,In_536);
and U2644 (N_2644,In_2052,In_1523);
or U2645 (N_2645,In_931,In_621);
nor U2646 (N_2646,In_35,In_652);
xor U2647 (N_2647,In_1142,In_988);
nand U2648 (N_2648,In_1633,In_917);
or U2649 (N_2649,In_979,In_2183);
nand U2650 (N_2650,In_1064,In_1666);
nand U2651 (N_2651,In_266,In_1083);
nor U2652 (N_2652,In_12,In_968);
xor U2653 (N_2653,In_613,In_2465);
nand U2654 (N_2654,In_981,In_1826);
nand U2655 (N_2655,In_864,In_215);
nor U2656 (N_2656,In_957,In_553);
nor U2657 (N_2657,In_1110,In_1338);
or U2658 (N_2658,In_1886,In_22);
nand U2659 (N_2659,In_1564,In_1761);
and U2660 (N_2660,In_611,In_1934);
or U2661 (N_2661,In_2048,In_1797);
or U2662 (N_2662,In_1108,In_582);
and U2663 (N_2663,In_2122,In_1811);
nand U2664 (N_2664,In_624,In_467);
and U2665 (N_2665,In_1687,In_1331);
nor U2666 (N_2666,In_1161,In_1194);
nor U2667 (N_2667,In_518,In_2402);
or U2668 (N_2668,In_1046,In_1884);
nor U2669 (N_2669,In_710,In_811);
nor U2670 (N_2670,In_62,In_558);
or U2671 (N_2671,In_2343,In_243);
nor U2672 (N_2672,In_1834,In_86);
or U2673 (N_2673,In_1281,In_2158);
and U2674 (N_2674,In_686,In_723);
nor U2675 (N_2675,In_823,In_2074);
nor U2676 (N_2676,In_2101,In_680);
nand U2677 (N_2677,In_591,In_970);
or U2678 (N_2678,In_2378,In_1258);
nand U2679 (N_2679,In_1955,In_1564);
and U2680 (N_2680,In_361,In_1023);
nand U2681 (N_2681,In_2431,In_830);
nand U2682 (N_2682,In_2035,In_2050);
or U2683 (N_2683,In_679,In_1843);
xor U2684 (N_2684,In_69,In_1358);
xnor U2685 (N_2685,In_684,In_124);
and U2686 (N_2686,In_2051,In_1504);
xnor U2687 (N_2687,In_1812,In_640);
xnor U2688 (N_2688,In_2393,In_1047);
or U2689 (N_2689,In_242,In_1192);
and U2690 (N_2690,In_2175,In_2215);
nor U2691 (N_2691,In_282,In_337);
nor U2692 (N_2692,In_2472,In_453);
nor U2693 (N_2693,In_471,In_495);
nand U2694 (N_2694,In_2427,In_822);
nand U2695 (N_2695,In_205,In_894);
nand U2696 (N_2696,In_245,In_535);
xnor U2697 (N_2697,In_1864,In_129);
and U2698 (N_2698,In_2397,In_448);
nor U2699 (N_2699,In_2352,In_1131);
xnor U2700 (N_2700,In_1780,In_2499);
and U2701 (N_2701,In_1377,In_1312);
or U2702 (N_2702,In_1441,In_1595);
or U2703 (N_2703,In_1585,In_2384);
nor U2704 (N_2704,In_1524,In_1631);
nor U2705 (N_2705,In_746,In_239);
nor U2706 (N_2706,In_850,In_1014);
nand U2707 (N_2707,In_2478,In_2027);
nand U2708 (N_2708,In_1582,In_1311);
and U2709 (N_2709,In_1926,In_1203);
and U2710 (N_2710,In_1534,In_861);
or U2711 (N_2711,In_965,In_1047);
nand U2712 (N_2712,In_1388,In_1725);
nand U2713 (N_2713,In_1425,In_276);
nand U2714 (N_2714,In_9,In_2240);
and U2715 (N_2715,In_1381,In_14);
nand U2716 (N_2716,In_1636,In_1611);
nor U2717 (N_2717,In_2070,In_1122);
and U2718 (N_2718,In_1488,In_2491);
nand U2719 (N_2719,In_554,In_1863);
nand U2720 (N_2720,In_1946,In_1614);
nor U2721 (N_2721,In_353,In_1862);
xor U2722 (N_2722,In_1125,In_1235);
nand U2723 (N_2723,In_121,In_161);
or U2724 (N_2724,In_1929,In_2213);
nand U2725 (N_2725,In_17,In_267);
and U2726 (N_2726,In_248,In_1373);
and U2727 (N_2727,In_877,In_304);
nor U2728 (N_2728,In_953,In_2340);
xnor U2729 (N_2729,In_515,In_1407);
nor U2730 (N_2730,In_1114,In_1965);
xnor U2731 (N_2731,In_684,In_1255);
or U2732 (N_2732,In_189,In_1246);
or U2733 (N_2733,In_2416,In_1606);
and U2734 (N_2734,In_1957,In_656);
and U2735 (N_2735,In_1024,In_1542);
nand U2736 (N_2736,In_959,In_1722);
or U2737 (N_2737,In_895,In_2235);
nand U2738 (N_2738,In_1372,In_759);
nor U2739 (N_2739,In_1283,In_371);
xnor U2740 (N_2740,In_1150,In_144);
or U2741 (N_2741,In_440,In_1779);
and U2742 (N_2742,In_661,In_2108);
or U2743 (N_2743,In_1661,In_1813);
nor U2744 (N_2744,In_748,In_1327);
nor U2745 (N_2745,In_568,In_189);
nor U2746 (N_2746,In_1089,In_317);
or U2747 (N_2747,In_2442,In_99);
nand U2748 (N_2748,In_668,In_558);
nor U2749 (N_2749,In_990,In_1146);
xor U2750 (N_2750,In_2254,In_957);
nor U2751 (N_2751,In_1118,In_343);
or U2752 (N_2752,In_1401,In_607);
nand U2753 (N_2753,In_1427,In_971);
and U2754 (N_2754,In_1579,In_202);
and U2755 (N_2755,In_159,In_2122);
or U2756 (N_2756,In_1890,In_832);
and U2757 (N_2757,In_1258,In_570);
nand U2758 (N_2758,In_2148,In_2341);
or U2759 (N_2759,In_1074,In_879);
or U2760 (N_2760,In_1233,In_2196);
and U2761 (N_2761,In_838,In_408);
and U2762 (N_2762,In_1215,In_1983);
nor U2763 (N_2763,In_912,In_1667);
or U2764 (N_2764,In_674,In_1426);
xor U2765 (N_2765,In_1564,In_2057);
nor U2766 (N_2766,In_1124,In_545);
and U2767 (N_2767,In_487,In_1874);
or U2768 (N_2768,In_2160,In_2047);
nand U2769 (N_2769,In_1607,In_1936);
nand U2770 (N_2770,In_2322,In_389);
nor U2771 (N_2771,In_2401,In_1066);
or U2772 (N_2772,In_597,In_1246);
and U2773 (N_2773,In_736,In_795);
and U2774 (N_2774,In_2233,In_104);
xnor U2775 (N_2775,In_501,In_2498);
nand U2776 (N_2776,In_2267,In_1948);
nor U2777 (N_2777,In_1024,In_1029);
xnor U2778 (N_2778,In_1115,In_2172);
nand U2779 (N_2779,In_2496,In_526);
or U2780 (N_2780,In_1946,In_1133);
nand U2781 (N_2781,In_1520,In_2318);
or U2782 (N_2782,In_287,In_1732);
nor U2783 (N_2783,In_1726,In_2444);
nor U2784 (N_2784,In_2020,In_1309);
or U2785 (N_2785,In_149,In_594);
xnor U2786 (N_2786,In_224,In_482);
nand U2787 (N_2787,In_2318,In_874);
or U2788 (N_2788,In_1601,In_1045);
and U2789 (N_2789,In_2053,In_1998);
and U2790 (N_2790,In_1394,In_1266);
nor U2791 (N_2791,In_1088,In_2196);
and U2792 (N_2792,In_1475,In_1197);
nor U2793 (N_2793,In_993,In_1177);
nand U2794 (N_2794,In_2314,In_797);
and U2795 (N_2795,In_778,In_2373);
and U2796 (N_2796,In_2430,In_1370);
nand U2797 (N_2797,In_1076,In_412);
nand U2798 (N_2798,In_1524,In_2003);
or U2799 (N_2799,In_2484,In_1536);
and U2800 (N_2800,In_1303,In_1285);
nand U2801 (N_2801,In_785,In_186);
or U2802 (N_2802,In_2264,In_243);
or U2803 (N_2803,In_1626,In_1019);
nand U2804 (N_2804,In_1587,In_490);
nor U2805 (N_2805,In_1082,In_289);
nor U2806 (N_2806,In_1078,In_973);
nor U2807 (N_2807,In_1913,In_608);
xnor U2808 (N_2808,In_75,In_1278);
xnor U2809 (N_2809,In_358,In_1898);
and U2810 (N_2810,In_1127,In_2322);
nor U2811 (N_2811,In_2402,In_495);
and U2812 (N_2812,In_1098,In_2275);
and U2813 (N_2813,In_1651,In_2209);
nor U2814 (N_2814,In_1325,In_1523);
nand U2815 (N_2815,In_723,In_641);
or U2816 (N_2816,In_2318,In_1786);
xnor U2817 (N_2817,In_1102,In_2472);
xor U2818 (N_2818,In_1694,In_1057);
or U2819 (N_2819,In_1340,In_987);
and U2820 (N_2820,In_861,In_2224);
nand U2821 (N_2821,In_1774,In_2113);
nand U2822 (N_2822,In_721,In_2237);
and U2823 (N_2823,In_1255,In_1758);
or U2824 (N_2824,In_1807,In_2088);
nand U2825 (N_2825,In_1199,In_25);
nand U2826 (N_2826,In_1032,In_1458);
nand U2827 (N_2827,In_735,In_1544);
and U2828 (N_2828,In_1263,In_2360);
xnor U2829 (N_2829,In_1208,In_581);
xnor U2830 (N_2830,In_2449,In_2199);
nand U2831 (N_2831,In_788,In_2303);
and U2832 (N_2832,In_2194,In_392);
nand U2833 (N_2833,In_2041,In_1108);
nor U2834 (N_2834,In_1131,In_1674);
or U2835 (N_2835,In_2133,In_788);
nor U2836 (N_2836,In_814,In_1267);
or U2837 (N_2837,In_1430,In_1273);
nor U2838 (N_2838,In_987,In_1917);
and U2839 (N_2839,In_2225,In_1288);
xnor U2840 (N_2840,In_1469,In_1034);
nor U2841 (N_2841,In_289,In_885);
nor U2842 (N_2842,In_392,In_1031);
nor U2843 (N_2843,In_1257,In_2332);
nor U2844 (N_2844,In_1451,In_1567);
nand U2845 (N_2845,In_2225,In_72);
or U2846 (N_2846,In_480,In_947);
or U2847 (N_2847,In_1878,In_189);
or U2848 (N_2848,In_541,In_886);
or U2849 (N_2849,In_885,In_936);
nand U2850 (N_2850,In_37,In_730);
nand U2851 (N_2851,In_139,In_168);
nand U2852 (N_2852,In_519,In_2444);
or U2853 (N_2853,In_528,In_2220);
and U2854 (N_2854,In_1247,In_2038);
or U2855 (N_2855,In_1027,In_1263);
nor U2856 (N_2856,In_303,In_2465);
and U2857 (N_2857,In_1504,In_1292);
nor U2858 (N_2858,In_1399,In_1820);
and U2859 (N_2859,In_1769,In_2239);
or U2860 (N_2860,In_568,In_1618);
or U2861 (N_2861,In_1260,In_397);
and U2862 (N_2862,In_266,In_324);
nand U2863 (N_2863,In_2304,In_1477);
or U2864 (N_2864,In_814,In_2220);
nor U2865 (N_2865,In_1053,In_1291);
nor U2866 (N_2866,In_2410,In_772);
or U2867 (N_2867,In_1484,In_1372);
and U2868 (N_2868,In_1376,In_364);
nand U2869 (N_2869,In_1458,In_293);
nor U2870 (N_2870,In_1825,In_158);
nor U2871 (N_2871,In_1413,In_1173);
and U2872 (N_2872,In_2019,In_1976);
nor U2873 (N_2873,In_1802,In_840);
nand U2874 (N_2874,In_1394,In_321);
and U2875 (N_2875,In_2452,In_2064);
nand U2876 (N_2876,In_2215,In_1492);
nor U2877 (N_2877,In_332,In_665);
or U2878 (N_2878,In_1657,In_1607);
nor U2879 (N_2879,In_2185,In_239);
nor U2880 (N_2880,In_235,In_1307);
and U2881 (N_2881,In_857,In_527);
and U2882 (N_2882,In_2185,In_1237);
nor U2883 (N_2883,In_316,In_2413);
nor U2884 (N_2884,In_2225,In_233);
and U2885 (N_2885,In_1176,In_1017);
nor U2886 (N_2886,In_516,In_2483);
and U2887 (N_2887,In_1146,In_1553);
nor U2888 (N_2888,In_1341,In_1992);
nand U2889 (N_2889,In_1280,In_2343);
nor U2890 (N_2890,In_1086,In_1412);
and U2891 (N_2891,In_2416,In_1203);
and U2892 (N_2892,In_728,In_722);
and U2893 (N_2893,In_912,In_1959);
and U2894 (N_2894,In_1167,In_1494);
or U2895 (N_2895,In_1614,In_1298);
nand U2896 (N_2896,In_2318,In_157);
and U2897 (N_2897,In_1123,In_1561);
or U2898 (N_2898,In_113,In_2345);
nor U2899 (N_2899,In_94,In_573);
nand U2900 (N_2900,In_2154,In_1001);
or U2901 (N_2901,In_1161,In_1713);
xnor U2902 (N_2902,In_2147,In_2284);
or U2903 (N_2903,In_1777,In_2053);
and U2904 (N_2904,In_875,In_2000);
nor U2905 (N_2905,In_2076,In_1177);
or U2906 (N_2906,In_965,In_891);
and U2907 (N_2907,In_155,In_1816);
and U2908 (N_2908,In_441,In_1902);
nand U2909 (N_2909,In_1751,In_2448);
xor U2910 (N_2910,In_1072,In_716);
nand U2911 (N_2911,In_705,In_154);
nor U2912 (N_2912,In_740,In_2489);
nor U2913 (N_2913,In_607,In_969);
and U2914 (N_2914,In_2068,In_2465);
xor U2915 (N_2915,In_842,In_1089);
and U2916 (N_2916,In_1560,In_671);
nand U2917 (N_2917,In_1313,In_708);
nor U2918 (N_2918,In_557,In_2182);
nor U2919 (N_2919,In_983,In_182);
nor U2920 (N_2920,In_1782,In_899);
xor U2921 (N_2921,In_1626,In_953);
nor U2922 (N_2922,In_2163,In_1744);
and U2923 (N_2923,In_94,In_1842);
nand U2924 (N_2924,In_2301,In_519);
xnor U2925 (N_2925,In_286,In_919);
and U2926 (N_2926,In_1229,In_1084);
nor U2927 (N_2927,In_1635,In_1230);
nor U2928 (N_2928,In_1041,In_1722);
xnor U2929 (N_2929,In_1665,In_1052);
xor U2930 (N_2930,In_1970,In_430);
nand U2931 (N_2931,In_2221,In_609);
nand U2932 (N_2932,In_2083,In_1271);
and U2933 (N_2933,In_484,In_312);
and U2934 (N_2934,In_2443,In_776);
nand U2935 (N_2935,In_1639,In_1051);
and U2936 (N_2936,In_2043,In_266);
nand U2937 (N_2937,In_1402,In_1642);
or U2938 (N_2938,In_1874,In_2229);
or U2939 (N_2939,In_1331,In_1972);
nor U2940 (N_2940,In_1672,In_1171);
xor U2941 (N_2941,In_1746,In_1893);
nand U2942 (N_2942,In_1221,In_2118);
or U2943 (N_2943,In_1541,In_345);
or U2944 (N_2944,In_2173,In_1382);
nand U2945 (N_2945,In_2219,In_2332);
nand U2946 (N_2946,In_192,In_1517);
or U2947 (N_2947,In_412,In_239);
nand U2948 (N_2948,In_420,In_2152);
nor U2949 (N_2949,In_1283,In_1673);
nand U2950 (N_2950,In_623,In_255);
xor U2951 (N_2951,In_1285,In_1611);
nand U2952 (N_2952,In_185,In_1199);
nand U2953 (N_2953,In_1715,In_766);
nor U2954 (N_2954,In_1173,In_1738);
and U2955 (N_2955,In_1546,In_609);
and U2956 (N_2956,In_1054,In_875);
or U2957 (N_2957,In_81,In_2346);
or U2958 (N_2958,In_1145,In_121);
nor U2959 (N_2959,In_1484,In_72);
and U2960 (N_2960,In_544,In_1798);
nor U2961 (N_2961,In_1159,In_2161);
xnor U2962 (N_2962,In_797,In_434);
nor U2963 (N_2963,In_552,In_1426);
xnor U2964 (N_2964,In_1912,In_355);
nand U2965 (N_2965,In_2441,In_1290);
xnor U2966 (N_2966,In_1920,In_1298);
or U2967 (N_2967,In_498,In_1056);
nand U2968 (N_2968,In_2360,In_1544);
nor U2969 (N_2969,In_966,In_361);
nand U2970 (N_2970,In_41,In_187);
or U2971 (N_2971,In_1227,In_248);
nand U2972 (N_2972,In_957,In_1611);
xnor U2973 (N_2973,In_1015,In_872);
nor U2974 (N_2974,In_1214,In_1992);
nor U2975 (N_2975,In_1078,In_2376);
and U2976 (N_2976,In_829,In_1492);
and U2977 (N_2977,In_2277,In_1447);
or U2978 (N_2978,In_1932,In_2485);
nand U2979 (N_2979,In_2492,In_1573);
nand U2980 (N_2980,In_647,In_2144);
xor U2981 (N_2981,In_317,In_1536);
and U2982 (N_2982,In_972,In_1967);
and U2983 (N_2983,In_1722,In_2253);
xnor U2984 (N_2984,In_800,In_510);
and U2985 (N_2985,In_807,In_245);
nand U2986 (N_2986,In_641,In_2307);
nor U2987 (N_2987,In_140,In_1250);
nor U2988 (N_2988,In_104,In_1222);
nor U2989 (N_2989,In_563,In_1394);
nand U2990 (N_2990,In_1835,In_628);
nor U2991 (N_2991,In_30,In_79);
and U2992 (N_2992,In_2189,In_371);
xnor U2993 (N_2993,In_1845,In_817);
nor U2994 (N_2994,In_776,In_1315);
or U2995 (N_2995,In_970,In_2156);
and U2996 (N_2996,In_2264,In_1359);
and U2997 (N_2997,In_1114,In_312);
xnor U2998 (N_2998,In_628,In_1065);
nor U2999 (N_2999,In_927,In_280);
xnor U3000 (N_3000,In_1038,In_1311);
or U3001 (N_3001,In_1085,In_1376);
nor U3002 (N_3002,In_136,In_606);
or U3003 (N_3003,In_1933,In_1992);
nor U3004 (N_3004,In_2462,In_322);
nand U3005 (N_3005,In_1459,In_1289);
nand U3006 (N_3006,In_1783,In_2087);
or U3007 (N_3007,In_764,In_1713);
nand U3008 (N_3008,In_853,In_1303);
and U3009 (N_3009,In_2216,In_561);
or U3010 (N_3010,In_1408,In_2064);
nand U3011 (N_3011,In_1705,In_2176);
xor U3012 (N_3012,In_2316,In_226);
and U3013 (N_3013,In_2263,In_759);
or U3014 (N_3014,In_1857,In_2274);
nor U3015 (N_3015,In_1339,In_350);
nand U3016 (N_3016,In_2127,In_2169);
and U3017 (N_3017,In_366,In_1646);
and U3018 (N_3018,In_1955,In_2157);
and U3019 (N_3019,In_826,In_976);
xnor U3020 (N_3020,In_1720,In_787);
nor U3021 (N_3021,In_270,In_2222);
nand U3022 (N_3022,In_1408,In_2224);
nand U3023 (N_3023,In_80,In_1188);
and U3024 (N_3024,In_1747,In_2290);
nor U3025 (N_3025,In_2057,In_1291);
or U3026 (N_3026,In_2200,In_2435);
or U3027 (N_3027,In_100,In_816);
nor U3028 (N_3028,In_1928,In_2441);
and U3029 (N_3029,In_663,In_38);
nand U3030 (N_3030,In_1953,In_2303);
nor U3031 (N_3031,In_226,In_582);
nor U3032 (N_3032,In_1336,In_1441);
or U3033 (N_3033,In_1630,In_2326);
nand U3034 (N_3034,In_843,In_2365);
nor U3035 (N_3035,In_802,In_1862);
nand U3036 (N_3036,In_1461,In_137);
or U3037 (N_3037,In_3,In_2091);
and U3038 (N_3038,In_251,In_855);
nor U3039 (N_3039,In_2228,In_820);
and U3040 (N_3040,In_949,In_1667);
and U3041 (N_3041,In_863,In_415);
nand U3042 (N_3042,In_383,In_177);
and U3043 (N_3043,In_489,In_2246);
or U3044 (N_3044,In_1635,In_642);
and U3045 (N_3045,In_948,In_423);
nand U3046 (N_3046,In_1110,In_80);
nor U3047 (N_3047,In_1214,In_219);
xor U3048 (N_3048,In_1979,In_1774);
or U3049 (N_3049,In_1305,In_1571);
nand U3050 (N_3050,In_1599,In_1708);
or U3051 (N_3051,In_1600,In_1790);
and U3052 (N_3052,In_1711,In_732);
and U3053 (N_3053,In_1939,In_936);
or U3054 (N_3054,In_1229,In_46);
xor U3055 (N_3055,In_1818,In_1128);
or U3056 (N_3056,In_1310,In_2205);
nor U3057 (N_3057,In_2013,In_1348);
xor U3058 (N_3058,In_442,In_1668);
nor U3059 (N_3059,In_817,In_1770);
or U3060 (N_3060,In_114,In_815);
or U3061 (N_3061,In_998,In_413);
or U3062 (N_3062,In_364,In_1474);
or U3063 (N_3063,In_442,In_1720);
and U3064 (N_3064,In_2258,In_1037);
and U3065 (N_3065,In_67,In_760);
or U3066 (N_3066,In_1853,In_1758);
or U3067 (N_3067,In_1241,In_1337);
and U3068 (N_3068,In_628,In_2288);
nand U3069 (N_3069,In_1199,In_1176);
nand U3070 (N_3070,In_1987,In_1700);
nor U3071 (N_3071,In_984,In_370);
or U3072 (N_3072,In_2479,In_216);
xnor U3073 (N_3073,In_1757,In_972);
nor U3074 (N_3074,In_118,In_956);
and U3075 (N_3075,In_292,In_286);
and U3076 (N_3076,In_1322,In_1978);
nor U3077 (N_3077,In_269,In_393);
nand U3078 (N_3078,In_479,In_348);
nand U3079 (N_3079,In_346,In_1186);
nor U3080 (N_3080,In_1391,In_2238);
nor U3081 (N_3081,In_884,In_1896);
nor U3082 (N_3082,In_1525,In_929);
xor U3083 (N_3083,In_1793,In_1640);
nand U3084 (N_3084,In_2061,In_2354);
or U3085 (N_3085,In_1220,In_240);
nand U3086 (N_3086,In_108,In_2125);
nor U3087 (N_3087,In_2400,In_141);
or U3088 (N_3088,In_1068,In_641);
nand U3089 (N_3089,In_1705,In_1358);
nand U3090 (N_3090,In_1426,In_575);
nand U3091 (N_3091,In_786,In_35);
or U3092 (N_3092,In_63,In_2302);
or U3093 (N_3093,In_1852,In_2142);
nor U3094 (N_3094,In_1097,In_1468);
and U3095 (N_3095,In_1798,In_579);
nor U3096 (N_3096,In_1825,In_909);
nor U3097 (N_3097,In_2190,In_1146);
or U3098 (N_3098,In_973,In_1697);
nand U3099 (N_3099,In_179,In_408);
or U3100 (N_3100,In_2001,In_2037);
and U3101 (N_3101,In_2094,In_2108);
nand U3102 (N_3102,In_2444,In_1377);
or U3103 (N_3103,In_650,In_764);
nand U3104 (N_3104,In_346,In_67);
and U3105 (N_3105,In_719,In_708);
and U3106 (N_3106,In_2458,In_1901);
and U3107 (N_3107,In_545,In_602);
and U3108 (N_3108,In_186,In_1232);
or U3109 (N_3109,In_883,In_2163);
nand U3110 (N_3110,In_454,In_1037);
and U3111 (N_3111,In_2204,In_1746);
or U3112 (N_3112,In_2437,In_194);
and U3113 (N_3113,In_2020,In_1492);
and U3114 (N_3114,In_1311,In_696);
nand U3115 (N_3115,In_1320,In_2195);
nand U3116 (N_3116,In_2097,In_686);
or U3117 (N_3117,In_1948,In_96);
nand U3118 (N_3118,In_111,In_2051);
nor U3119 (N_3119,In_56,In_1981);
nand U3120 (N_3120,In_871,In_1497);
or U3121 (N_3121,In_903,In_2472);
or U3122 (N_3122,In_219,In_1187);
xnor U3123 (N_3123,In_1389,In_2282);
xnor U3124 (N_3124,In_2151,In_89);
nand U3125 (N_3125,In_2345,In_837);
nor U3126 (N_3126,In_2209,In_1225);
or U3127 (N_3127,In_1451,In_1909);
or U3128 (N_3128,In_2475,In_480);
or U3129 (N_3129,In_1978,In_1945);
or U3130 (N_3130,In_1060,In_745);
nand U3131 (N_3131,In_2489,In_1487);
or U3132 (N_3132,In_1413,In_784);
and U3133 (N_3133,In_2476,In_833);
nand U3134 (N_3134,In_969,In_2177);
nand U3135 (N_3135,In_2054,In_911);
xnor U3136 (N_3136,In_1253,In_1809);
nor U3137 (N_3137,In_2434,In_704);
or U3138 (N_3138,In_169,In_1467);
nor U3139 (N_3139,In_2479,In_949);
nand U3140 (N_3140,In_1665,In_999);
nand U3141 (N_3141,In_2158,In_618);
xnor U3142 (N_3142,In_1270,In_1080);
nand U3143 (N_3143,In_794,In_1316);
or U3144 (N_3144,In_2329,In_1280);
or U3145 (N_3145,In_2277,In_1375);
or U3146 (N_3146,In_1928,In_728);
nand U3147 (N_3147,In_1429,In_1075);
and U3148 (N_3148,In_1566,In_1747);
and U3149 (N_3149,In_1005,In_2227);
nor U3150 (N_3150,In_1611,In_1333);
nand U3151 (N_3151,In_2117,In_1053);
nand U3152 (N_3152,In_444,In_2248);
and U3153 (N_3153,In_2201,In_1948);
nand U3154 (N_3154,In_1187,In_860);
or U3155 (N_3155,In_2245,In_2007);
or U3156 (N_3156,In_415,In_2382);
or U3157 (N_3157,In_1350,In_453);
and U3158 (N_3158,In_941,In_712);
xor U3159 (N_3159,In_533,In_996);
and U3160 (N_3160,In_1825,In_1053);
nand U3161 (N_3161,In_1314,In_2431);
and U3162 (N_3162,In_774,In_841);
nor U3163 (N_3163,In_1965,In_2009);
nor U3164 (N_3164,In_2054,In_1067);
nor U3165 (N_3165,In_1291,In_1701);
nor U3166 (N_3166,In_442,In_2412);
or U3167 (N_3167,In_1967,In_799);
nor U3168 (N_3168,In_1148,In_222);
and U3169 (N_3169,In_1852,In_1424);
nand U3170 (N_3170,In_1991,In_1782);
nand U3171 (N_3171,In_758,In_1485);
nor U3172 (N_3172,In_92,In_539);
nor U3173 (N_3173,In_260,In_2141);
xor U3174 (N_3174,In_746,In_794);
and U3175 (N_3175,In_1494,In_117);
xor U3176 (N_3176,In_2372,In_663);
or U3177 (N_3177,In_594,In_1064);
and U3178 (N_3178,In_1634,In_557);
nand U3179 (N_3179,In_1116,In_1884);
nor U3180 (N_3180,In_1504,In_1319);
nor U3181 (N_3181,In_476,In_2395);
or U3182 (N_3182,In_2153,In_1569);
nor U3183 (N_3183,In_2125,In_179);
nand U3184 (N_3184,In_1433,In_1520);
and U3185 (N_3185,In_972,In_1516);
and U3186 (N_3186,In_934,In_2138);
nand U3187 (N_3187,In_2173,In_1940);
and U3188 (N_3188,In_1890,In_50);
or U3189 (N_3189,In_1459,In_1403);
xor U3190 (N_3190,In_148,In_2242);
nor U3191 (N_3191,In_1993,In_1575);
nand U3192 (N_3192,In_1778,In_1409);
or U3193 (N_3193,In_2074,In_1019);
and U3194 (N_3194,In_405,In_632);
xor U3195 (N_3195,In_1158,In_238);
and U3196 (N_3196,In_1571,In_1460);
nand U3197 (N_3197,In_1367,In_1918);
nand U3198 (N_3198,In_537,In_2350);
and U3199 (N_3199,In_1470,In_2079);
nand U3200 (N_3200,In_1875,In_81);
or U3201 (N_3201,In_417,In_1548);
nor U3202 (N_3202,In_1589,In_985);
nand U3203 (N_3203,In_123,In_2410);
and U3204 (N_3204,In_1738,In_139);
nor U3205 (N_3205,In_1518,In_1931);
nor U3206 (N_3206,In_1807,In_305);
nand U3207 (N_3207,In_2002,In_1363);
nand U3208 (N_3208,In_1057,In_150);
and U3209 (N_3209,In_1955,In_1862);
nor U3210 (N_3210,In_1581,In_849);
nor U3211 (N_3211,In_98,In_1688);
xnor U3212 (N_3212,In_1545,In_161);
xor U3213 (N_3213,In_200,In_1236);
or U3214 (N_3214,In_2354,In_1715);
and U3215 (N_3215,In_138,In_1787);
nand U3216 (N_3216,In_1841,In_676);
xnor U3217 (N_3217,In_722,In_559);
or U3218 (N_3218,In_112,In_632);
nor U3219 (N_3219,In_2291,In_414);
nand U3220 (N_3220,In_1819,In_1269);
xnor U3221 (N_3221,In_657,In_2264);
nand U3222 (N_3222,In_418,In_982);
and U3223 (N_3223,In_748,In_1232);
or U3224 (N_3224,In_1081,In_1405);
xnor U3225 (N_3225,In_942,In_1990);
or U3226 (N_3226,In_1951,In_644);
nand U3227 (N_3227,In_1760,In_810);
nor U3228 (N_3228,In_283,In_1559);
and U3229 (N_3229,In_1515,In_218);
nand U3230 (N_3230,In_517,In_1023);
nor U3231 (N_3231,In_1297,In_934);
nand U3232 (N_3232,In_528,In_1466);
xor U3233 (N_3233,In_2141,In_141);
nor U3234 (N_3234,In_57,In_840);
and U3235 (N_3235,In_1092,In_2406);
xnor U3236 (N_3236,In_462,In_1070);
and U3237 (N_3237,In_2493,In_2148);
and U3238 (N_3238,In_1416,In_1604);
xor U3239 (N_3239,In_306,In_2197);
nand U3240 (N_3240,In_1306,In_666);
and U3241 (N_3241,In_173,In_1792);
nor U3242 (N_3242,In_214,In_1450);
xnor U3243 (N_3243,In_1847,In_812);
nor U3244 (N_3244,In_1958,In_805);
nor U3245 (N_3245,In_2196,In_1799);
or U3246 (N_3246,In_1688,In_523);
nor U3247 (N_3247,In_1801,In_2056);
nand U3248 (N_3248,In_1450,In_1788);
nand U3249 (N_3249,In_827,In_1213);
nand U3250 (N_3250,In_1887,In_2078);
xor U3251 (N_3251,In_97,In_2322);
and U3252 (N_3252,In_2043,In_409);
nor U3253 (N_3253,In_341,In_1900);
nor U3254 (N_3254,In_1512,In_941);
nor U3255 (N_3255,In_794,In_22);
nor U3256 (N_3256,In_744,In_998);
nand U3257 (N_3257,In_628,In_2478);
nor U3258 (N_3258,In_1537,In_614);
xor U3259 (N_3259,In_679,In_1745);
nand U3260 (N_3260,In_1385,In_161);
and U3261 (N_3261,In_1900,In_290);
nand U3262 (N_3262,In_1044,In_496);
xnor U3263 (N_3263,In_1532,In_2156);
nand U3264 (N_3264,In_139,In_924);
or U3265 (N_3265,In_1320,In_2124);
nor U3266 (N_3266,In_1794,In_2144);
nor U3267 (N_3267,In_1927,In_775);
nand U3268 (N_3268,In_147,In_1665);
and U3269 (N_3269,In_1812,In_972);
nand U3270 (N_3270,In_634,In_982);
or U3271 (N_3271,In_47,In_1482);
nor U3272 (N_3272,In_641,In_139);
xor U3273 (N_3273,In_306,In_1965);
or U3274 (N_3274,In_1743,In_1871);
nor U3275 (N_3275,In_1034,In_1785);
and U3276 (N_3276,In_907,In_1186);
nand U3277 (N_3277,In_1322,In_2249);
or U3278 (N_3278,In_489,In_177);
nand U3279 (N_3279,In_142,In_828);
nor U3280 (N_3280,In_1409,In_1078);
nor U3281 (N_3281,In_199,In_1759);
nor U3282 (N_3282,In_101,In_1098);
xnor U3283 (N_3283,In_2241,In_230);
xnor U3284 (N_3284,In_1498,In_321);
nor U3285 (N_3285,In_479,In_553);
nand U3286 (N_3286,In_176,In_638);
and U3287 (N_3287,In_983,In_2276);
and U3288 (N_3288,In_277,In_1259);
nand U3289 (N_3289,In_2361,In_366);
or U3290 (N_3290,In_1879,In_2270);
nand U3291 (N_3291,In_583,In_2098);
nand U3292 (N_3292,In_581,In_1303);
xor U3293 (N_3293,In_989,In_1252);
xor U3294 (N_3294,In_1664,In_1662);
nor U3295 (N_3295,In_2257,In_1226);
and U3296 (N_3296,In_2159,In_2413);
nand U3297 (N_3297,In_1211,In_1568);
nand U3298 (N_3298,In_213,In_1716);
or U3299 (N_3299,In_1182,In_2248);
nand U3300 (N_3300,In_453,In_2296);
and U3301 (N_3301,In_2012,In_338);
nand U3302 (N_3302,In_2352,In_1315);
nor U3303 (N_3303,In_1512,In_2274);
or U3304 (N_3304,In_2125,In_1017);
or U3305 (N_3305,In_954,In_509);
or U3306 (N_3306,In_1019,In_152);
xor U3307 (N_3307,In_2094,In_1022);
and U3308 (N_3308,In_1570,In_1063);
nand U3309 (N_3309,In_2333,In_1052);
xor U3310 (N_3310,In_2341,In_788);
nor U3311 (N_3311,In_460,In_503);
or U3312 (N_3312,In_2022,In_1163);
nand U3313 (N_3313,In_2129,In_728);
nand U3314 (N_3314,In_365,In_329);
or U3315 (N_3315,In_2171,In_2089);
nand U3316 (N_3316,In_50,In_533);
nand U3317 (N_3317,In_1974,In_150);
and U3318 (N_3318,In_1671,In_626);
nand U3319 (N_3319,In_2113,In_525);
and U3320 (N_3320,In_1706,In_112);
or U3321 (N_3321,In_586,In_403);
or U3322 (N_3322,In_1426,In_2388);
nor U3323 (N_3323,In_2241,In_13);
nor U3324 (N_3324,In_1277,In_1347);
nor U3325 (N_3325,In_655,In_216);
or U3326 (N_3326,In_2080,In_2400);
or U3327 (N_3327,In_2437,In_1667);
and U3328 (N_3328,In_1525,In_2114);
or U3329 (N_3329,In_979,In_2338);
nand U3330 (N_3330,In_170,In_1753);
nand U3331 (N_3331,In_1178,In_845);
and U3332 (N_3332,In_199,In_346);
nor U3333 (N_3333,In_1809,In_715);
nand U3334 (N_3334,In_758,In_1039);
or U3335 (N_3335,In_1576,In_2362);
nor U3336 (N_3336,In_338,In_2330);
nor U3337 (N_3337,In_2480,In_1981);
and U3338 (N_3338,In_793,In_2374);
nor U3339 (N_3339,In_347,In_2287);
nor U3340 (N_3340,In_29,In_2076);
nor U3341 (N_3341,In_2382,In_2103);
nand U3342 (N_3342,In_939,In_1163);
or U3343 (N_3343,In_1216,In_1135);
or U3344 (N_3344,In_1628,In_177);
nor U3345 (N_3345,In_399,In_763);
nand U3346 (N_3346,In_2266,In_832);
nor U3347 (N_3347,In_59,In_683);
xor U3348 (N_3348,In_940,In_2207);
and U3349 (N_3349,In_1283,In_972);
nand U3350 (N_3350,In_1490,In_1548);
or U3351 (N_3351,In_537,In_1150);
nand U3352 (N_3352,In_631,In_2033);
or U3353 (N_3353,In_1067,In_175);
nand U3354 (N_3354,In_393,In_832);
nor U3355 (N_3355,In_1132,In_1702);
and U3356 (N_3356,In_1945,In_1306);
or U3357 (N_3357,In_916,In_2454);
and U3358 (N_3358,In_2208,In_2087);
nand U3359 (N_3359,In_2030,In_2050);
and U3360 (N_3360,In_198,In_1363);
nand U3361 (N_3361,In_1466,In_51);
or U3362 (N_3362,In_2233,In_1009);
nor U3363 (N_3363,In_1332,In_2017);
or U3364 (N_3364,In_302,In_1943);
and U3365 (N_3365,In_1362,In_25);
or U3366 (N_3366,In_1509,In_886);
and U3367 (N_3367,In_1216,In_205);
nand U3368 (N_3368,In_1643,In_112);
nand U3369 (N_3369,In_1032,In_613);
nor U3370 (N_3370,In_84,In_282);
nor U3371 (N_3371,In_487,In_311);
xor U3372 (N_3372,In_2125,In_2306);
nor U3373 (N_3373,In_870,In_1154);
or U3374 (N_3374,In_1259,In_1526);
nor U3375 (N_3375,In_1721,In_226);
xor U3376 (N_3376,In_2302,In_1111);
or U3377 (N_3377,In_928,In_322);
nor U3378 (N_3378,In_707,In_2141);
nor U3379 (N_3379,In_83,In_2005);
nor U3380 (N_3380,In_1055,In_239);
or U3381 (N_3381,In_2378,In_1491);
nor U3382 (N_3382,In_2274,In_1933);
or U3383 (N_3383,In_2180,In_1012);
xor U3384 (N_3384,In_1788,In_1044);
nand U3385 (N_3385,In_2013,In_84);
or U3386 (N_3386,In_1742,In_1508);
nor U3387 (N_3387,In_472,In_2063);
and U3388 (N_3388,In_1873,In_1789);
and U3389 (N_3389,In_2254,In_1000);
nor U3390 (N_3390,In_924,In_1209);
nor U3391 (N_3391,In_1690,In_1200);
and U3392 (N_3392,In_854,In_1386);
and U3393 (N_3393,In_1214,In_1829);
and U3394 (N_3394,In_1978,In_962);
and U3395 (N_3395,In_1871,In_563);
and U3396 (N_3396,In_2241,In_731);
and U3397 (N_3397,In_1784,In_2293);
nand U3398 (N_3398,In_2176,In_474);
nor U3399 (N_3399,In_141,In_2027);
nor U3400 (N_3400,In_1581,In_92);
nor U3401 (N_3401,In_539,In_2096);
xor U3402 (N_3402,In_1213,In_2215);
xnor U3403 (N_3403,In_2180,In_2219);
and U3404 (N_3404,In_780,In_788);
nor U3405 (N_3405,In_927,In_214);
or U3406 (N_3406,In_627,In_1726);
nand U3407 (N_3407,In_2352,In_1088);
nand U3408 (N_3408,In_613,In_2400);
or U3409 (N_3409,In_1437,In_1392);
and U3410 (N_3410,In_1284,In_1258);
xnor U3411 (N_3411,In_1839,In_509);
nand U3412 (N_3412,In_2119,In_2020);
nor U3413 (N_3413,In_1955,In_1339);
and U3414 (N_3414,In_1185,In_2202);
or U3415 (N_3415,In_2293,In_932);
or U3416 (N_3416,In_2352,In_795);
and U3417 (N_3417,In_1514,In_2081);
nand U3418 (N_3418,In_1181,In_1403);
or U3419 (N_3419,In_795,In_732);
nor U3420 (N_3420,In_973,In_758);
nand U3421 (N_3421,In_541,In_1487);
or U3422 (N_3422,In_1958,In_1035);
nor U3423 (N_3423,In_1012,In_1135);
nor U3424 (N_3424,In_472,In_400);
nor U3425 (N_3425,In_1452,In_741);
or U3426 (N_3426,In_336,In_1154);
xor U3427 (N_3427,In_1640,In_1650);
nand U3428 (N_3428,In_353,In_2348);
and U3429 (N_3429,In_2462,In_2449);
nand U3430 (N_3430,In_1755,In_1543);
nand U3431 (N_3431,In_2406,In_2255);
and U3432 (N_3432,In_1753,In_1171);
nor U3433 (N_3433,In_547,In_2138);
nand U3434 (N_3434,In_692,In_352);
or U3435 (N_3435,In_2168,In_248);
xnor U3436 (N_3436,In_1866,In_1711);
nand U3437 (N_3437,In_878,In_801);
and U3438 (N_3438,In_1234,In_433);
nor U3439 (N_3439,In_1379,In_744);
nor U3440 (N_3440,In_922,In_2347);
or U3441 (N_3441,In_2141,In_1454);
nand U3442 (N_3442,In_1666,In_1987);
nand U3443 (N_3443,In_1073,In_2267);
nor U3444 (N_3444,In_1389,In_69);
and U3445 (N_3445,In_259,In_73);
nand U3446 (N_3446,In_1495,In_958);
nand U3447 (N_3447,In_1124,In_1784);
nand U3448 (N_3448,In_681,In_1553);
nand U3449 (N_3449,In_1559,In_1904);
xor U3450 (N_3450,In_2128,In_936);
nand U3451 (N_3451,In_487,In_1721);
and U3452 (N_3452,In_2180,In_1408);
or U3453 (N_3453,In_1577,In_1160);
or U3454 (N_3454,In_548,In_2295);
nor U3455 (N_3455,In_426,In_278);
and U3456 (N_3456,In_613,In_2132);
xnor U3457 (N_3457,In_447,In_67);
nand U3458 (N_3458,In_1851,In_520);
or U3459 (N_3459,In_643,In_1998);
or U3460 (N_3460,In_2107,In_1753);
xnor U3461 (N_3461,In_957,In_2133);
nor U3462 (N_3462,In_504,In_2462);
nand U3463 (N_3463,In_1441,In_505);
nor U3464 (N_3464,In_167,In_2323);
or U3465 (N_3465,In_592,In_1572);
or U3466 (N_3466,In_2029,In_2138);
nand U3467 (N_3467,In_1211,In_1275);
nand U3468 (N_3468,In_115,In_1178);
and U3469 (N_3469,In_1379,In_656);
nor U3470 (N_3470,In_2268,In_454);
xor U3471 (N_3471,In_907,In_939);
xnor U3472 (N_3472,In_314,In_1172);
and U3473 (N_3473,In_1562,In_2052);
and U3474 (N_3474,In_583,In_192);
and U3475 (N_3475,In_1695,In_1142);
nor U3476 (N_3476,In_2147,In_1441);
and U3477 (N_3477,In_1603,In_2143);
or U3478 (N_3478,In_654,In_499);
and U3479 (N_3479,In_1034,In_1794);
nor U3480 (N_3480,In_391,In_1480);
nor U3481 (N_3481,In_1094,In_2060);
and U3482 (N_3482,In_1156,In_94);
nor U3483 (N_3483,In_1454,In_1116);
nor U3484 (N_3484,In_335,In_169);
or U3485 (N_3485,In_2064,In_912);
nor U3486 (N_3486,In_198,In_1624);
and U3487 (N_3487,In_811,In_2496);
nor U3488 (N_3488,In_736,In_1182);
nand U3489 (N_3489,In_894,In_449);
or U3490 (N_3490,In_786,In_1804);
xor U3491 (N_3491,In_332,In_1839);
nand U3492 (N_3492,In_1108,In_1194);
or U3493 (N_3493,In_671,In_2358);
nand U3494 (N_3494,In_89,In_814);
or U3495 (N_3495,In_1159,In_1609);
xnor U3496 (N_3496,In_157,In_241);
and U3497 (N_3497,In_2390,In_1808);
or U3498 (N_3498,In_1605,In_337);
and U3499 (N_3499,In_347,In_1077);
or U3500 (N_3500,In_588,In_498);
xnor U3501 (N_3501,In_2243,In_1809);
or U3502 (N_3502,In_1720,In_2207);
nand U3503 (N_3503,In_1361,In_1394);
nand U3504 (N_3504,In_2487,In_1226);
or U3505 (N_3505,In_151,In_887);
nand U3506 (N_3506,In_540,In_1986);
or U3507 (N_3507,In_958,In_668);
nand U3508 (N_3508,In_1380,In_1151);
nand U3509 (N_3509,In_1595,In_2416);
nand U3510 (N_3510,In_633,In_1116);
nand U3511 (N_3511,In_2447,In_672);
and U3512 (N_3512,In_907,In_2347);
nor U3513 (N_3513,In_14,In_1880);
xnor U3514 (N_3514,In_2026,In_1013);
and U3515 (N_3515,In_504,In_805);
and U3516 (N_3516,In_2346,In_1961);
nor U3517 (N_3517,In_1156,In_1291);
or U3518 (N_3518,In_1397,In_1659);
xnor U3519 (N_3519,In_2230,In_156);
or U3520 (N_3520,In_2145,In_1529);
xnor U3521 (N_3521,In_140,In_658);
or U3522 (N_3522,In_686,In_1656);
nand U3523 (N_3523,In_106,In_595);
nor U3524 (N_3524,In_767,In_375);
nor U3525 (N_3525,In_2203,In_1808);
nand U3526 (N_3526,In_2294,In_816);
or U3527 (N_3527,In_482,In_1336);
nand U3528 (N_3528,In_1257,In_1934);
or U3529 (N_3529,In_2281,In_2175);
and U3530 (N_3530,In_137,In_1442);
nand U3531 (N_3531,In_1493,In_820);
nand U3532 (N_3532,In_1220,In_2361);
nand U3533 (N_3533,In_874,In_2398);
or U3534 (N_3534,In_2356,In_1019);
or U3535 (N_3535,In_712,In_1859);
nand U3536 (N_3536,In_2356,In_1453);
and U3537 (N_3537,In_2068,In_185);
and U3538 (N_3538,In_492,In_2090);
nor U3539 (N_3539,In_949,In_2068);
nand U3540 (N_3540,In_2305,In_126);
or U3541 (N_3541,In_2321,In_172);
and U3542 (N_3542,In_1913,In_41);
xor U3543 (N_3543,In_45,In_257);
nor U3544 (N_3544,In_1891,In_289);
nand U3545 (N_3545,In_997,In_514);
and U3546 (N_3546,In_1675,In_240);
nor U3547 (N_3547,In_103,In_261);
nand U3548 (N_3548,In_1030,In_201);
or U3549 (N_3549,In_207,In_716);
xnor U3550 (N_3550,In_2144,In_2399);
xnor U3551 (N_3551,In_707,In_1670);
or U3552 (N_3552,In_1211,In_1368);
nor U3553 (N_3553,In_360,In_1805);
xnor U3554 (N_3554,In_410,In_1224);
nand U3555 (N_3555,In_243,In_208);
xnor U3556 (N_3556,In_2151,In_456);
and U3557 (N_3557,In_2108,In_1440);
and U3558 (N_3558,In_2121,In_565);
nand U3559 (N_3559,In_769,In_815);
nand U3560 (N_3560,In_957,In_889);
and U3561 (N_3561,In_119,In_856);
nor U3562 (N_3562,In_348,In_2171);
and U3563 (N_3563,In_2351,In_1728);
nand U3564 (N_3564,In_1889,In_2128);
xnor U3565 (N_3565,In_1324,In_566);
and U3566 (N_3566,In_2213,In_57);
or U3567 (N_3567,In_1406,In_1787);
nand U3568 (N_3568,In_943,In_70);
nor U3569 (N_3569,In_1051,In_898);
nand U3570 (N_3570,In_2204,In_2127);
and U3571 (N_3571,In_403,In_1447);
nor U3572 (N_3572,In_1814,In_2135);
and U3573 (N_3573,In_269,In_856);
nand U3574 (N_3574,In_1263,In_1571);
or U3575 (N_3575,In_768,In_628);
nand U3576 (N_3576,In_2159,In_372);
nand U3577 (N_3577,In_854,In_674);
or U3578 (N_3578,In_804,In_387);
nand U3579 (N_3579,In_1397,In_891);
xor U3580 (N_3580,In_1085,In_399);
nand U3581 (N_3581,In_1290,In_917);
and U3582 (N_3582,In_1931,In_105);
and U3583 (N_3583,In_1549,In_1093);
and U3584 (N_3584,In_2429,In_2057);
nor U3585 (N_3585,In_2490,In_1104);
nor U3586 (N_3586,In_1922,In_1794);
or U3587 (N_3587,In_1168,In_2090);
and U3588 (N_3588,In_2209,In_1322);
nand U3589 (N_3589,In_1682,In_371);
nor U3590 (N_3590,In_119,In_871);
or U3591 (N_3591,In_1756,In_738);
and U3592 (N_3592,In_1558,In_131);
xnor U3593 (N_3593,In_1096,In_2248);
nor U3594 (N_3594,In_401,In_1063);
and U3595 (N_3595,In_455,In_87);
nand U3596 (N_3596,In_1292,In_581);
nand U3597 (N_3597,In_582,In_1218);
or U3598 (N_3598,In_1598,In_2056);
or U3599 (N_3599,In_2268,In_327);
nor U3600 (N_3600,In_2367,In_961);
and U3601 (N_3601,In_1067,In_1622);
xnor U3602 (N_3602,In_1022,In_96);
nor U3603 (N_3603,In_612,In_1046);
or U3604 (N_3604,In_164,In_1278);
nor U3605 (N_3605,In_1568,In_1296);
and U3606 (N_3606,In_75,In_1235);
nand U3607 (N_3607,In_2429,In_1600);
or U3608 (N_3608,In_856,In_1877);
nand U3609 (N_3609,In_1266,In_1306);
nor U3610 (N_3610,In_839,In_2391);
xnor U3611 (N_3611,In_106,In_1952);
and U3612 (N_3612,In_447,In_1202);
nand U3613 (N_3613,In_909,In_1869);
nand U3614 (N_3614,In_1700,In_1812);
or U3615 (N_3615,In_2332,In_1554);
nor U3616 (N_3616,In_1976,In_2189);
and U3617 (N_3617,In_2309,In_2479);
and U3618 (N_3618,In_973,In_692);
xnor U3619 (N_3619,In_2136,In_924);
nand U3620 (N_3620,In_991,In_447);
nand U3621 (N_3621,In_848,In_327);
or U3622 (N_3622,In_2145,In_1057);
nand U3623 (N_3623,In_2038,In_56);
nor U3624 (N_3624,In_1342,In_1553);
xor U3625 (N_3625,In_758,In_1820);
and U3626 (N_3626,In_91,In_2135);
or U3627 (N_3627,In_596,In_77);
or U3628 (N_3628,In_2137,In_2352);
and U3629 (N_3629,In_657,In_904);
nor U3630 (N_3630,In_1883,In_852);
nand U3631 (N_3631,In_1946,In_1163);
nor U3632 (N_3632,In_419,In_551);
or U3633 (N_3633,In_1070,In_1554);
nand U3634 (N_3634,In_798,In_1402);
and U3635 (N_3635,In_1581,In_1418);
or U3636 (N_3636,In_1030,In_2300);
nor U3637 (N_3637,In_961,In_849);
nor U3638 (N_3638,In_1867,In_435);
and U3639 (N_3639,In_2239,In_646);
xnor U3640 (N_3640,In_1755,In_1551);
and U3641 (N_3641,In_1750,In_1198);
and U3642 (N_3642,In_2463,In_1874);
nand U3643 (N_3643,In_1022,In_712);
or U3644 (N_3644,In_1389,In_337);
nand U3645 (N_3645,In_1726,In_1510);
and U3646 (N_3646,In_2339,In_900);
nor U3647 (N_3647,In_1888,In_36);
nand U3648 (N_3648,In_2082,In_1850);
xor U3649 (N_3649,In_2262,In_1323);
nor U3650 (N_3650,In_1890,In_1627);
and U3651 (N_3651,In_1706,In_811);
nor U3652 (N_3652,In_1246,In_2000);
nor U3653 (N_3653,In_2343,In_948);
or U3654 (N_3654,In_1497,In_2421);
or U3655 (N_3655,In_1730,In_1874);
or U3656 (N_3656,In_781,In_1067);
nand U3657 (N_3657,In_1572,In_54);
or U3658 (N_3658,In_1714,In_839);
xnor U3659 (N_3659,In_813,In_334);
or U3660 (N_3660,In_85,In_2057);
nor U3661 (N_3661,In_478,In_195);
nor U3662 (N_3662,In_2457,In_783);
and U3663 (N_3663,In_2140,In_671);
and U3664 (N_3664,In_155,In_2028);
or U3665 (N_3665,In_875,In_68);
nand U3666 (N_3666,In_2207,In_1153);
and U3667 (N_3667,In_646,In_878);
nand U3668 (N_3668,In_2113,In_578);
nand U3669 (N_3669,In_358,In_309);
nor U3670 (N_3670,In_1462,In_1849);
nand U3671 (N_3671,In_1558,In_309);
nand U3672 (N_3672,In_1244,In_2124);
xnor U3673 (N_3673,In_1080,In_145);
nand U3674 (N_3674,In_1178,In_946);
xor U3675 (N_3675,In_613,In_1528);
and U3676 (N_3676,In_1065,In_2038);
and U3677 (N_3677,In_2293,In_1147);
xnor U3678 (N_3678,In_359,In_1782);
or U3679 (N_3679,In_2256,In_1954);
xor U3680 (N_3680,In_363,In_49);
and U3681 (N_3681,In_1729,In_52);
xnor U3682 (N_3682,In_1465,In_2353);
and U3683 (N_3683,In_272,In_1218);
or U3684 (N_3684,In_990,In_2374);
and U3685 (N_3685,In_352,In_1483);
or U3686 (N_3686,In_1186,In_2394);
nand U3687 (N_3687,In_59,In_2243);
nor U3688 (N_3688,In_940,In_927);
or U3689 (N_3689,In_1113,In_1862);
nand U3690 (N_3690,In_1883,In_1961);
nor U3691 (N_3691,In_1525,In_589);
nand U3692 (N_3692,In_1285,In_565);
nand U3693 (N_3693,In_1744,In_2395);
or U3694 (N_3694,In_1137,In_1604);
and U3695 (N_3695,In_1760,In_9);
or U3696 (N_3696,In_2190,In_1448);
nand U3697 (N_3697,In_161,In_249);
nand U3698 (N_3698,In_1828,In_369);
nor U3699 (N_3699,In_255,In_289);
nand U3700 (N_3700,In_1055,In_1474);
nor U3701 (N_3701,In_1345,In_1261);
and U3702 (N_3702,In_25,In_1196);
nand U3703 (N_3703,In_1164,In_1250);
and U3704 (N_3704,In_536,In_2251);
and U3705 (N_3705,In_1569,In_183);
nand U3706 (N_3706,In_1986,In_617);
nand U3707 (N_3707,In_1740,In_1951);
or U3708 (N_3708,In_1449,In_1443);
nand U3709 (N_3709,In_565,In_1369);
or U3710 (N_3710,In_2466,In_2374);
and U3711 (N_3711,In_1130,In_2359);
nand U3712 (N_3712,In_130,In_1134);
and U3713 (N_3713,In_99,In_348);
nand U3714 (N_3714,In_700,In_2099);
or U3715 (N_3715,In_1610,In_8);
xnor U3716 (N_3716,In_1935,In_1970);
nor U3717 (N_3717,In_657,In_774);
and U3718 (N_3718,In_678,In_2295);
nor U3719 (N_3719,In_1673,In_1178);
and U3720 (N_3720,In_1055,In_1241);
nand U3721 (N_3721,In_1998,In_1937);
or U3722 (N_3722,In_2204,In_402);
or U3723 (N_3723,In_178,In_776);
or U3724 (N_3724,In_2467,In_1048);
nor U3725 (N_3725,In_984,In_971);
and U3726 (N_3726,In_496,In_1399);
or U3727 (N_3727,In_1138,In_274);
nand U3728 (N_3728,In_647,In_835);
or U3729 (N_3729,In_592,In_2131);
xor U3730 (N_3730,In_91,In_2471);
and U3731 (N_3731,In_1119,In_2042);
nand U3732 (N_3732,In_2013,In_1368);
or U3733 (N_3733,In_1490,In_2247);
and U3734 (N_3734,In_877,In_2190);
and U3735 (N_3735,In_226,In_2143);
or U3736 (N_3736,In_935,In_20);
xnor U3737 (N_3737,In_2303,In_2416);
nand U3738 (N_3738,In_2238,In_1513);
and U3739 (N_3739,In_1277,In_1150);
xor U3740 (N_3740,In_606,In_2455);
nand U3741 (N_3741,In_1365,In_608);
or U3742 (N_3742,In_1750,In_1814);
nand U3743 (N_3743,In_379,In_2313);
or U3744 (N_3744,In_92,In_1242);
and U3745 (N_3745,In_2122,In_221);
or U3746 (N_3746,In_1973,In_777);
nor U3747 (N_3747,In_1840,In_1798);
or U3748 (N_3748,In_169,In_520);
nand U3749 (N_3749,In_167,In_1242);
or U3750 (N_3750,In_1917,In_1633);
nand U3751 (N_3751,In_2043,In_281);
nand U3752 (N_3752,In_1962,In_316);
nor U3753 (N_3753,In_2118,In_40);
or U3754 (N_3754,In_2004,In_275);
and U3755 (N_3755,In_542,In_2202);
nand U3756 (N_3756,In_523,In_992);
xnor U3757 (N_3757,In_1009,In_1562);
or U3758 (N_3758,In_294,In_1152);
and U3759 (N_3759,In_203,In_1466);
and U3760 (N_3760,In_905,In_1049);
xor U3761 (N_3761,In_1777,In_1001);
nand U3762 (N_3762,In_2133,In_213);
nand U3763 (N_3763,In_2080,In_2325);
or U3764 (N_3764,In_2424,In_833);
xnor U3765 (N_3765,In_1735,In_1244);
nor U3766 (N_3766,In_2242,In_1438);
or U3767 (N_3767,In_858,In_1887);
and U3768 (N_3768,In_1676,In_1864);
nor U3769 (N_3769,In_1038,In_281);
or U3770 (N_3770,In_254,In_2483);
nand U3771 (N_3771,In_1904,In_924);
nand U3772 (N_3772,In_1308,In_1202);
nand U3773 (N_3773,In_1947,In_1370);
or U3774 (N_3774,In_2478,In_533);
or U3775 (N_3775,In_1159,In_555);
nand U3776 (N_3776,In_2083,In_1517);
and U3777 (N_3777,In_615,In_729);
or U3778 (N_3778,In_499,In_2074);
or U3779 (N_3779,In_2002,In_1470);
and U3780 (N_3780,In_1320,In_994);
nor U3781 (N_3781,In_1210,In_1321);
and U3782 (N_3782,In_600,In_734);
nor U3783 (N_3783,In_1000,In_247);
or U3784 (N_3784,In_2089,In_164);
or U3785 (N_3785,In_1421,In_568);
nand U3786 (N_3786,In_1370,In_1953);
nor U3787 (N_3787,In_1569,In_1711);
nor U3788 (N_3788,In_2460,In_609);
nor U3789 (N_3789,In_1122,In_1984);
and U3790 (N_3790,In_1831,In_442);
xor U3791 (N_3791,In_1954,In_121);
and U3792 (N_3792,In_16,In_606);
nand U3793 (N_3793,In_2365,In_2016);
nor U3794 (N_3794,In_819,In_1277);
nand U3795 (N_3795,In_113,In_1841);
or U3796 (N_3796,In_1292,In_2077);
nor U3797 (N_3797,In_1952,In_1773);
xnor U3798 (N_3798,In_320,In_647);
and U3799 (N_3799,In_878,In_943);
nor U3800 (N_3800,In_2034,In_750);
nand U3801 (N_3801,In_372,In_1763);
or U3802 (N_3802,In_808,In_185);
or U3803 (N_3803,In_1710,In_1657);
xor U3804 (N_3804,In_2434,In_1631);
xnor U3805 (N_3805,In_347,In_1869);
nor U3806 (N_3806,In_1934,In_197);
nand U3807 (N_3807,In_1409,In_2207);
xor U3808 (N_3808,In_547,In_444);
xor U3809 (N_3809,In_521,In_1257);
nor U3810 (N_3810,In_746,In_166);
and U3811 (N_3811,In_1472,In_1759);
nand U3812 (N_3812,In_726,In_252);
xnor U3813 (N_3813,In_2482,In_2322);
nand U3814 (N_3814,In_246,In_1873);
and U3815 (N_3815,In_1407,In_35);
nand U3816 (N_3816,In_1575,In_2327);
or U3817 (N_3817,In_241,In_1909);
and U3818 (N_3818,In_2074,In_1988);
nand U3819 (N_3819,In_211,In_172);
xor U3820 (N_3820,In_1863,In_406);
nor U3821 (N_3821,In_117,In_1616);
and U3822 (N_3822,In_1531,In_853);
or U3823 (N_3823,In_74,In_2139);
and U3824 (N_3824,In_1766,In_2093);
nor U3825 (N_3825,In_1259,In_1809);
and U3826 (N_3826,In_1655,In_288);
and U3827 (N_3827,In_1997,In_1580);
nand U3828 (N_3828,In_2239,In_2192);
xnor U3829 (N_3829,In_2334,In_2345);
xnor U3830 (N_3830,In_660,In_464);
nor U3831 (N_3831,In_1891,In_166);
nand U3832 (N_3832,In_678,In_2275);
nand U3833 (N_3833,In_1092,In_1129);
and U3834 (N_3834,In_69,In_1634);
and U3835 (N_3835,In_697,In_1908);
nand U3836 (N_3836,In_1609,In_1511);
and U3837 (N_3837,In_1602,In_1101);
or U3838 (N_3838,In_1903,In_2041);
and U3839 (N_3839,In_1746,In_241);
nand U3840 (N_3840,In_2393,In_1840);
nor U3841 (N_3841,In_2428,In_2248);
xnor U3842 (N_3842,In_1391,In_1973);
nor U3843 (N_3843,In_611,In_2004);
xnor U3844 (N_3844,In_445,In_2468);
nand U3845 (N_3845,In_15,In_1271);
nand U3846 (N_3846,In_55,In_1601);
xor U3847 (N_3847,In_1625,In_1924);
nor U3848 (N_3848,In_889,In_2027);
or U3849 (N_3849,In_895,In_1977);
and U3850 (N_3850,In_512,In_957);
xor U3851 (N_3851,In_20,In_186);
nor U3852 (N_3852,In_1736,In_1270);
nor U3853 (N_3853,In_553,In_726);
nand U3854 (N_3854,In_2250,In_1030);
and U3855 (N_3855,In_1611,In_313);
and U3856 (N_3856,In_739,In_2419);
nand U3857 (N_3857,In_2231,In_129);
and U3858 (N_3858,In_1072,In_297);
or U3859 (N_3859,In_1217,In_269);
and U3860 (N_3860,In_754,In_1120);
nor U3861 (N_3861,In_491,In_770);
nor U3862 (N_3862,In_1493,In_9);
xor U3863 (N_3863,In_1456,In_1343);
nand U3864 (N_3864,In_89,In_76);
xor U3865 (N_3865,In_462,In_148);
or U3866 (N_3866,In_1277,In_2070);
nor U3867 (N_3867,In_1789,In_2407);
nand U3868 (N_3868,In_1843,In_610);
nor U3869 (N_3869,In_1648,In_1788);
and U3870 (N_3870,In_745,In_1888);
or U3871 (N_3871,In_1101,In_2409);
nor U3872 (N_3872,In_650,In_1488);
nand U3873 (N_3873,In_1204,In_521);
or U3874 (N_3874,In_951,In_1846);
and U3875 (N_3875,In_549,In_2484);
or U3876 (N_3876,In_796,In_1943);
nor U3877 (N_3877,In_280,In_1350);
nand U3878 (N_3878,In_1640,In_1853);
nor U3879 (N_3879,In_1660,In_2106);
nand U3880 (N_3880,In_920,In_1353);
nand U3881 (N_3881,In_579,In_685);
nand U3882 (N_3882,In_2230,In_1815);
and U3883 (N_3883,In_1929,In_2246);
or U3884 (N_3884,In_443,In_2302);
or U3885 (N_3885,In_516,In_637);
xnor U3886 (N_3886,In_451,In_1913);
and U3887 (N_3887,In_2424,In_492);
and U3888 (N_3888,In_810,In_1856);
and U3889 (N_3889,In_198,In_2174);
nand U3890 (N_3890,In_440,In_693);
nor U3891 (N_3891,In_1996,In_1182);
or U3892 (N_3892,In_2361,In_1172);
nor U3893 (N_3893,In_1944,In_2354);
or U3894 (N_3894,In_2167,In_1112);
nor U3895 (N_3895,In_575,In_965);
or U3896 (N_3896,In_223,In_606);
xor U3897 (N_3897,In_1410,In_906);
and U3898 (N_3898,In_165,In_187);
nor U3899 (N_3899,In_402,In_459);
nor U3900 (N_3900,In_1515,In_1465);
nor U3901 (N_3901,In_1829,In_1538);
nor U3902 (N_3902,In_2250,In_67);
nor U3903 (N_3903,In_56,In_1678);
or U3904 (N_3904,In_1751,In_300);
or U3905 (N_3905,In_195,In_1040);
nor U3906 (N_3906,In_122,In_26);
nor U3907 (N_3907,In_770,In_2069);
and U3908 (N_3908,In_341,In_1246);
nand U3909 (N_3909,In_307,In_1309);
and U3910 (N_3910,In_1274,In_2432);
and U3911 (N_3911,In_1095,In_752);
xor U3912 (N_3912,In_1626,In_2392);
nand U3913 (N_3913,In_2032,In_1249);
nor U3914 (N_3914,In_1002,In_2163);
or U3915 (N_3915,In_16,In_2268);
or U3916 (N_3916,In_1332,In_2230);
nand U3917 (N_3917,In_2253,In_1846);
nand U3918 (N_3918,In_964,In_732);
and U3919 (N_3919,In_1838,In_185);
or U3920 (N_3920,In_425,In_508);
and U3921 (N_3921,In_441,In_360);
nand U3922 (N_3922,In_1635,In_2063);
nand U3923 (N_3923,In_2228,In_2323);
or U3924 (N_3924,In_1481,In_1315);
or U3925 (N_3925,In_1625,In_887);
xnor U3926 (N_3926,In_396,In_436);
or U3927 (N_3927,In_947,In_52);
or U3928 (N_3928,In_947,In_2278);
nor U3929 (N_3929,In_1360,In_1293);
or U3930 (N_3930,In_2266,In_156);
nor U3931 (N_3931,In_1442,In_2164);
nand U3932 (N_3932,In_1205,In_1032);
and U3933 (N_3933,In_1464,In_1608);
or U3934 (N_3934,In_90,In_1120);
and U3935 (N_3935,In_1319,In_2327);
xor U3936 (N_3936,In_1578,In_469);
and U3937 (N_3937,In_1615,In_1228);
and U3938 (N_3938,In_1820,In_2197);
nand U3939 (N_3939,In_893,In_73);
nor U3940 (N_3940,In_268,In_534);
and U3941 (N_3941,In_353,In_1809);
xor U3942 (N_3942,In_314,In_373);
or U3943 (N_3943,In_1079,In_2058);
xor U3944 (N_3944,In_1811,In_1803);
and U3945 (N_3945,In_998,In_1);
or U3946 (N_3946,In_966,In_608);
or U3947 (N_3947,In_977,In_289);
nor U3948 (N_3948,In_1780,In_1630);
nor U3949 (N_3949,In_2374,In_1782);
nor U3950 (N_3950,In_1753,In_942);
nor U3951 (N_3951,In_1307,In_1795);
or U3952 (N_3952,In_2103,In_2135);
and U3953 (N_3953,In_64,In_2215);
nand U3954 (N_3954,In_1611,In_2094);
and U3955 (N_3955,In_2018,In_916);
or U3956 (N_3956,In_1437,In_1382);
nor U3957 (N_3957,In_2227,In_1108);
nand U3958 (N_3958,In_2377,In_940);
xor U3959 (N_3959,In_512,In_1562);
nand U3960 (N_3960,In_1861,In_2365);
or U3961 (N_3961,In_292,In_1626);
nand U3962 (N_3962,In_1751,In_1051);
or U3963 (N_3963,In_2011,In_573);
nor U3964 (N_3964,In_614,In_1245);
and U3965 (N_3965,In_1325,In_689);
and U3966 (N_3966,In_27,In_1958);
nand U3967 (N_3967,In_2208,In_221);
and U3968 (N_3968,In_1793,In_165);
xor U3969 (N_3969,In_1794,In_1088);
nor U3970 (N_3970,In_1153,In_2150);
or U3971 (N_3971,In_1288,In_868);
nor U3972 (N_3972,In_2309,In_2440);
or U3973 (N_3973,In_1358,In_419);
and U3974 (N_3974,In_1450,In_1830);
nand U3975 (N_3975,In_582,In_2353);
or U3976 (N_3976,In_770,In_1683);
nor U3977 (N_3977,In_1942,In_1863);
nand U3978 (N_3978,In_2393,In_1769);
nor U3979 (N_3979,In_831,In_2478);
nor U3980 (N_3980,In_93,In_1063);
nor U3981 (N_3981,In_1097,In_2197);
and U3982 (N_3982,In_374,In_280);
and U3983 (N_3983,In_1178,In_677);
nand U3984 (N_3984,In_1567,In_149);
and U3985 (N_3985,In_2173,In_1591);
xor U3986 (N_3986,In_416,In_1328);
nand U3987 (N_3987,In_937,In_1492);
xnor U3988 (N_3988,In_1197,In_120);
nand U3989 (N_3989,In_2120,In_703);
or U3990 (N_3990,In_496,In_2497);
or U3991 (N_3991,In_391,In_1262);
nor U3992 (N_3992,In_1252,In_2252);
nor U3993 (N_3993,In_1342,In_549);
and U3994 (N_3994,In_1589,In_716);
and U3995 (N_3995,In_1402,In_1883);
nor U3996 (N_3996,In_1300,In_120);
and U3997 (N_3997,In_2022,In_1359);
and U3998 (N_3998,In_1468,In_2397);
nor U3999 (N_3999,In_712,In_2433);
nor U4000 (N_4000,In_1698,In_1185);
nor U4001 (N_4001,In_1500,In_1896);
xnor U4002 (N_4002,In_276,In_92);
or U4003 (N_4003,In_978,In_2449);
nand U4004 (N_4004,In_239,In_1538);
and U4005 (N_4005,In_851,In_87);
and U4006 (N_4006,In_1473,In_339);
and U4007 (N_4007,In_1613,In_2460);
and U4008 (N_4008,In_40,In_591);
nand U4009 (N_4009,In_981,In_298);
or U4010 (N_4010,In_2146,In_2104);
nand U4011 (N_4011,In_642,In_992);
and U4012 (N_4012,In_2477,In_561);
or U4013 (N_4013,In_2248,In_196);
and U4014 (N_4014,In_1603,In_1984);
and U4015 (N_4015,In_1886,In_1001);
or U4016 (N_4016,In_1871,In_240);
and U4017 (N_4017,In_1128,In_1901);
and U4018 (N_4018,In_709,In_100);
and U4019 (N_4019,In_2499,In_1446);
or U4020 (N_4020,In_2317,In_1863);
or U4021 (N_4021,In_2423,In_483);
nand U4022 (N_4022,In_642,In_1511);
and U4023 (N_4023,In_557,In_839);
and U4024 (N_4024,In_2276,In_2152);
or U4025 (N_4025,In_2419,In_137);
or U4026 (N_4026,In_1969,In_845);
nor U4027 (N_4027,In_1724,In_244);
nor U4028 (N_4028,In_1592,In_1859);
nand U4029 (N_4029,In_1391,In_387);
nor U4030 (N_4030,In_582,In_171);
nor U4031 (N_4031,In_852,In_2203);
and U4032 (N_4032,In_186,In_2013);
nor U4033 (N_4033,In_248,In_1316);
nor U4034 (N_4034,In_627,In_2051);
and U4035 (N_4035,In_400,In_2032);
nor U4036 (N_4036,In_526,In_1053);
or U4037 (N_4037,In_541,In_1497);
nand U4038 (N_4038,In_766,In_681);
or U4039 (N_4039,In_1927,In_379);
or U4040 (N_4040,In_1444,In_1788);
nand U4041 (N_4041,In_696,In_884);
nand U4042 (N_4042,In_2376,In_1562);
nand U4043 (N_4043,In_67,In_266);
and U4044 (N_4044,In_2262,In_239);
nor U4045 (N_4045,In_2273,In_1988);
and U4046 (N_4046,In_2389,In_2194);
or U4047 (N_4047,In_2042,In_1670);
and U4048 (N_4048,In_810,In_1714);
nor U4049 (N_4049,In_1527,In_2202);
or U4050 (N_4050,In_596,In_1743);
nand U4051 (N_4051,In_511,In_2010);
xor U4052 (N_4052,In_970,In_2472);
or U4053 (N_4053,In_349,In_1462);
nor U4054 (N_4054,In_1329,In_424);
nor U4055 (N_4055,In_1760,In_701);
and U4056 (N_4056,In_2296,In_2020);
or U4057 (N_4057,In_742,In_1397);
or U4058 (N_4058,In_1990,In_927);
xnor U4059 (N_4059,In_641,In_1204);
or U4060 (N_4060,In_2369,In_19);
and U4061 (N_4061,In_1986,In_1498);
nor U4062 (N_4062,In_1122,In_1772);
or U4063 (N_4063,In_896,In_1832);
nand U4064 (N_4064,In_2158,In_281);
nor U4065 (N_4065,In_2001,In_1610);
and U4066 (N_4066,In_662,In_2412);
or U4067 (N_4067,In_276,In_521);
xor U4068 (N_4068,In_1840,In_1483);
or U4069 (N_4069,In_457,In_2025);
xnor U4070 (N_4070,In_1936,In_524);
nand U4071 (N_4071,In_2101,In_233);
nor U4072 (N_4072,In_2292,In_1402);
xnor U4073 (N_4073,In_1776,In_400);
or U4074 (N_4074,In_2428,In_1454);
nor U4075 (N_4075,In_60,In_523);
or U4076 (N_4076,In_961,In_1678);
nor U4077 (N_4077,In_1258,In_1610);
nand U4078 (N_4078,In_2320,In_922);
nor U4079 (N_4079,In_2453,In_975);
nand U4080 (N_4080,In_938,In_2231);
or U4081 (N_4081,In_321,In_1003);
nand U4082 (N_4082,In_1621,In_1168);
or U4083 (N_4083,In_1641,In_2215);
nor U4084 (N_4084,In_224,In_1261);
or U4085 (N_4085,In_2456,In_988);
xnor U4086 (N_4086,In_2222,In_104);
nand U4087 (N_4087,In_1393,In_1191);
nor U4088 (N_4088,In_201,In_1346);
nand U4089 (N_4089,In_1194,In_766);
nand U4090 (N_4090,In_729,In_2313);
nor U4091 (N_4091,In_1495,In_1832);
or U4092 (N_4092,In_772,In_1740);
nand U4093 (N_4093,In_2124,In_884);
nor U4094 (N_4094,In_1860,In_1559);
nand U4095 (N_4095,In_623,In_722);
nor U4096 (N_4096,In_485,In_2457);
nor U4097 (N_4097,In_1705,In_1958);
and U4098 (N_4098,In_1873,In_1904);
or U4099 (N_4099,In_1660,In_1029);
or U4100 (N_4100,In_1287,In_809);
nor U4101 (N_4101,In_1960,In_2282);
nand U4102 (N_4102,In_1828,In_632);
nor U4103 (N_4103,In_2078,In_425);
nor U4104 (N_4104,In_2356,In_2174);
or U4105 (N_4105,In_377,In_589);
xnor U4106 (N_4106,In_1877,In_226);
or U4107 (N_4107,In_1371,In_1100);
and U4108 (N_4108,In_1352,In_610);
or U4109 (N_4109,In_264,In_180);
and U4110 (N_4110,In_2133,In_2494);
and U4111 (N_4111,In_271,In_968);
nand U4112 (N_4112,In_767,In_1698);
or U4113 (N_4113,In_830,In_1638);
nand U4114 (N_4114,In_430,In_6);
or U4115 (N_4115,In_1701,In_966);
xor U4116 (N_4116,In_553,In_1122);
or U4117 (N_4117,In_864,In_590);
nand U4118 (N_4118,In_749,In_1722);
nand U4119 (N_4119,In_2221,In_2456);
xor U4120 (N_4120,In_985,In_2024);
nand U4121 (N_4121,In_186,In_2454);
nand U4122 (N_4122,In_2079,In_2267);
nand U4123 (N_4123,In_2129,In_2198);
nor U4124 (N_4124,In_466,In_2156);
or U4125 (N_4125,In_1725,In_2267);
and U4126 (N_4126,In_2367,In_1311);
nor U4127 (N_4127,In_2251,In_1688);
nor U4128 (N_4128,In_2079,In_1851);
nor U4129 (N_4129,In_1088,In_552);
nand U4130 (N_4130,In_1212,In_676);
xnor U4131 (N_4131,In_2387,In_1520);
or U4132 (N_4132,In_562,In_1472);
or U4133 (N_4133,In_2321,In_415);
nor U4134 (N_4134,In_2155,In_2266);
or U4135 (N_4135,In_88,In_1454);
nand U4136 (N_4136,In_1258,In_888);
or U4137 (N_4137,In_1541,In_320);
or U4138 (N_4138,In_2435,In_1369);
and U4139 (N_4139,In_1306,In_412);
nand U4140 (N_4140,In_632,In_2484);
and U4141 (N_4141,In_528,In_886);
nand U4142 (N_4142,In_904,In_1126);
or U4143 (N_4143,In_5,In_2130);
nor U4144 (N_4144,In_1060,In_853);
nor U4145 (N_4145,In_388,In_1750);
nor U4146 (N_4146,In_1216,In_528);
or U4147 (N_4147,In_290,In_1248);
nor U4148 (N_4148,In_704,In_1503);
or U4149 (N_4149,In_2376,In_1757);
and U4150 (N_4150,In_319,In_291);
nand U4151 (N_4151,In_2452,In_2257);
nand U4152 (N_4152,In_2135,In_1345);
nor U4153 (N_4153,In_992,In_160);
or U4154 (N_4154,In_1871,In_2217);
or U4155 (N_4155,In_1378,In_1197);
nand U4156 (N_4156,In_443,In_585);
and U4157 (N_4157,In_672,In_585);
and U4158 (N_4158,In_275,In_888);
and U4159 (N_4159,In_1910,In_933);
or U4160 (N_4160,In_187,In_251);
nor U4161 (N_4161,In_1028,In_1854);
xnor U4162 (N_4162,In_1304,In_226);
or U4163 (N_4163,In_578,In_63);
or U4164 (N_4164,In_1285,In_472);
xor U4165 (N_4165,In_2325,In_1831);
nor U4166 (N_4166,In_710,In_112);
nand U4167 (N_4167,In_697,In_1122);
nand U4168 (N_4168,In_1436,In_1647);
or U4169 (N_4169,In_1365,In_1928);
nor U4170 (N_4170,In_87,In_931);
and U4171 (N_4171,In_2192,In_2288);
and U4172 (N_4172,In_1019,In_60);
nand U4173 (N_4173,In_837,In_361);
and U4174 (N_4174,In_1603,In_160);
nor U4175 (N_4175,In_207,In_1545);
xnor U4176 (N_4176,In_1377,In_426);
nand U4177 (N_4177,In_533,In_534);
or U4178 (N_4178,In_1426,In_2135);
and U4179 (N_4179,In_706,In_156);
nand U4180 (N_4180,In_853,In_1097);
or U4181 (N_4181,In_1320,In_1911);
or U4182 (N_4182,In_1556,In_2190);
nor U4183 (N_4183,In_261,In_878);
nor U4184 (N_4184,In_12,In_2204);
xor U4185 (N_4185,In_781,In_1182);
or U4186 (N_4186,In_720,In_1375);
and U4187 (N_4187,In_365,In_1089);
xor U4188 (N_4188,In_1002,In_335);
nand U4189 (N_4189,In_1998,In_1361);
nand U4190 (N_4190,In_52,In_202);
nor U4191 (N_4191,In_2146,In_2400);
and U4192 (N_4192,In_1223,In_718);
xor U4193 (N_4193,In_619,In_2134);
or U4194 (N_4194,In_1583,In_115);
nor U4195 (N_4195,In_37,In_393);
or U4196 (N_4196,In_2164,In_320);
nand U4197 (N_4197,In_2338,In_1373);
nand U4198 (N_4198,In_1513,In_1547);
nor U4199 (N_4199,In_273,In_1721);
nor U4200 (N_4200,In_1467,In_1807);
or U4201 (N_4201,In_1630,In_1741);
nor U4202 (N_4202,In_1890,In_824);
and U4203 (N_4203,In_2277,In_1315);
or U4204 (N_4204,In_846,In_382);
nor U4205 (N_4205,In_2036,In_328);
and U4206 (N_4206,In_861,In_2202);
and U4207 (N_4207,In_904,In_598);
nand U4208 (N_4208,In_967,In_1570);
nand U4209 (N_4209,In_299,In_1495);
nor U4210 (N_4210,In_279,In_462);
or U4211 (N_4211,In_1728,In_918);
nor U4212 (N_4212,In_2403,In_859);
nand U4213 (N_4213,In_1446,In_265);
and U4214 (N_4214,In_1023,In_1195);
xor U4215 (N_4215,In_1417,In_1151);
nor U4216 (N_4216,In_2055,In_1202);
and U4217 (N_4217,In_1581,In_1835);
and U4218 (N_4218,In_1826,In_457);
and U4219 (N_4219,In_1142,In_1425);
or U4220 (N_4220,In_782,In_755);
nand U4221 (N_4221,In_1304,In_830);
and U4222 (N_4222,In_2088,In_463);
and U4223 (N_4223,In_1156,In_1889);
nand U4224 (N_4224,In_1398,In_1732);
nor U4225 (N_4225,In_1936,In_2049);
xnor U4226 (N_4226,In_1920,In_1131);
nor U4227 (N_4227,In_1632,In_2251);
nor U4228 (N_4228,In_1784,In_1603);
nor U4229 (N_4229,In_1566,In_1255);
nor U4230 (N_4230,In_524,In_1009);
xnor U4231 (N_4231,In_1931,In_1830);
xor U4232 (N_4232,In_1367,In_1470);
or U4233 (N_4233,In_365,In_2068);
and U4234 (N_4234,In_2419,In_1051);
nand U4235 (N_4235,In_1170,In_2055);
nand U4236 (N_4236,In_1000,In_1559);
nor U4237 (N_4237,In_1936,In_2237);
nand U4238 (N_4238,In_634,In_1706);
nand U4239 (N_4239,In_1794,In_741);
nand U4240 (N_4240,In_439,In_591);
nand U4241 (N_4241,In_57,In_1410);
or U4242 (N_4242,In_545,In_1774);
nor U4243 (N_4243,In_477,In_2120);
or U4244 (N_4244,In_403,In_1696);
nor U4245 (N_4245,In_1355,In_1691);
nand U4246 (N_4246,In_2148,In_2249);
nor U4247 (N_4247,In_1217,In_2361);
nand U4248 (N_4248,In_807,In_1509);
nand U4249 (N_4249,In_1490,In_1130);
or U4250 (N_4250,In_151,In_1989);
or U4251 (N_4251,In_1214,In_1139);
or U4252 (N_4252,In_1242,In_657);
or U4253 (N_4253,In_1965,In_1154);
nor U4254 (N_4254,In_1110,In_816);
or U4255 (N_4255,In_1440,In_643);
and U4256 (N_4256,In_1012,In_999);
or U4257 (N_4257,In_876,In_40);
and U4258 (N_4258,In_1734,In_1539);
and U4259 (N_4259,In_824,In_2493);
and U4260 (N_4260,In_2092,In_227);
and U4261 (N_4261,In_750,In_1255);
and U4262 (N_4262,In_359,In_155);
nand U4263 (N_4263,In_2149,In_1415);
nand U4264 (N_4264,In_1752,In_2001);
and U4265 (N_4265,In_869,In_264);
or U4266 (N_4266,In_1838,In_1784);
and U4267 (N_4267,In_1248,In_89);
or U4268 (N_4268,In_1147,In_832);
nand U4269 (N_4269,In_149,In_1071);
or U4270 (N_4270,In_369,In_2370);
nand U4271 (N_4271,In_184,In_1796);
and U4272 (N_4272,In_915,In_692);
xor U4273 (N_4273,In_413,In_1757);
or U4274 (N_4274,In_2381,In_43);
or U4275 (N_4275,In_2267,In_1635);
and U4276 (N_4276,In_2224,In_364);
nor U4277 (N_4277,In_1454,In_2404);
nor U4278 (N_4278,In_2064,In_76);
nor U4279 (N_4279,In_1636,In_2398);
xor U4280 (N_4280,In_1698,In_1925);
or U4281 (N_4281,In_428,In_1427);
xor U4282 (N_4282,In_2185,In_45);
nand U4283 (N_4283,In_1588,In_1561);
nor U4284 (N_4284,In_469,In_1750);
nand U4285 (N_4285,In_2048,In_1527);
or U4286 (N_4286,In_56,In_64);
or U4287 (N_4287,In_1596,In_77);
nor U4288 (N_4288,In_1574,In_1968);
nor U4289 (N_4289,In_1152,In_407);
xor U4290 (N_4290,In_2499,In_853);
and U4291 (N_4291,In_1856,In_378);
or U4292 (N_4292,In_86,In_352);
xor U4293 (N_4293,In_2444,In_676);
nor U4294 (N_4294,In_2494,In_259);
nor U4295 (N_4295,In_2083,In_1373);
nor U4296 (N_4296,In_564,In_143);
nor U4297 (N_4297,In_2164,In_374);
and U4298 (N_4298,In_1750,In_695);
nor U4299 (N_4299,In_246,In_1377);
and U4300 (N_4300,In_1669,In_2129);
and U4301 (N_4301,In_606,In_2353);
nand U4302 (N_4302,In_1932,In_1500);
nor U4303 (N_4303,In_1001,In_84);
nand U4304 (N_4304,In_1384,In_827);
xnor U4305 (N_4305,In_1356,In_2288);
nand U4306 (N_4306,In_1054,In_1768);
and U4307 (N_4307,In_2066,In_13);
nor U4308 (N_4308,In_589,In_1258);
nor U4309 (N_4309,In_150,In_1537);
and U4310 (N_4310,In_1633,In_568);
xnor U4311 (N_4311,In_574,In_897);
nor U4312 (N_4312,In_1875,In_934);
xnor U4313 (N_4313,In_2322,In_31);
nor U4314 (N_4314,In_1312,In_2324);
nand U4315 (N_4315,In_1450,In_884);
nand U4316 (N_4316,In_1715,In_1309);
nor U4317 (N_4317,In_1174,In_2079);
and U4318 (N_4318,In_111,In_586);
or U4319 (N_4319,In_485,In_131);
nand U4320 (N_4320,In_708,In_2078);
and U4321 (N_4321,In_1300,In_1969);
xor U4322 (N_4322,In_950,In_957);
nor U4323 (N_4323,In_1577,In_1398);
or U4324 (N_4324,In_813,In_763);
nand U4325 (N_4325,In_1926,In_904);
or U4326 (N_4326,In_1704,In_1610);
nor U4327 (N_4327,In_2214,In_1158);
or U4328 (N_4328,In_71,In_531);
or U4329 (N_4329,In_733,In_1673);
and U4330 (N_4330,In_262,In_1288);
and U4331 (N_4331,In_1789,In_791);
and U4332 (N_4332,In_1297,In_1008);
and U4333 (N_4333,In_1097,In_2415);
and U4334 (N_4334,In_292,In_1915);
or U4335 (N_4335,In_1761,In_402);
or U4336 (N_4336,In_2110,In_1948);
and U4337 (N_4337,In_852,In_1914);
xor U4338 (N_4338,In_525,In_163);
xnor U4339 (N_4339,In_93,In_1141);
xnor U4340 (N_4340,In_1228,In_1859);
xnor U4341 (N_4341,In_949,In_5);
or U4342 (N_4342,In_1118,In_1121);
and U4343 (N_4343,In_1005,In_2370);
or U4344 (N_4344,In_677,In_1922);
nand U4345 (N_4345,In_932,In_846);
or U4346 (N_4346,In_2189,In_997);
nor U4347 (N_4347,In_2134,In_925);
nor U4348 (N_4348,In_1695,In_1378);
nor U4349 (N_4349,In_1968,In_425);
or U4350 (N_4350,In_1357,In_1843);
or U4351 (N_4351,In_2181,In_645);
or U4352 (N_4352,In_657,In_264);
nand U4353 (N_4353,In_1943,In_925);
or U4354 (N_4354,In_549,In_1912);
xnor U4355 (N_4355,In_902,In_1169);
and U4356 (N_4356,In_970,In_1882);
xnor U4357 (N_4357,In_1760,In_2298);
and U4358 (N_4358,In_1123,In_2472);
nand U4359 (N_4359,In_240,In_799);
xnor U4360 (N_4360,In_1775,In_1875);
or U4361 (N_4361,In_303,In_1389);
and U4362 (N_4362,In_1870,In_1397);
nand U4363 (N_4363,In_193,In_326);
nor U4364 (N_4364,In_1582,In_716);
or U4365 (N_4365,In_2042,In_2177);
nand U4366 (N_4366,In_2345,In_556);
or U4367 (N_4367,In_1435,In_1815);
or U4368 (N_4368,In_1151,In_1949);
or U4369 (N_4369,In_809,In_103);
xnor U4370 (N_4370,In_2314,In_442);
xnor U4371 (N_4371,In_2064,In_936);
xnor U4372 (N_4372,In_606,In_1938);
nor U4373 (N_4373,In_1313,In_755);
nand U4374 (N_4374,In_1580,In_1323);
or U4375 (N_4375,In_724,In_1618);
nor U4376 (N_4376,In_648,In_1933);
nor U4377 (N_4377,In_1727,In_676);
or U4378 (N_4378,In_2092,In_740);
and U4379 (N_4379,In_2202,In_1973);
nand U4380 (N_4380,In_1312,In_1680);
nor U4381 (N_4381,In_700,In_334);
or U4382 (N_4382,In_266,In_933);
or U4383 (N_4383,In_773,In_419);
or U4384 (N_4384,In_2372,In_582);
nand U4385 (N_4385,In_431,In_645);
and U4386 (N_4386,In_1379,In_1995);
and U4387 (N_4387,In_2076,In_986);
nand U4388 (N_4388,In_1986,In_843);
or U4389 (N_4389,In_784,In_727);
or U4390 (N_4390,In_2071,In_414);
nor U4391 (N_4391,In_675,In_1349);
nor U4392 (N_4392,In_2420,In_1365);
xnor U4393 (N_4393,In_1474,In_1778);
nor U4394 (N_4394,In_1184,In_2336);
nand U4395 (N_4395,In_701,In_42);
or U4396 (N_4396,In_2123,In_2420);
xnor U4397 (N_4397,In_550,In_1362);
nand U4398 (N_4398,In_468,In_1904);
nor U4399 (N_4399,In_1534,In_11);
nor U4400 (N_4400,In_2024,In_856);
nand U4401 (N_4401,In_1761,In_261);
nand U4402 (N_4402,In_1510,In_907);
or U4403 (N_4403,In_2397,In_1669);
nor U4404 (N_4404,In_1815,In_1939);
nand U4405 (N_4405,In_2460,In_662);
nand U4406 (N_4406,In_2114,In_1349);
and U4407 (N_4407,In_1105,In_699);
or U4408 (N_4408,In_1344,In_453);
nand U4409 (N_4409,In_2241,In_756);
xor U4410 (N_4410,In_2366,In_1146);
or U4411 (N_4411,In_234,In_1512);
or U4412 (N_4412,In_1740,In_583);
nand U4413 (N_4413,In_1586,In_37);
xor U4414 (N_4414,In_1597,In_1136);
xor U4415 (N_4415,In_794,In_977);
nand U4416 (N_4416,In_2075,In_969);
nor U4417 (N_4417,In_1698,In_1502);
and U4418 (N_4418,In_312,In_2237);
nand U4419 (N_4419,In_646,In_456);
and U4420 (N_4420,In_1329,In_1497);
nand U4421 (N_4421,In_1426,In_1384);
or U4422 (N_4422,In_132,In_2306);
nor U4423 (N_4423,In_1919,In_40);
and U4424 (N_4424,In_2030,In_1582);
nand U4425 (N_4425,In_617,In_563);
nand U4426 (N_4426,In_741,In_1854);
and U4427 (N_4427,In_86,In_211);
or U4428 (N_4428,In_192,In_1285);
or U4429 (N_4429,In_2230,In_703);
xnor U4430 (N_4430,In_542,In_1624);
nand U4431 (N_4431,In_48,In_2417);
or U4432 (N_4432,In_1571,In_211);
or U4433 (N_4433,In_549,In_2137);
nand U4434 (N_4434,In_860,In_211);
or U4435 (N_4435,In_1565,In_1786);
and U4436 (N_4436,In_353,In_2343);
and U4437 (N_4437,In_2274,In_1081);
or U4438 (N_4438,In_264,In_215);
or U4439 (N_4439,In_2375,In_397);
xor U4440 (N_4440,In_868,In_1954);
and U4441 (N_4441,In_1639,In_2092);
and U4442 (N_4442,In_1499,In_1651);
nand U4443 (N_4443,In_2019,In_1495);
and U4444 (N_4444,In_671,In_2337);
nor U4445 (N_4445,In_2403,In_1785);
xor U4446 (N_4446,In_1241,In_96);
nand U4447 (N_4447,In_185,In_537);
nor U4448 (N_4448,In_1841,In_341);
nor U4449 (N_4449,In_207,In_416);
and U4450 (N_4450,In_1405,In_1799);
nor U4451 (N_4451,In_651,In_993);
and U4452 (N_4452,In_583,In_1027);
or U4453 (N_4453,In_905,In_1041);
xor U4454 (N_4454,In_1360,In_271);
xnor U4455 (N_4455,In_271,In_880);
or U4456 (N_4456,In_1324,In_1812);
xor U4457 (N_4457,In_32,In_2132);
nor U4458 (N_4458,In_1898,In_1370);
and U4459 (N_4459,In_921,In_1308);
or U4460 (N_4460,In_2277,In_509);
and U4461 (N_4461,In_1620,In_692);
nor U4462 (N_4462,In_2279,In_1492);
and U4463 (N_4463,In_1953,In_2131);
or U4464 (N_4464,In_530,In_2132);
or U4465 (N_4465,In_2443,In_262);
nand U4466 (N_4466,In_1184,In_1636);
nor U4467 (N_4467,In_471,In_638);
nor U4468 (N_4468,In_2108,In_854);
and U4469 (N_4469,In_2456,In_1475);
nand U4470 (N_4470,In_1916,In_1329);
nand U4471 (N_4471,In_1494,In_1341);
or U4472 (N_4472,In_943,In_1252);
nor U4473 (N_4473,In_2008,In_1086);
and U4474 (N_4474,In_858,In_234);
and U4475 (N_4475,In_578,In_840);
nand U4476 (N_4476,In_344,In_522);
xor U4477 (N_4477,In_1218,In_2183);
nand U4478 (N_4478,In_51,In_2087);
xor U4479 (N_4479,In_2295,In_1018);
nand U4480 (N_4480,In_341,In_2271);
nor U4481 (N_4481,In_1778,In_545);
nor U4482 (N_4482,In_1364,In_318);
nor U4483 (N_4483,In_2032,In_264);
and U4484 (N_4484,In_1705,In_1359);
and U4485 (N_4485,In_1829,In_61);
xnor U4486 (N_4486,In_360,In_404);
and U4487 (N_4487,In_1254,In_202);
and U4488 (N_4488,In_766,In_1244);
or U4489 (N_4489,In_1381,In_1139);
nor U4490 (N_4490,In_1178,In_1360);
nand U4491 (N_4491,In_603,In_1950);
or U4492 (N_4492,In_776,In_1591);
nor U4493 (N_4493,In_2187,In_1410);
nor U4494 (N_4494,In_2193,In_1611);
nor U4495 (N_4495,In_1539,In_1242);
nand U4496 (N_4496,In_1450,In_1812);
nand U4497 (N_4497,In_932,In_2491);
nor U4498 (N_4498,In_61,In_1222);
or U4499 (N_4499,In_1389,In_421);
nor U4500 (N_4500,In_1931,In_809);
nor U4501 (N_4501,In_2097,In_1278);
nor U4502 (N_4502,In_228,In_2423);
or U4503 (N_4503,In_1235,In_1660);
xor U4504 (N_4504,In_2269,In_1812);
or U4505 (N_4505,In_2123,In_1387);
and U4506 (N_4506,In_95,In_369);
nor U4507 (N_4507,In_1629,In_563);
and U4508 (N_4508,In_963,In_2351);
xor U4509 (N_4509,In_2351,In_1891);
or U4510 (N_4510,In_48,In_755);
nor U4511 (N_4511,In_881,In_1419);
nand U4512 (N_4512,In_94,In_1557);
nor U4513 (N_4513,In_1078,In_2135);
and U4514 (N_4514,In_137,In_1526);
and U4515 (N_4515,In_2456,In_2140);
and U4516 (N_4516,In_79,In_1913);
and U4517 (N_4517,In_260,In_2282);
and U4518 (N_4518,In_2429,In_46);
and U4519 (N_4519,In_1130,In_752);
and U4520 (N_4520,In_536,In_1669);
and U4521 (N_4521,In_707,In_71);
nand U4522 (N_4522,In_1728,In_2034);
nor U4523 (N_4523,In_2341,In_9);
nand U4524 (N_4524,In_649,In_336);
xnor U4525 (N_4525,In_1590,In_511);
and U4526 (N_4526,In_176,In_1838);
nand U4527 (N_4527,In_1480,In_602);
and U4528 (N_4528,In_1168,In_1237);
nand U4529 (N_4529,In_1506,In_1617);
or U4530 (N_4530,In_401,In_1455);
or U4531 (N_4531,In_702,In_2200);
and U4532 (N_4532,In_606,In_1166);
nor U4533 (N_4533,In_1709,In_834);
nand U4534 (N_4534,In_875,In_1346);
nand U4535 (N_4535,In_25,In_562);
nor U4536 (N_4536,In_356,In_1140);
nor U4537 (N_4537,In_1523,In_1776);
xor U4538 (N_4538,In_435,In_1066);
nor U4539 (N_4539,In_2183,In_498);
or U4540 (N_4540,In_305,In_1191);
nand U4541 (N_4541,In_1093,In_175);
or U4542 (N_4542,In_1169,In_1449);
or U4543 (N_4543,In_195,In_1661);
or U4544 (N_4544,In_991,In_1598);
xnor U4545 (N_4545,In_323,In_1639);
or U4546 (N_4546,In_222,In_2347);
xor U4547 (N_4547,In_1292,In_1129);
or U4548 (N_4548,In_118,In_804);
or U4549 (N_4549,In_1386,In_2182);
nand U4550 (N_4550,In_587,In_2435);
or U4551 (N_4551,In_2018,In_1457);
or U4552 (N_4552,In_2246,In_1566);
and U4553 (N_4553,In_1711,In_1071);
nand U4554 (N_4554,In_2427,In_453);
or U4555 (N_4555,In_39,In_1337);
nand U4556 (N_4556,In_712,In_463);
or U4557 (N_4557,In_982,In_704);
and U4558 (N_4558,In_2348,In_1549);
and U4559 (N_4559,In_7,In_118);
nand U4560 (N_4560,In_297,In_1214);
and U4561 (N_4561,In_995,In_1210);
nand U4562 (N_4562,In_281,In_2434);
and U4563 (N_4563,In_2048,In_1447);
nand U4564 (N_4564,In_2457,In_2124);
and U4565 (N_4565,In_698,In_2050);
xnor U4566 (N_4566,In_2262,In_1142);
xnor U4567 (N_4567,In_538,In_2305);
nor U4568 (N_4568,In_104,In_1779);
nand U4569 (N_4569,In_846,In_1975);
and U4570 (N_4570,In_2264,In_1492);
nand U4571 (N_4571,In_100,In_1051);
nand U4572 (N_4572,In_386,In_1090);
nand U4573 (N_4573,In_1075,In_1752);
or U4574 (N_4574,In_1674,In_2045);
nor U4575 (N_4575,In_1969,In_2309);
xor U4576 (N_4576,In_860,In_1023);
xor U4577 (N_4577,In_1397,In_1319);
or U4578 (N_4578,In_711,In_1686);
nor U4579 (N_4579,In_797,In_1709);
or U4580 (N_4580,In_2274,In_1334);
or U4581 (N_4581,In_2005,In_1749);
and U4582 (N_4582,In_976,In_1553);
nand U4583 (N_4583,In_1231,In_38);
nor U4584 (N_4584,In_688,In_185);
and U4585 (N_4585,In_1317,In_1485);
or U4586 (N_4586,In_669,In_390);
nand U4587 (N_4587,In_1876,In_829);
or U4588 (N_4588,In_1341,In_64);
nand U4589 (N_4589,In_297,In_932);
nand U4590 (N_4590,In_1052,In_1609);
nand U4591 (N_4591,In_581,In_2207);
or U4592 (N_4592,In_2036,In_727);
nand U4593 (N_4593,In_807,In_44);
or U4594 (N_4594,In_1450,In_1213);
and U4595 (N_4595,In_1598,In_1623);
and U4596 (N_4596,In_694,In_2411);
and U4597 (N_4597,In_829,In_1540);
nand U4598 (N_4598,In_228,In_2277);
nand U4599 (N_4599,In_1960,In_173);
and U4600 (N_4600,In_1792,In_1658);
nor U4601 (N_4601,In_1204,In_1714);
nor U4602 (N_4602,In_2164,In_2198);
and U4603 (N_4603,In_375,In_91);
nor U4604 (N_4604,In_1031,In_819);
xor U4605 (N_4605,In_161,In_755);
and U4606 (N_4606,In_1107,In_612);
or U4607 (N_4607,In_1498,In_1435);
or U4608 (N_4608,In_2108,In_414);
or U4609 (N_4609,In_1357,In_2186);
nor U4610 (N_4610,In_1745,In_535);
nor U4611 (N_4611,In_856,In_226);
nor U4612 (N_4612,In_1405,In_1472);
or U4613 (N_4613,In_5,In_1287);
and U4614 (N_4614,In_2016,In_1490);
nand U4615 (N_4615,In_902,In_492);
nand U4616 (N_4616,In_1744,In_2326);
and U4617 (N_4617,In_2399,In_1621);
nor U4618 (N_4618,In_1045,In_776);
nor U4619 (N_4619,In_2184,In_588);
xor U4620 (N_4620,In_2099,In_2279);
nor U4621 (N_4621,In_2244,In_2064);
xnor U4622 (N_4622,In_1184,In_1178);
or U4623 (N_4623,In_93,In_136);
nand U4624 (N_4624,In_1973,In_1087);
nand U4625 (N_4625,In_825,In_235);
nor U4626 (N_4626,In_1331,In_705);
nand U4627 (N_4627,In_2350,In_183);
and U4628 (N_4628,In_543,In_1089);
and U4629 (N_4629,In_1756,In_2009);
or U4630 (N_4630,In_2484,In_2228);
or U4631 (N_4631,In_1806,In_2409);
or U4632 (N_4632,In_2194,In_2045);
and U4633 (N_4633,In_1532,In_987);
xor U4634 (N_4634,In_226,In_2187);
or U4635 (N_4635,In_444,In_1252);
and U4636 (N_4636,In_1031,In_2106);
and U4637 (N_4637,In_1150,In_1773);
nand U4638 (N_4638,In_989,In_1137);
nand U4639 (N_4639,In_2080,In_1373);
nor U4640 (N_4640,In_1846,In_2036);
or U4641 (N_4641,In_269,In_514);
and U4642 (N_4642,In_698,In_2478);
and U4643 (N_4643,In_2211,In_1303);
and U4644 (N_4644,In_2120,In_1177);
and U4645 (N_4645,In_2163,In_191);
nand U4646 (N_4646,In_1713,In_1128);
xor U4647 (N_4647,In_1874,In_1518);
and U4648 (N_4648,In_549,In_541);
nand U4649 (N_4649,In_103,In_946);
nor U4650 (N_4650,In_1355,In_1003);
nand U4651 (N_4651,In_1931,In_2104);
nor U4652 (N_4652,In_123,In_694);
nand U4653 (N_4653,In_665,In_1380);
nor U4654 (N_4654,In_1048,In_2425);
nor U4655 (N_4655,In_1970,In_489);
nor U4656 (N_4656,In_1231,In_448);
nand U4657 (N_4657,In_2373,In_1768);
and U4658 (N_4658,In_358,In_2381);
nand U4659 (N_4659,In_1949,In_1538);
nor U4660 (N_4660,In_2028,In_1395);
and U4661 (N_4661,In_2158,In_600);
nor U4662 (N_4662,In_1228,In_847);
or U4663 (N_4663,In_1460,In_1639);
and U4664 (N_4664,In_2487,In_1354);
or U4665 (N_4665,In_776,In_2284);
nand U4666 (N_4666,In_1005,In_2441);
xor U4667 (N_4667,In_1150,In_742);
or U4668 (N_4668,In_2078,In_336);
nor U4669 (N_4669,In_471,In_282);
nor U4670 (N_4670,In_580,In_1025);
nand U4671 (N_4671,In_936,In_925);
nor U4672 (N_4672,In_850,In_2077);
and U4673 (N_4673,In_610,In_2390);
xor U4674 (N_4674,In_128,In_1040);
nor U4675 (N_4675,In_1857,In_1530);
nand U4676 (N_4676,In_2367,In_749);
nand U4677 (N_4677,In_940,In_1060);
xnor U4678 (N_4678,In_156,In_1618);
or U4679 (N_4679,In_497,In_1068);
nand U4680 (N_4680,In_194,In_709);
or U4681 (N_4681,In_1771,In_953);
nand U4682 (N_4682,In_2343,In_531);
and U4683 (N_4683,In_202,In_1397);
nor U4684 (N_4684,In_666,In_117);
nand U4685 (N_4685,In_2177,In_587);
nor U4686 (N_4686,In_2320,In_652);
or U4687 (N_4687,In_2229,In_1512);
or U4688 (N_4688,In_310,In_12);
nor U4689 (N_4689,In_2332,In_891);
xor U4690 (N_4690,In_699,In_230);
xnor U4691 (N_4691,In_323,In_1290);
or U4692 (N_4692,In_581,In_2373);
nand U4693 (N_4693,In_1776,In_707);
nand U4694 (N_4694,In_816,In_1155);
and U4695 (N_4695,In_691,In_2419);
xor U4696 (N_4696,In_1134,In_235);
nand U4697 (N_4697,In_640,In_116);
or U4698 (N_4698,In_212,In_361);
or U4699 (N_4699,In_1259,In_2060);
nand U4700 (N_4700,In_1981,In_212);
and U4701 (N_4701,In_0,In_456);
and U4702 (N_4702,In_1030,In_1035);
or U4703 (N_4703,In_2109,In_2341);
or U4704 (N_4704,In_718,In_727);
and U4705 (N_4705,In_1762,In_1782);
nand U4706 (N_4706,In_1851,In_1839);
or U4707 (N_4707,In_1776,In_2057);
nor U4708 (N_4708,In_252,In_643);
nor U4709 (N_4709,In_1256,In_1369);
and U4710 (N_4710,In_1517,In_809);
and U4711 (N_4711,In_1981,In_1595);
xor U4712 (N_4712,In_1511,In_919);
xnor U4713 (N_4713,In_2194,In_212);
nor U4714 (N_4714,In_1860,In_2068);
xor U4715 (N_4715,In_1628,In_390);
and U4716 (N_4716,In_1585,In_2412);
nor U4717 (N_4717,In_1476,In_541);
or U4718 (N_4718,In_1032,In_1778);
or U4719 (N_4719,In_1961,In_385);
nor U4720 (N_4720,In_1314,In_1664);
and U4721 (N_4721,In_752,In_233);
nor U4722 (N_4722,In_1818,In_2484);
nor U4723 (N_4723,In_93,In_327);
and U4724 (N_4724,In_2453,In_472);
nand U4725 (N_4725,In_2255,In_1804);
and U4726 (N_4726,In_745,In_2152);
or U4727 (N_4727,In_1730,In_2117);
and U4728 (N_4728,In_2499,In_1830);
and U4729 (N_4729,In_1170,In_2288);
nand U4730 (N_4730,In_2082,In_818);
xor U4731 (N_4731,In_472,In_1856);
or U4732 (N_4732,In_2069,In_897);
nor U4733 (N_4733,In_1567,In_202);
or U4734 (N_4734,In_323,In_967);
and U4735 (N_4735,In_1436,In_1737);
and U4736 (N_4736,In_1657,In_2147);
nor U4737 (N_4737,In_1289,In_2293);
or U4738 (N_4738,In_827,In_1241);
or U4739 (N_4739,In_1629,In_1319);
and U4740 (N_4740,In_2256,In_552);
nand U4741 (N_4741,In_2316,In_1866);
or U4742 (N_4742,In_2179,In_1091);
nor U4743 (N_4743,In_1725,In_883);
or U4744 (N_4744,In_2058,In_254);
nor U4745 (N_4745,In_65,In_2225);
nand U4746 (N_4746,In_2110,In_1476);
xnor U4747 (N_4747,In_2097,In_1147);
nor U4748 (N_4748,In_413,In_2391);
nor U4749 (N_4749,In_1056,In_243);
and U4750 (N_4750,In_505,In_517);
and U4751 (N_4751,In_2494,In_240);
or U4752 (N_4752,In_1461,In_290);
or U4753 (N_4753,In_1519,In_235);
or U4754 (N_4754,In_46,In_1069);
or U4755 (N_4755,In_2189,In_903);
and U4756 (N_4756,In_1273,In_1296);
xor U4757 (N_4757,In_2222,In_1902);
nor U4758 (N_4758,In_2259,In_650);
nor U4759 (N_4759,In_432,In_1118);
nand U4760 (N_4760,In_2033,In_1382);
or U4761 (N_4761,In_982,In_776);
and U4762 (N_4762,In_174,In_1444);
nor U4763 (N_4763,In_1664,In_1366);
nand U4764 (N_4764,In_446,In_916);
nand U4765 (N_4765,In_2052,In_2412);
or U4766 (N_4766,In_189,In_1429);
nand U4767 (N_4767,In_90,In_622);
nand U4768 (N_4768,In_1917,In_1942);
and U4769 (N_4769,In_1754,In_58);
or U4770 (N_4770,In_182,In_1710);
or U4771 (N_4771,In_2235,In_1996);
or U4772 (N_4772,In_61,In_75);
nand U4773 (N_4773,In_1246,In_1409);
or U4774 (N_4774,In_554,In_2257);
nand U4775 (N_4775,In_1451,In_2106);
or U4776 (N_4776,In_126,In_2218);
nor U4777 (N_4777,In_766,In_2284);
nand U4778 (N_4778,In_1918,In_2310);
and U4779 (N_4779,In_49,In_16);
and U4780 (N_4780,In_298,In_1782);
nand U4781 (N_4781,In_2145,In_1055);
nand U4782 (N_4782,In_2109,In_1070);
or U4783 (N_4783,In_1543,In_2204);
nor U4784 (N_4784,In_1243,In_2485);
nand U4785 (N_4785,In_2379,In_2404);
or U4786 (N_4786,In_907,In_2437);
or U4787 (N_4787,In_176,In_991);
nor U4788 (N_4788,In_1741,In_990);
nor U4789 (N_4789,In_60,In_2322);
and U4790 (N_4790,In_863,In_856);
or U4791 (N_4791,In_1836,In_1688);
nand U4792 (N_4792,In_1457,In_951);
xnor U4793 (N_4793,In_901,In_2004);
or U4794 (N_4794,In_1940,In_1038);
xnor U4795 (N_4795,In_1137,In_114);
and U4796 (N_4796,In_1481,In_761);
nand U4797 (N_4797,In_806,In_2317);
nand U4798 (N_4798,In_818,In_1726);
and U4799 (N_4799,In_994,In_1276);
nand U4800 (N_4800,In_900,In_195);
or U4801 (N_4801,In_1763,In_1556);
nor U4802 (N_4802,In_485,In_1419);
or U4803 (N_4803,In_140,In_641);
nor U4804 (N_4804,In_1056,In_1526);
and U4805 (N_4805,In_859,In_325);
nor U4806 (N_4806,In_1746,In_667);
or U4807 (N_4807,In_786,In_2065);
or U4808 (N_4808,In_96,In_1873);
nor U4809 (N_4809,In_1796,In_1281);
and U4810 (N_4810,In_296,In_2018);
nor U4811 (N_4811,In_1533,In_2305);
xor U4812 (N_4812,In_169,In_1023);
nand U4813 (N_4813,In_1475,In_1826);
nand U4814 (N_4814,In_485,In_1565);
nand U4815 (N_4815,In_1839,In_993);
nor U4816 (N_4816,In_267,In_1950);
xor U4817 (N_4817,In_693,In_795);
and U4818 (N_4818,In_2326,In_1031);
or U4819 (N_4819,In_793,In_522);
nor U4820 (N_4820,In_117,In_440);
nor U4821 (N_4821,In_2397,In_460);
nor U4822 (N_4822,In_1946,In_1440);
nor U4823 (N_4823,In_546,In_996);
and U4824 (N_4824,In_934,In_2450);
and U4825 (N_4825,In_1322,In_1153);
nor U4826 (N_4826,In_1588,In_1116);
and U4827 (N_4827,In_1237,In_2305);
or U4828 (N_4828,In_587,In_1379);
and U4829 (N_4829,In_336,In_904);
and U4830 (N_4830,In_1028,In_1568);
and U4831 (N_4831,In_396,In_113);
nor U4832 (N_4832,In_399,In_674);
and U4833 (N_4833,In_204,In_607);
or U4834 (N_4834,In_306,In_782);
or U4835 (N_4835,In_761,In_2338);
and U4836 (N_4836,In_839,In_1991);
nor U4837 (N_4837,In_69,In_1312);
or U4838 (N_4838,In_1912,In_2161);
nor U4839 (N_4839,In_588,In_2120);
or U4840 (N_4840,In_314,In_1475);
nor U4841 (N_4841,In_771,In_202);
nand U4842 (N_4842,In_1404,In_1033);
or U4843 (N_4843,In_673,In_168);
nand U4844 (N_4844,In_1381,In_2471);
and U4845 (N_4845,In_2224,In_1957);
nor U4846 (N_4846,In_466,In_577);
nor U4847 (N_4847,In_1732,In_1185);
or U4848 (N_4848,In_1741,In_1199);
nand U4849 (N_4849,In_2461,In_1429);
or U4850 (N_4850,In_1807,In_324);
or U4851 (N_4851,In_431,In_144);
and U4852 (N_4852,In_1615,In_904);
and U4853 (N_4853,In_950,In_15);
and U4854 (N_4854,In_1571,In_1585);
xnor U4855 (N_4855,In_709,In_713);
and U4856 (N_4856,In_281,In_129);
nand U4857 (N_4857,In_1049,In_1754);
and U4858 (N_4858,In_949,In_1021);
and U4859 (N_4859,In_194,In_1602);
or U4860 (N_4860,In_1617,In_1941);
nor U4861 (N_4861,In_630,In_2316);
nand U4862 (N_4862,In_1198,In_1029);
and U4863 (N_4863,In_706,In_1271);
nand U4864 (N_4864,In_1295,In_2462);
nand U4865 (N_4865,In_1379,In_1916);
nor U4866 (N_4866,In_1005,In_234);
or U4867 (N_4867,In_1458,In_2413);
or U4868 (N_4868,In_517,In_1885);
nand U4869 (N_4869,In_218,In_1609);
nor U4870 (N_4870,In_2248,In_1541);
nand U4871 (N_4871,In_1516,In_156);
nor U4872 (N_4872,In_1827,In_1405);
or U4873 (N_4873,In_2241,In_229);
and U4874 (N_4874,In_692,In_998);
and U4875 (N_4875,In_1865,In_840);
nor U4876 (N_4876,In_1452,In_1389);
or U4877 (N_4877,In_1903,In_2162);
or U4878 (N_4878,In_10,In_235);
xor U4879 (N_4879,In_2266,In_1384);
xnor U4880 (N_4880,In_1815,In_2218);
or U4881 (N_4881,In_2220,In_2189);
nor U4882 (N_4882,In_1154,In_974);
and U4883 (N_4883,In_1064,In_2495);
nand U4884 (N_4884,In_1688,In_1598);
xor U4885 (N_4885,In_2418,In_683);
or U4886 (N_4886,In_593,In_829);
and U4887 (N_4887,In_521,In_1452);
or U4888 (N_4888,In_2312,In_2333);
and U4889 (N_4889,In_1461,In_470);
and U4890 (N_4890,In_2387,In_2127);
and U4891 (N_4891,In_914,In_1009);
or U4892 (N_4892,In_2081,In_648);
and U4893 (N_4893,In_1447,In_857);
nand U4894 (N_4894,In_1258,In_1270);
nand U4895 (N_4895,In_366,In_1282);
or U4896 (N_4896,In_1423,In_1720);
xor U4897 (N_4897,In_2194,In_1274);
or U4898 (N_4898,In_252,In_2240);
and U4899 (N_4899,In_1902,In_1247);
and U4900 (N_4900,In_2231,In_2148);
nor U4901 (N_4901,In_936,In_1952);
or U4902 (N_4902,In_227,In_526);
and U4903 (N_4903,In_1661,In_949);
and U4904 (N_4904,In_1633,In_1411);
nand U4905 (N_4905,In_1446,In_432);
and U4906 (N_4906,In_1505,In_756);
and U4907 (N_4907,In_1828,In_968);
and U4908 (N_4908,In_84,In_1354);
nor U4909 (N_4909,In_908,In_461);
and U4910 (N_4910,In_1595,In_319);
nand U4911 (N_4911,In_12,In_1855);
xor U4912 (N_4912,In_1266,In_1874);
and U4913 (N_4913,In_2161,In_765);
nand U4914 (N_4914,In_94,In_648);
xnor U4915 (N_4915,In_617,In_806);
nor U4916 (N_4916,In_971,In_2171);
nor U4917 (N_4917,In_404,In_892);
nand U4918 (N_4918,In_1299,In_1992);
or U4919 (N_4919,In_1155,In_545);
or U4920 (N_4920,In_1477,In_1453);
or U4921 (N_4921,In_1746,In_1854);
and U4922 (N_4922,In_819,In_1452);
xor U4923 (N_4923,In_16,In_163);
nand U4924 (N_4924,In_1435,In_2004);
or U4925 (N_4925,In_2174,In_1358);
nand U4926 (N_4926,In_2123,In_2179);
nand U4927 (N_4927,In_2030,In_1439);
nand U4928 (N_4928,In_931,In_1791);
nand U4929 (N_4929,In_2025,In_1441);
xnor U4930 (N_4930,In_1643,In_1233);
nor U4931 (N_4931,In_1233,In_1794);
or U4932 (N_4932,In_1715,In_2377);
and U4933 (N_4933,In_519,In_611);
xor U4934 (N_4934,In_157,In_2336);
nand U4935 (N_4935,In_367,In_546);
and U4936 (N_4936,In_1622,In_457);
xnor U4937 (N_4937,In_470,In_422);
and U4938 (N_4938,In_608,In_1959);
and U4939 (N_4939,In_1436,In_466);
or U4940 (N_4940,In_1116,In_2406);
nor U4941 (N_4941,In_1715,In_75);
nand U4942 (N_4942,In_1175,In_138);
or U4943 (N_4943,In_1790,In_982);
and U4944 (N_4944,In_176,In_255);
or U4945 (N_4945,In_976,In_2303);
xnor U4946 (N_4946,In_2136,In_826);
or U4947 (N_4947,In_695,In_1677);
nand U4948 (N_4948,In_77,In_2164);
or U4949 (N_4949,In_607,In_1524);
xnor U4950 (N_4950,In_1093,In_1908);
or U4951 (N_4951,In_1153,In_1253);
nand U4952 (N_4952,In_511,In_1803);
nor U4953 (N_4953,In_2291,In_220);
nor U4954 (N_4954,In_1533,In_269);
nand U4955 (N_4955,In_2314,In_2184);
nor U4956 (N_4956,In_174,In_1097);
nand U4957 (N_4957,In_1704,In_506);
nor U4958 (N_4958,In_159,In_139);
and U4959 (N_4959,In_378,In_1717);
nor U4960 (N_4960,In_257,In_772);
nand U4961 (N_4961,In_2457,In_535);
or U4962 (N_4962,In_1738,In_763);
or U4963 (N_4963,In_2012,In_808);
nand U4964 (N_4964,In_1444,In_746);
or U4965 (N_4965,In_800,In_2095);
and U4966 (N_4966,In_961,In_1731);
or U4967 (N_4967,In_1338,In_1253);
or U4968 (N_4968,In_269,In_808);
and U4969 (N_4969,In_335,In_1688);
nor U4970 (N_4970,In_66,In_219);
nand U4971 (N_4971,In_1039,In_323);
nor U4972 (N_4972,In_1941,In_255);
and U4973 (N_4973,In_295,In_725);
or U4974 (N_4974,In_985,In_863);
and U4975 (N_4975,In_5,In_2497);
or U4976 (N_4976,In_923,In_1027);
xnor U4977 (N_4977,In_1614,In_374);
nand U4978 (N_4978,In_426,In_2055);
nand U4979 (N_4979,In_97,In_945);
and U4980 (N_4980,In_1049,In_331);
or U4981 (N_4981,In_1826,In_1233);
xnor U4982 (N_4982,In_153,In_1716);
xor U4983 (N_4983,In_78,In_1640);
or U4984 (N_4984,In_1292,In_1506);
and U4985 (N_4985,In_1657,In_874);
nand U4986 (N_4986,In_1194,In_2495);
nor U4987 (N_4987,In_1414,In_505);
nand U4988 (N_4988,In_357,In_169);
nand U4989 (N_4989,In_2278,In_1409);
or U4990 (N_4990,In_713,In_1756);
nor U4991 (N_4991,In_885,In_1936);
nor U4992 (N_4992,In_1663,In_1305);
nor U4993 (N_4993,In_2247,In_658);
nand U4994 (N_4994,In_2239,In_2230);
xor U4995 (N_4995,In_656,In_1618);
nand U4996 (N_4996,In_2090,In_1752);
nand U4997 (N_4997,In_122,In_805);
nor U4998 (N_4998,In_1821,In_1740);
or U4999 (N_4999,In_581,In_1872);
or U5000 (N_5000,N_1493,N_3514);
nand U5001 (N_5001,N_2026,N_3013);
and U5002 (N_5002,N_918,N_3958);
or U5003 (N_5003,N_2337,N_4382);
nor U5004 (N_5004,N_2396,N_2761);
or U5005 (N_5005,N_2320,N_526);
nor U5006 (N_5006,N_926,N_1204);
and U5007 (N_5007,N_2294,N_1758);
nor U5008 (N_5008,N_2005,N_2766);
nand U5009 (N_5009,N_3446,N_1475);
nand U5010 (N_5010,N_2328,N_3154);
or U5011 (N_5011,N_2774,N_3584);
nor U5012 (N_5012,N_4394,N_1642);
and U5013 (N_5013,N_4234,N_1282);
nand U5014 (N_5014,N_1084,N_574);
nand U5015 (N_5015,N_555,N_2075);
and U5016 (N_5016,N_1167,N_4468);
and U5017 (N_5017,N_2933,N_4342);
nand U5018 (N_5018,N_1507,N_2148);
or U5019 (N_5019,N_826,N_4918);
nand U5020 (N_5020,N_751,N_3189);
nand U5021 (N_5021,N_54,N_3690);
nor U5022 (N_5022,N_4528,N_4529);
nand U5023 (N_5023,N_4521,N_4741);
nand U5024 (N_5024,N_395,N_4229);
or U5025 (N_5025,N_3065,N_2715);
and U5026 (N_5026,N_1653,N_4497);
xor U5027 (N_5027,N_4130,N_3837);
nand U5028 (N_5028,N_2441,N_4862);
nor U5029 (N_5029,N_2356,N_4732);
nand U5030 (N_5030,N_3671,N_2563);
nand U5031 (N_5031,N_625,N_2288);
xnor U5032 (N_5032,N_2016,N_2713);
and U5033 (N_5033,N_4375,N_286);
or U5034 (N_5034,N_2595,N_2044);
and U5035 (N_5035,N_3447,N_1576);
and U5036 (N_5036,N_424,N_2014);
and U5037 (N_5037,N_717,N_2090);
or U5038 (N_5038,N_4718,N_3249);
nand U5039 (N_5039,N_3565,N_2584);
and U5040 (N_5040,N_4074,N_1625);
nand U5041 (N_5041,N_1601,N_4395);
and U5042 (N_5042,N_403,N_1651);
and U5043 (N_5043,N_1694,N_1911);
nor U5044 (N_5044,N_313,N_3334);
and U5045 (N_5045,N_3324,N_1114);
and U5046 (N_5046,N_2657,N_2366);
or U5047 (N_5047,N_4948,N_1745);
nor U5048 (N_5048,N_3450,N_3346);
xor U5049 (N_5049,N_2027,N_3053);
nor U5050 (N_5050,N_20,N_271);
nor U5051 (N_5051,N_2346,N_1858);
nor U5052 (N_5052,N_2438,N_1034);
and U5053 (N_5053,N_4205,N_4813);
and U5054 (N_5054,N_3380,N_4594);
and U5055 (N_5055,N_3612,N_45);
xnor U5056 (N_5056,N_2447,N_4654);
xnor U5057 (N_5057,N_301,N_2219);
nand U5058 (N_5058,N_1174,N_2154);
nor U5059 (N_5059,N_4501,N_3772);
nand U5060 (N_5060,N_3498,N_1140);
nand U5061 (N_5061,N_617,N_834);
nand U5062 (N_5062,N_4330,N_3451);
nor U5063 (N_5063,N_3820,N_3091);
and U5064 (N_5064,N_3385,N_3859);
xnor U5065 (N_5065,N_3113,N_1272);
and U5066 (N_5066,N_360,N_1192);
nand U5067 (N_5067,N_3864,N_4290);
and U5068 (N_5068,N_3836,N_4142);
nand U5069 (N_5069,N_806,N_3972);
xnor U5070 (N_5070,N_1000,N_199);
nand U5071 (N_5071,N_1336,N_1088);
or U5072 (N_5072,N_2706,N_3829);
or U5073 (N_5073,N_829,N_4751);
nor U5074 (N_5074,N_3771,N_303);
or U5075 (N_5075,N_805,N_2735);
and U5076 (N_5076,N_3683,N_902);
nor U5077 (N_5077,N_4505,N_1721);
nand U5078 (N_5078,N_138,N_3449);
and U5079 (N_5079,N_537,N_1112);
nand U5080 (N_5080,N_595,N_962);
and U5081 (N_5081,N_3174,N_1409);
nor U5082 (N_5082,N_3074,N_2196);
and U5083 (N_5083,N_289,N_2551);
nor U5084 (N_5084,N_487,N_4009);
nand U5085 (N_5085,N_1636,N_2296);
and U5086 (N_5086,N_366,N_3098);
and U5087 (N_5087,N_1367,N_787);
or U5088 (N_5088,N_4867,N_57);
and U5089 (N_5089,N_4160,N_2646);
nor U5090 (N_5090,N_3060,N_1005);
or U5091 (N_5091,N_3581,N_4281);
nand U5092 (N_5092,N_668,N_4301);
nand U5093 (N_5093,N_4136,N_1699);
xor U5094 (N_5094,N_2381,N_3602);
nand U5095 (N_5095,N_3196,N_3577);
and U5096 (N_5096,N_1186,N_4615);
xor U5097 (N_5097,N_3250,N_3102);
xor U5098 (N_5098,N_4806,N_3178);
or U5099 (N_5099,N_4581,N_4688);
nor U5100 (N_5100,N_3945,N_3603);
or U5101 (N_5101,N_3230,N_4117);
and U5102 (N_5102,N_1797,N_295);
nor U5103 (N_5103,N_66,N_3898);
nand U5104 (N_5104,N_2591,N_278);
nor U5105 (N_5105,N_1395,N_1226);
nor U5106 (N_5106,N_139,N_1437);
nand U5107 (N_5107,N_608,N_1345);
nand U5108 (N_5108,N_2237,N_316);
nand U5109 (N_5109,N_4620,N_4910);
nor U5110 (N_5110,N_3630,N_4148);
nor U5111 (N_5111,N_2379,N_2433);
nor U5112 (N_5112,N_2932,N_2564);
and U5113 (N_5113,N_3543,N_2544);
nand U5114 (N_5114,N_3918,N_1203);
nor U5115 (N_5115,N_1033,N_453);
or U5116 (N_5116,N_655,N_4020);
xnor U5117 (N_5117,N_2351,N_937);
nor U5118 (N_5118,N_2202,N_713);
nand U5119 (N_5119,N_120,N_1212);
or U5120 (N_5120,N_1840,N_1945);
nand U5121 (N_5121,N_2530,N_408);
nand U5122 (N_5122,N_4149,N_1944);
nand U5123 (N_5123,N_2034,N_2493);
and U5124 (N_5124,N_3253,N_837);
or U5125 (N_5125,N_3199,N_1236);
or U5126 (N_5126,N_3648,N_1393);
or U5127 (N_5127,N_198,N_1574);
nor U5128 (N_5128,N_1251,N_686);
nor U5129 (N_5129,N_3519,N_2704);
and U5130 (N_5130,N_3860,N_2736);
nand U5131 (N_5131,N_4001,N_1179);
and U5132 (N_5132,N_320,N_2352);
nor U5133 (N_5133,N_34,N_3542);
and U5134 (N_5134,N_4412,N_3057);
nand U5135 (N_5135,N_944,N_2822);
nand U5136 (N_5136,N_447,N_3287);
nand U5137 (N_5137,N_1971,N_2084);
and U5138 (N_5138,N_4269,N_3079);
nor U5139 (N_5139,N_4010,N_4036);
xor U5140 (N_5140,N_4690,N_648);
or U5141 (N_5141,N_3695,N_521);
nand U5142 (N_5142,N_3654,N_637);
and U5143 (N_5143,N_559,N_744);
nor U5144 (N_5144,N_1221,N_756);
nor U5145 (N_5145,N_1963,N_2069);
and U5146 (N_5146,N_1878,N_1731);
or U5147 (N_5147,N_1935,N_4479);
nor U5148 (N_5148,N_3786,N_4173);
nor U5149 (N_5149,N_3442,N_4331);
or U5150 (N_5150,N_211,N_997);
nand U5151 (N_5151,N_461,N_508);
nand U5152 (N_5152,N_179,N_292);
nand U5153 (N_5153,N_4339,N_4220);
nand U5154 (N_5154,N_1967,N_4122);
and U5155 (N_5155,N_1394,N_4843);
nand U5156 (N_5156,N_4379,N_3248);
or U5157 (N_5157,N_641,N_3201);
and U5158 (N_5158,N_2787,N_2889);
nand U5159 (N_5159,N_2740,N_3353);
nand U5160 (N_5160,N_3355,N_3609);
or U5161 (N_5161,N_4304,N_1372);
nor U5162 (N_5162,N_1590,N_4374);
xnor U5163 (N_5163,N_1444,N_2502);
nand U5164 (N_5164,N_3107,N_4707);
nor U5165 (N_5165,N_928,N_892);
or U5166 (N_5166,N_443,N_3061);
nor U5167 (N_5167,N_1629,N_4438);
or U5168 (N_5168,N_536,N_4798);
nand U5169 (N_5169,N_1741,N_3681);
and U5170 (N_5170,N_1952,N_1924);
and U5171 (N_5171,N_2392,N_4228);
nor U5172 (N_5172,N_4733,N_3626);
or U5173 (N_5173,N_1119,N_1687);
nor U5174 (N_5174,N_4264,N_182);
nand U5175 (N_5175,N_1499,N_1368);
nor U5176 (N_5176,N_906,N_1925);
nor U5177 (N_5177,N_2236,N_4039);
and U5178 (N_5178,N_3822,N_4763);
nor U5179 (N_5179,N_724,N_1785);
nand U5180 (N_5180,N_3224,N_2183);
xor U5181 (N_5181,N_2639,N_4437);
or U5182 (N_5182,N_502,N_128);
nand U5183 (N_5183,N_3322,N_1616);
nand U5184 (N_5184,N_1158,N_2605);
nor U5185 (N_5185,N_1920,N_2881);
or U5186 (N_5186,N_478,N_2846);
or U5187 (N_5187,N_1706,N_2238);
nor U5188 (N_5188,N_2962,N_2669);
xnor U5189 (N_5189,N_2828,N_4182);
or U5190 (N_5190,N_977,N_2149);
and U5191 (N_5191,N_904,N_4302);
xnor U5192 (N_5192,N_1051,N_4928);
nor U5193 (N_5193,N_2156,N_4013);
or U5194 (N_5194,N_1001,N_675);
and U5195 (N_5195,N_2764,N_3692);
nor U5196 (N_5196,N_1579,N_1264);
or U5197 (N_5197,N_3598,N_252);
and U5198 (N_5198,N_4087,N_3724);
and U5199 (N_5199,N_3459,N_1916);
nand U5200 (N_5200,N_1985,N_2663);
nand U5201 (N_5201,N_2063,N_1965);
nand U5202 (N_5202,N_3597,N_634);
or U5203 (N_5203,N_2291,N_2282);
xnor U5204 (N_5204,N_302,N_2698);
or U5205 (N_5205,N_4196,N_1894);
nand U5206 (N_5206,N_4223,N_3960);
nand U5207 (N_5207,N_3878,N_2520);
nor U5208 (N_5208,N_373,N_3435);
and U5209 (N_5209,N_3088,N_3509);
or U5210 (N_5210,N_2902,N_4195);
nand U5211 (N_5211,N_178,N_2925);
or U5212 (N_5212,N_650,N_43);
or U5213 (N_5213,N_4586,N_2592);
nor U5214 (N_5214,N_89,N_3875);
nand U5215 (N_5215,N_4666,N_4317);
xnor U5216 (N_5216,N_3448,N_4463);
nand U5217 (N_5217,N_3425,N_784);
nor U5218 (N_5218,N_4099,N_2485);
or U5219 (N_5219,N_3774,N_1974);
nor U5220 (N_5220,N_1,N_3005);
nor U5221 (N_5221,N_4473,N_4729);
nor U5222 (N_5222,N_218,N_3001);
nor U5223 (N_5223,N_4389,N_476);
and U5224 (N_5224,N_579,N_3138);
nand U5225 (N_5225,N_3910,N_3793);
nand U5226 (N_5226,N_3012,N_2786);
nand U5227 (N_5227,N_3210,N_2519);
xor U5228 (N_5228,N_3545,N_851);
and U5229 (N_5229,N_1973,N_1388);
nor U5230 (N_5230,N_3378,N_771);
xor U5231 (N_5231,N_4323,N_881);
nor U5232 (N_5232,N_113,N_1157);
or U5233 (N_5233,N_1181,N_2087);
or U5234 (N_5234,N_3342,N_2949);
nand U5235 (N_5235,N_4315,N_4810);
or U5236 (N_5236,N_2424,N_3920);
nor U5237 (N_5237,N_2675,N_661);
and U5238 (N_5238,N_3949,N_1602);
and U5239 (N_5239,N_2964,N_1242);
or U5240 (N_5240,N_3348,N_3538);
nand U5241 (N_5241,N_1729,N_1068);
or U5242 (N_5242,N_1657,N_2092);
or U5243 (N_5243,N_1627,N_4728);
or U5244 (N_5244,N_4974,N_898);
nor U5245 (N_5245,N_3593,N_4559);
xor U5246 (N_5246,N_4678,N_3198);
nand U5247 (N_5247,N_1232,N_3413);
or U5248 (N_5248,N_4704,N_2710);
nor U5249 (N_5249,N_4980,N_1299);
or U5250 (N_5250,N_3722,N_533);
and U5251 (N_5251,N_3313,N_3532);
nor U5252 (N_5252,N_3047,N_2823);
and U5253 (N_5253,N_3564,N_3606);
and U5254 (N_5254,N_3482,N_1717);
and U5255 (N_5255,N_2406,N_2097);
nand U5256 (N_5256,N_4695,N_4);
and U5257 (N_5257,N_227,N_1392);
nand U5258 (N_5258,N_1734,N_251);
nor U5259 (N_5259,N_2220,N_4185);
and U5260 (N_5260,N_4760,N_3124);
and U5261 (N_5261,N_2340,N_2693);
and U5262 (N_5262,N_3486,N_2842);
nor U5263 (N_5263,N_255,N_3478);
nor U5264 (N_5264,N_4979,N_58);
and U5265 (N_5265,N_4628,N_3437);
nor U5266 (N_5266,N_4932,N_1171);
nand U5267 (N_5267,N_1554,N_1446);
or U5268 (N_5268,N_3309,N_4253);
or U5269 (N_5269,N_1077,N_50);
or U5270 (N_5270,N_1522,N_3844);
nor U5271 (N_5271,N_1802,N_712);
and U5272 (N_5272,N_1360,N_868);
and U5273 (N_5273,N_1006,N_2692);
and U5274 (N_5274,N_4899,N_187);
and U5275 (N_5275,N_4723,N_4855);
nand U5276 (N_5276,N_3158,N_1500);
nor U5277 (N_5277,N_3489,N_953);
and U5278 (N_5278,N_4702,N_1876);
or U5279 (N_5279,N_107,N_155);
nand U5280 (N_5280,N_2900,N_3664);
or U5281 (N_5281,N_274,N_4214);
nand U5282 (N_5282,N_4876,N_4293);
xnor U5283 (N_5283,N_3792,N_3420);
nand U5284 (N_5284,N_4057,N_532);
and U5285 (N_5285,N_1608,N_2694);
and U5286 (N_5286,N_2309,N_44);
or U5287 (N_5287,N_1723,N_4607);
nor U5288 (N_5288,N_963,N_3691);
nor U5289 (N_5289,N_2897,N_1709);
or U5290 (N_5290,N_693,N_378);
nand U5291 (N_5291,N_1194,N_2143);
nand U5292 (N_5292,N_4267,N_4864);
nor U5293 (N_5293,N_4539,N_3140);
and U5294 (N_5294,N_3725,N_2456);
nor U5295 (N_5295,N_828,N_529);
nor U5296 (N_5296,N_2361,N_966);
xnor U5297 (N_5297,N_351,N_3948);
or U5298 (N_5298,N_518,N_3636);
xor U5299 (N_5299,N_2218,N_235);
xnor U5300 (N_5300,N_1777,N_2086);
and U5301 (N_5301,N_3915,N_4530);
and U5302 (N_5302,N_1010,N_716);
nor U5303 (N_5303,N_1124,N_1110);
or U5304 (N_5304,N_26,N_2680);
and U5305 (N_5305,N_2322,N_4610);
nor U5306 (N_5306,N_2719,N_4191);
nor U5307 (N_5307,N_4526,N_4243);
and U5308 (N_5308,N_4168,N_3812);
nor U5309 (N_5309,N_1793,N_2465);
or U5310 (N_5310,N_3137,N_967);
nand U5311 (N_5311,N_3267,N_3983);
nor U5312 (N_5312,N_3651,N_2660);
nand U5313 (N_5313,N_4840,N_1244);
and U5314 (N_5314,N_1754,N_3560);
or U5315 (N_5315,N_612,N_1559);
nor U5316 (N_5316,N_2797,N_832);
or U5317 (N_5317,N_785,N_2391);
and U5318 (N_5318,N_3291,N_798);
xor U5319 (N_5319,N_4477,N_4773);
xnor U5320 (N_5320,N_1126,N_2997);
and U5321 (N_5321,N_2550,N_4764);
nand U5322 (N_5322,N_4047,N_4805);
xor U5323 (N_5323,N_4664,N_3);
and U5324 (N_5324,N_4995,N_3687);
and U5325 (N_5325,N_2998,N_2369);
nand U5326 (N_5326,N_1640,N_2533);
nand U5327 (N_5327,N_2929,N_1866);
nor U5328 (N_5328,N_3000,N_4556);
nand U5329 (N_5329,N_517,N_2999);
nor U5330 (N_5330,N_2690,N_672);
xor U5331 (N_5331,N_124,N_3292);
and U5332 (N_5332,N_2865,N_4675);
nor U5333 (N_5333,N_1565,N_3665);
and U5334 (N_5334,N_878,N_3706);
and U5335 (N_5335,N_889,N_879);
or U5336 (N_5336,N_2877,N_2631);
nand U5337 (N_5337,N_229,N_2370);
nor U5338 (N_5338,N_1122,N_1224);
nand U5339 (N_5339,N_1864,N_148);
nor U5340 (N_5340,N_995,N_3506);
nand U5341 (N_5341,N_2753,N_3685);
or U5342 (N_5342,N_4740,N_4721);
and U5343 (N_5343,N_1266,N_2166);
or U5344 (N_5344,N_221,N_2325);
nor U5345 (N_5345,N_3354,N_1028);
nand U5346 (N_5346,N_2099,N_1402);
and U5347 (N_5347,N_4488,N_669);
nor U5348 (N_5348,N_4513,N_1759);
or U5349 (N_5349,N_1199,N_3089);
xor U5350 (N_5350,N_2944,N_4015);
nor U5351 (N_5351,N_606,N_492);
and U5352 (N_5352,N_3390,N_106);
nor U5353 (N_5353,N_2228,N_2058);
and U5354 (N_5354,N_913,N_1502);
or U5355 (N_5355,N_1940,N_3381);
or U5356 (N_5356,N_3967,N_4857);
xnor U5357 (N_5357,N_2515,N_3017);
and U5358 (N_5358,N_3424,N_4930);
or U5359 (N_5359,N_109,N_690);
nand U5360 (N_5360,N_1190,N_1058);
or U5361 (N_5361,N_210,N_1626);
nand U5362 (N_5362,N_1770,N_547);
nand U5363 (N_5363,N_952,N_4247);
xnor U5364 (N_5364,N_1883,N_4515);
or U5365 (N_5365,N_4249,N_2979);
nor U5366 (N_5366,N_1298,N_3947);
nor U5367 (N_5367,N_3173,N_275);
and U5368 (N_5368,N_4490,N_758);
nor U5369 (N_5369,N_810,N_3139);
nand U5370 (N_5370,N_2714,N_2755);
or U5371 (N_5371,N_464,N_1279);
nand U5372 (N_5372,N_1850,N_3458);
and U5373 (N_5373,N_1738,N_1934);
xor U5374 (N_5374,N_2383,N_1867);
nand U5375 (N_5375,N_4426,N_1968);
nor U5376 (N_5376,N_1847,N_2807);
nor U5377 (N_5377,N_1466,N_1586);
nand U5378 (N_5378,N_2206,N_2686);
nor U5379 (N_5379,N_1455,N_2645);
xor U5380 (N_5380,N_3456,N_2744);
or U5381 (N_5381,N_3930,N_3374);
nor U5382 (N_5382,N_2908,N_3881);
and U5383 (N_5383,N_638,N_1914);
or U5384 (N_5384,N_582,N_1857);
or U5385 (N_5385,N_2231,N_3221);
xor U5386 (N_5386,N_1856,N_4931);
and U5387 (N_5387,N_1461,N_434);
and U5388 (N_5388,N_2720,N_4409);
and U5389 (N_5389,N_4563,N_79);
nor U5390 (N_5390,N_2562,N_1310);
nor U5391 (N_5391,N_2532,N_2338);
nor U5392 (N_5392,N_4255,N_2076);
nand U5393 (N_5393,N_2277,N_611);
xnor U5394 (N_5394,N_4259,N_3738);
nor U5395 (N_5395,N_3366,N_567);
xor U5396 (N_5396,N_2589,N_1156);
nand U5397 (N_5397,N_2610,N_4184);
nor U5398 (N_5398,N_2873,N_335);
or U5399 (N_5399,N_4672,N_3554);
xor U5400 (N_5400,N_264,N_1990);
nor U5401 (N_5401,N_1387,N_41);
or U5402 (N_5402,N_791,N_401);
nor U5403 (N_5403,N_4916,N_2467);
and U5404 (N_5404,N_3950,N_2619);
or U5405 (N_5405,N_2988,N_1730);
and U5406 (N_5406,N_988,N_1252);
nor U5407 (N_5407,N_640,N_4673);
and U5408 (N_5408,N_2286,N_4520);
nor U5409 (N_5409,N_2448,N_4440);
or U5410 (N_5410,N_48,N_3993);
or U5411 (N_5411,N_4052,N_4162);
nor U5412 (N_5412,N_4848,N_2718);
nor U5413 (N_5413,N_55,N_1460);
nor U5414 (N_5414,N_2576,N_4145);
nor U5415 (N_5415,N_4553,N_1659);
and U5416 (N_5416,N_2904,N_3803);
nor U5417 (N_5417,N_4703,N_1655);
nor U5418 (N_5418,N_2200,N_3641);
and U5419 (N_5419,N_1021,N_3419);
xor U5420 (N_5420,N_1353,N_939);
nand U5421 (N_5421,N_4197,N_2269);
nor U5422 (N_5422,N_3283,N_2725);
xor U5423 (N_5423,N_3481,N_1078);
and U5424 (N_5424,N_3764,N_2552);
nor U5425 (N_5425,N_2223,N_2644);
or U5426 (N_5426,N_1685,N_3816);
nor U5427 (N_5427,N_3443,N_1839);
nor U5428 (N_5428,N_4474,N_683);
nand U5429 (N_5429,N_1567,N_2227);
xnor U5430 (N_5430,N_1598,N_2976);
nand U5431 (N_5431,N_697,N_4088);
xnor U5432 (N_5432,N_3022,N_1744);
and U5433 (N_5433,N_2409,N_1188);
or U5434 (N_5434,N_3166,N_2580);
nand U5435 (N_5435,N_1217,N_1082);
or U5436 (N_5436,N_1281,N_733);
nand U5437 (N_5437,N_4606,N_3533);
nand U5438 (N_5438,N_4252,N_80);
or U5439 (N_5439,N_2954,N_3903);
nand U5440 (N_5440,N_4983,N_4970);
xor U5441 (N_5441,N_4770,N_678);
xnor U5442 (N_5442,N_984,N_954);
or U5443 (N_5443,N_4320,N_2358);
or U5444 (N_5444,N_654,N_4063);
or U5445 (N_5445,N_3059,N_1541);
nand U5446 (N_5446,N_3135,N_2763);
and U5447 (N_5447,N_348,N_763);
nor U5448 (N_5448,N_4893,N_332);
nand U5449 (N_5449,N_1441,N_232);
nor U5450 (N_5450,N_1843,N_162);
or U5451 (N_5451,N_4787,N_3999);
xnor U5452 (N_5452,N_2732,N_1781);
or U5453 (N_5453,N_2010,N_1373);
or U5454 (N_5454,N_1686,N_1755);
nand U5455 (N_5455,N_153,N_2127);
nand U5456 (N_5456,N_531,N_2969);
and U5457 (N_5457,N_1237,N_4984);
or U5458 (N_5458,N_2187,N_3904);
and U5459 (N_5459,N_3586,N_1947);
and U5460 (N_5460,N_4943,N_98);
and U5461 (N_5461,N_3808,N_3304);
or U5462 (N_5462,N_3026,N_4710);
xnor U5463 (N_5463,N_396,N_885);
and U5464 (N_5464,N_429,N_1516);
or U5465 (N_5465,N_2491,N_710);
or U5466 (N_5466,N_1648,N_4913);
and U5467 (N_5467,N_1427,N_2091);
nor U5468 (N_5468,N_2538,N_2668);
xor U5469 (N_5469,N_1287,N_268);
nor U5470 (N_5470,N_2751,N_731);
or U5471 (N_5471,N_1481,N_1988);
nand U5472 (N_5472,N_2770,N_2225);
xor U5473 (N_5473,N_4068,N_2845);
nor U5474 (N_5474,N_22,N_297);
nor U5475 (N_5475,N_4854,N_1246);
xor U5476 (N_5476,N_4580,N_3406);
and U5477 (N_5477,N_2537,N_312);
nor U5478 (N_5478,N_4744,N_580);
nor U5479 (N_5479,N_4150,N_4839);
xnor U5480 (N_5480,N_421,N_1415);
nor U5481 (N_5481,N_2184,N_4746);
nand U5482 (N_5482,N_1042,N_2995);
nor U5483 (N_5483,N_353,N_2053);
or U5484 (N_5484,N_3841,N_299);
nor U5485 (N_5485,N_1829,N_3160);
or U5486 (N_5486,N_4126,N_146);
nor U5487 (N_5487,N_4441,N_1634);
and U5488 (N_5488,N_2535,N_4124);
and U5489 (N_5489,N_4841,N_419);
xor U5490 (N_5490,N_942,N_1530);
nor U5491 (N_5491,N_3710,N_1575);
nor U5492 (N_5492,N_370,N_3625);
nand U5493 (N_5493,N_3633,N_564);
nor U5494 (N_5494,N_3117,N_2421);
nor U5495 (N_5495,N_633,N_728);
xnor U5496 (N_5496,N_820,N_1677);
and U5497 (N_5497,N_2212,N_3052);
nor U5498 (N_5498,N_1557,N_194);
nor U5499 (N_5499,N_2574,N_1424);
nor U5500 (N_5500,N_4903,N_4623);
and U5501 (N_5501,N_3400,N_2837);
xor U5502 (N_5502,N_2025,N_698);
nand U5503 (N_5503,N_1011,N_3511);
nor U5504 (N_5504,N_4187,N_2512);
and U5505 (N_5505,N_3835,N_2977);
or U5506 (N_5506,N_854,N_4000);
and U5507 (N_5507,N_919,N_2125);
and U5508 (N_5508,N_3976,N_1258);
nand U5509 (N_5509,N_774,N_1278);
and U5510 (N_5510,N_2510,N_3796);
or U5511 (N_5511,N_4006,N_2966);
nor U5512 (N_5512,N_3824,N_2702);
or U5513 (N_5513,N_623,N_2247);
and U5514 (N_5514,N_4878,N_4922);
or U5515 (N_5515,N_2321,N_2102);
nor U5516 (N_5516,N_2641,N_111);
or U5517 (N_5517,N_1683,N_1145);
or U5518 (N_5518,N_273,N_862);
or U5519 (N_5519,N_420,N_367);
and U5520 (N_5520,N_4527,N_3535);
nand U5521 (N_5521,N_1656,N_3770);
and U5522 (N_5522,N_2859,N_1503);
nor U5523 (N_5523,N_3645,N_976);
or U5524 (N_5524,N_2193,N_1644);
and U5525 (N_5525,N_3684,N_581);
and U5526 (N_5526,N_3848,N_3097);
nor U5527 (N_5527,N_4139,N_115);
nor U5528 (N_5528,N_317,N_3144);
and U5529 (N_5529,N_4357,N_2603);
nand U5530 (N_5530,N_1039,N_1477);
nor U5531 (N_5531,N_4151,N_2869);
and U5532 (N_5532,N_3044,N_1773);
or U5533 (N_5533,N_477,N_3714);
and U5534 (N_5534,N_496,N_3260);
xnor U5535 (N_5535,N_3150,N_4608);
and U5536 (N_5536,N_4398,N_2243);
or U5537 (N_5537,N_1195,N_3417);
nand U5538 (N_5538,N_4507,N_1820);
nand U5539 (N_5539,N_1772,N_1553);
and U5540 (N_5540,N_506,N_3078);
nor U5541 (N_5541,N_3051,N_1163);
nand U5542 (N_5542,N_4543,N_4804);
and U5543 (N_5543,N_4523,N_4343);
or U5544 (N_5544,N_1532,N_613);
nor U5545 (N_5545,N_735,N_1343);
nor U5546 (N_5546,N_3219,N_4383);
and U5547 (N_5547,N_1196,N_1177);
or U5548 (N_5548,N_432,N_577);
xor U5549 (N_5549,N_2386,N_797);
and U5550 (N_5550,N_4386,N_1735);
and U5551 (N_5551,N_1090,N_2569);
and U5552 (N_5552,N_2376,N_780);
xor U5553 (N_5553,N_2073,N_1453);
nand U5554 (N_5554,N_1561,N_454);
or U5555 (N_5555,N_1550,N_3761);
nor U5556 (N_5556,N_607,N_3525);
xor U5557 (N_5557,N_1780,N_2312);
or U5558 (N_5558,N_3444,N_2812);
and U5559 (N_5559,N_4595,N_4428);
xor U5560 (N_5560,N_4590,N_265);
nor U5561 (N_5561,N_4373,N_2983);
and U5562 (N_5562,N_2000,N_1547);
and U5563 (N_5563,N_945,N_748);
nor U5564 (N_5564,N_3579,N_4084);
nand U5565 (N_5565,N_1071,N_3002);
and U5566 (N_5566,N_3467,N_4929);
nand U5567 (N_5567,N_3077,N_4291);
or U5568 (N_5568,N_1125,N_544);
nand U5569 (N_5569,N_1015,N_884);
xor U5570 (N_5570,N_1442,N_1888);
xor U5571 (N_5571,N_3280,N_4612);
nor U5572 (N_5572,N_1540,N_69);
or U5573 (N_5573,N_4849,N_2004);
xor U5574 (N_5574,N_1505,N_2040);
nand U5575 (N_5575,N_853,N_2255);
or U5576 (N_5576,N_3454,N_3928);
nand U5577 (N_5577,N_4235,N_1794);
nor U5578 (N_5578,N_439,N_818);
and U5579 (N_5579,N_570,N_3951);
nand U5580 (N_5580,N_1172,N_4682);
or U5581 (N_5581,N_622,N_4626);
and U5582 (N_5582,N_3282,N_1357);
and U5583 (N_5583,N_2182,N_2142);
nor U5584 (N_5584,N_1091,N_3753);
nor U5585 (N_5585,N_4466,N_4942);
or U5586 (N_5586,N_2259,N_2656);
and U5587 (N_5587,N_509,N_2824);
nor U5588 (N_5588,N_3631,N_3888);
nor U5589 (N_5589,N_2132,N_4869);
nand U5590 (N_5590,N_2681,N_3739);
nor U5591 (N_5591,N_4277,N_983);
xor U5592 (N_5592,N_1714,N_1432);
xor U5593 (N_5593,N_3853,N_2170);
nand U5594 (N_5594,N_4092,N_4371);
or U5595 (N_5595,N_847,N_4800);
nand U5596 (N_5596,N_2293,N_3379);
and U5597 (N_5597,N_3320,N_203);
and U5598 (N_5598,N_4557,N_1542);
nand U5599 (N_5599,N_1892,N_1079);
and U5600 (N_5600,N_1340,N_3810);
nand U5601 (N_5601,N_1670,N_4042);
nand U5602 (N_5602,N_1067,N_1100);
nor U5603 (N_5603,N_1718,N_3715);
nand U5604 (N_5604,N_2559,N_169);
nor U5605 (N_5605,N_3152,N_1451);
or U5606 (N_5606,N_3858,N_3272);
and U5607 (N_5607,N_1874,N_4296);
and U5608 (N_5608,N_599,N_3122);
or U5609 (N_5609,N_409,N_171);
xnor U5610 (N_5610,N_3998,N_1457);
or U5611 (N_5611,N_1292,N_4167);
nand U5612 (N_5612,N_4336,N_119);
nor U5613 (N_5613,N_4542,N_1371);
and U5614 (N_5614,N_2662,N_3996);
or U5615 (N_5615,N_1375,N_2582);
xor U5616 (N_5616,N_1041,N_3369);
nor U5617 (N_5617,N_2522,N_3404);
and U5618 (N_5618,N_4879,N_3840);
xnor U5619 (N_5619,N_150,N_4021);
xnor U5620 (N_5620,N_4113,N_342);
nor U5621 (N_5621,N_3226,N_2960);
nor U5622 (N_5622,N_1235,N_2528);
and U5623 (N_5623,N_1356,N_3632);
nor U5624 (N_5624,N_3194,N_4725);
nor U5625 (N_5625,N_25,N_405);
nor U5626 (N_5626,N_781,N_3200);
xor U5627 (N_5627,N_1230,N_4444);
xor U5628 (N_5628,N_4778,N_431);
nor U5629 (N_5629,N_1767,N_1361);
nor U5630 (N_5630,N_3105,N_2009);
xor U5631 (N_5631,N_3751,N_1030);
or U5632 (N_5632,N_4079,N_4921);
nand U5633 (N_5633,N_3228,N_3592);
nor U5634 (N_5634,N_352,N_3084);
nor U5635 (N_5635,N_1907,N_2019);
nand U5636 (N_5636,N_507,N_1681);
and U5637 (N_5637,N_3465,N_2508);
and U5638 (N_5638,N_3795,N_1113);
nand U5639 (N_5639,N_542,N_1302);
nand U5640 (N_5640,N_1610,N_3741);
and U5641 (N_5641,N_1322,N_1096);
nand U5642 (N_5642,N_3595,N_3111);
and U5643 (N_5643,N_4588,N_2204);
nand U5644 (N_5644,N_3035,N_327);
and U5645 (N_5645,N_2108,N_2117);
and U5646 (N_5646,N_4183,N_208);
xnor U5647 (N_5647,N_37,N_701);
nand U5648 (N_5648,N_3109,N_2436);
nand U5649 (N_5649,N_4177,N_283);
or U5650 (N_5650,N_3336,N_383);
nand U5651 (N_5651,N_3916,N_4062);
nand U5652 (N_5652,N_1563,N_1498);
xor U5653 (N_5653,N_4356,N_4203);
and U5654 (N_5654,N_1248,N_3463);
and U5655 (N_5655,N_4446,N_1600);
nand U5656 (N_5656,N_1321,N_230);
nand U5657 (N_5657,N_1319,N_2327);
nand U5658 (N_5658,N_3719,N_3296);
or U5659 (N_5659,N_1756,N_760);
nand U5660 (N_5660,N_4550,N_4659);
or U5661 (N_5661,N_3070,N_430);
xnor U5662 (N_5662,N_4240,N_3112);
and U5663 (N_5663,N_2191,N_2267);
and U5664 (N_5664,N_2506,N_1293);
and U5665 (N_5665,N_894,N_2013);
or U5666 (N_5666,N_4981,N_2439);
and U5667 (N_5667,N_2517,N_2119);
and U5668 (N_5668,N_3540,N_2074);
or U5669 (N_5669,N_3628,N_3672);
or U5670 (N_5670,N_2068,N_4890);
nor U5671 (N_5671,N_1109,N_3123);
or U5672 (N_5672,N_3697,N_2305);
and U5673 (N_5673,N_2899,N_3270);
nor U5674 (N_5674,N_849,N_3952);
xor U5675 (N_5675,N_3965,N_940);
nor U5676 (N_5676,N_715,N_1012);
nor U5677 (N_5677,N_3410,N_2443);
or U5678 (N_5678,N_1472,N_2323);
or U5679 (N_5679,N_2959,N_322);
or U5680 (N_5680,N_556,N_1496);
and U5681 (N_5681,N_3759,N_2279);
xor U5682 (N_5682,N_4757,N_2310);
and U5683 (N_5683,N_1560,N_4227);
nor U5684 (N_5684,N_1178,N_4081);
nand U5685 (N_5685,N_3939,N_845);
and U5686 (N_5686,N_4114,N_588);
nor U5687 (N_5687,N_591,N_1749);
and U5688 (N_5688,N_749,N_4961);
or U5689 (N_5689,N_4232,N_961);
and U5690 (N_5690,N_934,N_3452);
nand U5691 (N_5691,N_3003,N_2487);
nand U5692 (N_5692,N_2417,N_129);
nor U5693 (N_5693,N_3266,N_4239);
or U5694 (N_5694,N_4990,N_1450);
xor U5695 (N_5695,N_3775,N_3961);
nor U5696 (N_5696,N_442,N_3922);
or U5697 (N_5697,N_1527,N_512);
or U5698 (N_5698,N_1848,N_1660);
nand U5699 (N_5699,N_3235,N_2303);
and U5700 (N_5700,N_1700,N_3676);
nor U5701 (N_5701,N_4158,N_191);
or U5702 (N_5702,N_1531,N_441);
nor U5703 (N_5703,N_673,N_62);
nand U5704 (N_5704,N_3382,N_1430);
or U5705 (N_5705,N_1768,N_4155);
xor U5706 (N_5706,N_912,N_4436);
nand U5707 (N_5707,N_451,N_3982);
nor U5708 (N_5708,N_3286,N_2233);
nand U5709 (N_5709,N_3180,N_4404);
nor U5710 (N_5710,N_4292,N_3395);
xor U5711 (N_5711,N_1471,N_1853);
nand U5712 (N_5712,N_4923,N_3015);
nor U5713 (N_5713,N_4012,N_1223);
or U5714 (N_5714,N_2198,N_39);
nand U5715 (N_5715,N_3956,N_3365);
xnor U5716 (N_5716,N_4135,N_3042);
or U5717 (N_5717,N_1976,N_193);
nor U5718 (N_5718,N_3556,N_4193);
and U5719 (N_5719,N_4946,N_3407);
and U5720 (N_5720,N_1087,N_4889);
or U5721 (N_5721,N_1483,N_244);
and U5722 (N_5722,N_2665,N_2144);
or U5723 (N_5723,N_3211,N_3350);
nor U5724 (N_5724,N_1510,N_1253);
nand U5725 (N_5725,N_2141,N_176);
and U5726 (N_5726,N_4517,N_2453);
or U5727 (N_5727,N_4055,N_4211);
nand U5728 (N_5728,N_1407,N_2364);
nand U5729 (N_5729,N_3071,N_2971);
nand U5730 (N_5730,N_1981,N_3298);
xor U5731 (N_5731,N_871,N_4962);
nand U5732 (N_5732,N_2471,N_2133);
or U5733 (N_5733,N_844,N_3828);
nor U5734 (N_5734,N_2295,N_1020);
or U5735 (N_5735,N_3573,N_1632);
or U5736 (N_5736,N_1072,N_2221);
or U5737 (N_5737,N_2466,N_4144);
or U5738 (N_5738,N_566,N_1026);
nand U5739 (N_5739,N_1915,N_2926);
and U5740 (N_5740,N_2799,N_569);
nor U5741 (N_5741,N_1057,N_706);
and U5742 (N_5742,N_708,N_1497);
or U5743 (N_5743,N_59,N_1875);
xnor U5744 (N_5744,N_3995,N_4905);
or U5745 (N_5745,N_4749,N_695);
or U5746 (N_5746,N_3698,N_2111);
and U5747 (N_5747,N_4603,N_1899);
and U5748 (N_5748,N_4248,N_1389);
and U5749 (N_5749,N_3788,N_2779);
or U5750 (N_5750,N_2951,N_1953);
and U5751 (N_5751,N_793,N_4391);
or U5752 (N_5752,N_643,N_979);
nor U5753 (N_5753,N_12,N_2608);
or U5754 (N_5754,N_2333,N_1671);
nor U5755 (N_5755,N_3126,N_1946);
nand U5756 (N_5756,N_475,N_1654);
xnor U5757 (N_5757,N_552,N_876);
or U5758 (N_5758,N_1504,N_3500);
nand U5759 (N_5759,N_4482,N_11);
nor U5760 (N_5760,N_296,N_2938);
nor U5761 (N_5761,N_2691,N_2882);
or U5762 (N_5762,N_3553,N_4026);
and U5763 (N_5763,N_2128,N_1599);
or U5764 (N_5764,N_1103,N_3028);
and U5765 (N_5765,N_4960,N_2430);
nor U5766 (N_5766,N_4572,N_3942);
or U5767 (N_5767,N_3217,N_4069);
xnor U5768 (N_5768,N_4478,N_1080);
or U5769 (N_5769,N_4260,N_644);
or U5770 (N_5770,N_1351,N_2819);
xnor U5771 (N_5771,N_2916,N_40);
nand U5772 (N_5772,N_825,N_3790);
or U5773 (N_5773,N_1693,N_561);
and U5774 (N_5774,N_2395,N_3401);
and U5775 (N_5775,N_4888,N_1349);
nand U5776 (N_5776,N_2367,N_1438);
or U5777 (N_5777,N_3128,N_4341);
or U5778 (N_5778,N_94,N_4988);
nand U5779 (N_5779,N_4376,N_2568);
or U5780 (N_5780,N_1470,N_4319);
or U5781 (N_5781,N_4172,N_850);
and U5782 (N_5782,N_2834,N_4587);
and U5783 (N_5783,N_3677,N_260);
nand U5784 (N_5784,N_2637,N_3752);
nor U5785 (N_5785,N_3798,N_1154);
nand U5786 (N_5786,N_4189,N_1790);
or U5787 (N_5787,N_3978,N_1007);
nand U5788 (N_5788,N_2776,N_2804);
nand U5789 (N_5789,N_134,N_761);
xor U5790 (N_5790,N_2425,N_2792);
nor U5791 (N_5791,N_4655,N_1674);
and U5792 (N_5792,N_1835,N_3935);
and U5793 (N_5793,N_4362,N_2205);
and U5794 (N_5794,N_3257,N_4775);
or U5795 (N_5795,N_1465,N_3034);
nand U5796 (N_5796,N_1017,N_3073);
nand U5797 (N_5797,N_1330,N_2628);
and U5798 (N_5798,N_3081,N_2531);
xnor U5799 (N_5799,N_1692,N_3530);
nor U5800 (N_5800,N_2181,N_1400);
nor U5801 (N_5801,N_3103,N_1467);
nand U5802 (N_5802,N_3254,N_4454);
nor U5803 (N_5803,N_3897,N_3206);
nand U5804 (N_5804,N_2072,N_576);
and U5805 (N_5805,N_482,N_3136);
and U5806 (N_5806,N_1213,N_2134);
or U5807 (N_5807,N_201,N_406);
and U5808 (N_5808,N_4900,N_535);
or U5809 (N_5809,N_4531,N_1877);
xnor U5810 (N_5810,N_1774,N_4705);
nand U5811 (N_5811,N_4875,N_1379);
and U5812 (N_5812,N_3583,N_2114);
nor U5813 (N_5813,N_2581,N_2311);
or U5814 (N_5814,N_1492,N_3329);
nand U5815 (N_5815,N_1309,N_1120);
and U5816 (N_5816,N_4200,N_4322);
nor U5817 (N_5817,N_2958,N_4540);
nor U5818 (N_5818,N_279,N_4639);
nand U5819 (N_5819,N_992,N_3362);
or U5820 (N_5820,N_1307,N_4427);
nand U5821 (N_5821,N_2650,N_4262);
xnor U5822 (N_5822,N_4392,N_4582);
or U5823 (N_5823,N_2726,N_1146);
nand U5824 (N_5824,N_1479,N_2145);
and U5825 (N_5825,N_3373,N_2672);
and U5826 (N_5826,N_718,N_1900);
nand U5827 (N_5827,N_1410,N_4866);
nor U5828 (N_5828,N_3384,N_315);
nand U5829 (N_5829,N_1615,N_2573);
nand U5830 (N_5830,N_1134,N_436);
and U5831 (N_5831,N_493,N_2319);
and U5832 (N_5832,N_2419,N_1055);
and U5833 (N_5833,N_1228,N_4976);
nor U5834 (N_5834,N_813,N_2635);
or U5835 (N_5835,N_930,N_4968);
or U5836 (N_5836,N_3911,N_1269);
xor U5837 (N_5837,N_4525,N_1619);
nor U5838 (N_5838,N_38,N_3580);
or U5839 (N_5839,N_456,N_1301);
or U5840 (N_5840,N_2521,N_4263);
and U5841 (N_5841,N_3590,N_3163);
nor U5842 (N_5842,N_1396,N_1431);
or U5843 (N_5843,N_3367,N_4352);
and U5844 (N_5844,N_2384,N_247);
and U5845 (N_5845,N_4643,N_4396);
nand U5846 (N_5846,N_1306,N_4644);
or U5847 (N_5847,N_4538,N_4279);
and U5848 (N_5848,N_1672,N_2712);
or U5849 (N_5849,N_4093,N_3239);
nor U5850 (N_5850,N_4665,N_1796);
nand U5851 (N_5851,N_4827,N_4868);
or U5852 (N_5852,N_3149,N_1612);
xnor U5853 (N_5853,N_2942,N_4072);
or U5854 (N_5854,N_4792,N_2116);
nor U5855 (N_5855,N_4536,N_415);
xor U5856 (N_5856,N_2492,N_1037);
and U5857 (N_5857,N_4640,N_4186);
nand U5858 (N_5858,N_1288,N_127);
or U5859 (N_5859,N_2138,N_2336);
xor U5860 (N_5860,N_4268,N_3285);
nor U5861 (N_5861,N_3574,N_4681);
and U5862 (N_5862,N_2606,N_2727);
or U5863 (N_5863,N_4121,N_97);
nand U5864 (N_5864,N_2451,N_1895);
nor U5865 (N_5865,N_3183,N_631);
or U5866 (N_5866,N_3723,N_3669);
nand U5867 (N_5867,N_4048,N_2936);
xor U5868 (N_5868,N_3843,N_4499);
and U5869 (N_5869,N_3050,N_3393);
or U5870 (N_5870,N_1948,N_3155);
nor U5871 (N_5871,N_4700,N_729);
or U5872 (N_5872,N_866,N_2922);
nand U5873 (N_5873,N_3162,N_1684);
and U5874 (N_5874,N_242,N_1555);
nor U5875 (N_5875,N_2782,N_2554);
nand U5876 (N_5876,N_2462,N_2131);
nor U5877 (N_5877,N_3213,N_2118);
and U5878 (N_5878,N_4471,N_727);
nor U5879 (N_5879,N_2452,N_3319);
xnor U5880 (N_5880,N_4095,N_2129);
nand U5881 (N_5881,N_4327,N_3392);
nand U5882 (N_5882,N_2788,N_1517);
and U5883 (N_5883,N_1609,N_3259);
and U5884 (N_5884,N_2250,N_3234);
nor U5885 (N_5885,N_2440,N_450);
or U5886 (N_5886,N_14,N_4340);
nand U5887 (N_5887,N_4101,N_2410);
nand U5888 (N_5888,N_3438,N_1635);
or U5889 (N_5889,N_2095,N_1129);
and U5890 (N_5890,N_437,N_2561);
nor U5891 (N_5891,N_4115,N_3883);
nor U5892 (N_5892,N_4360,N_3216);
or U5893 (N_5893,N_2653,N_2841);
or U5894 (N_5894,N_2136,N_1207);
nor U5895 (N_5895,N_635,N_3936);
xnor U5896 (N_5896,N_1209,N_1871);
or U5897 (N_5897,N_4585,N_4258);
xnor U5898 (N_5898,N_3080,N_1903);
xnor U5899 (N_5899,N_3893,N_233);
and U5900 (N_5900,N_1513,N_4311);
xor U5901 (N_5901,N_4118,N_598);
nand U5902 (N_5902,N_4198,N_2306);
and U5903 (N_5903,N_363,N_1658);
and U5904 (N_5904,N_3572,N_501);
nand U5905 (N_5905,N_777,N_3275);
or U5906 (N_5906,N_4564,N_4236);
and U5907 (N_5907,N_254,N_177);
or U5908 (N_5908,N_4722,N_4653);
or U5909 (N_5909,N_3125,N_3954);
nand U5910 (N_5910,N_1215,N_1523);
xnor U5911 (N_5911,N_3258,N_1184);
or U5912 (N_5912,N_3361,N_75);
nor U5913 (N_5913,N_605,N_2302);
nand U5914 (N_5914,N_389,N_1727);
nand U5915 (N_5915,N_2785,N_1234);
or U5916 (N_5916,N_3383,N_433);
and U5917 (N_5917,N_1161,N_4073);
and U5918 (N_5918,N_4750,N_337);
xnor U5919 (N_5919,N_3223,N_67);
and U5920 (N_5920,N_3072,N_4202);
nand U5921 (N_5921,N_1844,N_1816);
nand U5922 (N_5922,N_4887,N_2281);
or U5923 (N_5923,N_1901,N_269);
and U5924 (N_5924,N_1558,N_4381);
nand U5925 (N_5925,N_3726,N_4716);
nor U5926 (N_5926,N_4632,N_789);
or U5927 (N_5927,N_3118,N_1211);
and U5928 (N_5928,N_1689,N_74);
nor U5929 (N_5929,N_4742,N_1419);
and U5930 (N_5930,N_416,N_682);
nand U5931 (N_5931,N_3487,N_1805);
nor U5932 (N_5932,N_486,N_2071);
nand U5933 (N_5933,N_1663,N_938);
nand U5934 (N_5934,N_872,N_4966);
nand U5935 (N_5935,N_4107,N_3058);
xnor U5936 (N_5936,N_2739,N_3908);
and U5937 (N_5937,N_1294,N_3919);
nor U5938 (N_5938,N_4355,N_1135);
nand U5939 (N_5939,N_2978,N_287);
or U5940 (N_5940,N_3508,N_4971);
nand U5941 (N_5941,N_3119,N_4794);
nand U5942 (N_5942,N_4503,N_1426);
or U5943 (N_5943,N_3475,N_298);
nor U5944 (N_5944,N_1999,N_3143);
or U5945 (N_5945,N_4761,N_4891);
nor U5946 (N_5946,N_2986,N_3480);
nor U5947 (N_5947,N_1908,N_1164);
nor U5948 (N_5948,N_440,N_2213);
nand U5949 (N_5949,N_2630,N_2849);
or U5950 (N_5950,N_1412,N_1795);
or U5951 (N_5951,N_1778,N_782);
or U5952 (N_5952,N_1369,N_924);
or U5953 (N_5953,N_1494,N_3188);
nor U5954 (N_5954,N_3627,N_4920);
or U5955 (N_5955,N_3794,N_4777);
nor U5956 (N_5956,N_993,N_3231);
and U5957 (N_5957,N_860,N_505);
xnor U5958 (N_5958,N_2464,N_471);
and U5959 (N_5959,N_1715,N_3578);
and U5960 (N_5960,N_3861,N_4658);
nor U5961 (N_5961,N_2700,N_42);
and U5962 (N_5962,N_207,N_1896);
or U5963 (N_5963,N_1958,N_594);
or U5964 (N_5964,N_2085,N_1374);
nor U5965 (N_5965,N_1913,N_1180);
nor U5966 (N_5966,N_883,N_2699);
nand U5967 (N_5967,N_1633,N_2817);
nand U5968 (N_5968,N_2473,N_1992);
and U5969 (N_5969,N_736,N_572);
nor U5970 (N_5970,N_2290,N_3701);
xor U5971 (N_5971,N_4103,N_1696);
nor U5972 (N_5972,N_494,N_2100);
and U5973 (N_5973,N_2586,N_753);
nor U5974 (N_5974,N_1886,N_3754);
nand U5975 (N_5975,N_1956,N_2616);
nand U5976 (N_5976,N_2879,N_2163);
nor U5977 (N_5977,N_2850,N_372);
or U5978 (N_5978,N_4333,N_3377);
nand U5979 (N_5979,N_794,N_101);
nand U5980 (N_5980,N_2408,N_1249);
or U5981 (N_5981,N_4755,N_1585);
xnor U5982 (N_5982,N_1324,N_835);
nand U5983 (N_5983,N_1480,N_1752);
and U5984 (N_5984,N_2968,N_1551);
or U5985 (N_5985,N_1247,N_4877);
and U5986 (N_5986,N_3232,N_1488);
nand U5987 (N_5987,N_3779,N_2178);
or U5988 (N_5988,N_4669,N_3570);
and U5989 (N_5989,N_4024,N_4070);
and U5990 (N_5990,N_2211,N_4554);
and U5991 (N_5991,N_10,N_4280);
xnor U5992 (N_5992,N_4397,N_4030);
and U5993 (N_5993,N_1624,N_2651);
nor U5994 (N_5994,N_1245,N_4363);
nor U5995 (N_5995,N_3650,N_2778);
xor U5996 (N_5996,N_4860,N_1596);
nor U5997 (N_5997,N_2609,N_1106);
and U5998 (N_5998,N_2284,N_1830);
nand U5999 (N_5999,N_873,N_2411);
nor U6000 (N_6000,N_4067,N_2696);
nand U6001 (N_6001,N_3559,N_2874);
nand U6002 (N_6002,N_2935,N_769);
nor U6003 (N_6003,N_2708,N_4128);
nand U6004 (N_6004,N_1509,N_1150);
nand U6005 (N_6005,N_1564,N_4991);
nand U6006 (N_6006,N_3568,N_3518);
nand U6007 (N_6007,N_2224,N_248);
and U6008 (N_6008,N_4305,N_3929);
nor U6009 (N_6009,N_1529,N_1725);
nand U6010 (N_6010,N_3643,N_3007);
nand U6011 (N_6011,N_241,N_4561);
nor U6012 (N_6012,N_2209,N_4685);
or U6013 (N_6013,N_168,N_1227);
nand U6014 (N_6014,N_4119,N_1666);
or U6015 (N_6015,N_1023,N_1440);
or U6016 (N_6016,N_2018,N_1520);
nand U6017 (N_6017,N_985,N_2402);
nor U6018 (N_6018,N_3994,N_935);
or U6019 (N_6019,N_4056,N_1823);
nand U6020 (N_6020,N_1092,N_2130);
nand U6021 (N_6021,N_2442,N_2388);
and U6022 (N_6022,N_3616,N_3190);
or U6023 (N_6023,N_1315,N_3622);
xor U6024 (N_6024,N_3889,N_3944);
or U6025 (N_6025,N_114,N_1678);
xor U6026 (N_6026,N_2992,N_323);
nor U6027 (N_6027,N_2343,N_618);
and U6028 (N_6028,N_2615,N_540);
and U6029 (N_6029,N_2950,N_280);
or U6030 (N_6030,N_2529,N_2516);
or U6031 (N_6031,N_1139,N_1370);
or U6032 (N_6032,N_2765,N_601);
nor U6033 (N_6033,N_1546,N_343);
nor U6034 (N_6034,N_754,N_2596);
nand U6035 (N_6035,N_2499,N_3746);
nor U6036 (N_6036,N_2093,N_776);
and U6037 (N_6037,N_2676,N_929);
xnor U6038 (N_6038,N_4537,N_330);
or U6039 (N_6039,N_2359,N_4314);
and U6040 (N_6040,N_3315,N_4287);
or U6041 (N_6041,N_3647,N_4736);
and U6042 (N_6042,N_554,N_1902);
nor U6043 (N_6043,N_1909,N_1036);
and U6044 (N_6044,N_3433,N_1928);
or U6045 (N_6045,N_3116,N_4617);
or U6046 (N_6046,N_4023,N_3094);
or U6047 (N_6047,N_3423,N_1476);
nand U6048 (N_6048,N_2489,N_4410);
or U6049 (N_6049,N_3845,N_4388);
or U6050 (N_6050,N_284,N_4209);
or U6051 (N_6051,N_4719,N_1311);
nand U6052 (N_6052,N_3782,N_3411);
nor U6053 (N_6053,N_4218,N_1214);
and U6054 (N_6054,N_410,N_3364);
nor U6055 (N_6055,N_2836,N_1580);
and U6056 (N_6056,N_1420,N_911);
xnor U6057 (N_6057,N_2054,N_4345);
and U6058 (N_6058,N_1791,N_228);
xor U6059 (N_6059,N_4698,N_2659);
nand U6060 (N_6060,N_1720,N_3279);
and U6061 (N_6061,N_2906,N_2371);
nor U6062 (N_6062,N_994,N_374);
or U6063 (N_6063,N_2970,N_4668);
nand U6064 (N_6064,N_3192,N_3986);
xnor U6065 (N_6065,N_4754,N_656);
nor U6066 (N_6066,N_2155,N_3469);
and U6067 (N_6067,N_1308,N_375);
or U6068 (N_6068,N_4677,N_2077);
or U6069 (N_6069,N_4043,N_691);
and U6070 (N_6070,N_3049,N_1831);
or U6071 (N_6071,N_1506,N_2748);
nor U6072 (N_6072,N_2083,N_2810);
nand U6073 (N_6073,N_3943,N_1153);
xor U6074 (N_6074,N_0,N_3521);
nand U6075 (N_6075,N_411,N_2903);
and U6076 (N_6076,N_3085,N_2543);
nor U6077 (N_6077,N_3611,N_2614);
nand U6078 (N_6078,N_2230,N_1665);
or U6079 (N_6079,N_2820,N_2854);
nor U6080 (N_6080,N_1265,N_1263);
nor U6081 (N_6081,N_858,N_4842);
and U6082 (N_6082,N_4651,N_4367);
and U6083 (N_6083,N_95,N_488);
and U6084 (N_6084,N_548,N_16);
nor U6085 (N_6085,N_1912,N_3517);
nor U6086 (N_6086,N_1168,N_841);
nand U6087 (N_6087,N_3600,N_2887);
nor U6088 (N_6088,N_65,N_1448);
or U6089 (N_6089,N_3515,N_4029);
nand U6090 (N_6090,N_3037,N_2957);
nand U6091 (N_6091,N_412,N_3721);
nor U6092 (N_6092,N_2857,N_350);
xnor U6093 (N_6093,N_2422,N_1809);
nor U6094 (N_6094,N_2683,N_2943);
and U6095 (N_6095,N_3735,N_4892);
nor U6096 (N_6096,N_4989,N_3204);
nor U6097 (N_6097,N_190,N_2444);
or U6098 (N_6098,N_2459,N_1291);
nand U6099 (N_6099,N_4624,N_4154);
or U6100 (N_6100,N_901,N_272);
and U6101 (N_6101,N_4992,N_1380);
or U6102 (N_6102,N_2001,N_4282);
or U6103 (N_6103,N_1458,N_3018);
xor U6104 (N_6104,N_4385,N_1049);
and U6105 (N_6105,N_1416,N_1059);
or U6106 (N_6106,N_4299,N_2214);
or U6107 (N_6107,N_3096,N_4210);
and U6108 (N_6108,N_4307,N_3032);
nand U6109 (N_6109,N_291,N_3985);
nand U6110 (N_6110,N_2082,N_2851);
xor U6111 (N_6111,N_3783,N_2339);
xor U6112 (N_6112,N_3914,N_344);
nand U6113 (N_6113,N_2566,N_282);
nand U6114 (N_6114,N_4506,N_3356);
nor U6115 (N_6115,N_4491,N_3937);
nor U6116 (N_6116,N_3264,N_3990);
or U6117 (N_6117,N_1508,N_3876);
nor U6118 (N_6118,N_562,N_4694);
nor U6119 (N_6119,N_510,N_2035);
nor U6120 (N_6120,N_2172,N_2345);
nor U6121 (N_6121,N_1885,N_2146);
and U6122 (N_6122,N_388,N_3295);
xor U6123 (N_6123,N_539,N_481);
or U6124 (N_6124,N_2045,N_3571);
and U6125 (N_6125,N_393,N_4512);
xor U6126 (N_6126,N_2813,N_3901);
or U6127 (N_6127,N_524,N_473);
and U6128 (N_6128,N_3818,N_1341);
xor U6129 (N_6129,N_2975,N_2171);
nand U6130 (N_6130,N_956,N_694);
nand U6131 (N_6131,N_907,N_1760);
nand U6132 (N_6132,N_2789,N_4208);
xor U6133 (N_6133,N_2655,N_2329);
and U6134 (N_6134,N_3867,N_35);
nand U6135 (N_6135,N_1025,N_1344);
nor U6136 (N_6136,N_2385,N_156);
or U6137 (N_6137,N_1675,N_4445);
xor U6138 (N_6138,N_2658,N_4222);
xnor U6139 (N_6139,N_4452,N_4123);
or U6140 (N_6140,N_1239,N_4938);
and U6141 (N_6141,N_4434,N_1350);
nor U6142 (N_6142,N_4965,N_3493);
and U6143 (N_6143,N_2611,N_1358);
and U6144 (N_6144,N_2278,N_1982);
nor U6145 (N_6145,N_1337,N_4027);
nand U6146 (N_6146,N_3197,N_4957);
nand U6147 (N_6147,N_2203,N_2705);
nor U6148 (N_6148,N_802,N_1151);
nand U6149 (N_6149,N_3932,N_4745);
nand U6150 (N_6150,N_1501,N_349);
and U6151 (N_6151,N_3161,N_2298);
and U6152 (N_6152,N_8,N_4519);
xnor U6153 (N_6153,N_692,N_4256);
and U6154 (N_6154,N_1664,N_2524);
and U6155 (N_6155,N_2752,N_1014);
xor U6156 (N_6156,N_4771,N_2217);
nor U6157 (N_6157,N_4106,N_3326);
or U6158 (N_6158,N_339,N_36);
nor U6159 (N_6159,N_2734,N_1991);
and U6160 (N_6160,N_2816,N_1690);
xor U6161 (N_6161,N_2382,N_1929);
and U6162 (N_6162,N_3704,N_2195);
nor U6163 (N_6163,N_980,N_3069);
nand U6164 (N_6164,N_4851,N_1993);
or U6165 (N_6165,N_249,N_653);
nand U6166 (N_6166,N_4618,N_3090);
nor U6167 (N_6167,N_4045,N_2891);
nor U6168 (N_6168,N_4605,N_1771);
and U6169 (N_6169,N_1111,N_1906);
and U6170 (N_6170,N_1711,N_1428);
and U6171 (N_6171,N_1149,N_2853);
or U6172 (N_6172,N_2494,N_1846);
xnor U6173 (N_6173,N_4077,N_626);
and U6174 (N_6174,N_2268,N_83);
or U6175 (N_6175,N_4708,N_558);
and U6176 (N_6176,N_865,N_4429);
or U6177 (N_6177,N_1792,N_84);
nand U6178 (N_6178,N_3973,N_1972);
or U6179 (N_6179,N_4735,N_2357);
and U6180 (N_6180,N_1786,N_2894);
or U6181 (N_6181,N_1987,N_3130);
and U6182 (N_6182,N_597,N_1611);
or U6183 (N_6183,N_3496,N_1101);
xor U6184 (N_6184,N_3582,N_2081);
nor U6185 (N_6185,N_3387,N_663);
and U6186 (N_6186,N_909,N_3968);
nor U6187 (N_6187,N_4261,N_513);
nor U6188 (N_6188,N_2275,N_364);
nand U6189 (N_6189,N_4411,N_4847);
nand U6190 (N_6190,N_4737,N_4038);
or U6191 (N_6191,N_3668,N_4648);
or U6192 (N_6192,N_4390,N_1782);
xor U6193 (N_6193,N_2162,N_1219);
or U6194 (N_6194,N_1519,N_767);
or U6195 (N_6195,N_4837,N_4730);
nand U6196 (N_6196,N_1841,N_3909);
or U6197 (N_6197,N_2159,N_311);
nand U6198 (N_6198,N_2982,N_2940);
or U6199 (N_6199,N_809,N_2640);
and U6200 (N_6200,N_1966,N_362);
and U6201 (N_6201,N_3386,N_2909);
nor U6202 (N_6202,N_1631,N_1962);
xnor U6203 (N_6203,N_2945,N_3008);
or U6204 (N_6204,N_53,N_2558);
or U6205 (N_6205,N_485,N_511);
nor U6206 (N_6206,N_3767,N_4181);
nand U6207 (N_6207,N_2387,N_4687);
nor U6208 (N_6208,N_4844,N_3240);
and U6209 (N_6209,N_915,N_4836);
nand U6210 (N_6210,N_2434,N_807);
nand U6211 (N_6211,N_1889,N_4621);
nand U6212 (N_6212,N_2415,N_2241);
nor U6213 (N_6213,N_368,N_4575);
nor U6214 (N_6214,N_770,N_4784);
nand U6215 (N_6215,N_4285,N_3359);
and U6216 (N_6216,N_1818,N_803);
and U6217 (N_6217,N_2347,N_2829);
xor U6218 (N_6218,N_2479,N_4028);
xnor U6219 (N_6219,N_4720,N_2612);
and U6220 (N_6220,N_3601,N_1193);
or U6221 (N_6221,N_340,N_4809);
and U6222 (N_6222,N_2602,N_474);
nor U6223 (N_6223,N_2547,N_2109);
nor U6224 (N_6224,N_1868,N_224);
nor U6225 (N_6225,N_4347,N_2883);
xnor U6226 (N_6226,N_1813,N_2831);
and U6227 (N_6227,N_933,N_3699);
and U6228 (N_6228,N_4592,N_60);
nor U6229 (N_6229,N_1937,N_4692);
nor U6230 (N_6230,N_4883,N_2029);
nand U6231 (N_6231,N_2416,N_2021);
nand U6232 (N_6232,N_2350,N_1031);
nand U6233 (N_6233,N_1183,N_1750);
xor U6234 (N_6234,N_122,N_2017);
nand U6235 (N_6235,N_3934,N_4300);
and U6236 (N_6236,N_1724,N_3718);
or U6237 (N_6237,N_3763,N_1810);
nor U6238 (N_6238,N_4856,N_258);
and U6239 (N_6239,N_3660,N_2876);
or U6240 (N_6240,N_2256,N_1035);
xnor U6241 (N_6241,N_864,N_3917);
or U6242 (N_6242,N_3814,N_4895);
or U6243 (N_6243,N_3151,N_4823);
and U6244 (N_6244,N_1128,N_3054);
and U6245 (N_6245,N_4584,N_1572);
nand U6246 (N_6246,N_538,N_1603);
nand U6247 (N_6247,N_1063,N_1425);
or U6248 (N_6248,N_3460,N_3331);
nand U6249 (N_6249,N_689,N_2449);
or U6250 (N_6250,N_3288,N_2811);
and U6251 (N_6251,N_4005,N_140);
nand U6252 (N_6252,N_329,N_1489);
xor U6253 (N_6253,N_3045,N_3663);
xor U6254 (N_6254,N_3756,N_4711);
or U6255 (N_6255,N_4271,N_3027);
and U6256 (N_6256,N_1702,N_2793);
xnor U6257 (N_6257,N_4486,N_2261);
nand U6258 (N_6258,N_680,N_1605);
nor U6259 (N_6259,N_973,N_3159);
nor U6260 (N_6260,N_739,N_4169);
and U6261 (N_6261,N_4485,N_2481);
or U6262 (N_6262,N_964,N_709);
nor U6263 (N_6263,N_1175,N_237);
or U6264 (N_6264,N_3963,N_1710);
nor U6265 (N_6265,N_3422,N_3953);
and U6266 (N_6266,N_4912,N_2838);
nor U6267 (N_6267,N_1801,N_1986);
nor U6268 (N_6268,N_2607,N_3312);
nand U6269 (N_6269,N_4053,N_2041);
nand U6270 (N_6270,N_2781,N_831);
or U6271 (N_6271,N_4050,N_3229);
and U6272 (N_6272,N_386,N_1571);
and U6273 (N_6273,N_699,N_3921);
nand U6274 (N_6274,N_3311,N_3247);
and U6275 (N_6275,N_1404,N_3613);
nand U6276 (N_6276,N_890,N_3524);
or U6277 (N_6277,N_1573,N_917);
and U6278 (N_6278,N_4270,N_3262);
nand U6279 (N_6279,N_1065,N_1828);
or U6280 (N_6280,N_143,N_2673);
and U6281 (N_6281,N_4638,N_369);
or U6282 (N_6282,N_674,N_632);
nor U6283 (N_6283,N_3659,N_4846);
or U6284 (N_6284,N_2600,N_658);
nor U6285 (N_6285,N_1515,N_2796);
nor U6286 (N_6286,N_1002,N_4977);
nand U6287 (N_6287,N_4738,N_2930);
and U6288 (N_6288,N_1189,N_833);
nor U6289 (N_6289,N_4364,N_2783);
or U6290 (N_6290,N_3591,N_4650);
and U6291 (N_6291,N_2190,N_3177);
and U6292 (N_6292,N_1027,N_1403);
or U6293 (N_6293,N_3483,N_3225);
nand U6294 (N_6294,N_799,N_4734);
nor U6295 (N_6295,N_4313,N_2038);
or U6296 (N_6296,N_288,N_3440);
or U6297 (N_6297,N_2078,N_3870);
and U6298 (N_6298,N_4637,N_3453);
xor U6299 (N_6299,N_49,N_2721);
xor U6300 (N_6300,N_4213,N_3302);
nand U6301 (N_6301,N_4358,N_3256);
xnor U6302 (N_6302,N_1406,N_1581);
and U6303 (N_6303,N_1821,N_3838);
or U6304 (N_6304,N_4377,N_1383);
xnor U6305 (N_6305,N_4054,N_56);
xnor U6306 (N_6306,N_2617,N_861);
nor U6307 (N_6307,N_2741,N_4408);
and U6308 (N_6308,N_1148,N_212);
xnor U6309 (N_6309,N_2226,N_703);
nor U6310 (N_6310,N_217,N_225);
and U6311 (N_6311,N_2826,N_4475);
nand U6312 (N_6312,N_1105,N_4940);
nor U6313 (N_6313,N_2096,N_2638);
nor U6314 (N_6314,N_721,N_4096);
nor U6315 (N_6315,N_4245,N_3679);
nand U6316 (N_6316,N_2285,N_4780);
and U6317 (N_6317,N_1478,N_1649);
and U6318 (N_6318,N_1882,N_3977);
and U6319 (N_6319,N_2549,N_3271);
and U6320 (N_6320,N_64,N_1943);
and U6321 (N_6321,N_1751,N_385);
or U6322 (N_6322,N_1832,N_3341);
and U6323 (N_6323,N_2047,N_33);
xor U6324 (N_6324,N_719,N_2546);
xnor U6325 (N_6325,N_3971,N_4489);
xnor U6326 (N_6326,N_575,N_3702);
nand U6327 (N_6327,N_1166,N_4689);
or U6328 (N_6328,N_2707,N_4500);
nor U6329 (N_6329,N_1621,N_3550);
nor U6330 (N_6330,N_2801,N_3429);
nand U6331 (N_6331,N_1697,N_4146);
or U6332 (N_6332,N_3906,N_4803);
and U6333 (N_6333,N_4421,N_3363);
nand U6334 (N_6334,N_3705,N_1048);
nor U6335 (N_6335,N_1348,N_600);
or U6336 (N_6336,N_2299,N_1147);
nand U6337 (N_6337,N_479,N_4602);
nor U6338 (N_6338,N_262,N_4326);
and U6339 (N_6339,N_823,N_1955);
nor U6340 (N_6340,N_1443,N_2652);
xnor U6341 (N_6341,N_3913,N_1740);
nand U6342 (N_6342,N_916,N_4825);
nand U6343 (N_6343,N_1800,N_914);
or U6344 (N_6344,N_2825,N_4599);
nand U6345 (N_6345,N_2733,N_4199);
nor U6346 (N_6346,N_1243,N_4451);
nand U6347 (N_6347,N_1347,N_586);
nand U6348 (N_6348,N_4882,N_4834);
or U6349 (N_6349,N_77,N_3873);
nand U6350 (N_6350,N_4509,N_157);
nor U6351 (N_6351,N_856,N_2112);
xor U6352 (N_6352,N_3833,N_947);
nor U6353 (N_6353,N_3505,N_29);
and U6354 (N_6354,N_462,N_341);
nand U6355 (N_6355,N_2896,N_170);
nand U6356 (N_6356,N_3299,N_3263);
nor U6357 (N_6357,N_110,N_3132);
or U6358 (N_6358,N_1185,N_811);
and U6359 (N_6359,N_620,N_4776);
or U6360 (N_6360,N_78,N_85);
nand U6361 (N_6361,N_1932,N_2773);
and U6362 (N_6362,N_1977,N_3491);
nor U6363 (N_6363,N_3807,N_497);
nand U6364 (N_6364,N_3499,N_4008);
and U6365 (N_6365,N_404,N_445);
or U6366 (N_6366,N_4295,N_206);
nor U6367 (N_6367,N_3399,N_4458);
or U6368 (N_6368,N_3115,N_816);
nand U6369 (N_6369,N_3175,N_3748);
or U6370 (N_6370,N_1918,N_4956);
nor U6371 (N_6371,N_2301,N_1312);
nand U6372 (N_6372,N_553,N_974);
or U6373 (N_6373,N_4964,N_2898);
nand U6374 (N_6374,N_636,N_1003);
nand U6375 (N_6375,N_730,N_855);
or U6376 (N_6376,N_4852,N_4472);
and U6377 (N_6377,N_4748,N_571);
or U6378 (N_6378,N_159,N_2098);
xor U6379 (N_6379,N_4696,N_4829);
nor U6380 (N_6380,N_2814,N_2579);
or U6381 (N_6381,N_3310,N_3343);
and U6382 (N_6382,N_3607,N_3278);
xnor U6383 (N_6383,N_4573,N_4947);
and U6384 (N_6384,N_2750,N_1719);
and U6385 (N_6385,N_1452,N_3757);
nand U6386 (N_6386,N_2886,N_815);
nand U6387 (N_6387,N_3877,N_2137);
nand U6388 (N_6388,N_2394,N_1118);
or U6389 (N_6389,N_4433,N_1381);
nand U6390 (N_6390,N_1436,N_174);
nand U6391 (N_6391,N_2208,N_2666);
xnor U6392 (N_6392,N_3426,N_2947);
nand U6393 (N_6393,N_2180,N_2107);
and U6394 (N_6394,N_1628,N_1366);
nand U6395 (N_6395,N_931,N_4897);
nor U6396 (N_6396,N_4975,N_2273);
nor U6397 (N_6397,N_1798,N_4125);
nand U6398 (N_6398,N_4286,N_425);
nand U6399 (N_6399,N_647,N_1064);
nand U6400 (N_6400,N_2856,N_3799);
nor U6401 (N_6401,N_887,N_4464);
and U6402 (N_6402,N_2215,N_4171);
and U6403 (N_6403,N_1075,N_2488);
and U6404 (N_6404,N_3874,N_652);
nor U6405 (N_6405,N_4547,N_3405);
xnor U6406 (N_6406,N_2613,N_3629);
nand U6407 (N_6407,N_3021,N_3485);
xnor U6408 (N_6408,N_4993,N_2830);
nand U6409 (N_6409,N_2872,N_1491);
nor U6410 (N_6410,N_543,N_1769);
xnor U6411 (N_6411,N_1787,N_398);
nor U6412 (N_6412,N_3100,N_3274);
nor U6413 (N_6413,N_1208,N_3209);
or U6414 (N_6414,N_4188,N_764);
or U6415 (N_6415,N_253,N_1652);
nand U6416 (N_6416,N_2525,N_3237);
and U6417 (N_6417,N_1824,N_1747);
nand U6418 (N_6418,N_3821,N_2818);
nor U6419 (N_6419,N_1533,N_4297);
or U6420 (N_6420,N_243,N_1682);
and U6421 (N_6421,N_1004,N_4715);
nor U6422 (N_6422,N_1645,N_2767);
nand U6423 (N_6423,N_4680,N_4799);
nor U6424 (N_6424,N_2428,N_3618);
nor U6425 (N_6425,N_3179,N_1385);
nor U6426 (N_6426,N_3700,N_2264);
nor U6427 (N_6427,N_5,N_1274);
or U6428 (N_6428,N_3842,N_3923);
and U6429 (N_6429,N_1701,N_214);
nor U6430 (N_6430,N_2398,N_3445);
or U6431 (N_6431,N_2588,N_3145);
nand U6432 (N_6432,N_4288,N_392);
nand U6433 (N_6433,N_1618,N_2928);
nor U6434 (N_6434,N_4817,N_4945);
nor U6435 (N_6435,N_1604,N_1704);
or U6436 (N_6436,N_3528,N_1588);
nor U6437 (N_6437,N_4353,N_4717);
nor U6438 (N_6438,N_4372,N_869);
or U6439 (N_6439,N_4752,N_141);
xnor U6440 (N_6440,N_325,N_204);
xor U6441 (N_6441,N_4086,N_1422);
xor U6442 (N_6442,N_426,N_859);
nor U6443 (N_6443,N_4636,N_1046);
nor U6444 (N_6444,N_2967,N_4461);
and U6445 (N_6445,N_2747,N_3964);
nor U6446 (N_6446,N_3164,N_2414);
or U6447 (N_6447,N_4165,N_1435);
nand U6448 (N_6448,N_1317,N_863);
and U6449 (N_6449,N_239,N_4163);
and U6450 (N_6450,N_1329,N_2317);
nor U6451 (N_6451,N_2062,N_3418);
nor U6452 (N_6452,N_4318,N_152);
nor U6453 (N_6453,N_4808,N_998);
and U6454 (N_6454,N_1942,N_4275);
nor U6455 (N_6455,N_2509,N_1765);
or U6456 (N_6456,N_2152,N_812);
or U6457 (N_6457,N_1202,N_2186);
nor U6458 (N_6458,N_3344,N_2827);
or U6459 (N_6459,N_3776,N_3871);
nor U6460 (N_6460,N_1753,N_3068);
or U6461 (N_6461,N_277,N_1804);
nor U6462 (N_6462,N_3339,N_1468);
and U6463 (N_6463,N_3884,N_70);
and U6464 (N_6464,N_3062,N_2289);
nand U6465 (N_6465,N_3186,N_734);
or U6466 (N_6466,N_4896,N_1198);
xnor U6467 (N_6467,N_3854,N_732);
or U6468 (N_6468,N_3110,N_3809);
nand U6469 (N_6469,N_1884,N_1698);
or U6470 (N_6470,N_2560,N_867);
or U6471 (N_6471,N_4040,N_3502);
nor U6472 (N_6472,N_2685,N_2331);
nor U6473 (N_6473,N_465,N_2033);
nand U6474 (N_6474,N_3412,N_616);
nand U6475 (N_6475,N_4303,N_1905);
nor U6476 (N_6476,N_2946,N_1095);
or U6477 (N_6477,N_246,N_4656);
nand U6478 (N_6478,N_1930,N_309);
nor U6479 (N_6479,N_3712,N_3030);
nor U6480 (N_6480,N_3800,N_2548);
nand U6481 (N_6481,N_602,N_2094);
xnor U6482 (N_6482,N_4818,N_1029);
nor U6483 (N_6483,N_982,N_4998);
nor U6484 (N_6484,N_4276,N_3218);
or U6485 (N_6485,N_1676,N_3293);
nor U6486 (N_6486,N_4853,N_4174);
nor U6487 (N_6487,N_4830,N_116);
or U6488 (N_6488,N_2407,N_1880);
nand U6489 (N_6489,N_824,N_2972);
xnor U6490 (N_6490,N_3227,N_371);
nor U6491 (N_6491,N_2984,N_4127);
nor U6492 (N_6492,N_1984,N_446);
nor U6493 (N_6493,N_2342,N_4870);
nor U6494 (N_6494,N_4051,N_2571);
nand U6495 (N_6495,N_3031,N_2348);
and U6496 (N_6496,N_4642,N_1855);
nand U6497 (N_6497,N_1117,N_3169);
nand U6498 (N_6498,N_1314,N_4157);
and U6499 (N_6499,N_903,N_4894);
nand U6500 (N_6500,N_4871,N_2037);
nand U6501 (N_6501,N_1842,N_1764);
nand U6502 (N_6502,N_2110,N_3208);
nor U6503 (N_6503,N_4978,N_2252);
nand U6504 (N_6504,N_4634,N_3093);
nor U6505 (N_6505,N_3940,N_4619);
or U6506 (N_6506,N_1893,N_2374);
nand U6507 (N_6507,N_3734,N_4413);
nand U6508 (N_6508,N_3620,N_1849);
or U6509 (N_6509,N_2667,N_1280);
or U6510 (N_6510,N_4743,N_1009);
xnor U6511 (N_6511,N_3969,N_1045);
nor U6512 (N_6512,N_72,N_28);
nor U6513 (N_6513,N_1641,N_4601);
and U6514 (N_6514,N_2042,N_4663);
nand U6515 (N_6515,N_3709,N_772);
and U6516 (N_6516,N_166,N_1270);
nand U6517 (N_6517,N_24,N_943);
and U6518 (N_6518,N_4574,N_4387);
nor U6519 (N_6519,N_2101,N_1066);
nand U6520 (N_6520,N_4972,N_4826);
xor U6521 (N_6521,N_3222,N_2618);
or U6522 (N_6522,N_2624,N_790);
xor U6523 (N_6523,N_897,N_3504);
or U6524 (N_6524,N_1931,N_936);
or U6525 (N_6525,N_2679,N_895);
nand U6526 (N_6526,N_2780,N_4924);
xnor U6527 (N_6527,N_3522,N_2393);
or U6528 (N_6528,N_4589,N_1326);
or U6529 (N_6529,N_3127,N_908);
nand U6530 (N_6530,N_4031,N_2032);
xnor U6531 (N_6531,N_3797,N_3281);
xnor U6532 (N_6532,N_2833,N_2437);
nand U6533 (N_6533,N_546,N_3033);
and U6534 (N_6534,N_3020,N_2174);
nand U6535 (N_6535,N_3762,N_842);
nand U6536 (N_6536,N_2514,N_628);
and U6537 (N_6537,N_3652,N_4219);
or U6538 (N_6538,N_3314,N_4987);
nand U6539 (N_6539,N_3358,N_2808);
and U6540 (N_6540,N_259,N_1225);
nor U6541 (N_6541,N_3585,N_2884);
or U6542 (N_6542,N_3104,N_2875);
and U6543 (N_6543,N_702,N_1591);
nand U6544 (N_6544,N_4958,N_4111);
nor U6545 (N_6545,N_1382,N_4693);
nor U6546 (N_6546,N_2643,N_3191);
or U6547 (N_6547,N_516,N_2066);
or U6548 (N_6548,N_1418,N_1887);
nand U6549 (N_6549,N_1811,N_2703);
xor U6550 (N_6550,N_4907,N_2809);
nand U6551 (N_6551,N_627,N_236);
and U6552 (N_6552,N_1464,N_4504);
and U6553 (N_6553,N_2210,N_347);
or U6554 (N_6554,N_996,N_725);
nand U6555 (N_6555,N_522,N_4204);
or U6556 (N_6556,N_2620,N_4973);
or U6557 (N_6557,N_3825,N_2915);
nand U6558 (N_6558,N_583,N_2399);
or U6559 (N_6559,N_2866,N_4552);
nand U6560 (N_6560,N_3791,N_685);
nand U6561 (N_6561,N_3941,N_2762);
nand U6562 (N_6562,N_2478,N_3321);
or U6563 (N_6563,N_435,N_1260);
nand U6564 (N_6564,N_4453,N_3717);
or U6565 (N_6565,N_2513,N_1016);
nand U6566 (N_6566,N_1784,N_665);
or U6567 (N_6567,N_1606,N_4583);
and U6568 (N_6568,N_3290,N_4679);
xnor U6569 (N_6569,N_307,N_1261);
or U6570 (N_6570,N_4631,N_1668);
and U6571 (N_6571,N_2122,N_2746);
or U6572 (N_6572,N_773,N_778);
nand U6573 (N_6573,N_380,N_1789);
xnor U6574 (N_6574,N_3891,N_184);
and U6575 (N_6575,N_960,N_3157);
and U6576 (N_6576,N_1108,N_2880);
and U6577 (N_6577,N_3902,N_3466);
and U6578 (N_6578,N_1073,N_3185);
xor U6579 (N_6579,N_2536,N_2860);
nand U6580 (N_6580,N_1401,N_2855);
or U6581 (N_6581,N_99,N_4548);
and U6582 (N_6582,N_6,N_165);
xor U6583 (N_6583,N_1405,N_4289);
and U6584 (N_6584,N_3277,N_1865);
nor U6585 (N_6585,N_830,N_4078);
nand U6586 (N_6586,N_1662,N_2353);
and U6587 (N_6587,N_4442,N_1331);
and U6588 (N_6588,N_3370,N_2973);
nor U6589 (N_6589,N_4369,N_4058);
or U6590 (N_6590,N_951,N_989);
or U6591 (N_6591,N_1620,N_23);
and U6592 (N_6592,N_4120,N_2545);
and U6593 (N_6593,N_1526,N_792);
nor U6594 (N_6594,N_460,N_1860);
and U6595 (N_6595,N_4788,N_1736);
nand U6596 (N_6596,N_2455,N_2201);
and U6597 (N_6597,N_444,N_1647);
and U6598 (N_6598,N_3925,N_1939);
or U6599 (N_6599,N_1669,N_3708);
and U6600 (N_6600,N_1688,N_1983);
nand U6601 (N_6601,N_1484,N_1143);
and U6602 (N_6602,N_4298,N_2728);
nor U6603 (N_6603,N_2015,N_838);
nor U6604 (N_6604,N_2377,N_4811);
nor U6605 (N_6605,N_4494,N_3375);
nor U6606 (N_6606,N_1739,N_1584);
nand U6607 (N_6607,N_1200,N_4231);
and U6608 (N_6608,N_1229,N_3403);
nand U6609 (N_6609,N_4100,N_1679);
nor U6610 (N_6610,N_132,N_2862);
nor U6611 (N_6611,N_1141,N_4629);
nor U6612 (N_6612,N_4579,N_4934);
nor U6613 (N_6613,N_3414,N_2895);
and U6614 (N_6614,N_381,N_1138);
nor U6615 (N_6615,N_3066,N_160);
nor U6616 (N_6616,N_92,N_765);
and U6617 (N_6617,N_491,N_827);
nand U6618 (N_6618,N_3896,N_651);
and U6619 (N_6619,N_3548,N_3707);
and U6620 (N_6620,N_1743,N_1881);
or U6621 (N_6621,N_1822,N_467);
and U6622 (N_6622,N_796,N_1592);
and U6623 (N_6623,N_136,N_755);
and U6624 (N_6624,N_4487,N_3131);
nand U6625 (N_6625,N_4614,N_1097);
or U6626 (N_6626,N_711,N_2454);
nand U6627 (N_6627,N_2088,N_4683);
nand U6628 (N_6628,N_4140,N_4927);
and U6629 (N_6629,N_172,N_614);
nand U6630 (N_6630,N_1277,N_4143);
nand U6631 (N_6631,N_4457,N_4566);
and U6632 (N_6632,N_2800,N_3010);
or U6633 (N_6633,N_4807,N_4604);
nor U6634 (N_6634,N_3472,N_2070);
and U6635 (N_6635,N_2089,N_2360);
or U6636 (N_6636,N_2365,N_2759);
and U6637 (N_6637,N_2795,N_3980);
or U6638 (N_6638,N_596,N_3484);
nor U6639 (N_6639,N_4046,N_2400);
and U6640 (N_6640,N_1170,N_4952);
nand U6641 (N_6641,N_4577,N_2234);
or U6642 (N_6642,N_4007,N_3529);
xor U6643 (N_6643,N_1362,N_2498);
nand U6644 (N_6644,N_3768,N_4071);
and U6645 (N_6645,N_137,N_1485);
or U6646 (N_6646,N_2232,N_4533);
or U6647 (N_6647,N_2240,N_3009);
xnor U6648 (N_6648,N_950,N_3890);
or U6649 (N_6649,N_4066,N_2578);
nor U6650 (N_6650,N_3900,N_4201);
nor U6651 (N_6651,N_4014,N_1568);
nand U6652 (N_6652,N_2738,N_2684);
nand U6653 (N_6653,N_154,N_1613);
xnor U6654 (N_6654,N_1303,N_3987);
nand U6655 (N_6655,N_848,N_800);
nor U6656 (N_6656,N_4156,N_1047);
or U6657 (N_6657,N_1474,N_2287);
and U6658 (N_6658,N_4797,N_3255);
xor U6659 (N_6659,N_768,N_3476);
and U6660 (N_6660,N_2907,N_4767);
nor U6661 (N_6661,N_200,N_4518);
and U6662 (N_6662,N_3245,N_2405);
nor U6663 (N_6663,N_2623,N_1365);
nor U6664 (N_6664,N_88,N_1201);
nand U6665 (N_6665,N_2486,N_2996);
nor U6666 (N_6666,N_51,N_3984);
nor U6667 (N_6667,N_4801,N_925);
nor U6668 (N_6668,N_4332,N_1570);
or U6669 (N_6669,N_4061,N_2890);
xor U6670 (N_6670,N_4483,N_3389);
nand U6671 (N_6671,N_1061,N_71);
or U6672 (N_6672,N_2835,N_4443);
xor U6673 (N_6673,N_490,N_2324);
nand U6674 (N_6674,N_1639,N_3703);
and U6675 (N_6675,N_358,N_3345);
nor U6676 (N_6676,N_2446,N_4448);
nand U6677 (N_6677,N_400,N_2113);
and U6678 (N_6678,N_1098,N_1726);
nor U6679 (N_6679,N_968,N_1259);
or U6680 (N_6680,N_3236,N_4821);
xnor U6681 (N_6681,N_4546,N_469);
or U6682 (N_6682,N_1233,N_3397);
nor U6683 (N_6683,N_183,N_1398);
and U6684 (N_6684,N_4762,N_2540);
nand U6685 (N_6685,N_1019,N_4598);
or U6686 (N_6686,N_4447,N_257);
and U6687 (N_6687,N_1273,N_671);
or U6688 (N_6688,N_4510,N_4091);
or U6689 (N_6689,N_2008,N_4254);
nand U6690 (N_6690,N_216,N_4025);
xor U6691 (N_6691,N_4233,N_2265);
nand U6692 (N_6692,N_747,N_514);
xnor U6693 (N_6693,N_4759,N_4278);
nor U6694 (N_6694,N_2948,N_2420);
and U6695 (N_6695,N_1240,N_238);
nor U6696 (N_6696,N_1391,N_2080);
and U6697 (N_6697,N_4237,N_3108);
nand U6698 (N_6698,N_4083,N_4886);
and U6699 (N_6699,N_4180,N_1032);
or U6700 (N_6700,N_4484,N_1638);
and U6701 (N_6701,N_4105,N_2235);
nor U6702 (N_6702,N_4003,N_3488);
or U6703 (N_6703,N_4884,N_4791);
and U6704 (N_6704,N_4691,N_1182);
and U6705 (N_6705,N_3766,N_1176);
xor U6706 (N_6706,N_746,N_3905);
and U6707 (N_6707,N_4450,N_4425);
nor U6708 (N_6708,N_3220,N_2067);
nor U6709 (N_6709,N_294,N_1783);
nor U6710 (N_6710,N_1283,N_2164);
and U6711 (N_6711,N_4465,N_3711);
nor U6712 (N_6712,N_3594,N_3004);
and U6713 (N_6713,N_1250,N_4467);
and U6714 (N_6714,N_1222,N_3243);
and U6715 (N_6715,N_4469,N_3461);
nand U6716 (N_6716,N_3959,N_1998);
and U6717 (N_6717,N_2555,N_649);
or U6718 (N_6718,N_3760,N_3492);
nand U6719 (N_6719,N_2534,N_3376);
and U6720 (N_6720,N_4845,N_104);
nor U6721 (N_6721,N_2843,N_4724);
nor U6722 (N_6722,N_2539,N_1989);
or U6723 (N_6723,N_4865,N_4354);
nand U6724 (N_6724,N_1776,N_3750);
nand U6725 (N_6725,N_1761,N_4789);
nor U6726 (N_6726,N_4999,N_108);
or U6727 (N_6727,N_3558,N_2496);
nor U6728 (N_6728,N_2695,N_382);
xor U6729 (N_6729,N_3147,N_4161);
and U6730 (N_6730,N_2939,N_1439);
xnor U6731 (N_6731,N_1964,N_3815);
and U6732 (N_6732,N_4449,N_4306);
nand U6733 (N_6733,N_3882,N_3023);
nand U6734 (N_6734,N_4089,N_4176);
nor U6735 (N_6735,N_2412,N_1359);
nand U6736 (N_6736,N_3765,N_3388);
nor U6737 (N_6737,N_2031,N_135);
nor U6738 (N_6738,N_3817,N_3674);
or U6739 (N_6739,N_197,N_324);
nand U6740 (N_6740,N_1997,N_4316);
and U6741 (N_6741,N_4498,N_4206);
and U6742 (N_6742,N_3720,N_1970);
or U6743 (N_6743,N_1454,N_4850);
xor U6744 (N_6744,N_3830,N_2177);
nand U6745 (N_6745,N_4881,N_707);
nor U6746 (N_6746,N_3894,N_181);
nor U6747 (N_6747,N_4551,N_1969);
or U6748 (N_6748,N_1904,N_3537);
nand U6749 (N_6749,N_2500,N_2821);
or U6750 (N_6750,N_3557,N_2974);
nor U6751 (N_6751,N_3634,N_3546);
xor U6752 (N_6752,N_1115,N_63);
or U6753 (N_6753,N_1469,N_4802);
and U6754 (N_6754,N_972,N_2980);
and U6755 (N_6755,N_3541,N_3172);
xor U6756 (N_6756,N_2313,N_2730);
nor U6757 (N_6757,N_2495,N_4783);
and U6758 (N_6758,N_376,N_1411);
and U6759 (N_6759,N_4192,N_1926);
nor U6760 (N_6760,N_2065,N_1421);
xor U6761 (N_6761,N_1923,N_3184);
nand U6762 (N_6762,N_1364,N_1099);
or U6763 (N_6763,N_3430,N_4129);
or U6764 (N_6764,N_2953,N_2036);
nand U6765 (N_6765,N_2249,N_1712);
nor U6766 (N_6766,N_2372,N_1957);
and U6767 (N_6767,N_1022,N_1043);
or U6768 (N_6768,N_4701,N_3495);
xnor U6769 (N_6769,N_880,N_1456);
nand U6770 (N_6770,N_3244,N_888);
or U6771 (N_6771,N_1910,N_2754);
xnor U6772 (N_6772,N_896,N_563);
xor U6773 (N_6773,N_361,N_2844);
nor U6774 (N_6774,N_4190,N_922);
nor U6775 (N_6775,N_788,N_3907);
nand U6776 (N_6776,N_1933,N_2870);
and U6777 (N_6777,N_986,N_4674);
or U6778 (N_6778,N_2427,N_4422);
nand U6779 (N_6779,N_3531,N_2274);
nand U6780 (N_6780,N_1384,N_3886);
or U6781 (N_6781,N_2079,N_1622);
nand U6782 (N_6782,N_3333,N_3428);
nand U6783 (N_6783,N_2266,N_3667);
nand U6784 (N_6784,N_590,N_991);
nand U6785 (N_6785,N_1834,N_3372);
and U6786 (N_6786,N_1511,N_4439);
or U6787 (N_6787,N_2802,N_4481);
and U6788 (N_6788,N_987,N_4645);
nand U6789 (N_6789,N_1136,N_2594);
or U6790 (N_6790,N_4244,N_2664);
and U6791 (N_6791,N_1757,N_3927);
or U6792 (N_6792,N_1296,N_3656);
or U6793 (N_6793,N_1050,N_3924);
nor U6794 (N_6794,N_2022,N_3658);
nor U6795 (N_6795,N_1267,N_2771);
or U6796 (N_6796,N_3610,N_4613);
and U6797 (N_6797,N_457,N_2621);
nor U6798 (N_6798,N_3512,N_4939);
nand U6799 (N_6799,N_1917,N_4835);
and U6800 (N_6800,N_390,N_2262);
or U6801 (N_6801,N_3831,N_2931);
nand U6802 (N_6802,N_1623,N_219);
nor U6803 (N_6803,N_459,N_3335);
xor U6804 (N_6804,N_2482,N_2222);
nor U6805 (N_6805,N_4230,N_3318);
nor U6806 (N_6806,N_1545,N_397);
nor U6807 (N_6807,N_3813,N_3464);
nor U6808 (N_6808,N_1667,N_3471);
and U6809 (N_6809,N_1705,N_2304);
nand U6810 (N_6810,N_4350,N_3121);
xor U6811 (N_6811,N_1323,N_2649);
or U6812 (N_6812,N_480,N_738);
nand U6813 (N_6813,N_2475,N_149);
or U6814 (N_6814,N_2020,N_3252);
or U6815 (N_6815,N_726,N_3046);
nor U6816 (N_6816,N_2729,N_1076);
nand U6817 (N_6817,N_4969,N_1429);
nand U6818 (N_6818,N_4257,N_1377);
and U6819 (N_6819,N_1486,N_3981);
nor U6820 (N_6820,N_4824,N_276);
and U6821 (N_6821,N_3957,N_2300);
and U6822 (N_6822,N_3306,N_4097);
or U6823 (N_6823,N_515,N_4926);
nor U6824 (N_6824,N_2007,N_3297);
nand U6825 (N_6825,N_4022,N_1950);
nor U6826 (N_6826,N_534,N_2160);
xnor U6827 (N_6827,N_245,N_4321);
or U6828 (N_6828,N_2490,N_3006);
and U6829 (N_6829,N_2397,N_3133);
nor U6830 (N_6830,N_173,N_321);
or U6831 (N_6831,N_2484,N_1514);
nand U6832 (N_6832,N_2688,N_2927);
and U6833 (N_6833,N_1013,N_1869);
nand U6834 (N_6834,N_1703,N_2168);
nor U6835 (N_6835,N_2052,N_4456);
or U6836 (N_6836,N_528,N_1803);
or U6837 (N_6837,N_1826,N_123);
xor U6838 (N_6838,N_2061,N_4378);
or U6839 (N_6839,N_205,N_2179);
or U6840 (N_6840,N_1630,N_338);
nand U6841 (N_6841,N_3784,N_1595);
xnor U6842 (N_6842,N_4772,N_4765);
nand U6843 (N_6843,N_958,N_359);
nor U6844 (N_6844,N_504,N_3644);
and U6845 (N_6845,N_2924,N_2901);
xor U6846 (N_6846,N_2991,N_2642);
nand U6847 (N_6847,N_2910,N_4611);
and U6848 (N_6848,N_2167,N_2648);
nand U6849 (N_6849,N_1060,N_1390);
nor U6850 (N_6850,N_2893,N_2633);
nor U6851 (N_6851,N_2476,N_2711);
nor U6852 (N_6852,N_9,N_1231);
nor U6853 (N_6853,N_1938,N_1872);
xnor U6854 (N_6854,N_3555,N_2918);
nor U6855 (N_6855,N_3575,N_3289);
nor U6856 (N_6856,N_1806,N_2963);
xnor U6857 (N_6857,N_3394,N_417);
xnor U6858 (N_6858,N_1691,N_3855);
nor U6859 (N_6859,N_2483,N_4049);
xor U6860 (N_6860,N_1332,N_2671);
or U6861 (N_6861,N_1335,N_3212);
nand U6862 (N_6862,N_3477,N_1127);
or U6863 (N_6863,N_2315,N_2570);
nor U6864 (N_6864,N_4351,N_68);
and U6865 (N_6865,N_142,N_4212);
nor U6866 (N_6866,N_4756,N_2176);
and U6867 (N_6867,N_4407,N_1355);
nand U6868 (N_6868,N_3129,N_2497);
nor U6869 (N_6869,N_2604,N_1814);
nand U6870 (N_6870,N_2460,N_1297);
and U6871 (N_6871,N_1083,N_971);
nand U6872 (N_6872,N_133,N_2798);
nand U6873 (N_6873,N_949,N_3029);
nand U6874 (N_6874,N_3729,N_4963);
or U6875 (N_6875,N_662,N_145);
or U6876 (N_6876,N_76,N_1187);
xor U6877 (N_6877,N_2064,N_1339);
or U6878 (N_6878,N_852,N_240);
xor U6879 (N_6879,N_3811,N_2188);
nor U6880 (N_6880,N_2678,N_3276);
or U6881 (N_6881,N_1397,N_319);
and U6882 (N_6882,N_4159,N_4796);
or U6883 (N_6883,N_2777,N_1328);
or U6884 (N_6884,N_1262,N_4423);
xor U6885 (N_6885,N_688,N_4652);
xor U6886 (N_6886,N_4085,N_2923);
xnor U6887 (N_6887,N_1742,N_2981);
or U6888 (N_6888,N_3520,N_3802);
nor U6889 (N_6889,N_4116,N_1086);
nor U6890 (N_6890,N_1320,N_4102);
nor U6891 (N_6891,N_3823,N_920);
and U6892 (N_6892,N_3758,N_2335);
xor U6893 (N_6893,N_3785,N_4141);
nand U6894 (N_6894,N_105,N_3827);
nor U6895 (N_6895,N_4508,N_2677);
or U6896 (N_6896,N_541,N_281);
and U6897 (N_6897,N_3604,N_4815);
or U6898 (N_6898,N_3207,N_61);
and U6899 (N_6899,N_3846,N_3747);
or U6900 (N_6900,N_3640,N_585);
nand U6901 (N_6901,N_3623,N_2888);
and U6902 (N_6902,N_4925,N_4545);
or U6903 (N_6903,N_1116,N_3617);
xor U6904 (N_6904,N_1713,N_4831);
nor U6905 (N_6905,N_4037,N_527);
nand U6906 (N_6906,N_4670,N_750);
and U6907 (N_6907,N_3562,N_4793);
nor U6908 (N_6908,N_3675,N_2363);
or U6909 (N_6909,N_3730,N_3215);
and U6910 (N_6910,N_1543,N_468);
or U6911 (N_6911,N_2805,N_1275);
and U6912 (N_6912,N_3563,N_3552);
or U6913 (N_6913,N_196,N_1155);
xnor U6914 (N_6914,N_3892,N_2355);
or U6915 (N_6915,N_3832,N_3801);
and U6916 (N_6916,N_2161,N_1539);
xor U6917 (N_6917,N_3857,N_3946);
and U6918 (N_6918,N_3468,N_4384);
or U6919 (N_6919,N_3268,N_4955);
and U6920 (N_6920,N_2585,N_121);
nor U6921 (N_6921,N_4137,N_3176);
or U6922 (N_6922,N_192,N_759);
and U6923 (N_6923,N_2028,N_2197);
nand U6924 (N_6924,N_4933,N_2380);
nor U6925 (N_6925,N_300,N_4686);
nand U6926 (N_6926,N_1762,N_2276);
nor U6927 (N_6927,N_3099,N_2687);
and U6928 (N_6928,N_1159,N_3142);
xnor U6929 (N_6929,N_4492,N_4996);
or U6930 (N_6930,N_365,N_4224);
and U6931 (N_6931,N_1459,N_4359);
nand U6932 (N_6932,N_3865,N_959);
nor U6933 (N_6933,N_4324,N_737);
and U6934 (N_6934,N_2985,N_2913);
and U6935 (N_6935,N_4739,N_1463);
xnor U6936 (N_6936,N_4622,N_3181);
nand U6937 (N_6937,N_2011,N_4676);
and U6938 (N_6938,N_1433,N_3561);
and U6939 (N_6939,N_3317,N_2597);
or U6940 (N_6940,N_4569,N_3536);
nor U6941 (N_6941,N_3975,N_4082);
nand U6942 (N_6942,N_3351,N_4935);
or U6943 (N_6943,N_2280,N_4684);
nor U6944 (N_6944,N_1722,N_1825);
nor U6945 (N_6945,N_1535,N_1854);
or U6946 (N_6946,N_2242,N_2124);
and U6947 (N_6947,N_3666,N_499);
nand U6948 (N_6948,N_2625,N_4901);
xor U6949 (N_6949,N_4075,N_2012);
xnor U6950 (N_6950,N_1052,N_195);
xnor U6951 (N_6951,N_603,N_2057);
nand U6952 (N_6952,N_2185,N_326);
nand U6953 (N_6953,N_3396,N_1870);
nor U6954 (N_6954,N_3639,N_2254);
nor U6955 (N_6955,N_1414,N_4661);
and U6956 (N_6956,N_1352,N_2106);
and U6957 (N_6957,N_3847,N_3856);
or U6958 (N_6958,N_3043,N_814);
nand U6959 (N_6959,N_4779,N_2737);
xor U6960 (N_6960,N_3544,N_213);
or U6961 (N_6961,N_90,N_2431);
or U6962 (N_6962,N_4919,N_4534);
or U6963 (N_6963,N_4904,N_4401);
xnor U6964 (N_6964,N_2334,N_2993);
nor U6965 (N_6965,N_955,N_3398);
or U6966 (N_6966,N_3649,N_3141);
nand U6967 (N_6967,N_3238,N_557);
and U6968 (N_6968,N_2914,N_4562);
xnor U6969 (N_6969,N_4568,N_449);
and U6970 (N_6970,N_786,N_3462);
and U6971 (N_6971,N_3391,N_2140);
and U6972 (N_6972,N_293,N_3657);
nand U6973 (N_6973,N_3241,N_2760);
and U6974 (N_6974,N_4902,N_2622);
and U6975 (N_6975,N_3308,N_584);
or U6976 (N_6976,N_2023,N_4625);
xor U6977 (N_6977,N_126,N_666);
xnor U6978 (N_6978,N_1862,N_455);
and U6979 (N_6979,N_3989,N_32);
and U6980 (N_6980,N_1833,N_4986);
and U6981 (N_6981,N_3576,N_1334);
nand U6982 (N_6982,N_3503,N_458);
nor U6983 (N_6983,N_377,N_2472);
xor U6984 (N_6984,N_3479,N_1646);
nor U6985 (N_6985,N_4153,N_1799);
and U6986 (N_6986,N_2832,N_1325);
or U6987 (N_6987,N_3686,N_1815);
nand U6988 (N_6988,N_592,N_2840);
and U6989 (N_6989,N_2598,N_18);
or U6990 (N_6990,N_3431,N_1286);
nand U6991 (N_6991,N_1040,N_3165);
and U6992 (N_6992,N_687,N_345);
or U6993 (N_6993,N_4997,N_2871);
and U6994 (N_6994,N_4950,N_3300);
and U6995 (N_6995,N_3805,N_4368);
nor U6996 (N_6996,N_2952,N_3307);
and U6997 (N_6997,N_4110,N_466);
and U6998 (N_6998,N_610,N_4080);
xor U6999 (N_6999,N_1975,N_1643);
and U7000 (N_7000,N_1255,N_2297);
nor U7001 (N_7001,N_4430,N_4819);
and U7002 (N_7002,N_2435,N_1996);
nand U7003 (N_7003,N_1732,N_3294);
or U7004 (N_7004,N_4002,N_2271);
or U7005 (N_7005,N_1473,N_3740);
or U7006 (N_7006,N_2150,N_3086);
and U7007 (N_7007,N_2458,N_2885);
or U7008 (N_7008,N_4334,N_1979);
nor U7009 (N_7009,N_757,N_3067);
or U7010 (N_7010,N_523,N_2682);
and U7011 (N_7011,N_1423,N_4493);
nor U7012 (N_7012,N_3167,N_4402);
or U7013 (N_7013,N_3773,N_664);
nor U7014 (N_7014,N_4238,N_4880);
and U7015 (N_7015,N_2246,N_2474);
or U7016 (N_7016,N_2919,N_331);
or U7017 (N_7017,N_1413,N_3284);
nand U7018 (N_7018,N_2565,N_1827);
nand U7019 (N_7019,N_93,N_2390);
nor U7020 (N_7020,N_2769,N_2861);
nand U7021 (N_7021,N_2260,N_2429);
nor U7022 (N_7022,N_3064,N_1995);
nand U7023 (N_7023,N_3899,N_3962);
nand U7024 (N_7024,N_3731,N_7);
xor U7025 (N_7025,N_3328,N_1949);
or U7026 (N_7026,N_1534,N_4207);
and U7027 (N_7027,N_4194,N_2505);
and U7028 (N_7028,N_4786,N_3992);
xor U7029 (N_7029,N_4600,N_2314);
nor U7030 (N_7030,N_103,N_1577);
and U7031 (N_7031,N_310,N_4630);
and U7032 (N_7032,N_407,N_720);
nand U7033 (N_7033,N_3780,N_2135);
nand U7034 (N_7034,N_819,N_1218);
or U7035 (N_7035,N_2858,N_4414);
nor U7036 (N_7036,N_1399,N_1449);
nor U7037 (N_7037,N_1069,N_346);
xnor U7038 (N_7038,N_452,N_4164);
and U7039 (N_7039,N_422,N_4179);
or U7040 (N_7040,N_4828,N_4747);
xor U7041 (N_7041,N_1053,N_4544);
or U7042 (N_7042,N_503,N_2994);
nor U7043 (N_7043,N_4985,N_1838);
and U7044 (N_7044,N_4785,N_3120);
and U7045 (N_7045,N_4994,N_500);
nand U7046 (N_7046,N_836,N_927);
and U7047 (N_7047,N_2504,N_4713);
nand U7048 (N_7048,N_387,N_4170);
nand U7049 (N_7049,N_676,N_186);
or U7050 (N_7050,N_3168,N_413);
or U7051 (N_7051,N_4004,N_3203);
nand U7052 (N_7052,N_3696,N_1318);
xor U7053 (N_7053,N_3360,N_4863);
nor U7054 (N_7054,N_1954,N_2572);
nor U7055 (N_7055,N_4936,N_2934);
nor U7056 (N_7056,N_1637,N_846);
or U7057 (N_7057,N_3673,N_801);
nand U7058 (N_7058,N_1216,N_4647);
nand U7059 (N_7059,N_379,N_2541);
nand U7060 (N_7060,N_857,N_1205);
and U7061 (N_7061,N_1837,N_1417);
or U7062 (N_7062,N_2815,N_266);
nor U7063 (N_7063,N_31,N_899);
nor U7064 (N_7064,N_1941,N_1617);
or U7065 (N_7065,N_2344,N_1386);
xnor U7066 (N_7066,N_2244,N_519);
xor U7067 (N_7067,N_308,N_3036);
nor U7068 (N_7068,N_3744,N_3970);
or U7069 (N_7069,N_1487,N_645);
and U7070 (N_7070,N_3974,N_2567);
nand U7071 (N_7071,N_1891,N_2511);
or U7072 (N_7072,N_1056,N_2723);
nand U7073 (N_7073,N_2921,N_3879);
nand U7074 (N_7074,N_1994,N_1062);
nand U7075 (N_7075,N_2245,N_696);
and U7076 (N_7076,N_3777,N_448);
nor U7077 (N_7077,N_2480,N_3933);
nand U7078 (N_7078,N_659,N_3547);
or U7079 (N_7079,N_2316,N_52);
or U7080 (N_7080,N_1363,N_1873);
and U7081 (N_7081,N_4104,N_4225);
and U7082 (N_7082,N_4108,N_677);
and U7083 (N_7083,N_3614,N_875);
or U7084 (N_7084,N_1169,N_4016);
nand U7085 (N_7085,N_1024,N_1354);
nor U7086 (N_7086,N_1673,N_923);
xor U7087 (N_7087,N_3527,N_2373);
nand U7088 (N_7088,N_4065,N_3432);
nand U7089 (N_7089,N_4059,N_3106);
and U7090 (N_7090,N_4832,N_3195);
or U7091 (N_7091,N_705,N_4032);
nand U7092 (N_7092,N_2697,N_4951);
and U7093 (N_7093,N_4349,N_4671);
nor U7094 (N_7094,N_4616,N_3156);
and U7095 (N_7095,N_2583,N_4329);
or U7096 (N_7096,N_222,N_3202);
nor U7097 (N_7097,N_4873,N_3041);
nand U7098 (N_7098,N_1346,N_3733);
nand U7099 (N_7099,N_4712,N_3534);
and U7100 (N_7100,N_3416,N_3850);
nor U7101 (N_7101,N_3434,N_2867);
xor U7102 (N_7102,N_2002,N_1305);
xor U7103 (N_7103,N_3693,N_4132);
nor U7104 (N_7104,N_263,N_2175);
and U7105 (N_7105,N_1462,N_2674);
or U7106 (N_7106,N_4019,N_752);
xnor U7107 (N_7107,N_4949,N_1552);
or U7108 (N_7108,N_3588,N_2006);
xor U7109 (N_7109,N_2375,N_642);
and U7110 (N_7110,N_4731,N_2401);
nor U7111 (N_7111,N_1447,N_1819);
nand U7112 (N_7112,N_3549,N_2158);
or U7113 (N_7113,N_2892,N_4758);
nor U7114 (N_7114,N_2987,N_202);
nor U7115 (N_7115,N_4060,N_2059);
or U7116 (N_7116,N_2632,N_2139);
or U7117 (N_7117,N_969,N_1008);
nor U7118 (N_7118,N_4549,N_1817);
or U7119 (N_7119,N_1085,N_1763);
nand U7120 (N_7120,N_2368,N_4405);
nor U7121 (N_7121,N_2418,N_3839);
nor U7122 (N_7122,N_2024,N_2501);
xnor U7123 (N_7123,N_3187,N_2039);
xor U7124 (N_7124,N_1583,N_1716);
or U7125 (N_7125,N_2121,N_2587);
and U7126 (N_7126,N_4578,N_4399);
and U7127 (N_7127,N_1482,N_86);
xor U7128 (N_7128,N_1537,N_4076);
or U7129 (N_7129,N_4455,N_3193);
and U7130 (N_7130,N_3605,N_3016);
nor U7131 (N_7131,N_3569,N_2362);
nand U7132 (N_7132,N_17,N_4781);
xnor U7133 (N_7133,N_4338,N_2292);
nor U7134 (N_7134,N_4178,N_783);
nor U7135 (N_7135,N_3153,N_4812);
nand U7136 (N_7136,N_1737,N_4898);
or U7137 (N_7137,N_3330,N_1316);
or U7138 (N_7138,N_4567,N_4906);
and U7139 (N_7139,N_1960,N_3014);
and U7140 (N_7140,N_2701,N_1528);
nand U7141 (N_7141,N_1959,N_1131);
and U7142 (N_7142,N_2527,N_2912);
and U7143 (N_7143,N_15,N_4858);
nand U7144 (N_7144,N_1338,N_2239);
and U7145 (N_7145,N_305,N_3170);
nor U7146 (N_7146,N_384,N_3337);
or U7147 (N_7147,N_1695,N_565);
nand U7148 (N_7148,N_3171,N_681);
or U7149 (N_7149,N_4953,N_1094);
and U7150 (N_7150,N_2756,N_2463);
or U7151 (N_7151,N_3114,N_2043);
or U7152 (N_7152,N_821,N_4597);
nand U7153 (N_7153,N_2248,N_3095);
xnor U7154 (N_7154,N_4874,N_3473);
nor U7155 (N_7155,N_965,N_1490);
nand U7156 (N_7156,N_3852,N_839);
nor U7157 (N_7157,N_1206,N_96);
nor U7158 (N_7158,N_4348,N_306);
and U7159 (N_7159,N_4699,N_2852);
nor U7160 (N_7160,N_2105,N_2432);
and U7161 (N_7161,N_822,N_2263);
nor U7162 (N_7162,N_355,N_3332);
nor U7163 (N_7163,N_587,N_657);
or U7164 (N_7164,N_4496,N_4462);
xor U7165 (N_7165,N_498,N_3076);
nand U7166 (N_7166,N_3826,N_1081);
nand U7167 (N_7167,N_102,N_3455);
and U7168 (N_7168,N_4131,N_3635);
or U7169 (N_7169,N_4294,N_4657);
nor U7170 (N_7170,N_1521,N_4560);
and U7171 (N_7171,N_4576,N_3408);
and U7172 (N_7172,N_1589,N_4941);
and U7173 (N_7173,N_4366,N_3075);
and U7174 (N_7174,N_1859,N_4766);
nor U7175 (N_7175,N_3261,N_1569);
xor U7176 (N_7176,N_2557,N_1845);
nor U7177 (N_7177,N_1133,N_3402);
nor U7178 (N_7178,N_91,N_4416);
nand U7179 (N_7179,N_2731,N_1650);
nor U7180 (N_7180,N_762,N_629);
or U7181 (N_7181,N_639,N_660);
and U7182 (N_7182,N_3716,N_2216);
and U7183 (N_7183,N_2503,N_3713);
nand U7184 (N_7184,N_2169,N_4034);
or U7185 (N_7185,N_1160,N_551);
nand U7186 (N_7186,N_2868,N_3834);
xnor U7187 (N_7187,N_394,N_2689);
nand U7188 (N_7188,N_4335,N_1300);
nand U7189 (N_7189,N_4175,N_2445);
nor U7190 (N_7190,N_2507,N_1775);
or U7191 (N_7191,N_3510,N_1130);
xnor U7192 (N_7192,N_722,N_3056);
nor U7193 (N_7193,N_2937,N_4709);
or U7194 (N_7194,N_882,N_1289);
and U7195 (N_7195,N_1102,N_4753);
nor U7196 (N_7196,N_2775,N_399);
or U7197 (N_7197,N_593,N_4418);
nand U7198 (N_7198,N_3441,N_4424);
or U7199 (N_7199,N_568,N_4816);
nand U7200 (N_7200,N_1927,N_525);
and U7201 (N_7201,N_4308,N_4782);
nor U7202 (N_7202,N_163,N_3863);
nand U7203 (N_7203,N_4982,N_817);
nand U7204 (N_7204,N_4310,N_2864);
and U7205 (N_7205,N_624,N_808);
nor U7206 (N_7206,N_4134,N_3819);
and U7207 (N_7207,N_1897,N_1524);
nor U7208 (N_7208,N_2389,N_1607);
nor U7209 (N_7209,N_3849,N_2593);
nor U7210 (N_7210,N_3551,N_13);
nor U7211 (N_7211,N_2403,N_2423);
or U7212 (N_7212,N_130,N_3251);
nand U7213 (N_7213,N_1173,N_2553);
nor U7214 (N_7214,N_2577,N_2863);
or U7215 (N_7215,N_3680,N_4706);
nand U7216 (N_7216,N_3966,N_4361);
nand U7217 (N_7217,N_3670,N_1614);
nand U7218 (N_7218,N_4166,N_3737);
or U7219 (N_7219,N_1093,N_226);
nor U7220 (N_7220,N_2590,N_290);
nand U7221 (N_7221,N_3516,N_2469);
nor U7222 (N_7222,N_4774,N_1165);
nand U7223 (N_7223,N_3745,N_3727);
nor U7224 (N_7224,N_2961,N_1733);
and U7225 (N_7225,N_550,N_4872);
nor U7226 (N_7226,N_1578,N_714);
and U7227 (N_7227,N_185,N_2920);
nand U7228 (N_7228,N_2104,N_4309);
or U7229 (N_7229,N_4909,N_2404);
or U7230 (N_7230,N_3624,N_4266);
nand U7231 (N_7231,N_314,N_3615);
or U7232 (N_7232,N_231,N_3415);
or U7233 (N_7233,N_2151,N_4649);
nand U7234 (N_7234,N_4535,N_4727);
or U7235 (N_7235,N_4133,N_2965);
and U7236 (N_7236,N_2654,N_4822);
and U7237 (N_7237,N_3997,N_2046);
nand U7238 (N_7238,N_1536,N_893);
nand U7239 (N_7239,N_2049,N_2332);
xnor U7240 (N_7240,N_4273,N_4646);
xor U7241 (N_7241,N_357,N_4814);
xnor U7242 (N_7242,N_3325,N_3769);
and U7243 (N_7243,N_3955,N_2626);
or U7244 (N_7244,N_4502,N_3497);
and U7245 (N_7245,N_545,N_4726);
nor U7246 (N_7246,N_1566,N_1863);
nor U7247 (N_7247,N_4911,N_4859);
nand U7248 (N_7248,N_1890,N_2030);
nor U7249 (N_7249,N_2470,N_472);
or U7250 (N_7250,N_4609,N_1162);
nand U7251 (N_7251,N_2636,N_4274);
or U7252 (N_7252,N_270,N_3642);
or U7253 (N_7253,N_2194,N_1518);
and U7254 (N_7254,N_3246,N_3025);
nand U7255 (N_7255,N_1593,N_3205);
nand U7256 (N_7256,N_941,N_4495);
nor U7257 (N_7257,N_4944,N_1378);
or U7258 (N_7258,N_125,N_3728);
nor U7259 (N_7259,N_4011,N_3868);
nand U7260 (N_7260,N_3087,N_1512);
and U7261 (N_7261,N_3490,N_147);
or U7262 (N_7262,N_4627,N_1919);
or U7263 (N_7263,N_2542,N_3566);
nand U7264 (N_7264,N_745,N_3608);
xor U7265 (N_7265,N_4591,N_2);
or U7266 (N_7266,N_3567,N_4633);
or U7267 (N_7267,N_1708,N_3869);
or U7268 (N_7268,N_621,N_900);
and U7269 (N_7269,N_1327,N_3991);
and U7270 (N_7270,N_423,N_3301);
or U7271 (N_7271,N_4370,N_1256);
nor U7272 (N_7272,N_3887,N_2661);
or U7273 (N_7273,N_4272,N_2257);
nand U7274 (N_7274,N_2601,N_2941);
xnor U7275 (N_7275,N_2051,N_4098);
nor U7276 (N_7276,N_3273,N_530);
or U7277 (N_7277,N_3092,N_1342);
or U7278 (N_7278,N_2173,N_1220);
nor U7279 (N_7279,N_886,N_2126);
and U7280 (N_7280,N_3755,N_2468);
nor U7281 (N_7281,N_3789,N_1271);
nand U7282 (N_7282,N_3040,N_4596);
nor U7283 (N_7283,N_220,N_3926);
and U7284 (N_7284,N_2341,N_3682);
nand U7285 (N_7285,N_3637,N_27);
and U7286 (N_7286,N_1313,N_3019);
nand U7287 (N_7287,N_1121,N_4820);
and U7288 (N_7288,N_573,N_223);
nor U7289 (N_7289,N_489,N_4417);
nor U7290 (N_7290,N_2056,N_4403);
nand U7291 (N_7291,N_3182,N_3688);
nand U7292 (N_7292,N_3352,N_1544);
nor U7293 (N_7293,N_3134,N_250);
nand U7294 (N_7294,N_234,N_3661);
and U7295 (N_7295,N_3368,N_840);
nor U7296 (N_7296,N_4283,N_670);
and U7297 (N_7297,N_2749,N_3409);
nand U7298 (N_7298,N_3470,N_549);
nor U7299 (N_7299,N_2153,N_1807);
nand U7300 (N_7300,N_1748,N_1445);
nor U7301 (N_7301,N_2634,N_4861);
nor U7302 (N_7302,N_1808,N_2048);
or U7303 (N_7303,N_560,N_2847);
and U7304 (N_7304,N_4033,N_3083);
and U7305 (N_7305,N_2791,N_684);
nor U7306 (N_7306,N_4044,N_4516);
xor U7307 (N_7307,N_1728,N_4524);
and U7308 (N_7308,N_438,N_4460);
nand U7309 (N_7309,N_495,N_843);
nor U7310 (N_7310,N_1587,N_743);
or U7311 (N_7311,N_2717,N_1556);
nor U7312 (N_7312,N_1191,N_285);
xnor U7313 (N_7313,N_4435,N_630);
xor U7314 (N_7314,N_175,N_4138);
or U7315 (N_7315,N_2283,N_3214);
and U7316 (N_7316,N_2189,N_4246);
and U7317 (N_7317,N_4147,N_4215);
nand U7318 (N_7318,N_82,N_3303);
and U7319 (N_7319,N_4325,N_4833);
nand U7320 (N_7320,N_4152,N_3316);
nor U7321 (N_7321,N_742,N_1788);
or U7322 (N_7322,N_4838,N_1922);
nor U7323 (N_7323,N_3589,N_2526);
nor U7324 (N_7324,N_874,N_667);
nand U7325 (N_7325,N_2670,N_4431);
or U7326 (N_7326,N_4284,N_2956);
nor U7327 (N_7327,N_1152,N_3749);
and U7328 (N_7328,N_428,N_2055);
and U7329 (N_7329,N_4917,N_1538);
xor U7330 (N_7330,N_4662,N_2103);
nand U7331 (N_7331,N_1879,N_189);
xnor U7332 (N_7332,N_2270,N_118);
or U7333 (N_7333,N_151,N_4959);
xor U7334 (N_7334,N_2848,N_333);
nor U7335 (N_7335,N_870,N_4522);
nand U7336 (N_7336,N_3507,N_3063);
or U7337 (N_7337,N_1132,N_2378);
or U7338 (N_7338,N_2165,N_4094);
or U7339 (N_7339,N_4795,N_877);
xor U7340 (N_7340,N_1137,N_2743);
nor U7341 (N_7341,N_4406,N_4459);
nor U7342 (N_7342,N_4432,N_3357);
nor U7343 (N_7343,N_4555,N_2253);
nand U7344 (N_7344,N_578,N_334);
nor U7345 (N_7345,N_1238,N_1290);
nand U7346 (N_7346,N_4064,N_3806);
or U7347 (N_7347,N_470,N_2251);
or U7348 (N_7348,N_2003,N_336);
nand U7349 (N_7349,N_4558,N_1376);
nor U7350 (N_7350,N_1921,N_609);
xor U7351 (N_7351,N_4641,N_1107);
and U7352 (N_7352,N_999,N_2716);
or U7353 (N_7353,N_3323,N_1333);
and U7354 (N_7354,N_4419,N_1104);
or U7355 (N_7355,N_215,N_4476);
or U7356 (N_7356,N_604,N_990);
nor U7357 (N_7357,N_3621,N_679);
nor U7358 (N_7358,N_3885,N_318);
nor U7359 (N_7359,N_4035,N_87);
or U7360 (N_7360,N_4380,N_910);
or U7361 (N_7361,N_1257,N_1898);
and U7362 (N_7362,N_2955,N_209);
xnor U7363 (N_7363,N_4241,N_4885);
or U7364 (N_7364,N_1284,N_779);
and U7365 (N_7365,N_2147,N_483);
and U7366 (N_7366,N_1070,N_1408);
and U7367 (N_7367,N_2123,N_4908);
and U7368 (N_7368,N_891,N_356);
nor U7369 (N_7369,N_1812,N_4565);
nand U7370 (N_7370,N_3269,N_3638);
nand U7371 (N_7371,N_3371,N_2349);
nor U7372 (N_7372,N_3646,N_2575);
nor U7373 (N_7373,N_2629,N_3938);
and U7374 (N_7374,N_21,N_4667);
nand U7375 (N_7375,N_2790,N_4217);
and U7376 (N_7376,N_3233,N_1144);
or U7377 (N_7377,N_1495,N_3349);
and U7378 (N_7378,N_414,N_1861);
and U7379 (N_7379,N_1582,N_4514);
xor U7380 (N_7380,N_2120,N_905);
or U7381 (N_7381,N_484,N_3781);
nand U7382 (N_7382,N_932,N_354);
or U7383 (N_7383,N_4312,N_1525);
or U7384 (N_7384,N_4635,N_2757);
or U7385 (N_7385,N_3146,N_3655);
nand U7386 (N_7386,N_946,N_180);
nor U7387 (N_7387,N_3526,N_1304);
and U7388 (N_7388,N_795,N_2647);
nor U7389 (N_7389,N_81,N_700);
or U7390 (N_7390,N_3587,N_978);
and U7391 (N_7391,N_3678,N_3340);
and U7392 (N_7392,N_2229,N_164);
nor U7393 (N_7393,N_3024,N_1961);
and U7394 (N_7394,N_2330,N_3082);
nand U7395 (N_7395,N_1044,N_4790);
or U7396 (N_7396,N_2413,N_3880);
and U7397 (N_7397,N_1980,N_2477);
nor U7398 (N_7398,N_256,N_4344);
nor U7399 (N_7399,N_3539,N_391);
xnor U7400 (N_7400,N_1197,N_1210);
nor U7401 (N_7401,N_1597,N_1562);
or U7402 (N_7402,N_3778,N_2426);
nand U7403 (N_7403,N_3931,N_1295);
and U7404 (N_7404,N_3148,N_1746);
and U7405 (N_7405,N_1851,N_4480);
nor U7406 (N_7406,N_2556,N_723);
nand U7407 (N_7407,N_4365,N_4265);
and U7408 (N_7408,N_3501,N_4216);
nor U7409 (N_7409,N_418,N_4242);
nand U7410 (N_7410,N_4570,N_3787);
and U7411 (N_7411,N_3872,N_1241);
xor U7412 (N_7412,N_2060,N_4420);
or U7413 (N_7413,N_1978,N_981);
nand U7414 (N_7414,N_2199,N_4415);
nor U7415 (N_7415,N_4041,N_4697);
and U7416 (N_7416,N_4954,N_2709);
or U7417 (N_7417,N_4967,N_3039);
xor U7418 (N_7418,N_3523,N_2518);
and U7419 (N_7419,N_463,N_2157);
or U7420 (N_7420,N_957,N_4914);
nand U7421 (N_7421,N_3427,N_2758);
nor U7422 (N_7422,N_30,N_1434);
nor U7423 (N_7423,N_3599,N_2911);
nor U7424 (N_7424,N_3596,N_3988);
or U7425 (N_7425,N_1594,N_3011);
nor U7426 (N_7426,N_73,N_2839);
nand U7427 (N_7427,N_3895,N_1852);
and U7428 (N_7428,N_2905,N_2990);
or U7429 (N_7429,N_1779,N_4937);
and U7430 (N_7430,N_2192,N_2258);
and U7431 (N_7431,N_1549,N_948);
or U7432 (N_7432,N_304,N_3862);
or U7433 (N_7433,N_4112,N_3979);
xor U7434 (N_7434,N_3619,N_3101);
nor U7435 (N_7435,N_3421,N_2722);
and U7436 (N_7436,N_3347,N_2354);
or U7437 (N_7437,N_2742,N_2050);
nand U7438 (N_7438,N_3242,N_2724);
or U7439 (N_7439,N_4018,N_117);
nor U7440 (N_7440,N_47,N_1766);
and U7441 (N_7441,N_1142,N_3474);
and U7442 (N_7442,N_520,N_704);
and U7443 (N_7443,N_741,N_3436);
nand U7444 (N_7444,N_2794,N_3327);
or U7445 (N_7445,N_3851,N_2450);
nor U7446 (N_7446,N_921,N_1018);
or U7447 (N_7447,N_3866,N_4017);
nor U7448 (N_7448,N_2318,N_4337);
or U7449 (N_7449,N_1951,N_4400);
nand U7450 (N_7450,N_1276,N_3743);
nor U7451 (N_7451,N_131,N_589);
nor U7452 (N_7452,N_4393,N_1089);
or U7453 (N_7453,N_2207,N_1285);
and U7454 (N_7454,N_3265,N_402);
nor U7455 (N_7455,N_2272,N_3494);
nand U7456 (N_7456,N_804,N_1254);
or U7457 (N_7457,N_4660,N_4769);
xor U7458 (N_7458,N_4532,N_2768);
or U7459 (N_7459,N_2989,N_970);
or U7460 (N_7460,N_2307,N_3513);
nand U7461 (N_7461,N_4328,N_775);
and U7462 (N_7462,N_100,N_2599);
and U7463 (N_7463,N_3912,N_3653);
nor U7464 (N_7464,N_3305,N_4250);
nand U7465 (N_7465,N_4221,N_112);
nand U7466 (N_7466,N_4714,N_3662);
xor U7467 (N_7467,N_975,N_1123);
xnor U7468 (N_7468,N_328,N_2308);
nor U7469 (N_7469,N_4571,N_4346);
xnor U7470 (N_7470,N_3804,N_161);
nand U7471 (N_7471,N_144,N_2627);
nand U7472 (N_7472,N_766,N_2878);
and U7473 (N_7473,N_1548,N_619);
or U7474 (N_7474,N_3732,N_2326);
or U7475 (N_7475,N_46,N_2806);
and U7476 (N_7476,N_4226,N_4109);
and U7477 (N_7477,N_3338,N_4768);
and U7478 (N_7478,N_261,N_1268);
xor U7479 (N_7479,N_158,N_1038);
or U7480 (N_7480,N_646,N_2745);
and U7481 (N_7481,N_1936,N_188);
and U7482 (N_7482,N_267,N_2772);
nor U7483 (N_7483,N_4251,N_2784);
or U7484 (N_7484,N_1707,N_4470);
nor U7485 (N_7485,N_2115,N_3055);
or U7486 (N_7486,N_2917,N_1680);
and U7487 (N_7487,N_427,N_3457);
nand U7488 (N_7488,N_2461,N_1054);
and U7489 (N_7489,N_3742,N_1661);
or U7490 (N_7490,N_4090,N_3689);
nor U7491 (N_7491,N_3038,N_3694);
and U7492 (N_7492,N_2457,N_4511);
nor U7493 (N_7493,N_167,N_2803);
xnor U7494 (N_7494,N_3439,N_1836);
nand U7495 (N_7495,N_4915,N_3736);
xor U7496 (N_7496,N_2523,N_4593);
xnor U7497 (N_7497,N_19,N_740);
and U7498 (N_7498,N_3048,N_1074);
xnor U7499 (N_7499,N_615,N_4541);
nor U7500 (N_7500,N_2207,N_1708);
and U7501 (N_7501,N_3467,N_2517);
nor U7502 (N_7502,N_2723,N_2505);
or U7503 (N_7503,N_1699,N_3180);
and U7504 (N_7504,N_1023,N_3261);
and U7505 (N_7505,N_424,N_516);
or U7506 (N_7506,N_2120,N_2779);
nand U7507 (N_7507,N_1789,N_63);
and U7508 (N_7508,N_1323,N_2972);
or U7509 (N_7509,N_4919,N_1768);
or U7510 (N_7510,N_3537,N_2457);
nor U7511 (N_7511,N_4703,N_1788);
nand U7512 (N_7512,N_588,N_3562);
nor U7513 (N_7513,N_1435,N_2694);
and U7514 (N_7514,N_3204,N_4140);
or U7515 (N_7515,N_1822,N_4692);
nand U7516 (N_7516,N_1189,N_1463);
and U7517 (N_7517,N_2359,N_354);
nand U7518 (N_7518,N_4039,N_2726);
or U7519 (N_7519,N_726,N_4900);
or U7520 (N_7520,N_1357,N_2132);
nand U7521 (N_7521,N_761,N_3294);
nand U7522 (N_7522,N_3580,N_3243);
nand U7523 (N_7523,N_3744,N_1748);
and U7524 (N_7524,N_514,N_3337);
nand U7525 (N_7525,N_833,N_1852);
nand U7526 (N_7526,N_4362,N_2730);
and U7527 (N_7527,N_1533,N_1750);
or U7528 (N_7528,N_4889,N_988);
nand U7529 (N_7529,N_1927,N_2843);
or U7530 (N_7530,N_742,N_4251);
and U7531 (N_7531,N_4033,N_3622);
nand U7532 (N_7532,N_3437,N_2686);
and U7533 (N_7533,N_1888,N_574);
and U7534 (N_7534,N_2202,N_4012);
xor U7535 (N_7535,N_1598,N_2177);
nand U7536 (N_7536,N_4656,N_4969);
xnor U7537 (N_7537,N_986,N_186);
nor U7538 (N_7538,N_731,N_651);
nor U7539 (N_7539,N_3260,N_2909);
and U7540 (N_7540,N_1081,N_2488);
xnor U7541 (N_7541,N_4450,N_4667);
nor U7542 (N_7542,N_3787,N_3411);
nand U7543 (N_7543,N_2633,N_2889);
nand U7544 (N_7544,N_2786,N_1449);
or U7545 (N_7545,N_1035,N_2541);
and U7546 (N_7546,N_4153,N_4002);
and U7547 (N_7547,N_2964,N_165);
nor U7548 (N_7548,N_1296,N_2539);
and U7549 (N_7549,N_448,N_3245);
nand U7550 (N_7550,N_1874,N_3013);
and U7551 (N_7551,N_4415,N_821);
or U7552 (N_7552,N_4567,N_1912);
nand U7553 (N_7553,N_3483,N_2560);
nor U7554 (N_7554,N_3801,N_2);
xnor U7555 (N_7555,N_4765,N_248);
nand U7556 (N_7556,N_3640,N_2495);
and U7557 (N_7557,N_3855,N_3589);
and U7558 (N_7558,N_452,N_1312);
and U7559 (N_7559,N_1496,N_1827);
and U7560 (N_7560,N_3277,N_3666);
nand U7561 (N_7561,N_3415,N_1685);
and U7562 (N_7562,N_1178,N_2052);
or U7563 (N_7563,N_2816,N_2235);
nor U7564 (N_7564,N_3410,N_157);
xor U7565 (N_7565,N_982,N_4327);
xor U7566 (N_7566,N_4255,N_3004);
or U7567 (N_7567,N_3517,N_2286);
and U7568 (N_7568,N_4987,N_4967);
xor U7569 (N_7569,N_3403,N_699);
or U7570 (N_7570,N_1203,N_114);
nor U7571 (N_7571,N_285,N_1046);
nand U7572 (N_7572,N_4695,N_4644);
and U7573 (N_7573,N_4440,N_3758);
nor U7574 (N_7574,N_421,N_935);
and U7575 (N_7575,N_3038,N_2917);
or U7576 (N_7576,N_2571,N_1962);
and U7577 (N_7577,N_4345,N_2917);
and U7578 (N_7578,N_3011,N_2115);
nor U7579 (N_7579,N_587,N_495);
xnor U7580 (N_7580,N_553,N_4350);
and U7581 (N_7581,N_149,N_2757);
and U7582 (N_7582,N_3659,N_1486);
nor U7583 (N_7583,N_4828,N_668);
and U7584 (N_7584,N_3987,N_1644);
or U7585 (N_7585,N_4818,N_4991);
and U7586 (N_7586,N_1488,N_4006);
nand U7587 (N_7587,N_2785,N_423);
and U7588 (N_7588,N_4906,N_1788);
nand U7589 (N_7589,N_4699,N_985);
nand U7590 (N_7590,N_4569,N_2970);
nor U7591 (N_7591,N_1088,N_859);
or U7592 (N_7592,N_985,N_1348);
or U7593 (N_7593,N_2762,N_4813);
nor U7594 (N_7594,N_3891,N_3522);
nand U7595 (N_7595,N_4216,N_1329);
nor U7596 (N_7596,N_842,N_2718);
xnor U7597 (N_7597,N_1331,N_1356);
xnor U7598 (N_7598,N_4937,N_4915);
nand U7599 (N_7599,N_230,N_3738);
xnor U7600 (N_7600,N_4581,N_4881);
xor U7601 (N_7601,N_1570,N_710);
or U7602 (N_7602,N_4400,N_670);
or U7603 (N_7603,N_597,N_2347);
and U7604 (N_7604,N_266,N_4003);
and U7605 (N_7605,N_1627,N_331);
xor U7606 (N_7606,N_1967,N_2059);
xnor U7607 (N_7607,N_4965,N_2676);
or U7608 (N_7608,N_4689,N_2837);
and U7609 (N_7609,N_550,N_3195);
nand U7610 (N_7610,N_3402,N_1753);
and U7611 (N_7611,N_2014,N_2587);
nand U7612 (N_7612,N_393,N_1913);
and U7613 (N_7613,N_3904,N_3485);
nor U7614 (N_7614,N_3585,N_3983);
nand U7615 (N_7615,N_2233,N_4333);
xor U7616 (N_7616,N_2222,N_1437);
nor U7617 (N_7617,N_4608,N_953);
nand U7618 (N_7618,N_3954,N_3115);
and U7619 (N_7619,N_1308,N_1289);
nor U7620 (N_7620,N_1751,N_1054);
xnor U7621 (N_7621,N_2346,N_3965);
nor U7622 (N_7622,N_1556,N_4920);
and U7623 (N_7623,N_769,N_4831);
xor U7624 (N_7624,N_881,N_4260);
or U7625 (N_7625,N_3018,N_3191);
nand U7626 (N_7626,N_2092,N_1677);
nor U7627 (N_7627,N_1907,N_4481);
nor U7628 (N_7628,N_2172,N_114);
or U7629 (N_7629,N_170,N_1143);
nor U7630 (N_7630,N_774,N_229);
or U7631 (N_7631,N_3245,N_1021);
xor U7632 (N_7632,N_4964,N_572);
and U7633 (N_7633,N_697,N_765);
xnor U7634 (N_7634,N_4600,N_1538);
nand U7635 (N_7635,N_1772,N_2372);
nand U7636 (N_7636,N_1997,N_3029);
and U7637 (N_7637,N_3641,N_3637);
nand U7638 (N_7638,N_4438,N_3456);
and U7639 (N_7639,N_2194,N_3595);
nand U7640 (N_7640,N_3453,N_137);
nand U7641 (N_7641,N_695,N_4276);
nor U7642 (N_7642,N_129,N_3199);
or U7643 (N_7643,N_129,N_1667);
and U7644 (N_7644,N_2649,N_3300);
or U7645 (N_7645,N_4662,N_4035);
nand U7646 (N_7646,N_1445,N_2225);
or U7647 (N_7647,N_4163,N_114);
and U7648 (N_7648,N_2327,N_2408);
and U7649 (N_7649,N_4204,N_884);
nor U7650 (N_7650,N_4899,N_2436);
nand U7651 (N_7651,N_3823,N_2597);
and U7652 (N_7652,N_2204,N_104);
or U7653 (N_7653,N_3586,N_3516);
or U7654 (N_7654,N_4898,N_265);
nor U7655 (N_7655,N_3905,N_2291);
and U7656 (N_7656,N_3962,N_1010);
and U7657 (N_7657,N_243,N_1607);
or U7658 (N_7658,N_4754,N_3877);
nor U7659 (N_7659,N_4560,N_533);
and U7660 (N_7660,N_2180,N_3356);
nor U7661 (N_7661,N_3356,N_3155);
nor U7662 (N_7662,N_2530,N_719);
nand U7663 (N_7663,N_4326,N_895);
and U7664 (N_7664,N_4741,N_1422);
xor U7665 (N_7665,N_4027,N_4943);
nor U7666 (N_7666,N_4038,N_1360);
and U7667 (N_7667,N_3582,N_4668);
or U7668 (N_7668,N_474,N_2463);
or U7669 (N_7669,N_1953,N_4034);
nor U7670 (N_7670,N_3630,N_2514);
nand U7671 (N_7671,N_3268,N_2770);
or U7672 (N_7672,N_116,N_3124);
or U7673 (N_7673,N_3614,N_4847);
or U7674 (N_7674,N_4417,N_1206);
nand U7675 (N_7675,N_1824,N_4362);
nand U7676 (N_7676,N_924,N_3508);
or U7677 (N_7677,N_3164,N_1767);
nor U7678 (N_7678,N_4286,N_2433);
nand U7679 (N_7679,N_2689,N_1910);
and U7680 (N_7680,N_3464,N_1901);
nand U7681 (N_7681,N_2700,N_4955);
and U7682 (N_7682,N_959,N_906);
xnor U7683 (N_7683,N_3513,N_937);
nor U7684 (N_7684,N_4152,N_230);
and U7685 (N_7685,N_4275,N_2648);
nand U7686 (N_7686,N_83,N_4487);
nand U7687 (N_7687,N_4,N_3504);
and U7688 (N_7688,N_2831,N_1753);
nor U7689 (N_7689,N_802,N_276);
and U7690 (N_7690,N_4592,N_4052);
nand U7691 (N_7691,N_945,N_3457);
and U7692 (N_7692,N_2701,N_1170);
nand U7693 (N_7693,N_521,N_3890);
nor U7694 (N_7694,N_1135,N_1010);
nand U7695 (N_7695,N_2379,N_3298);
nand U7696 (N_7696,N_2850,N_2336);
nand U7697 (N_7697,N_600,N_4422);
nand U7698 (N_7698,N_983,N_3455);
or U7699 (N_7699,N_4282,N_2569);
nand U7700 (N_7700,N_3275,N_4325);
and U7701 (N_7701,N_4706,N_413);
or U7702 (N_7702,N_1372,N_1189);
and U7703 (N_7703,N_1331,N_2608);
or U7704 (N_7704,N_3841,N_1170);
nor U7705 (N_7705,N_4889,N_618);
nand U7706 (N_7706,N_619,N_599);
nand U7707 (N_7707,N_1009,N_1894);
nand U7708 (N_7708,N_3365,N_4840);
or U7709 (N_7709,N_1558,N_2653);
or U7710 (N_7710,N_3849,N_1867);
nor U7711 (N_7711,N_1511,N_4512);
and U7712 (N_7712,N_2456,N_4573);
nand U7713 (N_7713,N_2321,N_568);
nand U7714 (N_7714,N_617,N_2941);
nor U7715 (N_7715,N_4954,N_2215);
nand U7716 (N_7716,N_339,N_2663);
or U7717 (N_7717,N_3763,N_1361);
nor U7718 (N_7718,N_2917,N_2204);
nand U7719 (N_7719,N_3448,N_1430);
nor U7720 (N_7720,N_666,N_2816);
xor U7721 (N_7721,N_4033,N_3536);
or U7722 (N_7722,N_4715,N_4252);
or U7723 (N_7723,N_3982,N_1287);
nand U7724 (N_7724,N_392,N_4547);
nand U7725 (N_7725,N_2789,N_2632);
or U7726 (N_7726,N_3646,N_1394);
nand U7727 (N_7727,N_3995,N_3931);
nor U7728 (N_7728,N_2757,N_3582);
or U7729 (N_7729,N_4022,N_2836);
and U7730 (N_7730,N_4620,N_2339);
or U7731 (N_7731,N_3811,N_2028);
or U7732 (N_7732,N_4321,N_2514);
and U7733 (N_7733,N_3316,N_3133);
nor U7734 (N_7734,N_2163,N_1426);
nor U7735 (N_7735,N_4178,N_1799);
or U7736 (N_7736,N_162,N_3060);
or U7737 (N_7737,N_2283,N_2015);
nor U7738 (N_7738,N_2612,N_1833);
nor U7739 (N_7739,N_2941,N_2679);
nor U7740 (N_7740,N_3342,N_1755);
and U7741 (N_7741,N_3844,N_1986);
or U7742 (N_7742,N_2228,N_4988);
or U7743 (N_7743,N_3407,N_1210);
or U7744 (N_7744,N_1137,N_1771);
or U7745 (N_7745,N_491,N_3559);
nor U7746 (N_7746,N_1608,N_2846);
xnor U7747 (N_7747,N_171,N_3417);
and U7748 (N_7748,N_784,N_3774);
and U7749 (N_7749,N_3521,N_1403);
or U7750 (N_7750,N_4137,N_486);
or U7751 (N_7751,N_688,N_4720);
nor U7752 (N_7752,N_3563,N_1504);
nor U7753 (N_7753,N_1894,N_4380);
nand U7754 (N_7754,N_3223,N_1056);
and U7755 (N_7755,N_750,N_1326);
and U7756 (N_7756,N_1803,N_2724);
and U7757 (N_7757,N_1896,N_3613);
and U7758 (N_7758,N_3842,N_349);
nand U7759 (N_7759,N_2668,N_4875);
nand U7760 (N_7760,N_727,N_4875);
nand U7761 (N_7761,N_3783,N_3299);
nor U7762 (N_7762,N_318,N_4546);
nor U7763 (N_7763,N_1940,N_4659);
nand U7764 (N_7764,N_2658,N_3906);
and U7765 (N_7765,N_1026,N_2996);
nand U7766 (N_7766,N_1540,N_1311);
xor U7767 (N_7767,N_586,N_2518);
and U7768 (N_7768,N_855,N_1024);
nand U7769 (N_7769,N_3656,N_3359);
nor U7770 (N_7770,N_4172,N_669);
nor U7771 (N_7771,N_4181,N_1085);
nand U7772 (N_7772,N_2554,N_2798);
or U7773 (N_7773,N_1026,N_869);
or U7774 (N_7774,N_4784,N_2583);
and U7775 (N_7775,N_1583,N_4041);
nor U7776 (N_7776,N_1105,N_3273);
nor U7777 (N_7777,N_441,N_3842);
nand U7778 (N_7778,N_2419,N_614);
and U7779 (N_7779,N_718,N_1491);
nor U7780 (N_7780,N_299,N_4975);
and U7781 (N_7781,N_3622,N_2784);
and U7782 (N_7782,N_3540,N_4695);
and U7783 (N_7783,N_4221,N_1957);
nor U7784 (N_7784,N_1639,N_4012);
xnor U7785 (N_7785,N_4047,N_1381);
xor U7786 (N_7786,N_2873,N_1638);
and U7787 (N_7787,N_299,N_4626);
nor U7788 (N_7788,N_2411,N_338);
or U7789 (N_7789,N_1857,N_486);
nor U7790 (N_7790,N_2286,N_1156);
or U7791 (N_7791,N_3487,N_7);
and U7792 (N_7792,N_1180,N_1150);
and U7793 (N_7793,N_2806,N_3972);
nor U7794 (N_7794,N_2711,N_2327);
nand U7795 (N_7795,N_4740,N_1667);
xor U7796 (N_7796,N_3769,N_2170);
and U7797 (N_7797,N_4553,N_857);
nor U7798 (N_7798,N_3758,N_3855);
or U7799 (N_7799,N_1137,N_940);
or U7800 (N_7800,N_486,N_4465);
and U7801 (N_7801,N_2660,N_3828);
xnor U7802 (N_7802,N_1644,N_3830);
and U7803 (N_7803,N_1884,N_3360);
nand U7804 (N_7804,N_4537,N_2166);
or U7805 (N_7805,N_2703,N_3865);
nor U7806 (N_7806,N_3859,N_983);
and U7807 (N_7807,N_1710,N_2260);
nand U7808 (N_7808,N_2749,N_3790);
xor U7809 (N_7809,N_4191,N_3563);
nand U7810 (N_7810,N_732,N_3524);
nor U7811 (N_7811,N_2272,N_2055);
nand U7812 (N_7812,N_410,N_4208);
nand U7813 (N_7813,N_3781,N_2267);
and U7814 (N_7814,N_730,N_417);
and U7815 (N_7815,N_2877,N_4534);
and U7816 (N_7816,N_3963,N_3394);
nor U7817 (N_7817,N_1582,N_3565);
and U7818 (N_7818,N_4447,N_1544);
and U7819 (N_7819,N_3662,N_1834);
or U7820 (N_7820,N_1687,N_1579);
and U7821 (N_7821,N_299,N_2576);
nor U7822 (N_7822,N_769,N_490);
or U7823 (N_7823,N_3835,N_1268);
nor U7824 (N_7824,N_4377,N_1642);
and U7825 (N_7825,N_364,N_3417);
nor U7826 (N_7826,N_1123,N_4038);
and U7827 (N_7827,N_4628,N_4632);
or U7828 (N_7828,N_478,N_1017);
or U7829 (N_7829,N_3886,N_4864);
or U7830 (N_7830,N_970,N_4755);
nand U7831 (N_7831,N_425,N_2459);
and U7832 (N_7832,N_37,N_1783);
and U7833 (N_7833,N_1017,N_4602);
nand U7834 (N_7834,N_3872,N_3357);
and U7835 (N_7835,N_1620,N_302);
nand U7836 (N_7836,N_4260,N_442);
nand U7837 (N_7837,N_1425,N_4265);
xor U7838 (N_7838,N_2900,N_2435);
nor U7839 (N_7839,N_415,N_4316);
nor U7840 (N_7840,N_4234,N_1262);
and U7841 (N_7841,N_3858,N_4979);
and U7842 (N_7842,N_1366,N_320);
xnor U7843 (N_7843,N_4102,N_3043);
nor U7844 (N_7844,N_1190,N_1353);
or U7845 (N_7845,N_1708,N_977);
nand U7846 (N_7846,N_3985,N_3504);
and U7847 (N_7847,N_2391,N_2027);
nand U7848 (N_7848,N_4148,N_378);
nand U7849 (N_7849,N_4076,N_210);
or U7850 (N_7850,N_545,N_328);
nand U7851 (N_7851,N_1025,N_2732);
nor U7852 (N_7852,N_1451,N_679);
nand U7853 (N_7853,N_3288,N_1663);
nor U7854 (N_7854,N_4596,N_1351);
and U7855 (N_7855,N_2306,N_2332);
nand U7856 (N_7856,N_1158,N_4258);
and U7857 (N_7857,N_2750,N_1338);
or U7858 (N_7858,N_4340,N_4694);
or U7859 (N_7859,N_4298,N_2570);
and U7860 (N_7860,N_1578,N_2619);
nand U7861 (N_7861,N_2727,N_872);
or U7862 (N_7862,N_2568,N_3433);
nor U7863 (N_7863,N_238,N_2686);
nor U7864 (N_7864,N_3043,N_1320);
nand U7865 (N_7865,N_2582,N_2679);
nor U7866 (N_7866,N_4522,N_3652);
nand U7867 (N_7867,N_853,N_4311);
nor U7868 (N_7868,N_3376,N_3554);
nor U7869 (N_7869,N_1167,N_897);
and U7870 (N_7870,N_3070,N_4263);
and U7871 (N_7871,N_4731,N_3769);
or U7872 (N_7872,N_465,N_2510);
and U7873 (N_7873,N_739,N_1220);
or U7874 (N_7874,N_3243,N_4050);
or U7875 (N_7875,N_3823,N_3635);
or U7876 (N_7876,N_1543,N_3641);
nor U7877 (N_7877,N_128,N_1859);
nor U7878 (N_7878,N_2068,N_2722);
xor U7879 (N_7879,N_4753,N_4445);
or U7880 (N_7880,N_3515,N_1082);
or U7881 (N_7881,N_2939,N_3692);
and U7882 (N_7882,N_4720,N_3863);
and U7883 (N_7883,N_1679,N_3164);
or U7884 (N_7884,N_2897,N_1577);
or U7885 (N_7885,N_2300,N_4547);
nand U7886 (N_7886,N_4773,N_2661);
and U7887 (N_7887,N_884,N_1523);
xnor U7888 (N_7888,N_4760,N_143);
or U7889 (N_7889,N_4408,N_2997);
nor U7890 (N_7890,N_4274,N_2531);
nor U7891 (N_7891,N_2033,N_3750);
and U7892 (N_7892,N_2099,N_3836);
and U7893 (N_7893,N_4313,N_19);
nand U7894 (N_7894,N_1100,N_3902);
and U7895 (N_7895,N_3769,N_4162);
nand U7896 (N_7896,N_3915,N_3034);
nand U7897 (N_7897,N_4605,N_3505);
xor U7898 (N_7898,N_348,N_2322);
and U7899 (N_7899,N_1005,N_687);
nor U7900 (N_7900,N_3019,N_3236);
or U7901 (N_7901,N_2515,N_644);
nand U7902 (N_7902,N_627,N_2652);
nand U7903 (N_7903,N_1687,N_2253);
and U7904 (N_7904,N_4069,N_3971);
nor U7905 (N_7905,N_3314,N_3745);
nand U7906 (N_7906,N_974,N_1747);
nor U7907 (N_7907,N_2332,N_3304);
and U7908 (N_7908,N_4547,N_3413);
or U7909 (N_7909,N_3163,N_4593);
nor U7910 (N_7910,N_3232,N_4353);
and U7911 (N_7911,N_738,N_3531);
and U7912 (N_7912,N_1906,N_1771);
xnor U7913 (N_7913,N_3340,N_860);
and U7914 (N_7914,N_3480,N_4288);
xor U7915 (N_7915,N_1929,N_3730);
nand U7916 (N_7916,N_2040,N_4985);
nor U7917 (N_7917,N_1512,N_823);
nand U7918 (N_7918,N_1025,N_1162);
or U7919 (N_7919,N_100,N_1316);
xnor U7920 (N_7920,N_763,N_1613);
or U7921 (N_7921,N_2846,N_1754);
and U7922 (N_7922,N_4976,N_3429);
or U7923 (N_7923,N_2412,N_4194);
nand U7924 (N_7924,N_194,N_2233);
nand U7925 (N_7925,N_256,N_3924);
nand U7926 (N_7926,N_1228,N_3546);
nand U7927 (N_7927,N_3076,N_4222);
nor U7928 (N_7928,N_4539,N_1573);
nor U7929 (N_7929,N_1735,N_2679);
and U7930 (N_7930,N_401,N_1229);
and U7931 (N_7931,N_4382,N_1574);
nor U7932 (N_7932,N_2560,N_1269);
or U7933 (N_7933,N_1079,N_2219);
nand U7934 (N_7934,N_1025,N_3482);
nand U7935 (N_7935,N_4646,N_4258);
xor U7936 (N_7936,N_2283,N_1067);
nor U7937 (N_7937,N_2450,N_3681);
or U7938 (N_7938,N_1923,N_4381);
or U7939 (N_7939,N_2604,N_2360);
and U7940 (N_7940,N_710,N_3371);
nor U7941 (N_7941,N_3542,N_2067);
nor U7942 (N_7942,N_2865,N_3508);
or U7943 (N_7943,N_1226,N_2059);
or U7944 (N_7944,N_2950,N_4508);
or U7945 (N_7945,N_4440,N_3389);
nand U7946 (N_7946,N_1031,N_2371);
or U7947 (N_7947,N_2932,N_422);
nor U7948 (N_7948,N_4784,N_1306);
or U7949 (N_7949,N_695,N_2809);
nor U7950 (N_7950,N_1296,N_242);
and U7951 (N_7951,N_4214,N_2385);
and U7952 (N_7952,N_2789,N_4201);
nor U7953 (N_7953,N_1716,N_2993);
nand U7954 (N_7954,N_2199,N_3987);
and U7955 (N_7955,N_3511,N_1839);
and U7956 (N_7956,N_4675,N_3458);
xor U7957 (N_7957,N_3117,N_3816);
or U7958 (N_7958,N_4602,N_4553);
or U7959 (N_7959,N_1084,N_2375);
nor U7960 (N_7960,N_2221,N_205);
and U7961 (N_7961,N_569,N_4048);
and U7962 (N_7962,N_4790,N_4172);
nor U7963 (N_7963,N_2989,N_4327);
or U7964 (N_7964,N_2359,N_2214);
and U7965 (N_7965,N_3976,N_2168);
and U7966 (N_7966,N_4510,N_1535);
and U7967 (N_7967,N_1810,N_4588);
nor U7968 (N_7968,N_4049,N_4);
nor U7969 (N_7969,N_2650,N_3048);
or U7970 (N_7970,N_803,N_4060);
or U7971 (N_7971,N_4045,N_235);
nand U7972 (N_7972,N_2786,N_2410);
nand U7973 (N_7973,N_206,N_1343);
and U7974 (N_7974,N_3969,N_1104);
or U7975 (N_7975,N_3165,N_368);
and U7976 (N_7976,N_539,N_1902);
or U7977 (N_7977,N_3094,N_1875);
nand U7978 (N_7978,N_1175,N_449);
and U7979 (N_7979,N_1655,N_43);
nand U7980 (N_7980,N_4796,N_3999);
nor U7981 (N_7981,N_3273,N_1047);
xnor U7982 (N_7982,N_3344,N_4502);
or U7983 (N_7983,N_3897,N_1786);
nand U7984 (N_7984,N_1261,N_4535);
or U7985 (N_7985,N_2305,N_4042);
nand U7986 (N_7986,N_4801,N_4393);
or U7987 (N_7987,N_4167,N_263);
nand U7988 (N_7988,N_3976,N_2337);
and U7989 (N_7989,N_4263,N_3423);
and U7990 (N_7990,N_925,N_3012);
and U7991 (N_7991,N_3287,N_1742);
nor U7992 (N_7992,N_4101,N_2982);
nor U7993 (N_7993,N_180,N_1958);
nand U7994 (N_7994,N_326,N_4944);
nor U7995 (N_7995,N_3071,N_520);
or U7996 (N_7996,N_2199,N_2930);
nor U7997 (N_7997,N_1210,N_1550);
xor U7998 (N_7998,N_1681,N_1112);
and U7999 (N_7999,N_2247,N_366);
nor U8000 (N_8000,N_3551,N_266);
nand U8001 (N_8001,N_1923,N_1306);
nor U8002 (N_8002,N_2032,N_212);
or U8003 (N_8003,N_3918,N_142);
nor U8004 (N_8004,N_1549,N_2926);
or U8005 (N_8005,N_4458,N_525);
xnor U8006 (N_8006,N_3118,N_2889);
nand U8007 (N_8007,N_1725,N_3720);
and U8008 (N_8008,N_3669,N_2567);
nand U8009 (N_8009,N_116,N_2053);
nand U8010 (N_8010,N_2807,N_2591);
or U8011 (N_8011,N_2989,N_4613);
or U8012 (N_8012,N_2576,N_4260);
xnor U8013 (N_8013,N_305,N_740);
nor U8014 (N_8014,N_3570,N_843);
or U8015 (N_8015,N_2066,N_1278);
and U8016 (N_8016,N_4266,N_2623);
nor U8017 (N_8017,N_2191,N_470);
nor U8018 (N_8018,N_2310,N_21);
xor U8019 (N_8019,N_811,N_1952);
xnor U8020 (N_8020,N_4718,N_2933);
or U8021 (N_8021,N_4244,N_237);
nor U8022 (N_8022,N_4236,N_1103);
nor U8023 (N_8023,N_264,N_1068);
nand U8024 (N_8024,N_1592,N_596);
nor U8025 (N_8025,N_3346,N_1339);
nor U8026 (N_8026,N_39,N_265);
or U8027 (N_8027,N_527,N_4486);
nand U8028 (N_8028,N_320,N_1874);
or U8029 (N_8029,N_4018,N_2717);
and U8030 (N_8030,N_4451,N_762);
or U8031 (N_8031,N_504,N_1886);
nand U8032 (N_8032,N_334,N_1227);
xor U8033 (N_8033,N_3427,N_3678);
xor U8034 (N_8034,N_4553,N_1505);
nand U8035 (N_8035,N_3035,N_2803);
nand U8036 (N_8036,N_3729,N_2501);
nand U8037 (N_8037,N_2993,N_716);
and U8038 (N_8038,N_784,N_3095);
nand U8039 (N_8039,N_2424,N_1894);
or U8040 (N_8040,N_4787,N_4393);
or U8041 (N_8041,N_3443,N_4439);
nand U8042 (N_8042,N_4957,N_4620);
and U8043 (N_8043,N_79,N_3929);
or U8044 (N_8044,N_2847,N_1182);
xor U8045 (N_8045,N_3796,N_3221);
nand U8046 (N_8046,N_423,N_4555);
xnor U8047 (N_8047,N_1054,N_3101);
and U8048 (N_8048,N_504,N_3501);
and U8049 (N_8049,N_4380,N_3426);
and U8050 (N_8050,N_4911,N_2827);
and U8051 (N_8051,N_1248,N_4809);
xor U8052 (N_8052,N_4571,N_2506);
and U8053 (N_8053,N_3580,N_771);
and U8054 (N_8054,N_2584,N_1683);
nor U8055 (N_8055,N_1896,N_435);
xor U8056 (N_8056,N_4584,N_2096);
nand U8057 (N_8057,N_4837,N_1450);
and U8058 (N_8058,N_4643,N_1506);
nor U8059 (N_8059,N_4799,N_2621);
nand U8060 (N_8060,N_4379,N_3761);
or U8061 (N_8061,N_4238,N_3209);
xnor U8062 (N_8062,N_2084,N_2016);
and U8063 (N_8063,N_208,N_4240);
or U8064 (N_8064,N_3570,N_2064);
or U8065 (N_8065,N_4107,N_1305);
or U8066 (N_8066,N_955,N_2692);
xor U8067 (N_8067,N_2976,N_4936);
or U8068 (N_8068,N_3350,N_1601);
or U8069 (N_8069,N_4257,N_1251);
nand U8070 (N_8070,N_678,N_1933);
or U8071 (N_8071,N_632,N_270);
nand U8072 (N_8072,N_4034,N_2758);
nand U8073 (N_8073,N_2715,N_1407);
xnor U8074 (N_8074,N_3407,N_912);
or U8075 (N_8075,N_3855,N_3437);
or U8076 (N_8076,N_1886,N_2881);
nor U8077 (N_8077,N_4294,N_171);
xnor U8078 (N_8078,N_2484,N_90);
xor U8079 (N_8079,N_3321,N_3441);
and U8080 (N_8080,N_3916,N_253);
xnor U8081 (N_8081,N_2476,N_3466);
nand U8082 (N_8082,N_1048,N_600);
and U8083 (N_8083,N_241,N_2036);
or U8084 (N_8084,N_2805,N_4379);
nand U8085 (N_8085,N_270,N_4027);
and U8086 (N_8086,N_4033,N_1491);
nand U8087 (N_8087,N_3172,N_591);
and U8088 (N_8088,N_2861,N_199);
nor U8089 (N_8089,N_1932,N_4091);
and U8090 (N_8090,N_1714,N_2852);
and U8091 (N_8091,N_2293,N_1125);
and U8092 (N_8092,N_562,N_4179);
nand U8093 (N_8093,N_3110,N_2074);
nand U8094 (N_8094,N_3262,N_3878);
nand U8095 (N_8095,N_1559,N_2989);
nor U8096 (N_8096,N_4278,N_3755);
or U8097 (N_8097,N_2387,N_4016);
or U8098 (N_8098,N_3436,N_589);
and U8099 (N_8099,N_2166,N_4006);
nand U8100 (N_8100,N_1121,N_3476);
or U8101 (N_8101,N_1922,N_1646);
nand U8102 (N_8102,N_378,N_4283);
nor U8103 (N_8103,N_3165,N_3956);
and U8104 (N_8104,N_4226,N_1378);
and U8105 (N_8105,N_1817,N_3736);
and U8106 (N_8106,N_1797,N_860);
or U8107 (N_8107,N_3119,N_794);
and U8108 (N_8108,N_1175,N_1183);
or U8109 (N_8109,N_2684,N_3834);
or U8110 (N_8110,N_4433,N_3350);
nand U8111 (N_8111,N_4095,N_567);
and U8112 (N_8112,N_343,N_1189);
or U8113 (N_8113,N_243,N_3032);
or U8114 (N_8114,N_567,N_2490);
or U8115 (N_8115,N_3459,N_3632);
nor U8116 (N_8116,N_1557,N_1298);
or U8117 (N_8117,N_1466,N_3220);
xor U8118 (N_8118,N_3161,N_4028);
or U8119 (N_8119,N_3695,N_2395);
and U8120 (N_8120,N_2628,N_2370);
nor U8121 (N_8121,N_2356,N_948);
nand U8122 (N_8122,N_3382,N_4936);
nor U8123 (N_8123,N_2406,N_591);
nor U8124 (N_8124,N_378,N_1135);
nor U8125 (N_8125,N_4858,N_324);
nor U8126 (N_8126,N_2204,N_1530);
nand U8127 (N_8127,N_3965,N_2975);
nand U8128 (N_8128,N_2447,N_3310);
nand U8129 (N_8129,N_105,N_4280);
xnor U8130 (N_8130,N_82,N_3444);
nor U8131 (N_8131,N_4345,N_2770);
nor U8132 (N_8132,N_4208,N_2196);
nand U8133 (N_8133,N_4028,N_1859);
and U8134 (N_8134,N_2270,N_3747);
and U8135 (N_8135,N_4105,N_2442);
nor U8136 (N_8136,N_2424,N_1059);
or U8137 (N_8137,N_2708,N_21);
nand U8138 (N_8138,N_4301,N_2557);
xor U8139 (N_8139,N_1158,N_1542);
or U8140 (N_8140,N_1567,N_3757);
xor U8141 (N_8141,N_1966,N_2031);
or U8142 (N_8142,N_1056,N_780);
nand U8143 (N_8143,N_2351,N_1754);
xnor U8144 (N_8144,N_2408,N_76);
nor U8145 (N_8145,N_1682,N_951);
xnor U8146 (N_8146,N_1763,N_1303);
nand U8147 (N_8147,N_3285,N_3173);
nor U8148 (N_8148,N_4094,N_2595);
or U8149 (N_8149,N_1740,N_4816);
and U8150 (N_8150,N_2748,N_4691);
and U8151 (N_8151,N_610,N_2747);
or U8152 (N_8152,N_3144,N_2245);
nand U8153 (N_8153,N_788,N_4964);
nor U8154 (N_8154,N_1502,N_370);
and U8155 (N_8155,N_3080,N_4185);
and U8156 (N_8156,N_1023,N_4046);
nand U8157 (N_8157,N_3654,N_2772);
and U8158 (N_8158,N_4616,N_1703);
and U8159 (N_8159,N_2504,N_3630);
and U8160 (N_8160,N_1318,N_2891);
xor U8161 (N_8161,N_830,N_309);
nor U8162 (N_8162,N_4054,N_1044);
nor U8163 (N_8163,N_859,N_4507);
or U8164 (N_8164,N_4095,N_158);
xor U8165 (N_8165,N_2924,N_2736);
and U8166 (N_8166,N_211,N_4642);
nand U8167 (N_8167,N_1268,N_1902);
or U8168 (N_8168,N_2969,N_1844);
or U8169 (N_8169,N_4414,N_3997);
nor U8170 (N_8170,N_2013,N_658);
nor U8171 (N_8171,N_2110,N_4428);
and U8172 (N_8172,N_2816,N_3865);
nor U8173 (N_8173,N_1967,N_786);
and U8174 (N_8174,N_4131,N_3364);
xnor U8175 (N_8175,N_4115,N_3409);
or U8176 (N_8176,N_3910,N_3447);
nand U8177 (N_8177,N_739,N_273);
nor U8178 (N_8178,N_630,N_1268);
nor U8179 (N_8179,N_3768,N_1913);
nor U8180 (N_8180,N_4842,N_3432);
or U8181 (N_8181,N_4807,N_4088);
nand U8182 (N_8182,N_3907,N_1741);
or U8183 (N_8183,N_3721,N_2291);
and U8184 (N_8184,N_1425,N_428);
nand U8185 (N_8185,N_3335,N_3047);
nand U8186 (N_8186,N_3487,N_564);
nand U8187 (N_8187,N_3562,N_3230);
nor U8188 (N_8188,N_1295,N_2651);
or U8189 (N_8189,N_3112,N_3946);
and U8190 (N_8190,N_149,N_274);
and U8191 (N_8191,N_2787,N_3104);
and U8192 (N_8192,N_1073,N_1318);
or U8193 (N_8193,N_626,N_1599);
or U8194 (N_8194,N_3591,N_1398);
nand U8195 (N_8195,N_4285,N_2283);
nor U8196 (N_8196,N_2790,N_4188);
and U8197 (N_8197,N_2952,N_4785);
or U8198 (N_8198,N_1605,N_4885);
or U8199 (N_8199,N_3202,N_754);
nor U8200 (N_8200,N_3402,N_3478);
nand U8201 (N_8201,N_840,N_1650);
nor U8202 (N_8202,N_1624,N_4097);
or U8203 (N_8203,N_169,N_4816);
xor U8204 (N_8204,N_2822,N_152);
and U8205 (N_8205,N_4154,N_1084);
or U8206 (N_8206,N_2091,N_1986);
or U8207 (N_8207,N_3403,N_2133);
or U8208 (N_8208,N_4863,N_1819);
and U8209 (N_8209,N_4850,N_785);
nand U8210 (N_8210,N_429,N_2255);
xnor U8211 (N_8211,N_3109,N_1717);
xnor U8212 (N_8212,N_3265,N_2909);
nor U8213 (N_8213,N_3482,N_1602);
and U8214 (N_8214,N_1368,N_761);
or U8215 (N_8215,N_3647,N_4311);
nand U8216 (N_8216,N_3302,N_4264);
nand U8217 (N_8217,N_1132,N_2021);
or U8218 (N_8218,N_537,N_3777);
nor U8219 (N_8219,N_3205,N_2831);
nand U8220 (N_8220,N_3271,N_1075);
nor U8221 (N_8221,N_3305,N_4118);
xnor U8222 (N_8222,N_788,N_3046);
nand U8223 (N_8223,N_2531,N_3163);
or U8224 (N_8224,N_178,N_2248);
or U8225 (N_8225,N_3854,N_1175);
nor U8226 (N_8226,N_3027,N_4560);
or U8227 (N_8227,N_603,N_3815);
xor U8228 (N_8228,N_2744,N_1052);
and U8229 (N_8229,N_59,N_3760);
and U8230 (N_8230,N_320,N_4764);
and U8231 (N_8231,N_4378,N_718);
or U8232 (N_8232,N_3798,N_4955);
or U8233 (N_8233,N_1841,N_701);
nor U8234 (N_8234,N_2666,N_3332);
nand U8235 (N_8235,N_4272,N_2615);
or U8236 (N_8236,N_1569,N_1157);
and U8237 (N_8237,N_1636,N_2715);
nor U8238 (N_8238,N_4651,N_4872);
nor U8239 (N_8239,N_4308,N_2897);
nor U8240 (N_8240,N_12,N_67);
nand U8241 (N_8241,N_2617,N_45);
nor U8242 (N_8242,N_1009,N_3399);
nor U8243 (N_8243,N_3746,N_615);
or U8244 (N_8244,N_1058,N_3450);
nand U8245 (N_8245,N_2581,N_2430);
or U8246 (N_8246,N_4340,N_4958);
or U8247 (N_8247,N_134,N_10);
or U8248 (N_8248,N_4331,N_3307);
or U8249 (N_8249,N_1008,N_2817);
nand U8250 (N_8250,N_3506,N_3865);
and U8251 (N_8251,N_305,N_1440);
and U8252 (N_8252,N_355,N_3283);
nor U8253 (N_8253,N_2305,N_1851);
nor U8254 (N_8254,N_4387,N_400);
nand U8255 (N_8255,N_105,N_4293);
nor U8256 (N_8256,N_2424,N_2789);
nand U8257 (N_8257,N_57,N_4054);
and U8258 (N_8258,N_4740,N_669);
or U8259 (N_8259,N_1322,N_2178);
or U8260 (N_8260,N_1790,N_2512);
nor U8261 (N_8261,N_1483,N_2158);
and U8262 (N_8262,N_3545,N_3919);
nand U8263 (N_8263,N_2222,N_1361);
nand U8264 (N_8264,N_2321,N_3661);
or U8265 (N_8265,N_3320,N_2068);
and U8266 (N_8266,N_4205,N_772);
nand U8267 (N_8267,N_3142,N_3252);
nor U8268 (N_8268,N_4188,N_4776);
and U8269 (N_8269,N_1318,N_1124);
or U8270 (N_8270,N_3280,N_1706);
and U8271 (N_8271,N_3330,N_1155);
or U8272 (N_8272,N_1911,N_4368);
nand U8273 (N_8273,N_4935,N_1965);
xor U8274 (N_8274,N_137,N_1475);
and U8275 (N_8275,N_1323,N_999);
or U8276 (N_8276,N_168,N_2778);
xnor U8277 (N_8277,N_3831,N_3961);
xor U8278 (N_8278,N_1339,N_2955);
nand U8279 (N_8279,N_1959,N_3275);
or U8280 (N_8280,N_3272,N_969);
nand U8281 (N_8281,N_2475,N_261);
and U8282 (N_8282,N_2525,N_3685);
nand U8283 (N_8283,N_386,N_457);
or U8284 (N_8284,N_2868,N_3680);
and U8285 (N_8285,N_3154,N_2199);
xor U8286 (N_8286,N_3069,N_1062);
nor U8287 (N_8287,N_75,N_4457);
and U8288 (N_8288,N_1164,N_3568);
nor U8289 (N_8289,N_2471,N_1622);
or U8290 (N_8290,N_2721,N_2521);
nand U8291 (N_8291,N_1438,N_4519);
nand U8292 (N_8292,N_3799,N_1706);
and U8293 (N_8293,N_4743,N_286);
nor U8294 (N_8294,N_4634,N_1782);
nand U8295 (N_8295,N_1395,N_4151);
nand U8296 (N_8296,N_2612,N_4683);
nor U8297 (N_8297,N_1940,N_964);
and U8298 (N_8298,N_4030,N_2089);
or U8299 (N_8299,N_1062,N_669);
nor U8300 (N_8300,N_3672,N_2324);
or U8301 (N_8301,N_4088,N_2354);
nor U8302 (N_8302,N_1009,N_4974);
and U8303 (N_8303,N_1543,N_922);
nand U8304 (N_8304,N_4853,N_2461);
nor U8305 (N_8305,N_76,N_2959);
nor U8306 (N_8306,N_1491,N_4100);
nand U8307 (N_8307,N_4706,N_3719);
and U8308 (N_8308,N_3269,N_1569);
nor U8309 (N_8309,N_3854,N_4551);
and U8310 (N_8310,N_3748,N_1193);
nor U8311 (N_8311,N_893,N_4303);
or U8312 (N_8312,N_4119,N_4711);
nand U8313 (N_8313,N_1143,N_4263);
nor U8314 (N_8314,N_4227,N_3455);
or U8315 (N_8315,N_974,N_3213);
nand U8316 (N_8316,N_3674,N_1480);
nand U8317 (N_8317,N_1025,N_3576);
nor U8318 (N_8318,N_4316,N_3568);
nor U8319 (N_8319,N_2330,N_3825);
or U8320 (N_8320,N_3810,N_2419);
nor U8321 (N_8321,N_340,N_418);
nand U8322 (N_8322,N_299,N_451);
nor U8323 (N_8323,N_4484,N_2418);
and U8324 (N_8324,N_2656,N_4030);
or U8325 (N_8325,N_4205,N_1544);
nor U8326 (N_8326,N_3276,N_4817);
or U8327 (N_8327,N_2446,N_2349);
and U8328 (N_8328,N_77,N_973);
or U8329 (N_8329,N_3031,N_1729);
nand U8330 (N_8330,N_1312,N_774);
nor U8331 (N_8331,N_3725,N_1650);
and U8332 (N_8332,N_3683,N_1967);
and U8333 (N_8333,N_2895,N_4931);
nand U8334 (N_8334,N_2084,N_4269);
nor U8335 (N_8335,N_1240,N_1011);
and U8336 (N_8336,N_1009,N_4408);
and U8337 (N_8337,N_3183,N_1971);
nor U8338 (N_8338,N_1300,N_803);
or U8339 (N_8339,N_3527,N_2287);
or U8340 (N_8340,N_3059,N_4157);
and U8341 (N_8341,N_1539,N_3859);
or U8342 (N_8342,N_4815,N_4476);
nand U8343 (N_8343,N_837,N_4670);
or U8344 (N_8344,N_302,N_4179);
nand U8345 (N_8345,N_3321,N_3650);
nand U8346 (N_8346,N_299,N_2150);
xnor U8347 (N_8347,N_2813,N_453);
and U8348 (N_8348,N_1116,N_2646);
nor U8349 (N_8349,N_977,N_661);
xnor U8350 (N_8350,N_2296,N_2814);
and U8351 (N_8351,N_1733,N_3407);
xnor U8352 (N_8352,N_4626,N_576);
or U8353 (N_8353,N_3297,N_2418);
and U8354 (N_8354,N_3258,N_4000);
and U8355 (N_8355,N_1299,N_219);
and U8356 (N_8356,N_4109,N_1831);
and U8357 (N_8357,N_789,N_2118);
and U8358 (N_8358,N_1222,N_4202);
nor U8359 (N_8359,N_1276,N_2454);
nand U8360 (N_8360,N_2484,N_4909);
or U8361 (N_8361,N_4369,N_199);
or U8362 (N_8362,N_1192,N_2986);
nand U8363 (N_8363,N_2677,N_889);
and U8364 (N_8364,N_4200,N_2007);
nor U8365 (N_8365,N_2712,N_4385);
and U8366 (N_8366,N_503,N_4723);
nor U8367 (N_8367,N_292,N_4851);
nor U8368 (N_8368,N_561,N_220);
nor U8369 (N_8369,N_1801,N_531);
nand U8370 (N_8370,N_2319,N_2763);
nand U8371 (N_8371,N_3360,N_1750);
or U8372 (N_8372,N_3542,N_3530);
and U8373 (N_8373,N_1759,N_2516);
nor U8374 (N_8374,N_1309,N_992);
and U8375 (N_8375,N_1658,N_475);
and U8376 (N_8376,N_3710,N_3041);
nor U8377 (N_8377,N_3413,N_2912);
or U8378 (N_8378,N_4990,N_2893);
xor U8379 (N_8379,N_992,N_3600);
nor U8380 (N_8380,N_3858,N_4964);
and U8381 (N_8381,N_1812,N_1676);
nor U8382 (N_8382,N_174,N_2556);
and U8383 (N_8383,N_1701,N_1603);
or U8384 (N_8384,N_2475,N_3949);
nor U8385 (N_8385,N_2157,N_3455);
or U8386 (N_8386,N_1936,N_4052);
or U8387 (N_8387,N_1352,N_1287);
and U8388 (N_8388,N_4525,N_2998);
or U8389 (N_8389,N_4249,N_2665);
or U8390 (N_8390,N_3997,N_107);
xnor U8391 (N_8391,N_624,N_359);
nor U8392 (N_8392,N_2042,N_3706);
and U8393 (N_8393,N_3289,N_3073);
nand U8394 (N_8394,N_3873,N_4530);
or U8395 (N_8395,N_3960,N_3137);
or U8396 (N_8396,N_2053,N_2598);
and U8397 (N_8397,N_704,N_1739);
and U8398 (N_8398,N_2613,N_2351);
nor U8399 (N_8399,N_1186,N_4769);
nor U8400 (N_8400,N_1924,N_4793);
nor U8401 (N_8401,N_4910,N_2054);
nor U8402 (N_8402,N_1812,N_1618);
and U8403 (N_8403,N_3570,N_144);
and U8404 (N_8404,N_3719,N_2763);
and U8405 (N_8405,N_4660,N_1217);
or U8406 (N_8406,N_3809,N_3173);
nand U8407 (N_8407,N_3988,N_4727);
or U8408 (N_8408,N_4174,N_4656);
and U8409 (N_8409,N_2433,N_1050);
and U8410 (N_8410,N_3608,N_1142);
xnor U8411 (N_8411,N_2775,N_2522);
or U8412 (N_8412,N_4227,N_1434);
or U8413 (N_8413,N_3191,N_521);
nor U8414 (N_8414,N_4868,N_1086);
nor U8415 (N_8415,N_2793,N_4887);
or U8416 (N_8416,N_4089,N_3289);
and U8417 (N_8417,N_323,N_170);
or U8418 (N_8418,N_3841,N_3663);
nor U8419 (N_8419,N_2968,N_3637);
nand U8420 (N_8420,N_3534,N_3049);
and U8421 (N_8421,N_2461,N_974);
or U8422 (N_8422,N_1945,N_1707);
nand U8423 (N_8423,N_454,N_546);
or U8424 (N_8424,N_2510,N_4076);
nor U8425 (N_8425,N_2536,N_1376);
xnor U8426 (N_8426,N_3622,N_3308);
nand U8427 (N_8427,N_1055,N_4894);
or U8428 (N_8428,N_1090,N_3219);
nand U8429 (N_8429,N_1318,N_744);
xnor U8430 (N_8430,N_1705,N_3959);
nor U8431 (N_8431,N_837,N_1757);
nor U8432 (N_8432,N_4635,N_3484);
nand U8433 (N_8433,N_4435,N_4958);
or U8434 (N_8434,N_1492,N_2313);
nand U8435 (N_8435,N_2012,N_711);
nor U8436 (N_8436,N_2976,N_3242);
or U8437 (N_8437,N_4876,N_4029);
and U8438 (N_8438,N_1519,N_2786);
or U8439 (N_8439,N_2762,N_3255);
nand U8440 (N_8440,N_3307,N_322);
or U8441 (N_8441,N_3725,N_4527);
or U8442 (N_8442,N_1496,N_3477);
and U8443 (N_8443,N_62,N_909);
nand U8444 (N_8444,N_1522,N_3477);
or U8445 (N_8445,N_257,N_2615);
nand U8446 (N_8446,N_1782,N_4503);
or U8447 (N_8447,N_3234,N_39);
and U8448 (N_8448,N_671,N_3254);
and U8449 (N_8449,N_93,N_4533);
nor U8450 (N_8450,N_4273,N_942);
nor U8451 (N_8451,N_4217,N_3184);
and U8452 (N_8452,N_1158,N_1791);
or U8453 (N_8453,N_4341,N_4674);
or U8454 (N_8454,N_2753,N_3172);
xnor U8455 (N_8455,N_2948,N_2228);
nor U8456 (N_8456,N_4658,N_2453);
or U8457 (N_8457,N_4630,N_1625);
or U8458 (N_8458,N_4229,N_345);
nand U8459 (N_8459,N_2235,N_4075);
nand U8460 (N_8460,N_1772,N_4845);
nand U8461 (N_8461,N_2355,N_3299);
nand U8462 (N_8462,N_785,N_3118);
nor U8463 (N_8463,N_483,N_3586);
nand U8464 (N_8464,N_740,N_2042);
and U8465 (N_8465,N_2927,N_2458);
nand U8466 (N_8466,N_1896,N_4895);
and U8467 (N_8467,N_3937,N_3753);
and U8468 (N_8468,N_2716,N_2786);
xor U8469 (N_8469,N_395,N_2067);
nor U8470 (N_8470,N_137,N_2795);
or U8471 (N_8471,N_2237,N_562);
or U8472 (N_8472,N_1333,N_259);
xor U8473 (N_8473,N_1210,N_1665);
and U8474 (N_8474,N_3767,N_1069);
or U8475 (N_8475,N_1612,N_4944);
or U8476 (N_8476,N_1113,N_2423);
nor U8477 (N_8477,N_4777,N_478);
and U8478 (N_8478,N_3541,N_1263);
or U8479 (N_8479,N_3249,N_106);
or U8480 (N_8480,N_927,N_4093);
or U8481 (N_8481,N_1146,N_3966);
and U8482 (N_8482,N_4470,N_2952);
or U8483 (N_8483,N_4488,N_1982);
or U8484 (N_8484,N_3648,N_2455);
or U8485 (N_8485,N_4830,N_4164);
and U8486 (N_8486,N_1684,N_1650);
nand U8487 (N_8487,N_1575,N_3236);
or U8488 (N_8488,N_835,N_4802);
nand U8489 (N_8489,N_4809,N_4814);
nor U8490 (N_8490,N_2715,N_1941);
nor U8491 (N_8491,N_4272,N_590);
or U8492 (N_8492,N_800,N_1179);
xnor U8493 (N_8493,N_357,N_3667);
or U8494 (N_8494,N_4853,N_3593);
or U8495 (N_8495,N_3182,N_3303);
nor U8496 (N_8496,N_1547,N_3598);
nor U8497 (N_8497,N_4406,N_2979);
nor U8498 (N_8498,N_2502,N_4790);
xnor U8499 (N_8499,N_4512,N_4999);
nand U8500 (N_8500,N_3357,N_718);
nand U8501 (N_8501,N_2518,N_2833);
or U8502 (N_8502,N_2643,N_368);
or U8503 (N_8503,N_3436,N_1520);
nor U8504 (N_8504,N_3221,N_2904);
nor U8505 (N_8505,N_61,N_1358);
nor U8506 (N_8506,N_1362,N_1147);
and U8507 (N_8507,N_4030,N_3798);
nand U8508 (N_8508,N_4354,N_2784);
nor U8509 (N_8509,N_1984,N_169);
and U8510 (N_8510,N_2690,N_286);
nand U8511 (N_8511,N_4614,N_1771);
and U8512 (N_8512,N_2230,N_4604);
or U8513 (N_8513,N_1618,N_1090);
or U8514 (N_8514,N_521,N_1691);
or U8515 (N_8515,N_4246,N_989);
nand U8516 (N_8516,N_1874,N_1);
nand U8517 (N_8517,N_3902,N_3856);
and U8518 (N_8518,N_1099,N_4268);
nand U8519 (N_8519,N_4635,N_1027);
or U8520 (N_8520,N_4237,N_69);
or U8521 (N_8521,N_1955,N_2065);
nand U8522 (N_8522,N_4833,N_1305);
nor U8523 (N_8523,N_3882,N_4165);
and U8524 (N_8524,N_984,N_4702);
nor U8525 (N_8525,N_4227,N_1118);
or U8526 (N_8526,N_4751,N_1138);
nor U8527 (N_8527,N_3554,N_2818);
or U8528 (N_8528,N_4617,N_1968);
nor U8529 (N_8529,N_1264,N_1230);
nand U8530 (N_8530,N_3268,N_2179);
nor U8531 (N_8531,N_2350,N_1729);
nor U8532 (N_8532,N_3160,N_529);
and U8533 (N_8533,N_626,N_972);
and U8534 (N_8534,N_4473,N_808);
or U8535 (N_8535,N_2061,N_944);
nand U8536 (N_8536,N_2195,N_229);
nor U8537 (N_8537,N_4117,N_2761);
nor U8538 (N_8538,N_1532,N_2961);
xnor U8539 (N_8539,N_2099,N_4860);
nor U8540 (N_8540,N_4672,N_4515);
nand U8541 (N_8541,N_2164,N_424);
nand U8542 (N_8542,N_1658,N_1096);
or U8543 (N_8543,N_1870,N_2602);
nor U8544 (N_8544,N_4968,N_1028);
and U8545 (N_8545,N_724,N_487);
nor U8546 (N_8546,N_3793,N_1932);
nor U8547 (N_8547,N_3834,N_1058);
and U8548 (N_8548,N_2431,N_3047);
or U8549 (N_8549,N_1308,N_4822);
and U8550 (N_8550,N_4541,N_2084);
nor U8551 (N_8551,N_179,N_3533);
or U8552 (N_8552,N_2521,N_2414);
or U8553 (N_8553,N_2259,N_1809);
nand U8554 (N_8554,N_4772,N_2750);
nor U8555 (N_8555,N_4149,N_517);
or U8556 (N_8556,N_423,N_2496);
and U8557 (N_8557,N_3787,N_2217);
nand U8558 (N_8558,N_109,N_4185);
or U8559 (N_8559,N_687,N_1017);
nand U8560 (N_8560,N_2839,N_3327);
and U8561 (N_8561,N_93,N_3726);
nor U8562 (N_8562,N_3379,N_2188);
nor U8563 (N_8563,N_4042,N_1827);
nand U8564 (N_8564,N_4855,N_2009);
nor U8565 (N_8565,N_4172,N_1989);
xor U8566 (N_8566,N_430,N_4229);
nand U8567 (N_8567,N_3870,N_4728);
and U8568 (N_8568,N_3088,N_1182);
and U8569 (N_8569,N_2211,N_4710);
xnor U8570 (N_8570,N_2225,N_2232);
or U8571 (N_8571,N_531,N_2726);
or U8572 (N_8572,N_378,N_3067);
or U8573 (N_8573,N_2715,N_1291);
nor U8574 (N_8574,N_1131,N_800);
and U8575 (N_8575,N_839,N_3460);
and U8576 (N_8576,N_2314,N_2788);
nor U8577 (N_8577,N_1720,N_1665);
nor U8578 (N_8578,N_4523,N_1598);
or U8579 (N_8579,N_4138,N_3692);
xnor U8580 (N_8580,N_817,N_4831);
or U8581 (N_8581,N_1409,N_3748);
and U8582 (N_8582,N_2136,N_2433);
nand U8583 (N_8583,N_1455,N_4307);
nor U8584 (N_8584,N_3380,N_1943);
and U8585 (N_8585,N_54,N_2762);
or U8586 (N_8586,N_3138,N_1809);
nor U8587 (N_8587,N_3271,N_2465);
nor U8588 (N_8588,N_769,N_2808);
xor U8589 (N_8589,N_1731,N_2310);
or U8590 (N_8590,N_3995,N_687);
or U8591 (N_8591,N_2111,N_366);
xor U8592 (N_8592,N_777,N_4543);
nor U8593 (N_8593,N_1401,N_3347);
nand U8594 (N_8594,N_827,N_2707);
nor U8595 (N_8595,N_2305,N_1554);
and U8596 (N_8596,N_1024,N_1760);
and U8597 (N_8597,N_3316,N_4093);
or U8598 (N_8598,N_377,N_994);
or U8599 (N_8599,N_3302,N_93);
nand U8600 (N_8600,N_370,N_4707);
nor U8601 (N_8601,N_4068,N_1727);
nand U8602 (N_8602,N_1770,N_1592);
and U8603 (N_8603,N_70,N_3168);
nand U8604 (N_8604,N_322,N_1103);
or U8605 (N_8605,N_1793,N_1932);
or U8606 (N_8606,N_1116,N_95);
or U8607 (N_8607,N_4447,N_3279);
nand U8608 (N_8608,N_4507,N_3279);
xnor U8609 (N_8609,N_4680,N_2397);
and U8610 (N_8610,N_608,N_2050);
nor U8611 (N_8611,N_2051,N_2214);
or U8612 (N_8612,N_1317,N_3326);
nand U8613 (N_8613,N_4118,N_2052);
or U8614 (N_8614,N_268,N_1837);
nand U8615 (N_8615,N_3164,N_2574);
or U8616 (N_8616,N_1210,N_2632);
or U8617 (N_8617,N_2285,N_3005);
and U8618 (N_8618,N_343,N_2038);
nor U8619 (N_8619,N_2846,N_1022);
nand U8620 (N_8620,N_3079,N_4807);
xor U8621 (N_8621,N_4707,N_990);
nand U8622 (N_8622,N_4240,N_3216);
and U8623 (N_8623,N_1244,N_3399);
nor U8624 (N_8624,N_3529,N_2122);
or U8625 (N_8625,N_3525,N_2085);
and U8626 (N_8626,N_2569,N_1856);
nand U8627 (N_8627,N_3805,N_955);
and U8628 (N_8628,N_2127,N_2463);
nand U8629 (N_8629,N_3216,N_2026);
nand U8630 (N_8630,N_418,N_3858);
nand U8631 (N_8631,N_167,N_2965);
xnor U8632 (N_8632,N_3896,N_4741);
or U8633 (N_8633,N_343,N_829);
nand U8634 (N_8634,N_1629,N_385);
nor U8635 (N_8635,N_3755,N_2686);
nor U8636 (N_8636,N_4226,N_2035);
nor U8637 (N_8637,N_3115,N_504);
nand U8638 (N_8638,N_1671,N_2951);
nand U8639 (N_8639,N_1648,N_80);
or U8640 (N_8640,N_391,N_3151);
nand U8641 (N_8641,N_318,N_581);
nor U8642 (N_8642,N_392,N_2750);
nand U8643 (N_8643,N_2026,N_1481);
nor U8644 (N_8644,N_4668,N_4390);
and U8645 (N_8645,N_4923,N_4548);
or U8646 (N_8646,N_2360,N_1832);
or U8647 (N_8647,N_241,N_3286);
and U8648 (N_8648,N_457,N_2491);
nand U8649 (N_8649,N_4800,N_4378);
and U8650 (N_8650,N_4974,N_1786);
xor U8651 (N_8651,N_2272,N_490);
nor U8652 (N_8652,N_460,N_3783);
nor U8653 (N_8653,N_4606,N_2395);
and U8654 (N_8654,N_209,N_4388);
nor U8655 (N_8655,N_4889,N_462);
or U8656 (N_8656,N_3448,N_3887);
nor U8657 (N_8657,N_4955,N_4597);
nor U8658 (N_8658,N_3468,N_1093);
nor U8659 (N_8659,N_2687,N_3358);
xor U8660 (N_8660,N_3185,N_2014);
or U8661 (N_8661,N_2451,N_2432);
nor U8662 (N_8662,N_17,N_3071);
and U8663 (N_8663,N_1334,N_1469);
and U8664 (N_8664,N_602,N_504);
or U8665 (N_8665,N_2567,N_1379);
nand U8666 (N_8666,N_2614,N_672);
and U8667 (N_8667,N_4993,N_3812);
nand U8668 (N_8668,N_1792,N_2692);
and U8669 (N_8669,N_2156,N_4769);
xor U8670 (N_8670,N_21,N_2195);
nand U8671 (N_8671,N_1346,N_674);
xor U8672 (N_8672,N_4910,N_1250);
nand U8673 (N_8673,N_4849,N_4377);
nor U8674 (N_8674,N_421,N_2061);
nand U8675 (N_8675,N_661,N_930);
nor U8676 (N_8676,N_1293,N_3531);
or U8677 (N_8677,N_3483,N_1008);
nor U8678 (N_8678,N_4698,N_4848);
nor U8679 (N_8679,N_3535,N_2101);
and U8680 (N_8680,N_31,N_2733);
nor U8681 (N_8681,N_3813,N_2094);
or U8682 (N_8682,N_65,N_3033);
or U8683 (N_8683,N_1258,N_3719);
nand U8684 (N_8684,N_902,N_158);
nand U8685 (N_8685,N_4197,N_3607);
and U8686 (N_8686,N_2096,N_4405);
or U8687 (N_8687,N_2844,N_4673);
xnor U8688 (N_8688,N_1691,N_3130);
nor U8689 (N_8689,N_3432,N_2013);
or U8690 (N_8690,N_929,N_481);
nand U8691 (N_8691,N_4560,N_2301);
nand U8692 (N_8692,N_2261,N_4576);
and U8693 (N_8693,N_1320,N_2813);
or U8694 (N_8694,N_1272,N_3096);
or U8695 (N_8695,N_1588,N_93);
nor U8696 (N_8696,N_1370,N_4652);
or U8697 (N_8697,N_822,N_1536);
nor U8698 (N_8698,N_1334,N_1489);
or U8699 (N_8699,N_3245,N_2881);
nand U8700 (N_8700,N_1478,N_4777);
or U8701 (N_8701,N_3695,N_4136);
nor U8702 (N_8702,N_612,N_1153);
nor U8703 (N_8703,N_2048,N_2329);
nand U8704 (N_8704,N_1020,N_2464);
or U8705 (N_8705,N_267,N_4814);
nand U8706 (N_8706,N_2868,N_2779);
and U8707 (N_8707,N_3740,N_38);
nor U8708 (N_8708,N_4970,N_1386);
and U8709 (N_8709,N_1767,N_517);
nor U8710 (N_8710,N_3389,N_214);
xor U8711 (N_8711,N_2015,N_376);
or U8712 (N_8712,N_3276,N_3561);
nor U8713 (N_8713,N_4982,N_4014);
and U8714 (N_8714,N_3284,N_260);
nand U8715 (N_8715,N_2983,N_1629);
and U8716 (N_8716,N_3292,N_4233);
nand U8717 (N_8717,N_1595,N_679);
nor U8718 (N_8718,N_320,N_1684);
or U8719 (N_8719,N_4672,N_1241);
or U8720 (N_8720,N_254,N_2375);
xor U8721 (N_8721,N_2185,N_1728);
xnor U8722 (N_8722,N_1787,N_4368);
nor U8723 (N_8723,N_1702,N_775);
nand U8724 (N_8724,N_1488,N_2510);
or U8725 (N_8725,N_2197,N_1241);
and U8726 (N_8726,N_939,N_4696);
nand U8727 (N_8727,N_266,N_4425);
nor U8728 (N_8728,N_3266,N_4962);
nor U8729 (N_8729,N_3932,N_795);
nor U8730 (N_8730,N_1398,N_315);
or U8731 (N_8731,N_2805,N_3147);
and U8732 (N_8732,N_4658,N_2326);
nor U8733 (N_8733,N_3029,N_2874);
nand U8734 (N_8734,N_3600,N_3395);
xor U8735 (N_8735,N_1905,N_4958);
nand U8736 (N_8736,N_4155,N_4434);
and U8737 (N_8737,N_4245,N_134);
nand U8738 (N_8738,N_4041,N_362);
nand U8739 (N_8739,N_74,N_2249);
and U8740 (N_8740,N_3336,N_4484);
nand U8741 (N_8741,N_2165,N_1354);
nand U8742 (N_8742,N_2872,N_1154);
nor U8743 (N_8743,N_3361,N_2349);
nand U8744 (N_8744,N_4808,N_4402);
and U8745 (N_8745,N_1050,N_4824);
nor U8746 (N_8746,N_3859,N_4795);
nor U8747 (N_8747,N_1297,N_482);
xnor U8748 (N_8748,N_2718,N_4940);
nor U8749 (N_8749,N_2941,N_1160);
and U8750 (N_8750,N_2730,N_2502);
nor U8751 (N_8751,N_2924,N_3809);
nand U8752 (N_8752,N_1218,N_1659);
and U8753 (N_8753,N_1838,N_4042);
nor U8754 (N_8754,N_1015,N_3185);
nand U8755 (N_8755,N_4752,N_1398);
and U8756 (N_8756,N_3108,N_2311);
nand U8757 (N_8757,N_2406,N_795);
nor U8758 (N_8758,N_2698,N_2659);
and U8759 (N_8759,N_3069,N_1012);
nor U8760 (N_8760,N_4020,N_2031);
and U8761 (N_8761,N_4051,N_1740);
xor U8762 (N_8762,N_322,N_2374);
nor U8763 (N_8763,N_4408,N_957);
and U8764 (N_8764,N_2618,N_1373);
nor U8765 (N_8765,N_2973,N_1783);
nand U8766 (N_8766,N_4569,N_2123);
nor U8767 (N_8767,N_986,N_1450);
nor U8768 (N_8768,N_1250,N_2483);
nand U8769 (N_8769,N_417,N_2712);
xnor U8770 (N_8770,N_3508,N_1671);
and U8771 (N_8771,N_1283,N_4520);
nor U8772 (N_8772,N_4102,N_4267);
and U8773 (N_8773,N_2507,N_2256);
nor U8774 (N_8774,N_1465,N_4930);
xnor U8775 (N_8775,N_3123,N_2232);
nand U8776 (N_8776,N_2284,N_4078);
nand U8777 (N_8777,N_3340,N_1519);
or U8778 (N_8778,N_751,N_3962);
and U8779 (N_8779,N_3976,N_1519);
nand U8780 (N_8780,N_1018,N_4145);
nor U8781 (N_8781,N_819,N_2612);
nor U8782 (N_8782,N_2197,N_3194);
or U8783 (N_8783,N_3488,N_4658);
nand U8784 (N_8784,N_3969,N_910);
nand U8785 (N_8785,N_921,N_84);
nand U8786 (N_8786,N_2164,N_4253);
and U8787 (N_8787,N_679,N_1635);
nor U8788 (N_8788,N_2874,N_3210);
nor U8789 (N_8789,N_2062,N_1714);
nor U8790 (N_8790,N_4388,N_249);
nand U8791 (N_8791,N_2891,N_3011);
or U8792 (N_8792,N_4798,N_1447);
nor U8793 (N_8793,N_798,N_2504);
nand U8794 (N_8794,N_1408,N_4649);
or U8795 (N_8795,N_2839,N_4272);
and U8796 (N_8796,N_4558,N_81);
and U8797 (N_8797,N_2599,N_4348);
and U8798 (N_8798,N_2064,N_2349);
xnor U8799 (N_8799,N_3301,N_2602);
nand U8800 (N_8800,N_2414,N_4668);
nor U8801 (N_8801,N_3166,N_3646);
and U8802 (N_8802,N_1518,N_1651);
and U8803 (N_8803,N_4590,N_4713);
nor U8804 (N_8804,N_575,N_1928);
xor U8805 (N_8805,N_4223,N_1172);
and U8806 (N_8806,N_4612,N_1568);
or U8807 (N_8807,N_806,N_1943);
or U8808 (N_8808,N_2187,N_3589);
nor U8809 (N_8809,N_4380,N_3174);
nand U8810 (N_8810,N_4100,N_877);
nor U8811 (N_8811,N_1529,N_2164);
xnor U8812 (N_8812,N_618,N_2888);
nand U8813 (N_8813,N_2249,N_29);
nand U8814 (N_8814,N_3190,N_3569);
nor U8815 (N_8815,N_3304,N_2471);
and U8816 (N_8816,N_2563,N_966);
nor U8817 (N_8817,N_3214,N_410);
and U8818 (N_8818,N_3691,N_4272);
and U8819 (N_8819,N_1440,N_379);
or U8820 (N_8820,N_1337,N_2264);
nor U8821 (N_8821,N_4819,N_1060);
and U8822 (N_8822,N_4974,N_2803);
nand U8823 (N_8823,N_835,N_4365);
nand U8824 (N_8824,N_739,N_545);
nand U8825 (N_8825,N_3632,N_724);
nand U8826 (N_8826,N_97,N_2582);
and U8827 (N_8827,N_291,N_2513);
nor U8828 (N_8828,N_1129,N_4794);
nand U8829 (N_8829,N_306,N_90);
nand U8830 (N_8830,N_2975,N_920);
nor U8831 (N_8831,N_263,N_1384);
and U8832 (N_8832,N_2960,N_324);
and U8833 (N_8833,N_309,N_1822);
nand U8834 (N_8834,N_868,N_3389);
xnor U8835 (N_8835,N_1883,N_3454);
nand U8836 (N_8836,N_2997,N_2345);
xor U8837 (N_8837,N_2748,N_4134);
xnor U8838 (N_8838,N_4937,N_232);
xnor U8839 (N_8839,N_2812,N_2954);
or U8840 (N_8840,N_4907,N_605);
nand U8841 (N_8841,N_1825,N_2824);
nand U8842 (N_8842,N_1251,N_1605);
nand U8843 (N_8843,N_265,N_1042);
nor U8844 (N_8844,N_3737,N_563);
nor U8845 (N_8845,N_191,N_4730);
nand U8846 (N_8846,N_3742,N_2533);
xnor U8847 (N_8847,N_1773,N_1276);
xnor U8848 (N_8848,N_1828,N_2708);
and U8849 (N_8849,N_1147,N_2837);
or U8850 (N_8850,N_3782,N_999);
nand U8851 (N_8851,N_2601,N_109);
and U8852 (N_8852,N_3162,N_1066);
xor U8853 (N_8853,N_2310,N_4686);
nor U8854 (N_8854,N_2694,N_3773);
and U8855 (N_8855,N_2909,N_625);
and U8856 (N_8856,N_2695,N_31);
xor U8857 (N_8857,N_3049,N_559);
or U8858 (N_8858,N_2156,N_4734);
and U8859 (N_8859,N_783,N_3811);
nand U8860 (N_8860,N_204,N_2189);
xnor U8861 (N_8861,N_4470,N_1149);
or U8862 (N_8862,N_2332,N_2640);
or U8863 (N_8863,N_2915,N_3637);
nand U8864 (N_8864,N_3503,N_2686);
xor U8865 (N_8865,N_747,N_2486);
nor U8866 (N_8866,N_104,N_3086);
xor U8867 (N_8867,N_4593,N_4905);
nand U8868 (N_8868,N_4766,N_334);
and U8869 (N_8869,N_1839,N_3801);
nand U8870 (N_8870,N_939,N_1243);
xor U8871 (N_8871,N_4349,N_4946);
or U8872 (N_8872,N_4039,N_2958);
or U8873 (N_8873,N_3530,N_3415);
nand U8874 (N_8874,N_1331,N_3932);
and U8875 (N_8875,N_2184,N_3624);
nor U8876 (N_8876,N_821,N_883);
or U8877 (N_8877,N_3657,N_1742);
nor U8878 (N_8878,N_1319,N_288);
nor U8879 (N_8879,N_2075,N_3262);
nand U8880 (N_8880,N_2769,N_3271);
or U8881 (N_8881,N_344,N_2971);
or U8882 (N_8882,N_3255,N_2905);
and U8883 (N_8883,N_3573,N_2660);
and U8884 (N_8884,N_4227,N_1162);
or U8885 (N_8885,N_658,N_650);
and U8886 (N_8886,N_124,N_2989);
and U8887 (N_8887,N_4193,N_2864);
nand U8888 (N_8888,N_132,N_3833);
and U8889 (N_8889,N_1565,N_2534);
and U8890 (N_8890,N_1649,N_4818);
nor U8891 (N_8891,N_1014,N_962);
or U8892 (N_8892,N_3216,N_4829);
and U8893 (N_8893,N_2436,N_1241);
nand U8894 (N_8894,N_4572,N_955);
nor U8895 (N_8895,N_1199,N_3401);
and U8896 (N_8896,N_45,N_4007);
nand U8897 (N_8897,N_2025,N_4915);
nor U8898 (N_8898,N_4955,N_77);
or U8899 (N_8899,N_3749,N_2697);
or U8900 (N_8900,N_3594,N_3286);
nor U8901 (N_8901,N_4552,N_4218);
and U8902 (N_8902,N_2339,N_2367);
and U8903 (N_8903,N_979,N_3086);
and U8904 (N_8904,N_202,N_1489);
or U8905 (N_8905,N_2517,N_3168);
or U8906 (N_8906,N_1209,N_2374);
nor U8907 (N_8907,N_846,N_2843);
and U8908 (N_8908,N_2799,N_335);
and U8909 (N_8909,N_760,N_63);
nand U8910 (N_8910,N_2064,N_332);
xnor U8911 (N_8911,N_3747,N_640);
or U8912 (N_8912,N_293,N_2778);
and U8913 (N_8913,N_2559,N_1459);
or U8914 (N_8914,N_3849,N_4255);
nand U8915 (N_8915,N_469,N_862);
or U8916 (N_8916,N_2261,N_426);
xnor U8917 (N_8917,N_1462,N_4978);
xor U8918 (N_8918,N_3718,N_1558);
nor U8919 (N_8919,N_138,N_2283);
xnor U8920 (N_8920,N_1490,N_53);
and U8921 (N_8921,N_4060,N_665);
nor U8922 (N_8922,N_634,N_643);
nor U8923 (N_8923,N_4796,N_3133);
nor U8924 (N_8924,N_55,N_291);
or U8925 (N_8925,N_2159,N_2478);
or U8926 (N_8926,N_2794,N_3612);
nand U8927 (N_8927,N_3796,N_2311);
nand U8928 (N_8928,N_4384,N_2129);
or U8929 (N_8929,N_2952,N_1674);
and U8930 (N_8930,N_1334,N_2263);
or U8931 (N_8931,N_4287,N_4339);
xnor U8932 (N_8932,N_3630,N_260);
or U8933 (N_8933,N_3708,N_799);
nor U8934 (N_8934,N_1406,N_2172);
or U8935 (N_8935,N_3659,N_37);
nand U8936 (N_8936,N_3130,N_200);
nor U8937 (N_8937,N_1077,N_4443);
and U8938 (N_8938,N_684,N_3806);
nand U8939 (N_8939,N_1103,N_1046);
or U8940 (N_8940,N_745,N_3327);
nand U8941 (N_8941,N_188,N_1505);
or U8942 (N_8942,N_2016,N_3201);
nand U8943 (N_8943,N_4072,N_4599);
or U8944 (N_8944,N_742,N_700);
and U8945 (N_8945,N_3757,N_287);
nor U8946 (N_8946,N_566,N_4957);
and U8947 (N_8947,N_3777,N_2823);
and U8948 (N_8948,N_3368,N_1394);
nand U8949 (N_8949,N_246,N_2922);
or U8950 (N_8950,N_1550,N_4113);
xor U8951 (N_8951,N_4800,N_2774);
or U8952 (N_8952,N_4717,N_3472);
nor U8953 (N_8953,N_908,N_714);
or U8954 (N_8954,N_2401,N_1634);
or U8955 (N_8955,N_2665,N_13);
nor U8956 (N_8956,N_862,N_953);
or U8957 (N_8957,N_514,N_2078);
or U8958 (N_8958,N_1977,N_317);
nor U8959 (N_8959,N_2813,N_4793);
and U8960 (N_8960,N_570,N_3214);
nor U8961 (N_8961,N_2623,N_1243);
nor U8962 (N_8962,N_3201,N_2433);
and U8963 (N_8963,N_3661,N_1997);
nor U8964 (N_8964,N_2486,N_2522);
xor U8965 (N_8965,N_2460,N_4564);
and U8966 (N_8966,N_821,N_1546);
and U8967 (N_8967,N_2028,N_3671);
nor U8968 (N_8968,N_3909,N_1466);
nand U8969 (N_8969,N_2440,N_11);
xnor U8970 (N_8970,N_2043,N_2312);
and U8971 (N_8971,N_3074,N_4553);
xor U8972 (N_8972,N_4449,N_4122);
nor U8973 (N_8973,N_3583,N_1);
or U8974 (N_8974,N_1249,N_2248);
and U8975 (N_8975,N_840,N_878);
or U8976 (N_8976,N_4007,N_4861);
nand U8977 (N_8977,N_3770,N_986);
xnor U8978 (N_8978,N_3773,N_2557);
nand U8979 (N_8979,N_4241,N_4314);
nand U8980 (N_8980,N_1912,N_504);
nor U8981 (N_8981,N_508,N_4529);
nand U8982 (N_8982,N_1893,N_231);
nor U8983 (N_8983,N_159,N_2636);
nand U8984 (N_8984,N_4942,N_1322);
nand U8985 (N_8985,N_907,N_796);
nor U8986 (N_8986,N_2955,N_2345);
xnor U8987 (N_8987,N_3254,N_2870);
nor U8988 (N_8988,N_3118,N_4042);
nand U8989 (N_8989,N_3242,N_1117);
and U8990 (N_8990,N_3404,N_4578);
and U8991 (N_8991,N_67,N_965);
and U8992 (N_8992,N_2189,N_4164);
nand U8993 (N_8993,N_3435,N_1563);
xnor U8994 (N_8994,N_1087,N_4951);
nor U8995 (N_8995,N_2050,N_4779);
or U8996 (N_8996,N_4067,N_498);
and U8997 (N_8997,N_3026,N_4058);
and U8998 (N_8998,N_2222,N_2731);
nand U8999 (N_8999,N_973,N_4635);
nand U9000 (N_9000,N_3491,N_1383);
and U9001 (N_9001,N_1895,N_4284);
xor U9002 (N_9002,N_4534,N_1813);
nor U9003 (N_9003,N_4138,N_4245);
or U9004 (N_9004,N_4512,N_3712);
or U9005 (N_9005,N_192,N_412);
nand U9006 (N_9006,N_176,N_4047);
nor U9007 (N_9007,N_3918,N_2487);
xor U9008 (N_9008,N_2422,N_1833);
nand U9009 (N_9009,N_3545,N_1732);
or U9010 (N_9010,N_2223,N_3569);
xnor U9011 (N_9011,N_3755,N_4014);
nand U9012 (N_9012,N_3017,N_4033);
or U9013 (N_9013,N_4659,N_852);
or U9014 (N_9014,N_177,N_2838);
or U9015 (N_9015,N_649,N_1702);
or U9016 (N_9016,N_4731,N_3363);
and U9017 (N_9017,N_2966,N_2033);
nor U9018 (N_9018,N_35,N_91);
and U9019 (N_9019,N_2306,N_3339);
and U9020 (N_9020,N_363,N_443);
nor U9021 (N_9021,N_2193,N_808);
or U9022 (N_9022,N_1513,N_200);
and U9023 (N_9023,N_1061,N_1611);
nand U9024 (N_9024,N_3247,N_4738);
nor U9025 (N_9025,N_1787,N_419);
nor U9026 (N_9026,N_3254,N_2145);
nor U9027 (N_9027,N_630,N_4970);
nand U9028 (N_9028,N_1213,N_3097);
or U9029 (N_9029,N_43,N_4307);
nand U9030 (N_9030,N_3935,N_3628);
and U9031 (N_9031,N_1647,N_3834);
nor U9032 (N_9032,N_4257,N_42);
xnor U9033 (N_9033,N_2226,N_2814);
or U9034 (N_9034,N_2285,N_4029);
nand U9035 (N_9035,N_800,N_2077);
nor U9036 (N_9036,N_113,N_4169);
xnor U9037 (N_9037,N_3226,N_3888);
or U9038 (N_9038,N_521,N_4265);
and U9039 (N_9039,N_1057,N_4256);
nand U9040 (N_9040,N_1898,N_2343);
nor U9041 (N_9041,N_2533,N_1034);
or U9042 (N_9042,N_3698,N_2156);
nand U9043 (N_9043,N_1321,N_150);
xnor U9044 (N_9044,N_449,N_3947);
nor U9045 (N_9045,N_4085,N_212);
nor U9046 (N_9046,N_3177,N_1496);
and U9047 (N_9047,N_877,N_2528);
xnor U9048 (N_9048,N_4290,N_3896);
or U9049 (N_9049,N_1950,N_3940);
or U9050 (N_9050,N_1636,N_2444);
xor U9051 (N_9051,N_4497,N_1383);
nand U9052 (N_9052,N_1478,N_2077);
nand U9053 (N_9053,N_2558,N_1320);
and U9054 (N_9054,N_2388,N_2406);
nand U9055 (N_9055,N_4045,N_1878);
xor U9056 (N_9056,N_2131,N_4951);
nor U9057 (N_9057,N_57,N_818);
nand U9058 (N_9058,N_2542,N_4159);
or U9059 (N_9059,N_3677,N_2911);
and U9060 (N_9060,N_3421,N_4560);
and U9061 (N_9061,N_3536,N_4343);
nand U9062 (N_9062,N_1415,N_4341);
nand U9063 (N_9063,N_4185,N_3023);
or U9064 (N_9064,N_4166,N_4536);
nand U9065 (N_9065,N_1684,N_1765);
nand U9066 (N_9066,N_4587,N_1861);
and U9067 (N_9067,N_4960,N_2958);
nand U9068 (N_9068,N_2466,N_4824);
nor U9069 (N_9069,N_4745,N_308);
and U9070 (N_9070,N_1900,N_1134);
or U9071 (N_9071,N_4020,N_1889);
nor U9072 (N_9072,N_85,N_787);
nand U9073 (N_9073,N_695,N_4523);
and U9074 (N_9074,N_2019,N_2351);
nand U9075 (N_9075,N_161,N_2033);
nor U9076 (N_9076,N_1990,N_2141);
or U9077 (N_9077,N_2119,N_600);
nor U9078 (N_9078,N_4109,N_3257);
nand U9079 (N_9079,N_2485,N_4778);
or U9080 (N_9080,N_3676,N_4746);
nand U9081 (N_9081,N_798,N_2375);
and U9082 (N_9082,N_3714,N_1567);
and U9083 (N_9083,N_4491,N_4601);
nand U9084 (N_9084,N_4431,N_1654);
and U9085 (N_9085,N_2138,N_4625);
nor U9086 (N_9086,N_870,N_1651);
nand U9087 (N_9087,N_2582,N_2878);
and U9088 (N_9088,N_3506,N_4042);
nor U9089 (N_9089,N_584,N_3331);
and U9090 (N_9090,N_1669,N_939);
nor U9091 (N_9091,N_4108,N_3784);
or U9092 (N_9092,N_3239,N_4187);
nand U9093 (N_9093,N_3557,N_3907);
nand U9094 (N_9094,N_1703,N_3217);
or U9095 (N_9095,N_2325,N_1688);
and U9096 (N_9096,N_1525,N_2782);
xnor U9097 (N_9097,N_1307,N_2936);
and U9098 (N_9098,N_400,N_624);
nand U9099 (N_9099,N_4982,N_2009);
or U9100 (N_9100,N_3501,N_2016);
nor U9101 (N_9101,N_4137,N_468);
or U9102 (N_9102,N_173,N_4140);
nand U9103 (N_9103,N_1965,N_2992);
nor U9104 (N_9104,N_266,N_853);
nand U9105 (N_9105,N_4007,N_1827);
and U9106 (N_9106,N_4442,N_1577);
nor U9107 (N_9107,N_4246,N_2155);
nor U9108 (N_9108,N_4581,N_4696);
or U9109 (N_9109,N_1263,N_3637);
and U9110 (N_9110,N_3299,N_2383);
nor U9111 (N_9111,N_4647,N_1708);
and U9112 (N_9112,N_3261,N_2470);
nor U9113 (N_9113,N_37,N_1946);
nand U9114 (N_9114,N_3853,N_366);
and U9115 (N_9115,N_1682,N_3508);
and U9116 (N_9116,N_3896,N_3874);
xor U9117 (N_9117,N_2331,N_3659);
and U9118 (N_9118,N_181,N_3957);
xnor U9119 (N_9119,N_208,N_2544);
and U9120 (N_9120,N_4604,N_2070);
nand U9121 (N_9121,N_3805,N_1877);
nand U9122 (N_9122,N_1117,N_602);
nand U9123 (N_9123,N_3853,N_1723);
nand U9124 (N_9124,N_3857,N_1150);
and U9125 (N_9125,N_1420,N_1676);
or U9126 (N_9126,N_4200,N_2005);
nand U9127 (N_9127,N_3579,N_3702);
nand U9128 (N_9128,N_3401,N_4325);
or U9129 (N_9129,N_3877,N_2164);
nor U9130 (N_9130,N_1077,N_4911);
or U9131 (N_9131,N_3019,N_3540);
nor U9132 (N_9132,N_3231,N_4424);
and U9133 (N_9133,N_2458,N_2615);
nor U9134 (N_9134,N_2846,N_763);
nand U9135 (N_9135,N_257,N_2893);
nor U9136 (N_9136,N_157,N_2784);
and U9137 (N_9137,N_2215,N_2667);
nand U9138 (N_9138,N_3029,N_1823);
xnor U9139 (N_9139,N_3727,N_2699);
nand U9140 (N_9140,N_2484,N_4519);
nor U9141 (N_9141,N_550,N_2871);
nand U9142 (N_9142,N_147,N_169);
or U9143 (N_9143,N_2769,N_4294);
and U9144 (N_9144,N_4268,N_1000);
or U9145 (N_9145,N_625,N_516);
and U9146 (N_9146,N_1958,N_2593);
nor U9147 (N_9147,N_1700,N_1014);
and U9148 (N_9148,N_3583,N_1272);
nor U9149 (N_9149,N_2561,N_3555);
and U9150 (N_9150,N_968,N_1926);
nand U9151 (N_9151,N_520,N_228);
nor U9152 (N_9152,N_2574,N_1985);
nor U9153 (N_9153,N_347,N_3780);
nand U9154 (N_9154,N_3627,N_909);
nor U9155 (N_9155,N_4218,N_2224);
and U9156 (N_9156,N_2869,N_4140);
nand U9157 (N_9157,N_1610,N_66);
and U9158 (N_9158,N_4875,N_2157);
and U9159 (N_9159,N_4727,N_611);
nand U9160 (N_9160,N_152,N_3893);
and U9161 (N_9161,N_330,N_3105);
nor U9162 (N_9162,N_2411,N_4760);
xnor U9163 (N_9163,N_1329,N_2870);
nand U9164 (N_9164,N_3272,N_2711);
nor U9165 (N_9165,N_1174,N_54);
nand U9166 (N_9166,N_2841,N_1377);
or U9167 (N_9167,N_1617,N_4457);
nor U9168 (N_9168,N_430,N_2320);
or U9169 (N_9169,N_1506,N_4613);
nand U9170 (N_9170,N_1240,N_3651);
and U9171 (N_9171,N_4618,N_3490);
xnor U9172 (N_9172,N_3624,N_2947);
or U9173 (N_9173,N_3920,N_1780);
or U9174 (N_9174,N_4343,N_98);
and U9175 (N_9175,N_4237,N_1821);
nand U9176 (N_9176,N_3071,N_1750);
and U9177 (N_9177,N_4876,N_499);
nand U9178 (N_9178,N_30,N_4136);
nor U9179 (N_9179,N_918,N_1825);
nor U9180 (N_9180,N_4231,N_1925);
and U9181 (N_9181,N_3612,N_2575);
and U9182 (N_9182,N_3244,N_1353);
or U9183 (N_9183,N_2413,N_3534);
nor U9184 (N_9184,N_663,N_3899);
or U9185 (N_9185,N_1605,N_912);
or U9186 (N_9186,N_1228,N_126);
or U9187 (N_9187,N_2014,N_4384);
nor U9188 (N_9188,N_2894,N_2146);
xnor U9189 (N_9189,N_1904,N_4701);
or U9190 (N_9190,N_3169,N_3089);
xor U9191 (N_9191,N_3215,N_981);
or U9192 (N_9192,N_1910,N_2076);
nand U9193 (N_9193,N_1156,N_1227);
or U9194 (N_9194,N_1117,N_4067);
and U9195 (N_9195,N_2116,N_1196);
and U9196 (N_9196,N_3783,N_3453);
or U9197 (N_9197,N_1534,N_1131);
nor U9198 (N_9198,N_3703,N_4294);
nor U9199 (N_9199,N_251,N_1231);
or U9200 (N_9200,N_395,N_3382);
or U9201 (N_9201,N_506,N_4333);
and U9202 (N_9202,N_2449,N_518);
xor U9203 (N_9203,N_2874,N_4374);
or U9204 (N_9204,N_3629,N_3312);
and U9205 (N_9205,N_4164,N_3212);
nand U9206 (N_9206,N_2175,N_2171);
nand U9207 (N_9207,N_451,N_1639);
nand U9208 (N_9208,N_558,N_4562);
nand U9209 (N_9209,N_928,N_355);
nand U9210 (N_9210,N_984,N_4388);
or U9211 (N_9211,N_1158,N_707);
or U9212 (N_9212,N_1047,N_2673);
nor U9213 (N_9213,N_1776,N_232);
or U9214 (N_9214,N_4665,N_1628);
nor U9215 (N_9215,N_2228,N_3361);
nand U9216 (N_9216,N_147,N_4806);
or U9217 (N_9217,N_1276,N_3337);
or U9218 (N_9218,N_2851,N_3241);
or U9219 (N_9219,N_230,N_3162);
xor U9220 (N_9220,N_2597,N_3419);
and U9221 (N_9221,N_457,N_2369);
and U9222 (N_9222,N_4526,N_4217);
and U9223 (N_9223,N_312,N_1838);
xor U9224 (N_9224,N_1669,N_4040);
nand U9225 (N_9225,N_801,N_1768);
or U9226 (N_9226,N_0,N_1906);
and U9227 (N_9227,N_267,N_3477);
and U9228 (N_9228,N_1034,N_2618);
and U9229 (N_9229,N_4952,N_190);
nand U9230 (N_9230,N_3602,N_1757);
or U9231 (N_9231,N_1417,N_2933);
xnor U9232 (N_9232,N_2164,N_4189);
xnor U9233 (N_9233,N_4931,N_2731);
nor U9234 (N_9234,N_4930,N_3274);
or U9235 (N_9235,N_442,N_4471);
nand U9236 (N_9236,N_1309,N_3786);
or U9237 (N_9237,N_4663,N_3739);
or U9238 (N_9238,N_1041,N_2880);
nor U9239 (N_9239,N_1151,N_2814);
or U9240 (N_9240,N_2440,N_4576);
xnor U9241 (N_9241,N_2988,N_4863);
nand U9242 (N_9242,N_1976,N_4244);
nor U9243 (N_9243,N_3321,N_3001);
xnor U9244 (N_9244,N_78,N_2865);
nand U9245 (N_9245,N_4011,N_716);
and U9246 (N_9246,N_4745,N_562);
nand U9247 (N_9247,N_434,N_449);
or U9248 (N_9248,N_4910,N_2675);
nor U9249 (N_9249,N_106,N_2427);
and U9250 (N_9250,N_2941,N_3622);
nor U9251 (N_9251,N_3246,N_1487);
nand U9252 (N_9252,N_109,N_4921);
nor U9253 (N_9253,N_1707,N_4341);
or U9254 (N_9254,N_2752,N_539);
nand U9255 (N_9255,N_382,N_1822);
nor U9256 (N_9256,N_24,N_736);
and U9257 (N_9257,N_2308,N_1615);
and U9258 (N_9258,N_3048,N_252);
or U9259 (N_9259,N_2259,N_2739);
or U9260 (N_9260,N_1472,N_4850);
or U9261 (N_9261,N_973,N_606);
nand U9262 (N_9262,N_1217,N_357);
nand U9263 (N_9263,N_898,N_1728);
xnor U9264 (N_9264,N_4413,N_665);
nor U9265 (N_9265,N_1678,N_4552);
nor U9266 (N_9266,N_3670,N_2712);
xor U9267 (N_9267,N_707,N_4670);
nor U9268 (N_9268,N_4505,N_4888);
nand U9269 (N_9269,N_2013,N_2238);
nor U9270 (N_9270,N_3357,N_4426);
or U9271 (N_9271,N_1061,N_364);
xor U9272 (N_9272,N_4231,N_1170);
nand U9273 (N_9273,N_4995,N_1814);
and U9274 (N_9274,N_3828,N_1826);
nor U9275 (N_9275,N_2676,N_417);
nor U9276 (N_9276,N_4425,N_345);
xor U9277 (N_9277,N_3959,N_4573);
and U9278 (N_9278,N_988,N_4901);
nand U9279 (N_9279,N_1743,N_1477);
and U9280 (N_9280,N_3678,N_1917);
or U9281 (N_9281,N_2548,N_4078);
nor U9282 (N_9282,N_3289,N_2301);
or U9283 (N_9283,N_2031,N_4769);
nor U9284 (N_9284,N_2515,N_174);
and U9285 (N_9285,N_254,N_4990);
and U9286 (N_9286,N_3044,N_3556);
nand U9287 (N_9287,N_3940,N_3337);
nor U9288 (N_9288,N_1160,N_4616);
nor U9289 (N_9289,N_4625,N_46);
xor U9290 (N_9290,N_1449,N_611);
nand U9291 (N_9291,N_3453,N_1868);
or U9292 (N_9292,N_3792,N_2393);
nand U9293 (N_9293,N_4009,N_2908);
nor U9294 (N_9294,N_3948,N_3383);
xnor U9295 (N_9295,N_4566,N_4535);
nor U9296 (N_9296,N_3456,N_1784);
nor U9297 (N_9297,N_1889,N_3084);
nand U9298 (N_9298,N_869,N_81);
nand U9299 (N_9299,N_1793,N_4997);
nor U9300 (N_9300,N_936,N_1546);
and U9301 (N_9301,N_4853,N_3627);
and U9302 (N_9302,N_90,N_3710);
nand U9303 (N_9303,N_1894,N_3493);
nor U9304 (N_9304,N_3163,N_2787);
nand U9305 (N_9305,N_4977,N_1472);
nor U9306 (N_9306,N_4324,N_4814);
nand U9307 (N_9307,N_173,N_32);
or U9308 (N_9308,N_255,N_1367);
nand U9309 (N_9309,N_2699,N_4364);
nand U9310 (N_9310,N_2480,N_2466);
or U9311 (N_9311,N_4023,N_900);
or U9312 (N_9312,N_448,N_1430);
and U9313 (N_9313,N_1300,N_4789);
and U9314 (N_9314,N_1504,N_4515);
nor U9315 (N_9315,N_4227,N_4980);
and U9316 (N_9316,N_2721,N_992);
or U9317 (N_9317,N_3370,N_3452);
or U9318 (N_9318,N_3387,N_206);
and U9319 (N_9319,N_896,N_3400);
nor U9320 (N_9320,N_1277,N_3218);
nand U9321 (N_9321,N_764,N_4670);
nand U9322 (N_9322,N_87,N_97);
or U9323 (N_9323,N_4418,N_630);
or U9324 (N_9324,N_3749,N_2703);
or U9325 (N_9325,N_2731,N_3856);
nor U9326 (N_9326,N_1629,N_3520);
xnor U9327 (N_9327,N_694,N_3498);
nor U9328 (N_9328,N_1714,N_1932);
nand U9329 (N_9329,N_1641,N_2224);
or U9330 (N_9330,N_2717,N_551);
or U9331 (N_9331,N_2780,N_4479);
nor U9332 (N_9332,N_1954,N_4345);
xor U9333 (N_9333,N_697,N_338);
xor U9334 (N_9334,N_4537,N_2493);
xor U9335 (N_9335,N_2169,N_721);
and U9336 (N_9336,N_2232,N_1488);
nand U9337 (N_9337,N_2751,N_3816);
nor U9338 (N_9338,N_2085,N_2625);
nor U9339 (N_9339,N_1960,N_4908);
nand U9340 (N_9340,N_1511,N_1001);
nor U9341 (N_9341,N_2825,N_3788);
and U9342 (N_9342,N_432,N_3561);
nor U9343 (N_9343,N_1828,N_1026);
or U9344 (N_9344,N_2385,N_3564);
or U9345 (N_9345,N_2604,N_900);
nand U9346 (N_9346,N_4838,N_4996);
nand U9347 (N_9347,N_583,N_3678);
nor U9348 (N_9348,N_2074,N_2299);
nand U9349 (N_9349,N_1004,N_1103);
or U9350 (N_9350,N_842,N_2088);
nand U9351 (N_9351,N_4173,N_3643);
nand U9352 (N_9352,N_341,N_3373);
and U9353 (N_9353,N_2494,N_1560);
and U9354 (N_9354,N_3094,N_126);
nor U9355 (N_9355,N_3548,N_2673);
or U9356 (N_9356,N_307,N_1850);
or U9357 (N_9357,N_1526,N_1472);
nand U9358 (N_9358,N_4530,N_1778);
nand U9359 (N_9359,N_395,N_1548);
or U9360 (N_9360,N_1051,N_494);
xor U9361 (N_9361,N_2736,N_288);
nor U9362 (N_9362,N_3099,N_1447);
nand U9363 (N_9363,N_2036,N_2922);
nor U9364 (N_9364,N_1650,N_244);
or U9365 (N_9365,N_2311,N_4507);
nand U9366 (N_9366,N_4168,N_4344);
nand U9367 (N_9367,N_1919,N_4874);
nor U9368 (N_9368,N_2070,N_925);
and U9369 (N_9369,N_585,N_1267);
or U9370 (N_9370,N_1278,N_2364);
nor U9371 (N_9371,N_190,N_2201);
and U9372 (N_9372,N_4932,N_2150);
or U9373 (N_9373,N_1475,N_2428);
nand U9374 (N_9374,N_3732,N_4246);
and U9375 (N_9375,N_2269,N_1151);
nand U9376 (N_9376,N_1851,N_3895);
nor U9377 (N_9377,N_2602,N_2423);
nor U9378 (N_9378,N_2049,N_3107);
nor U9379 (N_9379,N_3725,N_3820);
and U9380 (N_9380,N_521,N_652);
or U9381 (N_9381,N_1254,N_3957);
nor U9382 (N_9382,N_4807,N_3956);
nand U9383 (N_9383,N_4394,N_3721);
or U9384 (N_9384,N_4935,N_996);
nand U9385 (N_9385,N_689,N_3867);
nor U9386 (N_9386,N_2938,N_4266);
nand U9387 (N_9387,N_1575,N_3195);
nor U9388 (N_9388,N_4416,N_2125);
and U9389 (N_9389,N_388,N_2635);
nand U9390 (N_9390,N_4735,N_4203);
or U9391 (N_9391,N_2811,N_3120);
nor U9392 (N_9392,N_2939,N_824);
or U9393 (N_9393,N_595,N_4556);
nand U9394 (N_9394,N_388,N_2362);
xnor U9395 (N_9395,N_4642,N_425);
and U9396 (N_9396,N_1278,N_1335);
nor U9397 (N_9397,N_2066,N_4580);
or U9398 (N_9398,N_4961,N_4762);
nand U9399 (N_9399,N_1793,N_1951);
nor U9400 (N_9400,N_4297,N_3591);
nor U9401 (N_9401,N_4690,N_3415);
xnor U9402 (N_9402,N_331,N_1842);
nor U9403 (N_9403,N_304,N_4990);
nand U9404 (N_9404,N_4558,N_192);
or U9405 (N_9405,N_188,N_3026);
or U9406 (N_9406,N_4392,N_395);
or U9407 (N_9407,N_1147,N_3296);
and U9408 (N_9408,N_2350,N_2776);
xnor U9409 (N_9409,N_2052,N_3093);
nand U9410 (N_9410,N_2980,N_2468);
nand U9411 (N_9411,N_2033,N_910);
nor U9412 (N_9412,N_763,N_1250);
and U9413 (N_9413,N_983,N_398);
nand U9414 (N_9414,N_789,N_3310);
or U9415 (N_9415,N_1921,N_4419);
or U9416 (N_9416,N_4346,N_3705);
and U9417 (N_9417,N_3982,N_4862);
nor U9418 (N_9418,N_810,N_3983);
nand U9419 (N_9419,N_4819,N_2081);
or U9420 (N_9420,N_2200,N_1831);
nand U9421 (N_9421,N_60,N_2289);
nor U9422 (N_9422,N_980,N_2311);
xnor U9423 (N_9423,N_959,N_2002);
nor U9424 (N_9424,N_3971,N_1434);
and U9425 (N_9425,N_3832,N_3793);
and U9426 (N_9426,N_1936,N_4140);
xor U9427 (N_9427,N_2780,N_3921);
nand U9428 (N_9428,N_4824,N_1953);
and U9429 (N_9429,N_1405,N_2944);
and U9430 (N_9430,N_1910,N_1552);
or U9431 (N_9431,N_4116,N_126);
nor U9432 (N_9432,N_3408,N_777);
or U9433 (N_9433,N_1969,N_4466);
xnor U9434 (N_9434,N_1605,N_4463);
xnor U9435 (N_9435,N_1029,N_4176);
or U9436 (N_9436,N_4800,N_4532);
or U9437 (N_9437,N_4845,N_981);
or U9438 (N_9438,N_3513,N_80);
or U9439 (N_9439,N_4981,N_1988);
or U9440 (N_9440,N_4398,N_4525);
nor U9441 (N_9441,N_2876,N_4060);
or U9442 (N_9442,N_1316,N_786);
xor U9443 (N_9443,N_3289,N_2029);
nand U9444 (N_9444,N_510,N_1803);
xnor U9445 (N_9445,N_1165,N_4021);
nand U9446 (N_9446,N_842,N_4196);
or U9447 (N_9447,N_2809,N_1094);
or U9448 (N_9448,N_80,N_2912);
nor U9449 (N_9449,N_4350,N_1135);
nor U9450 (N_9450,N_4487,N_3876);
nor U9451 (N_9451,N_3189,N_4741);
nand U9452 (N_9452,N_2739,N_1709);
xor U9453 (N_9453,N_920,N_4322);
and U9454 (N_9454,N_3518,N_2370);
nor U9455 (N_9455,N_4927,N_3875);
or U9456 (N_9456,N_4188,N_2356);
or U9457 (N_9457,N_3860,N_3856);
and U9458 (N_9458,N_1211,N_3423);
nor U9459 (N_9459,N_239,N_3292);
and U9460 (N_9460,N_4562,N_2514);
and U9461 (N_9461,N_4863,N_944);
nand U9462 (N_9462,N_3476,N_137);
and U9463 (N_9463,N_4313,N_786);
nor U9464 (N_9464,N_4641,N_2290);
nor U9465 (N_9465,N_96,N_808);
or U9466 (N_9466,N_293,N_2254);
or U9467 (N_9467,N_3364,N_3185);
or U9468 (N_9468,N_4160,N_673);
nand U9469 (N_9469,N_2260,N_2766);
or U9470 (N_9470,N_2771,N_540);
nand U9471 (N_9471,N_1501,N_2388);
and U9472 (N_9472,N_3404,N_3451);
or U9473 (N_9473,N_2242,N_927);
xnor U9474 (N_9474,N_4550,N_320);
and U9475 (N_9475,N_1623,N_3737);
and U9476 (N_9476,N_1419,N_715);
nand U9477 (N_9477,N_1896,N_4821);
nor U9478 (N_9478,N_4922,N_697);
xnor U9479 (N_9479,N_53,N_47);
or U9480 (N_9480,N_3757,N_1325);
or U9481 (N_9481,N_2819,N_798);
and U9482 (N_9482,N_1769,N_2676);
nand U9483 (N_9483,N_4283,N_4821);
nand U9484 (N_9484,N_1770,N_1497);
nor U9485 (N_9485,N_859,N_2767);
nand U9486 (N_9486,N_2680,N_1366);
and U9487 (N_9487,N_3405,N_539);
nor U9488 (N_9488,N_2943,N_3016);
or U9489 (N_9489,N_1258,N_2679);
nand U9490 (N_9490,N_4552,N_4818);
nor U9491 (N_9491,N_3794,N_4362);
and U9492 (N_9492,N_1504,N_990);
or U9493 (N_9493,N_1307,N_2407);
or U9494 (N_9494,N_1275,N_318);
nor U9495 (N_9495,N_4964,N_3889);
nor U9496 (N_9496,N_2724,N_457);
nor U9497 (N_9497,N_3956,N_3745);
and U9498 (N_9498,N_1430,N_855);
and U9499 (N_9499,N_781,N_2048);
nand U9500 (N_9500,N_1316,N_2064);
nand U9501 (N_9501,N_1677,N_816);
or U9502 (N_9502,N_209,N_1389);
or U9503 (N_9503,N_2745,N_4824);
xnor U9504 (N_9504,N_1294,N_4057);
xnor U9505 (N_9505,N_2669,N_553);
nand U9506 (N_9506,N_3538,N_4740);
nor U9507 (N_9507,N_4414,N_772);
nor U9508 (N_9508,N_4312,N_325);
or U9509 (N_9509,N_596,N_4545);
and U9510 (N_9510,N_4722,N_3002);
xnor U9511 (N_9511,N_2844,N_1558);
nand U9512 (N_9512,N_4611,N_2082);
nor U9513 (N_9513,N_4225,N_2290);
nand U9514 (N_9514,N_160,N_1948);
or U9515 (N_9515,N_1836,N_4669);
xor U9516 (N_9516,N_4443,N_459);
or U9517 (N_9517,N_470,N_4340);
or U9518 (N_9518,N_3631,N_2377);
nor U9519 (N_9519,N_3017,N_2135);
nor U9520 (N_9520,N_522,N_4544);
xnor U9521 (N_9521,N_4549,N_3721);
nor U9522 (N_9522,N_1949,N_4659);
and U9523 (N_9523,N_1430,N_4576);
nand U9524 (N_9524,N_3924,N_4729);
and U9525 (N_9525,N_1272,N_1668);
nor U9526 (N_9526,N_2217,N_4984);
nand U9527 (N_9527,N_1898,N_3088);
or U9528 (N_9528,N_1884,N_534);
nand U9529 (N_9529,N_50,N_2189);
nand U9530 (N_9530,N_3168,N_1650);
xnor U9531 (N_9531,N_768,N_3149);
xor U9532 (N_9532,N_3709,N_1473);
and U9533 (N_9533,N_3163,N_1364);
nand U9534 (N_9534,N_998,N_2841);
nand U9535 (N_9535,N_382,N_2911);
xnor U9536 (N_9536,N_2720,N_4509);
and U9537 (N_9537,N_2345,N_1535);
and U9538 (N_9538,N_361,N_3079);
or U9539 (N_9539,N_1606,N_3512);
nor U9540 (N_9540,N_203,N_1307);
or U9541 (N_9541,N_2722,N_4459);
nor U9542 (N_9542,N_132,N_2419);
or U9543 (N_9543,N_4957,N_3498);
nand U9544 (N_9544,N_907,N_491);
and U9545 (N_9545,N_1833,N_634);
nand U9546 (N_9546,N_3928,N_4624);
nand U9547 (N_9547,N_3545,N_1267);
and U9548 (N_9548,N_1217,N_3904);
nand U9549 (N_9549,N_3017,N_2168);
xor U9550 (N_9550,N_4769,N_2875);
and U9551 (N_9551,N_3720,N_3444);
or U9552 (N_9552,N_1704,N_3486);
nand U9553 (N_9553,N_1424,N_4520);
or U9554 (N_9554,N_3578,N_4749);
nor U9555 (N_9555,N_1189,N_3254);
nor U9556 (N_9556,N_4838,N_3669);
nor U9557 (N_9557,N_4780,N_2261);
nand U9558 (N_9558,N_612,N_2555);
and U9559 (N_9559,N_727,N_1604);
nor U9560 (N_9560,N_3524,N_470);
and U9561 (N_9561,N_2830,N_2034);
or U9562 (N_9562,N_454,N_1086);
or U9563 (N_9563,N_3,N_2937);
nor U9564 (N_9564,N_4131,N_4705);
nand U9565 (N_9565,N_1689,N_2149);
or U9566 (N_9566,N_1847,N_1667);
or U9567 (N_9567,N_2191,N_3520);
nor U9568 (N_9568,N_722,N_4451);
or U9569 (N_9569,N_1570,N_2799);
nand U9570 (N_9570,N_2979,N_1865);
and U9571 (N_9571,N_3960,N_306);
and U9572 (N_9572,N_562,N_2911);
or U9573 (N_9573,N_4769,N_510);
nand U9574 (N_9574,N_961,N_2632);
nor U9575 (N_9575,N_1043,N_2473);
nand U9576 (N_9576,N_217,N_3097);
nor U9577 (N_9577,N_4284,N_2237);
nor U9578 (N_9578,N_3696,N_2345);
nand U9579 (N_9579,N_3473,N_2128);
nand U9580 (N_9580,N_3263,N_1142);
nor U9581 (N_9581,N_3078,N_4688);
or U9582 (N_9582,N_3132,N_4997);
nor U9583 (N_9583,N_114,N_1891);
nand U9584 (N_9584,N_3323,N_2342);
xor U9585 (N_9585,N_1543,N_3543);
nand U9586 (N_9586,N_419,N_3045);
or U9587 (N_9587,N_4908,N_2766);
xor U9588 (N_9588,N_4467,N_1231);
or U9589 (N_9589,N_4516,N_1776);
or U9590 (N_9590,N_4828,N_830);
or U9591 (N_9591,N_3574,N_1653);
nor U9592 (N_9592,N_1592,N_3158);
and U9593 (N_9593,N_3187,N_4481);
or U9594 (N_9594,N_2669,N_1314);
nor U9595 (N_9595,N_3794,N_920);
or U9596 (N_9596,N_3675,N_2471);
nand U9597 (N_9597,N_3841,N_3961);
or U9598 (N_9598,N_4570,N_1567);
nor U9599 (N_9599,N_2940,N_2643);
nand U9600 (N_9600,N_2377,N_4425);
nand U9601 (N_9601,N_1890,N_3933);
and U9602 (N_9602,N_671,N_4230);
and U9603 (N_9603,N_1096,N_1137);
or U9604 (N_9604,N_3993,N_4478);
xor U9605 (N_9605,N_4347,N_3829);
or U9606 (N_9606,N_2816,N_887);
or U9607 (N_9607,N_1106,N_3010);
nor U9608 (N_9608,N_4247,N_1077);
nor U9609 (N_9609,N_3354,N_3668);
nor U9610 (N_9610,N_4972,N_4809);
xor U9611 (N_9611,N_1132,N_1485);
nand U9612 (N_9612,N_3053,N_1483);
nand U9613 (N_9613,N_2207,N_10);
or U9614 (N_9614,N_2697,N_183);
nor U9615 (N_9615,N_3983,N_889);
xnor U9616 (N_9616,N_3856,N_2398);
and U9617 (N_9617,N_4424,N_4266);
and U9618 (N_9618,N_240,N_1055);
nand U9619 (N_9619,N_3649,N_3444);
and U9620 (N_9620,N_3810,N_688);
and U9621 (N_9621,N_2098,N_3267);
or U9622 (N_9622,N_2889,N_585);
xor U9623 (N_9623,N_3456,N_3686);
or U9624 (N_9624,N_2637,N_1042);
nor U9625 (N_9625,N_3011,N_2893);
and U9626 (N_9626,N_2065,N_1685);
nand U9627 (N_9627,N_1509,N_489);
and U9628 (N_9628,N_754,N_1038);
nand U9629 (N_9629,N_67,N_782);
xor U9630 (N_9630,N_1594,N_999);
or U9631 (N_9631,N_700,N_202);
nor U9632 (N_9632,N_132,N_3355);
and U9633 (N_9633,N_1922,N_2090);
nand U9634 (N_9634,N_1857,N_1382);
or U9635 (N_9635,N_3073,N_2042);
nand U9636 (N_9636,N_372,N_2687);
and U9637 (N_9637,N_3514,N_307);
or U9638 (N_9638,N_4127,N_3548);
and U9639 (N_9639,N_3045,N_2500);
and U9640 (N_9640,N_4571,N_2882);
and U9641 (N_9641,N_4453,N_4729);
nand U9642 (N_9642,N_4161,N_3083);
xnor U9643 (N_9643,N_2987,N_4977);
nor U9644 (N_9644,N_1662,N_4249);
nand U9645 (N_9645,N_2244,N_4746);
nor U9646 (N_9646,N_3468,N_209);
nand U9647 (N_9647,N_1551,N_3477);
nor U9648 (N_9648,N_709,N_2695);
and U9649 (N_9649,N_205,N_2651);
nor U9650 (N_9650,N_1317,N_2056);
nor U9651 (N_9651,N_1761,N_4158);
or U9652 (N_9652,N_184,N_2014);
nand U9653 (N_9653,N_2129,N_2221);
nor U9654 (N_9654,N_2662,N_60);
nand U9655 (N_9655,N_3316,N_4772);
and U9656 (N_9656,N_3390,N_1643);
nand U9657 (N_9657,N_1639,N_2523);
nand U9658 (N_9658,N_4817,N_2877);
nand U9659 (N_9659,N_810,N_4290);
nand U9660 (N_9660,N_4756,N_574);
or U9661 (N_9661,N_1563,N_4297);
xor U9662 (N_9662,N_893,N_2898);
and U9663 (N_9663,N_1367,N_1910);
xor U9664 (N_9664,N_1680,N_68);
and U9665 (N_9665,N_3851,N_917);
and U9666 (N_9666,N_2676,N_144);
nand U9667 (N_9667,N_2885,N_2958);
nand U9668 (N_9668,N_3811,N_1312);
or U9669 (N_9669,N_27,N_241);
nand U9670 (N_9670,N_3466,N_2306);
and U9671 (N_9671,N_1994,N_616);
and U9672 (N_9672,N_1170,N_501);
xnor U9673 (N_9673,N_3036,N_1145);
or U9674 (N_9674,N_106,N_4278);
nand U9675 (N_9675,N_1918,N_4269);
xor U9676 (N_9676,N_1849,N_2496);
nand U9677 (N_9677,N_1450,N_2731);
or U9678 (N_9678,N_4919,N_2530);
nor U9679 (N_9679,N_1277,N_2587);
or U9680 (N_9680,N_4877,N_4508);
nor U9681 (N_9681,N_701,N_2075);
nor U9682 (N_9682,N_1611,N_2825);
and U9683 (N_9683,N_2826,N_4414);
nor U9684 (N_9684,N_3572,N_3977);
xor U9685 (N_9685,N_3725,N_821);
or U9686 (N_9686,N_3088,N_4338);
nand U9687 (N_9687,N_3124,N_2306);
nand U9688 (N_9688,N_149,N_3840);
and U9689 (N_9689,N_3988,N_1820);
and U9690 (N_9690,N_59,N_4201);
xnor U9691 (N_9691,N_3290,N_1517);
nor U9692 (N_9692,N_2085,N_650);
nand U9693 (N_9693,N_4042,N_3433);
nand U9694 (N_9694,N_4861,N_4200);
and U9695 (N_9695,N_4278,N_109);
or U9696 (N_9696,N_4708,N_4994);
nand U9697 (N_9697,N_1438,N_2260);
nor U9698 (N_9698,N_1114,N_1341);
or U9699 (N_9699,N_3953,N_762);
nand U9700 (N_9700,N_3894,N_1944);
nor U9701 (N_9701,N_4814,N_3015);
and U9702 (N_9702,N_4624,N_3227);
xor U9703 (N_9703,N_1906,N_1120);
and U9704 (N_9704,N_892,N_1416);
nand U9705 (N_9705,N_133,N_4584);
or U9706 (N_9706,N_3617,N_2815);
xor U9707 (N_9707,N_2966,N_3754);
or U9708 (N_9708,N_1190,N_3590);
nand U9709 (N_9709,N_501,N_3545);
nand U9710 (N_9710,N_3879,N_838);
nand U9711 (N_9711,N_2121,N_3767);
and U9712 (N_9712,N_4567,N_712);
nor U9713 (N_9713,N_3198,N_5);
and U9714 (N_9714,N_3219,N_364);
xnor U9715 (N_9715,N_2519,N_4408);
or U9716 (N_9716,N_4450,N_4191);
or U9717 (N_9717,N_2452,N_4484);
xor U9718 (N_9718,N_516,N_2183);
and U9719 (N_9719,N_1987,N_3912);
nor U9720 (N_9720,N_1643,N_4057);
xnor U9721 (N_9721,N_2149,N_1751);
nor U9722 (N_9722,N_4250,N_573);
nand U9723 (N_9723,N_3008,N_3613);
nand U9724 (N_9724,N_3988,N_291);
xor U9725 (N_9725,N_1976,N_4856);
xnor U9726 (N_9726,N_2968,N_1544);
and U9727 (N_9727,N_1612,N_3884);
and U9728 (N_9728,N_4047,N_2210);
and U9729 (N_9729,N_3736,N_4587);
or U9730 (N_9730,N_2146,N_2569);
xnor U9731 (N_9731,N_3733,N_2639);
nor U9732 (N_9732,N_4099,N_34);
or U9733 (N_9733,N_2796,N_162);
xor U9734 (N_9734,N_4932,N_1829);
or U9735 (N_9735,N_102,N_4566);
nand U9736 (N_9736,N_1378,N_2454);
and U9737 (N_9737,N_4526,N_4912);
and U9738 (N_9738,N_1825,N_3036);
nand U9739 (N_9739,N_381,N_1853);
and U9740 (N_9740,N_593,N_3030);
nor U9741 (N_9741,N_3930,N_4884);
xor U9742 (N_9742,N_3369,N_2831);
nand U9743 (N_9743,N_2375,N_980);
nand U9744 (N_9744,N_85,N_1397);
and U9745 (N_9745,N_3909,N_369);
nand U9746 (N_9746,N_3855,N_4194);
nor U9747 (N_9747,N_3064,N_972);
or U9748 (N_9748,N_3582,N_3631);
nor U9749 (N_9749,N_3284,N_4676);
nand U9750 (N_9750,N_1866,N_3334);
nand U9751 (N_9751,N_1988,N_2556);
or U9752 (N_9752,N_3874,N_2521);
nand U9753 (N_9753,N_764,N_1114);
nor U9754 (N_9754,N_3899,N_923);
and U9755 (N_9755,N_1564,N_1425);
nor U9756 (N_9756,N_4964,N_3893);
nand U9757 (N_9757,N_3819,N_34);
and U9758 (N_9758,N_1714,N_2536);
nor U9759 (N_9759,N_4061,N_4462);
nand U9760 (N_9760,N_1284,N_4404);
or U9761 (N_9761,N_2924,N_2086);
or U9762 (N_9762,N_1414,N_2920);
nand U9763 (N_9763,N_4383,N_3337);
nand U9764 (N_9764,N_4272,N_1166);
or U9765 (N_9765,N_2729,N_4648);
nor U9766 (N_9766,N_4484,N_3543);
nand U9767 (N_9767,N_210,N_4438);
or U9768 (N_9768,N_1134,N_2265);
nor U9769 (N_9769,N_1494,N_4130);
nor U9770 (N_9770,N_4033,N_3347);
and U9771 (N_9771,N_2113,N_872);
nor U9772 (N_9772,N_2771,N_714);
nor U9773 (N_9773,N_1009,N_283);
nand U9774 (N_9774,N_2634,N_2248);
and U9775 (N_9775,N_1202,N_4647);
nor U9776 (N_9776,N_2009,N_3899);
nand U9777 (N_9777,N_3686,N_3959);
nand U9778 (N_9778,N_602,N_548);
nor U9779 (N_9779,N_1017,N_4489);
and U9780 (N_9780,N_2955,N_2939);
and U9781 (N_9781,N_3133,N_3430);
and U9782 (N_9782,N_1683,N_2878);
or U9783 (N_9783,N_3604,N_1483);
nor U9784 (N_9784,N_4075,N_3630);
or U9785 (N_9785,N_2583,N_4720);
nor U9786 (N_9786,N_3718,N_3110);
nor U9787 (N_9787,N_2997,N_4455);
xor U9788 (N_9788,N_2459,N_1720);
and U9789 (N_9789,N_2926,N_3158);
and U9790 (N_9790,N_3182,N_2582);
or U9791 (N_9791,N_1347,N_2576);
xor U9792 (N_9792,N_2543,N_4982);
and U9793 (N_9793,N_1892,N_3211);
and U9794 (N_9794,N_109,N_4512);
nand U9795 (N_9795,N_3162,N_237);
nand U9796 (N_9796,N_3914,N_807);
xnor U9797 (N_9797,N_4212,N_1582);
nor U9798 (N_9798,N_4201,N_518);
nor U9799 (N_9799,N_2858,N_3528);
or U9800 (N_9800,N_31,N_4807);
or U9801 (N_9801,N_264,N_2175);
or U9802 (N_9802,N_8,N_3869);
or U9803 (N_9803,N_4722,N_2657);
and U9804 (N_9804,N_760,N_3218);
and U9805 (N_9805,N_1472,N_3347);
nand U9806 (N_9806,N_1317,N_769);
or U9807 (N_9807,N_134,N_3681);
nor U9808 (N_9808,N_1480,N_2456);
or U9809 (N_9809,N_2745,N_4909);
nand U9810 (N_9810,N_4280,N_2450);
nor U9811 (N_9811,N_3602,N_2665);
nand U9812 (N_9812,N_4443,N_522);
nand U9813 (N_9813,N_737,N_1267);
and U9814 (N_9814,N_2903,N_661);
or U9815 (N_9815,N_3068,N_1182);
or U9816 (N_9816,N_3057,N_412);
nor U9817 (N_9817,N_577,N_3588);
nand U9818 (N_9818,N_2062,N_2925);
or U9819 (N_9819,N_1795,N_1752);
nor U9820 (N_9820,N_2307,N_1725);
and U9821 (N_9821,N_4928,N_4748);
or U9822 (N_9822,N_4713,N_3620);
or U9823 (N_9823,N_587,N_3470);
nand U9824 (N_9824,N_3148,N_505);
nor U9825 (N_9825,N_3347,N_3548);
nor U9826 (N_9826,N_1948,N_4335);
nand U9827 (N_9827,N_1649,N_4984);
or U9828 (N_9828,N_787,N_3958);
and U9829 (N_9829,N_4873,N_3990);
nand U9830 (N_9830,N_1533,N_2302);
nor U9831 (N_9831,N_3610,N_2741);
nand U9832 (N_9832,N_769,N_4694);
nand U9833 (N_9833,N_4154,N_2053);
nor U9834 (N_9834,N_2051,N_763);
and U9835 (N_9835,N_906,N_3170);
nor U9836 (N_9836,N_2681,N_3563);
nor U9837 (N_9837,N_2744,N_2139);
nand U9838 (N_9838,N_445,N_4652);
nor U9839 (N_9839,N_3406,N_3041);
and U9840 (N_9840,N_1398,N_2407);
xor U9841 (N_9841,N_1821,N_1037);
nand U9842 (N_9842,N_4940,N_3340);
or U9843 (N_9843,N_3946,N_1820);
nor U9844 (N_9844,N_778,N_3853);
nand U9845 (N_9845,N_3684,N_3226);
and U9846 (N_9846,N_4345,N_2460);
nand U9847 (N_9847,N_1279,N_2514);
and U9848 (N_9848,N_3249,N_2520);
nand U9849 (N_9849,N_133,N_384);
or U9850 (N_9850,N_2476,N_3124);
and U9851 (N_9851,N_3993,N_4008);
xnor U9852 (N_9852,N_1621,N_3515);
nor U9853 (N_9853,N_347,N_441);
and U9854 (N_9854,N_3223,N_2346);
nor U9855 (N_9855,N_751,N_2003);
or U9856 (N_9856,N_3321,N_4803);
and U9857 (N_9857,N_2566,N_2980);
nor U9858 (N_9858,N_242,N_1441);
and U9859 (N_9859,N_4197,N_717);
and U9860 (N_9860,N_1035,N_3383);
nand U9861 (N_9861,N_2939,N_4599);
nand U9862 (N_9862,N_1269,N_1734);
nand U9863 (N_9863,N_1433,N_1139);
and U9864 (N_9864,N_2176,N_1565);
nand U9865 (N_9865,N_3951,N_114);
nor U9866 (N_9866,N_3084,N_24);
nor U9867 (N_9867,N_4432,N_1383);
xnor U9868 (N_9868,N_1657,N_4962);
and U9869 (N_9869,N_959,N_244);
nand U9870 (N_9870,N_4071,N_810);
and U9871 (N_9871,N_3614,N_3583);
xnor U9872 (N_9872,N_4837,N_2282);
nand U9873 (N_9873,N_1176,N_3018);
or U9874 (N_9874,N_3532,N_4988);
or U9875 (N_9875,N_4134,N_2907);
or U9876 (N_9876,N_3645,N_4740);
or U9877 (N_9877,N_2530,N_4215);
and U9878 (N_9878,N_248,N_4252);
or U9879 (N_9879,N_495,N_4554);
xor U9880 (N_9880,N_4413,N_162);
nand U9881 (N_9881,N_3602,N_3135);
and U9882 (N_9882,N_4490,N_1286);
nor U9883 (N_9883,N_860,N_1814);
or U9884 (N_9884,N_3730,N_3197);
nand U9885 (N_9885,N_1699,N_355);
nand U9886 (N_9886,N_2968,N_749);
or U9887 (N_9887,N_3799,N_4718);
nand U9888 (N_9888,N_3549,N_3765);
nor U9889 (N_9889,N_3842,N_3300);
nand U9890 (N_9890,N_4011,N_452);
or U9891 (N_9891,N_1259,N_3986);
nor U9892 (N_9892,N_4844,N_3343);
and U9893 (N_9893,N_509,N_393);
nor U9894 (N_9894,N_2518,N_1206);
xor U9895 (N_9895,N_3442,N_1688);
nor U9896 (N_9896,N_3498,N_1973);
and U9897 (N_9897,N_4275,N_2433);
and U9898 (N_9898,N_3270,N_1642);
and U9899 (N_9899,N_3722,N_3915);
and U9900 (N_9900,N_131,N_3430);
nand U9901 (N_9901,N_470,N_650);
or U9902 (N_9902,N_3771,N_1267);
nand U9903 (N_9903,N_4371,N_2855);
nand U9904 (N_9904,N_4951,N_4333);
nand U9905 (N_9905,N_2371,N_2092);
or U9906 (N_9906,N_2874,N_2271);
nand U9907 (N_9907,N_2097,N_3135);
nor U9908 (N_9908,N_537,N_253);
nor U9909 (N_9909,N_14,N_4428);
or U9910 (N_9910,N_2370,N_2475);
nand U9911 (N_9911,N_1065,N_2187);
and U9912 (N_9912,N_3040,N_3566);
nand U9913 (N_9913,N_2696,N_3675);
or U9914 (N_9914,N_3450,N_4970);
nor U9915 (N_9915,N_158,N_2714);
and U9916 (N_9916,N_4940,N_3157);
or U9917 (N_9917,N_2982,N_4850);
and U9918 (N_9918,N_2087,N_66);
nor U9919 (N_9919,N_825,N_4510);
xor U9920 (N_9920,N_1694,N_732);
and U9921 (N_9921,N_4703,N_3160);
and U9922 (N_9922,N_4625,N_2225);
or U9923 (N_9923,N_3456,N_4563);
nand U9924 (N_9924,N_4475,N_1700);
xor U9925 (N_9925,N_4259,N_4130);
nand U9926 (N_9926,N_1836,N_1891);
nor U9927 (N_9927,N_3099,N_2645);
nand U9928 (N_9928,N_2251,N_4181);
and U9929 (N_9929,N_1312,N_3094);
nand U9930 (N_9930,N_4628,N_2985);
nand U9931 (N_9931,N_4342,N_398);
nor U9932 (N_9932,N_4064,N_785);
or U9933 (N_9933,N_3478,N_3508);
nand U9934 (N_9934,N_1456,N_4523);
nand U9935 (N_9935,N_4113,N_428);
and U9936 (N_9936,N_2770,N_3336);
nor U9937 (N_9937,N_3928,N_2301);
nor U9938 (N_9938,N_1127,N_1066);
nor U9939 (N_9939,N_652,N_3122);
nor U9940 (N_9940,N_370,N_4437);
nor U9941 (N_9941,N_4598,N_83);
nand U9942 (N_9942,N_4479,N_1244);
nor U9943 (N_9943,N_2649,N_843);
or U9944 (N_9944,N_2454,N_3369);
and U9945 (N_9945,N_1059,N_4679);
nor U9946 (N_9946,N_4821,N_4150);
xnor U9947 (N_9947,N_1912,N_3649);
or U9948 (N_9948,N_1758,N_3000);
or U9949 (N_9949,N_3581,N_3544);
xor U9950 (N_9950,N_287,N_4985);
or U9951 (N_9951,N_4749,N_2470);
or U9952 (N_9952,N_4173,N_2441);
nand U9953 (N_9953,N_4152,N_3033);
or U9954 (N_9954,N_4570,N_1385);
nor U9955 (N_9955,N_1319,N_3695);
and U9956 (N_9956,N_3726,N_1270);
and U9957 (N_9957,N_1602,N_1357);
nor U9958 (N_9958,N_3319,N_2736);
nand U9959 (N_9959,N_3077,N_458);
nand U9960 (N_9960,N_2407,N_4385);
and U9961 (N_9961,N_3745,N_652);
or U9962 (N_9962,N_2441,N_3069);
xor U9963 (N_9963,N_4253,N_552);
nor U9964 (N_9964,N_35,N_3480);
or U9965 (N_9965,N_4718,N_907);
and U9966 (N_9966,N_207,N_1278);
nand U9967 (N_9967,N_1378,N_43);
nor U9968 (N_9968,N_4692,N_882);
nor U9969 (N_9969,N_2136,N_4722);
or U9970 (N_9970,N_3191,N_4474);
or U9971 (N_9971,N_2431,N_1144);
nor U9972 (N_9972,N_902,N_228);
or U9973 (N_9973,N_2700,N_768);
nor U9974 (N_9974,N_4001,N_2924);
nand U9975 (N_9975,N_2480,N_4157);
nand U9976 (N_9976,N_4074,N_4859);
and U9977 (N_9977,N_21,N_1398);
nand U9978 (N_9978,N_2140,N_2636);
nor U9979 (N_9979,N_2282,N_4354);
or U9980 (N_9980,N_3406,N_1976);
and U9981 (N_9981,N_1431,N_1644);
or U9982 (N_9982,N_167,N_1227);
and U9983 (N_9983,N_1603,N_4400);
and U9984 (N_9984,N_171,N_4500);
nand U9985 (N_9985,N_1052,N_4323);
or U9986 (N_9986,N_2895,N_4755);
xnor U9987 (N_9987,N_2486,N_1816);
nand U9988 (N_9988,N_1815,N_2406);
or U9989 (N_9989,N_4028,N_4889);
and U9990 (N_9990,N_1405,N_716);
or U9991 (N_9991,N_2226,N_3415);
nor U9992 (N_9992,N_3443,N_2523);
nand U9993 (N_9993,N_2591,N_3583);
nor U9994 (N_9994,N_1718,N_4356);
or U9995 (N_9995,N_589,N_2550);
and U9996 (N_9996,N_2237,N_1878);
xnor U9997 (N_9997,N_3198,N_3418);
and U9998 (N_9998,N_1696,N_4386);
nor U9999 (N_9999,N_576,N_714);
nand U10000 (N_10000,N_9121,N_5658);
or U10001 (N_10001,N_7443,N_9340);
xnor U10002 (N_10002,N_6666,N_8096);
or U10003 (N_10003,N_9600,N_6803);
or U10004 (N_10004,N_5892,N_9046);
nor U10005 (N_10005,N_8535,N_7576);
nand U10006 (N_10006,N_7411,N_8059);
and U10007 (N_10007,N_6584,N_8428);
or U10008 (N_10008,N_7047,N_5619);
nand U10009 (N_10009,N_7695,N_9903);
and U10010 (N_10010,N_8087,N_5463);
xnor U10011 (N_10011,N_9495,N_5546);
or U10012 (N_10012,N_9252,N_6651);
or U10013 (N_10013,N_7090,N_8607);
or U10014 (N_10014,N_5062,N_9801);
and U10015 (N_10015,N_9517,N_5755);
nor U10016 (N_10016,N_9604,N_9124);
or U10017 (N_10017,N_7463,N_8361);
nand U10018 (N_10018,N_5814,N_7597);
or U10019 (N_10019,N_7376,N_7113);
nand U10020 (N_10020,N_9730,N_7383);
or U10021 (N_10021,N_5374,N_6608);
and U10022 (N_10022,N_8606,N_5567);
nor U10023 (N_10023,N_6984,N_9746);
or U10024 (N_10024,N_7401,N_6829);
nand U10025 (N_10025,N_8523,N_9872);
nor U10026 (N_10026,N_8730,N_7241);
nor U10027 (N_10027,N_9650,N_7628);
and U10028 (N_10028,N_7889,N_5236);
or U10029 (N_10029,N_6824,N_9159);
nor U10030 (N_10030,N_5703,N_9295);
or U10031 (N_10031,N_8734,N_9427);
or U10032 (N_10032,N_9097,N_9843);
nor U10033 (N_10033,N_6508,N_6444);
and U10034 (N_10034,N_6971,N_8802);
and U10035 (N_10035,N_6115,N_6462);
or U10036 (N_10036,N_7467,N_7344);
nand U10037 (N_10037,N_9363,N_8633);
and U10038 (N_10038,N_9163,N_7537);
or U10039 (N_10039,N_5327,N_5110);
nor U10040 (N_10040,N_6669,N_6967);
and U10041 (N_10041,N_8954,N_5121);
and U10042 (N_10042,N_5444,N_8638);
nor U10043 (N_10043,N_7130,N_9251);
or U10044 (N_10044,N_6946,N_7895);
nand U10045 (N_10045,N_8257,N_9615);
nor U10046 (N_10046,N_7894,N_6964);
nor U10047 (N_10047,N_6606,N_7266);
nand U10048 (N_10048,N_9051,N_7201);
or U10049 (N_10049,N_5272,N_7722);
nor U10050 (N_10050,N_7534,N_8726);
xnor U10051 (N_10051,N_7669,N_7989);
xnor U10052 (N_10052,N_6996,N_7002);
nor U10053 (N_10053,N_8360,N_8993);
or U10054 (N_10054,N_9726,N_9132);
or U10055 (N_10055,N_9911,N_5557);
or U10056 (N_10056,N_5773,N_7625);
nand U10057 (N_10057,N_8975,N_6215);
nor U10058 (N_10058,N_7461,N_9940);
and U10059 (N_10059,N_6063,N_5894);
nand U10060 (N_10060,N_9313,N_9620);
nor U10061 (N_10061,N_6693,N_6661);
nor U10062 (N_10062,N_5537,N_6092);
xor U10063 (N_10063,N_7439,N_8671);
or U10064 (N_10064,N_5378,N_9575);
and U10065 (N_10065,N_9810,N_5438);
nor U10066 (N_10066,N_5138,N_8787);
and U10067 (N_10067,N_8599,N_7585);
or U10068 (N_10068,N_7706,N_8461);
nor U10069 (N_10069,N_9795,N_6592);
nand U10070 (N_10070,N_8981,N_6286);
and U10071 (N_10071,N_6079,N_6764);
nand U10072 (N_10072,N_5606,N_7063);
nor U10073 (N_10073,N_8171,N_8422);
nand U10074 (N_10074,N_7984,N_5257);
and U10075 (N_10075,N_9497,N_8868);
and U10076 (N_10076,N_7572,N_9745);
nand U10077 (N_10077,N_8340,N_5972);
nor U10078 (N_10078,N_9640,N_6474);
xnor U10079 (N_10079,N_8610,N_6129);
and U10080 (N_10080,N_7492,N_6894);
and U10081 (N_10081,N_9212,N_9174);
or U10082 (N_10082,N_9892,N_5761);
or U10083 (N_10083,N_8399,N_6436);
nand U10084 (N_10084,N_8534,N_6516);
or U10085 (N_10085,N_5441,N_5298);
nor U10086 (N_10086,N_5900,N_7213);
nor U10087 (N_10087,N_5700,N_9529);
nand U10088 (N_10088,N_7876,N_6380);
or U10089 (N_10089,N_8646,N_5399);
nor U10090 (N_10090,N_6117,N_9400);
or U10091 (N_10091,N_5548,N_5277);
nand U10092 (N_10092,N_9564,N_7645);
or U10093 (N_10093,N_8500,N_9868);
or U10094 (N_10094,N_9963,N_7678);
nor U10095 (N_10095,N_6571,N_9602);
nand U10096 (N_10096,N_9853,N_8942);
nand U10097 (N_10097,N_6817,N_7565);
or U10098 (N_10098,N_5230,N_9239);
or U10099 (N_10099,N_6968,N_7956);
xor U10100 (N_10100,N_9469,N_6379);
nand U10101 (N_10101,N_7041,N_8409);
or U10102 (N_10102,N_9571,N_6952);
nand U10103 (N_10103,N_7126,N_5018);
xnor U10104 (N_10104,N_8652,N_6249);
nand U10105 (N_10105,N_7745,N_5917);
xor U10106 (N_10106,N_7407,N_5304);
or U10107 (N_10107,N_7164,N_6056);
or U10108 (N_10108,N_7215,N_6480);
nor U10109 (N_10109,N_9583,N_7869);
xnor U10110 (N_10110,N_6231,N_6599);
nand U10111 (N_10111,N_9009,N_9706);
and U10112 (N_10112,N_5223,N_5310);
or U10113 (N_10113,N_5100,N_5586);
nand U10114 (N_10114,N_5642,N_9857);
or U10115 (N_10115,N_6048,N_9769);
or U10116 (N_10116,N_8886,N_7342);
and U10117 (N_10117,N_8751,N_5422);
or U10118 (N_10118,N_5930,N_6538);
nand U10119 (N_10119,N_8386,N_5860);
nor U10120 (N_10120,N_8163,N_5686);
or U10121 (N_10121,N_7018,N_9783);
or U10122 (N_10122,N_7781,N_8739);
nand U10123 (N_10123,N_7615,N_9950);
or U10124 (N_10124,N_6326,N_5580);
nor U10125 (N_10125,N_7578,N_9173);
nor U10126 (N_10126,N_7371,N_8401);
nor U10127 (N_10127,N_9765,N_9542);
xor U10128 (N_10128,N_6321,N_5987);
nand U10129 (N_10129,N_6161,N_9737);
and U10130 (N_10130,N_6526,N_8898);
nand U10131 (N_10131,N_6145,N_6642);
nand U10132 (N_10132,N_9433,N_8324);
nand U10133 (N_10133,N_7767,N_6674);
nor U10134 (N_10134,N_7449,N_6522);
nor U10135 (N_10135,N_9064,N_5626);
xor U10136 (N_10136,N_9019,N_8063);
and U10137 (N_10137,N_5093,N_8547);
and U10138 (N_10138,N_9000,N_9189);
nor U10139 (N_10139,N_7805,N_7554);
and U10140 (N_10140,N_6871,N_8336);
and U10141 (N_10141,N_9597,N_8771);
xnor U10142 (N_10142,N_9557,N_5063);
nor U10143 (N_10143,N_5662,N_6327);
or U10144 (N_10144,N_5682,N_6768);
or U10145 (N_10145,N_6421,N_6104);
xnor U10146 (N_10146,N_6080,N_7623);
and U10147 (N_10147,N_5565,N_7389);
nor U10148 (N_10148,N_7286,N_8541);
or U10149 (N_10149,N_8425,N_6368);
nand U10150 (N_10150,N_6409,N_7274);
nor U10151 (N_10151,N_9405,N_7234);
nand U10152 (N_10152,N_9191,N_8165);
or U10153 (N_10153,N_8433,N_6266);
or U10154 (N_10154,N_6841,N_9863);
xor U10155 (N_10155,N_8432,N_5324);
nand U10156 (N_10156,N_9120,N_9490);
and U10157 (N_10157,N_5156,N_8838);
or U10158 (N_10158,N_9739,N_8764);
nand U10159 (N_10159,N_5307,N_9105);
nor U10160 (N_10160,N_7135,N_8892);
and U10161 (N_10161,N_6398,N_7074);
or U10162 (N_10162,N_9807,N_8497);
xnor U10163 (N_10163,N_9154,N_8840);
and U10164 (N_10164,N_7363,N_9976);
and U10165 (N_10165,N_6396,N_5424);
xor U10166 (N_10166,N_6430,N_6188);
and U10167 (N_10167,N_6448,N_9435);
or U10168 (N_10168,N_9862,N_7847);
nor U10169 (N_10169,N_9088,N_7823);
or U10170 (N_10170,N_9354,N_6366);
and U10171 (N_10171,N_8965,N_5340);
and U10172 (N_10172,N_8183,N_7990);
nand U10173 (N_10173,N_5620,N_6856);
nand U10174 (N_10174,N_8142,N_9869);
nand U10175 (N_10175,N_6918,N_7832);
nor U10176 (N_10176,N_6323,N_6741);
nand U10177 (N_10177,N_9358,N_8265);
and U10178 (N_10178,N_6844,N_9210);
nand U10179 (N_10179,N_5633,N_5437);
and U10180 (N_10180,N_7302,N_6002);
or U10181 (N_10181,N_9279,N_8385);
and U10182 (N_10182,N_7038,N_5410);
nand U10183 (N_10183,N_8192,N_5800);
nor U10184 (N_10184,N_6458,N_5820);
nor U10185 (N_10185,N_5713,N_8139);
nor U10186 (N_10186,N_6122,N_8679);
or U10187 (N_10187,N_8862,N_7983);
nand U10188 (N_10188,N_6032,N_7151);
nor U10189 (N_10189,N_7907,N_5060);
nor U10190 (N_10190,N_5585,N_8978);
and U10191 (N_10191,N_5885,N_9042);
xor U10192 (N_10192,N_5980,N_7644);
nor U10193 (N_10193,N_7854,N_8817);
and U10194 (N_10194,N_9790,N_7473);
and U10195 (N_10195,N_7023,N_7934);
and U10196 (N_10196,N_9499,N_7009);
and U10197 (N_10197,N_7691,N_6437);
nand U10198 (N_10198,N_7616,N_9933);
xor U10199 (N_10199,N_5690,N_5041);
nor U10200 (N_10200,N_8143,N_8395);
and U10201 (N_10201,N_5080,N_6037);
nand U10202 (N_10202,N_7109,N_9375);
nor U10203 (N_10203,N_8448,N_9621);
nor U10204 (N_10204,N_6251,N_5765);
xnor U10205 (N_10205,N_9696,N_9095);
nand U10206 (N_10206,N_7161,N_5948);
nor U10207 (N_10207,N_5837,N_6465);
nand U10208 (N_10208,N_9603,N_8666);
nor U10209 (N_10209,N_5570,N_7702);
nor U10210 (N_10210,N_5815,N_9909);
nand U10211 (N_10211,N_9357,N_6673);
and U10212 (N_10212,N_8016,N_9574);
or U10213 (N_10213,N_9618,N_8267);
nor U10214 (N_10214,N_7501,N_9260);
nand U10215 (N_10215,N_5017,N_9293);
or U10216 (N_10216,N_5213,N_7533);
or U10217 (N_10217,N_5808,N_6356);
or U10218 (N_10218,N_8998,N_7558);
nand U10219 (N_10219,N_7422,N_6210);
or U10220 (N_10220,N_6186,N_8130);
nand U10221 (N_10221,N_9970,N_9187);
nand U10222 (N_10222,N_6410,N_6101);
nand U10223 (N_10223,N_9034,N_7082);
or U10224 (N_10224,N_5641,N_8443);
nor U10225 (N_10225,N_6176,N_6858);
and U10226 (N_10226,N_6505,N_6887);
nand U10227 (N_10227,N_9073,N_5650);
or U10228 (N_10228,N_9102,N_9185);
and U10229 (N_10229,N_7667,N_8634);
nand U10230 (N_10230,N_9249,N_7536);
nand U10231 (N_10231,N_7535,N_6730);
nand U10232 (N_10232,N_7765,N_9014);
nand U10233 (N_10233,N_6974,N_5443);
or U10234 (N_10234,N_5912,N_9192);
and U10235 (N_10235,N_9043,N_6011);
and U10236 (N_10236,N_5893,N_5037);
or U10237 (N_10237,N_7887,N_7177);
nand U10238 (N_10238,N_5043,N_6100);
nor U10239 (N_10239,N_5189,N_8974);
nor U10240 (N_10240,N_7693,N_6959);
or U10241 (N_10241,N_8774,N_5668);
nor U10242 (N_10242,N_5931,N_8036);
or U10243 (N_10243,N_7881,N_9084);
and U10244 (N_10244,N_5175,N_7620);
or U10245 (N_10245,N_7013,N_5589);
or U10246 (N_10246,N_9425,N_7060);
and U10247 (N_10247,N_9733,N_9563);
and U10248 (N_10248,N_5745,N_6120);
nand U10249 (N_10249,N_8293,N_6752);
or U10250 (N_10250,N_8184,N_5433);
nand U10251 (N_10251,N_9871,N_9415);
nand U10252 (N_10252,N_9325,N_9076);
xnor U10253 (N_10253,N_7520,N_7970);
or U10254 (N_10254,N_8961,N_9685);
nor U10255 (N_10255,N_7316,N_9642);
nor U10256 (N_10256,N_5095,N_5924);
or U10257 (N_10257,N_9462,N_5042);
and U10258 (N_10258,N_6236,N_8731);
or U10259 (N_10259,N_7836,N_7381);
and U10260 (N_10260,N_8587,N_7602);
and U10261 (N_10261,N_9989,N_9488);
xor U10262 (N_10262,N_6053,N_5217);
xnor U10263 (N_10263,N_7313,N_6413);
nor U10264 (N_10264,N_5986,N_9480);
nor U10265 (N_10265,N_9553,N_9297);
nor U10266 (N_10266,N_9244,N_9952);
and U10267 (N_10267,N_7944,N_7664);
nand U10268 (N_10268,N_8876,N_5036);
xnor U10269 (N_10269,N_8746,N_6914);
or U10270 (N_10270,N_6006,N_9668);
nor U10271 (N_10271,N_7810,N_6611);
xor U10272 (N_10272,N_5556,N_5573);
nand U10273 (N_10273,N_9964,N_6322);
nor U10274 (N_10274,N_6456,N_6027);
or U10275 (N_10275,N_6965,N_7795);
and U10276 (N_10276,N_5376,N_5791);
xor U10277 (N_10277,N_7773,N_7042);
nor U10278 (N_10278,N_8678,N_7006);
and U10279 (N_10279,N_7608,N_7684);
or U10280 (N_10280,N_5144,N_7149);
and U10281 (N_10281,N_8176,N_6239);
nand U10282 (N_10282,N_7415,N_9516);
nor U10283 (N_10283,N_5993,N_7140);
and U10284 (N_10284,N_5717,N_8147);
and U10285 (N_10285,N_5430,N_5191);
and U10286 (N_10286,N_7392,N_6167);
or U10287 (N_10287,N_5311,N_6753);
or U10288 (N_10288,N_9002,N_9356);
and U10289 (N_10289,N_7067,N_9037);
and U10290 (N_10290,N_9712,N_6885);
nand U10291 (N_10291,N_5051,N_5373);
nor U10292 (N_10292,N_7502,N_9478);
xor U10293 (N_10293,N_5178,N_5188);
or U10294 (N_10294,N_5541,N_7262);
nand U10295 (N_10295,N_7900,N_8806);
nor U10296 (N_10296,N_5563,N_9158);
or U10297 (N_10297,N_9925,N_8614);
and U10298 (N_10298,N_6043,N_7996);
nand U10299 (N_10299,N_6739,N_5994);
nand U10300 (N_10300,N_6232,N_7249);
or U10301 (N_10301,N_8513,N_8322);
nand U10302 (N_10302,N_6678,N_7146);
and U10303 (N_10303,N_6684,N_6221);
nand U10304 (N_10304,N_9001,N_9673);
nor U10305 (N_10305,N_8721,N_8134);
and U10306 (N_10306,N_9866,N_6487);
and U10307 (N_10307,N_6285,N_5957);
or U10308 (N_10308,N_6041,N_8732);
nor U10309 (N_10309,N_9110,N_9893);
and U10310 (N_10310,N_7864,N_9011);
and U10311 (N_10311,N_5243,N_9704);
or U10312 (N_10312,N_5052,N_8278);
nand U10313 (N_10313,N_8249,N_6438);
and U10314 (N_10314,N_7959,N_8420);
nand U10315 (N_10315,N_7681,N_6718);
nand U10316 (N_10316,N_8514,N_5528);
xnor U10317 (N_10317,N_7486,N_8826);
nand U10318 (N_10318,N_7911,N_7718);
nand U10319 (N_10319,N_8430,N_8054);
nor U10320 (N_10320,N_7081,N_5698);
nand U10321 (N_10321,N_8262,N_6537);
nor U10322 (N_10322,N_5952,N_8571);
nand U10323 (N_10323,N_8531,N_5780);
nor U10324 (N_10324,N_7890,N_8704);
nand U10325 (N_10325,N_6158,N_6524);
and U10326 (N_10326,N_5498,N_5325);
or U10327 (N_10327,N_5462,N_9694);
or U10328 (N_10328,N_8067,N_6951);
nand U10329 (N_10329,N_8848,N_9116);
nor U10330 (N_10330,N_6300,N_7357);
and U10331 (N_10331,N_5360,N_7477);
or U10332 (N_10332,N_6575,N_5262);
nor U10333 (N_10333,N_8248,N_7598);
or U10334 (N_10334,N_5148,N_8752);
nor U10335 (N_10335,N_7163,N_7750);
nand U10336 (N_10336,N_7282,N_8077);
nand U10337 (N_10337,N_7657,N_9459);
nand U10338 (N_10338,N_7778,N_5855);
and U10339 (N_10339,N_5845,N_9364);
and U10340 (N_10340,N_7001,N_7325);
and U10341 (N_10341,N_7014,N_7402);
nand U10342 (N_10342,N_6010,N_5558);
nor U10343 (N_10343,N_6907,N_6633);
nand U10344 (N_10344,N_8814,N_9859);
nor U10345 (N_10345,N_7057,N_5264);
or U10346 (N_10346,N_6415,N_6828);
nand U10347 (N_10347,N_9355,N_7464);
nand U10348 (N_10348,N_6758,N_8072);
nor U10349 (N_10349,N_6573,N_8894);
nor U10350 (N_10350,N_6531,N_6510);
nor U10351 (N_10351,N_9498,N_9389);
or U10352 (N_10352,N_7721,N_5335);
or U10353 (N_10353,N_5237,N_7043);
nand U10354 (N_10354,N_6111,N_9629);
nor U10355 (N_10355,N_8622,N_6755);
nand U10356 (N_10356,N_6066,N_8877);
or U10357 (N_10357,N_7749,N_8872);
and U10358 (N_10358,N_5027,N_5165);
or U10359 (N_10359,N_5807,N_6688);
nand U10360 (N_10360,N_5390,N_8237);
nand U10361 (N_10361,N_7328,N_8778);
and U10362 (N_10362,N_9331,N_8925);
or U10363 (N_10363,N_7817,N_5081);
nand U10364 (N_10364,N_9987,N_6605);
xor U10365 (N_10365,N_8818,N_7731);
nor U10366 (N_10366,N_5830,N_7539);
nand U10367 (N_10367,N_7430,N_9670);
nand U10368 (N_10368,N_8266,N_5181);
nand U10369 (N_10369,N_5946,N_7931);
nand U10370 (N_10370,N_9554,N_9020);
or U10371 (N_10371,N_7878,N_9350);
nor U10372 (N_10372,N_5829,N_7727);
and U10373 (N_10373,N_6785,N_8719);
and U10374 (N_10374,N_8781,N_5754);
nand U10375 (N_10375,N_5832,N_9840);
or U10376 (N_10376,N_7480,N_6625);
or U10377 (N_10377,N_5786,N_8871);
or U10378 (N_10378,N_7021,N_8844);
and U10379 (N_10379,N_8651,N_6915);
nand U10380 (N_10380,N_5884,N_5870);
nand U10381 (N_10381,N_6963,N_6941);
and U10382 (N_10382,N_7076,N_8010);
or U10383 (N_10383,N_8899,N_8645);
nor U10384 (N_10384,N_6767,N_6036);
or U10385 (N_10385,N_7757,N_6149);
or U10386 (N_10386,N_8929,N_5802);
or U10387 (N_10387,N_8594,N_6019);
and U10388 (N_10388,N_8517,N_6093);
or U10389 (N_10389,N_8109,N_5566);
nor U10390 (N_10390,N_5320,N_6384);
nor U10391 (N_10391,N_8103,N_9703);
nor U10392 (N_10392,N_9936,N_7115);
or U10393 (N_10393,N_6013,N_8129);
xnor U10394 (N_10394,N_5420,N_5076);
and U10395 (N_10395,N_7378,N_6742);
or U10396 (N_10396,N_9953,N_9521);
and U10397 (N_10397,N_5219,N_5628);
or U10398 (N_10398,N_9537,N_9788);
nor U10399 (N_10399,N_5742,N_8735);
or U10400 (N_10400,N_8714,N_9981);
or U10401 (N_10401,N_5218,N_8186);
nor U10402 (N_10402,N_9791,N_9077);
nand U10403 (N_10403,N_7816,N_9570);
or U10404 (N_10404,N_7362,N_5798);
nor U10405 (N_10405,N_5479,N_7515);
nor U10406 (N_10406,N_5795,N_9416);
and U10407 (N_10407,N_8026,N_8480);
and U10408 (N_10408,N_6426,N_9535);
nand U10409 (N_10409,N_6391,N_6819);
nor U10410 (N_10410,N_7094,N_7396);
and U10411 (N_10411,N_7677,N_6948);
nor U10412 (N_10412,N_5260,N_8455);
xnor U10413 (N_10413,N_8776,N_8354);
nand U10414 (N_10414,N_9927,N_6827);
or U10415 (N_10415,N_5848,N_9023);
nand U10416 (N_10416,N_6141,N_8426);
or U10417 (N_10417,N_5029,N_5920);
nor U10418 (N_10418,N_7049,N_9320);
or U10419 (N_10419,N_6703,N_8987);
nor U10420 (N_10420,N_9594,N_5550);
nand U10421 (N_10421,N_6071,N_9311);
nand U10422 (N_10422,N_5590,N_9216);
or U10423 (N_10423,N_7438,N_7085);
nor U10424 (N_10424,N_7545,N_5512);
nand U10425 (N_10425,N_7360,N_6033);
nor U10426 (N_10426,N_7519,N_8117);
and U10427 (N_10427,N_8672,N_7860);
nor U10428 (N_10428,N_9306,N_9348);
nand U10429 (N_10429,N_7101,N_8860);
and U10430 (N_10430,N_8973,N_7237);
or U10431 (N_10431,N_8081,N_8511);
nor U10432 (N_10432,N_8417,N_5197);
and U10433 (N_10433,N_9487,N_6750);
xor U10434 (N_10434,N_9017,N_6256);
nor U10435 (N_10435,N_5890,N_6960);
xor U10436 (N_10436,N_6357,N_5105);
nand U10437 (N_10437,N_6657,N_9214);
nor U10438 (N_10438,N_9441,N_7924);
xnor U10439 (N_10439,N_8613,N_6497);
and U10440 (N_10440,N_8619,N_7525);
nor U10441 (N_10441,N_5921,N_9901);
nand U10442 (N_10442,N_9898,N_7037);
nand U10443 (N_10443,N_8995,N_8926);
nor U10444 (N_10444,N_8024,N_7715);
nor U10445 (N_10445,N_8858,N_8585);
and U10446 (N_10446,N_5804,N_5889);
or U10447 (N_10447,N_9920,N_8166);
nand U10448 (N_10448,N_7409,N_5851);
and U10449 (N_10449,N_6724,N_6190);
nor U10450 (N_10450,N_8021,N_7334);
and U10451 (N_10451,N_8940,N_5818);
or U10452 (N_10452,N_9420,N_6795);
nand U10453 (N_10453,N_6270,N_7888);
or U10454 (N_10454,N_9395,N_8512);
or U10455 (N_10455,N_5097,N_5710);
nand U10456 (N_10456,N_6875,N_6148);
or U10457 (N_10457,N_8226,N_7447);
or U10458 (N_10458,N_7954,N_8048);
nor U10459 (N_10459,N_7406,N_8621);
nand U10460 (N_10460,N_9267,N_7338);
nand U10461 (N_10461,N_8617,N_8241);
xnor U10462 (N_10462,N_7416,N_9732);
or U10463 (N_10463,N_5024,N_7004);
or U10464 (N_10464,N_6906,N_9772);
or U10465 (N_10465,N_8456,N_5533);
nand U10466 (N_10466,N_6617,N_9681);
and U10467 (N_10467,N_7446,N_8034);
nand U10468 (N_10468,N_5869,N_7379);
nand U10469 (N_10469,N_5640,N_5785);
xor U10470 (N_10470,N_9774,N_6021);
nor U10471 (N_10471,N_9198,N_8675);
nand U10472 (N_10472,N_6893,N_8173);
nor U10473 (N_10473,N_7133,N_5267);
nand U10474 (N_10474,N_8588,N_7943);
and U10475 (N_10475,N_7772,N_6889);
nor U10476 (N_10476,N_7165,N_8145);
and U10477 (N_10477,N_9491,N_6892);
nand U10478 (N_10478,N_9101,N_8641);
or U10479 (N_10479,N_6520,N_7459);
and U10480 (N_10480,N_5778,N_9399);
nor U10481 (N_10481,N_9138,N_7512);
nand U10482 (N_10482,N_5466,N_7180);
and U10483 (N_10483,N_7560,N_5469);
and U10484 (N_10484,N_7828,N_5897);
and U10485 (N_10485,N_9837,N_8841);
nor U10486 (N_10486,N_8558,N_7754);
nor U10487 (N_10487,N_7630,N_6801);
nand U10488 (N_10488,N_6826,N_8687);
xor U10489 (N_10489,N_8032,N_5910);
xor U10490 (N_10490,N_5193,N_5244);
or U10491 (N_10491,N_8039,N_9476);
nor U10492 (N_10492,N_8210,N_9820);
nand U10493 (N_10493,N_8592,N_8174);
nand U10494 (N_10494,N_5607,N_5622);
nor U10495 (N_10495,N_5402,N_6466);
or U10496 (N_10496,N_7619,N_9429);
xnor U10497 (N_10497,N_5248,N_5015);
xor U10498 (N_10498,N_5667,N_6776);
and U10499 (N_10499,N_6782,N_5927);
or U10500 (N_10500,N_9265,N_9309);
nor U10501 (N_10501,N_8252,N_5699);
or U10502 (N_10502,N_8479,N_9304);
nor U10503 (N_10503,N_8126,N_9735);
or U10504 (N_10504,N_7910,N_6902);
or U10505 (N_10505,N_9514,N_7730);
or U10506 (N_10506,N_8969,N_8794);
nor U10507 (N_10507,N_9691,N_6314);
nand U10508 (N_10508,N_7185,N_9287);
and U10509 (N_10509,N_8955,N_8028);
nor U10510 (N_10510,N_5693,N_7641);
and U10511 (N_10511,N_8037,N_9305);
and U10512 (N_10512,N_8911,N_9928);
or U10513 (N_10513,N_9748,N_8712);
and U10514 (N_10514,N_5407,N_6973);
xnor U10515 (N_10515,N_6935,N_8156);
and U10516 (N_10516,N_7867,N_7909);
and U10517 (N_10517,N_6351,N_6763);
nand U10518 (N_10518,N_5679,N_8316);
nand U10519 (N_10519,N_9995,N_9028);
and U10520 (N_10520,N_9882,N_5751);
and U10521 (N_10521,N_6586,N_6796);
and U10522 (N_10522,N_9687,N_7839);
and U10523 (N_10523,N_6185,N_8753);
and U10524 (N_10524,N_9858,N_8582);
nor U10525 (N_10525,N_9572,N_5152);
or U10526 (N_10526,N_7264,N_5337);
or U10527 (N_10527,N_7963,N_7245);
and U10528 (N_10528,N_6252,N_7420);
nor U10529 (N_10529,N_7574,N_8280);
nand U10530 (N_10530,N_9232,N_7656);
nand U10531 (N_10531,N_8356,N_9635);
or U10532 (N_10532,N_9654,N_6942);
nand U10533 (N_10533,N_7892,N_8348);
nand U10534 (N_10534,N_9272,N_9506);
or U10535 (N_10535,N_8355,N_9947);
nand U10536 (N_10536,N_7927,N_9453);
xor U10537 (N_10537,N_7550,N_5734);
or U10538 (N_10538,N_6435,N_9261);
and U10539 (N_10539,N_9494,N_7327);
nand U10540 (N_10540,N_7882,N_9749);
and U10541 (N_10541,N_5527,N_9247);
nand U10542 (N_10542,N_9758,N_8740);
or U10543 (N_10543,N_9460,N_5935);
xor U10544 (N_10544,N_9122,N_6220);
nor U10545 (N_10545,N_9467,N_6457);
and U10546 (N_10546,N_9850,N_7066);
and U10547 (N_10547,N_7640,N_7377);
nand U10548 (N_10548,N_6751,N_7526);
and U10549 (N_10549,N_8827,N_7247);
nand U10550 (N_10550,N_6123,N_7248);
xnor U10551 (N_10551,N_8550,N_8082);
and U10552 (N_10552,N_6070,N_5465);
nor U10553 (N_10553,N_9513,N_8100);
nand U10554 (N_10554,N_8928,N_9273);
and U10555 (N_10555,N_8365,N_9446);
nand U10556 (N_10556,N_7462,N_9581);
or U10557 (N_10557,N_5266,N_7766);
and U10558 (N_10558,N_6088,N_7712);
nor U10559 (N_10559,N_9802,N_6132);
and U10560 (N_10560,N_5453,N_9372);
nor U10561 (N_10561,N_5711,N_7981);
nor U10562 (N_10562,N_5284,N_8887);
or U10563 (N_10563,N_6569,N_9576);
nand U10564 (N_10564,N_5261,N_9886);
nor U10565 (N_10565,N_6588,N_8364);
or U10566 (N_10566,N_8821,N_8083);
or U10567 (N_10567,N_5398,N_6969);
nand U10568 (N_10568,N_9870,N_7064);
or U10569 (N_10569,N_6057,N_7150);
nand U10570 (N_10570,N_8389,N_8854);
nand U10571 (N_10571,N_5221,N_7364);
xnor U10572 (N_10572,N_6955,N_5123);
nand U10573 (N_10573,N_8206,N_7777);
nand U10574 (N_10574,N_8391,N_7744);
and U10575 (N_10575,N_9103,N_5631);
or U10576 (N_10576,N_6094,N_8490);
and U10577 (N_10577,N_5083,N_6151);
or U10578 (N_10578,N_9710,N_6540);
or U10579 (N_10579,N_8539,N_5281);
nor U10580 (N_10580,N_9148,N_9151);
nor U10581 (N_10581,N_9968,N_8378);
or U10582 (N_10582,N_9983,N_9692);
or U10583 (N_10583,N_6392,N_6985);
and U10584 (N_10584,N_5763,N_8482);
or U10585 (N_10585,N_9534,N_7780);
and U10586 (N_10586,N_5998,N_9456);
or U10587 (N_10587,N_5947,N_5678);
and U10588 (N_10588,N_8832,N_8813);
nand U10589 (N_10589,N_7472,N_8901);
or U10590 (N_10590,N_9024,N_5823);
or U10591 (N_10591,N_9775,N_8935);
nand U10592 (N_10592,N_7005,N_7969);
nor U10593 (N_10593,N_9319,N_6572);
nor U10594 (N_10594,N_8201,N_8392);
nand U10595 (N_10595,N_8367,N_8467);
nand U10596 (N_10596,N_9130,N_8457);
xnor U10597 (N_10597,N_6972,N_6098);
or U10598 (N_10598,N_5824,N_9152);
or U10599 (N_10599,N_9721,N_9268);
or U10600 (N_10600,N_6355,N_5587);
and U10601 (N_10601,N_9161,N_8572);
and U10602 (N_10602,N_9326,N_7221);
xor U10603 (N_10603,N_7295,N_8334);
and U10604 (N_10604,N_5155,N_9182);
or U10605 (N_10605,N_9049,N_9894);
nand U10606 (N_10606,N_9167,N_6336);
nand U10607 (N_10607,N_6274,N_9624);
xnor U10608 (N_10608,N_6991,N_6701);
nand U10609 (N_10609,N_7257,N_7813);
nand U10610 (N_10610,N_9891,N_8628);
or U10611 (N_10611,N_6558,N_9264);
and U10612 (N_10612,N_7891,N_9457);
and U10613 (N_10613,N_7095,N_9057);
and U10614 (N_10614,N_8956,N_5560);
xor U10615 (N_10615,N_8586,N_5645);
and U10616 (N_10616,N_8309,N_9330);
or U10617 (N_10617,N_7428,N_9114);
or U10618 (N_10618,N_5396,N_5124);
nand U10619 (N_10619,N_9519,N_9236);
or U10620 (N_10620,N_8211,N_6720);
nor U10621 (N_10621,N_8300,N_8908);
or U10622 (N_10622,N_7450,N_7307);
nand U10623 (N_10623,N_6677,N_6008);
xor U10624 (N_10624,N_7523,N_6280);
nor U10625 (N_10625,N_8435,N_5199);
or U10626 (N_10626,N_9335,N_6282);
and U10627 (N_10627,N_9492,N_9177);
nand U10628 (N_10628,N_8728,N_6883);
nor U10629 (N_10629,N_6848,N_8194);
and U10630 (N_10630,N_7908,N_9369);
and U10631 (N_10631,N_9253,N_9021);
or U10632 (N_10632,N_5934,N_5954);
and U10633 (N_10633,N_6460,N_8382);
xor U10634 (N_10634,N_6483,N_5502);
nor U10635 (N_10635,N_6241,N_6125);
or U10636 (N_10636,N_8664,N_7674);
and U10637 (N_10637,N_9373,N_8312);
nor U10638 (N_10638,N_5813,N_6975);
or U10639 (N_10639,N_7193,N_8717);
nand U10640 (N_10640,N_5484,N_6276);
and U10641 (N_10641,N_8014,N_8444);
and U10642 (N_10642,N_5534,N_6331);
nor U10643 (N_10643,N_9845,N_5482);
and U10644 (N_10644,N_5790,N_5021);
xnor U10645 (N_10645,N_9256,N_6212);
xor U10646 (N_10646,N_6812,N_8834);
xnor U10647 (N_10647,N_8127,N_6277);
nor U10648 (N_10648,N_8476,N_5085);
and U10649 (N_10649,N_9170,N_7849);
nor U10650 (N_10650,N_7125,N_9742);
or U10651 (N_10651,N_8519,N_5545);
or U10652 (N_10652,N_6291,N_9149);
nor U10653 (N_10653,N_7685,N_7884);
or U10654 (N_10654,N_7465,N_7575);
or U10655 (N_10655,N_6956,N_8275);
xor U10656 (N_10656,N_8258,N_7010);
or U10657 (N_10657,N_8372,N_9217);
or U10658 (N_10658,N_7776,N_6077);
or U10659 (N_10659,N_6699,N_9353);
nand U10660 (N_10660,N_5073,N_6075);
and U10661 (N_10661,N_7824,N_8379);
or U10662 (N_10662,N_5660,N_7807);
nand U10663 (N_10663,N_6590,N_9489);
nor U10664 (N_10664,N_6700,N_9698);
or U10665 (N_10665,N_6987,N_7367);
or U10666 (N_10666,N_7559,N_9986);
and U10667 (N_10667,N_9796,N_8358);
nor U10668 (N_10668,N_5833,N_5718);
xnor U10669 (N_10669,N_5819,N_7687);
and U10670 (N_10670,N_9951,N_6174);
nand U10671 (N_10671,N_5704,N_7877);
nor U10672 (N_10672,N_7541,N_6566);
nor U10673 (N_10673,N_8842,N_8296);
and U10674 (N_10674,N_5341,N_6626);
nor U10675 (N_10675,N_5293,N_6648);
or U10676 (N_10676,N_8750,N_8363);
nand U10677 (N_10677,N_8069,N_7859);
xnor U10678 (N_10678,N_5522,N_8164);
nor U10679 (N_10679,N_5300,N_7758);
or U10680 (N_10680,N_6361,N_7434);
nand U10681 (N_10681,N_9835,N_7736);
or U10682 (N_10682,N_5505,N_9966);
xnor U10683 (N_10683,N_7242,N_7636);
and U10684 (N_10684,N_9370,N_9179);
nor U10685 (N_10685,N_5435,N_8503);
or U10686 (N_10686,N_8994,N_8880);
nor U10687 (N_10687,N_6183,N_5624);
nor U10688 (N_10688,N_5369,N_5740);
nor U10689 (N_10689,N_9825,N_5385);
nor U10690 (N_10690,N_6017,N_7284);
or U10691 (N_10691,N_6929,N_8092);
xnor U10692 (N_10692,N_5339,N_6170);
nor U10693 (N_10693,N_8182,N_7114);
nor U10694 (N_10694,N_9376,N_9258);
and U10695 (N_10695,N_6622,N_9345);
and U10696 (N_10696,N_6792,N_5542);
nor U10697 (N_10697,N_7470,N_6719);
or U10698 (N_10698,N_5203,N_7827);
and U10699 (N_10699,N_7782,N_7053);
and U10700 (N_10700,N_9281,N_9780);
and U10701 (N_10701,N_5874,N_7663);
nor U10702 (N_10702,N_6453,N_8720);
and U10703 (N_10703,N_5372,N_9384);
nor U10704 (N_10704,N_9921,N_9455);
xnor U10705 (N_10705,N_5447,N_8041);
xnor U10706 (N_10706,N_8162,N_8376);
or U10707 (N_10707,N_7490,N_6200);
nor U10708 (N_10708,N_7617,N_8875);
nand U10709 (N_10709,N_6610,N_8219);
nor U10710 (N_10710,N_8815,N_6512);
and U10711 (N_10711,N_8900,N_6403);
nand U10712 (N_10712,N_6294,N_7179);
nor U10713 (N_10713,N_9799,N_5737);
and U10714 (N_10714,N_9708,N_5997);
or U10715 (N_10715,N_9510,N_5334);
or U10716 (N_10716,N_6653,N_6364);
xor U10717 (N_10717,N_5368,N_9263);
nand U10718 (N_10718,N_9098,N_5523);
and U10719 (N_10719,N_6087,N_6962);
nor U10720 (N_10720,N_6867,N_9419);
nor U10721 (N_10721,N_9548,N_6908);
or U10722 (N_10722,N_6461,N_9653);
and U10723 (N_10723,N_6770,N_6257);
nor U10724 (N_10724,N_6432,N_6401);
xnor U10725 (N_10725,N_9481,N_5992);
nor U10726 (N_10726,N_7137,N_9522);
nor U10727 (N_10727,N_8798,N_9711);
nand U10728 (N_10728,N_7746,N_7937);
and U10729 (N_10729,N_6723,N_6095);
and U10730 (N_10730,N_7016,N_8536);
nand U10731 (N_10731,N_9552,N_8498);
or U10732 (N_10732,N_9382,N_8057);
nor U10733 (N_10733,N_9162,N_8847);
nand U10734 (N_10734,N_8140,N_9770);
nor U10735 (N_10735,N_8629,N_9689);
nand U10736 (N_10736,N_5349,N_7369);
or U10737 (N_10737,N_8603,N_5359);
nand U10738 (N_10738,N_9631,N_9533);
nand U10739 (N_10739,N_8205,N_5302);
nand U10740 (N_10740,N_6338,N_9463);
and U10741 (N_10741,N_7982,N_5627);
and U10742 (N_10742,N_5245,N_9686);
xnor U10743 (N_10743,N_8650,N_9752);
nor U10744 (N_10744,N_6861,N_9421);
xor U10745 (N_10745,N_8795,N_9381);
or U10746 (N_10746,N_9220,N_6523);
or U10747 (N_10747,N_7848,N_6090);
nor U10748 (N_10748,N_6121,N_8505);
and U10749 (N_10749,N_5480,N_9242);
nor U10750 (N_10750,N_5045,N_7948);
nor U10751 (N_10751,N_6916,N_8377);
xnor U10752 (N_10752,N_7348,N_9632);
xnor U10753 (N_10753,N_7099,N_6855);
and U10754 (N_10754,N_7157,N_6717);
xor U10755 (N_10755,N_7279,N_7468);
nor U10756 (N_10756,N_7609,N_9816);
nor U10757 (N_10757,N_7414,N_6993);
nor U10758 (N_10758,N_8458,N_8649);
nor U10759 (N_10759,N_7408,N_9003);
nand U10760 (N_10760,N_5675,N_7003);
and U10761 (N_10761,N_9137,N_9811);
and U10762 (N_10762,N_8502,N_6822);
and U10763 (N_10763,N_7254,N_9334);
nor U10764 (N_10764,N_6157,N_9079);
nor U10765 (N_10765,N_8927,N_5046);
nand U10766 (N_10766,N_8953,N_5132);
or U10767 (N_10767,N_7170,N_7147);
and U10768 (N_10768,N_5473,N_8369);
and U10769 (N_10769,N_6631,N_5578);
nor U10770 (N_10770,N_8397,N_8351);
or U10771 (N_10771,N_8161,N_6708);
nand U10772 (N_10772,N_6337,N_6542);
nor U10773 (N_10773,N_7903,N_9822);
and U10774 (N_10774,N_7770,N_8313);
nor U10775 (N_10775,N_8091,N_5478);
and U10776 (N_10776,N_8484,N_6900);
xor U10777 (N_10777,N_6307,N_8729);
and U10778 (N_10778,N_8522,N_8786);
and U10779 (N_10779,N_5316,N_9080);
or U10780 (N_10780,N_8980,N_8023);
nand U10781 (N_10781,N_9643,N_7380);
nand U10782 (N_10782,N_8910,N_9906);
nor U10783 (N_10783,N_7372,N_6813);
nand U10784 (N_10784,N_6582,N_7946);
nor U10785 (N_10785,N_7724,N_7240);
nor U10786 (N_10786,N_9226,N_8406);
xnor U10787 (N_10787,N_6811,N_6732);
and U10788 (N_10788,N_8620,N_8870);
nor U10789 (N_10789,N_6756,N_7322);
and U10790 (N_10790,N_9904,N_7263);
nand U10791 (N_10791,N_6888,N_5732);
nand U10792 (N_10792,N_6255,N_7662);
nand U10793 (N_10793,N_7084,N_5028);
or U10794 (N_10794,N_5914,N_8557);
nand U10795 (N_10795,N_7977,N_8328);
or U10796 (N_10796,N_7917,N_8709);
or U10797 (N_10797,N_8495,N_8769);
xnor U10798 (N_10798,N_8035,N_9885);
nor U10799 (N_10799,N_5981,N_7072);
and U10800 (N_10800,N_9215,N_7134);
or U10801 (N_10801,N_7155,N_6377);
and U10802 (N_10802,N_6922,N_9008);
and U10803 (N_10803,N_7755,N_7521);
xor U10804 (N_10804,N_6615,N_9541);
or U10805 (N_10805,N_8170,N_7740);
nor U10806 (N_10806,N_5336,N_5928);
nand U10807 (N_10807,N_9679,N_5853);
nor U10808 (N_10808,N_7935,N_9994);
xnor U10809 (N_10809,N_9972,N_5180);
or U10810 (N_10810,N_5880,N_8080);
or U10811 (N_10811,N_5697,N_6802);
or U10812 (N_10812,N_5695,N_9377);
and U10813 (N_10813,N_6097,N_5071);
and U10814 (N_10814,N_8642,N_9644);
and U10815 (N_10815,N_6535,N_9688);
nand U10816 (N_10816,N_8469,N_5468);
nand U10817 (N_10817,N_6722,N_9666);
and U10818 (N_10818,N_6304,N_8780);
nand U10819 (N_10819,N_8005,N_8255);
nor U10820 (N_10820,N_9282,N_8064);
nor U10821 (N_10821,N_9766,N_5458);
nor U10822 (N_10822,N_7967,N_9299);
nand U10823 (N_10823,N_9543,N_9662);
nor U10824 (N_10824,N_8232,N_5485);
nand U10825 (N_10825,N_9005,N_9619);
and U10826 (N_10826,N_7643,N_9408);
nor U10827 (N_10827,N_7022,N_9196);
nand U10828 (N_10828,N_6054,N_9231);
and U10829 (N_10829,N_5591,N_5065);
and U10830 (N_10830,N_9477,N_5716);
and U10831 (N_10831,N_7083,N_9536);
and U10832 (N_10832,N_8785,N_6731);
or U10833 (N_10833,N_9155,N_5209);
nand U10834 (N_10834,N_6568,N_7920);
nor U10835 (N_10835,N_8180,N_6464);
or U10836 (N_10836,N_6630,N_6716);
or U10837 (N_10837,N_8475,N_5665);
nand U10838 (N_10838,N_9942,N_9136);
nor U10839 (N_10839,N_5552,N_7299);
or U10840 (N_10840,N_5852,N_8703);
or U10841 (N_10841,N_6921,N_8883);
and U10842 (N_10842,N_9329,N_6961);
nand U10843 (N_10843,N_5099,N_5945);
and U10844 (N_10844,N_6830,N_6242);
nor U10845 (N_10845,N_6292,N_7232);
nand U10846 (N_10846,N_6085,N_6570);
or U10847 (N_10847,N_7748,N_6350);
or U10848 (N_10848,N_6533,N_6074);
and U10849 (N_10849,N_6193,N_5531);
or U10850 (N_10850,N_7672,N_8837);
and U10851 (N_10851,N_6905,N_5635);
nand U10852 (N_10852,N_9050,N_6560);
and U10853 (N_10853,N_9479,N_7582);
nor U10854 (N_10854,N_5269,N_7291);
and U10855 (N_10855,N_5383,N_8440);
and U10856 (N_10856,N_5120,N_5600);
nand U10857 (N_10857,N_6517,N_5417);
nand U10858 (N_10858,N_8964,N_9013);
nor U10859 (N_10859,N_8460,N_5781);
and U10860 (N_10860,N_5423,N_7802);
and U10861 (N_10861,N_9086,N_9234);
or U10862 (N_10862,N_9555,N_9744);
nor U10863 (N_10863,N_6515,N_8310);
nor U10864 (N_10864,N_6378,N_7222);
nor U10865 (N_10865,N_8215,N_5268);
and U10866 (N_10866,N_9428,N_8611);
and U10867 (N_10867,N_8724,N_8463);
or U10868 (N_10868,N_7131,N_6139);
nor U10869 (N_10869,N_6496,N_6447);
xnor U10870 (N_10870,N_8970,N_8823);
or U10871 (N_10871,N_9803,N_6406);
or U10872 (N_10872,N_6788,N_8869);
and U10873 (N_10873,N_5895,N_7424);
and U10874 (N_10874,N_9082,N_7162);
nor U10875 (N_10875,N_5170,N_5938);
nor U10876 (N_10876,N_5006,N_9006);
nand U10877 (N_10877,N_5812,N_6052);
and U10878 (N_10878,N_8895,N_8197);
and U10879 (N_10879,N_7187,N_5964);
nor U10880 (N_10880,N_5190,N_6901);
and U10881 (N_10881,N_5741,N_9714);
nand U10882 (N_10882,N_6353,N_5210);
nor U10883 (N_10883,N_8453,N_9797);
nor U10884 (N_10884,N_9181,N_6621);
nand U10885 (N_10885,N_6546,N_8058);
nor U10886 (N_10886,N_8452,N_6192);
nor U10887 (N_10887,N_9166,N_6994);
xnor U10888 (N_10888,N_9647,N_5771);
nand U10889 (N_10889,N_5503,N_8193);
or U10890 (N_10890,N_5318,N_9145);
and U10891 (N_10891,N_8093,N_6073);
nor U10892 (N_10892,N_7595,N_5164);
and U10893 (N_10893,N_6851,N_9307);
nand U10894 (N_10894,N_7280,N_6387);
nand U10895 (N_10895,N_8368,N_6832);
and U10896 (N_10896,N_9842,N_5836);
nand U10897 (N_10897,N_9975,N_7505);
nor U10898 (N_10898,N_5357,N_5403);
nor U10899 (N_10899,N_9768,N_5612);
nand U10900 (N_10900,N_7457,N_7331);
nor U10901 (N_10901,N_6933,N_6498);
nor U10902 (N_10902,N_8345,N_8119);
nand U10903 (N_10903,N_8756,N_5249);
xnor U10904 (N_10904,N_8544,N_6408);
and U10905 (N_10905,N_6857,N_5881);
nor U10906 (N_10906,N_7144,N_6671);
nand U10907 (N_10907,N_8242,N_9627);
nor U10908 (N_10908,N_6479,N_5706);
or U10909 (N_10909,N_5515,N_5902);
and U10910 (N_10910,N_7399,N_8902);
and U10911 (N_10911,N_8615,N_8335);
or U10912 (N_10912,N_6644,N_9411);
nand U10913 (N_10913,N_6038,N_8144);
nand U10914 (N_10914,N_8481,N_6172);
and U10915 (N_10915,N_8264,N_8019);
nor U10916 (N_10916,N_6947,N_9424);
and U10917 (N_10917,N_7862,N_6284);
or U10918 (N_10918,N_8782,N_5953);
xor U10919 (N_10919,N_5883,N_7661);
xor U10920 (N_10920,N_7289,N_9385);
xnor U10921 (N_10921,N_5247,N_8945);
xor U10922 (N_10922,N_5375,N_7606);
nand U10923 (N_10923,N_9846,N_6219);
nor U10924 (N_10924,N_9278,N_5206);
xor U10925 (N_10925,N_6216,N_8631);
nor U10926 (N_10926,N_7797,N_9702);
and U10927 (N_10927,N_6562,N_7425);
or U10928 (N_10928,N_5387,N_9085);
nand U10929 (N_10929,N_6076,N_5632);
nor U10930 (N_10930,N_9406,N_8828);
or U10931 (N_10931,N_7825,N_9777);
or U10932 (N_10932,N_8137,N_7719);
and U10933 (N_10933,N_6445,N_5561);
and U10934 (N_10934,N_6596,N_5140);
xor U10935 (N_10935,N_9074,N_7528);
nand U10936 (N_10936,N_6204,N_6040);
xor U10937 (N_10937,N_9511,N_6715);
nor U10938 (N_10938,N_9454,N_5530);
nor U10939 (N_10939,N_8598,N_8578);
nand U10940 (N_10940,N_7872,N_8321);
nor U10941 (N_10941,N_6676,N_5618);
and U10942 (N_10942,N_9407,N_8716);
xor U10943 (N_10943,N_7479,N_7922);
nand U10944 (N_10944,N_9549,N_5471);
nand U10945 (N_10945,N_7930,N_7929);
or U10946 (N_10946,N_6668,N_5016);
or U10947 (N_10947,N_5308,N_8233);
nor U10948 (N_10948,N_5283,N_6769);
nand U10949 (N_10949,N_9143,N_7793);
nand U10950 (N_10950,N_9100,N_7239);
xnor U10951 (N_10951,N_7236,N_5225);
or U10952 (N_10952,N_9343,N_8859);
and U10953 (N_10953,N_8333,N_8499);
nor U10954 (N_10954,N_5362,N_7775);
xor U10955 (N_10955,N_8464,N_8958);
nor U10956 (N_10956,N_5898,N_8102);
nand U10957 (N_10957,N_5366,N_5661);
nand U10958 (N_10958,N_9945,N_8494);
or U10959 (N_10959,N_7653,N_7974);
xnor U10960 (N_10960,N_7143,N_7205);
or U10961 (N_10961,N_8124,N_6912);
or U10962 (N_10962,N_5228,N_5979);
nand U10963 (N_10963,N_7548,N_5594);
or U10964 (N_10964,N_9365,N_5803);
nor U10965 (N_10965,N_8200,N_7806);
nor U10966 (N_10966,N_6108,N_7812);
and U10967 (N_10967,N_8985,N_5271);
nand U10968 (N_10968,N_6602,N_9684);
nor U10969 (N_10969,N_9342,N_8772);
nor U10970 (N_10970,N_6001,N_9394);
or U10971 (N_10971,N_9473,N_9351);
and U10972 (N_10972,N_8757,N_9030);
or U10973 (N_10973,N_7091,N_6127);
nand U10974 (N_10974,N_5416,N_8566);
nand U10975 (N_10975,N_7216,N_9436);
and U10976 (N_10976,N_6113,N_6799);
nor U10977 (N_10977,N_5822,N_6686);
or U10978 (N_10978,N_8259,N_7349);
nand U10979 (N_10979,N_7660,N_6205);
or U10980 (N_10980,N_8698,N_7985);
xor U10981 (N_10981,N_5776,N_6689);
or U10982 (N_10982,N_7395,N_5192);
nor U10983 (N_10983,N_8864,N_5194);
nor U10984 (N_10984,N_9289,N_7017);
nor U10985 (N_10985,N_6484,N_5371);
nand U10986 (N_10986,N_7330,N_9486);
nand U10987 (N_10987,N_6587,N_7132);
and U10988 (N_10988,N_9482,N_5182);
nand U10989 (N_10989,N_8381,N_5265);
and U10990 (N_10990,N_9889,N_8287);
nand U10991 (N_10991,N_8533,N_7271);
or U10992 (N_10992,N_8670,N_9778);
nand U10993 (N_10993,N_9736,N_7080);
xor U10994 (N_10994,N_6976,N_7044);
or U10995 (N_10995,N_6289,N_9729);
and U10996 (N_10996,N_6529,N_7252);
nor U10997 (N_10997,N_7863,N_5436);
and U10998 (N_10998,N_9109,N_8612);
or U10999 (N_10999,N_8284,N_8167);
or U11000 (N_11000,N_5995,N_7426);
or U11001 (N_11001,N_6287,N_7166);
or U11002 (N_11002,N_6428,N_8966);
nor U11003 (N_11003,N_5577,N_9208);
nor U11004 (N_11004,N_6427,N_8874);
and U11005 (N_11005,N_6009,N_7814);
or U11006 (N_11006,N_7659,N_6998);
or U11007 (N_11007,N_6332,N_7738);
nor U11008 (N_11008,N_5177,N_7139);
or U11009 (N_11009,N_8038,N_9207);
nor U11010 (N_11010,N_6169,N_7329);
and U11011 (N_11011,N_9960,N_9907);
or U11012 (N_11012,N_9332,N_8518);
or U11013 (N_11013,N_6182,N_6275);
xor U11014 (N_11014,N_7522,N_5730);
or U11015 (N_11015,N_6016,N_6203);
or U11016 (N_11016,N_9038,N_9924);
or U11017 (N_11017,N_9387,N_7107);
or U11018 (N_11018,N_6816,N_8933);
nand U11019 (N_11019,N_7586,N_5918);
or U11020 (N_11020,N_8577,N_8225);
and U11021 (N_11021,N_6565,N_5518);
and U11022 (N_11022,N_7476,N_9700);
xnor U11023 (N_11023,N_5034,N_6635);
nor U11024 (N_11024,N_6263,N_9880);
xor U11025 (N_11025,N_9771,N_7158);
or U11026 (N_11026,N_8789,N_7495);
nand U11027 (N_11027,N_5239,N_8168);
and U11028 (N_11028,N_5529,N_9403);
nand U11029 (N_11029,N_8196,N_5520);
xnor U11030 (N_11030,N_8273,N_9682);
and U11031 (N_11031,N_7033,N_5207);
nor U11032 (N_11032,N_6370,N_9178);
or U11033 (N_11033,N_6402,N_7012);
nand U11034 (N_11034,N_9923,N_5971);
and U11035 (N_11035,N_9926,N_9707);
and U11036 (N_11036,N_7304,N_8107);
nand U11037 (N_11037,N_8690,N_5201);
and U11038 (N_11038,N_5117,N_7198);
and U11039 (N_11039,N_5939,N_9262);
or U11040 (N_11040,N_7441,N_7673);
nand U11041 (N_11041,N_8349,N_6604);
or U11042 (N_11042,N_7051,N_5096);
nand U11043 (N_11043,N_6110,N_8625);
and U11044 (N_11044,N_9422,N_7552);
or U11045 (N_11045,N_8122,N_9397);
nor U11046 (N_11046,N_8227,N_8290);
nor U11047 (N_11047,N_9622,N_5879);
and U11048 (N_11048,N_7992,N_5722);
nor U11049 (N_11049,N_8889,N_5241);
or U11050 (N_11050,N_5347,N_8011);
nand U11051 (N_11051,N_5449,N_9565);
nand U11052 (N_11052,N_9579,N_9300);
nor U11053 (N_11053,N_5227,N_8260);
or U11054 (N_11054,N_5000,N_6980);
or U11055 (N_11055,N_9505,N_8263);
nor U11056 (N_11056,N_8076,N_5871);
and U11057 (N_11057,N_8357,N_8410);
or U11058 (N_11058,N_5493,N_7932);
nand U11059 (N_11059,N_5162,N_9333);
nor U11060 (N_11060,N_7259,N_8532);
and U11061 (N_11061,N_5739,N_8281);
or U11062 (N_11062,N_9727,N_5370);
nand U11063 (N_11063,N_7484,N_5514);
or U11064 (N_11064,N_7366,N_5970);
nand U11065 (N_11065,N_7056,N_7783);
and U11066 (N_11066,N_6358,N_9641);
nand U11067 (N_11067,N_5250,N_9111);
nand U11068 (N_11068,N_8699,N_6779);
nand U11069 (N_11069,N_9776,N_6577);
and U11070 (N_11070,N_5608,N_9931);
and U11071 (N_11071,N_8976,N_9832);
xor U11072 (N_11072,N_6876,N_8553);
nand U11073 (N_11073,N_7953,N_9512);
nand U11074 (N_11074,N_5174,N_5625);
nand U11075 (N_11075,N_9118,N_8204);
nand U11076 (N_11076,N_5673,N_6989);
and U11077 (N_11077,N_8856,N_8579);
and U11078 (N_11078,N_6842,N_5816);
nand U11079 (N_11079,N_9916,N_9860);
nand U11080 (N_11080,N_5501,N_6594);
nor U11081 (N_11081,N_7513,N_7926);
nor U11082 (N_11082,N_8748,N_8002);
and U11083 (N_11083,N_8074,N_9275);
or U11084 (N_11084,N_6078,N_7385);
nor U11085 (N_11085,N_7893,N_5011);
nand U11086 (N_11086,N_8643,N_5906);
or U11087 (N_11087,N_7448,N_9715);
nand U11088 (N_11088,N_8554,N_5652);
nor U11089 (N_11089,N_6924,N_9659);
nand U11090 (N_11090,N_7729,N_9445);
and U11091 (N_11091,N_6754,N_9709);
nor U11092 (N_11092,N_5489,N_9633);
and U11093 (N_11093,N_9625,N_7627);
and U11094 (N_11094,N_5128,N_6690);
nand U11095 (N_11095,N_9831,N_7658);
nor U11096 (N_11096,N_5025,N_6441);
or U11097 (N_11097,N_9793,N_7054);
or U11098 (N_11098,N_9248,N_7032);
and U11099 (N_11099,N_9125,N_7826);
nand U11100 (N_11100,N_5145,N_6878);
nor U11101 (N_11101,N_7747,N_7214);
nor U11102 (N_11102,N_5184,N_5825);
nor U11103 (N_11103,N_5401,N_9649);
or U11104 (N_11104,N_9753,N_9312);
nand U11105 (N_11105,N_6808,N_9190);
nand U11106 (N_11106,N_7688,N_5198);
nor U11107 (N_11107,N_6886,N_8308);
or U11108 (N_11108,N_7709,N_8658);
xnor U11109 (N_11109,N_8094,N_7454);
or U11110 (N_11110,N_5610,N_7319);
xor U11111 (N_11111,N_8530,N_7880);
nand U11112 (N_11112,N_8542,N_5176);
nand U11113 (N_11113,N_6244,N_6949);
and U11114 (N_11114,N_7675,N_7571);
or U11115 (N_11115,N_9458,N_5013);
xnor U11116 (N_11116,N_9219,N_7752);
nand U11117 (N_11117,N_6736,N_9808);
or U11118 (N_11118,N_6919,N_5297);
and U11119 (N_11119,N_6777,N_5779);
and U11120 (N_11120,N_5715,N_7561);
or U11121 (N_11121,N_6748,N_6018);
xnor U11122 (N_11122,N_7276,N_5057);
xor U11123 (N_11123,N_5012,N_7855);
xor U11124 (N_11124,N_7923,N_7800);
xor U11125 (N_11125,N_6226,N_7391);
or U11126 (N_11126,N_9359,N_8459);
nand U11127 (N_11127,N_7404,N_5838);
or U11128 (N_11128,N_9139,N_9438);
xnor U11129 (N_11129,N_9461,N_5146);
nand U11130 (N_11130,N_9269,N_6446);
xnor U11131 (N_11131,N_8657,N_8185);
or U11132 (N_11132,N_5158,N_5032);
nand U11133 (N_11133,N_8411,N_8865);
nor U11134 (N_11134,N_8819,N_5154);
nand U11135 (N_11135,N_6225,N_8879);
nor U11136 (N_11136,N_7741,N_8507);
or U11137 (N_11137,N_6091,N_7726);
nor U11138 (N_11138,N_7145,N_6660);
nand U11139 (N_11139,N_6360,N_9186);
or U11140 (N_11140,N_9150,N_5574);
and U11141 (N_11141,N_8903,N_8804);
nand U11142 (N_11142,N_7318,N_7335);
and U11143 (N_11143,N_6267,N_5671);
nand U11144 (N_11144,N_5434,N_5303);
or U11145 (N_11145,N_8466,N_9915);
or U11146 (N_11146,N_9977,N_5139);
and U11147 (N_11147,N_6222,N_7845);
or U11148 (N_11148,N_7710,N_7031);
nand U11149 (N_11149,N_9961,N_6390);
nand U11150 (N_11150,N_6429,N_8383);
nor U11151 (N_11151,N_7343,N_6896);
and U11152 (N_11152,N_7444,N_5766);
nor U11153 (N_11153,N_5130,N_8405);
nand U11154 (N_11154,N_5638,N_5555);
nand U11155 (N_11155,N_5978,N_7650);
nand U11156 (N_11156,N_5002,N_5400);
nor U11157 (N_11157,N_8822,N_5654);
and U11158 (N_11158,N_9881,N_9270);
nor U11159 (N_11159,N_7008,N_5084);
and U11160 (N_11160,N_5497,N_9773);
nor U11161 (N_11161,N_5050,N_7566);
nand U11162 (N_11162,N_7489,N_9999);
nor U11163 (N_11163,N_7808,N_7160);
nand U11164 (N_11164,N_9131,N_7030);
or U11165 (N_11165,N_6729,N_7652);
and U11166 (N_11166,N_6992,N_6329);
and U11167 (N_11167,N_7370,N_8727);
nand U11168 (N_11168,N_6805,N_6804);
nor U11169 (N_11169,N_9838,N_5942);
nand U11170 (N_11170,N_8468,N_5689);
or U11171 (N_11171,N_8169,N_5391);
xnor U11172 (N_11172,N_7666,N_6060);
and U11173 (N_11173,N_5617,N_9096);
or U11174 (N_11174,N_5386,N_7050);
and U11175 (N_11175,N_9129,N_9526);
nor U11176 (N_11176,N_5762,N_8637);
nor U11177 (N_11177,N_8668,N_7394);
or U11178 (N_11178,N_6679,N_5470);
and U11179 (N_11179,N_8946,N_9750);
xnor U11180 (N_11180,N_5415,N_8559);
xor U11181 (N_11181,N_8857,N_9280);
nor U11182 (N_11182,N_5648,N_7714);
or U11183 (N_11183,N_6007,N_8695);
nor U11184 (N_11184,N_7061,N_7701);
nand U11185 (N_11185,N_5406,N_7600);
or U11186 (N_11186,N_5160,N_5490);
xnor U11187 (N_11187,N_7059,N_6554);
nand U11188 (N_11188,N_5279,N_9271);
nor U11189 (N_11189,N_6862,N_7184);
nor U11190 (N_11190,N_8454,N_8835);
nor U11191 (N_11191,N_9104,N_7886);
nand U11192 (N_11192,N_5809,N_7194);
and U11193 (N_11193,N_7906,N_8775);
and U11194 (N_11194,N_9718,N_7980);
and U11195 (N_11195,N_6654,N_5344);
xor U11196 (N_11196,N_8234,N_9813);
nand U11197 (N_11197,N_7790,N_7756);
and U11198 (N_11198,N_6899,N_9588);
nor U11199 (N_11199,N_9955,N_7296);
or U11200 (N_11200,N_7698,N_8086);
and U11201 (N_11201,N_5101,N_7432);
and U11202 (N_11202,N_6772,N_7469);
and U11203 (N_11203,N_6774,N_9391);
and U11204 (N_11204,N_6603,N_7062);
nand U11205 (N_11205,N_8701,N_9204);
and U11206 (N_11206,N_8150,N_5238);
or U11207 (N_11207,N_8590,N_9743);
or U11208 (N_11208,N_7837,N_7306);
nor U11209 (N_11209,N_5759,N_6455);
nor U11210 (N_11210,N_6870,N_7442);
and U11211 (N_11211,N_9176,N_5064);
nor U11212 (N_11212,N_9225,N_9701);
or U11213 (N_11213,N_9873,N_7562);
nor U11214 (N_11214,N_8685,N_8158);
and U11215 (N_11215,N_9447,N_5151);
nand U11216 (N_11216,N_7947,N_8568);
and U11217 (N_11217,N_7312,N_7352);
nand U11218 (N_11218,N_6641,N_6296);
and U11219 (N_11219,N_6099,N_7423);
or U11220 (N_11220,N_5526,N_8851);
nand U11221 (N_11221,N_9876,N_9589);
nor U11222 (N_11222,N_7865,N_6614);
nand U11223 (N_11223,N_5549,N_6397);
or U11224 (N_11224,N_9959,N_5951);
or U11225 (N_11225,N_7195,N_8489);
nand U11226 (N_11226,N_9418,N_7605);
nor U11227 (N_11227,N_7332,N_6163);
nor U11228 (N_11228,N_6389,N_9318);
nand U11229 (N_11229,N_6629,N_6310);
or U11230 (N_11230,N_6181,N_6260);
and U11231 (N_11231,N_5601,N_8253);
nand U11232 (N_11232,N_7873,N_9895);
nor U11233 (N_11233,N_9091,N_7784);
and U11234 (N_11234,N_8640,N_5168);
nor U11235 (N_11235,N_6107,N_5750);
or U11236 (N_11236,N_6618,N_8220);
nor U11237 (N_11237,N_7078,N_9203);
nand U11238 (N_11238,N_8362,N_8836);
nor U11239 (N_11239,N_5353,N_6904);
nand U11240 (N_11240,N_6620,N_5442);
nand U11241 (N_11241,N_7156,N_5429);
nor U11242 (N_11242,N_8218,N_6045);
or U11243 (N_11243,N_5404,N_7181);
and U11244 (N_11244,N_8477,N_9782);
nor U11245 (N_11245,N_9720,N_8151);
nand U11246 (N_11246,N_7358,N_7485);
or U11247 (N_11247,N_5694,N_7393);
xnor U11248 (N_11248,N_8623,N_5454);
and U11249 (N_11249,N_9062,N_6055);
or U11250 (N_11250,N_6986,N_9812);
or U11251 (N_11251,N_5215,N_8339);
nand U11252 (N_11252,N_6778,N_9222);
xor U11253 (N_11253,N_8562,N_7692);
nand U11254 (N_11254,N_9665,N_7188);
nor U11255 (N_11255,N_7086,N_9848);
nand U11256 (N_11256,N_5643,N_6272);
xnor U11257 (N_11257,N_6814,N_6815);
or U11258 (N_11258,N_5983,N_5891);
xnor U11259 (N_11259,N_5559,N_6175);
or U11260 (N_11260,N_5226,N_5285);
nor U11261 (N_11261,N_6334,N_9443);
nor U11262 (N_11262,N_7921,N_6065);
nor U11263 (N_11263,N_5651,N_9444);
and U11264 (N_11264,N_6585,N_5166);
or U11265 (N_11265,N_8153,N_8992);
nand U11266 (N_11266,N_8449,N_9971);
and U11267 (N_11267,N_8172,N_9556);
or U11268 (N_11268,N_6394,N_6541);
nor U11269 (N_11269,N_5278,N_9956);
or U11270 (N_11270,N_8244,N_9439);
and U11271 (N_11271,N_5646,N_5440);
nor U11272 (N_11272,N_6561,N_6781);
and U11273 (N_11273,N_8766,N_9468);
xnor U11274 (N_11274,N_5613,N_8066);
nand U11275 (N_11275,N_5873,N_9398);
nand U11276 (N_11276,N_5653,N_5692);
and U11277 (N_11277,N_8230,N_5296);
nand U11278 (N_11278,N_9760,N_7870);
or U11279 (N_11279,N_8761,N_8673);
xor U11280 (N_11280,N_8758,N_6910);
or U11281 (N_11281,N_5088,N_7497);
nor U11282 (N_11282,N_8332,N_8485);
and U11283 (N_11283,N_5882,N_5077);
xor U11284 (N_11284,N_6405,N_6034);
and U11285 (N_11285,N_5459,N_9747);
nor U11286 (N_11286,N_8323,N_9317);
nor U11287 (N_11287,N_5135,N_7594);
or U11288 (N_11288,N_6514,N_8111);
or U11289 (N_11289,N_7382,N_5621);
or U11290 (N_11290,N_5630,N_6670);
nor U11291 (N_11291,N_7883,N_8277);
nor U11292 (N_11292,N_5974,N_7831);
and U11293 (N_11293,N_6218,N_6258);
and U11294 (N_11294,N_8861,N_5909);
and U11295 (N_11295,N_8982,N_5875);
nand U11296 (N_11296,N_6940,N_7629);
and U11297 (N_11297,N_6838,N_5389);
nand U11298 (N_11298,N_6983,N_8920);
nand U11299 (N_11299,N_5738,N_9115);
or U11300 (N_11300,N_7235,N_9657);
nand U11301 (N_11301,N_6412,N_5112);
nand U11302 (N_11302,N_7093,N_5222);
and U11303 (N_11303,N_5211,N_5163);
nor U11304 (N_11304,N_9322,N_5872);
and U11305 (N_11305,N_9044,N_5849);
nand U11306 (N_11306,N_9221,N_5963);
nor U11307 (N_11307,N_6798,N_6318);
nand U11308 (N_11308,N_7716,N_7456);
nand U11309 (N_11309,N_8708,N_6168);
and U11310 (N_11310,N_5295,N_5426);
nand U11311 (N_11311,N_7840,N_7019);
xnor U11312 (N_11312,N_5614,N_5862);
nand U11313 (N_11313,N_7212,N_8988);
xor U11314 (N_11314,N_6126,N_9943);
xnor U11315 (N_11315,N_9613,N_9559);
xor U11316 (N_11316,N_8918,N_6521);
nand U11317 (N_11317,N_5543,N_7759);
nor U11318 (N_11318,N_9277,N_8510);
and U11319 (N_11319,N_8285,N_9228);
or U11320 (N_11320,N_9417,N_8904);
xor U11321 (N_11321,N_8984,N_8235);
nand U11322 (N_11322,N_8279,N_8943);
nand U11323 (N_11323,N_5907,N_7994);
or U11324 (N_11324,N_7610,N_6990);
nand U11325 (N_11325,N_6476,N_7621);
or U11326 (N_11326,N_5676,N_5109);
nand U11327 (N_11327,N_7487,N_6765);
and U11328 (N_11328,N_7117,N_7524);
nand U11329 (N_11329,N_6553,N_5451);
or U11330 (N_11330,N_7314,N_6649);
nor U11331 (N_11331,N_6313,N_6369);
or U11332 (N_11332,N_9540,N_6233);
and U11333 (N_11333,N_8749,N_7915);
nand U11334 (N_11334,N_6264,N_9366);
and U11335 (N_11335,N_7321,N_9284);
xor U11336 (N_11336,N_5195,N_8556);
nor U11337 (N_11337,N_8488,N_9680);
or U11338 (N_11338,N_9500,N_9525);
or U11339 (N_11339,N_6488,N_9393);
or U11340 (N_11340,N_8972,N_8013);
or U11341 (N_11341,N_5602,N_8108);
xor U11342 (N_11342,N_7191,N_7711);
xnor U11343 (N_11343,N_8261,N_5421);
or U11344 (N_11344,N_9171,N_9847);
nor U11345 (N_11345,N_8149,N_5171);
xnor U11346 (N_11346,N_5364,N_6925);
and U11347 (N_11347,N_5936,N_8979);
and U11348 (N_11348,N_8202,N_5554);
or U11349 (N_11349,N_8326,N_9875);
nand U11350 (N_11350,N_7118,N_9029);
or U11351 (N_11351,N_7589,N_5106);
nand U11352 (N_11352,N_5220,N_8046);
or U11353 (N_11353,N_6342,N_8656);
and U11354 (N_11354,N_8674,N_8855);
nor U11355 (N_11355,N_6201,N_5916);
nor U11356 (N_11356,N_8128,N_5538);
or U11357 (N_11357,N_6187,N_5286);
nor U11358 (N_11358,N_9722,N_5233);
and U11359 (N_11359,N_9874,N_5958);
or U11360 (N_11360,N_7904,N_9636);
or U11361 (N_11361,N_5127,N_9056);
nor U11362 (N_11362,N_9630,N_6852);
nor U11363 (N_11363,N_9674,N_8713);
nor U11364 (N_11364,N_8415,N_5683);
nand U11365 (N_11365,N_9601,N_6235);
nand U11366 (N_11366,N_9361,N_9538);
nor U11367 (N_11367,N_5167,N_7703);
xor U11368 (N_11368,N_5540,N_5735);
and U11369 (N_11369,N_6191,N_8846);
or U11370 (N_11370,N_6416,N_6189);
xnor U11371 (N_11371,N_6373,N_5582);
nand U11372 (N_11372,N_5092,N_9205);
xnor U11373 (N_11373,N_8564,N_5605);
nor U11374 (N_11374,N_7103,N_9193);
nand U11375 (N_11375,N_6662,N_5342);
nand U11376 (N_11376,N_7168,N_6180);
nor U11377 (N_11377,N_9695,N_6936);
nand U11378 (N_11378,N_5393,N_6146);
nor U11379 (N_11379,N_5955,N_6014);
or U11380 (N_11380,N_9844,N_5456);
nor U11381 (N_11381,N_5273,N_8291);
nand U11382 (N_11382,N_7821,N_7015);
or U11383 (N_11383,N_6083,N_5597);
nand U11384 (N_11384,N_9218,N_6388);
nand U11385 (N_11385,N_8315,N_7665);
and U11386 (N_11386,N_7148,N_5014);
nor U11387 (N_11387,N_6548,N_8239);
nor U11388 (N_11388,N_6144,N_7787);
and U11389 (N_11389,N_9824,N_6375);
nand U11390 (N_11390,N_8120,N_6124);
nand U11391 (N_11391,N_7287,N_9910);
and U11392 (N_11392,N_8947,N_7070);
xor U11393 (N_11393,N_6999,N_8070);
and U11394 (N_11394,N_9346,N_7690);
or U11395 (N_11395,N_7189,N_5817);
and U11396 (N_11396,N_5495,N_5294);
nor U11397 (N_11397,N_5450,N_8247);
or U11398 (N_11398,N_7374,N_8692);
nand U11399 (N_11399,N_9294,N_5363);
nor U11400 (N_11400,N_5961,N_9310);
and U11401 (N_11401,N_5758,N_8655);
and U11402 (N_11402,N_7460,N_8001);
nand U11403 (N_11403,N_6543,N_8106);
xnor U11404 (N_11404,N_8589,N_9841);
xor U11405 (N_11405,N_6834,N_5475);
nand U11406 (N_11406,N_5655,N_6847);
and U11407 (N_11407,N_7250,N_6012);
or U11408 (N_11408,N_5333,N_6567);
nand U11409 (N_11409,N_5125,N_6695);
nand U11410 (N_11410,N_5365,N_8809);
or U11411 (N_11411,N_5707,N_8304);
and U11412 (N_11412,N_9123,N_7427);
or U11413 (N_11413,N_8404,N_8922);
nor U11414 (N_11414,N_7707,N_7901);
nand U11415 (N_11415,N_5748,N_9344);
or U11416 (N_11416,N_8537,N_7581);
nand U11417 (N_11417,N_7283,N_5147);
xnor U11418 (N_11418,N_7898,N_8936);
nand U11419 (N_11419,N_8540,N_8950);
nand U11420 (N_11420,N_6791,N_7875);
and U11421 (N_11421,N_5476,N_7088);
nor U11422 (N_11422,N_5315,N_6903);
and U11423 (N_11423,N_9867,N_7647);
and U11424 (N_11424,N_6647,N_9106);
and U11425 (N_11425,N_9015,N_6820);
or U11426 (N_11426,N_6114,N_9448);
nor U11427 (N_11427,N_7587,N_7683);
or U11428 (N_11428,N_7400,N_7273);
nand U11429 (N_11429,N_6897,N_5200);
and U11430 (N_11430,N_5187,N_6727);
or U11431 (N_11431,N_9180,N_5380);
xnor U11432 (N_11432,N_5544,N_9223);
or U11433 (N_11433,N_8526,N_9741);
and U11434 (N_11434,N_6330,N_5317);
or U11435 (N_11435,N_6234,N_8593);
or U11436 (N_11436,N_7517,N_5413);
nand U11437 (N_11437,N_8604,N_5086);
nand U11438 (N_11438,N_6367,N_8250);
and U11439 (N_11439,N_5103,N_7933);
or U11440 (N_11440,N_5115,N_9230);
nor U11441 (N_11441,N_9751,N_5196);
and U11442 (N_11442,N_8609,N_7359);
nand U11443 (N_11443,N_8240,N_6711);
nor U11444 (N_11444,N_7508,N_5967);
and U11445 (N_11445,N_6173,N_5305);
and U11446 (N_11446,N_6086,N_6335);
or U11447 (N_11447,N_6555,N_5098);
nor U11448 (N_11448,N_6957,N_7029);
or U11449 (N_11449,N_7988,N_8914);
nor U11450 (N_11450,N_5169,N_6082);
nand U11451 (N_11451,N_7918,N_8473);
xor U11452 (N_11452,N_5432,N_5975);
and U11453 (N_11453,N_5772,N_5256);
and U11454 (N_11454,N_8520,N_6290);
nand U11455 (N_11455,N_9616,N_7301);
nand U11456 (N_11456,N_8689,N_7337);
nand U11457 (N_11457,N_9466,N_8767);
or U11458 (N_11458,N_8960,N_8783);
and U11459 (N_11459,N_5888,N_9996);
nor U11460 (N_11460,N_9547,N_6783);
nor U11461 (N_11461,N_6382,N_5395);
nand U11462 (N_11462,N_7183,N_9092);
nor U11463 (N_11463,N_9128,N_7739);
xor U11464 (N_11464,N_8567,N_8683);
nor U11465 (N_11465,N_5886,N_8548);
and U11466 (N_11466,N_7220,N_9973);
xor U11467 (N_11467,N_8115,N_5757);
and U11468 (N_11468,N_8375,N_7563);
nor U11469 (N_11469,N_7437,N_9699);
and U11470 (N_11470,N_6288,N_6821);
and U11471 (N_11471,N_8040,N_5102);
nand U11472 (N_11472,N_6818,N_7549);
nand U11473 (N_11473,N_8043,N_8866);
nand U11474 (N_11474,N_5186,N_5532);
or U11475 (N_11475,N_6026,N_8320);
and U11476 (N_11476,N_7708,N_7341);
nand U11477 (N_11477,N_8653,N_8181);
and U11478 (N_11478,N_5571,N_5122);
and U11479 (N_11479,N_7995,N_9974);
nor U11480 (N_11480,N_7822,N_5510);
or U11481 (N_11481,N_8214,N_5005);
nor U11482 (N_11482,N_8508,N_5575);
xor U11483 (N_11483,N_5496,N_7612);
or U11484 (N_11484,N_7323,N_8483);
nor U11485 (N_11485,N_7555,N_9484);
or U11486 (N_11486,N_9637,N_6627);
or U11487 (N_11487,N_6709,N_5519);
nand U11488 (N_11488,N_6866,N_9551);
nand U11489 (N_11489,N_6557,N_7228);
xnor U11490 (N_11490,N_9229,N_5685);
and U11491 (N_11491,N_6872,N_9804);
nor U11492 (N_11492,N_6319,N_6268);
nand U11493 (N_11493,N_9172,N_5568);
nand U11494 (N_11494,N_5856,N_8684);
nor U11495 (N_11495,N_8471,N_6574);
and U11496 (N_11496,N_7246,N_8231);
and U11497 (N_11497,N_5843,N_9518);
nor U11498 (N_11498,N_8990,N_9059);
nor U11499 (N_11499,N_6869,N_8849);
nand U11500 (N_11500,N_6762,N_6491);
or U11501 (N_11501,N_5231,N_6845);
or U11502 (N_11502,N_8015,N_7818);
or U11503 (N_11503,N_7159,N_6166);
nor U11504 (N_11504,N_9865,N_8419);
nor U11505 (N_11505,N_6058,N_6271);
nor U11506 (N_11506,N_8999,N_5725);
nand U11507 (N_11507,N_5394,N_9089);
or U11508 (N_11508,N_8254,N_6344);
and U11509 (N_11509,N_6840,N_8045);
nand U11510 (N_11510,N_6105,N_8521);
nand U11511 (N_11511,N_6434,N_5599);
nand U11512 (N_11512,N_8380,N_5990);
nand U11513 (N_11513,N_6152,N_8575);
nor U11514 (N_11514,N_6787,N_5991);
nand U11515 (N_11515,N_6044,N_5901);
or U11516 (N_11516,N_7642,N_6381);
or U11517 (N_11517,N_8060,N_7857);
nor U11518 (N_11518,N_9053,N_9016);
nand U11519 (N_11519,N_8423,N_6042);
nand U11520 (N_11520,N_9127,N_7799);
xor U11521 (N_11521,N_5356,N_5039);
and U11522 (N_11522,N_7588,N_9200);
and U11523 (N_11523,N_9902,N_8831);
nand U11524 (N_11524,N_5777,N_8957);
nor U11525 (N_11525,N_7491,N_9759);
and U11526 (N_11526,N_6261,N_8759);
and U11527 (N_11527,N_7413,N_5656);
or U11528 (N_11528,N_6081,N_9827);
nor U11529 (N_11529,N_6072,N_8812);
or U11530 (N_11530,N_9380,N_7345);
nand U11531 (N_11531,N_7260,N_8088);
nor U11532 (N_11532,N_5944,N_5345);
or U11533 (N_11533,N_9890,N_6578);
nand U11534 (N_11534,N_6917,N_9612);
nor U11535 (N_11535,N_7186,N_5989);
and U11536 (N_11536,N_8907,N_8431);
nand U11537 (N_11537,N_6227,N_9819);
nor U11538 (N_11538,N_8268,N_8686);
or U11539 (N_11539,N_6860,N_6064);
nand U11540 (N_11540,N_8402,N_6623);
nand U11541 (N_11541,N_6362,N_8543);
nand U11542 (N_11542,N_5149,N_8131);
nand U11543 (N_11543,N_5322,N_8199);
or U11544 (N_11544,N_8888,N_9141);
nor U11545 (N_11545,N_8222,N_8852);
nor U11546 (N_11546,N_8693,N_9164);
nor U11547 (N_11547,N_5133,N_9784);
xnor U11548 (N_11548,N_9126,N_7269);
or U11549 (N_11549,N_7999,N_9591);
nor U11550 (N_11550,N_9705,N_5806);
nand U11551 (N_11551,N_8790,N_6927);
nand U11552 (N_11552,N_8799,N_5878);
or U11553 (N_11553,N_6492,N_6469);
and U11554 (N_11554,N_6706,N_7720);
and U11555 (N_11555,N_5134,N_8329);
nor U11556 (N_11556,N_9918,N_7851);
nand U11557 (N_11557,N_6029,N_5634);
xor U11558 (N_11558,N_8694,N_5314);
and U11559 (N_11559,N_6472,N_6519);
and U11560 (N_11560,N_9474,N_6663);
or U11561 (N_11561,N_5031,N_8779);
or U11562 (N_11562,N_6463,N_9301);
and U11563 (N_11563,N_7705,N_8971);
nor U11564 (N_11564,N_7987,N_7027);
and U11565 (N_11565,N_5828,N_7351);
and U11566 (N_11566,N_5329,N_6704);
nand U11567 (N_11567,N_7071,N_6682);
and U11568 (N_11568,N_6640,N_5326);
or U11569 (N_11569,N_5008,N_8347);
nor U11570 (N_11570,N_7686,N_6003);
nor U11571 (N_11571,N_7483,N_6658);
or U11572 (N_11572,N_6775,N_9672);
nor U11573 (N_11573,N_6025,N_9914);
nand U11574 (N_11574,N_5709,N_9676);
or U11575 (N_11575,N_5242,N_6735);
or U11576 (N_11576,N_8596,N_7311);
xnor U11577 (N_11577,N_7190,N_6773);
nor U11578 (N_11578,N_6084,N_6943);
and U11579 (N_11579,N_9531,N_5214);
nor U11580 (N_11580,N_5313,N_6854);
nand U11581 (N_11581,N_7046,N_9754);
nor U11582 (N_11582,N_6197,N_9426);
nand U11583 (N_11583,N_8427,N_9502);
or U11584 (N_11584,N_6672,N_9645);
xor U11585 (N_11585,N_9093,N_8118);
nand U11586 (N_11586,N_9303,N_6184);
nand U11587 (N_11587,N_8595,N_9821);
nand U11588 (N_11588,N_8881,N_6154);
nand U11589 (N_11589,N_7879,N_8796);
and U11590 (N_11590,N_9887,N_6850);
nand U11591 (N_11591,N_8891,N_7830);
nand U11592 (N_11592,N_7387,N_9036);
nor U11593 (N_11593,N_6414,N_5976);
or U11594 (N_11594,N_7278,N_8916);
nor U11595 (N_11595,N_5714,N_6807);
nor U11596 (N_11596,N_5185,N_8545);
and U11597 (N_11597,N_6513,N_9292);
nor U11598 (N_11598,N_9560,N_6995);
nor U11599 (N_11599,N_6024,N_9590);
and U11600 (N_11600,N_8125,N_5418);
nand U11601 (N_11601,N_9290,N_5691);
or U11602 (N_11602,N_7803,N_6022);
nand U11603 (N_11603,N_8421,N_6138);
nor U11604 (N_11604,N_9285,N_9958);
or U11605 (N_11605,N_8915,N_6502);
or U11606 (N_11606,N_6895,N_6481);
nand U11607 (N_11607,N_9716,N_7511);
and U11608 (N_11608,N_8504,N_9233);
or U11609 (N_11609,N_7938,N_6733);
or U11610 (N_11610,N_5040,N_5061);
or U11611 (N_11611,N_8989,N_6051);
or U11612 (N_11612,N_5782,N_5504);
nor U11613 (N_11613,N_7153,N_9605);
and U11614 (N_11614,N_5746,N_5428);
or U11615 (N_11615,N_6299,N_5205);
nand U11616 (N_11616,N_8647,N_9800);
or U11617 (N_11617,N_7026,N_6937);
nand U11618 (N_11618,N_7123,N_9609);
nor U11619 (N_11619,N_9108,N_5933);
or U11620 (N_11620,N_5381,N_9368);
nand U11621 (N_11621,N_5681,N_5687);
and U11622 (N_11622,N_8370,N_9787);
nor U11623 (N_11623,N_5966,N_5826);
and U11624 (N_11624,N_6046,N_6655);
nand U11625 (N_11625,N_7651,N_8919);
nor U11626 (N_11626,N_6552,N_9238);
or U11627 (N_11627,N_6551,N_6400);
or U11628 (N_11628,N_7573,N_8020);
or U11629 (N_11629,N_5598,N_9794);
and U11630 (N_11630,N_7696,N_6643);
or U11631 (N_11631,N_6135,N_8387);
xor U11632 (N_11632,N_5023,N_7303);
nand U11633 (N_11633,N_7792,N_5677);
or U11634 (N_11634,N_6761,N_9504);
nand U11635 (N_11635,N_9697,N_6619);
nor U11636 (N_11636,N_8788,N_7025);
nand U11637 (N_11637,N_8997,N_9298);
nand U11638 (N_11638,N_8697,N_8374);
nand U11639 (N_11639,N_6705,N_6507);
and U11640 (N_11640,N_5461,N_6328);
xor U11641 (N_11641,N_9324,N_8853);
nand U11642 (N_11642,N_6297,N_8867);
and U11643 (N_11643,N_8065,N_9007);
and U11644 (N_11644,N_9501,N_8765);
nor U11645 (N_11645,N_6831,N_6853);
nor U11646 (N_11646,N_7841,N_9068);
and U11647 (N_11647,N_6797,N_6131);
nand U11648 (N_11648,N_6363,N_6423);
or U11649 (N_11649,N_5769,N_6207);
nor U11650 (N_11650,N_6103,N_9169);
and U11651 (N_11651,N_5547,N_8830);
nor U11652 (N_11652,N_9792,N_8055);
nor U11653 (N_11653,N_9877,N_7543);
nand U11654 (N_11654,N_6988,N_6549);
or U11655 (N_11655,N_9201,N_7290);
nor U11656 (N_11656,N_8366,N_7225);
nor U11657 (N_11657,N_7694,N_6580);
nor U11658 (N_11658,N_6130,N_6944);
nor U11659 (N_11659,N_5956,N_7569);
nor U11660 (N_11660,N_7531,N_8725);
nand U11661 (N_11661,N_6354,N_8905);
nor U11662 (N_11662,N_6395,N_8718);
nand U11663 (N_11663,N_8189,N_6503);
nor U11664 (N_11664,N_7068,N_5439);
or U11665 (N_11665,N_8148,N_6386);
nand U11666 (N_11666,N_8952,N_6243);
or U11667 (N_11667,N_5136,N_6440);
or U11668 (N_11668,N_5596,N_6638);
and U11669 (N_11669,N_8413,N_5521);
nand U11670 (N_11670,N_8390,N_7121);
nor U11671 (N_11671,N_6953,N_9849);
xnor U11672 (N_11672,N_7209,N_6525);
nand U11673 (N_11673,N_5108,N_7611);
and U11674 (N_11674,N_5488,N_7671);
and U11675 (N_11675,N_7648,N_5850);
nor U11676 (N_11676,N_9663,N_5143);
nand U11677 (N_11677,N_8179,N_5183);
or U11678 (N_11678,N_7077,N_5020);
and U11679 (N_11679,N_5841,N_7052);
nor U11680 (N_11680,N_9414,N_8414);
nor U11681 (N_11681,N_6536,N_9567);
and U11682 (N_11682,N_9058,N_8546);
nand U11683 (N_11683,N_8436,N_5419);
and U11684 (N_11684,N_9194,N_9764);
nor U11685 (N_11685,N_7244,N_5731);
nor U11686 (N_11686,N_8825,N_9078);
xor U11687 (N_11687,N_6539,N_6877);
xor U11688 (N_11688,N_8101,N_9071);
xor U11689 (N_11689,N_5282,N_7866);
or U11690 (N_11690,N_7958,N_9634);
and U11691 (N_11691,N_8191,N_8710);
or U11692 (N_11692,N_8722,N_5111);
nor U11693 (N_11693,N_8135,N_8501);
nand U11694 (N_11694,N_6913,N_7649);
nand U11695 (N_11695,N_7120,N_6224);
nand U11696 (N_11696,N_8229,N_9140);
nor U11697 (N_11697,N_8762,N_6891);
nand U11698 (N_11698,N_5309,N_8317);
xnor U11699 (N_11699,N_6766,N_5793);
nand U11700 (N_11700,N_5846,N_9815);
nor U11701 (N_11701,N_5865,N_8408);
and U11702 (N_11702,N_8667,N_5384);
and U11703 (N_11703,N_8371,N_5932);
or U11704 (N_11704,N_8654,N_5009);
xor U11705 (N_11705,N_9052,N_5609);
and U11706 (N_11706,N_7435,N_6881);
or U11707 (N_11707,N_8095,N_5235);
nor U11708 (N_11708,N_7518,N_6005);
nor U11709 (N_11709,N_9509,N_8217);
nand U11710 (N_11710,N_8245,N_5377);
and U11711 (N_11711,N_5069,N_9675);
nor U11712 (N_11712,N_8882,N_9944);
nor U11713 (N_11713,N_9135,N_8133);
nor U11714 (N_11714,N_5965,N_8073);
nand U11715 (N_11715,N_6333,N_8863);
nor U11716 (N_11716,N_9388,N_7365);
nand U11717 (N_11717,N_7789,N_8295);
xnor U11718 (N_11718,N_9734,N_9327);
and U11719 (N_11719,N_7210,N_6134);
xor U11720 (N_11720,N_9026,N_5744);
or U11721 (N_11721,N_9814,N_7682);
nor U11722 (N_11722,N_9065,N_9740);
nor U11723 (N_11723,N_8912,N_9266);
and U11724 (N_11724,N_6966,N_9651);
or U11725 (N_11725,N_9569,N_7544);
nor U11726 (N_11726,N_6734,N_6303);
or U11727 (N_11727,N_6597,N_8583);
or U11728 (N_11728,N_5919,N_9941);
xnor U11729 (N_11729,N_5350,N_9639);
nor U11730 (N_11730,N_8676,N_9805);
and U11731 (N_11731,N_7433,N_9339);
and U11732 (N_11732,N_5584,N_5173);
or U11733 (N_11733,N_6047,N_5984);
and U11734 (N_11734,N_5588,N_9045);
or U11735 (N_11735,N_7482,N_5212);
nand U11736 (N_11736,N_5026,N_9241);
nor U11737 (N_11737,N_6712,N_5623);
and U11738 (N_11738,N_5764,N_7065);
and U11739 (N_11739,N_7105,N_9090);
and U11740 (N_11740,N_6223,N_8967);
nor U11741 (N_11741,N_5960,N_7717);
nor U11742 (N_11742,N_8465,N_8307);
and U11743 (N_11743,N_9954,N_8246);
nand U11744 (N_11744,N_7353,N_8597);
or U11745 (N_11745,N_8605,N_9939);
nand U11746 (N_11746,N_8330,N_7949);
nor U11747 (N_11747,N_5457,N_9184);
or U11748 (N_11748,N_9410,N_9828);
nand U11749 (N_11749,N_6645,N_8977);
or U11750 (N_11750,N_8003,N_9449);
nor U11751 (N_11751,N_8745,N_6931);
xor U11752 (N_11752,N_7622,N_7368);
nand U11753 (N_11753,N_7494,N_6443);
nor U11754 (N_11754,N_6062,N_6743);
or U11755 (N_11755,N_6245,N_6691);
and U11756 (N_11756,N_8175,N_9900);
or U11757 (N_11757,N_8302,N_5664);
or U11758 (N_11758,N_8644,N_7939);
or U11759 (N_11759,N_8816,N_8025);
and U11760 (N_11760,N_8635,N_9879);
nor U11761 (N_11761,N_7538,N_9544);
nor U11762 (N_11762,N_9107,N_5204);
nand U11763 (N_11763,N_7124,N_6102);
or U11764 (N_11764,N_9896,N_7285);
xnor U11765 (N_11765,N_5905,N_6020);
and U11766 (N_11766,N_8276,N_5068);
nand U11767 (N_11767,N_5908,N_5788);
or U11768 (N_11768,N_5539,N_9188);
or U11769 (N_11769,N_8618,N_6835);
and U11770 (N_11770,N_7275,N_5367);
nand U11771 (N_11771,N_8047,N_9496);
nand U11772 (N_11772,N_9763,N_5868);
nand U11773 (N_11773,N_8344,N_7229);
nor U11774 (N_11774,N_6309,N_8941);
nand U11775 (N_11775,N_8662,N_6109);
or U11776 (N_11776,N_6509,N_7676);
or U11777 (N_11777,N_9767,N_8008);
and U11778 (N_11778,N_9235,N_5072);
and U11779 (N_11779,N_5925,N_9033);
nand U11780 (N_11780,N_8791,N_9724);
and U11781 (N_11781,N_5208,N_8509);
nand U11782 (N_11782,N_9781,N_8581);
nor U11783 (N_11783,N_8412,N_7596);
nand U11784 (N_11784,N_5669,N_7791);
nand U11785 (N_11785,N_9423,N_7098);
nand U11786 (N_11786,N_5232,N_6118);
nor U11787 (N_11787,N_9060,N_7200);
nand U11788 (N_11788,N_8996,N_6530);
and U11789 (N_11789,N_8478,N_7011);
or U11790 (N_11790,N_8707,N_6349);
and U11791 (N_11791,N_6532,N_9566);
nand U11792 (N_11792,N_7466,N_8053);
and U11793 (N_11793,N_6665,N_9401);
and U11794 (N_11794,N_6147,N_5775);
or U11795 (N_11795,N_5361,N_9830);
nand U11796 (N_11796,N_6471,N_6343);
nand U11797 (N_11797,N_7618,N_8286);
and U11798 (N_11798,N_8042,N_8777);
or U11799 (N_11799,N_9861,N_9117);
and U11800 (N_11800,N_8188,N_7950);
and U11801 (N_11801,N_7173,N_6612);
nand U11802 (N_11802,N_5352,N_5743);
nand U11803 (N_11803,N_7208,N_8763);
nand U11804 (N_11804,N_8665,N_6348);
and U11805 (N_11805,N_5973,N_7961);
nand U11806 (N_11806,N_6837,N_9165);
and U11807 (N_11807,N_8688,N_8027);
and U11808 (N_11808,N_5604,N_6143);
nor U11809 (N_11809,N_6486,N_5035);
nand U11810 (N_11810,N_8737,N_8552);
or U11811 (N_11811,N_8272,N_8742);
nand U11812 (N_11812,N_5705,N_5896);
nor U11813 (N_11813,N_9655,N_6874);
nand U11814 (N_11814,N_7256,N_9568);
and U11815 (N_11815,N_9658,N_5774);
nor U11816 (N_11816,N_8394,N_5941);
and U11817 (N_11817,N_7347,N_6067);
and U11818 (N_11818,N_7333,N_5330);
nor U11819 (N_11819,N_6547,N_6789);
nand U11820 (N_11820,N_9227,N_6710);
nor U11821 (N_11821,N_7219,N_9144);
nor U11822 (N_11822,N_6898,N_5576);
nor U11823 (N_11823,N_5611,N_8327);
nor U11824 (N_11824,N_7308,N_6470);
nor U11825 (N_11825,N_8626,N_5864);
nand U11826 (N_11826,N_9211,N_9652);
and U11827 (N_11827,N_6112,N_7028);
and U11828 (N_11828,N_6475,N_5663);
and U11829 (N_11829,N_9113,N_5801);
nand U11830 (N_11830,N_8207,N_7829);
nor U11831 (N_11831,N_6316,N_7801);
nor U11832 (N_11832,N_8012,N_6581);
nor U11833 (N_11833,N_9628,N_6563);
nor U11834 (N_11834,N_5926,N_5796);
and U11835 (N_11835,N_6150,N_9723);
nand U11836 (N_11836,N_7218,N_8447);
nor U11837 (N_11837,N_6680,N_7564);
nor U11838 (N_11838,N_8885,N_7281);
nor U11839 (N_11839,N_5397,N_8403);
or U11840 (N_11840,N_8353,N_9099);
xnor U11841 (N_11841,N_7136,N_8030);
nor U11842 (N_11842,N_7583,N_8050);
nand U11843 (N_11843,N_8084,N_8991);
nand U11844 (N_11844,N_7167,N_6544);
and U11845 (N_11845,N_7390,N_8105);
or U11846 (N_11846,N_9878,N_9785);
or U11847 (N_11847,N_7638,N_6119);
and U11848 (N_11848,N_8934,N_5913);
xor U11849 (N_11849,N_9464,N_8031);
nand U11850 (N_11850,N_7725,N_7418);
and U11851 (N_11851,N_6600,N_8491);
and U11852 (N_11852,N_9646,N_8516);
nand U11853 (N_11853,N_9855,N_6393);
nor U11854 (N_11854,N_8318,N_8549);
nand U11855 (N_11855,N_8033,N_8434);
or U11856 (N_11856,N_9988,N_8152);
or U11857 (N_11857,N_7073,N_7036);
and U11858 (N_11858,N_5408,N_5999);
nand U11859 (N_11859,N_7850,N_9341);
xnor U11860 (N_11860,N_9913,N_8829);
nor U11861 (N_11861,N_9493,N_8416);
xor U11862 (N_11862,N_9762,N_9069);
or U11863 (N_11863,N_9580,N_7431);
nand U11864 (N_11864,N_6760,N_6564);
nor U11865 (N_11865,N_8890,N_6153);
or U11866 (N_11866,N_5253,N_6646);
nand U11867 (N_11867,N_8303,N_9592);
nand U11868 (N_11868,N_7614,N_5259);
nor U11869 (N_11869,N_5508,N_6909);
nor U11870 (N_11870,N_7668,N_5049);
and U11871 (N_11871,N_5047,N_7224);
nand U11872 (N_11872,N_8209,N_7728);
nor U11873 (N_11873,N_7819,N_7945);
nand U11874 (N_11874,N_7633,N_8017);
xor U11875 (N_11875,N_9452,N_9626);
or U11876 (N_11876,N_9296,N_5355);
and U11877 (N_11877,N_9728,N_5583);
nor U11878 (N_11878,N_8146,N_6346);
nand U11879 (N_11879,N_5674,N_9386);
nand U11880 (N_11880,N_8407,N_9347);
and U11881 (N_11881,N_8963,N_9321);
and U11882 (N_11882,N_9991,N_7110);
nor U11883 (N_11883,N_9067,N_6345);
nor U11884 (N_11884,N_7227,N_5922);
xor U11885 (N_11885,N_8801,N_7634);
or U11886 (N_11886,N_6000,N_5409);
or U11887 (N_11887,N_5224,N_8114);
and U11888 (N_11888,N_8439,N_6039);
and U11889 (N_11889,N_7503,N_8474);
and U11890 (N_11890,N_6238,N_8800);
nor U11891 (N_11891,N_5950,N_9094);
nor U11892 (N_11892,N_7488,N_8155);
nand U11893 (N_11893,N_9240,N_9992);
nor U11894 (N_11894,N_9465,N_5727);
and U11895 (N_11895,N_6028,N_5001);
nor U11896 (N_11896,N_6958,N_6833);
or U11897 (N_11897,N_6230,N_7292);
or U11898 (N_11898,N_6454,N_6459);
xor U11899 (N_11899,N_5114,N_7119);
nand U11900 (N_11900,N_9047,N_6749);
or U11901 (N_11901,N_6371,N_7211);
and U11902 (N_11902,N_7529,N_8314);
and U11903 (N_11903,N_5616,N_6880);
and U11904 (N_11904,N_5354,N_8007);
and U11905 (N_11905,N_9035,N_8529);
and U11906 (N_11906,N_8660,N_5647);
or U11907 (N_11907,N_8630,N_5464);
and U11908 (N_11908,N_7905,N_5481);
and U11909 (N_11909,N_7000,N_9690);
and U11910 (N_11910,N_8190,N_9738);
nor U11911 (N_11911,N_7751,N_5794);
nand U11912 (N_11912,N_5923,N_6031);
or U11913 (N_11913,N_6116,N_8569);
nand U11914 (N_11914,N_5499,N_7516);
or U11915 (N_11915,N_8138,N_5680);
nor U11916 (N_11916,N_9153,N_6250);
nand U11917 (N_11917,N_6593,N_5075);
nand U11918 (N_11918,N_8706,N_7753);
nand U11919 (N_11919,N_7127,N_9561);
nor U11920 (N_11920,N_9081,N_8681);
and U11921 (N_11921,N_5581,N_9213);
nor U11922 (N_11922,N_6155,N_5044);
and U11923 (N_11923,N_6702,N_6209);
or U11924 (N_11924,N_5787,N_6579);
nand U11925 (N_11925,N_6656,N_9175);
nor U11926 (N_11926,N_6746,N_6865);
nor U11927 (N_11927,N_5911,N_5290);
or U11928 (N_11928,N_6675,N_9948);
or U11929 (N_11929,N_8450,N_7646);
nor U11930 (N_11930,N_6639,N_8493);
and U11931 (N_11931,N_9147,N_8051);
nor U11932 (N_11932,N_7106,N_8018);
and U11933 (N_11933,N_8661,N_9157);
or U11934 (N_11934,N_5840,N_5863);
or U11935 (N_11935,N_6247,N_9577);
xor U11936 (N_11936,N_6793,N_5629);
xor U11937 (N_11937,N_7700,N_5887);
nand U11938 (N_11938,N_7723,N_9962);
nand U11939 (N_11939,N_6713,N_8238);
nand U11940 (N_11940,N_8044,N_8492);
and U11941 (N_11941,N_6449,N_9237);
and U11942 (N_11942,N_8755,N_6836);
and U11943 (N_11943,N_8663,N_6849);
and U11944 (N_11944,N_5414,N_6311);
and U11945 (N_11945,N_7339,N_7542);
nand U11946 (N_11946,N_5472,N_8930);
xor U11947 (N_11947,N_6451,N_9508);
or U11948 (N_11948,N_8221,N_5107);
and U11949 (N_11949,N_5202,N_6372);
xor U11950 (N_11950,N_5455,N_6305);
or U11951 (N_11951,N_7842,N_5003);
nand U11952 (N_11952,N_9503,N_5649);
or U11953 (N_11953,N_7384,N_9352);
and U11954 (N_11954,N_7785,N_8298);
xor U11955 (N_11955,N_6159,N_9596);
and U11956 (N_11956,N_9982,N_7310);
nor U11957 (N_11957,N_6930,N_8319);
or U11958 (N_11958,N_5770,N_8896);
xor U11959 (N_11959,N_7217,N_8301);
nand U11960 (N_11960,N_6598,N_5131);
nand U11961 (N_11961,N_8269,N_9507);
nor U11962 (N_11962,N_8682,N_6868);
or U11963 (N_11963,N_5004,N_6534);
nand U11964 (N_11964,N_9713,N_6425);
nor U11965 (N_11965,N_9937,N_6527);
nand U11966 (N_11966,N_9055,N_7942);
xor U11967 (N_11967,N_9922,N_6433);
nand U11968 (N_11968,N_8393,N_9027);
nand U11969 (N_11969,N_5595,N_6237);
or U11970 (N_11970,N_6714,N_6283);
xor U11971 (N_11971,N_6576,N_5509);
nand U11972 (N_11972,N_8948,N_8292);
nand U11973 (N_11973,N_7499,N_5551);
or U11974 (N_11974,N_8560,N_9437);
nand U11975 (N_11975,N_6171,N_8733);
and U11976 (N_11976,N_9450,N_5810);
nand U11977 (N_11977,N_7230,N_7902);
and U11978 (N_11978,N_5708,N_7599);
nand U11979 (N_11979,N_5977,N_6911);
or U11980 (N_11980,N_8331,N_7493);
or U11981 (N_11981,N_6685,N_6950);
xnor U11982 (N_11982,N_7272,N_9010);
nor U11983 (N_11983,N_6890,N_7858);
nand U11984 (N_11984,N_7579,N_7231);
nand U11985 (N_11985,N_5799,N_7637);
or U11986 (N_11986,N_7355,N_6374);
nand U11987 (N_11987,N_7471,N_5258);
or U11988 (N_11988,N_5491,N_7294);
nand U11989 (N_11989,N_7768,N_6140);
and U11990 (N_11990,N_9834,N_7199);
and U11991 (N_11991,N_9717,N_9378);
nand U11992 (N_11992,N_5720,N_9611);
or U11993 (N_11993,N_9402,N_8810);
nor U11994 (N_11994,N_9836,N_7577);
and U11995 (N_11995,N_5536,N_8893);
nand U11996 (N_11996,N_9614,N_7734);
xnor U11997 (N_11997,N_8384,N_6312);
nor U11998 (N_11998,N_9888,N_5159);
nor U11999 (N_11999,N_8121,N_9669);
or U12000 (N_12000,N_9809,N_6339);
nand U12001 (N_12001,N_7925,N_9578);
xnor U12002 (N_12002,N_5569,N_5644);
nand U12003 (N_12003,N_5288,N_6589);
nor U12004 (N_12004,N_6106,N_7631);
xor U12005 (N_12005,N_7451,N_7978);
nor U12006 (N_12006,N_8624,N_6468);
nor U12007 (N_12007,N_7820,N_8446);
and U12008 (N_12008,N_6740,N_5985);
nand U12009 (N_12009,N_6240,N_6214);
and U12010 (N_12010,N_9683,N_9022);
and U12011 (N_12011,N_6273,N_8177);
nand U12012 (N_12012,N_6794,N_6721);
nand U12013 (N_12013,N_7584,N_8524);
or U12014 (N_12014,N_7474,N_5877);
or U12015 (N_12015,N_7089,N_7979);
nor U12016 (N_12016,N_5726,N_8085);
nand U12017 (N_12017,N_7169,N_6591);
and U12018 (N_12018,N_7305,N_9997);
or U12019 (N_12019,N_5572,N_7815);
and U12020 (N_12020,N_8195,N_8909);
or U12021 (N_12021,N_9731,N_7197);
or U12022 (N_12022,N_5696,N_5263);
or U12023 (N_12023,N_8429,N_5494);
nor U12024 (N_12024,N_6325,N_8616);
nor U12025 (N_12025,N_5789,N_5603);
nand U12026 (N_12026,N_9276,N_5312);
nor U12027 (N_12027,N_6306,N_7635);
or U12028 (N_12028,N_7699,N_6738);
xnor U12029 (N_12029,N_7324,N_6926);
xnor U12030 (N_12030,N_6745,N_6308);
nor U12031 (N_12031,N_5382,N_7771);
nand U12032 (N_12032,N_6198,N_7277);
nand U12033 (N_12033,N_8198,N_6156);
and U12034 (N_12034,N_7196,N_6725);
nand U12035 (N_12035,N_7680,N_7079);
xnor U12036 (N_12036,N_8938,N_7251);
or U12037 (N_12037,N_5321,N_9349);
nand U12038 (N_12038,N_8538,N_7991);
nor U12039 (N_12039,N_5179,N_6365);
nor U12040 (N_12040,N_9638,N_6347);
nor U12041 (N_12041,N_9283,N_7604);
nor U12042 (N_12042,N_7172,N_9040);
nor U12043 (N_12043,N_5805,N_7852);
nor U12044 (N_12044,N_6399,N_9546);
and U12045 (N_12045,N_5446,N_6298);
or U12046 (N_12046,N_8884,N_9031);
nand U12047 (N_12047,N_7833,N_7639);
or U12048 (N_12048,N_7613,N_5332);
and U12049 (N_12049,N_8754,N_6341);
nand U12050 (N_12050,N_6683,N_5637);
and U12051 (N_12051,N_5056,N_6359);
xor U12052 (N_12052,N_7514,N_5988);
and U12053 (N_12053,N_8784,N_6265);
and U12054 (N_12054,N_6757,N_5427);
and U12055 (N_12055,N_8075,N_9206);
nand U12056 (N_12056,N_7993,N_9558);
or U12057 (N_12057,N_7547,N_5728);
and U12058 (N_12058,N_8216,N_9374);
and U12059 (N_12059,N_6420,N_5066);
or U12060 (N_12060,N_8297,N_7069);
nand U12061 (N_12061,N_8438,N_6068);
or U12062 (N_12062,N_6004,N_7527);
nor U12063 (N_12063,N_5392,N_8565);
or U12064 (N_12064,N_8833,N_9671);
and U12065 (N_12065,N_6938,N_8878);
and U12066 (N_12066,N_5474,N_7971);
and U12067 (N_12067,N_5448,N_5701);
or U12068 (N_12068,N_7354,N_9032);
nor U12069 (N_12069,N_6790,N_7096);
nor U12070 (N_12070,N_8608,N_6069);
xor U12071 (N_12071,N_9360,N_5338);
and U12072 (N_12072,N_5767,N_5431);
nand U12073 (N_12073,N_9432,N_5657);
nor U12074 (N_12074,N_5723,N_8515);
nand U12075 (N_12075,N_8346,N_9199);
nor U12076 (N_12076,N_8212,N_7097);
and U12077 (N_12077,N_6061,N_9012);
nand U12078 (N_12078,N_9993,N_6253);
or U12079 (N_12079,N_5866,N_6494);
and U12080 (N_12080,N_5351,N_5733);
xnor U12081 (N_12081,N_7176,N_7315);
nor U12082 (N_12082,N_7452,N_5768);
nor U12083 (N_12083,N_7226,N_6843);
nand U12084 (N_12084,N_7632,N_6825);
xor U12085 (N_12085,N_8949,N_8418);
nand U12086 (N_12086,N_7510,N_7174);
or U12087 (N_12087,N_7421,N_8157);
nor U12088 (N_12088,N_5929,N_8359);
or U12089 (N_12089,N_6737,N_6030);
and U12090 (N_12090,N_7309,N_7697);
or U12091 (N_12091,N_7040,N_9146);
xnor U12092 (N_12092,N_5058,N_8398);
or U12093 (N_12093,N_9598,N_5467);
or U12094 (N_12094,N_6320,N_5251);
and U12095 (N_12095,N_9967,N_6506);
nor U12096 (N_12096,N_5712,N_8294);
and U12097 (N_12097,N_6687,N_9412);
xor U12098 (N_12098,N_6601,N_9573);
nand U12099 (N_12099,N_5858,N_7297);
nand U12100 (N_12100,N_5736,N_6759);
nand U12101 (N_12101,N_7233,N_9917);
and U12102 (N_12102,N_8299,N_6133);
or U12103 (N_12103,N_8251,N_8305);
nor U12104 (N_12104,N_7811,N_5055);
or U12105 (N_12105,N_9607,N_8525);
and U12106 (N_12106,N_5074,N_9593);
or U12107 (N_12107,N_8350,N_9978);
or U12108 (N_12108,N_7498,N_7972);
nand U12109 (N_12109,N_5949,N_8282);
nand U12110 (N_12110,N_7129,N_7732);
or U12111 (N_12111,N_7962,N_7679);
nor U12112 (N_12112,N_5854,N_6160);
or U12113 (N_12113,N_9930,N_8213);
and U12114 (N_12114,N_8897,N_5033);
nand U12115 (N_12115,N_7567,N_8141);
and U12116 (N_12116,N_7861,N_9779);
or U12117 (N_12117,N_7202,N_5113);
xnor U12118 (N_12118,N_5487,N_8396);
nand U12119 (N_12119,N_6295,N_9004);
nand U12120 (N_12120,N_8573,N_8803);
nand U12121 (N_12121,N_6692,N_8445);
nand U12122 (N_12122,N_6128,N_8741);
nor U12123 (N_12123,N_6556,N_9527);
nand U12124 (N_12124,N_5859,N_8288);
nor U12125 (N_12125,N_6634,N_5702);
nand U12126 (N_12126,N_6202,N_9883);
or U12127 (N_12127,N_6317,N_6806);
nor U12128 (N_12128,N_9545,N_7509);
nor U12129 (N_12129,N_9693,N_5425);
xor U12130 (N_12130,N_7912,N_7957);
and U12131 (N_12131,N_6015,N_5289);
nor U12132 (N_12132,N_5070,N_6489);
and U12133 (N_12133,N_5684,N_9156);
or U12134 (N_12134,N_9485,N_6784);
and U12135 (N_12135,N_5784,N_8079);
xnor U12136 (N_12136,N_7203,N_8123);
and U12137 (N_12137,N_8160,N_7336);
xnor U12138 (N_12138,N_9250,N_6607);
and U12139 (N_12139,N_9851,N_7506);
and U12140 (N_12140,N_8283,N_9379);
or U12141 (N_12141,N_6879,N_5216);
nand U12142 (N_12142,N_7838,N_7478);
xor U12143 (N_12143,N_9451,N_9786);
and U12144 (N_12144,N_5452,N_6934);
and U12145 (N_12145,N_7397,N_5839);
and U12146 (N_12146,N_6667,N_7936);
and U12147 (N_12147,N_8797,N_5615);
and U12148 (N_12148,N_9315,N_5753);
nor U12149 (N_12149,N_6780,N_9818);
and U12150 (N_12150,N_8223,N_6800);
nor U12151 (N_12151,N_7976,N_6501);
and U12152 (N_12152,N_6050,N_9667);
xor U12153 (N_12153,N_9938,N_7243);
nor U12154 (N_12154,N_8338,N_5511);
xor U12155 (N_12155,N_5749,N_5405);
nor U12156 (N_12156,N_5229,N_9523);
nor U12157 (N_12157,N_5346,N_5867);
and U12158 (N_12158,N_5500,N_8711);
and U12159 (N_12159,N_9934,N_8224);
and U12160 (N_12160,N_7532,N_8178);
nand U12161 (N_12161,N_6467,N_5535);
xnor U12162 (N_12162,N_5831,N_7340);
or U12163 (N_12163,N_8939,N_8913);
or U12164 (N_12164,N_7551,N_7445);
or U12165 (N_12165,N_7955,N_9854);
nor U12166 (N_12166,N_7055,N_8574);
or U12167 (N_12167,N_7986,N_6281);
nor U12168 (N_12168,N_9648,N_6217);
and U12169 (N_12169,N_6419,N_5516);
nor U12170 (N_12170,N_6982,N_7591);
nand U12171 (N_12171,N_5729,N_7346);
or U12172 (N_12172,N_7592,N_9587);
nand U12173 (N_12173,N_7540,N_6473);
and U12174 (N_12174,N_7966,N_9472);
or U12175 (N_12175,N_7580,N_8924);
and U12176 (N_12176,N_9025,N_9063);
or U12177 (N_12177,N_9338,N_8068);
and U12178 (N_12178,N_7874,N_9048);
nor U12179 (N_12179,N_8705,N_9833);
nor U12180 (N_12180,N_6179,N_6970);
nand U12181 (N_12181,N_8580,N_8243);
and U12182 (N_12182,N_5292,N_9409);
or U12183 (N_12183,N_7871,N_9990);
xor U12184 (N_12184,N_8563,N_5388);
nand U12185 (N_12185,N_8029,N_7436);
nor U12186 (N_12186,N_7128,N_5306);
and U12187 (N_12187,N_9134,N_8110);
or U12188 (N_12188,N_5579,N_5246);
or U12189 (N_12189,N_5792,N_5477);
nand U12190 (N_12190,N_5525,N_8968);
or U12191 (N_12191,N_7288,N_7624);
or U12192 (N_12192,N_9483,N_8486);
nand U12193 (N_12193,N_9884,N_9606);
and U12194 (N_12194,N_7207,N_8850);
and U12195 (N_12195,N_8743,N_9257);
or U12196 (N_12196,N_9946,N_5022);
nand U12197 (N_12197,N_6199,N_8451);
nor U12198 (N_12198,N_7265,N_5666);
or U12199 (N_12199,N_6954,N_6262);
or U12200 (N_12200,N_8584,N_7769);
or U12201 (N_12201,N_9719,N_5486);
xor U12202 (N_12202,N_9610,N_8921);
nand U12203 (N_12203,N_6279,N_6697);
nor U12204 (N_12204,N_6246,N_8099);
and U12205 (N_12205,N_7045,N_7941);
nand U12206 (N_12206,N_7356,N_8337);
nand U12207 (N_12207,N_6493,N_6707);
nand U12208 (N_12208,N_7419,N_8648);
nor U12209 (N_12209,N_8342,N_7733);
nor U12210 (N_12210,N_6162,N_9066);
xnor U12211 (N_12211,N_5274,N_5255);
or U12212 (N_12212,N_8388,N_9112);
and U12213 (N_12213,N_6206,N_6726);
nor U12214 (N_12214,N_5842,N_8061);
and U12215 (N_12215,N_6518,N_9586);
or U12216 (N_12216,N_6747,N_6839);
or U12217 (N_12217,N_8256,N_9530);
or U12218 (N_12218,N_6137,N_5118);
and U12219 (N_12219,N_7429,N_6978);
xor U12220 (N_12220,N_9980,N_5094);
and U12221 (N_12221,N_5719,N_5959);
nor U12222 (N_12222,N_6352,N_8052);
or U12223 (N_12223,N_9789,N_9656);
nand U12224 (N_12224,N_5079,N_7104);
or U12225 (N_12225,N_6049,N_9430);
nor U12226 (N_12226,N_7809,N_9314);
nor U12227 (N_12227,N_7704,N_5968);
or U12228 (N_12228,N_5821,N_5137);
or U12229 (N_12229,N_7914,N_8824);
and U12230 (N_12230,N_7761,N_8098);
nand U12231 (N_12231,N_7762,N_7258);
xnor U12232 (N_12232,N_6411,N_8639);
and U12233 (N_12233,N_5116,N_5348);
nand U12234 (N_12234,N_6632,N_9308);
or U12235 (N_12235,N_8677,N_7968);
nor U12236 (N_12236,N_6609,N_5089);
nand U12237 (N_12237,N_5564,N_7913);
nor U12238 (N_12238,N_5287,N_7152);
nand U12239 (N_12239,N_6208,N_6979);
nand U12240 (N_12240,N_9998,N_6977);
or U12241 (N_12241,N_5752,N_9817);
nand U12242 (N_12242,N_7742,N_6383);
nand U12243 (N_12243,N_6136,N_9072);
and U12244 (N_12244,N_5636,N_7100);
xnor U12245 (N_12245,N_9209,N_9018);
or U12246 (N_12246,N_6177,N_8768);
or U12247 (N_12247,N_5670,N_9475);
and U12248 (N_12248,N_8228,N_7238);
nor U12249 (N_12249,N_6559,N_7965);
nor U12250 (N_12250,N_7798,N_7417);
nand U12251 (N_12251,N_7440,N_5412);
or U12252 (N_12252,N_7654,N_5982);
nor U12253 (N_12253,N_8496,N_5319);
nor U12254 (N_12254,N_8136,N_7570);
or U12255 (N_12255,N_7896,N_5460);
xor U12256 (N_12256,N_8602,N_8770);
nor U12257 (N_12257,N_7034,N_9677);
and U12258 (N_12258,N_5150,N_7764);
and U12259 (N_12259,N_7670,N_7530);
nor U12260 (N_12260,N_8006,N_7178);
nor U12261 (N_12261,N_7507,N_7796);
or U12262 (N_12262,N_6254,N_8962);
nand U12263 (N_12263,N_8906,N_7897);
nor U12264 (N_12264,N_9336,N_8472);
or U12265 (N_12265,N_7398,N_8154);
nor U12266 (N_12266,N_8022,N_7763);
nor U12267 (N_12267,N_5524,N_8696);
and U12268 (N_12268,N_6636,N_8208);
or U12269 (N_12269,N_6404,N_9664);
or U12270 (N_12270,N_5411,N_7774);
nand U12271 (N_12271,N_8004,N_7834);
nand U12272 (N_12272,N_9224,N_7007);
xnor U12273 (N_12273,N_5331,N_7223);
xnor U12274 (N_12274,N_8159,N_9608);
and U12275 (N_12275,N_8636,N_8951);
nand U12276 (N_12276,N_9404,N_6997);
and U12277 (N_12277,N_6550,N_7481);
nor U12278 (N_12278,N_7386,N_6178);
or U12279 (N_12279,N_6424,N_9142);
xnor U12280 (N_12280,N_7919,N_9852);
xnor U12281 (N_12281,N_7261,N_9829);
or U12282 (N_12282,N_6945,N_6920);
nor U12283 (N_12283,N_7270,N_7175);
nand U12284 (N_12284,N_6324,N_7455);
nor U12285 (N_12285,N_6981,N_7317);
nor U12286 (N_12286,N_7737,N_9288);
nor U12287 (N_12287,N_8820,N_6499);
nand U12288 (N_12288,N_8561,N_6637);
or U12289 (N_12289,N_8944,N_7138);
or U12290 (N_12290,N_9202,N_8442);
or U12291 (N_12291,N_8090,N_6477);
and U12292 (N_12292,N_6495,N_8659);
nand U12293 (N_12293,N_9070,N_7556);
nand U12294 (N_12294,N_6511,N_5240);
nand U12295 (N_12295,N_8400,N_8274);
and U12296 (N_12296,N_5962,N_7403);
or U12297 (N_12297,N_9585,N_8576);
nand U12298 (N_12298,N_9316,N_5659);
xor U12299 (N_12299,N_7804,N_6694);
or U12300 (N_12300,N_9054,N_8843);
or U12301 (N_12301,N_9133,N_8112);
nor U12302 (N_12302,N_8986,N_6613);
nand U12303 (N_12303,N_7843,N_7846);
and U12304 (N_12304,N_7496,N_8113);
nor U12305 (N_12305,N_9471,N_9396);
and U12306 (N_12306,N_5593,N_5592);
xnor U12307 (N_12307,N_9470,N_6213);
xnor U12308 (N_12308,N_7788,N_8627);
nand U12309 (N_12309,N_7035,N_5747);
xor U12310 (N_12310,N_8600,N_5078);
xnor U12311 (N_12311,N_8760,N_7601);
or U12312 (N_12312,N_6194,N_6490);
nor U12313 (N_12313,N_9660,N_9195);
nor U12314 (N_12314,N_7141,N_9539);
xnor U12315 (N_12315,N_7590,N_6932);
nor U12316 (N_12316,N_9337,N_6229);
xor U12317 (N_12317,N_7500,N_6545);
and U12318 (N_12318,N_8773,N_7412);
xor U12319 (N_12319,N_8352,N_7298);
or U12320 (N_12320,N_6196,N_5445);
or U12321 (N_12321,N_5937,N_8343);
or U12322 (N_12322,N_9434,N_6478);
nand U12323 (N_12323,N_7689,N_9392);
xor U12324 (N_12324,N_9595,N_8506);
xnor U12325 (N_12325,N_5082,N_9119);
or U12326 (N_12326,N_9984,N_5301);
and U12327 (N_12327,N_8116,N_7300);
and U12328 (N_12328,N_7952,N_7326);
nand U12329 (N_12329,N_5783,N_6315);
or U12330 (N_12330,N_8632,N_6211);
or U12331 (N_12331,N_6269,N_8805);
nand U12332 (N_12332,N_8700,N_9761);
nand U12333 (N_12333,N_6302,N_5940);
nand U12334 (N_12334,N_9532,N_9323);
or U12335 (N_12335,N_7171,N_6728);
xnor U12336 (N_12336,N_8527,N_5358);
or U12337 (N_12337,N_5506,N_9617);
nand U12338 (N_12338,N_8691,N_8078);
xor U12339 (N_12339,N_7868,N_9383);
xor U12340 (N_12340,N_7075,N_6624);
and U12341 (N_12341,N_6450,N_5129);
or U12342 (N_12342,N_9839,N_6652);
xnor U12343 (N_12343,N_5067,N_8071);
nor U12344 (N_12344,N_6884,N_8917);
and U12345 (N_12345,N_9908,N_6583);
xnor U12346 (N_12346,N_9905,N_7182);
xnor U12347 (N_12347,N_6035,N_5059);
nand U12348 (N_12348,N_5760,N_8839);
and U12349 (N_12349,N_6482,N_8723);
nor U12350 (N_12350,N_9515,N_8702);
nor U12351 (N_12351,N_8462,N_6923);
nor U12352 (N_12352,N_5847,N_9431);
or U12353 (N_12353,N_7603,N_9083);
nor U12354 (N_12354,N_7475,N_7024);
or U12355 (N_12355,N_5090,N_8424);
or U12356 (N_12356,N_5904,N_7320);
nor U12357 (N_12357,N_8311,N_7102);
and U12358 (N_12358,N_7856,N_6771);
or U12359 (N_12359,N_5104,N_7048);
and U12360 (N_12360,N_9039,N_7504);
nand U12361 (N_12361,N_9864,N_7405);
nor U12362 (N_12362,N_5291,N_9929);
xnor U12363 (N_12363,N_7794,N_5157);
xnor U12364 (N_12364,N_6164,N_6696);
nand U12365 (N_12365,N_7453,N_5507);
or U12366 (N_12366,N_9274,N_6659);
nor U12367 (N_12367,N_5270,N_5639);
xor U12368 (N_12368,N_6846,N_6442);
xor U12369 (N_12369,N_8807,N_8715);
nor U12370 (N_12370,N_5054,N_8270);
and U12371 (N_12371,N_9623,N_7713);
nor U12372 (N_12372,N_6248,N_8931);
and U12373 (N_12373,N_5943,N_6301);
nand U12374 (N_12374,N_7568,N_8132);
and U12375 (N_12375,N_9755,N_7111);
nand U12376 (N_12376,N_6023,N_8441);
or U12377 (N_12377,N_9932,N_8062);
and U12378 (N_12378,N_7928,N_8736);
nor U12379 (N_12379,N_7388,N_5087);
or U12380 (N_12380,N_8793,N_7112);
or U12381 (N_12381,N_5721,N_7844);
nor U12382 (N_12382,N_6485,N_8570);
and U12383 (N_12383,N_7192,N_5513);
nor U12384 (N_12384,N_7626,N_5030);
nor U12385 (N_12385,N_7557,N_6616);
or U12386 (N_12386,N_9168,N_8744);
nor U12387 (N_12387,N_8000,N_9255);
nand U12388 (N_12388,N_5252,N_8551);
xor U12389 (N_12389,N_7293,N_6939);
nor U12390 (N_12390,N_6417,N_8373);
nor U12391 (N_12391,N_6228,N_9806);
or U12392 (N_12392,N_7743,N_8009);
or U12393 (N_12393,N_6376,N_6650);
xor U12394 (N_12394,N_6385,N_5299);
and U12395 (N_12395,N_8792,N_7964);
and U12396 (N_12396,N_6293,N_8811);
and U12397 (N_12397,N_5379,N_8049);
and U12398 (N_12398,N_6628,N_9912);
xor U12399 (N_12399,N_8937,N_9413);
nor U12400 (N_12400,N_9582,N_9328);
nand U12401 (N_12401,N_7204,N_9183);
and U12402 (N_12402,N_7607,N_6439);
or U12403 (N_12403,N_9362,N_9197);
or U12404 (N_12404,N_9798,N_5517);
xnor U12405 (N_12405,N_6863,N_6664);
and U12406 (N_12406,N_5903,N_8808);
nand U12407 (N_12407,N_6500,N_6873);
and U12408 (N_12408,N_9969,N_8289);
nand U12409 (N_12409,N_5857,N_9442);
and U12410 (N_12410,N_9897,N_7267);
or U12411 (N_12411,N_7853,N_6698);
xor U12412 (N_12412,N_7108,N_5834);
xnor U12413 (N_12413,N_6504,N_7835);
nor U12414 (N_12414,N_9550,N_7458);
or U12415 (N_12415,N_7655,N_9979);
or U12416 (N_12416,N_5119,N_6823);
nand U12417 (N_12417,N_9957,N_9678);
nor U12418 (N_12418,N_6278,N_7373);
nand U12419 (N_12419,N_9243,N_5038);
and U12420 (N_12420,N_8555,N_6418);
and U12421 (N_12421,N_5010,N_5899);
nor U12422 (N_12422,N_5172,N_5328);
nor U12423 (N_12423,N_7092,N_9245);
and U12424 (N_12424,N_6259,N_6864);
and U12425 (N_12425,N_8528,N_7087);
nand U12426 (N_12426,N_5019,N_6431);
nand U12427 (N_12427,N_8203,N_5053);
nand U12428 (N_12428,N_8669,N_9254);
xnor U12429 (N_12429,N_9286,N_5234);
nor U12430 (N_12430,N_6407,N_6809);
or U12431 (N_12431,N_7735,N_5483);
nand U12432 (N_12432,N_5827,N_5142);
nor U12433 (N_12433,N_8932,N_7973);
xnor U12434 (N_12434,N_5835,N_5672);
nor U12435 (N_12435,N_7951,N_9390);
xnor U12436 (N_12436,N_7253,N_5797);
nand U12437 (N_12437,N_6165,N_6142);
and U12438 (N_12438,N_5048,N_9160);
nor U12439 (N_12439,N_6340,N_8487);
or U12440 (N_12440,N_6786,N_9075);
and U12441 (N_12441,N_5153,N_7899);
nand U12442 (N_12442,N_9291,N_6422);
nor U12443 (N_12443,N_9826,N_8187);
nand U12444 (N_12444,N_7546,N_7350);
or U12445 (N_12445,N_5254,N_7255);
nand U12446 (N_12446,N_7593,N_9757);
or U12447 (N_12447,N_8236,N_9856);
and U12448 (N_12448,N_6452,N_7206);
nor U12449 (N_12449,N_9725,N_9061);
and U12450 (N_12450,N_9584,N_9965);
nor U12451 (N_12451,N_8089,N_5562);
and U12452 (N_12452,N_5323,N_5343);
xnor U12453 (N_12453,N_9899,N_8983);
or U12454 (N_12454,N_6882,N_7779);
nor U12455 (N_12455,N_9524,N_5007);
nor U12456 (N_12456,N_5969,N_8306);
nand U12457 (N_12457,N_9367,N_7960);
or U12458 (N_12458,N_6681,N_7786);
nor U12459 (N_12459,N_7058,N_7142);
or U12460 (N_12460,N_9259,N_8470);
nor U12461 (N_12461,N_5141,N_7410);
and U12462 (N_12462,N_5091,N_9246);
or U12463 (N_12463,N_8056,N_6096);
or U12464 (N_12464,N_8738,N_6595);
nand U12465 (N_12465,N_7122,N_8601);
xor U12466 (N_12466,N_8680,N_9520);
xnor U12467 (N_12467,N_9302,N_8747);
or U12468 (N_12468,N_8271,N_8923);
nor U12469 (N_12469,N_5275,N_9919);
and U12470 (N_12470,N_9041,N_5996);
nand U12471 (N_12471,N_7154,N_8341);
or U12472 (N_12472,N_7375,N_9985);
nand U12473 (N_12473,N_7940,N_5161);
nor U12474 (N_12474,N_8104,N_8437);
nand U12475 (N_12475,N_8591,N_5876);
nand U12476 (N_12476,N_7998,N_9823);
and U12477 (N_12477,N_6928,N_9661);
xor U12478 (N_12478,N_5756,N_5280);
nand U12479 (N_12479,N_9599,N_6528);
and U12480 (N_12480,N_9087,N_6859);
xor U12481 (N_12481,N_6810,N_7039);
nand U12482 (N_12482,N_5553,N_6059);
nand U12483 (N_12483,N_9562,N_7997);
and U12484 (N_12484,N_6195,N_9949);
nor U12485 (N_12485,N_5861,N_8097);
nor U12486 (N_12486,N_5492,N_5688);
and U12487 (N_12487,N_5811,N_8873);
and U12488 (N_12488,N_5276,N_7760);
nand U12489 (N_12489,N_9935,N_6089);
and U12490 (N_12490,N_9371,N_7885);
or U12491 (N_12491,N_6744,N_8959);
or U12492 (N_12492,N_7916,N_7975);
and U12493 (N_12493,N_9440,N_9756);
and U12494 (N_12494,N_5724,N_7116);
nor U12495 (N_12495,N_5915,N_5844);
or U12496 (N_12496,N_7268,N_7361);
nand U12497 (N_12497,N_8325,N_8845);
nand U12498 (N_12498,N_9528,N_7020);
nor U12499 (N_12499,N_5126,N_7553);
nand U12500 (N_12500,N_9497,N_9841);
nand U12501 (N_12501,N_5546,N_9316);
or U12502 (N_12502,N_8818,N_6344);
and U12503 (N_12503,N_7376,N_7110);
nand U12504 (N_12504,N_9670,N_6011);
xor U12505 (N_12505,N_8186,N_8893);
or U12506 (N_12506,N_9305,N_9484);
or U12507 (N_12507,N_7072,N_9430);
nand U12508 (N_12508,N_9640,N_6330);
nand U12509 (N_12509,N_6900,N_6799);
and U12510 (N_12510,N_7913,N_6773);
nor U12511 (N_12511,N_9196,N_8902);
nor U12512 (N_12512,N_8899,N_8641);
nor U12513 (N_12513,N_5338,N_8748);
or U12514 (N_12514,N_8652,N_5677);
and U12515 (N_12515,N_7701,N_6459);
and U12516 (N_12516,N_9655,N_8974);
and U12517 (N_12517,N_9091,N_7740);
nor U12518 (N_12518,N_8901,N_6456);
nand U12519 (N_12519,N_9707,N_8569);
and U12520 (N_12520,N_8886,N_6341);
and U12521 (N_12521,N_8963,N_9777);
and U12522 (N_12522,N_8159,N_5507);
and U12523 (N_12523,N_7404,N_6834);
nand U12524 (N_12524,N_9264,N_6782);
nand U12525 (N_12525,N_6219,N_7659);
nand U12526 (N_12526,N_6004,N_9201);
xnor U12527 (N_12527,N_8762,N_9923);
and U12528 (N_12528,N_9026,N_8638);
nor U12529 (N_12529,N_9964,N_8728);
nor U12530 (N_12530,N_6936,N_5396);
and U12531 (N_12531,N_9122,N_9526);
or U12532 (N_12532,N_5805,N_5853);
nor U12533 (N_12533,N_5566,N_6853);
nand U12534 (N_12534,N_7607,N_6048);
nor U12535 (N_12535,N_8227,N_9588);
xnor U12536 (N_12536,N_6562,N_8491);
and U12537 (N_12537,N_6380,N_9731);
nor U12538 (N_12538,N_9600,N_9992);
or U12539 (N_12539,N_8781,N_7547);
or U12540 (N_12540,N_7970,N_8752);
nand U12541 (N_12541,N_5922,N_7055);
nor U12542 (N_12542,N_6148,N_7044);
xor U12543 (N_12543,N_6830,N_9773);
nor U12544 (N_12544,N_9334,N_7413);
or U12545 (N_12545,N_8507,N_9739);
xor U12546 (N_12546,N_9085,N_7835);
and U12547 (N_12547,N_6846,N_6228);
and U12548 (N_12548,N_6195,N_7743);
xnor U12549 (N_12549,N_8415,N_7455);
and U12550 (N_12550,N_9091,N_5012);
nand U12551 (N_12551,N_5082,N_5205);
and U12552 (N_12552,N_9114,N_9349);
xor U12553 (N_12553,N_9317,N_9099);
nor U12554 (N_12554,N_6898,N_6525);
xnor U12555 (N_12555,N_9179,N_9965);
xor U12556 (N_12556,N_9355,N_5674);
xor U12557 (N_12557,N_5377,N_9854);
nand U12558 (N_12558,N_7483,N_9423);
and U12559 (N_12559,N_5517,N_5468);
nand U12560 (N_12560,N_5563,N_8579);
nand U12561 (N_12561,N_6517,N_5623);
or U12562 (N_12562,N_6242,N_9158);
or U12563 (N_12563,N_7276,N_6710);
or U12564 (N_12564,N_5444,N_6419);
and U12565 (N_12565,N_7130,N_7300);
or U12566 (N_12566,N_9646,N_8186);
nand U12567 (N_12567,N_8857,N_9338);
nand U12568 (N_12568,N_7418,N_9176);
or U12569 (N_12569,N_5178,N_5582);
nor U12570 (N_12570,N_9637,N_8365);
and U12571 (N_12571,N_9602,N_5211);
xnor U12572 (N_12572,N_6018,N_8264);
nor U12573 (N_12573,N_7038,N_9127);
nand U12574 (N_12574,N_8395,N_7402);
and U12575 (N_12575,N_6369,N_6546);
and U12576 (N_12576,N_7448,N_8582);
nor U12577 (N_12577,N_5513,N_5559);
nor U12578 (N_12578,N_6819,N_7854);
xor U12579 (N_12579,N_6168,N_5362);
or U12580 (N_12580,N_5759,N_8279);
nor U12581 (N_12581,N_9052,N_7416);
xnor U12582 (N_12582,N_5871,N_7909);
or U12583 (N_12583,N_9983,N_6004);
nand U12584 (N_12584,N_8808,N_5862);
nand U12585 (N_12585,N_9518,N_9781);
and U12586 (N_12586,N_9491,N_9182);
or U12587 (N_12587,N_9791,N_9221);
xnor U12588 (N_12588,N_5638,N_8093);
or U12589 (N_12589,N_5136,N_5636);
and U12590 (N_12590,N_6401,N_7311);
nand U12591 (N_12591,N_5965,N_9566);
nor U12592 (N_12592,N_7019,N_6432);
nor U12593 (N_12593,N_8040,N_5190);
xnor U12594 (N_12594,N_8639,N_5226);
nor U12595 (N_12595,N_7474,N_7133);
nor U12596 (N_12596,N_6049,N_9284);
nand U12597 (N_12597,N_8639,N_8270);
and U12598 (N_12598,N_5102,N_9710);
and U12599 (N_12599,N_6850,N_6338);
xnor U12600 (N_12600,N_6736,N_9618);
nand U12601 (N_12601,N_7708,N_7951);
nor U12602 (N_12602,N_9856,N_9502);
and U12603 (N_12603,N_6934,N_6054);
or U12604 (N_12604,N_9581,N_8145);
nand U12605 (N_12605,N_5001,N_7828);
nor U12606 (N_12606,N_9676,N_5769);
nor U12607 (N_12607,N_9754,N_5755);
nand U12608 (N_12608,N_6119,N_5887);
or U12609 (N_12609,N_8786,N_7780);
nand U12610 (N_12610,N_8663,N_8800);
and U12611 (N_12611,N_9786,N_5334);
and U12612 (N_12612,N_9849,N_9087);
nor U12613 (N_12613,N_8439,N_6651);
or U12614 (N_12614,N_9005,N_5805);
and U12615 (N_12615,N_6534,N_9862);
nor U12616 (N_12616,N_7469,N_9668);
or U12617 (N_12617,N_6790,N_5651);
xor U12618 (N_12618,N_5569,N_8952);
nand U12619 (N_12619,N_9570,N_5348);
nand U12620 (N_12620,N_8880,N_9630);
nand U12621 (N_12621,N_9401,N_5667);
nor U12622 (N_12622,N_7083,N_8465);
or U12623 (N_12623,N_6600,N_9526);
or U12624 (N_12624,N_8038,N_7366);
and U12625 (N_12625,N_8669,N_9193);
and U12626 (N_12626,N_9205,N_9823);
nor U12627 (N_12627,N_9723,N_7309);
and U12628 (N_12628,N_6105,N_7390);
nand U12629 (N_12629,N_9055,N_6951);
nor U12630 (N_12630,N_6351,N_7350);
or U12631 (N_12631,N_7611,N_5410);
nor U12632 (N_12632,N_6594,N_9586);
nand U12633 (N_12633,N_7552,N_7918);
xnor U12634 (N_12634,N_5390,N_8263);
and U12635 (N_12635,N_7765,N_7508);
nand U12636 (N_12636,N_5714,N_8732);
xnor U12637 (N_12637,N_5942,N_7164);
nand U12638 (N_12638,N_9536,N_7632);
nand U12639 (N_12639,N_6290,N_6139);
nand U12640 (N_12640,N_5949,N_5147);
and U12641 (N_12641,N_6457,N_6724);
nor U12642 (N_12642,N_8878,N_5878);
xor U12643 (N_12643,N_5764,N_7342);
xor U12644 (N_12644,N_9042,N_8514);
nand U12645 (N_12645,N_9702,N_8258);
xor U12646 (N_12646,N_6688,N_5234);
or U12647 (N_12647,N_7021,N_8482);
or U12648 (N_12648,N_8982,N_7580);
or U12649 (N_12649,N_6783,N_9471);
or U12650 (N_12650,N_5860,N_9497);
and U12651 (N_12651,N_9161,N_5303);
and U12652 (N_12652,N_6173,N_5435);
nand U12653 (N_12653,N_8904,N_7447);
and U12654 (N_12654,N_5972,N_8356);
nand U12655 (N_12655,N_5636,N_7551);
or U12656 (N_12656,N_7364,N_5358);
nor U12657 (N_12657,N_5596,N_9659);
and U12658 (N_12658,N_6424,N_7121);
nor U12659 (N_12659,N_5149,N_7882);
or U12660 (N_12660,N_8760,N_6325);
nor U12661 (N_12661,N_8586,N_7894);
nor U12662 (N_12662,N_9616,N_7226);
xnor U12663 (N_12663,N_5187,N_5598);
and U12664 (N_12664,N_9774,N_6101);
or U12665 (N_12665,N_9975,N_5688);
and U12666 (N_12666,N_9529,N_5221);
or U12667 (N_12667,N_7382,N_5554);
xnor U12668 (N_12668,N_5554,N_5832);
nor U12669 (N_12669,N_6425,N_8723);
or U12670 (N_12670,N_8603,N_9416);
xor U12671 (N_12671,N_6005,N_8667);
or U12672 (N_12672,N_6683,N_9994);
nand U12673 (N_12673,N_6599,N_5834);
nand U12674 (N_12674,N_5413,N_8384);
and U12675 (N_12675,N_8405,N_5619);
or U12676 (N_12676,N_9439,N_6661);
or U12677 (N_12677,N_6195,N_9707);
nand U12678 (N_12678,N_6285,N_5966);
nor U12679 (N_12679,N_8975,N_8429);
or U12680 (N_12680,N_7634,N_8108);
nor U12681 (N_12681,N_8868,N_9148);
and U12682 (N_12682,N_9190,N_9326);
and U12683 (N_12683,N_7472,N_9996);
xnor U12684 (N_12684,N_6234,N_5541);
or U12685 (N_12685,N_6572,N_7405);
and U12686 (N_12686,N_5383,N_8806);
and U12687 (N_12687,N_9195,N_5574);
nor U12688 (N_12688,N_5280,N_7716);
nand U12689 (N_12689,N_9738,N_8231);
nor U12690 (N_12690,N_8667,N_6061);
or U12691 (N_12691,N_6757,N_6959);
and U12692 (N_12692,N_9044,N_6239);
nand U12693 (N_12693,N_6785,N_9373);
or U12694 (N_12694,N_8914,N_8641);
and U12695 (N_12695,N_5282,N_5653);
nor U12696 (N_12696,N_5286,N_9255);
nor U12697 (N_12697,N_7006,N_6141);
xor U12698 (N_12698,N_8684,N_7210);
or U12699 (N_12699,N_7658,N_9742);
or U12700 (N_12700,N_8095,N_7579);
xor U12701 (N_12701,N_8986,N_5758);
and U12702 (N_12702,N_8281,N_5209);
or U12703 (N_12703,N_5785,N_9777);
nand U12704 (N_12704,N_7229,N_5458);
or U12705 (N_12705,N_6072,N_6347);
nor U12706 (N_12706,N_8815,N_8954);
nand U12707 (N_12707,N_5915,N_6247);
or U12708 (N_12708,N_7301,N_8471);
nor U12709 (N_12709,N_8752,N_7061);
or U12710 (N_12710,N_6332,N_7249);
and U12711 (N_12711,N_6985,N_7231);
xor U12712 (N_12712,N_8688,N_6081);
and U12713 (N_12713,N_7156,N_7955);
and U12714 (N_12714,N_7859,N_8724);
and U12715 (N_12715,N_9482,N_9327);
nand U12716 (N_12716,N_9633,N_6246);
nand U12717 (N_12717,N_7300,N_5995);
nand U12718 (N_12718,N_6735,N_5276);
nor U12719 (N_12719,N_6733,N_5296);
nand U12720 (N_12720,N_7850,N_7617);
or U12721 (N_12721,N_5142,N_9203);
and U12722 (N_12722,N_7450,N_8008);
nand U12723 (N_12723,N_5526,N_8327);
or U12724 (N_12724,N_6993,N_5994);
xor U12725 (N_12725,N_9065,N_6436);
nor U12726 (N_12726,N_8481,N_5069);
xor U12727 (N_12727,N_5691,N_5150);
nand U12728 (N_12728,N_7193,N_6233);
xor U12729 (N_12729,N_7382,N_8043);
and U12730 (N_12730,N_6789,N_5048);
nor U12731 (N_12731,N_6407,N_7124);
nor U12732 (N_12732,N_5641,N_7003);
and U12733 (N_12733,N_6594,N_7015);
or U12734 (N_12734,N_9286,N_7183);
and U12735 (N_12735,N_5162,N_5645);
or U12736 (N_12736,N_8484,N_7257);
and U12737 (N_12737,N_5339,N_5426);
xnor U12738 (N_12738,N_7154,N_7371);
nor U12739 (N_12739,N_5757,N_9092);
or U12740 (N_12740,N_6571,N_5831);
nand U12741 (N_12741,N_8842,N_6287);
nand U12742 (N_12742,N_5016,N_8687);
or U12743 (N_12743,N_6896,N_9556);
xnor U12744 (N_12744,N_8229,N_8564);
nor U12745 (N_12745,N_9036,N_6237);
nor U12746 (N_12746,N_7215,N_5677);
nand U12747 (N_12747,N_8911,N_7083);
or U12748 (N_12748,N_5373,N_9576);
xnor U12749 (N_12749,N_5338,N_9184);
nand U12750 (N_12750,N_6651,N_8581);
nor U12751 (N_12751,N_9328,N_5097);
xor U12752 (N_12752,N_9282,N_7959);
nand U12753 (N_12753,N_9781,N_7484);
nand U12754 (N_12754,N_6877,N_5107);
nor U12755 (N_12755,N_8159,N_5550);
nand U12756 (N_12756,N_7684,N_6811);
nor U12757 (N_12757,N_6952,N_7388);
and U12758 (N_12758,N_9991,N_5646);
xor U12759 (N_12759,N_8221,N_8515);
nand U12760 (N_12760,N_7520,N_7689);
nand U12761 (N_12761,N_9133,N_7403);
nand U12762 (N_12762,N_7057,N_7040);
nand U12763 (N_12763,N_5868,N_5270);
and U12764 (N_12764,N_7403,N_6930);
nand U12765 (N_12765,N_7118,N_8784);
nor U12766 (N_12766,N_5210,N_5220);
or U12767 (N_12767,N_5746,N_7725);
xnor U12768 (N_12768,N_9896,N_8051);
or U12769 (N_12769,N_6606,N_9350);
and U12770 (N_12770,N_6075,N_5333);
nand U12771 (N_12771,N_8637,N_9999);
and U12772 (N_12772,N_9885,N_8644);
and U12773 (N_12773,N_8489,N_7620);
nand U12774 (N_12774,N_7867,N_9653);
or U12775 (N_12775,N_9965,N_6142);
or U12776 (N_12776,N_7885,N_7352);
nand U12777 (N_12777,N_8039,N_5941);
and U12778 (N_12778,N_5971,N_9088);
xnor U12779 (N_12779,N_9010,N_8762);
and U12780 (N_12780,N_5567,N_7120);
nand U12781 (N_12781,N_9103,N_6065);
nor U12782 (N_12782,N_6878,N_7925);
and U12783 (N_12783,N_9728,N_6855);
nor U12784 (N_12784,N_9133,N_7721);
or U12785 (N_12785,N_6609,N_8065);
nand U12786 (N_12786,N_7634,N_8224);
nand U12787 (N_12787,N_7084,N_8244);
and U12788 (N_12788,N_9992,N_9207);
or U12789 (N_12789,N_6845,N_7755);
and U12790 (N_12790,N_7524,N_9682);
or U12791 (N_12791,N_8815,N_5682);
and U12792 (N_12792,N_8293,N_6578);
nor U12793 (N_12793,N_8350,N_6270);
nor U12794 (N_12794,N_7317,N_8107);
nand U12795 (N_12795,N_6288,N_6044);
and U12796 (N_12796,N_9701,N_6615);
nand U12797 (N_12797,N_7479,N_9035);
nor U12798 (N_12798,N_6607,N_6106);
xnor U12799 (N_12799,N_7108,N_8407);
or U12800 (N_12800,N_8820,N_6764);
or U12801 (N_12801,N_7847,N_7804);
xor U12802 (N_12802,N_8685,N_9161);
and U12803 (N_12803,N_5394,N_8607);
nand U12804 (N_12804,N_9287,N_8407);
and U12805 (N_12805,N_6117,N_5805);
nor U12806 (N_12806,N_7017,N_8924);
nor U12807 (N_12807,N_8015,N_8086);
nor U12808 (N_12808,N_6689,N_9799);
and U12809 (N_12809,N_9509,N_9587);
nor U12810 (N_12810,N_6112,N_7723);
nand U12811 (N_12811,N_7591,N_7078);
or U12812 (N_12812,N_9851,N_6579);
nand U12813 (N_12813,N_9302,N_8424);
and U12814 (N_12814,N_9508,N_6132);
and U12815 (N_12815,N_7426,N_7017);
xor U12816 (N_12816,N_9042,N_7040);
and U12817 (N_12817,N_8087,N_6573);
nor U12818 (N_12818,N_7002,N_6731);
nor U12819 (N_12819,N_8761,N_9467);
or U12820 (N_12820,N_7987,N_6302);
nor U12821 (N_12821,N_8808,N_9262);
nor U12822 (N_12822,N_9243,N_6808);
nor U12823 (N_12823,N_9074,N_7950);
and U12824 (N_12824,N_6459,N_5603);
nand U12825 (N_12825,N_7243,N_5708);
nand U12826 (N_12826,N_5524,N_5712);
or U12827 (N_12827,N_8485,N_8540);
or U12828 (N_12828,N_5886,N_6100);
nand U12829 (N_12829,N_8772,N_9514);
or U12830 (N_12830,N_5082,N_6417);
or U12831 (N_12831,N_9489,N_6540);
nand U12832 (N_12832,N_5986,N_9437);
and U12833 (N_12833,N_7029,N_8043);
and U12834 (N_12834,N_6100,N_7064);
and U12835 (N_12835,N_5781,N_5141);
nand U12836 (N_12836,N_5335,N_6101);
nand U12837 (N_12837,N_5259,N_8140);
nor U12838 (N_12838,N_9211,N_9180);
nand U12839 (N_12839,N_6114,N_5687);
nand U12840 (N_12840,N_9829,N_9895);
nor U12841 (N_12841,N_6502,N_5438);
and U12842 (N_12842,N_8540,N_9760);
nand U12843 (N_12843,N_9530,N_6300);
or U12844 (N_12844,N_6307,N_8392);
nand U12845 (N_12845,N_8917,N_8179);
nor U12846 (N_12846,N_9807,N_5923);
nand U12847 (N_12847,N_6355,N_8152);
or U12848 (N_12848,N_6375,N_7939);
or U12849 (N_12849,N_8444,N_9619);
nor U12850 (N_12850,N_6911,N_6848);
xor U12851 (N_12851,N_9031,N_7956);
nand U12852 (N_12852,N_5964,N_5006);
or U12853 (N_12853,N_7971,N_5700);
and U12854 (N_12854,N_6412,N_5824);
nand U12855 (N_12855,N_9813,N_5619);
xnor U12856 (N_12856,N_6991,N_9885);
nand U12857 (N_12857,N_9137,N_9526);
xnor U12858 (N_12858,N_7396,N_8414);
or U12859 (N_12859,N_6734,N_8664);
and U12860 (N_12860,N_7294,N_8916);
or U12861 (N_12861,N_7871,N_9952);
or U12862 (N_12862,N_8736,N_8808);
or U12863 (N_12863,N_7929,N_5303);
nand U12864 (N_12864,N_9076,N_9271);
and U12865 (N_12865,N_9592,N_5606);
and U12866 (N_12866,N_5338,N_5559);
nor U12867 (N_12867,N_9787,N_7528);
or U12868 (N_12868,N_8187,N_5833);
nor U12869 (N_12869,N_9060,N_6593);
nand U12870 (N_12870,N_5028,N_5460);
and U12871 (N_12871,N_5750,N_6794);
or U12872 (N_12872,N_6293,N_8540);
or U12873 (N_12873,N_8108,N_9395);
or U12874 (N_12874,N_6595,N_5268);
or U12875 (N_12875,N_8878,N_7798);
and U12876 (N_12876,N_9339,N_9505);
nor U12877 (N_12877,N_9178,N_7994);
nand U12878 (N_12878,N_6216,N_9295);
or U12879 (N_12879,N_7318,N_7173);
and U12880 (N_12880,N_5803,N_7903);
nand U12881 (N_12881,N_6416,N_9639);
and U12882 (N_12882,N_5939,N_5043);
nor U12883 (N_12883,N_7923,N_9287);
nor U12884 (N_12884,N_7316,N_7928);
xor U12885 (N_12885,N_9735,N_5421);
or U12886 (N_12886,N_6547,N_7560);
nand U12887 (N_12887,N_7141,N_5489);
xnor U12888 (N_12888,N_7735,N_7693);
or U12889 (N_12889,N_9148,N_8475);
nand U12890 (N_12890,N_6783,N_9101);
and U12891 (N_12891,N_8278,N_7647);
and U12892 (N_12892,N_6582,N_7666);
nand U12893 (N_12893,N_6749,N_9175);
nor U12894 (N_12894,N_7198,N_9426);
nand U12895 (N_12895,N_7915,N_8311);
xnor U12896 (N_12896,N_6223,N_6956);
or U12897 (N_12897,N_9227,N_6908);
nand U12898 (N_12898,N_6527,N_6782);
and U12899 (N_12899,N_5582,N_6154);
and U12900 (N_12900,N_8865,N_5239);
or U12901 (N_12901,N_5994,N_5871);
nand U12902 (N_12902,N_6198,N_6290);
and U12903 (N_12903,N_8681,N_9104);
nor U12904 (N_12904,N_9286,N_5117);
nand U12905 (N_12905,N_5857,N_7978);
or U12906 (N_12906,N_8839,N_5342);
xnor U12907 (N_12907,N_6610,N_8517);
or U12908 (N_12908,N_6019,N_8769);
or U12909 (N_12909,N_6082,N_9853);
and U12910 (N_12910,N_7347,N_6331);
or U12911 (N_12911,N_5849,N_9398);
nand U12912 (N_12912,N_5444,N_8175);
or U12913 (N_12913,N_9203,N_9524);
and U12914 (N_12914,N_6196,N_9034);
and U12915 (N_12915,N_7432,N_7881);
or U12916 (N_12916,N_5152,N_6714);
nand U12917 (N_12917,N_7318,N_9960);
or U12918 (N_12918,N_8163,N_7291);
nand U12919 (N_12919,N_8670,N_8240);
or U12920 (N_12920,N_6053,N_9340);
nor U12921 (N_12921,N_5589,N_6701);
or U12922 (N_12922,N_5001,N_5157);
nand U12923 (N_12923,N_8040,N_9045);
nand U12924 (N_12924,N_8676,N_6337);
nand U12925 (N_12925,N_6071,N_9857);
nor U12926 (N_12926,N_8953,N_6438);
or U12927 (N_12927,N_7468,N_8203);
nor U12928 (N_12928,N_9007,N_9027);
xor U12929 (N_12929,N_9310,N_8082);
and U12930 (N_12930,N_8927,N_9228);
nand U12931 (N_12931,N_5714,N_8419);
nor U12932 (N_12932,N_9174,N_5061);
and U12933 (N_12933,N_5529,N_6191);
xnor U12934 (N_12934,N_6680,N_5014);
nand U12935 (N_12935,N_7864,N_9127);
nor U12936 (N_12936,N_5404,N_9747);
and U12937 (N_12937,N_6189,N_7819);
nand U12938 (N_12938,N_8865,N_6326);
xor U12939 (N_12939,N_5382,N_7279);
and U12940 (N_12940,N_7259,N_5288);
nor U12941 (N_12941,N_5656,N_8725);
and U12942 (N_12942,N_5016,N_6941);
or U12943 (N_12943,N_9356,N_8062);
nor U12944 (N_12944,N_5285,N_5731);
or U12945 (N_12945,N_5822,N_9700);
or U12946 (N_12946,N_7501,N_8403);
nor U12947 (N_12947,N_5537,N_9721);
and U12948 (N_12948,N_5899,N_6166);
or U12949 (N_12949,N_6767,N_7857);
nor U12950 (N_12950,N_9511,N_9399);
nor U12951 (N_12951,N_6687,N_8904);
xor U12952 (N_12952,N_5442,N_8591);
and U12953 (N_12953,N_8934,N_8654);
nand U12954 (N_12954,N_8457,N_9807);
nand U12955 (N_12955,N_8216,N_7898);
xnor U12956 (N_12956,N_9982,N_9359);
and U12957 (N_12957,N_9498,N_7468);
and U12958 (N_12958,N_7419,N_7737);
or U12959 (N_12959,N_9513,N_5649);
and U12960 (N_12960,N_8111,N_5839);
or U12961 (N_12961,N_7902,N_7469);
nand U12962 (N_12962,N_8181,N_8272);
and U12963 (N_12963,N_5304,N_5602);
or U12964 (N_12964,N_7710,N_6102);
and U12965 (N_12965,N_7940,N_6056);
and U12966 (N_12966,N_5253,N_8009);
and U12967 (N_12967,N_7130,N_9207);
nor U12968 (N_12968,N_8114,N_8928);
nor U12969 (N_12969,N_7336,N_6939);
nor U12970 (N_12970,N_5926,N_5430);
or U12971 (N_12971,N_8272,N_9093);
nand U12972 (N_12972,N_5482,N_7293);
nand U12973 (N_12973,N_6114,N_5999);
nand U12974 (N_12974,N_8749,N_9872);
xor U12975 (N_12975,N_7069,N_7413);
xnor U12976 (N_12976,N_7978,N_9210);
or U12977 (N_12977,N_8470,N_9247);
nor U12978 (N_12978,N_9774,N_7071);
and U12979 (N_12979,N_7902,N_7149);
nand U12980 (N_12980,N_7436,N_6762);
xnor U12981 (N_12981,N_6552,N_5920);
and U12982 (N_12982,N_7025,N_8615);
or U12983 (N_12983,N_9715,N_6947);
nor U12984 (N_12984,N_6813,N_9423);
nor U12985 (N_12985,N_5758,N_9747);
and U12986 (N_12986,N_5198,N_9279);
and U12987 (N_12987,N_8572,N_5479);
nor U12988 (N_12988,N_9869,N_6928);
xnor U12989 (N_12989,N_5502,N_7066);
nor U12990 (N_12990,N_7517,N_8625);
or U12991 (N_12991,N_6249,N_8997);
or U12992 (N_12992,N_5365,N_7676);
nand U12993 (N_12993,N_5109,N_8374);
and U12994 (N_12994,N_9609,N_7186);
and U12995 (N_12995,N_9881,N_9107);
nor U12996 (N_12996,N_9925,N_7845);
and U12997 (N_12997,N_6870,N_9551);
nor U12998 (N_12998,N_6930,N_7692);
xor U12999 (N_12999,N_6352,N_7002);
nand U13000 (N_13000,N_7366,N_5993);
or U13001 (N_13001,N_9436,N_8400);
nor U13002 (N_13002,N_5190,N_7657);
xor U13003 (N_13003,N_8641,N_5281);
and U13004 (N_13004,N_6742,N_6678);
and U13005 (N_13005,N_5831,N_7581);
nor U13006 (N_13006,N_8518,N_5473);
nand U13007 (N_13007,N_7011,N_9430);
or U13008 (N_13008,N_5353,N_7599);
and U13009 (N_13009,N_6149,N_5866);
and U13010 (N_13010,N_5421,N_9527);
and U13011 (N_13011,N_8028,N_5425);
nor U13012 (N_13012,N_7289,N_7319);
nand U13013 (N_13013,N_6992,N_9560);
nand U13014 (N_13014,N_8417,N_6523);
and U13015 (N_13015,N_7914,N_5651);
nor U13016 (N_13016,N_6974,N_9539);
nor U13017 (N_13017,N_6616,N_6437);
and U13018 (N_13018,N_7273,N_5589);
nor U13019 (N_13019,N_8008,N_8034);
and U13020 (N_13020,N_8454,N_9039);
and U13021 (N_13021,N_8586,N_5939);
or U13022 (N_13022,N_8634,N_9659);
nor U13023 (N_13023,N_7072,N_5260);
nand U13024 (N_13024,N_6882,N_7730);
nand U13025 (N_13025,N_5680,N_6123);
nand U13026 (N_13026,N_7898,N_5943);
nand U13027 (N_13027,N_6939,N_9364);
nor U13028 (N_13028,N_6158,N_6806);
xor U13029 (N_13029,N_8319,N_8776);
and U13030 (N_13030,N_8021,N_5930);
and U13031 (N_13031,N_5873,N_9171);
and U13032 (N_13032,N_6716,N_6638);
or U13033 (N_13033,N_7298,N_8189);
nand U13034 (N_13034,N_7056,N_6765);
nand U13035 (N_13035,N_7857,N_9588);
or U13036 (N_13036,N_8005,N_9602);
and U13037 (N_13037,N_8640,N_9619);
xor U13038 (N_13038,N_8678,N_7903);
and U13039 (N_13039,N_8342,N_7325);
and U13040 (N_13040,N_6143,N_5373);
xnor U13041 (N_13041,N_5477,N_8705);
nor U13042 (N_13042,N_6597,N_8733);
or U13043 (N_13043,N_9654,N_8076);
and U13044 (N_13044,N_7244,N_5705);
and U13045 (N_13045,N_7211,N_9669);
and U13046 (N_13046,N_8923,N_6492);
nor U13047 (N_13047,N_6720,N_5263);
nand U13048 (N_13048,N_7378,N_5934);
or U13049 (N_13049,N_6273,N_7087);
or U13050 (N_13050,N_6894,N_9911);
nand U13051 (N_13051,N_5688,N_7558);
nand U13052 (N_13052,N_6844,N_6138);
xor U13053 (N_13053,N_7531,N_5711);
nor U13054 (N_13054,N_9417,N_8939);
xor U13055 (N_13055,N_7648,N_5765);
nor U13056 (N_13056,N_7550,N_5687);
nand U13057 (N_13057,N_9380,N_5625);
and U13058 (N_13058,N_8460,N_9298);
or U13059 (N_13059,N_9984,N_9027);
and U13060 (N_13060,N_5579,N_5488);
or U13061 (N_13061,N_7945,N_6470);
nor U13062 (N_13062,N_6560,N_9455);
nor U13063 (N_13063,N_8383,N_6754);
nor U13064 (N_13064,N_9533,N_9323);
or U13065 (N_13065,N_5494,N_5124);
nor U13066 (N_13066,N_8283,N_7929);
and U13067 (N_13067,N_5239,N_7414);
xnor U13068 (N_13068,N_7486,N_6724);
nor U13069 (N_13069,N_5431,N_8907);
nor U13070 (N_13070,N_6883,N_7072);
xnor U13071 (N_13071,N_9073,N_5090);
and U13072 (N_13072,N_7196,N_9813);
nand U13073 (N_13073,N_9013,N_5617);
xor U13074 (N_13074,N_9546,N_6362);
or U13075 (N_13075,N_9639,N_5387);
nand U13076 (N_13076,N_8776,N_9200);
and U13077 (N_13077,N_5619,N_8345);
nor U13078 (N_13078,N_5852,N_5389);
or U13079 (N_13079,N_9181,N_5156);
nand U13080 (N_13080,N_6190,N_8248);
nand U13081 (N_13081,N_7922,N_8630);
nor U13082 (N_13082,N_8830,N_9477);
or U13083 (N_13083,N_5180,N_8747);
nor U13084 (N_13084,N_7042,N_6430);
nand U13085 (N_13085,N_6755,N_6447);
or U13086 (N_13086,N_9150,N_6271);
nand U13087 (N_13087,N_9198,N_6461);
or U13088 (N_13088,N_7965,N_8440);
nand U13089 (N_13089,N_8258,N_6870);
and U13090 (N_13090,N_5823,N_8358);
or U13091 (N_13091,N_9177,N_6454);
nor U13092 (N_13092,N_7122,N_7083);
or U13093 (N_13093,N_9778,N_9418);
and U13094 (N_13094,N_5041,N_5321);
nor U13095 (N_13095,N_8111,N_6934);
and U13096 (N_13096,N_7462,N_9265);
nor U13097 (N_13097,N_9973,N_5015);
nor U13098 (N_13098,N_8484,N_8221);
nand U13099 (N_13099,N_7236,N_5357);
and U13100 (N_13100,N_7491,N_9865);
nor U13101 (N_13101,N_7081,N_7770);
or U13102 (N_13102,N_7628,N_9284);
nand U13103 (N_13103,N_8619,N_6972);
and U13104 (N_13104,N_8456,N_9280);
nor U13105 (N_13105,N_7818,N_9700);
and U13106 (N_13106,N_7119,N_7836);
nor U13107 (N_13107,N_9923,N_9415);
xnor U13108 (N_13108,N_9815,N_6731);
or U13109 (N_13109,N_5733,N_5208);
nor U13110 (N_13110,N_7602,N_6472);
nor U13111 (N_13111,N_7722,N_8246);
and U13112 (N_13112,N_9581,N_7128);
and U13113 (N_13113,N_8234,N_6372);
or U13114 (N_13114,N_6045,N_9063);
nor U13115 (N_13115,N_9282,N_8857);
and U13116 (N_13116,N_8294,N_9753);
or U13117 (N_13117,N_6040,N_5714);
or U13118 (N_13118,N_6281,N_8973);
nand U13119 (N_13119,N_5755,N_8154);
or U13120 (N_13120,N_5838,N_5478);
nand U13121 (N_13121,N_5191,N_8099);
nand U13122 (N_13122,N_6839,N_8179);
nor U13123 (N_13123,N_8996,N_7324);
nor U13124 (N_13124,N_5554,N_9972);
nor U13125 (N_13125,N_9728,N_7025);
and U13126 (N_13126,N_6541,N_5868);
nand U13127 (N_13127,N_7527,N_8378);
xnor U13128 (N_13128,N_8796,N_5486);
nor U13129 (N_13129,N_9069,N_6292);
nor U13130 (N_13130,N_7986,N_7757);
nor U13131 (N_13131,N_9476,N_8537);
nor U13132 (N_13132,N_5624,N_6755);
and U13133 (N_13133,N_6081,N_8663);
or U13134 (N_13134,N_9383,N_6430);
nand U13135 (N_13135,N_8096,N_8474);
or U13136 (N_13136,N_7669,N_9444);
xnor U13137 (N_13137,N_9140,N_6373);
or U13138 (N_13138,N_8787,N_9686);
nand U13139 (N_13139,N_6502,N_9210);
nand U13140 (N_13140,N_9031,N_6922);
nand U13141 (N_13141,N_8360,N_5634);
and U13142 (N_13142,N_9809,N_6882);
or U13143 (N_13143,N_5158,N_7828);
and U13144 (N_13144,N_6838,N_8618);
nor U13145 (N_13145,N_6574,N_5560);
nor U13146 (N_13146,N_8408,N_7609);
xor U13147 (N_13147,N_6018,N_6016);
nand U13148 (N_13148,N_7806,N_5508);
xor U13149 (N_13149,N_8825,N_6891);
xor U13150 (N_13150,N_8418,N_5438);
nor U13151 (N_13151,N_6875,N_7023);
xor U13152 (N_13152,N_6960,N_7383);
nor U13153 (N_13153,N_8072,N_5995);
nor U13154 (N_13154,N_7294,N_5714);
nand U13155 (N_13155,N_9998,N_9281);
or U13156 (N_13156,N_9913,N_5094);
xor U13157 (N_13157,N_7959,N_9740);
or U13158 (N_13158,N_8523,N_7853);
nor U13159 (N_13159,N_7560,N_6158);
nand U13160 (N_13160,N_6364,N_8054);
nor U13161 (N_13161,N_8643,N_5044);
nor U13162 (N_13162,N_7522,N_6083);
nor U13163 (N_13163,N_6287,N_9422);
nand U13164 (N_13164,N_8414,N_6489);
or U13165 (N_13165,N_5971,N_7922);
nand U13166 (N_13166,N_8068,N_9392);
nand U13167 (N_13167,N_6418,N_5448);
and U13168 (N_13168,N_7653,N_5369);
xnor U13169 (N_13169,N_9663,N_8584);
nand U13170 (N_13170,N_6139,N_9910);
and U13171 (N_13171,N_9280,N_8578);
and U13172 (N_13172,N_6459,N_6719);
xor U13173 (N_13173,N_7950,N_9664);
or U13174 (N_13174,N_9830,N_6873);
nand U13175 (N_13175,N_9349,N_5510);
and U13176 (N_13176,N_7596,N_6947);
nand U13177 (N_13177,N_7773,N_7424);
or U13178 (N_13178,N_8113,N_9950);
and U13179 (N_13179,N_9673,N_7371);
nor U13180 (N_13180,N_9214,N_7457);
and U13181 (N_13181,N_6372,N_6434);
or U13182 (N_13182,N_9929,N_5297);
and U13183 (N_13183,N_8364,N_5850);
nor U13184 (N_13184,N_6580,N_8686);
or U13185 (N_13185,N_8263,N_9393);
or U13186 (N_13186,N_9907,N_9074);
and U13187 (N_13187,N_8368,N_5031);
and U13188 (N_13188,N_5123,N_8594);
nand U13189 (N_13189,N_7311,N_8056);
or U13190 (N_13190,N_9675,N_5831);
nand U13191 (N_13191,N_9857,N_8538);
or U13192 (N_13192,N_9720,N_6798);
nand U13193 (N_13193,N_5078,N_7380);
nor U13194 (N_13194,N_7948,N_5677);
and U13195 (N_13195,N_8531,N_9648);
or U13196 (N_13196,N_7315,N_8345);
nor U13197 (N_13197,N_7053,N_7303);
xor U13198 (N_13198,N_6611,N_9684);
nand U13199 (N_13199,N_6277,N_9504);
nand U13200 (N_13200,N_6910,N_8172);
nor U13201 (N_13201,N_9793,N_6092);
or U13202 (N_13202,N_9003,N_5647);
xnor U13203 (N_13203,N_5217,N_6324);
nand U13204 (N_13204,N_6602,N_9802);
or U13205 (N_13205,N_7999,N_6955);
nand U13206 (N_13206,N_9504,N_9286);
nor U13207 (N_13207,N_9222,N_5671);
nor U13208 (N_13208,N_6967,N_7440);
or U13209 (N_13209,N_6489,N_8654);
nor U13210 (N_13210,N_5972,N_8987);
or U13211 (N_13211,N_8685,N_8946);
nand U13212 (N_13212,N_6735,N_7761);
or U13213 (N_13213,N_9934,N_5832);
nand U13214 (N_13214,N_6720,N_7124);
nor U13215 (N_13215,N_5907,N_6976);
nor U13216 (N_13216,N_6964,N_6705);
nor U13217 (N_13217,N_5411,N_8621);
and U13218 (N_13218,N_7870,N_6373);
xor U13219 (N_13219,N_8180,N_9977);
nand U13220 (N_13220,N_6576,N_9854);
nand U13221 (N_13221,N_5057,N_9949);
nor U13222 (N_13222,N_6664,N_9849);
nor U13223 (N_13223,N_8443,N_6516);
or U13224 (N_13224,N_8060,N_7903);
or U13225 (N_13225,N_7871,N_9370);
nor U13226 (N_13226,N_5661,N_5975);
and U13227 (N_13227,N_6317,N_8685);
nor U13228 (N_13228,N_7753,N_9494);
nor U13229 (N_13229,N_5838,N_6756);
or U13230 (N_13230,N_7663,N_5649);
or U13231 (N_13231,N_8336,N_8619);
and U13232 (N_13232,N_6512,N_8892);
and U13233 (N_13233,N_9955,N_8142);
nand U13234 (N_13234,N_9494,N_5492);
xnor U13235 (N_13235,N_8932,N_7721);
nand U13236 (N_13236,N_5480,N_7099);
nand U13237 (N_13237,N_9757,N_5620);
nand U13238 (N_13238,N_9864,N_5049);
xnor U13239 (N_13239,N_6416,N_7425);
nor U13240 (N_13240,N_7901,N_7103);
and U13241 (N_13241,N_8742,N_6188);
nor U13242 (N_13242,N_9241,N_5334);
nor U13243 (N_13243,N_6800,N_5731);
and U13244 (N_13244,N_6742,N_8923);
and U13245 (N_13245,N_8425,N_5795);
and U13246 (N_13246,N_8890,N_7635);
nor U13247 (N_13247,N_6767,N_7517);
nand U13248 (N_13248,N_6300,N_7135);
and U13249 (N_13249,N_9875,N_8372);
nor U13250 (N_13250,N_7963,N_6635);
nand U13251 (N_13251,N_7113,N_5400);
nand U13252 (N_13252,N_9063,N_7909);
and U13253 (N_13253,N_7352,N_5481);
nor U13254 (N_13254,N_6137,N_5336);
xor U13255 (N_13255,N_9020,N_5287);
nor U13256 (N_13256,N_6479,N_5766);
xor U13257 (N_13257,N_6446,N_5008);
nor U13258 (N_13258,N_5294,N_5145);
xor U13259 (N_13259,N_5643,N_8033);
or U13260 (N_13260,N_9707,N_8274);
or U13261 (N_13261,N_9771,N_6443);
nand U13262 (N_13262,N_9793,N_7443);
and U13263 (N_13263,N_5438,N_8868);
or U13264 (N_13264,N_7427,N_5805);
nor U13265 (N_13265,N_7520,N_9679);
nand U13266 (N_13266,N_5347,N_8796);
nand U13267 (N_13267,N_5692,N_7558);
or U13268 (N_13268,N_5530,N_8996);
nor U13269 (N_13269,N_8399,N_6598);
nand U13270 (N_13270,N_7764,N_9017);
or U13271 (N_13271,N_9679,N_9038);
nand U13272 (N_13272,N_6122,N_7897);
nor U13273 (N_13273,N_5359,N_8426);
nand U13274 (N_13274,N_9294,N_6810);
or U13275 (N_13275,N_8199,N_9017);
or U13276 (N_13276,N_6272,N_7406);
or U13277 (N_13277,N_5577,N_8038);
nor U13278 (N_13278,N_6456,N_8167);
or U13279 (N_13279,N_8427,N_9145);
nor U13280 (N_13280,N_5044,N_6971);
or U13281 (N_13281,N_6522,N_8741);
nand U13282 (N_13282,N_7153,N_8826);
or U13283 (N_13283,N_7974,N_6949);
nor U13284 (N_13284,N_9880,N_5399);
and U13285 (N_13285,N_9755,N_9753);
nor U13286 (N_13286,N_9199,N_9803);
or U13287 (N_13287,N_9080,N_9992);
nand U13288 (N_13288,N_6553,N_5014);
nor U13289 (N_13289,N_8008,N_9976);
and U13290 (N_13290,N_6110,N_7163);
or U13291 (N_13291,N_7365,N_8250);
or U13292 (N_13292,N_9655,N_6789);
and U13293 (N_13293,N_6380,N_5343);
xor U13294 (N_13294,N_6534,N_8165);
nand U13295 (N_13295,N_5941,N_5188);
and U13296 (N_13296,N_7613,N_7188);
and U13297 (N_13297,N_9984,N_6218);
nand U13298 (N_13298,N_5854,N_7251);
nand U13299 (N_13299,N_8846,N_9717);
nor U13300 (N_13300,N_6442,N_9066);
or U13301 (N_13301,N_8654,N_6259);
xnor U13302 (N_13302,N_9889,N_5899);
xnor U13303 (N_13303,N_8104,N_8143);
xor U13304 (N_13304,N_8706,N_6590);
or U13305 (N_13305,N_6811,N_6372);
or U13306 (N_13306,N_5297,N_7255);
xnor U13307 (N_13307,N_8136,N_5175);
nand U13308 (N_13308,N_7841,N_7761);
nand U13309 (N_13309,N_9758,N_6241);
and U13310 (N_13310,N_6251,N_6358);
nand U13311 (N_13311,N_5631,N_5355);
and U13312 (N_13312,N_6225,N_5980);
nor U13313 (N_13313,N_6937,N_8544);
or U13314 (N_13314,N_8204,N_8954);
nand U13315 (N_13315,N_7788,N_6350);
or U13316 (N_13316,N_5649,N_9349);
and U13317 (N_13317,N_9777,N_7879);
or U13318 (N_13318,N_6978,N_6504);
nand U13319 (N_13319,N_8832,N_7126);
and U13320 (N_13320,N_9013,N_8984);
xor U13321 (N_13321,N_5148,N_5975);
and U13322 (N_13322,N_7737,N_7616);
nor U13323 (N_13323,N_8307,N_9675);
nor U13324 (N_13324,N_8555,N_7036);
nor U13325 (N_13325,N_8044,N_6810);
or U13326 (N_13326,N_9430,N_6352);
nand U13327 (N_13327,N_8267,N_9021);
or U13328 (N_13328,N_9483,N_9545);
xnor U13329 (N_13329,N_6634,N_9651);
nand U13330 (N_13330,N_9981,N_7245);
and U13331 (N_13331,N_5293,N_5967);
or U13332 (N_13332,N_8987,N_9751);
and U13333 (N_13333,N_5323,N_6353);
nor U13334 (N_13334,N_9335,N_9974);
nand U13335 (N_13335,N_7631,N_8860);
or U13336 (N_13336,N_9673,N_6198);
and U13337 (N_13337,N_5240,N_7929);
and U13338 (N_13338,N_8478,N_7943);
xnor U13339 (N_13339,N_6459,N_7312);
or U13340 (N_13340,N_9249,N_9043);
nor U13341 (N_13341,N_5480,N_7505);
and U13342 (N_13342,N_6928,N_5163);
nor U13343 (N_13343,N_5934,N_6768);
and U13344 (N_13344,N_8573,N_6817);
or U13345 (N_13345,N_8920,N_6699);
xor U13346 (N_13346,N_7152,N_8712);
or U13347 (N_13347,N_6795,N_9753);
or U13348 (N_13348,N_8686,N_5448);
and U13349 (N_13349,N_5675,N_9432);
xor U13350 (N_13350,N_9722,N_7817);
nand U13351 (N_13351,N_5250,N_7364);
nor U13352 (N_13352,N_7566,N_9633);
nor U13353 (N_13353,N_6548,N_7289);
or U13354 (N_13354,N_8243,N_8949);
xnor U13355 (N_13355,N_8050,N_6948);
nand U13356 (N_13356,N_9044,N_8883);
nand U13357 (N_13357,N_8694,N_9428);
or U13358 (N_13358,N_8690,N_8865);
nand U13359 (N_13359,N_6293,N_8675);
and U13360 (N_13360,N_9927,N_6609);
nor U13361 (N_13361,N_7098,N_9846);
nor U13362 (N_13362,N_7904,N_6596);
nand U13363 (N_13363,N_5294,N_8520);
or U13364 (N_13364,N_9050,N_6213);
nand U13365 (N_13365,N_8343,N_6694);
nor U13366 (N_13366,N_7035,N_6688);
nand U13367 (N_13367,N_8616,N_9819);
or U13368 (N_13368,N_8719,N_8570);
xor U13369 (N_13369,N_7009,N_9826);
or U13370 (N_13370,N_7239,N_8492);
and U13371 (N_13371,N_6829,N_6290);
or U13372 (N_13372,N_7597,N_8433);
or U13373 (N_13373,N_9208,N_7144);
and U13374 (N_13374,N_7880,N_8013);
and U13375 (N_13375,N_6160,N_7710);
nand U13376 (N_13376,N_8185,N_8450);
or U13377 (N_13377,N_6192,N_9027);
nor U13378 (N_13378,N_7761,N_8706);
or U13379 (N_13379,N_7121,N_6243);
and U13380 (N_13380,N_8547,N_9852);
nor U13381 (N_13381,N_6336,N_6485);
nand U13382 (N_13382,N_5341,N_9311);
or U13383 (N_13383,N_9244,N_9182);
nor U13384 (N_13384,N_6408,N_7439);
or U13385 (N_13385,N_5606,N_9117);
and U13386 (N_13386,N_6402,N_5740);
xor U13387 (N_13387,N_8789,N_7421);
and U13388 (N_13388,N_8129,N_7614);
nor U13389 (N_13389,N_8703,N_8038);
and U13390 (N_13390,N_5244,N_9282);
nand U13391 (N_13391,N_6445,N_7744);
and U13392 (N_13392,N_5986,N_6040);
and U13393 (N_13393,N_5333,N_8607);
or U13394 (N_13394,N_6405,N_7636);
or U13395 (N_13395,N_6045,N_7017);
nand U13396 (N_13396,N_8117,N_5593);
and U13397 (N_13397,N_9340,N_6992);
nor U13398 (N_13398,N_9159,N_7735);
nor U13399 (N_13399,N_9260,N_9989);
nand U13400 (N_13400,N_9592,N_6990);
nand U13401 (N_13401,N_6216,N_9442);
nand U13402 (N_13402,N_5648,N_6177);
and U13403 (N_13403,N_6229,N_6836);
or U13404 (N_13404,N_5035,N_8121);
or U13405 (N_13405,N_6014,N_7542);
nor U13406 (N_13406,N_6183,N_5005);
and U13407 (N_13407,N_7468,N_7581);
or U13408 (N_13408,N_6516,N_6585);
nand U13409 (N_13409,N_9362,N_9814);
nor U13410 (N_13410,N_9289,N_9510);
or U13411 (N_13411,N_8513,N_7673);
xor U13412 (N_13412,N_6306,N_6350);
nor U13413 (N_13413,N_7411,N_8084);
nand U13414 (N_13414,N_5679,N_6571);
nand U13415 (N_13415,N_6830,N_8454);
nor U13416 (N_13416,N_6141,N_6491);
nand U13417 (N_13417,N_8474,N_5278);
nand U13418 (N_13418,N_8980,N_8876);
nor U13419 (N_13419,N_7523,N_6961);
nand U13420 (N_13420,N_7438,N_6634);
nor U13421 (N_13421,N_9053,N_8327);
or U13422 (N_13422,N_9527,N_8346);
and U13423 (N_13423,N_5474,N_9394);
nor U13424 (N_13424,N_9113,N_7057);
nor U13425 (N_13425,N_6694,N_8028);
and U13426 (N_13426,N_7493,N_6619);
nor U13427 (N_13427,N_6179,N_5405);
nand U13428 (N_13428,N_7629,N_6514);
nor U13429 (N_13429,N_6343,N_9951);
xor U13430 (N_13430,N_8417,N_8210);
nor U13431 (N_13431,N_6465,N_8769);
or U13432 (N_13432,N_8978,N_8330);
and U13433 (N_13433,N_6444,N_9226);
nor U13434 (N_13434,N_7214,N_7577);
or U13435 (N_13435,N_9945,N_9663);
and U13436 (N_13436,N_8813,N_6912);
and U13437 (N_13437,N_7586,N_8166);
nor U13438 (N_13438,N_7888,N_5058);
and U13439 (N_13439,N_5006,N_9347);
and U13440 (N_13440,N_9939,N_5497);
nor U13441 (N_13441,N_7369,N_8709);
or U13442 (N_13442,N_6757,N_5213);
nand U13443 (N_13443,N_7284,N_5118);
nor U13444 (N_13444,N_6152,N_7234);
and U13445 (N_13445,N_9347,N_6711);
nor U13446 (N_13446,N_9227,N_8913);
or U13447 (N_13447,N_8644,N_7924);
or U13448 (N_13448,N_6503,N_5721);
or U13449 (N_13449,N_9998,N_5285);
and U13450 (N_13450,N_5494,N_7538);
and U13451 (N_13451,N_9163,N_5445);
xnor U13452 (N_13452,N_8771,N_7367);
xnor U13453 (N_13453,N_5820,N_6552);
nand U13454 (N_13454,N_8915,N_6819);
or U13455 (N_13455,N_7718,N_7595);
nor U13456 (N_13456,N_8237,N_9079);
and U13457 (N_13457,N_9459,N_8164);
nand U13458 (N_13458,N_8192,N_9792);
xnor U13459 (N_13459,N_7125,N_7923);
xnor U13460 (N_13460,N_5793,N_9512);
and U13461 (N_13461,N_8175,N_5616);
nand U13462 (N_13462,N_8375,N_6281);
nor U13463 (N_13463,N_8134,N_9664);
and U13464 (N_13464,N_9992,N_6078);
nand U13465 (N_13465,N_6707,N_9437);
nand U13466 (N_13466,N_5010,N_8060);
and U13467 (N_13467,N_8775,N_8130);
nand U13468 (N_13468,N_6153,N_7460);
xor U13469 (N_13469,N_8491,N_7592);
and U13470 (N_13470,N_7750,N_6283);
xnor U13471 (N_13471,N_7067,N_5433);
and U13472 (N_13472,N_7685,N_9196);
nor U13473 (N_13473,N_7647,N_9201);
xnor U13474 (N_13474,N_8160,N_6458);
nor U13475 (N_13475,N_5358,N_7187);
nand U13476 (N_13476,N_9558,N_7379);
and U13477 (N_13477,N_6708,N_7850);
xor U13478 (N_13478,N_6297,N_6436);
nand U13479 (N_13479,N_9339,N_7619);
or U13480 (N_13480,N_6329,N_5033);
nand U13481 (N_13481,N_8356,N_7223);
and U13482 (N_13482,N_9935,N_9128);
or U13483 (N_13483,N_5148,N_7130);
nor U13484 (N_13484,N_8301,N_8164);
and U13485 (N_13485,N_9312,N_6021);
or U13486 (N_13486,N_5002,N_9939);
and U13487 (N_13487,N_5230,N_7343);
and U13488 (N_13488,N_9570,N_5503);
or U13489 (N_13489,N_5420,N_7067);
nor U13490 (N_13490,N_6871,N_7987);
and U13491 (N_13491,N_9659,N_7378);
or U13492 (N_13492,N_8054,N_8544);
and U13493 (N_13493,N_8963,N_9394);
or U13494 (N_13494,N_7519,N_9170);
nand U13495 (N_13495,N_7731,N_6954);
or U13496 (N_13496,N_5544,N_7601);
xnor U13497 (N_13497,N_7435,N_9846);
or U13498 (N_13498,N_9244,N_7262);
nand U13499 (N_13499,N_5965,N_5147);
or U13500 (N_13500,N_6425,N_6230);
nand U13501 (N_13501,N_9763,N_8949);
xnor U13502 (N_13502,N_6297,N_7545);
nor U13503 (N_13503,N_5160,N_5078);
xor U13504 (N_13504,N_6234,N_8645);
xnor U13505 (N_13505,N_7362,N_8276);
and U13506 (N_13506,N_9838,N_8344);
nor U13507 (N_13507,N_8771,N_9731);
nand U13508 (N_13508,N_7353,N_8244);
or U13509 (N_13509,N_8123,N_6299);
xnor U13510 (N_13510,N_8107,N_6273);
and U13511 (N_13511,N_8919,N_5803);
and U13512 (N_13512,N_7316,N_8552);
nor U13513 (N_13513,N_8396,N_6281);
and U13514 (N_13514,N_6035,N_7230);
nor U13515 (N_13515,N_5921,N_8783);
and U13516 (N_13516,N_8399,N_7742);
or U13517 (N_13517,N_8962,N_8977);
nand U13518 (N_13518,N_9306,N_6631);
nor U13519 (N_13519,N_8054,N_6568);
and U13520 (N_13520,N_9703,N_5172);
xnor U13521 (N_13521,N_7883,N_5110);
and U13522 (N_13522,N_8579,N_6698);
nor U13523 (N_13523,N_6133,N_8883);
or U13524 (N_13524,N_5992,N_5667);
xnor U13525 (N_13525,N_6886,N_9026);
nand U13526 (N_13526,N_6395,N_8292);
or U13527 (N_13527,N_5623,N_9554);
nor U13528 (N_13528,N_7657,N_8419);
nor U13529 (N_13529,N_5324,N_5705);
nand U13530 (N_13530,N_7538,N_8432);
and U13531 (N_13531,N_7011,N_5264);
and U13532 (N_13532,N_8935,N_6390);
or U13533 (N_13533,N_8758,N_5532);
nand U13534 (N_13534,N_5624,N_6613);
and U13535 (N_13535,N_8953,N_5003);
nor U13536 (N_13536,N_6668,N_6056);
nand U13537 (N_13537,N_7848,N_9849);
and U13538 (N_13538,N_5760,N_5284);
nand U13539 (N_13539,N_9793,N_6195);
nand U13540 (N_13540,N_7529,N_9405);
or U13541 (N_13541,N_9098,N_7682);
or U13542 (N_13542,N_6521,N_6784);
or U13543 (N_13543,N_6232,N_9629);
or U13544 (N_13544,N_9371,N_5752);
nand U13545 (N_13545,N_9907,N_5164);
xor U13546 (N_13546,N_9977,N_6537);
nor U13547 (N_13547,N_7282,N_9128);
nand U13548 (N_13548,N_5458,N_9888);
and U13549 (N_13549,N_9585,N_8171);
nor U13550 (N_13550,N_6433,N_8748);
nor U13551 (N_13551,N_5738,N_5678);
or U13552 (N_13552,N_7777,N_7344);
xnor U13553 (N_13553,N_8307,N_6423);
or U13554 (N_13554,N_7618,N_8610);
and U13555 (N_13555,N_6118,N_5166);
xnor U13556 (N_13556,N_5233,N_8632);
nand U13557 (N_13557,N_6125,N_9146);
and U13558 (N_13558,N_6885,N_7037);
nor U13559 (N_13559,N_9892,N_7620);
nor U13560 (N_13560,N_5978,N_7837);
or U13561 (N_13561,N_8987,N_8648);
nand U13562 (N_13562,N_7198,N_5909);
nor U13563 (N_13563,N_8831,N_6746);
nand U13564 (N_13564,N_7058,N_5670);
nand U13565 (N_13565,N_6381,N_7708);
nand U13566 (N_13566,N_7930,N_9627);
or U13567 (N_13567,N_7991,N_6971);
and U13568 (N_13568,N_8032,N_9050);
and U13569 (N_13569,N_6604,N_6034);
or U13570 (N_13570,N_8737,N_7249);
nor U13571 (N_13571,N_8805,N_7620);
nand U13572 (N_13572,N_9625,N_6051);
nand U13573 (N_13573,N_6437,N_8040);
nand U13574 (N_13574,N_7908,N_8467);
nor U13575 (N_13575,N_9472,N_5059);
nor U13576 (N_13576,N_5792,N_8638);
nand U13577 (N_13577,N_9601,N_8042);
nor U13578 (N_13578,N_9095,N_9804);
or U13579 (N_13579,N_9961,N_6142);
xnor U13580 (N_13580,N_6527,N_5773);
xor U13581 (N_13581,N_6626,N_6089);
and U13582 (N_13582,N_8502,N_5852);
nor U13583 (N_13583,N_9322,N_9360);
or U13584 (N_13584,N_5762,N_6108);
or U13585 (N_13585,N_9683,N_9735);
xor U13586 (N_13586,N_6056,N_7438);
or U13587 (N_13587,N_8486,N_9715);
nand U13588 (N_13588,N_5735,N_8423);
or U13589 (N_13589,N_9381,N_5725);
xnor U13590 (N_13590,N_9337,N_8347);
nor U13591 (N_13591,N_7264,N_5298);
or U13592 (N_13592,N_5182,N_8477);
and U13593 (N_13593,N_5850,N_6699);
nand U13594 (N_13594,N_8183,N_6359);
and U13595 (N_13595,N_6809,N_7964);
or U13596 (N_13596,N_5675,N_5663);
or U13597 (N_13597,N_8350,N_9740);
nor U13598 (N_13598,N_8914,N_5173);
or U13599 (N_13599,N_5526,N_6176);
nand U13600 (N_13600,N_9405,N_5572);
or U13601 (N_13601,N_9869,N_7523);
xnor U13602 (N_13602,N_8475,N_6024);
and U13603 (N_13603,N_8858,N_7892);
or U13604 (N_13604,N_6186,N_6618);
nand U13605 (N_13605,N_9040,N_6098);
or U13606 (N_13606,N_6979,N_5218);
and U13607 (N_13607,N_5604,N_8955);
or U13608 (N_13608,N_9069,N_6661);
or U13609 (N_13609,N_9919,N_8605);
nand U13610 (N_13610,N_7324,N_7896);
nor U13611 (N_13611,N_8756,N_7079);
nor U13612 (N_13612,N_5804,N_7579);
or U13613 (N_13613,N_8605,N_7352);
nand U13614 (N_13614,N_7949,N_8104);
nor U13615 (N_13615,N_7242,N_8750);
nor U13616 (N_13616,N_9287,N_9065);
or U13617 (N_13617,N_5623,N_6952);
or U13618 (N_13618,N_5211,N_5162);
nand U13619 (N_13619,N_7682,N_7098);
or U13620 (N_13620,N_7259,N_5743);
nor U13621 (N_13621,N_5191,N_5590);
and U13622 (N_13622,N_7975,N_5541);
nor U13623 (N_13623,N_8212,N_8064);
xor U13624 (N_13624,N_5135,N_6946);
or U13625 (N_13625,N_6977,N_9016);
nor U13626 (N_13626,N_8147,N_6490);
xor U13627 (N_13627,N_8846,N_5126);
or U13628 (N_13628,N_7658,N_8297);
nand U13629 (N_13629,N_8404,N_7486);
nand U13630 (N_13630,N_5582,N_8357);
nand U13631 (N_13631,N_6369,N_8568);
nor U13632 (N_13632,N_5117,N_9082);
and U13633 (N_13633,N_9997,N_7760);
xor U13634 (N_13634,N_8553,N_6208);
nand U13635 (N_13635,N_5489,N_6454);
nand U13636 (N_13636,N_5906,N_7878);
nor U13637 (N_13637,N_5956,N_9582);
and U13638 (N_13638,N_9912,N_5684);
and U13639 (N_13639,N_9077,N_7558);
xnor U13640 (N_13640,N_5256,N_5372);
nor U13641 (N_13641,N_5116,N_6616);
and U13642 (N_13642,N_7902,N_5479);
and U13643 (N_13643,N_8206,N_8303);
and U13644 (N_13644,N_7489,N_8209);
nand U13645 (N_13645,N_8250,N_5196);
nand U13646 (N_13646,N_7696,N_7172);
nand U13647 (N_13647,N_6447,N_6242);
or U13648 (N_13648,N_8463,N_9059);
or U13649 (N_13649,N_8116,N_7995);
or U13650 (N_13650,N_5434,N_5343);
xor U13651 (N_13651,N_6036,N_6507);
and U13652 (N_13652,N_8818,N_9176);
nand U13653 (N_13653,N_9070,N_7885);
nor U13654 (N_13654,N_8733,N_9439);
nor U13655 (N_13655,N_6015,N_7577);
nor U13656 (N_13656,N_9062,N_7258);
nor U13657 (N_13657,N_8947,N_7886);
or U13658 (N_13658,N_6710,N_5898);
and U13659 (N_13659,N_8542,N_8338);
or U13660 (N_13660,N_5547,N_6982);
or U13661 (N_13661,N_8703,N_6836);
nor U13662 (N_13662,N_8854,N_5963);
or U13663 (N_13663,N_8691,N_6664);
xnor U13664 (N_13664,N_7910,N_5167);
xnor U13665 (N_13665,N_5546,N_7001);
nand U13666 (N_13666,N_7308,N_8658);
nor U13667 (N_13667,N_9057,N_5859);
or U13668 (N_13668,N_8307,N_8623);
nand U13669 (N_13669,N_9274,N_7407);
nand U13670 (N_13670,N_6639,N_7249);
and U13671 (N_13671,N_7519,N_8677);
and U13672 (N_13672,N_9325,N_9009);
nand U13673 (N_13673,N_5293,N_7343);
nand U13674 (N_13674,N_9097,N_9716);
or U13675 (N_13675,N_7809,N_7803);
nor U13676 (N_13676,N_6310,N_8197);
nor U13677 (N_13677,N_5663,N_6232);
and U13678 (N_13678,N_5646,N_9705);
or U13679 (N_13679,N_6124,N_7928);
and U13680 (N_13680,N_5528,N_8491);
nand U13681 (N_13681,N_7255,N_7632);
or U13682 (N_13682,N_5036,N_9895);
nor U13683 (N_13683,N_6710,N_8080);
or U13684 (N_13684,N_7089,N_5338);
nor U13685 (N_13685,N_8069,N_6579);
and U13686 (N_13686,N_6148,N_8476);
nand U13687 (N_13687,N_5581,N_6451);
nor U13688 (N_13688,N_6111,N_6602);
or U13689 (N_13689,N_9419,N_8920);
nand U13690 (N_13690,N_9713,N_7114);
xor U13691 (N_13691,N_9725,N_8115);
or U13692 (N_13692,N_6261,N_9954);
or U13693 (N_13693,N_7015,N_5105);
nor U13694 (N_13694,N_5533,N_5948);
nor U13695 (N_13695,N_6619,N_5437);
nand U13696 (N_13696,N_8521,N_6193);
nor U13697 (N_13697,N_9770,N_9928);
or U13698 (N_13698,N_7035,N_5663);
or U13699 (N_13699,N_6668,N_5712);
nand U13700 (N_13700,N_8925,N_5467);
and U13701 (N_13701,N_9299,N_8023);
and U13702 (N_13702,N_7294,N_6288);
and U13703 (N_13703,N_5164,N_9503);
and U13704 (N_13704,N_7142,N_5106);
xnor U13705 (N_13705,N_8581,N_9243);
xnor U13706 (N_13706,N_7408,N_8957);
nor U13707 (N_13707,N_9698,N_7200);
or U13708 (N_13708,N_7653,N_7623);
xor U13709 (N_13709,N_5734,N_7373);
or U13710 (N_13710,N_6879,N_7129);
and U13711 (N_13711,N_7837,N_7571);
or U13712 (N_13712,N_6535,N_8640);
nand U13713 (N_13713,N_8868,N_6870);
and U13714 (N_13714,N_8462,N_7877);
or U13715 (N_13715,N_8650,N_8309);
and U13716 (N_13716,N_8188,N_7301);
and U13717 (N_13717,N_8793,N_8743);
or U13718 (N_13718,N_9355,N_9534);
xnor U13719 (N_13719,N_5725,N_6376);
nor U13720 (N_13720,N_5143,N_7179);
nand U13721 (N_13721,N_6497,N_9469);
nand U13722 (N_13722,N_7160,N_5407);
and U13723 (N_13723,N_7227,N_9136);
nand U13724 (N_13724,N_6641,N_8304);
nor U13725 (N_13725,N_7219,N_5582);
and U13726 (N_13726,N_5799,N_5967);
nand U13727 (N_13727,N_6278,N_8229);
or U13728 (N_13728,N_7249,N_9457);
nor U13729 (N_13729,N_5425,N_6325);
and U13730 (N_13730,N_8786,N_7051);
nand U13731 (N_13731,N_5785,N_6304);
and U13732 (N_13732,N_7787,N_7668);
or U13733 (N_13733,N_9617,N_6370);
and U13734 (N_13734,N_5502,N_8715);
or U13735 (N_13735,N_6610,N_8702);
nor U13736 (N_13736,N_9241,N_6054);
or U13737 (N_13737,N_5698,N_9828);
nor U13738 (N_13738,N_9497,N_9310);
nor U13739 (N_13739,N_8096,N_5960);
nand U13740 (N_13740,N_8488,N_8425);
nand U13741 (N_13741,N_9156,N_5423);
or U13742 (N_13742,N_6064,N_5059);
nor U13743 (N_13743,N_8804,N_5578);
nor U13744 (N_13744,N_9019,N_5452);
nand U13745 (N_13745,N_9442,N_6692);
and U13746 (N_13746,N_5613,N_5651);
nand U13747 (N_13747,N_7112,N_9728);
or U13748 (N_13748,N_9082,N_9594);
nand U13749 (N_13749,N_7382,N_8480);
and U13750 (N_13750,N_8228,N_5099);
xnor U13751 (N_13751,N_5348,N_5600);
or U13752 (N_13752,N_5118,N_9905);
nor U13753 (N_13753,N_7207,N_9567);
or U13754 (N_13754,N_5251,N_6340);
nand U13755 (N_13755,N_6539,N_5827);
nand U13756 (N_13756,N_6141,N_7546);
xnor U13757 (N_13757,N_7814,N_9874);
nor U13758 (N_13758,N_7535,N_6085);
xor U13759 (N_13759,N_7928,N_7100);
or U13760 (N_13760,N_8863,N_7914);
and U13761 (N_13761,N_8253,N_6034);
nand U13762 (N_13762,N_7184,N_8991);
nor U13763 (N_13763,N_8448,N_7384);
nor U13764 (N_13764,N_5550,N_8124);
nor U13765 (N_13765,N_7259,N_7930);
or U13766 (N_13766,N_5441,N_7143);
and U13767 (N_13767,N_6266,N_7537);
and U13768 (N_13768,N_8530,N_6068);
or U13769 (N_13769,N_6188,N_9854);
and U13770 (N_13770,N_5092,N_5729);
nand U13771 (N_13771,N_8431,N_8184);
nor U13772 (N_13772,N_9426,N_8635);
nor U13773 (N_13773,N_5701,N_7355);
nor U13774 (N_13774,N_8439,N_9514);
xor U13775 (N_13775,N_5344,N_8770);
or U13776 (N_13776,N_6880,N_9728);
nor U13777 (N_13777,N_9572,N_6852);
nor U13778 (N_13778,N_8750,N_5833);
or U13779 (N_13779,N_8801,N_8632);
xnor U13780 (N_13780,N_5329,N_5183);
xnor U13781 (N_13781,N_8876,N_9094);
or U13782 (N_13782,N_5001,N_8042);
and U13783 (N_13783,N_7559,N_9306);
and U13784 (N_13784,N_9984,N_7970);
nand U13785 (N_13785,N_6932,N_9115);
nand U13786 (N_13786,N_5651,N_9922);
xnor U13787 (N_13787,N_7397,N_6612);
nor U13788 (N_13788,N_5025,N_9721);
or U13789 (N_13789,N_8836,N_8077);
nand U13790 (N_13790,N_6553,N_9302);
nor U13791 (N_13791,N_8739,N_9438);
nor U13792 (N_13792,N_6114,N_7068);
nand U13793 (N_13793,N_9633,N_6173);
nand U13794 (N_13794,N_9042,N_6041);
nor U13795 (N_13795,N_6376,N_6359);
and U13796 (N_13796,N_5925,N_5586);
and U13797 (N_13797,N_5606,N_6679);
nor U13798 (N_13798,N_9919,N_7689);
xor U13799 (N_13799,N_7681,N_5984);
nor U13800 (N_13800,N_9363,N_6167);
nand U13801 (N_13801,N_9509,N_6938);
or U13802 (N_13802,N_9686,N_8128);
and U13803 (N_13803,N_8542,N_6370);
nor U13804 (N_13804,N_6244,N_5714);
nor U13805 (N_13805,N_7090,N_7020);
or U13806 (N_13806,N_8386,N_8908);
and U13807 (N_13807,N_8005,N_6898);
nor U13808 (N_13808,N_8664,N_9533);
xor U13809 (N_13809,N_8170,N_9177);
or U13810 (N_13810,N_5092,N_7944);
nor U13811 (N_13811,N_9674,N_8410);
nor U13812 (N_13812,N_6532,N_9621);
or U13813 (N_13813,N_8767,N_5315);
and U13814 (N_13814,N_5186,N_9821);
nand U13815 (N_13815,N_9214,N_6917);
nand U13816 (N_13816,N_6624,N_5053);
and U13817 (N_13817,N_9180,N_5998);
xnor U13818 (N_13818,N_6156,N_9288);
and U13819 (N_13819,N_5445,N_6447);
or U13820 (N_13820,N_7325,N_8694);
or U13821 (N_13821,N_8591,N_5441);
nand U13822 (N_13822,N_8326,N_9975);
nand U13823 (N_13823,N_9536,N_8795);
and U13824 (N_13824,N_5182,N_9556);
nand U13825 (N_13825,N_5207,N_5756);
nand U13826 (N_13826,N_7032,N_6936);
nor U13827 (N_13827,N_7223,N_6644);
xnor U13828 (N_13828,N_5421,N_9622);
xor U13829 (N_13829,N_8538,N_9036);
or U13830 (N_13830,N_5348,N_9944);
nor U13831 (N_13831,N_6135,N_8254);
nor U13832 (N_13832,N_5191,N_7657);
nand U13833 (N_13833,N_9275,N_5214);
nand U13834 (N_13834,N_5637,N_8634);
or U13835 (N_13835,N_7442,N_7643);
nand U13836 (N_13836,N_6405,N_6709);
nand U13837 (N_13837,N_8266,N_8489);
nor U13838 (N_13838,N_8745,N_8221);
or U13839 (N_13839,N_9484,N_5370);
xnor U13840 (N_13840,N_7170,N_6906);
nand U13841 (N_13841,N_5809,N_8189);
and U13842 (N_13842,N_5304,N_6877);
nor U13843 (N_13843,N_9323,N_8552);
and U13844 (N_13844,N_6456,N_8327);
nor U13845 (N_13845,N_9749,N_9857);
nor U13846 (N_13846,N_9659,N_6843);
and U13847 (N_13847,N_6963,N_9795);
and U13848 (N_13848,N_5215,N_6588);
nor U13849 (N_13849,N_5668,N_5313);
or U13850 (N_13850,N_8757,N_9096);
or U13851 (N_13851,N_7446,N_8078);
and U13852 (N_13852,N_9446,N_6224);
and U13853 (N_13853,N_7820,N_6589);
or U13854 (N_13854,N_5488,N_8802);
or U13855 (N_13855,N_8898,N_8240);
nor U13856 (N_13856,N_5371,N_5424);
and U13857 (N_13857,N_5545,N_9060);
nand U13858 (N_13858,N_5658,N_6859);
nor U13859 (N_13859,N_9982,N_7468);
nor U13860 (N_13860,N_9085,N_5645);
or U13861 (N_13861,N_6962,N_8056);
or U13862 (N_13862,N_7954,N_8696);
and U13863 (N_13863,N_7414,N_6562);
and U13864 (N_13864,N_6291,N_8750);
nand U13865 (N_13865,N_8090,N_9441);
or U13866 (N_13866,N_5267,N_6186);
nand U13867 (N_13867,N_8535,N_5485);
and U13868 (N_13868,N_6676,N_5951);
nand U13869 (N_13869,N_9850,N_9512);
nand U13870 (N_13870,N_7514,N_7153);
nor U13871 (N_13871,N_9487,N_5463);
nor U13872 (N_13872,N_8613,N_6318);
and U13873 (N_13873,N_9070,N_8927);
and U13874 (N_13874,N_6784,N_8644);
or U13875 (N_13875,N_6039,N_6447);
nand U13876 (N_13876,N_5033,N_9465);
nor U13877 (N_13877,N_7103,N_7045);
and U13878 (N_13878,N_8819,N_5778);
nand U13879 (N_13879,N_8607,N_7688);
xor U13880 (N_13880,N_9320,N_7814);
or U13881 (N_13881,N_5291,N_5568);
nand U13882 (N_13882,N_9693,N_5442);
and U13883 (N_13883,N_6170,N_8227);
nor U13884 (N_13884,N_7418,N_9347);
nor U13885 (N_13885,N_9967,N_9757);
nor U13886 (N_13886,N_9576,N_8221);
or U13887 (N_13887,N_7064,N_6076);
and U13888 (N_13888,N_7685,N_5129);
or U13889 (N_13889,N_5984,N_5492);
nor U13890 (N_13890,N_8841,N_6419);
or U13891 (N_13891,N_7061,N_6250);
or U13892 (N_13892,N_8500,N_6811);
xnor U13893 (N_13893,N_6364,N_8315);
or U13894 (N_13894,N_7876,N_5350);
nor U13895 (N_13895,N_9128,N_6198);
nor U13896 (N_13896,N_6304,N_9812);
nor U13897 (N_13897,N_5189,N_7166);
nand U13898 (N_13898,N_8123,N_9446);
nand U13899 (N_13899,N_7834,N_8222);
xnor U13900 (N_13900,N_6624,N_8653);
nand U13901 (N_13901,N_6510,N_9657);
and U13902 (N_13902,N_9119,N_7827);
or U13903 (N_13903,N_7958,N_6090);
and U13904 (N_13904,N_5422,N_5537);
nand U13905 (N_13905,N_7805,N_7053);
or U13906 (N_13906,N_8721,N_8560);
xor U13907 (N_13907,N_7523,N_8209);
nor U13908 (N_13908,N_7298,N_9000);
nand U13909 (N_13909,N_8508,N_6194);
nor U13910 (N_13910,N_7801,N_7238);
and U13911 (N_13911,N_9284,N_9985);
and U13912 (N_13912,N_9731,N_8322);
or U13913 (N_13913,N_6769,N_5505);
or U13914 (N_13914,N_9761,N_5570);
xnor U13915 (N_13915,N_7848,N_9709);
nand U13916 (N_13916,N_6094,N_9713);
nand U13917 (N_13917,N_9287,N_7083);
nor U13918 (N_13918,N_6869,N_8903);
nor U13919 (N_13919,N_7439,N_5808);
or U13920 (N_13920,N_9360,N_7654);
or U13921 (N_13921,N_8902,N_7618);
nor U13922 (N_13922,N_7907,N_7236);
xor U13923 (N_13923,N_6870,N_5100);
xnor U13924 (N_13924,N_8697,N_8217);
nor U13925 (N_13925,N_9405,N_6057);
nand U13926 (N_13926,N_5732,N_7379);
xnor U13927 (N_13927,N_7202,N_9976);
nor U13928 (N_13928,N_8248,N_7315);
nand U13929 (N_13929,N_6494,N_8100);
nor U13930 (N_13930,N_8643,N_5442);
nor U13931 (N_13931,N_9047,N_6731);
nor U13932 (N_13932,N_9309,N_6327);
nand U13933 (N_13933,N_5819,N_6817);
xor U13934 (N_13934,N_5089,N_5001);
nor U13935 (N_13935,N_6521,N_6991);
and U13936 (N_13936,N_8910,N_7720);
and U13937 (N_13937,N_9932,N_5869);
and U13938 (N_13938,N_8118,N_9294);
or U13939 (N_13939,N_6981,N_9771);
nand U13940 (N_13940,N_6305,N_9143);
nand U13941 (N_13941,N_6714,N_8766);
nand U13942 (N_13942,N_7004,N_5083);
and U13943 (N_13943,N_8823,N_5690);
nor U13944 (N_13944,N_7866,N_8469);
and U13945 (N_13945,N_6614,N_6513);
nor U13946 (N_13946,N_7226,N_5644);
nor U13947 (N_13947,N_9046,N_8790);
nand U13948 (N_13948,N_9156,N_5556);
xnor U13949 (N_13949,N_9526,N_5290);
nor U13950 (N_13950,N_5668,N_9217);
nand U13951 (N_13951,N_8139,N_9400);
nand U13952 (N_13952,N_7040,N_7490);
and U13953 (N_13953,N_8653,N_7390);
nor U13954 (N_13954,N_8928,N_6543);
nand U13955 (N_13955,N_5593,N_5564);
nor U13956 (N_13956,N_6115,N_5464);
or U13957 (N_13957,N_7212,N_8796);
nand U13958 (N_13958,N_8919,N_5502);
nor U13959 (N_13959,N_5781,N_7439);
nand U13960 (N_13960,N_8913,N_7154);
nand U13961 (N_13961,N_9960,N_6712);
and U13962 (N_13962,N_5046,N_6900);
nor U13963 (N_13963,N_9407,N_6620);
and U13964 (N_13964,N_6857,N_6505);
xnor U13965 (N_13965,N_7590,N_7996);
and U13966 (N_13966,N_9855,N_8337);
nor U13967 (N_13967,N_5013,N_5892);
nor U13968 (N_13968,N_7047,N_8295);
and U13969 (N_13969,N_8068,N_8477);
xnor U13970 (N_13970,N_5960,N_6194);
or U13971 (N_13971,N_7515,N_6120);
and U13972 (N_13972,N_9316,N_6713);
and U13973 (N_13973,N_8756,N_8915);
xnor U13974 (N_13974,N_6448,N_8779);
nor U13975 (N_13975,N_7619,N_8904);
or U13976 (N_13976,N_8307,N_8264);
xnor U13977 (N_13977,N_8123,N_5322);
nand U13978 (N_13978,N_6039,N_5507);
and U13979 (N_13979,N_9725,N_7514);
nor U13980 (N_13980,N_6747,N_5031);
or U13981 (N_13981,N_8940,N_9585);
nand U13982 (N_13982,N_8206,N_9247);
or U13983 (N_13983,N_9260,N_5726);
nor U13984 (N_13984,N_8402,N_6328);
nand U13985 (N_13985,N_6972,N_5336);
nor U13986 (N_13986,N_8984,N_7414);
or U13987 (N_13987,N_5699,N_8486);
nor U13988 (N_13988,N_8441,N_8986);
xnor U13989 (N_13989,N_9232,N_8302);
xor U13990 (N_13990,N_8926,N_5715);
or U13991 (N_13991,N_7365,N_8510);
nand U13992 (N_13992,N_9232,N_9784);
or U13993 (N_13993,N_7867,N_9592);
and U13994 (N_13994,N_8329,N_7085);
nand U13995 (N_13995,N_7005,N_5395);
or U13996 (N_13996,N_6410,N_9939);
nor U13997 (N_13997,N_5941,N_5626);
and U13998 (N_13998,N_5471,N_6234);
or U13999 (N_13999,N_5510,N_7434);
nand U14000 (N_14000,N_9644,N_7112);
or U14001 (N_14001,N_9589,N_9830);
nor U14002 (N_14002,N_7718,N_8514);
xor U14003 (N_14003,N_8586,N_7748);
nor U14004 (N_14004,N_8116,N_8347);
nor U14005 (N_14005,N_8816,N_5460);
nor U14006 (N_14006,N_6036,N_6688);
or U14007 (N_14007,N_6987,N_8559);
nor U14008 (N_14008,N_6556,N_9813);
nand U14009 (N_14009,N_5852,N_9571);
nand U14010 (N_14010,N_6533,N_5528);
nor U14011 (N_14011,N_6551,N_7645);
xor U14012 (N_14012,N_9431,N_7964);
or U14013 (N_14013,N_8279,N_7885);
and U14014 (N_14014,N_5607,N_8565);
xnor U14015 (N_14015,N_6293,N_9282);
nand U14016 (N_14016,N_7024,N_8285);
nand U14017 (N_14017,N_7752,N_5171);
and U14018 (N_14018,N_6163,N_7658);
or U14019 (N_14019,N_8369,N_9204);
and U14020 (N_14020,N_8886,N_8320);
nor U14021 (N_14021,N_5284,N_6197);
nor U14022 (N_14022,N_6397,N_8739);
and U14023 (N_14023,N_5068,N_6039);
xnor U14024 (N_14024,N_9361,N_7425);
nand U14025 (N_14025,N_9260,N_7782);
and U14026 (N_14026,N_9080,N_5217);
and U14027 (N_14027,N_6187,N_7320);
or U14028 (N_14028,N_8466,N_9641);
xor U14029 (N_14029,N_6214,N_9173);
nand U14030 (N_14030,N_6267,N_7324);
nand U14031 (N_14031,N_7373,N_9928);
and U14032 (N_14032,N_8762,N_8510);
or U14033 (N_14033,N_5522,N_6131);
and U14034 (N_14034,N_7451,N_6639);
and U14035 (N_14035,N_6264,N_7621);
and U14036 (N_14036,N_7872,N_6057);
nand U14037 (N_14037,N_5617,N_7918);
or U14038 (N_14038,N_7701,N_5925);
or U14039 (N_14039,N_5513,N_8174);
nand U14040 (N_14040,N_9552,N_9788);
nand U14041 (N_14041,N_8948,N_6731);
xor U14042 (N_14042,N_7056,N_5604);
and U14043 (N_14043,N_7699,N_7848);
or U14044 (N_14044,N_6636,N_6858);
or U14045 (N_14045,N_8708,N_5560);
and U14046 (N_14046,N_9449,N_5354);
xnor U14047 (N_14047,N_8235,N_8079);
or U14048 (N_14048,N_9812,N_8390);
and U14049 (N_14049,N_7873,N_6858);
xor U14050 (N_14050,N_8081,N_7487);
and U14051 (N_14051,N_7232,N_9699);
nor U14052 (N_14052,N_8624,N_7193);
and U14053 (N_14053,N_6346,N_7448);
or U14054 (N_14054,N_5521,N_6912);
and U14055 (N_14055,N_5500,N_7842);
and U14056 (N_14056,N_5240,N_7228);
or U14057 (N_14057,N_6879,N_5526);
nand U14058 (N_14058,N_9098,N_9673);
nand U14059 (N_14059,N_7756,N_8725);
or U14060 (N_14060,N_6905,N_8229);
xor U14061 (N_14061,N_5230,N_8173);
nand U14062 (N_14062,N_5878,N_7285);
nor U14063 (N_14063,N_6316,N_9377);
or U14064 (N_14064,N_6037,N_8439);
nor U14065 (N_14065,N_9160,N_8159);
or U14066 (N_14066,N_6024,N_8967);
or U14067 (N_14067,N_7182,N_7773);
xor U14068 (N_14068,N_6313,N_8851);
and U14069 (N_14069,N_9259,N_6612);
nor U14070 (N_14070,N_7560,N_5273);
nand U14071 (N_14071,N_5624,N_8263);
nor U14072 (N_14072,N_8232,N_5940);
nor U14073 (N_14073,N_8274,N_7285);
nor U14074 (N_14074,N_5927,N_6307);
nand U14075 (N_14075,N_6674,N_8689);
nand U14076 (N_14076,N_9982,N_6055);
or U14077 (N_14077,N_7606,N_5125);
or U14078 (N_14078,N_7912,N_7743);
nor U14079 (N_14079,N_9779,N_6398);
and U14080 (N_14080,N_9700,N_6369);
and U14081 (N_14081,N_6132,N_9470);
nor U14082 (N_14082,N_9690,N_6158);
nand U14083 (N_14083,N_7483,N_8611);
nand U14084 (N_14084,N_7565,N_6373);
and U14085 (N_14085,N_8730,N_6188);
or U14086 (N_14086,N_6350,N_9017);
and U14087 (N_14087,N_6274,N_5304);
nor U14088 (N_14088,N_5497,N_7648);
and U14089 (N_14089,N_7515,N_9967);
nand U14090 (N_14090,N_9172,N_8365);
or U14091 (N_14091,N_9121,N_6533);
or U14092 (N_14092,N_7247,N_6002);
and U14093 (N_14093,N_5482,N_5320);
or U14094 (N_14094,N_9264,N_7555);
xnor U14095 (N_14095,N_8854,N_8551);
or U14096 (N_14096,N_7687,N_7701);
and U14097 (N_14097,N_9361,N_5906);
and U14098 (N_14098,N_7375,N_7021);
or U14099 (N_14099,N_8621,N_8846);
and U14100 (N_14100,N_7076,N_5666);
nand U14101 (N_14101,N_6232,N_7536);
nor U14102 (N_14102,N_7925,N_6964);
nand U14103 (N_14103,N_6160,N_7119);
or U14104 (N_14104,N_5059,N_8677);
nor U14105 (N_14105,N_6124,N_8814);
nor U14106 (N_14106,N_8271,N_5894);
or U14107 (N_14107,N_5703,N_6073);
nand U14108 (N_14108,N_8255,N_5077);
nand U14109 (N_14109,N_9847,N_5082);
or U14110 (N_14110,N_5190,N_5183);
nand U14111 (N_14111,N_7952,N_9351);
nand U14112 (N_14112,N_8956,N_5790);
or U14113 (N_14113,N_7115,N_9843);
nor U14114 (N_14114,N_8449,N_8418);
and U14115 (N_14115,N_8422,N_8766);
xor U14116 (N_14116,N_7210,N_5050);
and U14117 (N_14117,N_8923,N_5345);
xor U14118 (N_14118,N_6830,N_7044);
nand U14119 (N_14119,N_8489,N_5286);
and U14120 (N_14120,N_5035,N_8597);
nor U14121 (N_14121,N_7769,N_7954);
or U14122 (N_14122,N_8835,N_5779);
and U14123 (N_14123,N_7736,N_7991);
xor U14124 (N_14124,N_6753,N_7037);
nor U14125 (N_14125,N_6796,N_7527);
or U14126 (N_14126,N_5540,N_7792);
or U14127 (N_14127,N_5713,N_9757);
or U14128 (N_14128,N_7322,N_6155);
and U14129 (N_14129,N_7071,N_7323);
nor U14130 (N_14130,N_8755,N_7836);
nand U14131 (N_14131,N_7252,N_5299);
or U14132 (N_14132,N_5522,N_7783);
and U14133 (N_14133,N_9410,N_9788);
and U14134 (N_14134,N_7814,N_6739);
and U14135 (N_14135,N_5938,N_5649);
nor U14136 (N_14136,N_7265,N_8472);
or U14137 (N_14137,N_5632,N_6878);
nor U14138 (N_14138,N_5161,N_6370);
and U14139 (N_14139,N_8342,N_7314);
nor U14140 (N_14140,N_9980,N_7915);
and U14141 (N_14141,N_7115,N_8672);
and U14142 (N_14142,N_7347,N_9720);
nor U14143 (N_14143,N_9596,N_6001);
and U14144 (N_14144,N_5243,N_8110);
and U14145 (N_14145,N_9756,N_5468);
nor U14146 (N_14146,N_9991,N_6858);
nor U14147 (N_14147,N_9434,N_9991);
or U14148 (N_14148,N_6374,N_5887);
and U14149 (N_14149,N_6414,N_9039);
nand U14150 (N_14150,N_6305,N_9757);
or U14151 (N_14151,N_8211,N_8968);
nor U14152 (N_14152,N_8436,N_9727);
and U14153 (N_14153,N_6792,N_5251);
nand U14154 (N_14154,N_8543,N_8625);
and U14155 (N_14155,N_5914,N_8830);
or U14156 (N_14156,N_8076,N_9821);
nand U14157 (N_14157,N_6742,N_5648);
or U14158 (N_14158,N_9200,N_9547);
nand U14159 (N_14159,N_9744,N_9579);
or U14160 (N_14160,N_7099,N_9048);
nand U14161 (N_14161,N_9448,N_7618);
nand U14162 (N_14162,N_5250,N_8195);
nor U14163 (N_14163,N_9576,N_9783);
nor U14164 (N_14164,N_8883,N_6881);
nor U14165 (N_14165,N_9025,N_6718);
and U14166 (N_14166,N_9654,N_7407);
nor U14167 (N_14167,N_6329,N_6953);
or U14168 (N_14168,N_7942,N_9393);
or U14169 (N_14169,N_5619,N_7420);
nor U14170 (N_14170,N_6455,N_5733);
and U14171 (N_14171,N_8049,N_7449);
nor U14172 (N_14172,N_7190,N_7419);
nor U14173 (N_14173,N_9612,N_6420);
xor U14174 (N_14174,N_5196,N_9516);
or U14175 (N_14175,N_9245,N_6837);
nor U14176 (N_14176,N_5270,N_9938);
or U14177 (N_14177,N_7566,N_6428);
nand U14178 (N_14178,N_6690,N_6318);
nand U14179 (N_14179,N_7915,N_8903);
nor U14180 (N_14180,N_6852,N_6738);
or U14181 (N_14181,N_9776,N_5090);
nor U14182 (N_14182,N_6249,N_8983);
and U14183 (N_14183,N_8060,N_8454);
and U14184 (N_14184,N_8213,N_9648);
and U14185 (N_14185,N_9561,N_7987);
and U14186 (N_14186,N_5811,N_5479);
or U14187 (N_14187,N_8875,N_6688);
nor U14188 (N_14188,N_7047,N_6121);
nor U14189 (N_14189,N_6237,N_7064);
xnor U14190 (N_14190,N_7891,N_8322);
and U14191 (N_14191,N_9216,N_5721);
and U14192 (N_14192,N_8016,N_7710);
nor U14193 (N_14193,N_6998,N_6517);
and U14194 (N_14194,N_9900,N_6701);
nand U14195 (N_14195,N_7805,N_8989);
nand U14196 (N_14196,N_8684,N_5715);
and U14197 (N_14197,N_9946,N_9437);
nor U14198 (N_14198,N_5844,N_5126);
or U14199 (N_14199,N_6278,N_6740);
and U14200 (N_14200,N_5798,N_5198);
nand U14201 (N_14201,N_7571,N_9247);
and U14202 (N_14202,N_9215,N_9113);
or U14203 (N_14203,N_6020,N_9078);
nor U14204 (N_14204,N_8823,N_9436);
or U14205 (N_14205,N_9482,N_6801);
xor U14206 (N_14206,N_7512,N_8357);
nand U14207 (N_14207,N_5473,N_8319);
and U14208 (N_14208,N_6795,N_9501);
nand U14209 (N_14209,N_6241,N_5492);
nand U14210 (N_14210,N_5411,N_8965);
and U14211 (N_14211,N_9460,N_7589);
and U14212 (N_14212,N_6947,N_9592);
and U14213 (N_14213,N_8018,N_9692);
nor U14214 (N_14214,N_7467,N_8744);
nand U14215 (N_14215,N_5384,N_6272);
and U14216 (N_14216,N_9030,N_9888);
nor U14217 (N_14217,N_8554,N_7960);
and U14218 (N_14218,N_9202,N_5230);
nor U14219 (N_14219,N_9395,N_6182);
xor U14220 (N_14220,N_9130,N_6465);
xnor U14221 (N_14221,N_9598,N_6865);
nand U14222 (N_14222,N_8562,N_6022);
and U14223 (N_14223,N_7367,N_6045);
nor U14224 (N_14224,N_6466,N_8629);
and U14225 (N_14225,N_7786,N_8125);
xor U14226 (N_14226,N_5063,N_9577);
nor U14227 (N_14227,N_9056,N_9944);
or U14228 (N_14228,N_7152,N_7863);
or U14229 (N_14229,N_9333,N_8736);
or U14230 (N_14230,N_6108,N_9681);
and U14231 (N_14231,N_7401,N_7603);
nor U14232 (N_14232,N_6459,N_6333);
and U14233 (N_14233,N_8090,N_7364);
or U14234 (N_14234,N_6568,N_9168);
and U14235 (N_14235,N_7238,N_6524);
or U14236 (N_14236,N_7655,N_6982);
nand U14237 (N_14237,N_6104,N_7313);
and U14238 (N_14238,N_7833,N_9007);
and U14239 (N_14239,N_9769,N_9549);
xnor U14240 (N_14240,N_5641,N_5594);
or U14241 (N_14241,N_9616,N_6157);
nor U14242 (N_14242,N_9295,N_7080);
nor U14243 (N_14243,N_7318,N_7174);
nand U14244 (N_14244,N_5894,N_5745);
nand U14245 (N_14245,N_5327,N_9050);
nor U14246 (N_14246,N_6726,N_9644);
or U14247 (N_14247,N_8026,N_9499);
and U14248 (N_14248,N_9355,N_5567);
nand U14249 (N_14249,N_8553,N_6650);
or U14250 (N_14250,N_5615,N_6543);
nand U14251 (N_14251,N_6670,N_8175);
nor U14252 (N_14252,N_7165,N_8046);
nor U14253 (N_14253,N_8656,N_5072);
and U14254 (N_14254,N_6478,N_6944);
or U14255 (N_14255,N_6575,N_8427);
and U14256 (N_14256,N_7957,N_6890);
and U14257 (N_14257,N_9170,N_9346);
or U14258 (N_14258,N_8458,N_8292);
and U14259 (N_14259,N_5987,N_5647);
nand U14260 (N_14260,N_7506,N_5739);
and U14261 (N_14261,N_9369,N_5328);
and U14262 (N_14262,N_9994,N_8165);
or U14263 (N_14263,N_6062,N_9958);
or U14264 (N_14264,N_5412,N_6798);
and U14265 (N_14265,N_7568,N_9274);
or U14266 (N_14266,N_6328,N_8265);
or U14267 (N_14267,N_5811,N_6919);
and U14268 (N_14268,N_5336,N_7227);
nand U14269 (N_14269,N_8330,N_8025);
nand U14270 (N_14270,N_8356,N_9988);
and U14271 (N_14271,N_7399,N_6346);
and U14272 (N_14272,N_6395,N_9976);
and U14273 (N_14273,N_8755,N_7082);
and U14274 (N_14274,N_9390,N_6115);
xnor U14275 (N_14275,N_6264,N_9761);
or U14276 (N_14276,N_5411,N_6300);
xor U14277 (N_14277,N_5601,N_9211);
xor U14278 (N_14278,N_5087,N_5965);
nor U14279 (N_14279,N_6498,N_7578);
nand U14280 (N_14280,N_6103,N_7215);
nor U14281 (N_14281,N_6274,N_6684);
nor U14282 (N_14282,N_5432,N_9638);
and U14283 (N_14283,N_7179,N_8544);
nor U14284 (N_14284,N_9539,N_7118);
and U14285 (N_14285,N_9256,N_5492);
nand U14286 (N_14286,N_6316,N_7493);
and U14287 (N_14287,N_9722,N_9857);
nand U14288 (N_14288,N_7574,N_9191);
and U14289 (N_14289,N_5606,N_8244);
or U14290 (N_14290,N_8994,N_7491);
nand U14291 (N_14291,N_5222,N_9941);
nand U14292 (N_14292,N_9333,N_8385);
nor U14293 (N_14293,N_5044,N_6591);
or U14294 (N_14294,N_5828,N_6550);
nor U14295 (N_14295,N_8712,N_7937);
nor U14296 (N_14296,N_5988,N_7331);
or U14297 (N_14297,N_9223,N_5025);
and U14298 (N_14298,N_7967,N_7630);
xnor U14299 (N_14299,N_7068,N_9754);
or U14300 (N_14300,N_5412,N_5570);
and U14301 (N_14301,N_8063,N_8637);
or U14302 (N_14302,N_5329,N_9902);
and U14303 (N_14303,N_9491,N_8594);
or U14304 (N_14304,N_8003,N_9906);
or U14305 (N_14305,N_6377,N_8136);
and U14306 (N_14306,N_6386,N_9621);
or U14307 (N_14307,N_6918,N_5926);
nand U14308 (N_14308,N_8061,N_5725);
or U14309 (N_14309,N_7418,N_9442);
or U14310 (N_14310,N_8244,N_8243);
xor U14311 (N_14311,N_7285,N_8493);
or U14312 (N_14312,N_7450,N_9645);
nand U14313 (N_14313,N_7292,N_5136);
xnor U14314 (N_14314,N_6304,N_8822);
and U14315 (N_14315,N_5386,N_7151);
nand U14316 (N_14316,N_6939,N_6924);
nor U14317 (N_14317,N_9763,N_7108);
nor U14318 (N_14318,N_9721,N_6002);
nor U14319 (N_14319,N_6157,N_6456);
nand U14320 (N_14320,N_9178,N_6008);
or U14321 (N_14321,N_8648,N_6311);
and U14322 (N_14322,N_6998,N_5306);
or U14323 (N_14323,N_6950,N_8287);
nand U14324 (N_14324,N_6009,N_9068);
xnor U14325 (N_14325,N_8815,N_7909);
nor U14326 (N_14326,N_6062,N_7819);
or U14327 (N_14327,N_5506,N_7751);
nand U14328 (N_14328,N_8544,N_8326);
and U14329 (N_14329,N_8459,N_7365);
nand U14330 (N_14330,N_9486,N_7401);
nand U14331 (N_14331,N_6209,N_5762);
nand U14332 (N_14332,N_6736,N_7111);
nor U14333 (N_14333,N_9775,N_6539);
nor U14334 (N_14334,N_8482,N_6874);
nand U14335 (N_14335,N_6612,N_6866);
or U14336 (N_14336,N_6734,N_5135);
nand U14337 (N_14337,N_6291,N_7598);
and U14338 (N_14338,N_9625,N_9480);
nand U14339 (N_14339,N_9227,N_6719);
nand U14340 (N_14340,N_9828,N_9802);
nor U14341 (N_14341,N_8714,N_9455);
and U14342 (N_14342,N_5182,N_9924);
nand U14343 (N_14343,N_5717,N_8449);
nor U14344 (N_14344,N_5746,N_9968);
xor U14345 (N_14345,N_8848,N_5905);
or U14346 (N_14346,N_8762,N_8336);
xor U14347 (N_14347,N_5672,N_5252);
nand U14348 (N_14348,N_5268,N_8788);
or U14349 (N_14349,N_9778,N_8289);
nor U14350 (N_14350,N_8868,N_9434);
or U14351 (N_14351,N_8564,N_6870);
or U14352 (N_14352,N_7445,N_5812);
nor U14353 (N_14353,N_9451,N_5588);
xnor U14354 (N_14354,N_6256,N_5705);
and U14355 (N_14355,N_6088,N_8520);
nand U14356 (N_14356,N_5782,N_6090);
nand U14357 (N_14357,N_6694,N_8018);
or U14358 (N_14358,N_8277,N_6575);
nand U14359 (N_14359,N_8372,N_7162);
xnor U14360 (N_14360,N_5543,N_8859);
nand U14361 (N_14361,N_9069,N_6169);
or U14362 (N_14362,N_8249,N_8459);
or U14363 (N_14363,N_7341,N_8304);
xor U14364 (N_14364,N_8752,N_9301);
nor U14365 (N_14365,N_5581,N_9547);
and U14366 (N_14366,N_7168,N_9476);
nor U14367 (N_14367,N_9070,N_5065);
nand U14368 (N_14368,N_6706,N_7557);
nor U14369 (N_14369,N_5746,N_8663);
or U14370 (N_14370,N_5430,N_9944);
or U14371 (N_14371,N_9501,N_8197);
xor U14372 (N_14372,N_7986,N_8445);
nor U14373 (N_14373,N_8901,N_7179);
xnor U14374 (N_14374,N_5673,N_5452);
xnor U14375 (N_14375,N_6268,N_7997);
nand U14376 (N_14376,N_5622,N_6906);
nand U14377 (N_14377,N_5936,N_9004);
nor U14378 (N_14378,N_7561,N_6441);
and U14379 (N_14379,N_8578,N_6081);
xor U14380 (N_14380,N_9177,N_8527);
nor U14381 (N_14381,N_5075,N_7075);
nor U14382 (N_14382,N_9766,N_6057);
and U14383 (N_14383,N_6707,N_9016);
or U14384 (N_14384,N_8196,N_8762);
and U14385 (N_14385,N_6463,N_7298);
or U14386 (N_14386,N_7548,N_6393);
or U14387 (N_14387,N_5932,N_6793);
xor U14388 (N_14388,N_8651,N_9443);
xnor U14389 (N_14389,N_9902,N_7048);
nand U14390 (N_14390,N_7876,N_5904);
or U14391 (N_14391,N_6074,N_7446);
or U14392 (N_14392,N_8527,N_8828);
and U14393 (N_14393,N_7647,N_7260);
nand U14394 (N_14394,N_9529,N_6084);
and U14395 (N_14395,N_6928,N_8280);
or U14396 (N_14396,N_8637,N_9928);
or U14397 (N_14397,N_8237,N_7968);
nand U14398 (N_14398,N_8860,N_5819);
and U14399 (N_14399,N_5101,N_9090);
and U14400 (N_14400,N_9431,N_8262);
and U14401 (N_14401,N_7920,N_8956);
or U14402 (N_14402,N_7640,N_9125);
and U14403 (N_14403,N_9059,N_5765);
nand U14404 (N_14404,N_5265,N_7408);
or U14405 (N_14405,N_8829,N_6389);
nand U14406 (N_14406,N_8000,N_8856);
or U14407 (N_14407,N_8338,N_9460);
and U14408 (N_14408,N_9512,N_5135);
nand U14409 (N_14409,N_6658,N_9294);
xnor U14410 (N_14410,N_5374,N_8947);
or U14411 (N_14411,N_7993,N_7670);
nor U14412 (N_14412,N_5229,N_9298);
or U14413 (N_14413,N_8393,N_9375);
or U14414 (N_14414,N_7848,N_7200);
nand U14415 (N_14415,N_7290,N_7249);
nand U14416 (N_14416,N_9131,N_7060);
xor U14417 (N_14417,N_9698,N_5225);
nand U14418 (N_14418,N_9293,N_6775);
and U14419 (N_14419,N_8642,N_6424);
xor U14420 (N_14420,N_6140,N_7503);
and U14421 (N_14421,N_8791,N_6045);
xor U14422 (N_14422,N_5138,N_8713);
or U14423 (N_14423,N_8908,N_9336);
and U14424 (N_14424,N_6668,N_6868);
nand U14425 (N_14425,N_6477,N_5679);
nand U14426 (N_14426,N_7054,N_5545);
nor U14427 (N_14427,N_9190,N_5993);
nand U14428 (N_14428,N_8655,N_8818);
nor U14429 (N_14429,N_6618,N_6046);
nor U14430 (N_14430,N_5420,N_6670);
or U14431 (N_14431,N_8332,N_6886);
nand U14432 (N_14432,N_9226,N_8382);
nand U14433 (N_14433,N_7142,N_5026);
or U14434 (N_14434,N_8260,N_7703);
or U14435 (N_14435,N_5473,N_9153);
or U14436 (N_14436,N_8720,N_5104);
and U14437 (N_14437,N_7068,N_9839);
or U14438 (N_14438,N_8031,N_9898);
or U14439 (N_14439,N_5339,N_6240);
xor U14440 (N_14440,N_9899,N_6748);
nand U14441 (N_14441,N_7813,N_9876);
nor U14442 (N_14442,N_9690,N_6118);
or U14443 (N_14443,N_5342,N_5419);
nor U14444 (N_14444,N_7956,N_5070);
xor U14445 (N_14445,N_9262,N_9336);
nand U14446 (N_14446,N_7571,N_6613);
and U14447 (N_14447,N_5985,N_8064);
nand U14448 (N_14448,N_9415,N_9722);
and U14449 (N_14449,N_5640,N_5239);
or U14450 (N_14450,N_6019,N_8129);
and U14451 (N_14451,N_6587,N_8124);
or U14452 (N_14452,N_5863,N_8996);
xnor U14453 (N_14453,N_5408,N_7743);
and U14454 (N_14454,N_7483,N_8147);
and U14455 (N_14455,N_8342,N_8337);
nand U14456 (N_14456,N_6303,N_5279);
and U14457 (N_14457,N_9214,N_5440);
nand U14458 (N_14458,N_7011,N_6193);
nor U14459 (N_14459,N_6523,N_5678);
xnor U14460 (N_14460,N_5859,N_7447);
or U14461 (N_14461,N_8111,N_7914);
nor U14462 (N_14462,N_8578,N_8631);
or U14463 (N_14463,N_9796,N_8723);
nand U14464 (N_14464,N_8574,N_7071);
nor U14465 (N_14465,N_8984,N_9821);
or U14466 (N_14466,N_6575,N_5103);
or U14467 (N_14467,N_7813,N_8381);
nand U14468 (N_14468,N_9894,N_6955);
and U14469 (N_14469,N_6233,N_8251);
nand U14470 (N_14470,N_7633,N_8992);
or U14471 (N_14471,N_7215,N_8283);
nand U14472 (N_14472,N_6559,N_7852);
and U14473 (N_14473,N_7619,N_9343);
or U14474 (N_14474,N_6197,N_9255);
nand U14475 (N_14475,N_8412,N_6132);
and U14476 (N_14476,N_6312,N_9706);
xnor U14477 (N_14477,N_9238,N_7950);
or U14478 (N_14478,N_5086,N_8176);
and U14479 (N_14479,N_8158,N_5407);
nor U14480 (N_14480,N_6809,N_9752);
xnor U14481 (N_14481,N_9567,N_5010);
or U14482 (N_14482,N_8606,N_7789);
or U14483 (N_14483,N_6945,N_8195);
nor U14484 (N_14484,N_6219,N_8273);
and U14485 (N_14485,N_8072,N_7043);
xor U14486 (N_14486,N_5776,N_6580);
or U14487 (N_14487,N_6083,N_8165);
xnor U14488 (N_14488,N_8774,N_7574);
or U14489 (N_14489,N_5769,N_8469);
or U14490 (N_14490,N_6063,N_5621);
xor U14491 (N_14491,N_9036,N_7648);
nand U14492 (N_14492,N_5565,N_9254);
nor U14493 (N_14493,N_8809,N_5960);
and U14494 (N_14494,N_6050,N_5412);
xor U14495 (N_14495,N_5480,N_5608);
nor U14496 (N_14496,N_6941,N_5874);
or U14497 (N_14497,N_6595,N_7390);
or U14498 (N_14498,N_6215,N_7242);
nand U14499 (N_14499,N_6108,N_5875);
nor U14500 (N_14500,N_8891,N_7205);
nand U14501 (N_14501,N_6110,N_7571);
or U14502 (N_14502,N_6890,N_9129);
nand U14503 (N_14503,N_6888,N_8227);
or U14504 (N_14504,N_8302,N_8778);
and U14505 (N_14505,N_8335,N_6961);
nand U14506 (N_14506,N_5866,N_5644);
and U14507 (N_14507,N_9976,N_7969);
or U14508 (N_14508,N_6039,N_7403);
or U14509 (N_14509,N_8200,N_6365);
or U14510 (N_14510,N_9262,N_6145);
xor U14511 (N_14511,N_8421,N_7175);
nor U14512 (N_14512,N_6720,N_7183);
or U14513 (N_14513,N_5160,N_7672);
or U14514 (N_14514,N_8341,N_7558);
nor U14515 (N_14515,N_9966,N_5078);
nor U14516 (N_14516,N_7640,N_6609);
or U14517 (N_14517,N_7021,N_7576);
or U14518 (N_14518,N_5362,N_7956);
nor U14519 (N_14519,N_8773,N_6959);
xnor U14520 (N_14520,N_8446,N_7316);
nor U14521 (N_14521,N_7825,N_9898);
or U14522 (N_14522,N_5235,N_9156);
and U14523 (N_14523,N_6699,N_9409);
nand U14524 (N_14524,N_5675,N_9874);
nand U14525 (N_14525,N_9338,N_8380);
and U14526 (N_14526,N_9779,N_5059);
nand U14527 (N_14527,N_7018,N_5698);
and U14528 (N_14528,N_7515,N_5618);
and U14529 (N_14529,N_7403,N_6269);
xor U14530 (N_14530,N_8367,N_7070);
and U14531 (N_14531,N_8093,N_9573);
nor U14532 (N_14532,N_5744,N_7693);
and U14533 (N_14533,N_7464,N_5728);
and U14534 (N_14534,N_6751,N_9610);
or U14535 (N_14535,N_6353,N_9039);
nor U14536 (N_14536,N_5853,N_7684);
and U14537 (N_14537,N_7959,N_6985);
xnor U14538 (N_14538,N_8002,N_9170);
nor U14539 (N_14539,N_6484,N_7986);
or U14540 (N_14540,N_8868,N_5076);
nand U14541 (N_14541,N_7076,N_9050);
nand U14542 (N_14542,N_7077,N_5946);
and U14543 (N_14543,N_8788,N_7625);
and U14544 (N_14544,N_9289,N_6909);
nand U14545 (N_14545,N_8320,N_6004);
or U14546 (N_14546,N_7559,N_7986);
xnor U14547 (N_14547,N_7590,N_6460);
nand U14548 (N_14548,N_5450,N_8030);
or U14549 (N_14549,N_8288,N_8520);
nand U14550 (N_14550,N_7876,N_9792);
nor U14551 (N_14551,N_7644,N_5159);
and U14552 (N_14552,N_7446,N_9106);
xor U14553 (N_14553,N_5827,N_5936);
nor U14554 (N_14554,N_7220,N_7185);
or U14555 (N_14555,N_9794,N_9820);
nor U14556 (N_14556,N_7346,N_6619);
or U14557 (N_14557,N_6330,N_9932);
or U14558 (N_14558,N_5748,N_7938);
or U14559 (N_14559,N_9701,N_8888);
and U14560 (N_14560,N_9565,N_9067);
nand U14561 (N_14561,N_8454,N_8134);
nand U14562 (N_14562,N_8907,N_7092);
nand U14563 (N_14563,N_6313,N_5696);
nor U14564 (N_14564,N_5672,N_8570);
nor U14565 (N_14565,N_8260,N_8161);
nand U14566 (N_14566,N_5053,N_8489);
nor U14567 (N_14567,N_8376,N_6591);
xor U14568 (N_14568,N_8226,N_5950);
nor U14569 (N_14569,N_8581,N_9470);
nor U14570 (N_14570,N_5276,N_5408);
nor U14571 (N_14571,N_5658,N_6956);
and U14572 (N_14572,N_9182,N_5910);
or U14573 (N_14573,N_8645,N_8379);
nand U14574 (N_14574,N_9073,N_6526);
or U14575 (N_14575,N_7400,N_5227);
nand U14576 (N_14576,N_7170,N_8461);
nand U14577 (N_14577,N_8536,N_5632);
and U14578 (N_14578,N_9639,N_5747);
xnor U14579 (N_14579,N_9478,N_9731);
nor U14580 (N_14580,N_7932,N_7504);
and U14581 (N_14581,N_6447,N_5389);
or U14582 (N_14582,N_6514,N_9229);
nand U14583 (N_14583,N_5297,N_6854);
xnor U14584 (N_14584,N_6016,N_8354);
nor U14585 (N_14585,N_8056,N_7014);
nor U14586 (N_14586,N_6140,N_7349);
or U14587 (N_14587,N_7219,N_8920);
nand U14588 (N_14588,N_8224,N_5177);
and U14589 (N_14589,N_8018,N_7908);
xor U14590 (N_14590,N_7076,N_5061);
and U14591 (N_14591,N_8001,N_5007);
or U14592 (N_14592,N_7280,N_5791);
or U14593 (N_14593,N_5630,N_9349);
nand U14594 (N_14594,N_8948,N_5055);
or U14595 (N_14595,N_7110,N_6236);
xor U14596 (N_14596,N_5810,N_7550);
nand U14597 (N_14597,N_9254,N_8569);
and U14598 (N_14598,N_6129,N_7137);
nor U14599 (N_14599,N_9346,N_7116);
and U14600 (N_14600,N_9454,N_5695);
nor U14601 (N_14601,N_9540,N_7824);
and U14602 (N_14602,N_5931,N_5800);
nand U14603 (N_14603,N_7714,N_7503);
nand U14604 (N_14604,N_8508,N_6643);
nor U14605 (N_14605,N_7956,N_5660);
or U14606 (N_14606,N_5001,N_6256);
or U14607 (N_14607,N_5069,N_9994);
nor U14608 (N_14608,N_8646,N_9720);
and U14609 (N_14609,N_7240,N_6172);
and U14610 (N_14610,N_8607,N_9098);
nand U14611 (N_14611,N_5233,N_7300);
and U14612 (N_14612,N_9381,N_8554);
nor U14613 (N_14613,N_6870,N_7976);
nor U14614 (N_14614,N_9934,N_5724);
or U14615 (N_14615,N_5918,N_7200);
or U14616 (N_14616,N_6922,N_6039);
nor U14617 (N_14617,N_6549,N_5823);
or U14618 (N_14618,N_5489,N_8652);
or U14619 (N_14619,N_6107,N_5687);
or U14620 (N_14620,N_7844,N_8917);
nand U14621 (N_14621,N_6648,N_7138);
nor U14622 (N_14622,N_9477,N_7059);
nor U14623 (N_14623,N_6655,N_5858);
and U14624 (N_14624,N_7589,N_6906);
or U14625 (N_14625,N_8929,N_7490);
nor U14626 (N_14626,N_8469,N_6310);
nor U14627 (N_14627,N_5999,N_6162);
and U14628 (N_14628,N_6526,N_6350);
and U14629 (N_14629,N_6827,N_9369);
and U14630 (N_14630,N_7122,N_5209);
nand U14631 (N_14631,N_5748,N_5207);
xor U14632 (N_14632,N_6527,N_9800);
and U14633 (N_14633,N_6397,N_5713);
nand U14634 (N_14634,N_6944,N_9846);
or U14635 (N_14635,N_5523,N_8056);
or U14636 (N_14636,N_8790,N_8185);
and U14637 (N_14637,N_6910,N_8974);
and U14638 (N_14638,N_8452,N_9426);
or U14639 (N_14639,N_6940,N_5142);
nor U14640 (N_14640,N_5056,N_5318);
nor U14641 (N_14641,N_7223,N_8101);
nor U14642 (N_14642,N_8207,N_5856);
and U14643 (N_14643,N_8105,N_9748);
nand U14644 (N_14644,N_5778,N_6510);
or U14645 (N_14645,N_7060,N_7570);
or U14646 (N_14646,N_5598,N_8795);
or U14647 (N_14647,N_7500,N_6778);
and U14648 (N_14648,N_7844,N_8307);
nand U14649 (N_14649,N_5410,N_6946);
and U14650 (N_14650,N_6805,N_5547);
and U14651 (N_14651,N_5644,N_5743);
nor U14652 (N_14652,N_6986,N_5974);
nor U14653 (N_14653,N_5558,N_5704);
or U14654 (N_14654,N_5112,N_5287);
nand U14655 (N_14655,N_8793,N_9568);
nand U14656 (N_14656,N_9911,N_9604);
or U14657 (N_14657,N_5048,N_5942);
or U14658 (N_14658,N_5823,N_6621);
or U14659 (N_14659,N_7519,N_8012);
and U14660 (N_14660,N_9348,N_5768);
and U14661 (N_14661,N_9862,N_8803);
or U14662 (N_14662,N_7074,N_8234);
nand U14663 (N_14663,N_8581,N_7909);
and U14664 (N_14664,N_8221,N_9924);
or U14665 (N_14665,N_8133,N_7487);
nand U14666 (N_14666,N_7268,N_9094);
nand U14667 (N_14667,N_6844,N_5956);
and U14668 (N_14668,N_7131,N_7227);
nand U14669 (N_14669,N_8183,N_9163);
or U14670 (N_14670,N_7458,N_6186);
nand U14671 (N_14671,N_7293,N_9631);
nor U14672 (N_14672,N_9691,N_6681);
nand U14673 (N_14673,N_7387,N_7714);
nand U14674 (N_14674,N_8035,N_6567);
or U14675 (N_14675,N_5152,N_6305);
nor U14676 (N_14676,N_6756,N_9859);
nand U14677 (N_14677,N_5082,N_7653);
nand U14678 (N_14678,N_6126,N_9516);
nand U14679 (N_14679,N_6064,N_8158);
or U14680 (N_14680,N_5915,N_5950);
nor U14681 (N_14681,N_8562,N_9326);
nor U14682 (N_14682,N_6039,N_5587);
nor U14683 (N_14683,N_5874,N_7044);
or U14684 (N_14684,N_7749,N_6703);
nand U14685 (N_14685,N_9127,N_6807);
nand U14686 (N_14686,N_5209,N_6795);
and U14687 (N_14687,N_6174,N_9534);
nand U14688 (N_14688,N_8472,N_9987);
xnor U14689 (N_14689,N_6652,N_9803);
or U14690 (N_14690,N_5332,N_6157);
nor U14691 (N_14691,N_5124,N_7454);
nand U14692 (N_14692,N_6594,N_5415);
xnor U14693 (N_14693,N_7232,N_8035);
nand U14694 (N_14694,N_8852,N_7740);
and U14695 (N_14695,N_9706,N_8533);
nand U14696 (N_14696,N_8987,N_7489);
or U14697 (N_14697,N_5460,N_9812);
and U14698 (N_14698,N_7960,N_7852);
nand U14699 (N_14699,N_7108,N_6289);
nand U14700 (N_14700,N_6597,N_8780);
nand U14701 (N_14701,N_5574,N_7695);
and U14702 (N_14702,N_6634,N_7990);
xnor U14703 (N_14703,N_8752,N_6757);
nand U14704 (N_14704,N_9419,N_7097);
or U14705 (N_14705,N_6294,N_6587);
nor U14706 (N_14706,N_9916,N_6315);
and U14707 (N_14707,N_8933,N_9409);
nor U14708 (N_14708,N_8513,N_8191);
and U14709 (N_14709,N_7910,N_9136);
nand U14710 (N_14710,N_8732,N_5785);
nor U14711 (N_14711,N_5201,N_8084);
nor U14712 (N_14712,N_5659,N_5763);
xor U14713 (N_14713,N_7139,N_8672);
and U14714 (N_14714,N_6501,N_6520);
or U14715 (N_14715,N_6430,N_7292);
nor U14716 (N_14716,N_7175,N_8031);
and U14717 (N_14717,N_5370,N_7765);
nor U14718 (N_14718,N_8879,N_7854);
and U14719 (N_14719,N_7317,N_8492);
and U14720 (N_14720,N_6182,N_8473);
nand U14721 (N_14721,N_8218,N_5199);
nand U14722 (N_14722,N_8351,N_6719);
nor U14723 (N_14723,N_6749,N_5279);
nand U14724 (N_14724,N_8378,N_7664);
and U14725 (N_14725,N_8697,N_9597);
nor U14726 (N_14726,N_9831,N_5010);
nor U14727 (N_14727,N_9436,N_8096);
and U14728 (N_14728,N_5410,N_8033);
or U14729 (N_14729,N_9063,N_6435);
nor U14730 (N_14730,N_5983,N_9219);
and U14731 (N_14731,N_8236,N_5874);
nand U14732 (N_14732,N_8785,N_8598);
or U14733 (N_14733,N_5962,N_6638);
and U14734 (N_14734,N_6220,N_8747);
or U14735 (N_14735,N_6641,N_9688);
and U14736 (N_14736,N_8075,N_6434);
or U14737 (N_14737,N_5649,N_5856);
xnor U14738 (N_14738,N_6162,N_6316);
nor U14739 (N_14739,N_8608,N_5727);
nand U14740 (N_14740,N_9307,N_5883);
nor U14741 (N_14741,N_7492,N_9860);
nor U14742 (N_14742,N_9970,N_8744);
nor U14743 (N_14743,N_6133,N_9815);
nand U14744 (N_14744,N_7523,N_6651);
nor U14745 (N_14745,N_6017,N_5986);
or U14746 (N_14746,N_8741,N_9167);
xor U14747 (N_14747,N_8164,N_5612);
nand U14748 (N_14748,N_8113,N_6655);
or U14749 (N_14749,N_5124,N_9415);
and U14750 (N_14750,N_9037,N_6002);
and U14751 (N_14751,N_7219,N_8372);
and U14752 (N_14752,N_6100,N_8563);
nor U14753 (N_14753,N_8921,N_6357);
or U14754 (N_14754,N_7178,N_6365);
and U14755 (N_14755,N_6417,N_9058);
nor U14756 (N_14756,N_9049,N_7654);
nand U14757 (N_14757,N_6626,N_7199);
nor U14758 (N_14758,N_7839,N_7174);
nand U14759 (N_14759,N_9200,N_7539);
or U14760 (N_14760,N_7827,N_6944);
nand U14761 (N_14761,N_8914,N_7651);
nor U14762 (N_14762,N_8256,N_9538);
nor U14763 (N_14763,N_7680,N_6717);
and U14764 (N_14764,N_7149,N_8406);
xor U14765 (N_14765,N_6843,N_8121);
nand U14766 (N_14766,N_7410,N_7860);
and U14767 (N_14767,N_5957,N_5228);
and U14768 (N_14768,N_9065,N_9333);
and U14769 (N_14769,N_9386,N_9858);
nand U14770 (N_14770,N_5907,N_5576);
nand U14771 (N_14771,N_5221,N_9252);
nand U14772 (N_14772,N_7495,N_7603);
nor U14773 (N_14773,N_9901,N_6503);
and U14774 (N_14774,N_7499,N_9156);
nor U14775 (N_14775,N_8136,N_9382);
nand U14776 (N_14776,N_7499,N_8679);
xor U14777 (N_14777,N_9000,N_8064);
nor U14778 (N_14778,N_9479,N_6942);
nand U14779 (N_14779,N_9176,N_7921);
nor U14780 (N_14780,N_8906,N_6903);
nand U14781 (N_14781,N_7330,N_6165);
nor U14782 (N_14782,N_6110,N_9108);
nand U14783 (N_14783,N_8606,N_5516);
nand U14784 (N_14784,N_8283,N_8685);
nand U14785 (N_14785,N_7940,N_6331);
and U14786 (N_14786,N_9537,N_6784);
nor U14787 (N_14787,N_8151,N_7067);
nor U14788 (N_14788,N_6181,N_5717);
or U14789 (N_14789,N_9737,N_9024);
nor U14790 (N_14790,N_9748,N_6917);
and U14791 (N_14791,N_5760,N_9688);
or U14792 (N_14792,N_6444,N_7501);
and U14793 (N_14793,N_8815,N_9294);
and U14794 (N_14794,N_9279,N_8694);
nand U14795 (N_14795,N_5261,N_6282);
or U14796 (N_14796,N_5418,N_8761);
nor U14797 (N_14797,N_8344,N_7946);
and U14798 (N_14798,N_5053,N_8445);
xnor U14799 (N_14799,N_6173,N_6624);
nand U14800 (N_14800,N_9537,N_9466);
nand U14801 (N_14801,N_7600,N_8513);
or U14802 (N_14802,N_7675,N_9750);
and U14803 (N_14803,N_5385,N_6094);
and U14804 (N_14804,N_5314,N_5582);
nor U14805 (N_14805,N_6382,N_5076);
and U14806 (N_14806,N_7951,N_6651);
or U14807 (N_14807,N_7858,N_7921);
and U14808 (N_14808,N_5903,N_9172);
nor U14809 (N_14809,N_9014,N_7241);
xor U14810 (N_14810,N_5274,N_7368);
xnor U14811 (N_14811,N_7781,N_8245);
or U14812 (N_14812,N_8389,N_9786);
nor U14813 (N_14813,N_9707,N_6138);
and U14814 (N_14814,N_7259,N_9342);
nor U14815 (N_14815,N_7238,N_6990);
and U14816 (N_14816,N_7396,N_8220);
or U14817 (N_14817,N_8101,N_6462);
or U14818 (N_14818,N_7544,N_7420);
nand U14819 (N_14819,N_5662,N_5140);
and U14820 (N_14820,N_7610,N_5689);
nand U14821 (N_14821,N_8298,N_6483);
xor U14822 (N_14822,N_5561,N_9354);
and U14823 (N_14823,N_8475,N_6954);
and U14824 (N_14824,N_7963,N_5079);
xor U14825 (N_14825,N_9516,N_6567);
nand U14826 (N_14826,N_8643,N_9828);
and U14827 (N_14827,N_6221,N_5658);
or U14828 (N_14828,N_6293,N_8873);
or U14829 (N_14829,N_7705,N_8759);
xnor U14830 (N_14830,N_5261,N_7451);
nand U14831 (N_14831,N_6358,N_5486);
xor U14832 (N_14832,N_6094,N_7064);
and U14833 (N_14833,N_6529,N_5527);
xor U14834 (N_14834,N_7814,N_7898);
nor U14835 (N_14835,N_9528,N_8294);
nor U14836 (N_14836,N_9429,N_6153);
and U14837 (N_14837,N_5545,N_7292);
nand U14838 (N_14838,N_9531,N_7433);
xnor U14839 (N_14839,N_9511,N_9682);
xor U14840 (N_14840,N_6732,N_5080);
nor U14841 (N_14841,N_6999,N_5705);
and U14842 (N_14842,N_8088,N_7588);
nor U14843 (N_14843,N_7003,N_9731);
or U14844 (N_14844,N_6148,N_7654);
nand U14845 (N_14845,N_6537,N_7606);
or U14846 (N_14846,N_5832,N_8617);
nand U14847 (N_14847,N_7143,N_6117);
xnor U14848 (N_14848,N_5602,N_8017);
or U14849 (N_14849,N_5004,N_5686);
and U14850 (N_14850,N_7761,N_8309);
nor U14851 (N_14851,N_7613,N_6005);
nor U14852 (N_14852,N_6377,N_6274);
and U14853 (N_14853,N_9447,N_6244);
or U14854 (N_14854,N_9530,N_5566);
or U14855 (N_14855,N_8728,N_6725);
nor U14856 (N_14856,N_8032,N_5771);
or U14857 (N_14857,N_7717,N_9769);
xnor U14858 (N_14858,N_6476,N_7034);
nand U14859 (N_14859,N_9725,N_8467);
nor U14860 (N_14860,N_9338,N_8243);
nand U14861 (N_14861,N_6556,N_9539);
nand U14862 (N_14862,N_7696,N_8251);
nor U14863 (N_14863,N_8074,N_6765);
nand U14864 (N_14864,N_5917,N_9824);
nand U14865 (N_14865,N_9785,N_8396);
nor U14866 (N_14866,N_9700,N_9274);
nand U14867 (N_14867,N_6827,N_5163);
and U14868 (N_14868,N_8483,N_6569);
nand U14869 (N_14869,N_7849,N_9548);
or U14870 (N_14870,N_8591,N_7720);
nor U14871 (N_14871,N_6438,N_5109);
and U14872 (N_14872,N_8264,N_9857);
or U14873 (N_14873,N_5905,N_9204);
nor U14874 (N_14874,N_6292,N_7466);
or U14875 (N_14875,N_5721,N_6554);
and U14876 (N_14876,N_7131,N_5109);
nand U14877 (N_14877,N_5451,N_7020);
or U14878 (N_14878,N_9158,N_9566);
nand U14879 (N_14879,N_8526,N_8060);
nor U14880 (N_14880,N_8065,N_6251);
nand U14881 (N_14881,N_7380,N_8882);
and U14882 (N_14882,N_6550,N_8695);
xnor U14883 (N_14883,N_7532,N_6798);
nor U14884 (N_14884,N_7694,N_7153);
nor U14885 (N_14885,N_8881,N_6115);
nor U14886 (N_14886,N_9225,N_5985);
or U14887 (N_14887,N_8661,N_9056);
xor U14888 (N_14888,N_8460,N_6468);
nor U14889 (N_14889,N_5029,N_9885);
nand U14890 (N_14890,N_9605,N_9646);
or U14891 (N_14891,N_5100,N_8696);
or U14892 (N_14892,N_6750,N_7189);
and U14893 (N_14893,N_6058,N_6448);
nor U14894 (N_14894,N_9609,N_5285);
nand U14895 (N_14895,N_7414,N_6600);
nor U14896 (N_14896,N_7094,N_5035);
or U14897 (N_14897,N_5976,N_6381);
and U14898 (N_14898,N_5148,N_8301);
nand U14899 (N_14899,N_5005,N_9300);
and U14900 (N_14900,N_9976,N_5246);
or U14901 (N_14901,N_7564,N_8293);
nor U14902 (N_14902,N_7974,N_7352);
nand U14903 (N_14903,N_9858,N_8330);
nor U14904 (N_14904,N_6816,N_7204);
nor U14905 (N_14905,N_6726,N_9820);
nand U14906 (N_14906,N_5050,N_5049);
xnor U14907 (N_14907,N_5684,N_6998);
or U14908 (N_14908,N_9617,N_7361);
nor U14909 (N_14909,N_9040,N_8884);
nor U14910 (N_14910,N_8889,N_7241);
nand U14911 (N_14911,N_7788,N_8087);
and U14912 (N_14912,N_8303,N_8320);
or U14913 (N_14913,N_9027,N_6033);
or U14914 (N_14914,N_9137,N_6551);
or U14915 (N_14915,N_9127,N_8508);
nor U14916 (N_14916,N_8040,N_9532);
nand U14917 (N_14917,N_9743,N_6135);
or U14918 (N_14918,N_5444,N_8045);
or U14919 (N_14919,N_7326,N_8030);
nand U14920 (N_14920,N_8618,N_8225);
nor U14921 (N_14921,N_9421,N_8359);
nor U14922 (N_14922,N_7633,N_7645);
or U14923 (N_14923,N_8905,N_7042);
and U14924 (N_14924,N_8420,N_5084);
and U14925 (N_14925,N_6321,N_6024);
nand U14926 (N_14926,N_6163,N_6211);
and U14927 (N_14927,N_9918,N_5609);
nor U14928 (N_14928,N_5540,N_9731);
xnor U14929 (N_14929,N_5620,N_8538);
and U14930 (N_14930,N_6293,N_8196);
and U14931 (N_14931,N_9635,N_6502);
nand U14932 (N_14932,N_5909,N_5890);
or U14933 (N_14933,N_9516,N_7518);
nand U14934 (N_14934,N_5848,N_7832);
nor U14935 (N_14935,N_6026,N_5062);
or U14936 (N_14936,N_6696,N_7241);
nor U14937 (N_14937,N_6336,N_9356);
nor U14938 (N_14938,N_8881,N_6798);
nor U14939 (N_14939,N_5789,N_9944);
nand U14940 (N_14940,N_8674,N_7788);
xnor U14941 (N_14941,N_9890,N_9565);
nand U14942 (N_14942,N_5009,N_8661);
or U14943 (N_14943,N_6581,N_8080);
nor U14944 (N_14944,N_6980,N_9290);
nand U14945 (N_14945,N_6983,N_8031);
and U14946 (N_14946,N_9871,N_6355);
nand U14947 (N_14947,N_7289,N_8745);
and U14948 (N_14948,N_7969,N_5797);
nand U14949 (N_14949,N_9629,N_5029);
and U14950 (N_14950,N_7266,N_8947);
or U14951 (N_14951,N_9242,N_6443);
nand U14952 (N_14952,N_9044,N_6366);
nand U14953 (N_14953,N_7735,N_6128);
and U14954 (N_14954,N_7474,N_7155);
and U14955 (N_14955,N_9192,N_8929);
xor U14956 (N_14956,N_5716,N_8629);
nor U14957 (N_14957,N_7549,N_9030);
and U14958 (N_14958,N_9269,N_8397);
nor U14959 (N_14959,N_7449,N_6948);
xnor U14960 (N_14960,N_7316,N_6640);
and U14961 (N_14961,N_9224,N_6619);
nand U14962 (N_14962,N_9177,N_6725);
nor U14963 (N_14963,N_6262,N_5258);
nand U14964 (N_14964,N_6984,N_9372);
nor U14965 (N_14965,N_9890,N_6542);
nor U14966 (N_14966,N_9138,N_9120);
xnor U14967 (N_14967,N_8224,N_7598);
and U14968 (N_14968,N_9138,N_6462);
and U14969 (N_14969,N_9353,N_7658);
nand U14970 (N_14970,N_6911,N_7072);
or U14971 (N_14971,N_9791,N_5418);
nor U14972 (N_14972,N_8160,N_8747);
or U14973 (N_14973,N_7795,N_6857);
nor U14974 (N_14974,N_8080,N_5296);
nor U14975 (N_14975,N_5200,N_6227);
nor U14976 (N_14976,N_5423,N_6756);
and U14977 (N_14977,N_8218,N_8289);
and U14978 (N_14978,N_8206,N_5383);
nor U14979 (N_14979,N_5815,N_5434);
nand U14980 (N_14980,N_7685,N_6231);
nand U14981 (N_14981,N_7484,N_7580);
nand U14982 (N_14982,N_5709,N_5588);
nor U14983 (N_14983,N_8830,N_9646);
nand U14984 (N_14984,N_7098,N_5056);
nand U14985 (N_14985,N_9793,N_7714);
or U14986 (N_14986,N_5449,N_7907);
and U14987 (N_14987,N_8646,N_7114);
or U14988 (N_14988,N_6075,N_5728);
or U14989 (N_14989,N_9892,N_9080);
nor U14990 (N_14990,N_8031,N_8274);
nor U14991 (N_14991,N_6208,N_5608);
nand U14992 (N_14992,N_8328,N_7498);
or U14993 (N_14993,N_9350,N_9130);
nand U14994 (N_14994,N_6147,N_6036);
xnor U14995 (N_14995,N_9624,N_8834);
nand U14996 (N_14996,N_7186,N_9569);
xor U14997 (N_14997,N_9584,N_9526);
nor U14998 (N_14998,N_7260,N_5929);
nand U14999 (N_14999,N_7970,N_8016);
and U15000 (N_15000,N_10384,N_11669);
or U15001 (N_15001,N_10709,N_13463);
or U15002 (N_15002,N_13954,N_14715);
nand U15003 (N_15003,N_11857,N_11768);
and U15004 (N_15004,N_11547,N_14824);
nor U15005 (N_15005,N_13788,N_11086);
nor U15006 (N_15006,N_14840,N_13158);
or U15007 (N_15007,N_14023,N_10262);
nand U15008 (N_15008,N_10554,N_14744);
nor U15009 (N_15009,N_14149,N_14243);
nor U15010 (N_15010,N_14263,N_11896);
and U15011 (N_15011,N_11729,N_13748);
xnor U15012 (N_15012,N_13919,N_12446);
nand U15013 (N_15013,N_10926,N_13208);
xnor U15014 (N_15014,N_12106,N_12600);
nand U15015 (N_15015,N_14865,N_11194);
nand U15016 (N_15016,N_13172,N_13493);
xor U15017 (N_15017,N_13107,N_11270);
xnor U15018 (N_15018,N_10513,N_14027);
xnor U15019 (N_15019,N_12779,N_11332);
or U15020 (N_15020,N_14348,N_13785);
nand U15021 (N_15021,N_10663,N_10334);
nand U15022 (N_15022,N_13519,N_10886);
and U15023 (N_15023,N_13189,N_11654);
nor U15024 (N_15024,N_14695,N_14942);
and U15025 (N_15025,N_14338,N_10620);
nor U15026 (N_15026,N_12558,N_12041);
or U15027 (N_15027,N_14567,N_12533);
and U15028 (N_15028,N_14789,N_11662);
nor U15029 (N_15029,N_10588,N_10163);
and U15030 (N_15030,N_10067,N_11381);
or U15031 (N_15031,N_12334,N_10996);
nor U15032 (N_15032,N_10829,N_14725);
xnor U15033 (N_15033,N_10786,N_14532);
nand U15034 (N_15034,N_11433,N_14677);
and U15035 (N_15035,N_13373,N_12011);
or U15036 (N_15036,N_11962,N_12190);
nand U15037 (N_15037,N_10153,N_11755);
xor U15038 (N_15038,N_13180,N_14980);
or U15039 (N_15039,N_10116,N_11293);
or U15040 (N_15040,N_13371,N_11369);
nor U15041 (N_15041,N_14370,N_10354);
nor U15042 (N_15042,N_12240,N_14788);
or U15043 (N_15043,N_14321,N_13324);
nor U15044 (N_15044,N_13016,N_10167);
xor U15045 (N_15045,N_12869,N_14174);
nor U15046 (N_15046,N_11720,N_10047);
and U15047 (N_15047,N_10240,N_13144);
or U15048 (N_15048,N_12871,N_11621);
and U15049 (N_15049,N_10161,N_12112);
nand U15050 (N_15050,N_11338,N_13163);
or U15051 (N_15051,N_11680,N_10946);
and U15052 (N_15052,N_10617,N_11747);
or U15053 (N_15053,N_12731,N_13966);
or U15054 (N_15054,N_14833,N_12413);
nand U15055 (N_15055,N_11358,N_13214);
nand U15056 (N_15056,N_14945,N_14047);
nand U15057 (N_15057,N_10186,N_11902);
and U15058 (N_15058,N_12813,N_10940);
nand U15059 (N_15059,N_12142,N_12031);
and U15060 (N_15060,N_10509,N_13083);
or U15061 (N_15061,N_14965,N_12003);
or U15062 (N_15062,N_14608,N_12107);
and U15063 (N_15063,N_12627,N_14057);
and U15064 (N_15064,N_12485,N_12867);
xor U15065 (N_15065,N_13804,N_11651);
or U15066 (N_15066,N_14182,N_13282);
or U15067 (N_15067,N_14576,N_10526);
and U15068 (N_15068,N_10405,N_12396);
nand U15069 (N_15069,N_13732,N_14249);
or U15070 (N_15070,N_12966,N_10607);
nand U15071 (N_15071,N_13186,N_13945);
nor U15072 (N_15072,N_11942,N_11596);
nand U15073 (N_15073,N_11757,N_11064);
or U15074 (N_15074,N_14946,N_13146);
nor U15075 (N_15075,N_10254,N_12455);
nand U15076 (N_15076,N_12035,N_11493);
nand U15077 (N_15077,N_12159,N_10202);
or U15078 (N_15078,N_13676,N_11703);
or U15079 (N_15079,N_10846,N_11920);
or U15080 (N_15080,N_11744,N_11916);
nand U15081 (N_15081,N_14271,N_13625);
or U15082 (N_15082,N_12501,N_10619);
nor U15083 (N_15083,N_11003,N_12006);
or U15084 (N_15084,N_12258,N_13195);
and U15085 (N_15085,N_13478,N_12808);
nor U15086 (N_15086,N_13179,N_13225);
nand U15087 (N_15087,N_11829,N_12936);
and U15088 (N_15088,N_13366,N_11665);
or U15089 (N_15089,N_12656,N_12453);
nand U15090 (N_15090,N_10099,N_13504);
nor U15091 (N_15091,N_10928,N_14184);
nand U15092 (N_15092,N_12757,N_14966);
nand U15093 (N_15093,N_10566,N_13080);
nor U15094 (N_15094,N_13209,N_12196);
nand U15095 (N_15095,N_10534,N_12059);
and U15096 (N_15096,N_13817,N_13101);
nor U15097 (N_15097,N_11572,N_14687);
nor U15098 (N_15098,N_13269,N_11664);
or U15099 (N_15099,N_12493,N_10417);
nor U15100 (N_15100,N_11310,N_14866);
or U15101 (N_15101,N_10224,N_12676);
nand U15102 (N_15102,N_10982,N_13599);
or U15103 (N_15103,N_12042,N_14076);
or U15104 (N_15104,N_14728,N_10913);
and U15105 (N_15105,N_10632,N_10877);
nand U15106 (N_15106,N_14591,N_12171);
or U15107 (N_15107,N_12657,N_14955);
or U15108 (N_15108,N_12482,N_11778);
or U15109 (N_15109,N_11924,N_12391);
nor U15110 (N_15110,N_12166,N_13693);
nor U15111 (N_15111,N_13702,N_13616);
nor U15112 (N_15112,N_13433,N_12748);
nand U15113 (N_15113,N_13746,N_12296);
or U15114 (N_15114,N_14969,N_10227);
nor U15115 (N_15115,N_11058,N_13823);
or U15116 (N_15116,N_13484,N_14910);
nor U15117 (N_15117,N_13018,N_13281);
and U15118 (N_15118,N_13509,N_10994);
or U15119 (N_15119,N_12535,N_12462);
xnor U15120 (N_15120,N_12180,N_13729);
xnor U15121 (N_15121,N_14599,N_14198);
or U15122 (N_15122,N_13297,N_13948);
and U15123 (N_15123,N_12194,N_13452);
or U15124 (N_15124,N_14492,N_11307);
nor U15125 (N_15125,N_14374,N_13791);
and U15126 (N_15126,N_13940,N_10676);
and U15127 (N_15127,N_14381,N_11971);
nor U15128 (N_15128,N_11503,N_12433);
nor U15129 (N_15129,N_12122,N_10909);
and U15130 (N_15130,N_13759,N_12038);
or U15131 (N_15131,N_14595,N_13125);
xnor U15132 (N_15132,N_13538,N_14500);
nor U15133 (N_15133,N_14311,N_11475);
nor U15134 (N_15134,N_12505,N_14220);
or U15135 (N_15135,N_12203,N_13622);
or U15136 (N_15136,N_13411,N_11106);
or U15137 (N_15137,N_14967,N_13550);
nor U15138 (N_15138,N_12751,N_14250);
nand U15139 (N_15139,N_11653,N_14424);
and U15140 (N_15140,N_10021,N_11590);
and U15141 (N_15141,N_13754,N_10009);
or U15142 (N_15142,N_14718,N_14861);
nand U15143 (N_15143,N_13082,N_12425);
nand U15144 (N_15144,N_10299,N_10689);
and U15145 (N_15145,N_10824,N_10594);
or U15146 (N_15146,N_12328,N_10847);
nand U15147 (N_15147,N_11983,N_10369);
or U15148 (N_15148,N_13191,N_14901);
and U15149 (N_15149,N_14863,N_13304);
nor U15150 (N_15150,N_13378,N_10226);
nand U15151 (N_15151,N_10213,N_11026);
or U15152 (N_15152,N_14887,N_13003);
and U15153 (N_15153,N_12688,N_10557);
nor U15154 (N_15154,N_11889,N_11607);
and U15155 (N_15155,N_13812,N_11907);
nor U15156 (N_15156,N_11181,N_12037);
or U15157 (N_15157,N_13956,N_12089);
or U15158 (N_15158,N_11922,N_13007);
nand U15159 (N_15159,N_12992,N_13000);
nor U15160 (N_15160,N_10025,N_14937);
and U15161 (N_15161,N_14556,N_13672);
and U15162 (N_15162,N_14644,N_10542);
nor U15163 (N_15163,N_13887,N_12617);
or U15164 (N_15164,N_10000,N_13457);
nor U15165 (N_15165,N_12877,N_13884);
and U15166 (N_15166,N_11758,N_12795);
and U15167 (N_15167,N_14804,N_11776);
and U15168 (N_15168,N_11806,N_12665);
nor U15169 (N_15169,N_12113,N_11028);
nand U15170 (N_15170,N_10861,N_14948);
nor U15171 (N_15171,N_12358,N_14899);
and U15172 (N_15172,N_12909,N_14136);
or U15173 (N_15173,N_10631,N_11501);
nor U15174 (N_15174,N_11589,N_11144);
xor U15175 (N_15175,N_13372,N_10400);
nor U15176 (N_15176,N_12385,N_10683);
or U15177 (N_15177,N_11648,N_13204);
nor U15178 (N_15178,N_11089,N_10980);
or U15179 (N_15179,N_14118,N_12933);
or U15180 (N_15180,N_12917,N_14818);
and U15181 (N_15181,N_12478,N_13274);
nand U15182 (N_15182,N_11336,N_11670);
nor U15183 (N_15183,N_10667,N_11390);
or U15184 (N_15184,N_11859,N_10235);
nor U15185 (N_15185,N_14814,N_12963);
and U15186 (N_15186,N_14077,N_13421);
nand U15187 (N_15187,N_10406,N_14900);
nand U15188 (N_15188,N_11795,N_12233);
and U15189 (N_15189,N_10165,N_11031);
xnor U15190 (N_15190,N_12508,N_14086);
xnor U15191 (N_15191,N_12002,N_12199);
and U15192 (N_15192,N_12283,N_11134);
or U15193 (N_15193,N_11903,N_10825);
or U15194 (N_15194,N_12791,N_14206);
or U15195 (N_15195,N_14098,N_12284);
and U15196 (N_15196,N_14628,N_14357);
and U15197 (N_15197,N_13430,N_14375);
or U15198 (N_15198,N_12388,N_12934);
xor U15199 (N_15199,N_11414,N_11274);
or U15200 (N_15200,N_11199,N_13054);
nor U15201 (N_15201,N_14440,N_13863);
nor U15202 (N_15202,N_11397,N_10200);
or U15203 (N_15203,N_11966,N_13439);
nand U15204 (N_15204,N_11818,N_10193);
or U15205 (N_15205,N_11769,N_10083);
nor U15206 (N_15206,N_12781,N_11399);
and U15207 (N_15207,N_12322,N_13357);
nor U15208 (N_15208,N_10291,N_13066);
and U15209 (N_15209,N_11571,N_10423);
nor U15210 (N_15210,N_14002,N_13454);
nor U15211 (N_15211,N_14892,N_13675);
and U15212 (N_15212,N_13109,N_13276);
xnor U15213 (N_15213,N_10256,N_10698);
nand U15214 (N_15214,N_12929,N_10457);
nor U15215 (N_15215,N_14257,N_10989);
and U15216 (N_15216,N_12613,N_13402);
nand U15217 (N_15217,N_11588,N_14663);
nand U15218 (N_15218,N_12070,N_12928);
and U15219 (N_15219,N_10640,N_14771);
nor U15220 (N_15220,N_14778,N_11716);
xnor U15221 (N_15221,N_11137,N_12824);
or U15222 (N_15222,N_14620,N_10465);
nor U15223 (N_15223,N_11512,N_13403);
and U15224 (N_15224,N_14868,N_11772);
nand U15225 (N_15225,N_11153,N_10654);
or U15226 (N_15226,N_14803,N_13329);
nor U15227 (N_15227,N_11961,N_14734);
nor U15228 (N_15228,N_13898,N_14109);
nor U15229 (N_15229,N_14507,N_12949);
xor U15230 (N_15230,N_11504,N_11832);
nor U15231 (N_15231,N_13999,N_12143);
or U15232 (N_15232,N_13166,N_13854);
and U15233 (N_15233,N_11939,N_14296);
nor U15234 (N_15234,N_10769,N_10724);
xnor U15235 (N_15235,N_12753,N_12269);
nor U15236 (N_15236,N_14819,N_11843);
or U15237 (N_15237,N_12092,N_10930);
nand U15238 (N_15238,N_14380,N_10629);
and U15239 (N_15239,N_13476,N_11861);
xor U15240 (N_15240,N_11204,N_13181);
nand U15241 (N_15241,N_11619,N_14878);
nor U15242 (N_15242,N_12156,N_14860);
and U15243 (N_15243,N_12486,N_13775);
and U15244 (N_15244,N_13792,N_13374);
nand U15245 (N_15245,N_10844,N_12368);
and U15246 (N_15246,N_13260,N_13810);
or U15247 (N_15247,N_11905,N_13316);
and U15248 (N_15248,N_10879,N_11364);
or U15249 (N_15249,N_13258,N_14986);
or U15250 (N_15250,N_11482,N_12880);
nor U15251 (N_15251,N_10263,N_11506);
nor U15252 (N_15252,N_12518,N_13703);
nand U15253 (N_15253,N_13952,N_13992);
nor U15254 (N_15254,N_12502,N_14735);
nand U15255 (N_15255,N_14767,N_12695);
or U15256 (N_15256,N_11249,N_11929);
nor U15257 (N_15257,N_12421,N_13577);
nor U15258 (N_15258,N_10293,N_11344);
or U15259 (N_15259,N_11917,N_12348);
nor U15260 (N_15260,N_13049,N_11262);
nand U15261 (N_15261,N_13198,N_14686);
nor U15262 (N_15262,N_13710,N_11033);
and U15263 (N_15263,N_12175,N_14512);
nand U15264 (N_15264,N_10304,N_11746);
or U15265 (N_15265,N_14753,N_11909);
and U15266 (N_15266,N_13699,N_10501);
nand U15267 (N_15267,N_13879,N_13974);
and U15268 (N_15268,N_12739,N_12874);
or U15269 (N_15269,N_11613,N_11250);
nand U15270 (N_15270,N_13882,N_12990);
nor U15271 (N_15271,N_13574,N_11492);
or U15272 (N_15272,N_12723,N_14630);
nor U15273 (N_15273,N_14506,N_13038);
nand U15274 (N_15274,N_13385,N_12735);
and U15275 (N_15275,N_12044,N_13668);
and U15276 (N_15276,N_14444,N_13313);
nor U15277 (N_15277,N_11645,N_10691);
or U15278 (N_15278,N_10138,N_11237);
xor U15279 (N_15279,N_12087,N_11277);
nor U15280 (N_15280,N_14823,N_11289);
nor U15281 (N_15281,N_10484,N_12666);
nor U15282 (N_15282,N_12655,N_12794);
and U15283 (N_15283,N_12353,N_10455);
nor U15284 (N_15284,N_11944,N_11330);
nor U15285 (N_15285,N_13980,N_10333);
xnor U15286 (N_15286,N_11544,N_14080);
and U15287 (N_15287,N_12120,N_10908);
and U15288 (N_15288,N_12093,N_14383);
or U15289 (N_15289,N_14536,N_11533);
or U15290 (N_15290,N_12318,N_13012);
and U15291 (N_15291,N_11117,N_12046);
nor U15292 (N_15292,N_13850,N_12335);
and U15293 (N_15293,N_10636,N_14487);
nor U15294 (N_15294,N_13436,N_14325);
and U15295 (N_15295,N_10098,N_12177);
xnor U15296 (N_15296,N_11174,N_11240);
xnor U15297 (N_15297,N_10581,N_12057);
or U15298 (N_15298,N_10223,N_12321);
nand U15299 (N_15299,N_14028,N_13609);
and U15300 (N_15300,N_10366,N_10221);
and U15301 (N_15301,N_11419,N_10968);
xor U15302 (N_15302,N_12875,N_12952);
nand U15303 (N_15303,N_11182,N_12708);
and U15304 (N_15304,N_10220,N_11269);
nor U15305 (N_15305,N_13299,N_13397);
or U15306 (N_15306,N_12821,N_10562);
or U15307 (N_15307,N_10558,N_10476);
nor U15308 (N_15308,N_13869,N_13184);
and U15309 (N_15309,N_12235,N_12223);
nand U15310 (N_15310,N_12658,N_11597);
and U15311 (N_15311,N_13858,N_10856);
nand U15312 (N_15312,N_10643,N_14331);
nand U15313 (N_15313,N_12069,N_14958);
and U15314 (N_15314,N_14982,N_11035);
nor U15315 (N_15315,N_10335,N_12690);
nand U15316 (N_15316,N_13190,N_10425);
nand U15317 (N_15317,N_12341,N_10037);
nand U15318 (N_15318,N_10267,N_11140);
and U15319 (N_15319,N_13072,N_10954);
xor U15320 (N_15320,N_14442,N_13853);
nand U15321 (N_15321,N_10489,N_10478);
xor U15322 (N_15322,N_13408,N_12573);
nand U15323 (N_15323,N_10156,N_14390);
nand U15324 (N_15324,N_11996,N_11207);
nand U15325 (N_15325,N_11147,N_12189);
nor U15326 (N_15326,N_11835,N_10041);
or U15327 (N_15327,N_14720,N_10231);
or U15328 (N_15328,N_14830,N_12123);
xor U15329 (N_15329,N_13314,N_10967);
or U15330 (N_15330,N_10814,N_14073);
or U15331 (N_15331,N_13935,N_14631);
nor U15332 (N_15332,N_12725,N_13936);
and U15333 (N_15333,N_13838,N_13218);
and U15334 (N_15334,N_12601,N_13857);
nand U15335 (N_15335,N_14196,N_14733);
nand U15336 (N_15336,N_10445,N_12458);
or U15337 (N_15337,N_11868,N_14333);
nor U15338 (N_15338,N_10007,N_10528);
or U15339 (N_15339,N_11688,N_10488);
nor U15340 (N_15340,N_10260,N_12526);
or U15341 (N_15341,N_14448,N_13247);
or U15342 (N_15342,N_12095,N_14617);
nor U15343 (N_15343,N_12820,N_14645);
nor U15344 (N_15344,N_14713,N_10976);
and U15345 (N_15345,N_13630,N_10898);
xor U15346 (N_15346,N_10702,N_14597);
xnor U15347 (N_15347,N_10031,N_11520);
and U15348 (N_15348,N_10670,N_10784);
xnor U15349 (N_15349,N_13645,N_12300);
or U15350 (N_15350,N_10661,N_11687);
nand U15351 (N_15351,N_13132,N_11188);
or U15352 (N_15352,N_12243,N_13238);
nand U15353 (N_15353,N_14015,N_14849);
and U15354 (N_15354,N_14805,N_11311);
xnor U15355 (N_15355,N_11771,N_14745);
or U15356 (N_15356,N_14267,N_10342);
or U15357 (N_15357,N_12540,N_13486);
xnor U15358 (N_15358,N_14402,N_10712);
and U15359 (N_15359,N_12027,N_13951);
and U15360 (N_15360,N_14766,N_13285);
nand U15361 (N_15361,N_14854,N_11566);
or U15362 (N_15362,N_11160,N_12800);
or U15363 (N_15363,N_13025,N_11745);
nor U15364 (N_15364,N_13819,N_11103);
nand U15365 (N_15365,N_13438,N_11075);
nand U15366 (N_15366,N_14163,N_14721);
and U15367 (N_15367,N_10816,N_10149);
or U15368 (N_15368,N_11488,N_14431);
and U15369 (N_15369,N_13920,N_14452);
and U15370 (N_15370,N_10807,N_10337);
nor U15371 (N_15371,N_10269,N_11792);
nor U15372 (N_15372,N_10531,N_13392);
or U15373 (N_15373,N_13152,N_12839);
nor U15374 (N_15374,N_13683,N_14238);
and U15375 (N_15375,N_12103,N_12705);
nor U15376 (N_15376,N_10664,N_11649);
and U15377 (N_15377,N_14498,N_11751);
nand U15378 (N_15378,N_14758,N_14592);
or U15379 (N_15379,N_11759,N_12392);
nand U15380 (N_15380,N_13878,N_13168);
nand U15381 (N_15381,N_10216,N_13926);
or U15382 (N_15382,N_11954,N_13727);
or U15383 (N_15383,N_12611,N_13808);
or U15384 (N_15384,N_11047,N_10541);
and U15385 (N_15385,N_12908,N_13291);
and U15386 (N_15386,N_11846,N_14276);
xor U15387 (N_15387,N_14575,N_10572);
nor U15388 (N_15388,N_12043,N_13239);
and U15389 (N_15389,N_14685,N_14699);
or U15390 (N_15390,N_12288,N_10027);
nand U15391 (N_15391,N_14670,N_10701);
nor U15392 (N_15392,N_10274,N_12568);
or U15393 (N_15393,N_14067,N_14843);
xnor U15394 (N_15394,N_13903,N_10307);
nor U15395 (N_15395,N_10377,N_13010);
nor U15396 (N_15396,N_13753,N_14459);
and U15397 (N_15397,N_13097,N_14682);
xnor U15398 (N_15398,N_13818,N_10834);
nor U15399 (N_15399,N_11581,N_14975);
and U15400 (N_15400,N_10345,N_12067);
nor U15401 (N_15401,N_14143,N_11908);
nand U15402 (N_15402,N_14129,N_14615);
nand U15403 (N_15403,N_14898,N_14283);
or U15404 (N_15404,N_12629,N_10907);
nor U15405 (N_15405,N_10111,N_13883);
or U15406 (N_15406,N_12538,N_12983);
xor U15407 (N_15407,N_14139,N_14223);
and U15408 (N_15408,N_14880,N_12221);
and U15409 (N_15409,N_10941,N_11368);
and U15410 (N_15410,N_14489,N_12303);
and U15411 (N_15411,N_10107,N_13626);
and U15412 (N_15412,N_14069,N_10830);
or U15413 (N_15413,N_12995,N_10325);
nand U15414 (N_15414,N_13388,N_14233);
xor U15415 (N_15415,N_14821,N_14499);
nand U15416 (N_15416,N_14688,N_11056);
and U15417 (N_15417,N_14648,N_10214);
nand U15418 (N_15418,N_12536,N_10507);
nand U15419 (N_15419,N_14280,N_13736);
xor U15420 (N_15420,N_10942,N_13073);
nor U15421 (N_15421,N_13221,N_11816);
nand U15422 (N_15422,N_11893,N_13071);
or U15423 (N_15423,N_13338,N_14398);
or U15424 (N_15424,N_12523,N_12596);
nor U15425 (N_15425,N_12620,N_11434);
nand U15426 (N_15426,N_13288,N_10132);
and U15427 (N_15427,N_14650,N_11214);
nand U15428 (N_15428,N_14405,N_11025);
or U15429 (N_15429,N_10438,N_12320);
or U15430 (N_15430,N_14160,N_10399);
nor U15431 (N_15431,N_10551,N_14672);
or U15432 (N_15432,N_11709,N_10641);
or U15433 (N_15433,N_11158,N_13053);
nand U15434 (N_15434,N_11387,N_11515);
xnor U15435 (N_15435,N_14722,N_14740);
xor U15436 (N_15436,N_11335,N_14943);
nor U15437 (N_15437,N_10746,N_12647);
nor U15438 (N_15438,N_14320,N_11932);
nor U15439 (N_15439,N_14540,N_11405);
and U15440 (N_15440,N_10560,N_12623);
nor U15441 (N_15441,N_11061,N_11694);
or U15442 (N_15442,N_10287,N_13498);
and U15443 (N_15443,N_10755,N_13489);
and U15444 (N_15444,N_14435,N_10963);
nor U15445 (N_15445,N_11781,N_14476);
and U15446 (N_15446,N_13289,N_13485);
or U15447 (N_15447,N_11317,N_13468);
or U15448 (N_15448,N_12740,N_10152);
and U15449 (N_15449,N_11647,N_14230);
nand U15450 (N_15450,N_12977,N_12152);
or U15451 (N_15451,N_12055,N_11513);
and U15452 (N_15452,N_13995,N_10756);
nor U15453 (N_15453,N_14853,N_14112);
nor U15454 (N_15454,N_12032,N_12273);
nor U15455 (N_15455,N_13658,N_12706);
nand U15456 (N_15456,N_14451,N_13922);
or U15457 (N_15457,N_10411,N_10800);
nor U15458 (N_15458,N_11725,N_13110);
and U15459 (N_15459,N_14949,N_13226);
xor U15460 (N_15460,N_14146,N_10114);
and U15461 (N_15461,N_11895,N_10385);
nand U15462 (N_15462,N_13119,N_13063);
nor U15463 (N_15463,N_12589,N_10753);
and U15464 (N_15464,N_14903,N_11398);
and U15465 (N_15465,N_11363,N_12479);
or U15466 (N_15466,N_10129,N_12039);
nand U15467 (N_15467,N_11287,N_12605);
nand U15468 (N_15468,N_12844,N_10833);
nor U15469 (N_15469,N_13350,N_12692);
or U15470 (N_15470,N_11360,N_11327);
nor U15471 (N_15471,N_14134,N_11637);
nor U15472 (N_15472,N_11611,N_14791);
and U15473 (N_15473,N_12270,N_13934);
nor U15474 (N_15474,N_11676,N_12772);
nand U15475 (N_15475,N_13345,N_13752);
nand U15476 (N_15476,N_13740,N_11455);
nand U15477 (N_15477,N_10196,N_13585);
nor U15478 (N_15478,N_14179,N_11068);
and U15479 (N_15479,N_11558,N_10920);
or U15480 (N_15480,N_12506,N_11638);
nor U15481 (N_15481,N_14428,N_12248);
nand U15482 (N_15482,N_10246,N_10778);
nor U15483 (N_15483,N_11518,N_11876);
nor U15484 (N_15484,N_13722,N_11690);
and U15485 (N_15485,N_14756,N_12846);
or U15486 (N_15486,N_14944,N_13986);
xnor U15487 (N_15487,N_10183,N_13985);
nand U15488 (N_15488,N_11490,N_11914);
or U15489 (N_15489,N_13603,N_14683);
xor U15490 (N_15490,N_12661,N_14546);
and U15491 (N_15491,N_14749,N_14570);
nor U15492 (N_15492,N_14344,N_11704);
xnor U15493 (N_15493,N_10840,N_10750);
and U15494 (N_15494,N_11367,N_13036);
xor U15495 (N_15495,N_14963,N_13462);
nand U15496 (N_15496,N_13892,N_10001);
nand U15497 (N_15497,N_12804,N_14054);
xnor U15498 (N_15498,N_13721,N_13904);
nand U15499 (N_15499,N_12153,N_11657);
nor U15500 (N_15500,N_12492,N_13881);
nor U15501 (N_15501,N_11842,N_12566);
and U15502 (N_15502,N_12681,N_14148);
nand U15503 (N_15503,N_10684,N_13091);
and U15504 (N_15504,N_12590,N_13346);
nor U15505 (N_15505,N_12197,N_11855);
nand U15506 (N_15506,N_14164,N_10229);
and U15507 (N_15507,N_13939,N_14173);
xnor U15508 (N_15508,N_12671,N_12733);
xor U15509 (N_15509,N_14404,N_12304);
and U15510 (N_15510,N_12521,N_13268);
or U15511 (N_15511,N_10441,N_10972);
or U15512 (N_15512,N_12884,N_14389);
nand U15513 (N_15513,N_10243,N_11601);
nand U15514 (N_15514,N_12554,N_14310);
nor U15515 (N_15515,N_13156,N_11883);
and U15516 (N_15516,N_10593,N_13773);
nand U15517 (N_15517,N_11984,N_13781);
nor U15518 (N_15518,N_11750,N_10300);
or U15519 (N_15519,N_12763,N_10681);
nor U15520 (N_15520,N_12634,N_13045);
nor U15521 (N_15521,N_12139,N_12991);
nand U15522 (N_15522,N_13787,N_14445);
nor U15523 (N_15523,N_12912,N_14484);
and U15524 (N_15524,N_14928,N_13094);
nand U15525 (N_15525,N_13507,N_13605);
and U15526 (N_15526,N_10845,N_10318);
nand U15527 (N_15527,N_13834,N_11784);
nor U15528 (N_15528,N_14577,N_12709);
or U15529 (N_15529,N_14183,N_14675);
nor U15530 (N_15530,N_14413,N_12097);
and U15531 (N_15531,N_12749,N_10969);
nand U15532 (N_15532,N_13634,N_11510);
or U15533 (N_15533,N_11472,N_13816);
xor U15534 (N_15534,N_11192,N_10276);
nor U15535 (N_15535,N_14780,N_10303);
nor U15536 (N_15536,N_12215,N_12593);
nor U15537 (N_15537,N_10789,N_10462);
nor U15538 (N_15538,N_14940,N_14613);
nand U15539 (N_15539,N_10705,N_12683);
nand U15540 (N_15540,N_12842,N_14053);
nand U15541 (N_15541,N_10207,N_11266);
or U15542 (N_15542,N_14342,N_12764);
and U15543 (N_15543,N_11881,N_12732);
xnor U15544 (N_15544,N_11673,N_11525);
nand U15545 (N_15545,N_13901,N_12459);
xnor U15546 (N_15546,N_11775,N_10956);
nor U15547 (N_15547,N_11685,N_10238);
nor U15548 (N_15548,N_11614,N_11275);
nand U15549 (N_15549,N_12911,N_10537);
and U15550 (N_15550,N_13306,N_12405);
nand U15551 (N_15551,N_14152,N_12220);
or U15552 (N_15552,N_13905,N_10865);
xnor U15553 (N_15553,N_11284,N_11319);
nand U15554 (N_15554,N_12803,N_13597);
or U15555 (N_15555,N_13294,N_11467);
nand U15556 (N_15556,N_14231,N_13113);
nand U15557 (N_15557,N_14065,N_13118);
nand U15558 (N_15558,N_10527,N_14317);
nand U15559 (N_15559,N_12294,N_14925);
and U15560 (N_15560,N_12347,N_12609);
and U15561 (N_15561,N_12150,N_11221);
or U15562 (N_15562,N_14711,N_13728);
nand U15563 (N_15563,N_13455,N_12470);
nor U15564 (N_15564,N_13050,N_10977);
and U15565 (N_15565,N_12339,N_10821);
nor U15566 (N_15566,N_11197,N_11162);
nand U15567 (N_15567,N_10352,N_13915);
nor U15568 (N_15568,N_12178,N_12342);
nor U15569 (N_15569,N_12583,N_10069);
or U15570 (N_15570,N_10854,N_12469);
and U15571 (N_15571,N_10812,N_10250);
xor U15572 (N_15572,N_13602,N_12149);
or U15573 (N_15573,N_11696,N_14364);
nor U15574 (N_15574,N_12274,N_11679);
nor U15575 (N_15575,N_12389,N_14995);
nor U15576 (N_15576,N_14488,N_11591);
xnor U15577 (N_15577,N_14355,N_14605);
nor U15578 (N_15578,N_13257,N_12841);
and U15579 (N_15579,N_11006,N_11788);
or U15580 (N_15580,N_13868,N_13275);
or U15581 (N_15581,N_12053,N_10410);
and U15582 (N_15582,N_10564,N_13309);
nor U15583 (N_15583,N_10095,N_14952);
or U15584 (N_15584,N_14318,N_10515);
nor U15585 (N_15585,N_12840,N_14478);
or U15586 (N_15586,N_11969,N_13972);
xnor U15587 (N_15587,N_11576,N_10780);
or U15588 (N_15588,N_10477,N_11109);
xnor U15589 (N_15589,N_14950,N_10835);
nand U15590 (N_15590,N_14578,N_12099);
or U15591 (N_15591,N_11051,N_14420);
and U15592 (N_15592,N_14561,N_11285);
and U15593 (N_15593,N_11667,N_14839);
nor U15594 (N_15594,N_11982,N_13328);
or U15595 (N_15595,N_11019,N_11113);
nand U15596 (N_15596,N_14792,N_10358);
nand U15597 (N_15597,N_10241,N_14759);
nand U15598 (N_15598,N_14956,N_12578);
nor U15599 (N_15599,N_10723,N_10890);
or U15600 (N_15600,N_13031,N_10815);
or U15601 (N_15601,N_12287,N_11149);
and U15602 (N_15602,N_11029,N_11957);
or U15603 (N_15603,N_14905,N_13444);
nor U15604 (N_15604,N_12997,N_12116);
nand U15605 (N_15605,N_13395,N_10894);
and U15606 (N_15606,N_11706,N_10210);
and U15607 (N_15607,N_10123,N_12360);
and U15608 (N_15608,N_11447,N_13687);
xor U15609 (N_15609,N_11574,N_11615);
and U15610 (N_15610,N_10888,N_11459);
nor U15611 (N_15611,N_12445,N_13930);
and U15612 (N_15612,N_13765,N_14837);
and U15613 (N_15613,N_13173,N_11339);
or U15614 (N_15614,N_13377,N_12336);
and U15615 (N_15615,N_14841,N_13011);
xnor U15616 (N_15616,N_13789,N_14889);
xor U15617 (N_15617,N_12560,N_14268);
nand U15618 (N_15618,N_12078,N_12693);
or U15619 (N_15619,N_12712,N_11371);
or U15620 (N_15620,N_13440,N_10586);
xnor U15621 (N_15621,N_13551,N_12192);
or U15622 (N_15622,N_10295,N_12514);
nor U15623 (N_15623,N_11139,N_13755);
and U15624 (N_15624,N_13565,N_14135);
nor U15625 (N_15625,N_11502,N_14014);
xnor U15626 (N_15626,N_14813,N_11392);
and U15627 (N_15627,N_11626,N_14794);
or U15628 (N_15628,N_11438,N_12982);
and U15629 (N_15629,N_10394,N_13213);
and U15630 (N_15630,N_12686,N_13825);
and U15631 (N_15631,N_10211,N_10265);
nand U15632 (N_15632,N_10370,N_14913);
and U15633 (N_15633,N_11427,N_10320);
and U15634 (N_15634,N_13692,N_12713);
or U15635 (N_15635,N_10868,N_14423);
and U15636 (N_15636,N_13733,N_11076);
nand U15637 (N_15637,N_12048,N_13977);
nor U15638 (N_15638,N_13685,N_12610);
or U15639 (N_15639,N_10233,N_11041);
or U15640 (N_15640,N_10321,N_12516);
nand U15641 (N_15641,N_11837,N_10759);
xnor U15642 (N_15642,N_14590,N_11494);
or U15643 (N_15643,N_14864,N_10360);
nor U15644 (N_15644,N_14292,N_10434);
nor U15645 (N_15645,N_11135,N_11489);
xnor U15646 (N_15646,N_11634,N_12016);
and U15647 (N_15647,N_12582,N_11044);
and U15648 (N_15648,N_14602,N_14563);
nand U15649 (N_15649,N_13876,N_13735);
or U15650 (N_15650,N_11904,N_11550);
or U15651 (N_15651,N_11925,N_10783);
or U15652 (N_15652,N_11879,N_12372);
or U15653 (N_15653,N_14643,N_13296);
and U15654 (N_15654,N_12102,N_11131);
xor U15655 (N_15655,N_12383,N_14291);
nand U15656 (N_15656,N_13279,N_13448);
nand U15657 (N_15657,N_12530,N_13480);
nor U15658 (N_15658,N_13143,N_11575);
nand U15659 (N_15659,N_13960,N_14553);
or U15660 (N_15660,N_13106,N_11717);
xor U15661 (N_15661,N_12571,N_13580);
nand U15662 (N_15662,N_10016,N_14657);
xor U15663 (N_15663,N_10311,N_10764);
and U15664 (N_15664,N_11431,N_12504);
nor U15665 (N_15665,N_14209,N_12562);
xnor U15666 (N_15666,N_12023,N_13908);
nor U15667 (N_15667,N_13386,N_13020);
xnor U15668 (N_15668,N_11660,N_13997);
or U15669 (N_15669,N_12823,N_12004);
and U15670 (N_15670,N_11440,N_11499);
nand U15671 (N_15671,N_10466,N_11623);
and U15672 (N_15672,N_10768,N_14137);
nand U15673 (N_15673,N_12984,N_10869);
nand U15674 (N_15674,N_10440,N_11543);
nor U15675 (N_15675,N_10014,N_10166);
and U15676 (N_15676,N_14464,N_12927);
xnor U15677 (N_15677,N_14379,N_12013);
nand U15678 (N_15678,N_11989,N_10960);
xor U15679 (N_15679,N_12956,N_12151);
nand U15680 (N_15680,N_10131,N_12170);
or U15681 (N_15681,N_14345,N_11733);
nor U15682 (N_15682,N_12071,N_14051);
nand U15683 (N_15683,N_10732,N_10727);
or U15684 (N_15684,N_11362,N_14585);
or U15685 (N_15685,N_11451,N_10912);
or U15686 (N_15686,N_10573,N_12338);
xor U15687 (N_15687,N_10585,N_12987);
or U15688 (N_15688,N_10657,N_11910);
or U15689 (N_15689,N_10426,N_11195);
nor U15690 (N_15690,N_12507,N_12637);
nand U15691 (N_15691,N_14165,N_14366);
and U15692 (N_15692,N_10073,N_12260);
xor U15693 (N_15693,N_14361,N_13375);
nor U15694 (N_15694,N_11196,N_11042);
xnor U15695 (N_15695,N_12423,N_11777);
nor U15696 (N_15696,N_10748,N_13414);
and U15697 (N_15697,N_11691,N_11477);
nor U15698 (N_15698,N_12866,N_10180);
xor U15699 (N_15699,N_10546,N_14679);
or U15700 (N_15700,N_12761,N_10822);
nand U15701 (N_15701,N_12265,N_14213);
and U15702 (N_15702,N_12268,N_13795);
and U15703 (N_15703,N_10737,N_14689);
xor U15704 (N_15704,N_10891,N_13569);
or U15705 (N_15705,N_12553,N_11994);
nor U15706 (N_15706,N_10916,N_12905);
nand U15707 (N_15707,N_10178,N_14646);
nand U15708 (N_15708,N_10015,N_10219);
nor U15709 (N_15709,N_11354,N_12612);
or U15710 (N_15710,N_12750,N_11830);
or U15711 (N_15711,N_14539,N_14772);
nand U15712 (N_15712,N_10962,N_10716);
and U15713 (N_15713,N_10085,N_13040);
and U15714 (N_15714,N_11450,N_14218);
and U15715 (N_15715,N_14096,N_13767);
and U15716 (N_15716,N_12014,N_12138);
or U15717 (N_15717,N_13250,N_10625);
or U15718 (N_15718,N_12836,N_14158);
or U15719 (N_15719,N_12052,N_14011);
and U15720 (N_15720,N_13065,N_13662);
nor U15721 (N_15721,N_11396,N_14960);
or U15722 (N_15722,N_14309,N_14285);
and U15723 (N_15723,N_13393,N_14612);
nand U15724 (N_15724,N_13192,N_11443);
or U15725 (N_15725,N_13093,N_13514);
nor U15726 (N_15726,N_11341,N_10029);
nand U15727 (N_15727,N_12483,N_11378);
nor U15728 (N_15728,N_13280,N_11290);
or U15729 (N_15729,N_10120,N_13177);
or U15730 (N_15730,N_12957,N_13679);
and U15731 (N_15731,N_11655,N_13128);
or U15732 (N_15732,N_13562,N_10185);
xnor U15733 (N_15733,N_12344,N_14166);
and U15734 (N_15734,N_14929,N_11542);
and U15735 (N_15735,N_11132,N_14094);
nor U15736 (N_15736,N_12255,N_10222);
xnor U15737 (N_15737,N_11748,N_11138);
nand U15738 (N_15738,N_14760,N_14706);
and U15739 (N_15739,N_13505,N_14300);
and U15740 (N_15740,N_11605,N_13861);
or U15741 (N_15741,N_14113,N_11177);
nor U15742 (N_15742,N_11684,N_10239);
and U15743 (N_15743,N_11951,N_13617);
and U15744 (N_15744,N_13358,N_10642);
or U15745 (N_15745,N_13586,N_13111);
nor U15746 (N_15746,N_14930,N_12088);
or U15747 (N_15747,N_11342,N_10595);
or U15748 (N_15748,N_10046,N_13990);
nor U15749 (N_15749,N_10981,N_10790);
xnor U15750 (N_15750,N_10674,N_10191);
nand U15751 (N_15751,N_13720,N_13557);
and U15752 (N_15752,N_10376,N_14520);
or U15753 (N_15753,N_14842,N_14013);
nor U15754 (N_15754,N_10703,N_11236);
nor U15755 (N_15755,N_14883,N_13983);
nand U15756 (N_15756,N_12094,N_13174);
or U15757 (N_15757,N_12913,N_12947);
or U15758 (N_15758,N_12818,N_11836);
nand U15759 (N_15759,N_14573,N_13413);
nand U15760 (N_15760,N_12182,N_13872);
xor U15761 (N_15761,N_12432,N_11404);
or U15762 (N_15762,N_12663,N_14251);
nand U15763 (N_15763,N_10288,N_12026);
or U15764 (N_15764,N_11541,N_10413);
nand U15765 (N_15765,N_12576,N_13591);
nor U15766 (N_15766,N_11231,N_12049);
nand U15767 (N_15767,N_12444,N_14221);
or U15768 (N_15768,N_11432,N_11858);
xor U15769 (N_15769,N_10497,N_12789);
and U15770 (N_15770,N_14629,N_13911);
nand U15771 (N_15771,N_13487,N_10378);
nor U15772 (N_15772,N_10372,N_11726);
nand U15773 (N_15773,N_12145,N_13263);
or U15774 (N_15774,N_13176,N_13417);
nand U15775 (N_15775,N_10953,N_13157);
nor U15776 (N_15776,N_12371,N_12250);
nor U15777 (N_15777,N_10524,N_13370);
nand U15778 (N_15778,N_12585,N_12948);
and U15779 (N_15779,N_10182,N_11585);
or U15780 (N_15780,N_13099,N_11785);
xor U15781 (N_15781,N_10802,N_12263);
or U15782 (N_15782,N_11524,N_11980);
nor U15783 (N_15783,N_13084,N_10957);
nor U15784 (N_15784,N_12525,N_12163);
nor U15785 (N_15785,N_14193,N_14660);
and U15786 (N_15786,N_11424,N_13167);
xor U15787 (N_15787,N_11583,N_10090);
and U15788 (N_15788,N_10452,N_13449);
or U15789 (N_15789,N_11241,N_13806);
nand U15790 (N_15790,N_14081,N_10831);
and U15791 (N_15791,N_10449,N_10395);
nand U15792 (N_15792,N_14527,N_14017);
nand U15793 (N_15793,N_13963,N_10547);
or U15794 (N_15794,N_12015,N_13637);
nor U15795 (N_15795,N_10600,N_10089);
xor U15796 (N_15796,N_12759,N_12330);
or U15797 (N_15797,N_14588,N_13653);
nand U15798 (N_15798,N_12548,N_11933);
nand U15799 (N_15799,N_10770,N_13148);
nor U15800 (N_15800,N_14964,N_14907);
nor U15801 (N_15801,N_11847,N_12958);
nor U15802 (N_15802,N_14664,N_13666);
or U15803 (N_15803,N_10901,N_13578);
nor U15804 (N_15804,N_12876,N_13691);
nor U15805 (N_15805,N_10146,N_13913);
nand U15806 (N_15806,N_12186,N_10419);
nor U15807 (N_15807,N_10382,N_14748);
xnor U15808 (N_15808,N_13886,N_14048);
and U15809 (N_15809,N_10284,N_10252);
xor U15810 (N_15810,N_11507,N_11213);
and U15811 (N_15811,N_11186,N_14084);
nand U15812 (N_15812,N_13632,N_13828);
and U15813 (N_15813,N_11620,N_14496);
and U15814 (N_15814,N_14996,N_13867);
nand U15815 (N_15815,N_13236,N_12137);
xor U15816 (N_15816,N_12500,N_11415);
xor U15817 (N_15817,N_13273,N_11172);
and U15818 (N_15818,N_11325,N_14426);
and U15819 (N_15819,N_10610,N_10195);
xor U15820 (N_15820,N_12664,N_14399);
or U15821 (N_15821,N_11953,N_13014);
nand U15822 (N_15822,N_11097,N_10057);
xnor U15823 (N_15823,N_10743,N_11331);
and U15824 (N_15824,N_12953,N_11435);
nor U15825 (N_15825,N_10777,N_14121);
or U15826 (N_15826,N_11445,N_10757);
nand U15827 (N_15827,N_10787,N_13984);
and U15828 (N_15828,N_13145,N_10164);
nand U15829 (N_15829,N_11255,N_12404);
or U15830 (N_15830,N_13394,N_13826);
nand U15831 (N_15831,N_10791,N_11294);
nand U15832 (N_15832,N_12855,N_10061);
nand U15833 (N_15833,N_13978,N_14003);
and U15834 (N_15834,N_11804,N_13535);
and U15835 (N_15835,N_10051,N_14055);
xnor U15836 (N_15836,N_11373,N_13559);
xnor U15837 (N_15837,N_13965,N_11412);
xnor U15838 (N_15838,N_12701,N_10647);
and U15839 (N_15839,N_10242,N_14639);
or U15840 (N_15840,N_13548,N_11663);
nor U15841 (N_15841,N_13103,N_14343);
and U15842 (N_15842,N_11538,N_10711);
and U15843 (N_15843,N_14684,N_14558);
xor U15844 (N_15844,N_11463,N_12411);
or U15845 (N_15845,N_13596,N_10719);
nor U15846 (N_15846,N_12403,N_11304);
and U15847 (N_15847,N_13379,N_14875);
xor U15848 (N_15848,N_14755,N_11299);
nand U15849 (N_15849,N_13220,N_13640);
and U15850 (N_15850,N_10583,N_13312);
or U15851 (N_15851,N_12440,N_10899);
nor U15852 (N_15852,N_11115,N_13416);
or U15853 (N_15853,N_11529,N_14265);
nand U15854 (N_15854,N_14882,N_11462);
and U15855 (N_15855,N_11024,N_10838);
and U15856 (N_15856,N_12136,N_14095);
or U15857 (N_15857,N_10003,N_14394);
nor U15858 (N_15858,N_11243,N_14990);
nor U15859 (N_15859,N_10843,N_12050);
and U15860 (N_15860,N_11272,N_14241);
or U15861 (N_15861,N_11532,N_14806);
and U15862 (N_15862,N_10172,N_12667);
nand U15863 (N_15863,N_12926,N_14535);
or U15864 (N_15864,N_11555,N_11245);
and U15865 (N_15865,N_12631,N_12534);
or U15866 (N_15866,N_11546,N_14812);
nand U15867 (N_15867,N_14407,N_11500);
or U15868 (N_15868,N_11636,N_11697);
xor U15869 (N_15869,N_10197,N_10579);
nor U15870 (N_15870,N_14462,N_10203);
xor U15871 (N_15871,N_12989,N_11854);
nand U15872 (N_15872,N_10611,N_12806);
nor U15873 (N_15873,N_12672,N_12278);
nor U15874 (N_15874,N_12760,N_14815);
xor U15875 (N_15875,N_12000,N_14119);
or U15876 (N_15876,N_11393,N_12972);
nor U15877 (N_15877,N_11111,N_13262);
and U15878 (N_15878,N_14302,N_12921);
nor U15879 (N_15879,N_10792,N_10604);
nor U15880 (N_15880,N_11129,N_12161);
xnor U15881 (N_15881,N_10959,N_13069);
nor U15882 (N_15882,N_11067,N_14978);
and U15883 (N_15883,N_11739,N_10020);
and U15884 (N_15884,N_10706,N_11514);
and U15885 (N_15885,N_11119,N_12352);
or U15886 (N_15886,N_14101,N_11761);
or U15887 (N_15887,N_11054,N_12259);
nor U15888 (N_15888,N_14176,N_11892);
xnor U15889 (N_15889,N_14784,N_13327);
nand U15890 (N_15890,N_10305,N_11023);
nand U15891 (N_15891,N_14341,N_14710);
nand U15892 (N_15892,N_11862,N_12639);
nand U15893 (N_15893,N_10379,N_13526);
and U15894 (N_15894,N_14807,N_10864);
or U15895 (N_15895,N_12965,N_13571);
or U15896 (N_15896,N_11598,N_13342);
nand U15897 (N_15897,N_10740,N_14836);
or U15898 (N_15898,N_13659,N_14151);
nor U15899 (N_15899,N_12295,N_12944);
or U15900 (N_15900,N_14680,N_13541);
and U15901 (N_15901,N_12930,N_14873);
nor U15902 (N_15902,N_12796,N_10308);
nor U15903 (N_15903,N_14754,N_13254);
nor U15904 (N_15904,N_14301,N_12447);
and U15905 (N_15905,N_11168,N_10474);
or U15906 (N_15906,N_12784,N_12346);
and U15907 (N_15907,N_12218,N_12091);
and U15908 (N_15908,N_13554,N_10599);
or U15909 (N_15909,N_10053,N_13193);
and U15910 (N_15910,N_10613,N_13739);
nor U15911 (N_15911,N_12906,N_11305);
or U15912 (N_15912,N_10762,N_14298);
and U15913 (N_15913,N_14850,N_10782);
nand U15914 (N_15914,N_12362,N_10741);
or U15915 (N_15915,N_12386,N_14768);
or U15916 (N_15916,N_10179,N_10422);
nand U15917 (N_15917,N_13361,N_12427);
and U15918 (N_15918,N_10092,N_11580);
and U15919 (N_15919,N_10577,N_10268);
and U15920 (N_15920,N_10685,N_12168);
or U15921 (N_15921,N_10301,N_14705);
nor U15922 (N_15922,N_10019,N_11814);
and U15923 (N_15923,N_10257,N_13932);
and U15924 (N_15924,N_11074,N_14382);
and U15925 (N_15925,N_12552,N_10074);
nor U15926 (N_15926,N_11350,N_12722);
and U15927 (N_15927,N_10633,N_11142);
and U15928 (N_15928,N_10232,N_14132);
and U15929 (N_15929,N_13584,N_13875);
nand U15930 (N_15930,N_14926,N_10206);
nor U15931 (N_15931,N_13267,N_10159);
or U15932 (N_15932,N_14441,N_11618);
and U15933 (N_15933,N_13398,N_10817);
or U15934 (N_15934,N_13654,N_14363);
nand U15935 (N_15935,N_13962,N_13587);
nand U15936 (N_15936,N_14315,N_11712);
or U15937 (N_15937,N_14035,N_13149);
nand U15938 (N_15938,N_11210,N_14820);
nor U15939 (N_15939,N_13914,N_12472);
and U15940 (N_15940,N_10772,N_14337);
nor U15941 (N_15941,N_11264,N_13424);
nor U15942 (N_15942,N_12860,N_13673);
or U15943 (N_15943,N_10112,N_11420);
or U15944 (N_15944,N_11508,N_13482);
nor U15945 (N_15945,N_11820,N_14007);
or U15946 (N_15946,N_14716,N_13228);
nor U15947 (N_15947,N_13764,N_14888);
nand U15948 (N_15948,N_14793,N_13757);
nand U15949 (N_15949,N_11860,N_13500);
nand U15950 (N_15950,N_10408,N_10935);
nand U15951 (N_15951,N_14308,N_14202);
nor U15952 (N_15952,N_14938,N_11206);
or U15953 (N_15953,N_14855,N_12565);
nor U15954 (N_15954,N_13820,N_14434);
or U15955 (N_15955,N_13716,N_10587);
or U15956 (N_15956,N_13367,N_14555);
nor U15957 (N_15957,N_13745,N_11004);
xnor U15958 (N_15958,N_13511,N_12768);
and U15959 (N_15959,N_11632,N_12679);
nand U15960 (N_15960,N_14124,N_11935);
and U15961 (N_15961,N_14447,N_13387);
or U15962 (N_15962,N_13957,N_14859);
xnor U15963 (N_15963,N_12466,N_14170);
and U15964 (N_15964,N_13002,N_14640);
or U15965 (N_15965,N_10649,N_12662);
and U15966 (N_15966,N_11256,N_13401);
and U15967 (N_15967,N_14802,N_10026);
nand U15968 (N_15968,N_14998,N_11040);
and U15969 (N_15969,N_10760,N_11554);
nand U15970 (N_15970,N_12729,N_14915);
nor U15971 (N_15971,N_11884,N_12310);
and U15972 (N_15972,N_12012,N_10364);
nand U15973 (N_15973,N_11901,N_12430);
xor U15974 (N_15974,N_12747,N_12297);
nor U15975 (N_15975,N_11321,N_11767);
and U15976 (N_15976,N_14801,N_14299);
nor U15977 (N_15977,N_13359,N_11595);
or U15978 (N_15978,N_14569,N_13953);
xor U15979 (N_15979,N_10323,N_14161);
nor U15980 (N_15980,N_11668,N_12282);
nor U15981 (N_15981,N_10277,N_14550);
or U15982 (N_15982,N_12234,N_13178);
nor U15983 (N_15983,N_13896,N_14732);
nand U15984 (N_15984,N_11802,N_14800);
nor U15985 (N_15985,N_10731,N_11090);
nor U15986 (N_15986,N_12442,N_12850);
nand U15987 (N_15987,N_12312,N_12211);
nor U15988 (N_15988,N_10150,N_14127);
or U15989 (N_15989,N_11848,N_14030);
and U15990 (N_15990,N_11267,N_10943);
and U15991 (N_15991,N_12141,N_12745);
nor U15992 (N_15992,N_11276,N_13095);
or U15993 (N_15993,N_12814,N_13062);
xnor U15994 (N_15994,N_13606,N_12649);
nor U15995 (N_15995,N_12480,N_14439);
xnor U15996 (N_15996,N_11978,N_12537);
nand U15997 (N_15997,N_13799,N_14473);
xnor U15998 (N_15998,N_12996,N_11975);
nand U15999 (N_15999,N_12101,N_10022);
and U16000 (N_16000,N_14449,N_10550);
or U16001 (N_16001,N_11394,N_11278);
nand U16002 (N_16002,N_14385,N_11165);
nand U16003 (N_16003,N_11167,N_14050);
xor U16004 (N_16004,N_11118,N_10034);
nand U16005 (N_16005,N_10752,N_13183);
or U16006 (N_16006,N_10561,N_14919);
and U16007 (N_16007,N_14971,N_14796);
or U16008 (N_16008,N_12154,N_14516);
nand U16009 (N_16009,N_11038,N_12420);
and U16010 (N_16010,N_12450,N_14225);
nor U16011 (N_16011,N_14319,N_12028);
or U16012 (N_16012,N_11468,N_13698);
or U16013 (N_16013,N_13390,N_11121);
nand U16014 (N_16014,N_13822,N_11987);
or U16015 (N_16015,N_11841,N_12797);
nand U16016 (N_16016,N_13098,N_11105);
nand U16017 (N_16017,N_11406,N_11166);
and U16018 (N_16018,N_11783,N_11055);
and U16019 (N_16019,N_12222,N_13406);
nand U16020 (N_16020,N_10435,N_11913);
nor U16021 (N_16021,N_13665,N_11408);
and U16022 (N_16022,N_11316,N_11812);
or U16023 (N_16023,N_14239,N_13690);
xnor U16024 (N_16024,N_10326,N_14153);
xor U16025 (N_16025,N_14205,N_12752);
nand U16026 (N_16026,N_10902,N_11261);
nor U16027 (N_16027,N_12890,N_10096);
nand U16028 (N_16028,N_14513,N_10900);
nand U16029 (N_16029,N_10896,N_11359);
or U16030 (N_16030,N_13202,N_10339);
nand U16031 (N_16031,N_10874,N_14568);
nor U16032 (N_16032,N_14125,N_13369);
and U16033 (N_16033,N_12726,N_10249);
and U16034 (N_16034,N_13418,N_11698);
and U16035 (N_16035,N_13339,N_11817);
and U16036 (N_16036,N_13138,N_10048);
xor U16037 (N_16037,N_14359,N_11169);
or U16038 (N_16038,N_14811,N_10696);
or U16039 (N_16039,N_13287,N_12212);
or U16040 (N_16040,N_14879,N_13321);
or U16041 (N_16041,N_13362,N_10811);
xor U16042 (N_16042,N_14626,N_12689);
nor U16043 (N_16043,N_10421,N_10454);
nor U16044 (N_16044,N_14845,N_13783);
nand U16045 (N_16045,N_11912,N_14304);
and U16046 (N_16046,N_10862,N_11564);
nor U16047 (N_16047,N_13465,N_13750);
nand U16048 (N_16048,N_14763,N_13052);
nand U16049 (N_16049,N_13490,N_10925);
and U16050 (N_16050,N_10949,N_11030);
or U16051 (N_16051,N_13944,N_11985);
nor U16052 (N_16052,N_14234,N_13349);
or U16053 (N_16053,N_13243,N_13206);
nand U16054 (N_16054,N_10645,N_12777);
nand U16055 (N_16055,N_14571,N_10125);
nand U16056 (N_16056,N_13761,N_14906);
nand U16057 (N_16057,N_13404,N_14229);
or U16058 (N_16058,N_13473,N_11050);
xor U16059 (N_16059,N_14614,N_12219);
nand U16060 (N_16060,N_10119,N_11686);
or U16061 (N_16061,N_10225,N_13918);
and U16062 (N_16062,N_12244,N_12707);
and U16063 (N_16063,N_12068,N_12074);
nand U16064 (N_16064,N_11509,N_13460);
nand U16065 (N_16065,N_12737,N_11898);
nor U16066 (N_16066,N_11184,N_12643);
or U16067 (N_16067,N_12873,N_12394);
xor U16068 (N_16068,N_11234,N_10929);
nand U16069 (N_16069,N_12931,N_14921);
nand U16070 (N_16070,N_14016,N_11179);
nor U16071 (N_16071,N_10571,N_12131);
and U16072 (N_16072,N_10248,N_13033);
nor U16073 (N_16073,N_14642,N_10294);
nand U16074 (N_16074,N_11382,N_10468);
and U16075 (N_16075,N_11322,N_12184);
nor U16076 (N_16076,N_12616,N_14432);
or U16077 (N_16077,N_12529,N_14199);
xor U16078 (N_16078,N_12673,N_12398);
xor U16079 (N_16079,N_12217,N_10553);
nand U16080 (N_16080,N_13677,N_14219);
and U16081 (N_16081,N_14180,N_13942);
nand U16082 (N_16082,N_14667,N_11674);
or U16083 (N_16083,N_14425,N_12494);
nor U16084 (N_16084,N_13331,N_14637);
xnor U16085 (N_16085,N_12835,N_12355);
nand U16086 (N_16086,N_11388,N_14583);
nor U16087 (N_16087,N_11136,N_14236);
and U16088 (N_16088,N_12422,N_10398);
nand U16089 (N_16089,N_10694,N_11226);
or U16090 (N_16090,N_12964,N_11384);
nor U16091 (N_16091,N_13747,N_11486);
nand U16092 (N_16092,N_10396,N_13227);
nand U16093 (N_16093,N_14922,N_12441);
and U16094 (N_16094,N_11300,N_10775);
or U16095 (N_16095,N_11334,N_13365);
nor U16096 (N_16096,N_14596,N_14918);
nor U16097 (N_16097,N_12146,N_11986);
nand U16098 (N_16098,N_12805,N_14693);
and U16099 (N_16099,N_13005,N_10306);
xnor U16100 (N_16100,N_14240,N_11794);
nand U16101 (N_16101,N_12100,N_11411);
and U16102 (N_16102,N_14480,N_13835);
nor U16103 (N_16103,N_12854,N_10059);
or U16104 (N_16104,N_10458,N_13949);
and U16105 (N_16105,N_11824,N_13368);
and U16106 (N_16106,N_14039,N_13777);
and U16107 (N_16107,N_10517,N_10505);
and U16108 (N_16108,N_10005,N_13725);
xor U16109 (N_16109,N_10987,N_11710);
and U16110 (N_16110,N_14795,N_11552);
nand U16111 (N_16111,N_11711,N_11870);
and U16112 (N_16112,N_11773,N_10160);
nand U16113 (N_16113,N_12711,N_13352);
and U16114 (N_16114,N_11754,N_13924);
nand U16115 (N_16115,N_12773,N_12515);
and U16116 (N_16116,N_12829,N_12408);
nor U16117 (N_16117,N_14409,N_10208);
or U16118 (N_16118,N_13196,N_13044);
xnor U16119 (N_16119,N_14346,N_10442);
nand U16120 (N_16120,N_14064,N_10145);
nand U16121 (N_16121,N_13866,N_13780);
or U16122 (N_16122,N_12799,N_13481);
nand U16123 (N_16123,N_11742,N_14256);
xnor U16124 (N_16124,N_13575,N_13224);
and U16125 (N_16125,N_10190,N_12428);
nor U16126 (N_16126,N_13461,N_14924);
nand U16127 (N_16127,N_11981,N_11380);
and U16128 (N_16128,N_10872,N_12524);
or U16129 (N_16129,N_13570,N_10919);
nor U16130 (N_16130,N_14021,N_11133);
nor U16131 (N_16131,N_11372,N_14350);
nand U16132 (N_16132,N_11005,N_13601);
nor U16133 (N_16133,N_13117,N_12471);
and U16134 (N_16134,N_14874,N_12225);
nor U16135 (N_16135,N_10271,N_11522);
nand U16136 (N_16136,N_14467,N_10317);
and U16137 (N_16137,N_10446,N_11242);
nand U16138 (N_16138,N_13542,N_12132);
or U16139 (N_16139,N_12306,N_11496);
xnor U16140 (N_16140,N_14128,N_12072);
or U16141 (N_16141,N_10479,N_14068);
nor U16142 (N_16142,N_14781,N_12785);
xor U16143 (N_16143,N_12550,N_12775);
or U16144 (N_16144,N_13150,N_12406);
nor U16145 (N_16145,N_12162,N_14111);
and U16146 (N_16146,N_10827,N_11225);
nor U16147 (N_16147,N_14226,N_12728);
and U16148 (N_16148,N_11279,N_12968);
nand U16149 (N_16149,N_14037,N_13188);
and U16150 (N_16150,N_10798,N_11872);
and U16151 (N_16151,N_10108,N_11559);
and U16152 (N_16152,N_12787,N_11156);
nor U16153 (N_16153,N_11343,N_13079);
nand U16154 (N_16154,N_11990,N_13684);
and U16155 (N_16155,N_10536,N_11998);
nand U16156 (N_16156,N_13235,N_10855);
nand U16157 (N_16157,N_11303,N_13778);
or U16158 (N_16158,N_13660,N_13847);
nor U16159 (N_16159,N_10416,N_13035);
nor U16160 (N_16160,N_11183,N_13623);
nand U16161 (N_16161,N_13649,N_10881);
xnor U16162 (N_16162,N_10947,N_10450);
and U16163 (N_16163,N_10175,N_14279);
nand U16164 (N_16164,N_14141,N_12889);
and U16165 (N_16165,N_12376,N_13425);
nand U16166 (N_16166,N_12539,N_14738);
or U16167 (N_16167,N_10065,N_12354);
and U16168 (N_16168,N_14201,N_14493);
xor U16169 (N_16169,N_10194,N_14461);
and U16170 (N_16170,N_13657,N_13900);
xnor U16171 (N_16171,N_12644,N_14494);
or U16172 (N_16172,N_11553,N_12369);
nand U16173 (N_16173,N_10735,N_11882);
and U16174 (N_16174,N_11107,N_12124);
or U16175 (N_16175,N_13779,N_13237);
and U16176 (N_16176,N_11780,N_12702);
xnor U16177 (N_16177,N_13902,N_14917);
or U16178 (N_16178,N_13696,N_10351);
or U16179 (N_16179,N_14548,N_11888);
nand U16180 (N_16180,N_14936,N_11705);
or U16181 (N_16181,N_14632,N_12698);
nand U16182 (N_16182,N_12872,N_13126);
nand U16183 (N_16183,N_10218,N_11254);
xor U16184 (N_16184,N_10860,N_11845);
or U16185 (N_16185,N_10522,N_13096);
and U16186 (N_16186,N_12058,N_13860);
and U16187 (N_16187,N_12434,N_12267);
and U16188 (N_16188,N_10582,N_13700);
or U16189 (N_16189,N_11066,N_13251);
nor U16190 (N_16190,N_14329,N_12810);
or U16191 (N_16191,N_13325,N_13981);
nor U16192 (N_16192,N_11020,N_14062);
xnor U16193 (N_16193,N_10118,N_13422);
nor U16194 (N_16194,N_10002,N_14034);
or U16195 (N_16195,N_11329,N_10184);
nand U16196 (N_16196,N_12574,N_10055);
nand U16197 (N_16197,N_10148,N_10341);
and U16198 (N_16198,N_10682,N_14175);
nand U16199 (N_16199,N_10013,N_14521);
nand U16200 (N_16200,N_11819,N_10402);
or U16201 (N_16201,N_11640,N_10915);
and U16202 (N_16202,N_14589,N_12741);
nor U16203 (N_16203,N_10461,N_13030);
or U16204 (N_16204,N_13909,N_12721);
and U16205 (N_16205,N_10851,N_10918);
or U16206 (N_16206,N_14103,N_12029);
and U16207 (N_16207,N_12716,N_14203);
nor U16208 (N_16208,N_14902,N_10285);
nor U16209 (N_16209,N_10136,N_10646);
and U16210 (N_16210,N_13305,N_13737);
nand U16211 (N_16211,N_11511,N_11087);
and U16212 (N_16212,N_11928,N_13277);
nor U16213 (N_16213,N_12668,N_13283);
or U16214 (N_16214,N_11070,N_13648);
and U16215 (N_16215,N_14747,N_12286);
nor U16216 (N_16216,N_12435,N_12367);
nand U16217 (N_16217,N_10420,N_10726);
nor U16218 (N_16218,N_14472,N_10502);
xnor U16219 (N_16219,N_12942,N_11001);
xnor U16220 (N_16220,N_11215,N_13216);
nor U16221 (N_16221,N_14525,N_10071);
or U16222 (N_16222,N_12924,N_10290);
and U16223 (N_16223,N_14627,N_13497);
nand U16224 (N_16224,N_14116,N_14551);
or U16225 (N_16225,N_13205,N_14411);
and U16226 (N_16226,N_14275,N_14541);
nand U16227 (N_16227,N_12868,N_10532);
nor U16228 (N_16228,N_12319,N_12762);
nor U16229 (N_16229,N_10045,N_11460);
xnor U16230 (N_16230,N_10128,N_12477);
and U16231 (N_16231,N_13888,N_12542);
xor U16232 (N_16232,N_13443,N_10773);
or U16233 (N_16233,N_14258,N_14968);
xnor U16234 (N_16234,N_14810,N_14244);
nand U16235 (N_16235,N_10081,N_14281);
nor U16236 (N_16236,N_13376,N_11796);
nor U16237 (N_16237,N_10064,N_13797);
and U16238 (N_16238,N_13032,N_11926);
xor U16239 (N_16239,N_14973,N_13199);
nor U16240 (N_16240,N_10799,N_13741);
and U16241 (N_16241,N_14038,N_13212);
xnor U16242 (N_16242,N_10397,N_13343);
nor U16243 (N_16243,N_12429,N_10758);
or U16244 (N_16244,N_11753,N_13088);
or U16245 (N_16245,N_10606,N_10841);
nand U16246 (N_16246,N_10332,N_11347);
nor U16247 (N_16247,N_13015,N_12241);
nand U16248 (N_16248,N_11718,N_10392);
or U16249 (N_16249,N_13970,N_10853);
or U16250 (N_16250,N_14019,N_10785);
and U16251 (N_16251,N_12817,N_13950);
and U16252 (N_16252,N_11079,N_12730);
and U16253 (N_16253,N_13363,N_10319);
nand U16254 (N_16254,N_14829,N_12412);
nand U16255 (N_16255,N_12738,N_14696);
and U16256 (N_16256,N_12065,N_11052);
nor U16257 (N_16257,N_10648,N_10330);
nor U16258 (N_16258,N_14470,N_12652);
nand U16259 (N_16259,N_10678,N_11631);
or U16260 (N_16260,N_13758,N_14574);
and U16261 (N_16261,N_14941,N_10472);
and U16262 (N_16262,N_13155,N_11826);
nor U16263 (N_16263,N_11852,N_13089);
or U16264 (N_16264,N_12118,N_10490);
nor U16265 (N_16265,N_11374,N_10596);
or U16266 (N_16266,N_13508,N_10945);
nand U16267 (N_16267,N_12324,N_13057);
and U16268 (N_16268,N_11517,N_10324);
nor U16269 (N_16269,N_10139,N_11603);
nor U16270 (N_16270,N_10028,N_14332);
or U16271 (N_16271,N_11423,N_11809);
nand U16272 (N_16272,N_10487,N_11154);
and U16273 (N_16273,N_11110,N_11937);
or U16274 (N_16274,N_12437,N_12758);
nor U16275 (N_16275,N_14851,N_14530);
or U16276 (N_16276,N_10545,N_10187);
and U16277 (N_16277,N_11972,N_12022);
or U16278 (N_16278,N_13531,N_11258);
or U16279 (N_16279,N_13553,N_12659);
nand U16280 (N_16280,N_11561,N_12580);
xor U16281 (N_16281,N_14959,N_12066);
or U16282 (N_16282,N_14045,N_13796);
nor U16283 (N_16283,N_12481,N_13081);
nand U16284 (N_16284,N_14607,N_11678);
or U16285 (N_16285,N_12967,N_13232);
and U16286 (N_16286,N_11059,N_14378);
and U16287 (N_16287,N_14032,N_10910);
and U16288 (N_16288,N_10494,N_11681);
nor U16289 (N_16289,N_10675,N_10806);
or U16290 (N_16290,N_10480,N_11439);
or U16291 (N_16291,N_11964,N_12782);
nor U16292 (N_16292,N_11856,N_14009);
and U16293 (N_16293,N_11722,N_11203);
or U16294 (N_16294,N_14102,N_12169);
or U16295 (N_16295,N_14897,N_13185);
or U16296 (N_16296,N_11407,N_14117);
and U16297 (N_16297,N_14197,N_10137);
nand U16298 (N_16298,N_12034,N_10174);
nand U16299 (N_16299,N_10141,N_11227);
xor U16300 (N_16300,N_11973,N_12082);
nand U16301 (N_16301,N_11060,N_13230);
or U16302 (N_16302,N_10110,N_10483);
xnor U16303 (N_16303,N_14356,N_14297);
or U16304 (N_16304,N_10936,N_10459);
and U16305 (N_16305,N_12718,N_12393);
nand U16306 (N_16306,N_11039,N_13301);
or U16307 (N_16307,N_11630,N_11866);
xor U16308 (N_16308,N_10715,N_14623);
and U16309 (N_16309,N_11244,N_14989);
and U16310 (N_16310,N_10516,N_13709);
and U16311 (N_16311,N_10870,N_13259);
and U16312 (N_16312,N_12848,N_11268);
and U16313 (N_16313,N_10430,N_12851);
nand U16314 (N_16314,N_13712,N_13008);
or U16315 (N_16315,N_10135,N_12864);
nor U16316 (N_16316,N_14579,N_12677);
nor U16317 (N_16317,N_11116,N_13061);
nor U16318 (N_16318,N_12792,N_13768);
or U16319 (N_16319,N_11877,N_13523);
nor U16320 (N_16320,N_10511,N_10032);
nor U16321 (N_16321,N_12257,N_10535);
and U16322 (N_16322,N_14858,N_12575);
nand U16323 (N_16323,N_10431,N_12311);
nor U16324 (N_16324,N_14322,N_10628);
or U16325 (N_16325,N_12252,N_10630);
and U16326 (N_16326,N_10658,N_13085);
xnor U16327 (N_16327,N_14410,N_12628);
nor U16328 (N_16328,N_14187,N_14005);
nand U16329 (N_16329,N_14259,N_12774);
nor U16330 (N_16330,N_12227,N_10813);
nand U16331 (N_16331,N_10875,N_13833);
nor U16332 (N_16332,N_12030,N_13652);
and U16333 (N_16333,N_13776,N_14367);
and U16334 (N_16334,N_13890,N_14211);
or U16335 (N_16335,N_10679,N_10017);
nand U16336 (N_16336,N_10043,N_11104);
or U16337 (N_16337,N_12879,N_13270);
or U16338 (N_16338,N_10103,N_11805);
or U16339 (N_16339,N_14647,N_14932);
and U16340 (N_16340,N_12134,N_12454);
nand U16341 (N_16341,N_14216,N_11516);
nor U16342 (N_16342,N_14894,N_12602);
nand U16343 (N_16343,N_10327,N_11955);
or U16344 (N_16344,N_12900,N_13092);
nor U16345 (N_16345,N_10882,N_12691);
xnor U16346 (N_16346,N_11741,N_10725);
xor U16347 (N_16347,N_13543,N_13333);
or U16348 (N_16348,N_14208,N_10289);
nor U16349 (N_16349,N_11828,N_14707);
nand U16350 (N_16350,N_11295,N_13730);
nand U16351 (N_16351,N_12981,N_13201);
and U16352 (N_16352,N_10204,N_13194);
nor U16353 (N_16353,N_11337,N_11170);
nand U16354 (N_16354,N_10133,N_11617);
nor U16355 (N_16355,N_14970,N_10567);
nand U16356 (N_16356,N_13600,N_12641);
nor U16357 (N_16357,N_11495,N_14676);
or U16358 (N_16358,N_10634,N_10990);
nand U16359 (N_16359,N_12127,N_14133);
and U16360 (N_16360,N_13885,N_10292);
nand U16361 (N_16361,N_13582,N_12418);
or U16362 (N_16362,N_12650,N_13701);
or U16363 (N_16363,N_13423,N_10858);
or U16364 (N_16364,N_10355,N_13751);
or U16365 (N_16365,N_10113,N_10722);
nor U16366 (N_16366,N_14287,N_12025);
and U16367 (N_16367,N_10077,N_11352);
nor U16368 (N_16368,N_13615,N_10451);
and U16369 (N_16369,N_12674,N_12316);
nand U16370 (N_16370,N_11349,N_14188);
and U16371 (N_16371,N_11454,N_11291);
nor U16372 (N_16372,N_14088,N_10721);
nor U16373 (N_16373,N_14455,N_13100);
xnor U16374 (N_16374,N_11094,N_14669);
nand U16375 (N_16375,N_14278,N_13877);
and U16376 (N_16376,N_11470,N_12586);
nor U16377 (N_16377,N_11164,N_14787);
or U16378 (N_16378,N_12648,N_10779);
or U16379 (N_16379,N_12114,N_13556);
and U16380 (N_16380,N_13348,N_10923);
or U16381 (N_16381,N_14603,N_12463);
nor U16382 (N_16382,N_11946,N_12767);
or U16383 (N_16383,N_13437,N_13159);
or U16384 (N_16384,N_10993,N_10575);
and U16385 (N_16385,N_13718,N_12359);
nand U16386 (N_16386,N_13459,N_12045);
or U16387 (N_16387,N_14469,N_10117);
nor U16388 (N_16388,N_10979,N_13364);
or U16389 (N_16389,N_12941,N_11150);
and U16390 (N_16390,N_14029,N_13495);
or U16391 (N_16391,N_10245,N_13116);
xnor U16392 (N_16392,N_10100,N_11642);
or U16393 (N_16393,N_13544,N_14757);
and U16394 (N_16394,N_14846,N_11416);
and U16395 (N_16395,N_14091,N_11426);
and U16396 (N_16396,N_12130,N_14914);
and U16397 (N_16397,N_12527,N_14075);
and U16398 (N_16398,N_12214,N_11478);
nand U16399 (N_16399,N_10742,N_12077);
and U16400 (N_16400,N_10278,N_10695);
and U16401 (N_16401,N_11013,N_11159);
and U16402 (N_16402,N_11444,N_14826);
nor U16403 (N_16403,N_10033,N_12815);
and U16404 (N_16404,N_11045,N_13530);
or U16405 (N_16405,N_14386,N_11801);
or U16406 (N_16406,N_11229,N_12834);
and U16407 (N_16407,N_12461,N_10623);
or U16408 (N_16408,N_12108,N_10142);
nor U16409 (N_16409,N_12176,N_14694);
and U16410 (N_16410,N_10205,N_14636);
nand U16411 (N_16411,N_11715,N_11081);
xor U16412 (N_16412,N_10012,N_10974);
and U16413 (N_16413,N_10795,N_11474);
nand U16414 (N_16414,N_14877,N_13078);
nand U16415 (N_16415,N_14698,N_11699);
and U16416 (N_16416,N_10668,N_14752);
nor U16417 (N_16417,N_12115,N_14147);
nor U16418 (N_16418,N_11222,N_10850);
and U16419 (N_16419,N_14939,N_11479);
and U16420 (N_16420,N_13955,N_11185);
and U16421 (N_16421,N_12531,N_10796);
nand U16422 (N_16422,N_12017,N_12110);
and U16423 (N_16423,N_14486,N_13975);
nand U16424 (N_16424,N_10036,N_14528);
nor U16425 (N_16425,N_10964,N_13355);
xor U16426 (N_16426,N_10140,N_12736);
and U16427 (N_16427,N_14106,N_14368);
nand U16428 (N_16428,N_10122,N_10444);
or U16429 (N_16429,N_11965,N_11383);
or U16430 (N_16430,N_12863,N_14862);
nand U16431 (N_16431,N_14450,N_11988);
and U16432 (N_16432,N_13041,N_11563);
nor U16433 (N_16433,N_13619,N_12438);
nor U16434 (N_16434,N_14869,N_13713);
or U16435 (N_16435,N_13051,N_13706);
nor U16436 (N_16436,N_12183,N_14290);
nand U16437 (N_16437,N_13539,N_12417);
nand U16438 (N_16438,N_13923,N_14786);
nor U16439 (N_16439,N_12468,N_10328);
nor U16440 (N_16440,N_13105,N_12232);
nand U16441 (N_16441,N_13598,N_11865);
or U16442 (N_16442,N_10448,N_11774);
nand U16443 (N_16443,N_14295,N_12878);
nand U16444 (N_16444,N_10404,N_13160);
nand U16445 (N_16445,N_12054,N_13893);
xor U16446 (N_16446,N_13023,N_13976);
or U16447 (N_16447,N_12188,N_11766);
and U16448 (N_16448,N_11840,N_13618);
nor U16449 (N_16449,N_10104,N_14782);
nor U16450 (N_16450,N_10988,N_11088);
or U16451 (N_16451,N_12802,N_11945);
or U16452 (N_16452,N_12419,N_12630);
and U16453 (N_16453,N_10079,N_13389);
and U16454 (N_16454,N_11692,N_12603);
nand U16455 (N_16455,N_13749,N_14008);
nand U16456 (N_16456,N_13506,N_11328);
or U16457 (N_16457,N_14523,N_13852);
nand U16458 (N_16458,N_11579,N_10744);
nand U16459 (N_16459,N_14951,N_13973);
nor U16460 (N_16460,N_14324,N_12198);
and U16461 (N_16461,N_11425,N_13859);
xor U16462 (N_16462,N_14870,N_14272);
or U16463 (N_16463,N_12308,N_12843);
and U16464 (N_16464,N_13197,N_14739);
or U16465 (N_16465,N_13917,N_10475);
nor U16466 (N_16466,N_10781,N_14044);
and U16467 (N_16467,N_13517,N_11296);
xnor U16468 (N_16468,N_11077,N_10523);
nand U16469 (N_16469,N_10393,N_10508);
nor U16470 (N_16470,N_12581,N_14282);
nor U16471 (N_16471,N_10794,N_13760);
or U16472 (N_16472,N_12923,N_12400);
nor U16473 (N_16473,N_13756,N_12520);
and U16474 (N_16474,N_11108,N_11421);
nand U16475 (N_16475,N_10383,N_10672);
and U16476 (N_16476,N_10309,N_14246);
nor U16477 (N_16477,N_14099,N_10880);
xor U16478 (N_16478,N_14115,N_10255);
or U16479 (N_16479,N_13211,N_12746);
nor U16480 (N_16480,N_11948,N_10415);
xor U16481 (N_16481,N_14171,N_12377);
or U16482 (N_16482,N_11323,N_14416);
xor U16483 (N_16483,N_12104,N_14560);
nor U16484 (N_16484,N_14071,N_12608);
and U16485 (N_16485,N_12155,N_11825);
nand U16486 (N_16486,N_13831,N_12208);
xor U16487 (N_16487,N_11915,N_10075);
or U16488 (N_16488,N_12084,N_13842);
or U16489 (N_16489,N_12597,N_12522);
xor U16490 (N_16490,N_14043,N_12464);
nand U16491 (N_16491,N_13524,N_13353);
and U16492 (N_16492,N_13532,N_10004);
nor U16493 (N_16493,N_14031,N_11312);
and U16494 (N_16494,N_14908,N_14000);
xnor U16495 (N_16495,N_12939,N_12845);
nand U16496 (N_16496,N_11288,N_12626);
or U16497 (N_16497,N_13527,N_12062);
xor U16498 (N_16498,N_10109,N_14708);
nand U16499 (N_16499,N_14495,N_12636);
nand U16500 (N_16500,N_12079,N_10346);
nand U16501 (N_16501,N_10520,N_13171);
nand U16502 (N_16502,N_12439,N_11202);
nand U16503 (N_16503,N_11790,N_13351);
xnor U16504 (N_16504,N_10496,N_14430);
nand U16505 (N_16505,N_12510,N_13865);
nand U16506 (N_16506,N_11764,N_10662);
or U16507 (N_16507,N_12224,N_11356);
nor U16508 (N_16508,N_11851,N_13431);
or U16509 (N_16509,N_12517,N_13558);
nand U16510 (N_16510,N_11943,N_14122);
or U16511 (N_16511,N_14262,N_13136);
or U16512 (N_16512,N_10897,N_11658);
or U16513 (N_16513,N_11095,N_10050);
and U16514 (N_16514,N_12961,N_11148);
or U16515 (N_16515,N_13241,N_14661);
nand U16516 (N_16516,N_12476,N_12856);
nor U16517 (N_16517,N_10965,N_13427);
and U16518 (N_16518,N_13814,N_10481);
or U16519 (N_16519,N_10538,N_14087);
nand U16520 (N_16520,N_10519,N_12696);
xor U16521 (N_16521,N_12625,N_10548);
nor U16522 (N_16522,N_10467,N_14519);
or U16523 (N_16523,N_13135,N_12594);
or U16524 (N_16524,N_13731,N_13114);
and U16525 (N_16525,N_10329,N_13680);
nor U16526 (N_16526,N_10921,N_11811);
nand U16527 (N_16527,N_10992,N_12886);
or U16528 (N_16528,N_14798,N_10911);
or U16529 (N_16529,N_12325,N_11436);
nor U16530 (N_16530,N_13821,N_14092);
and U16531 (N_16531,N_14580,N_14893);
xnor U16532 (N_16532,N_11557,N_14232);
xor U16533 (N_16533,N_14654,N_11143);
or U16534 (N_16534,N_12363,N_11015);
and U16535 (N_16535,N_10999,N_12165);
or U16536 (N_16536,N_14835,N_12950);
and U16537 (N_16537,N_12938,N_12891);
or U16538 (N_16538,N_13410,N_10124);
nand U16539 (N_16539,N_10044,N_10933);
and U16540 (N_16540,N_10984,N_13549);
or U16541 (N_16541,N_11689,N_11082);
xor U16542 (N_16542,N_14881,N_11894);
or U16543 (N_16543,N_11057,N_10543);
nand U16544 (N_16544,N_13631,N_11122);
xor U16545 (N_16545,N_10552,N_12994);
or U16546 (N_16546,N_13664,N_13994);
or U16547 (N_16547,N_11283,N_11639);
and U16548 (N_16548,N_14181,N_13001);
xnor U16549 (N_16549,N_12345,N_14429);
or U16550 (N_16550,N_14709,N_10549);
nor U16551 (N_16551,N_12063,N_13800);
and U16552 (N_16552,N_10035,N_12090);
nand U16553 (N_16553,N_14741,N_10767);
or U16554 (N_16554,N_14126,N_10728);
or U16555 (N_16555,N_11314,N_12451);
nor U16556 (N_16556,N_13246,N_13472);
nand U16557 (N_16557,N_14746,N_12307);
and U16558 (N_16558,N_11093,N_14463);
or U16559 (N_16559,N_13851,N_13638);
or U16560 (N_16560,N_10805,N_13572);
nand U16561 (N_16561,N_10867,N_12357);
and U16562 (N_16562,N_14026,N_14649);
xnor U16563 (N_16563,N_10754,N_11938);
or U16564 (N_16564,N_14481,N_11114);
and U16565 (N_16565,N_13027,N_11263);
and U16566 (N_16566,N_12937,N_11302);
or U16567 (N_16567,N_11779,N_13608);
nand U16568 (N_16568,N_12409,N_10154);
nand U16569 (N_16569,N_12174,N_10565);
nand U16570 (N_16570,N_11016,N_14991);
or U16571 (N_16571,N_14737,N_10414);
or U16572 (N_16572,N_13946,N_10343);
nor U16573 (N_16573,N_11102,N_11921);
and U16574 (N_16574,N_13811,N_14920);
or U16575 (N_16575,N_11301,N_13643);
and U16576 (N_16576,N_14060,N_11743);
and U16577 (N_16577,N_14909,N_14018);
nor U16578 (N_16578,N_12126,N_11190);
nand U16579 (N_16579,N_13104,N_11967);
nand U16580 (N_16580,N_13971,N_10887);
nor U16581 (N_16581,N_14621,N_12769);
or U16582 (N_16582,N_12943,N_12080);
and U16583 (N_16583,N_13391,N_12809);
nor U16584 (N_16584,N_13060,N_11230);
nor U16585 (N_16585,N_10839,N_10510);
nor U16586 (N_16586,N_14392,N_10409);
or U16587 (N_16587,N_13284,N_12426);
and U16588 (N_16588,N_12902,N_10264);
nand U16589 (N_16589,N_14545,N_11189);
nand U16590 (N_16590,N_10217,N_13766);
nand U16591 (N_16591,N_13064,N_13029);
nand U16592 (N_16592,N_13112,N_14327);
nor U16593 (N_16593,N_10922,N_13931);
nand U16594 (N_16594,N_12329,N_13793);
nor U16595 (N_16595,N_12414,N_14509);
xnor U16596 (N_16596,N_13134,N_14638);
or U16597 (N_16597,N_14742,N_13356);
and U16598 (N_16598,N_13629,N_12776);
and U16599 (N_16599,N_11573,N_14436);
nor U16600 (N_16600,N_10857,N_11584);
nor U16601 (N_16601,N_14983,N_14288);
and U16602 (N_16602,N_10749,N_10924);
nand U16603 (N_16603,N_11735,N_13845);
xnor U16604 (N_16604,N_12001,N_12021);
and U16605 (N_16605,N_11014,N_11085);
nand U16606 (N_16606,N_12496,N_14885);
xor U16607 (N_16607,N_13248,N_14475);
nand U16608 (N_16608,N_10810,N_11485);
nor U16609 (N_16609,N_14777,N_14089);
nor U16610 (N_16610,N_14736,N_12291);
nor U16611 (N_16611,N_11428,N_12633);
nor U16612 (N_16612,N_12619,N_11593);
xnor U16613 (N_16613,N_14107,N_11594);
or U16614 (N_16614,N_13512,N_11191);
nand U16615 (N_16615,N_12266,N_12254);
or U16616 (N_16616,N_12133,N_14678);
nor U16617 (N_16617,N_11007,N_14701);
or U16618 (N_16618,N_13479,N_11995);
nor U16619 (N_16619,N_11599,N_13568);
nor U16620 (N_16620,N_13344,N_12719);
nand U16621 (N_16621,N_12920,N_14785);
nor U16622 (N_16622,N_11652,N_11130);
or U16623 (N_16623,N_14144,N_11560);
and U16624 (N_16624,N_10350,N_13711);
and U16625 (N_16625,N_13874,N_13843);
or U16626 (N_16626,N_14994,N_10106);
or U16627 (N_16627,N_11049,N_12033);
and U16628 (N_16628,N_13717,N_12465);
or U16629 (N_16629,N_14652,N_13982);
and U16630 (N_16630,N_11018,N_11002);
nand U16631 (N_16631,N_12251,N_11413);
xnor U16632 (N_16632,N_13165,N_12778);
nand U16633 (N_16633,N_14156,N_14066);
xor U16634 (N_16634,N_13614,N_14587);
nand U16635 (N_16635,N_14562,N_11449);
and U16636 (N_16636,N_14857,N_11448);
and U16637 (N_16637,N_14235,N_11693);
nor U16638 (N_16638,N_10082,N_11760);
nand U16639 (N_16639,N_11782,N_12365);
nand U16640 (N_16640,N_12051,N_12473);
nor U16641 (N_16641,N_13122,N_10447);
nor U16642 (N_16642,N_14999,N_14261);
or U16643 (N_16643,N_10173,N_12765);
xor U16644 (N_16644,N_13039,N_10030);
nor U16645 (N_16645,N_12356,N_11155);
nand U16646 (N_16646,N_10176,N_10826);
and U16647 (N_16647,N_11570,N_14036);
nand U16648 (N_16648,N_10866,N_12343);
and U16649 (N_16649,N_14340,N_11389);
and U16650 (N_16650,N_13784,N_10143);
nor U16651 (N_16651,N_11223,N_11497);
xnor U16652 (N_16652,N_14606,N_13222);
nand U16653 (N_16653,N_11365,N_14761);
nand U16654 (N_16654,N_12678,N_13451);
and U16655 (N_16655,N_10540,N_14377);
xnor U16656 (N_16656,N_10072,N_11233);
nor U16657 (N_16657,N_12285,N_14834);
nand U16658 (N_16658,N_10054,N_11430);
and U16659 (N_16659,N_13108,N_13130);
nand U16660 (N_16660,N_13798,N_11875);
or U16661 (N_16661,N_11209,N_13499);
nand U16662 (N_16662,N_10597,N_14207);
and U16663 (N_16663,N_14554,N_10495);
nand U16664 (N_16664,N_13070,N_13827);
nor U16665 (N_16665,N_10801,N_14433);
nand U16666 (N_16666,N_11740,N_13678);
or U16667 (N_16667,N_13621,N_14890);
nor U16668 (N_16668,N_10639,N_12828);
nor U16669 (N_16669,N_11628,N_10914);
and U16670 (N_16670,N_13458,N_14619);
xor U16671 (N_16671,N_14248,N_13090);
nor U16672 (N_16672,N_10605,N_12970);
nand U16673 (N_16673,N_12882,N_13689);
nand U16674 (N_16674,N_13123,N_13938);
and U16675 (N_16675,N_11253,N_11124);
nor U16676 (N_16676,N_13300,N_11009);
nor U16677 (N_16677,N_12870,N_11306);
nor U16678 (N_16678,N_13612,N_14335);
xor U16679 (N_16679,N_13873,N_11519);
and U16680 (N_16680,N_13590,N_13026);
and U16681 (N_16681,N_14085,N_12826);
or U16682 (N_16682,N_13682,N_10313);
nand U16683 (N_16683,N_13993,N_11850);
or U16684 (N_16684,N_10201,N_14730);
and U16685 (N_16685,N_11979,N_10653);
nand U16686 (N_16686,N_14140,N_14517);
nand U16687 (N_16687,N_12487,N_13261);
nor U16688 (N_16688,N_11083,N_10971);
nor U16689 (N_16689,N_10237,N_11752);
nand U16690 (N_16690,N_14896,N_12687);
or U16691 (N_16691,N_12577,N_11798);
and U16692 (N_16692,N_12862,N_12280);
or U16693 (N_16693,N_11737,N_13501);
xor U16694 (N_16694,N_10525,N_11481);
nor U16695 (N_16695,N_13832,N_11803);
or U16696 (N_16696,N_10105,N_14284);
nand U16697 (N_16697,N_14273,N_14458);
nand U16698 (N_16698,N_13763,N_13844);
nand U16699 (N_16699,N_10955,N_10279);
and U16700 (N_16700,N_12556,N_11128);
and U16701 (N_16701,N_11656,N_11949);
nand U16702 (N_16702,N_10492,N_14104);
xnor U16703 (N_16703,N_10973,N_14090);
xnor U16704 (N_16704,N_10598,N_14195);
nand U16705 (N_16705,N_11228,N_14665);
and U16706 (N_16706,N_12205,N_14260);
and U16707 (N_16707,N_12734,N_12819);
and U16708 (N_16708,N_14582,N_11442);
xor U16709 (N_16709,N_11844,N_13330);
nor U16710 (N_16710,N_13705,N_13055);
and U16711 (N_16711,N_14884,N_14237);
nor U16712 (N_16712,N_13521,N_14731);
nor U16713 (N_16713,N_10893,N_11878);
nand U16714 (N_16714,N_12460,N_12129);
nor U16715 (N_16715,N_14025,N_12591);
nor U16716 (N_16716,N_13131,N_10340);
nand U16717 (N_16717,N_14403,N_11635);
xor U16718 (N_16718,N_10504,N_12572);
nor U16719 (N_16719,N_10997,N_10230);
or U16720 (N_16720,N_13317,N_13182);
and U16721 (N_16721,N_12395,N_11749);
and U16722 (N_16722,N_11890,N_11582);
and U16723 (N_16723,N_11246,N_14655);
and U16724 (N_16724,N_12378,N_10818);
nand U16725 (N_16725,N_13405,N_10078);
and U16726 (N_16726,N_14510,N_11587);
or U16727 (N_16727,N_14979,N_14911);
or U16728 (N_16728,N_14365,N_13916);
or U16729 (N_16729,N_14957,N_14537);
nand U16730 (N_16730,N_14572,N_13042);
nor U16731 (N_16731,N_12135,N_12206);
and U16732 (N_16732,N_11606,N_13450);
and U16733 (N_16733,N_10927,N_14286);
nand U16734 (N_16734,N_13907,N_11823);
nor U16735 (N_16735,N_12467,N_13894);
nor U16736 (N_16736,N_11395,N_11624);
or U16737 (N_16737,N_13409,N_12216);
nand U16738 (N_16738,N_13133,N_13906);
nor U16739 (N_16739,N_12551,N_12281);
or U16740 (N_16740,N_14779,N_10094);
and U16741 (N_16741,N_14497,N_13286);
xnor U16742 (N_16742,N_11218,N_10080);
nand U16743 (N_16743,N_12337,N_12085);
nand U16744 (N_16744,N_12061,N_12315);
nor U16745 (N_16745,N_14189,N_13442);
nand U16746 (N_16746,N_10361,N_13419);
nor U16747 (N_16747,N_13298,N_14157);
and U16748 (N_16748,N_14891,N_14977);
or U16749 (N_16749,N_14671,N_10315);
nor U16750 (N_16750,N_12898,N_13318);
nor U16751 (N_16751,N_10418,N_14831);
xor U16752 (N_16752,N_14100,N_13161);
and U16753 (N_16753,N_13187,N_11027);
nand U16754 (N_16754,N_13576,N_11535);
nor U16755 (N_16755,N_14191,N_11992);
nor U16756 (N_16756,N_11695,N_12654);
nor U16757 (N_16757,N_11375,N_14774);
or U16758 (N_16758,N_10093,N_11046);
and U16759 (N_16759,N_13332,N_10761);
xor U16760 (N_16760,N_12173,N_10464);
or U16761 (N_16761,N_11714,N_10659);
or U16762 (N_16762,N_14264,N_13836);
and U16763 (N_16763,N_14961,N_10439);
and U16764 (N_16764,N_12401,N_14414);
or U16765 (N_16765,N_14056,N_10374);
or U16766 (N_16766,N_10115,N_13996);
xor U16767 (N_16767,N_11911,N_12640);
nor U16768 (N_16768,N_14947,N_13272);
nand U16769 (N_16769,N_13453,N_13734);
and U16770 (N_16770,N_10666,N_13019);
xor U16771 (N_16771,N_13927,N_11956);
and U16772 (N_16772,N_10348,N_10878);
or U16773 (N_16773,N_14339,N_12073);
nand U16774 (N_16774,N_10060,N_11610);
and U16775 (N_16775,N_11171,N_11012);
or U16776 (N_16776,N_14723,N_13467);
nand U16777 (N_16777,N_12247,N_13943);
xor U16778 (N_16778,N_11437,N_14412);
nor U16779 (N_16779,N_12899,N_11292);
nand U16780 (N_16780,N_14253,N_13592);
nor U16781 (N_16781,N_11869,N_11198);
or U16782 (N_16782,N_14372,N_13829);
nor U16783 (N_16783,N_10720,N_14934);
nor U16784 (N_16784,N_12893,N_14916);
nor U16785 (N_16785,N_12588,N_10859);
nor U16786 (N_16786,N_11810,N_10934);
and U16787 (N_16787,N_10432,N_14097);
nor U16788 (N_16788,N_14289,N_10349);
and U16789 (N_16789,N_11491,N_13891);
nor U16790 (N_16790,N_14353,N_13774);
xor U16791 (N_16791,N_13794,N_10734);
or U16792 (N_16792,N_11821,N_10975);
or U16793 (N_16793,N_12684,N_13839);
and U16794 (N_16794,N_11469,N_10803);
nor U16795 (N_16795,N_10380,N_11834);
nor U16796 (N_16796,N_11487,N_12382);
nand U16797 (N_16797,N_12379,N_13947);
and U16798 (N_16798,N_10609,N_10503);
or U16799 (N_16799,N_14358,N_14691);
nand U16800 (N_16800,N_13769,N_12366);
or U16801 (N_16801,N_14714,N_12499);
or U16802 (N_16802,N_14593,N_14985);
and U16803 (N_16803,N_11682,N_12771);
and U16804 (N_16804,N_13483,N_13203);
nor U16805 (N_16805,N_12720,N_12825);
xor U16806 (N_16806,N_14511,N_12564);
or U16807 (N_16807,N_13545,N_11616);
nor U16808 (N_16808,N_11498,N_10189);
and U16809 (N_16809,N_14110,N_14293);
or U16810 (N_16810,N_14634,N_11123);
nor U16811 (N_16811,N_13564,N_11625);
nand U16812 (N_16812,N_13533,N_10228);
or U16813 (N_16813,N_13407,N_14600);
or U16814 (N_16814,N_13864,N_10932);
or U16815 (N_16815,N_14294,N_10283);
xor U16816 (N_16816,N_13959,N_13432);
or U16817 (N_16817,N_12622,N_10270);
nand U16818 (N_16818,N_14360,N_12475);
nand U16819 (N_16819,N_13837,N_10023);
or U16820 (N_16820,N_12332,N_13311);
or U16821 (N_16821,N_14674,N_10903);
nor U16822 (N_16822,N_11633,N_12682);
or U16823 (N_16823,N_13151,N_14465);
and U16824 (N_16824,N_10347,N_11466);
nor U16825 (N_16825,N_11880,N_12543);
or U16826 (N_16826,N_12940,N_10602);
or U16827 (N_16827,N_11545,N_11220);
and U16828 (N_16828,N_14330,N_14159);
or U16829 (N_16829,N_14852,N_14070);
or U16830 (N_16830,N_11787,N_12024);
or U16831 (N_16831,N_14204,N_11092);
nand U16832 (N_16832,N_14886,N_13762);
nand U16833 (N_16833,N_14145,N_10849);
or U16834 (N_16834,N_14212,N_13809);
or U16835 (N_16835,N_10344,N_10873);
or U16836 (N_16836,N_12229,N_11238);
and U16837 (N_16837,N_11078,N_10614);
nand U16838 (N_16838,N_11569,N_10390);
nand U16839 (N_16839,N_12714,N_12491);
xnor U16840 (N_16840,N_10876,N_10356);
and U16841 (N_16841,N_13534,N_13714);
and U16842 (N_16842,N_12140,N_10848);
nand U16843 (N_16843,N_14717,N_11281);
nor U16844 (N_16844,N_12988,N_14974);
and U16845 (N_16845,N_14518,N_10155);
xor U16846 (N_16846,N_11022,N_11157);
and U16847 (N_16847,N_14988,N_11540);
and U16848 (N_16848,N_12256,N_14305);
nand U16849 (N_16849,N_11770,N_12755);
or U16850 (N_16850,N_13169,N_12710);
and U16851 (N_16851,N_13670,N_14501);
nor U16852 (N_16852,N_11043,N_14604);
or U16853 (N_16853,N_13154,N_11930);
and U16854 (N_16854,N_13667,N_12857);
nor U16855 (N_16855,N_11308,N_14001);
xor U16856 (N_16856,N_14082,N_11728);
and U16857 (N_16857,N_12010,N_14004);
or U16858 (N_16858,N_10938,N_12350);
or U16859 (N_16859,N_10584,N_10368);
and U16860 (N_16860,N_12897,N_11578);
nor U16861 (N_16861,N_11011,N_14544);
nand U16862 (N_16862,N_11736,N_13726);
or U16863 (N_16863,N_14601,N_10895);
nor U16864 (N_16864,N_14040,N_14041);
or U16865 (N_16865,N_13249,N_13536);
nand U16866 (N_16866,N_12005,N_13074);
nand U16867 (N_16867,N_14168,N_12960);
nand U16868 (N_16868,N_14078,N_12096);
nor U16869 (N_16869,N_12980,N_12852);
xor U16870 (N_16870,N_13910,N_11568);
or U16871 (N_16871,N_13870,N_12109);
xnor U16872 (N_16872,N_13124,N_12788);
or U16873 (N_16873,N_10436,N_14114);
nor U16874 (N_16874,N_10771,N_13671);
or U16875 (N_16875,N_13595,N_12907);
and U16876 (N_16876,N_12694,N_11476);
xor U16877 (N_16877,N_12951,N_13142);
nor U16878 (N_16878,N_12448,N_10904);
nand U16879 (N_16879,N_13849,N_12301);
or U16880 (N_16880,N_11644,N_13636);
nand U16881 (N_16881,N_11565,N_14417);
and U16882 (N_16882,N_11000,N_14061);
nor U16883 (N_16883,N_10147,N_13593);
or U16884 (N_16884,N_10170,N_12837);
nand U16885 (N_16885,N_13695,N_13573);
nand U16886 (N_16886,N_10842,N_10482);
and U16887 (N_16887,N_11671,N_11385);
and U16888 (N_16888,N_12105,N_11683);
nand U16889 (N_16889,N_10521,N_10063);
nor U16890 (N_16890,N_14624,N_12827);
xor U16891 (N_16891,N_11297,N_11659);
nand U16892 (N_16892,N_14927,N_13307);
or U16893 (N_16893,N_12210,N_14751);
nand U16894 (N_16894,N_14635,N_13335);
nand U16895 (N_16895,N_11702,N_13651);
nand U16896 (N_16896,N_10038,N_12962);
or U16897 (N_16897,N_11480,N_14245);
or U16898 (N_16898,N_11073,N_13644);
nor U16899 (N_16899,N_11101,N_12020);
and U16900 (N_16900,N_13969,N_13037);
or U16901 (N_16901,N_13991,N_13141);
nor U16902 (N_16902,N_12201,N_12489);
nor U16903 (N_16903,N_11286,N_11813);
nand U16904 (N_16904,N_12888,N_11099);
nor U16905 (N_16905,N_13077,N_14093);
and U16906 (N_16906,N_10403,N_11906);
and U16907 (N_16907,N_12925,N_14270);
and U16908 (N_16908,N_14504,N_12457);
nand U16909 (N_16909,N_12858,N_13719);
or U16910 (N_16910,N_14856,N_12642);
nor U16911 (N_16911,N_11923,N_14352);
nand U16912 (N_16912,N_14765,N_12157);
xor U16913 (N_16913,N_10058,N_14006);
nor U16914 (N_16914,N_10906,N_11036);
or U16915 (N_16915,N_13474,N_10603);
nor U16916 (N_16916,N_13229,N_14217);
or U16917 (N_16917,N_13738,N_14702);
xor U16918 (N_16918,N_14020,N_13856);
nand U16919 (N_16919,N_12148,N_10804);
or U16920 (N_16920,N_11239,N_12892);
and U16921 (N_16921,N_11707,N_12309);
or U16922 (N_16922,N_13347,N_10687);
and U16923 (N_16923,N_12415,N_13255);
nand U16924 (N_16924,N_14215,N_13320);
and U16925 (N_16925,N_10499,N_14334);
nor U16926 (N_16926,N_12076,N_14252);
nand U16927 (N_16927,N_13415,N_13566);
nand U16928 (N_16928,N_13803,N_11458);
xnor U16929 (N_16929,N_12204,N_12399);
nand U16930 (N_16930,N_13302,N_12587);
and U16931 (N_16931,N_13628,N_10970);
nor U16932 (N_16932,N_10375,N_10991);
nor U16933 (N_16933,N_10514,N_12340);
nand U16934 (N_16934,N_14395,N_14729);
or U16935 (N_16935,N_14079,N_10428);
or U16936 (N_16936,N_13293,N_14700);
xnor U16937 (N_16937,N_10832,N_14393);
and U16938 (N_16938,N_12895,N_12579);
nand U16939 (N_16939,N_11874,N_14306);
nor U16940 (N_16940,N_13412,N_13492);
nand U16941 (N_16941,N_13813,N_10272);
or U16942 (N_16942,N_12503,N_12081);
nand U16943 (N_16943,N_14072,N_12275);
or U16944 (N_16944,N_12009,N_13048);
nor U16945 (N_16945,N_13242,N_11976);
or U16946 (N_16946,N_11608,N_12238);
nand U16947 (N_16947,N_10948,N_13929);
and U16948 (N_16948,N_11567,N_10453);
or U16949 (N_16949,N_10486,N_10765);
or U16950 (N_16950,N_10062,N_12111);
and U16951 (N_16951,N_14391,N_11808);
and U16952 (N_16952,N_12172,N_10443);
or U16953 (N_16953,N_10774,N_10388);
and U16954 (N_16954,N_12570,N_13515);
nand U16955 (N_16955,N_12117,N_13164);
nor U16956 (N_16956,N_10697,N_11173);
or U16957 (N_16957,N_12973,N_12424);
nand U16958 (N_16958,N_10863,N_13540);
or U16959 (N_16959,N_11457,N_14503);
and U16960 (N_16960,N_10788,N_13786);
nor U16961 (N_16961,N_11521,N_14838);
and U16962 (N_16962,N_12416,N_13723);
and U16963 (N_16963,N_14543,N_14155);
nand U16964 (N_16964,N_14533,N_11357);
nand U16965 (N_16965,N_10776,N_11793);
nand U16966 (N_16966,N_14058,N_11461);
nand U16967 (N_16967,N_10665,N_11219);
or U16968 (N_16968,N_14524,N_13588);
nand U16969 (N_16969,N_10621,N_12546);
nor U16970 (N_16970,N_12144,N_11853);
or U16971 (N_16971,N_11827,N_12584);
nor U16972 (N_16972,N_11797,N_10533);
or U16973 (N_16973,N_13646,N_12606);
and U16974 (N_16974,N_11864,N_14775);
and U16975 (N_16975,N_13941,N_14384);
or U16976 (N_16976,N_13633,N_11401);
or U16977 (N_16977,N_10236,N_13022);
or U16978 (N_16978,N_11484,N_11100);
nand U16979 (N_16979,N_12569,N_14681);
nand U16980 (N_16980,N_13503,N_12783);
nor U16981 (N_16981,N_13326,N_11586);
and U16982 (N_16982,N_14773,N_13477);
nand U16983 (N_16983,N_13295,N_12946);
nand U16984 (N_16984,N_11400,N_12567);
nand U16985 (N_16985,N_13607,N_14105);
or U16986 (N_16986,N_13656,N_14150);
nor U16987 (N_16987,N_13231,N_12685);
xnor U16988 (N_16988,N_12660,N_13961);
nand U16989 (N_16989,N_12807,N_10259);
and U16990 (N_16990,N_12861,N_12128);
nor U16991 (N_16991,N_14419,N_13115);
nor U16992 (N_16992,N_13102,N_14633);
nor U16993 (N_16993,N_12191,N_14690);
and U16994 (N_16994,N_11180,N_13271);
nand U16995 (N_16995,N_10717,N_13988);
nor U16996 (N_16996,N_12402,N_10669);
nor U16997 (N_16997,N_10555,N_14895);
and U16998 (N_16998,N_10944,N_12373);
nand U16999 (N_16999,N_10373,N_10819);
nand U17000 (N_17000,N_12528,N_11355);
and U17001 (N_17001,N_14466,N_12832);
xor U17002 (N_17002,N_12932,N_12853);
nor U17003 (N_17003,N_10939,N_11871);
and U17004 (N_17004,N_12207,N_11991);
nand U17005 (N_17005,N_12474,N_11609);
nand U17006 (N_17006,N_11537,N_10280);
and U17007 (N_17007,N_13967,N_13742);
nor U17008 (N_17008,N_14307,N_10018);
and U17009 (N_17009,N_10885,N_11271);
and U17010 (N_17010,N_11708,N_14042);
nand U17011 (N_17011,N_11366,N_12766);
and U17012 (N_17012,N_13469,N_11765);
nor U17013 (N_17013,N_10024,N_11831);
nor U17014 (N_17014,N_12036,N_11386);
nor U17015 (N_17015,N_12561,N_10387);
and U17016 (N_17016,N_12040,N_13862);
nand U17017 (N_17017,N_14692,N_10040);
nor U17018 (N_17018,N_11763,N_14274);
and U17019 (N_17019,N_13256,N_11999);
xnor U17020 (N_17020,N_13337,N_14063);
or U17021 (N_17021,N_11146,N_13013);
xor U17022 (N_17022,N_14923,N_10892);
nand U17023 (N_17023,N_14931,N_10637);
xor U17024 (N_17024,N_12901,N_11126);
nand U17025 (N_17025,N_14508,N_10437);
xor U17026 (N_17026,N_11017,N_13624);
nand U17027 (N_17027,N_14453,N_13428);
xnor U17028 (N_17028,N_11822,N_10157);
nor U17029 (N_17029,N_12271,N_13340);
nand U17030 (N_17030,N_14120,N_11734);
nor U17031 (N_17031,N_14549,N_13704);
nor U17032 (N_17032,N_14817,N_12604);
nand U17033 (N_17033,N_13360,N_10286);
xnor U17034 (N_17034,N_14200,N_10177);
or U17035 (N_17035,N_10680,N_14622);
nand U17036 (N_17036,N_10247,N_10162);
nor U17037 (N_17037,N_13471,N_11072);
xnor U17038 (N_17038,N_10088,N_14108);
or U17039 (N_17039,N_12292,N_14460);
or U17040 (N_17040,N_12833,N_14427);
and U17041 (N_17041,N_12276,N_10298);
nor U17042 (N_17042,N_14052,N_10056);
and U17043 (N_17043,N_12498,N_12179);
or U17044 (N_17044,N_13921,N_13841);
xor U17045 (N_17045,N_12915,N_10473);
and U17046 (N_17046,N_12333,N_13278);
and U17047 (N_17047,N_11968,N_14477);
nor U17048 (N_17048,N_13848,N_12699);
nor U17049 (N_17049,N_14953,N_13207);
or U17050 (N_17050,N_11251,N_13466);
nor U17051 (N_17051,N_14131,N_12064);
nand U17052 (N_17052,N_14349,N_14194);
or U17053 (N_17053,N_11528,N_14825);
and U17054 (N_17054,N_13252,N_13613);
nand U17055 (N_17055,N_14373,N_11873);
xnor U17056 (N_17056,N_11675,N_14269);
and U17057 (N_17057,N_14566,N_11807);
nand U17058 (N_17058,N_13137,N_11446);
and U17059 (N_17059,N_11096,N_13004);
or U17060 (N_17060,N_13244,N_14162);
or U17061 (N_17061,N_14538,N_10091);
nor U17062 (N_17062,N_13707,N_13964);
and U17063 (N_17063,N_14534,N_10365);
nand U17064 (N_17064,N_11886,N_13219);
and U17065 (N_17065,N_11815,N_10407);
nand U17066 (N_17066,N_11265,N_12119);
and U17067 (N_17067,N_13488,N_10121);
and U17068 (N_17068,N_10961,N_14369);
xor U17069 (N_17069,N_13447,N_11833);
or U17070 (N_17070,N_13336,N_10578);
or U17071 (N_17071,N_13240,N_14984);
or U17072 (N_17072,N_13265,N_10086);
xor U17073 (N_17073,N_10563,N_12919);
and U17074 (N_17074,N_12547,N_14847);
and U17075 (N_17075,N_11927,N_10367);
nand U17076 (N_17076,N_11536,N_11348);
and U17077 (N_17077,N_10127,N_10714);
and U17078 (N_17078,N_14547,N_11409);
nor U17079 (N_17079,N_12390,N_11600);
nor U17080 (N_17080,N_11549,N_10066);
or U17081 (N_17081,N_12314,N_10736);
and U17082 (N_17082,N_13434,N_11010);
and U17083 (N_17083,N_14438,N_14371);
nor U17084 (N_17084,N_10917,N_10738);
xnor U17085 (N_17085,N_12847,N_10297);
and U17086 (N_17086,N_14169,N_11069);
nand U17087 (N_17087,N_11789,N_12121);
and U17088 (N_17088,N_11974,N_14502);
or U17089 (N_17089,N_14656,N_13581);
nor U17090 (N_17090,N_11091,N_11313);
xnor U17091 (N_17091,N_14454,N_14992);
and U17092 (N_17092,N_14074,N_12249);
nand U17093 (N_17093,N_11391,N_12670);
and U17094 (N_17094,N_12653,N_10469);
xnor U17095 (N_17095,N_14559,N_13382);
nor U17096 (N_17096,N_12651,N_13139);
nor U17097 (N_17097,N_14083,N_14594);
nand U17098 (N_17098,N_13323,N_10244);
nor U17099 (N_17099,N_11483,N_12838);
nand U17100 (N_17100,N_13855,N_11084);
and U17101 (N_17101,N_13998,N_12544);
and U17102 (N_17102,N_12236,N_14186);
nor U17103 (N_17103,N_10097,N_12431);
or U17104 (N_17104,N_12646,N_13979);
nand U17105 (N_17105,N_13334,N_10708);
nand U17106 (N_17106,N_10686,N_12830);
or U17107 (N_17107,N_11353,N_14666);
nor U17108 (N_17108,N_13017,N_11539);
nand U17109 (N_17109,N_12754,N_13620);
nor U17110 (N_17110,N_11351,N_12264);
or U17111 (N_17111,N_11526,N_14010);
and U17112 (N_17112,N_11403,N_11326);
nand U17113 (N_17113,N_10718,N_11700);
nor U17114 (N_17114,N_11592,N_13456);
nor U17115 (N_17115,N_12541,N_12979);
nor U17116 (N_17116,N_10429,N_13396);
xnor U17117 (N_17117,N_10310,N_10952);
or U17118 (N_17118,N_14354,N_13510);
nor U17119 (N_17119,N_12798,N_14704);
nor U17120 (N_17120,N_11887,N_10506);
and U17121 (N_17121,N_13589,N_13987);
or U17122 (N_17122,N_14167,N_13563);
or U17123 (N_17123,N_10363,N_14912);
nand U17124 (N_17124,N_11672,N_10357);
and U17125 (N_17125,N_10463,N_10931);
and U17126 (N_17126,N_12904,N_12614);
or U17127 (N_17127,N_11410,N_11993);
xor U17128 (N_17128,N_10500,N_12621);
or U17129 (N_17129,N_13024,N_10690);
and U17130 (N_17130,N_14123,N_10371);
nor U17131 (N_17131,N_10985,N_14033);
or U17132 (N_17132,N_11053,N_11950);
or U17133 (N_17133,N_14362,N_14799);
or U17134 (N_17134,N_12407,N_12998);
and U17135 (N_17135,N_10673,N_13928);
nand U17136 (N_17136,N_11885,N_14483);
nand U17137 (N_17137,N_11934,N_14314);
or U17138 (N_17138,N_13175,N_11701);
nor U17139 (N_17139,N_12326,N_14255);
nor U17140 (N_17140,N_14142,N_11724);
and U17141 (N_17141,N_13560,N_14828);
or U17142 (N_17142,N_14046,N_13871);
nand U17143 (N_17143,N_10618,N_10008);
nand U17144 (N_17144,N_10739,N_13233);
xor U17145 (N_17145,N_13067,N_13567);
nor U17146 (N_17146,N_10733,N_13579);
or U17147 (N_17147,N_11315,N_10427);
nand U17148 (N_17148,N_10591,N_13805);
nor U17149 (N_17149,N_13491,N_11346);
or U17150 (N_17150,N_11259,N_10251);
nand U17151 (N_17151,N_10745,N_14797);
nand U17152 (N_17152,N_12018,N_11034);
or U17153 (N_17153,N_12384,N_11800);
nand U17154 (N_17154,N_14313,N_12331);
nand U17155 (N_17155,N_10793,N_13782);
xor U17156 (N_17156,N_14529,N_12903);
nand U17157 (N_17157,N_11152,N_13743);
and U17158 (N_17158,N_12743,N_12317);
and U17159 (N_17159,N_14972,N_14172);
or U17160 (N_17160,N_10809,N_12181);
nand U17161 (N_17161,N_14584,N_10302);
nor U17162 (N_17162,N_10671,N_11931);
xor U17163 (N_17163,N_10171,N_13009);
nor U17164 (N_17164,N_13647,N_11661);
nand U17165 (N_17165,N_11627,N_14336);
and U17166 (N_17166,N_12635,N_14658);
nor U17167 (N_17167,N_11471,N_12488);
and U17168 (N_17168,N_13245,N_13264);
nor U17169 (N_17169,N_10042,N_10568);
and U17170 (N_17170,N_12786,N_10966);
nor U17171 (N_17171,N_13470,N_12253);
nand U17172 (N_17172,N_14668,N_10889);
or U17173 (N_17173,N_14764,N_13537);
nand U17174 (N_17174,N_12632,N_11622);
nand U17175 (N_17175,N_10624,N_12410);
nor U17176 (N_17176,N_12618,N_13043);
nand U17177 (N_17177,N_12793,N_11732);
or U17178 (N_17178,N_13068,N_13223);
xor U17179 (N_17179,N_10937,N_14769);
nor U17180 (N_17180,N_11534,N_14962);
nand U17181 (N_17181,N_12727,N_14316);
xor U17182 (N_17182,N_12272,N_13034);
and U17183 (N_17183,N_14227,N_11959);
nor U17184 (N_17184,N_12187,N_14618);
nor U17185 (N_17185,N_10612,N_11527);
and U17186 (N_17186,N_13661,N_14491);
nand U17187 (N_17187,N_13641,N_11453);
xor U17188 (N_17188,N_10336,N_11127);
xor U17189 (N_17189,N_12008,N_10199);
and U17190 (N_17190,N_12896,N_10126);
and U17191 (N_17191,N_10635,N_10391);
and U17192 (N_17192,N_12289,N_11727);
nor U17193 (N_17193,N_11505,N_13968);
or U17194 (N_17194,N_13140,N_14437);
and U17195 (N_17195,N_12374,N_10314);
and U17196 (N_17196,N_12497,N_12242);
or U17197 (N_17197,N_14876,N_11723);
and U17198 (N_17198,N_14401,N_12261);
nor U17199 (N_17199,N_14490,N_13086);
and U17200 (N_17200,N_12060,N_11063);
nand U17201 (N_17201,N_11863,N_11208);
and U17202 (N_17202,N_10836,N_10626);
or U17203 (N_17203,N_12007,N_13933);
and U17204 (N_17204,N_13604,N_13642);
nand U17205 (N_17205,N_11867,N_10700);
nor U17206 (N_17206,N_11577,N_13502);
or U17207 (N_17207,N_12822,N_12313);
nor U17208 (N_17208,N_11212,N_14762);
and U17209 (N_17209,N_10471,N_13899);
nor U17210 (N_17210,N_13006,N_14351);
xnor U17211 (N_17211,N_10729,N_10530);
nand U17212 (N_17212,N_12724,N_10518);
xnor U17213 (N_17213,N_12974,N_11080);
and U17214 (N_17214,N_10713,N_13895);
nand U17215 (N_17215,N_11151,N_10151);
nand U17216 (N_17216,N_14190,N_10576);
xnor U17217 (N_17217,N_11791,N_11604);
nor U17218 (N_17218,N_12645,N_12277);
or U17219 (N_17219,N_14581,N_11252);
and U17220 (N_17220,N_12239,N_13840);
xnor U17221 (N_17221,N_11211,N_11548);
nor U17222 (N_17222,N_12894,N_10699);
xor U17223 (N_17223,N_12715,N_13650);
nand U17224 (N_17224,N_11176,N_12638);
nor U17225 (N_17225,N_13801,N_13681);
nor U17226 (N_17226,N_12780,N_12209);
xnor U17227 (N_17227,N_12955,N_12975);
nand U17228 (N_17228,N_13807,N_11958);
nand U17229 (N_17229,N_14443,N_14776);
nor U17230 (N_17230,N_10983,N_12697);
nand U17231 (N_17231,N_13162,N_14228);
or U17232 (N_17232,N_14326,N_13520);
nand U17233 (N_17233,N_11125,N_12592);
xor U17234 (N_17234,N_14750,N_12380);
and U17235 (N_17235,N_11201,N_10281);
nor U17236 (N_17236,N_14609,N_13475);
or U17237 (N_17237,N_14832,N_11612);
and U17238 (N_17238,N_12056,N_14210);
and U17239 (N_17239,N_11376,N_13076);
or U17240 (N_17240,N_10627,N_11429);
and U17241 (N_17241,N_14981,N_10498);
nand U17242 (N_17242,N_12756,N_13655);
nand U17243 (N_17243,N_13056,N_10353);
nand U17244 (N_17244,N_12351,N_10852);
or U17245 (N_17245,N_10460,N_12557);
or U17246 (N_17246,N_14565,N_11523);
or U17247 (N_17247,N_14485,N_12019);
or U17248 (N_17248,N_10169,N_13308);
or U17249 (N_17249,N_14564,N_14662);
or U17250 (N_17250,N_11112,N_14012);
xor U17251 (N_17251,N_11178,N_11402);
and U17252 (N_17252,N_11562,N_10456);
and U17253 (N_17253,N_10559,N_10359);
nor U17254 (N_17254,N_10102,N_11247);
or U17255 (N_17255,N_12098,N_13380);
or U17256 (N_17256,N_12669,N_10470);
nor U17257 (N_17257,N_13435,N_10084);
xor U17258 (N_17258,N_12279,N_13129);
or U17259 (N_17259,N_14816,N_12559);
nand U17260 (N_17260,N_14222,N_10529);
and U17261 (N_17261,N_10362,N_13639);
nand U17262 (N_17262,N_13210,N_10951);
nor U17263 (N_17263,N_11602,N_13846);
nor U17264 (N_17264,N_10978,N_11163);
nor U17265 (N_17265,N_12770,N_10322);
or U17266 (N_17266,N_12298,N_10837);
or U17267 (N_17267,N_14192,N_10766);
or U17268 (N_17268,N_14254,N_11940);
or U17269 (N_17269,N_11738,N_14049);
nand U17270 (N_17270,N_13290,N_11963);
nor U17271 (N_17271,N_13555,N_14214);
nand U17272 (N_17272,N_14531,N_10656);
and U17273 (N_17273,N_13087,N_11141);
and U17274 (N_17274,N_10282,N_14323);
nand U17275 (N_17275,N_12831,N_10006);
xnor U17276 (N_17276,N_13446,N_12555);
nor U17277 (N_17277,N_14059,N_13121);
or U17278 (N_17278,N_14542,N_11713);
and U17279 (N_17279,N_14770,N_14505);
and U17280 (N_17280,N_10209,N_11008);
xor U17281 (N_17281,N_11997,N_14783);
or U17282 (N_17282,N_14844,N_13120);
nor U17283 (N_17283,N_14471,N_14598);
and U17284 (N_17284,N_13426,N_14526);
or U17285 (N_17285,N_12811,N_10615);
nand U17286 (N_17286,N_12262,N_12293);
or U17287 (N_17287,N_11977,N_11970);
nor U17288 (N_17288,N_14933,N_11320);
nand U17289 (N_17289,N_10592,N_12158);
or U17290 (N_17290,N_12986,N_11899);
nor U17291 (N_17291,N_14397,N_14703);
or U17292 (N_17292,N_13830,N_14610);
nor U17293 (N_17293,N_14641,N_11370);
or U17294 (N_17294,N_12971,N_12323);
or U17295 (N_17295,N_14178,N_10485);
or U17296 (N_17296,N_11224,N_14673);
and U17297 (N_17297,N_10608,N_12700);
or U17298 (N_17298,N_12228,N_12381);
or U17299 (N_17299,N_13384,N_10590);
or U17300 (N_17300,N_12086,N_12075);
xnor U17301 (N_17301,N_10544,N_12164);
xor U17302 (N_17302,N_10134,N_14247);
and U17303 (N_17303,N_10747,N_12083);
or U17304 (N_17304,N_13522,N_12327);
or U17305 (N_17305,N_13744,N_14727);
and U17306 (N_17306,N_13889,N_11838);
or U17307 (N_17307,N_12993,N_10707);
or U17308 (N_17308,N_10763,N_12213);
nand U17309 (N_17309,N_10433,N_11417);
xor U17310 (N_17310,N_11161,N_13059);
xnor U17311 (N_17311,N_14653,N_11187);
xnor U17312 (N_17312,N_14719,N_13445);
or U17313 (N_17313,N_11556,N_13315);
nand U17314 (N_17314,N_14822,N_10011);
and U17315 (N_17315,N_12193,N_10052);
nor U17316 (N_17316,N_10168,N_11120);
nor U17317 (N_17317,N_10995,N_10660);
nand U17318 (N_17318,N_10424,N_13802);
nor U17319 (N_17319,N_11298,N_14408);
and U17320 (N_17320,N_13292,N_12387);
and U17321 (N_17321,N_10539,N_11551);
xor U17322 (N_17322,N_14421,N_12200);
nand U17323 (N_17323,N_10181,N_13021);
xnor U17324 (N_17324,N_14185,N_13880);
nand U17325 (N_17325,N_12849,N_14904);
nand U17326 (N_17326,N_12299,N_12302);
nand U17327 (N_17327,N_11918,N_13200);
nand U17328 (N_17328,N_13310,N_12999);
nand U17329 (N_17329,N_11021,N_14790);
and U17330 (N_17330,N_12436,N_13147);
nor U17331 (N_17331,N_13322,N_13669);
nor U17332 (N_17332,N_14514,N_14418);
nand U17333 (N_17333,N_12910,N_11282);
and U17334 (N_17334,N_13583,N_12443);
or U17335 (N_17335,N_10188,N_11730);
nand U17336 (N_17336,N_13824,N_11756);
nand U17337 (N_17337,N_12397,N_11919);
nor U17338 (N_17338,N_11677,N_12202);
or U17339 (N_17339,N_11248,N_10797);
nand U17340 (N_17340,N_12978,N_14993);
nand U17341 (N_17341,N_12703,N_10651);
xnor U17342 (N_17342,N_10275,N_11721);
nand U17343 (N_17343,N_10730,N_13610);
and U17344 (N_17344,N_13464,N_11200);
and U17345 (N_17345,N_10828,N_14726);
nor U17346 (N_17346,N_14697,N_12185);
or U17347 (N_17347,N_10638,N_13715);
xor U17348 (N_17348,N_11037,N_14659);
nor U17349 (N_17349,N_10601,N_14997);
nand U17350 (N_17350,N_11318,N_14328);
nor U17351 (N_17351,N_14712,N_14515);
nand U17352 (N_17352,N_13354,N_13529);
or U17353 (N_17353,N_11839,N_10688);
nor U17354 (N_17354,N_13513,N_12744);
nor U17355 (N_17355,N_13215,N_12680);
xor U17356 (N_17356,N_12922,N_12790);
and U17357 (N_17357,N_14415,N_13253);
nor U17358 (N_17358,N_13912,N_10192);
nor U17359 (N_17359,N_13217,N_12976);
nor U17360 (N_17360,N_10556,N_14557);
and U17361 (N_17361,N_13518,N_11719);
nand U17362 (N_17362,N_13127,N_11947);
nand U17363 (N_17363,N_12512,N_13047);
and U17364 (N_17364,N_12305,N_13937);
and U17365 (N_17365,N_13046,N_10871);
or U17366 (N_17366,N_13561,N_10261);
nand U17367 (N_17367,N_12985,N_11193);
or U17368 (N_17368,N_10039,N_10644);
and U17369 (N_17369,N_12954,N_13383);
and U17370 (N_17370,N_10401,N_13697);
nor U17371 (N_17371,N_10580,N_14867);
nor U17372 (N_17372,N_10296,N_14400);
nand U17373 (N_17373,N_10158,N_12511);
xor U17374 (N_17374,N_10010,N_13663);
nor U17375 (N_17375,N_10652,N_13496);
nor U17376 (N_17376,N_12969,N_14479);
nand U17377 (N_17377,N_12495,N_10589);
or U17378 (N_17378,N_13770,N_11891);
and U17379 (N_17379,N_13694,N_14809);
xor U17380 (N_17380,N_10883,N_13546);
or U17381 (N_17381,N_11324,N_11646);
nor U17382 (N_17382,N_10493,N_11379);
and U17383 (N_17383,N_11418,N_12147);
and U17384 (N_17384,N_13441,N_10823);
or U17385 (N_17385,N_12195,N_10212);
or U17386 (N_17386,N_11960,N_10312);
nor U17387 (N_17387,N_13771,N_13897);
xnor U17388 (N_17388,N_10950,N_13925);
and U17389 (N_17389,N_11473,N_13153);
and U17390 (N_17390,N_10512,N_13815);
and U17391 (N_17391,N_14224,N_14651);
nor U17392 (N_17392,N_14022,N_13429);
nand U17393 (N_17393,N_10381,N_12484);
or U17394 (N_17394,N_11531,N_13170);
nor U17395 (N_17395,N_10331,N_10569);
and U17396 (N_17396,N_10622,N_11422);
or U17397 (N_17397,N_11762,N_14154);
nand U17398 (N_17398,N_13341,N_13989);
nand U17399 (N_17399,N_10068,N_10087);
nand U17400 (N_17400,N_13594,N_14474);
and U17401 (N_17401,N_10491,N_12916);
or U17402 (N_17402,N_10704,N_11452);
nor U17403 (N_17403,N_14347,N_10258);
nand U17404 (N_17404,N_12364,N_12959);
nor U17405 (N_17405,N_13611,N_10650);
nand U17406 (N_17406,N_12914,N_12237);
xnor U17407 (N_17407,N_13708,N_13319);
or U17408 (N_17408,N_12452,N_14456);
nand U17409 (N_17409,N_11273,N_14935);
nand U17410 (N_17410,N_12598,N_12370);
nand U17411 (N_17411,N_12816,N_11145);
xnor U17412 (N_17412,N_11941,N_12742);
nor U17413 (N_17413,N_12883,N_12801);
nand U17414 (N_17414,N_13058,N_12881);
nor U17415 (N_17415,N_10338,N_14987);
and U17416 (N_17416,N_11465,N_11849);
or U17417 (N_17417,N_12519,N_14024);
nand U17418 (N_17418,N_11666,N_11175);
and U17419 (N_17419,N_14522,N_12231);
or U17420 (N_17420,N_11456,N_14724);
xnor U17421 (N_17421,N_14376,N_13266);
xor U17422 (N_17422,N_14388,N_12607);
nand U17423 (N_17423,N_14611,N_11260);
or U17424 (N_17424,N_10316,N_10986);
or U17425 (N_17425,N_14468,N_14586);
or U17426 (N_17426,N_13303,N_12859);
nor U17427 (N_17427,N_11952,N_12624);
nor U17428 (N_17428,N_14482,N_12449);
and U17429 (N_17429,N_14743,N_14871);
and U17430 (N_17430,N_13790,N_12615);
or U17431 (N_17431,N_11062,N_14625);
and U17432 (N_17432,N_12167,N_13420);
and U17433 (N_17433,N_10905,N_14976);
nor U17434 (N_17434,N_13400,N_11232);
nand U17435 (N_17435,N_12125,N_12047);
nor U17436 (N_17436,N_12230,N_10130);
and U17437 (N_17437,N_13399,N_12865);
and U17438 (N_17438,N_11098,N_11345);
nand U17439 (N_17439,N_14130,N_11340);
and U17440 (N_17440,N_14446,N_13635);
nand U17441 (N_17441,N_14242,N_11530);
xor U17442 (N_17442,N_10751,N_12226);
or U17443 (N_17443,N_12945,N_11048);
nor U17444 (N_17444,N_14312,N_12545);
nor U17445 (N_17445,N_11799,N_14954);
or U17446 (N_17446,N_11641,N_11071);
or U17447 (N_17447,N_14616,N_10198);
nor U17448 (N_17448,N_10958,N_12595);
nand U17449 (N_17449,N_11235,N_14872);
and U17450 (N_17450,N_11205,N_13686);
and U17451 (N_17451,N_11650,N_12490);
nor U17452 (N_17452,N_12887,N_11333);
nand U17453 (N_17453,N_13028,N_12160);
nand U17454 (N_17454,N_10616,N_12375);
nor U17455 (N_17455,N_14303,N_12918);
or U17456 (N_17456,N_13075,N_10101);
nand U17457 (N_17457,N_12456,N_11216);
or U17458 (N_17458,N_13674,N_13381);
or U17459 (N_17459,N_14552,N_10266);
or U17460 (N_17460,N_12246,N_11257);
and U17461 (N_17461,N_11897,N_12935);
or U17462 (N_17462,N_13516,N_13528);
nor U17463 (N_17463,N_11464,N_10070);
nand U17464 (N_17464,N_14266,N_11309);
and U17465 (N_17465,N_11900,N_11629);
nor U17466 (N_17466,N_12717,N_10253);
xor U17467 (N_17467,N_10820,N_14277);
or U17468 (N_17468,N_14422,N_10655);
or U17469 (N_17469,N_12532,N_10693);
and U17470 (N_17470,N_14406,N_12563);
nand U17471 (N_17471,N_12549,N_10234);
and U17472 (N_17472,N_10710,N_13724);
xor U17473 (N_17473,N_13958,N_14457);
and U17474 (N_17474,N_13627,N_12599);
or U17475 (N_17475,N_11217,N_10389);
or U17476 (N_17476,N_11441,N_11731);
or U17477 (N_17477,N_14808,N_11643);
nor U17478 (N_17478,N_14177,N_10570);
nand U17479 (N_17479,N_13525,N_10215);
nor U17480 (N_17480,N_13772,N_12513);
nor U17481 (N_17481,N_12509,N_11280);
and U17482 (N_17482,N_11936,N_12704);
nor U17483 (N_17483,N_11377,N_12245);
and U17484 (N_17484,N_12361,N_10144);
xor U17485 (N_17485,N_14848,N_10049);
or U17486 (N_17486,N_13552,N_12885);
or U17487 (N_17487,N_14138,N_14396);
nor U17488 (N_17488,N_12349,N_12675);
xor U17489 (N_17489,N_10574,N_12290);
nor U17490 (N_17490,N_10808,N_12812);
nand U17491 (N_17491,N_10884,N_11032);
and U17492 (N_17492,N_11361,N_14827);
or U17493 (N_17493,N_11786,N_14387);
or U17494 (N_17494,N_13234,N_10076);
xnor U17495 (N_17495,N_10273,N_13494);
and U17496 (N_17496,N_13547,N_10692);
nand U17497 (N_17497,N_10998,N_11065);
xnor U17498 (N_17498,N_10386,N_10677);
nor U17499 (N_17499,N_13688,N_10412);
nand U17500 (N_17500,N_12308,N_13840);
nor U17501 (N_17501,N_13879,N_12225);
or U17502 (N_17502,N_13263,N_14940);
nand U17503 (N_17503,N_14950,N_14456);
nor U17504 (N_17504,N_14064,N_11789);
or U17505 (N_17505,N_12246,N_11287);
nor U17506 (N_17506,N_10226,N_11671);
nor U17507 (N_17507,N_12172,N_13957);
nand U17508 (N_17508,N_10857,N_14382);
or U17509 (N_17509,N_12382,N_14787);
nor U17510 (N_17510,N_13162,N_11972);
or U17511 (N_17511,N_14566,N_11728);
nor U17512 (N_17512,N_13311,N_12335);
or U17513 (N_17513,N_11345,N_12150);
or U17514 (N_17514,N_14809,N_14906);
nand U17515 (N_17515,N_13404,N_11740);
xnor U17516 (N_17516,N_12328,N_12447);
nand U17517 (N_17517,N_10148,N_11269);
or U17518 (N_17518,N_14899,N_11985);
or U17519 (N_17519,N_10120,N_14373);
and U17520 (N_17520,N_14129,N_13900);
nand U17521 (N_17521,N_12813,N_14070);
or U17522 (N_17522,N_12135,N_11745);
nor U17523 (N_17523,N_12852,N_13614);
and U17524 (N_17524,N_14819,N_14289);
nor U17525 (N_17525,N_14622,N_11603);
and U17526 (N_17526,N_12736,N_12832);
nand U17527 (N_17527,N_10774,N_12104);
nand U17528 (N_17528,N_13852,N_14984);
nand U17529 (N_17529,N_13045,N_10230);
or U17530 (N_17530,N_11660,N_10980);
nor U17531 (N_17531,N_12187,N_10418);
nor U17532 (N_17532,N_10461,N_13150);
nor U17533 (N_17533,N_10279,N_12606);
nor U17534 (N_17534,N_12441,N_14100);
nand U17535 (N_17535,N_14299,N_10009);
and U17536 (N_17536,N_13300,N_14092);
nand U17537 (N_17537,N_10974,N_11318);
nor U17538 (N_17538,N_10819,N_11446);
or U17539 (N_17539,N_10616,N_13079);
nand U17540 (N_17540,N_10689,N_12790);
nor U17541 (N_17541,N_10666,N_12693);
nand U17542 (N_17542,N_14212,N_13856);
nand U17543 (N_17543,N_12056,N_11279);
nand U17544 (N_17544,N_14571,N_13860);
nor U17545 (N_17545,N_10838,N_13634);
or U17546 (N_17546,N_10295,N_11166);
nand U17547 (N_17547,N_13062,N_14524);
and U17548 (N_17548,N_14496,N_14323);
xnor U17549 (N_17549,N_14815,N_11770);
nor U17550 (N_17550,N_13997,N_11524);
and U17551 (N_17551,N_12979,N_10389);
nor U17552 (N_17552,N_11375,N_10068);
nor U17553 (N_17553,N_10025,N_13018);
or U17554 (N_17554,N_14668,N_14913);
and U17555 (N_17555,N_12226,N_13712);
or U17556 (N_17556,N_12436,N_10325);
nor U17557 (N_17557,N_13687,N_13517);
or U17558 (N_17558,N_12157,N_11198);
nand U17559 (N_17559,N_13423,N_14705);
nand U17560 (N_17560,N_10802,N_13323);
nor U17561 (N_17561,N_10281,N_12925);
nand U17562 (N_17562,N_13981,N_10927);
nor U17563 (N_17563,N_14263,N_13352);
nand U17564 (N_17564,N_11918,N_12588);
and U17565 (N_17565,N_12527,N_13326);
nor U17566 (N_17566,N_13904,N_13562);
or U17567 (N_17567,N_13663,N_12433);
nor U17568 (N_17568,N_11258,N_13825);
nand U17569 (N_17569,N_11495,N_10881);
and U17570 (N_17570,N_11420,N_13872);
nand U17571 (N_17571,N_10335,N_10557);
and U17572 (N_17572,N_14006,N_14845);
xor U17573 (N_17573,N_13722,N_12152);
nand U17574 (N_17574,N_13523,N_14889);
nor U17575 (N_17575,N_12150,N_13846);
and U17576 (N_17576,N_11305,N_10259);
xnor U17577 (N_17577,N_14332,N_10985);
or U17578 (N_17578,N_12800,N_12475);
nand U17579 (N_17579,N_10822,N_13248);
and U17580 (N_17580,N_12649,N_12150);
xor U17581 (N_17581,N_10139,N_12830);
and U17582 (N_17582,N_12614,N_11669);
and U17583 (N_17583,N_14045,N_13882);
nand U17584 (N_17584,N_11439,N_14058);
and U17585 (N_17585,N_12216,N_12497);
nand U17586 (N_17586,N_12435,N_10063);
nor U17587 (N_17587,N_10695,N_11924);
and U17588 (N_17588,N_14903,N_14661);
nor U17589 (N_17589,N_11244,N_13193);
nand U17590 (N_17590,N_14868,N_13893);
and U17591 (N_17591,N_13730,N_14351);
nor U17592 (N_17592,N_12106,N_13939);
and U17593 (N_17593,N_14471,N_12411);
nand U17594 (N_17594,N_12758,N_11628);
or U17595 (N_17595,N_13904,N_12164);
xor U17596 (N_17596,N_13863,N_11533);
nor U17597 (N_17597,N_13664,N_13801);
and U17598 (N_17598,N_13203,N_11382);
or U17599 (N_17599,N_11811,N_13548);
nand U17600 (N_17600,N_10915,N_12044);
and U17601 (N_17601,N_12716,N_11003);
nand U17602 (N_17602,N_11201,N_14454);
nand U17603 (N_17603,N_13357,N_13445);
xnor U17604 (N_17604,N_14674,N_12866);
nor U17605 (N_17605,N_12034,N_10573);
or U17606 (N_17606,N_14592,N_11137);
nand U17607 (N_17607,N_11487,N_12703);
nand U17608 (N_17608,N_14779,N_11793);
nor U17609 (N_17609,N_11894,N_11343);
and U17610 (N_17610,N_11405,N_11683);
and U17611 (N_17611,N_13237,N_12086);
and U17612 (N_17612,N_12757,N_14936);
nand U17613 (N_17613,N_10694,N_11573);
or U17614 (N_17614,N_12034,N_11630);
or U17615 (N_17615,N_10320,N_13399);
and U17616 (N_17616,N_12731,N_13961);
nand U17617 (N_17617,N_10367,N_11460);
nor U17618 (N_17618,N_13688,N_14540);
and U17619 (N_17619,N_11959,N_13784);
nand U17620 (N_17620,N_11108,N_13721);
nand U17621 (N_17621,N_11345,N_10999);
and U17622 (N_17622,N_14378,N_10656);
nor U17623 (N_17623,N_13925,N_12358);
nand U17624 (N_17624,N_11402,N_12778);
and U17625 (N_17625,N_14356,N_10041);
and U17626 (N_17626,N_13283,N_13188);
and U17627 (N_17627,N_13434,N_10570);
or U17628 (N_17628,N_12468,N_14082);
or U17629 (N_17629,N_11920,N_12636);
and U17630 (N_17630,N_10180,N_12521);
nor U17631 (N_17631,N_13507,N_11535);
or U17632 (N_17632,N_11919,N_10312);
and U17633 (N_17633,N_14637,N_10209);
nor U17634 (N_17634,N_13956,N_14256);
and U17635 (N_17635,N_11767,N_12408);
and U17636 (N_17636,N_14676,N_13533);
or U17637 (N_17637,N_10327,N_11177);
nand U17638 (N_17638,N_13153,N_11624);
and U17639 (N_17639,N_13225,N_12866);
and U17640 (N_17640,N_11394,N_13039);
nor U17641 (N_17641,N_13595,N_11228);
nand U17642 (N_17642,N_13199,N_11512);
nor U17643 (N_17643,N_10283,N_14062);
and U17644 (N_17644,N_12121,N_12492);
and U17645 (N_17645,N_11378,N_12941);
and U17646 (N_17646,N_10589,N_10743);
and U17647 (N_17647,N_12284,N_12023);
nor U17648 (N_17648,N_13244,N_14818);
nand U17649 (N_17649,N_13831,N_14092);
nand U17650 (N_17650,N_13025,N_10115);
nand U17651 (N_17651,N_11917,N_13724);
and U17652 (N_17652,N_10565,N_10125);
or U17653 (N_17653,N_13586,N_12344);
nand U17654 (N_17654,N_13342,N_12524);
or U17655 (N_17655,N_10765,N_10072);
or U17656 (N_17656,N_14133,N_11802);
nand U17657 (N_17657,N_11668,N_14808);
nand U17658 (N_17658,N_13989,N_11101);
nor U17659 (N_17659,N_10640,N_13265);
xnor U17660 (N_17660,N_13694,N_14037);
nand U17661 (N_17661,N_11076,N_13727);
and U17662 (N_17662,N_11278,N_13548);
nor U17663 (N_17663,N_10695,N_14083);
or U17664 (N_17664,N_10919,N_14835);
and U17665 (N_17665,N_13537,N_11303);
nor U17666 (N_17666,N_13880,N_10790);
nor U17667 (N_17667,N_10150,N_10576);
nand U17668 (N_17668,N_11359,N_11435);
or U17669 (N_17669,N_12737,N_12447);
and U17670 (N_17670,N_13461,N_10639);
nand U17671 (N_17671,N_12662,N_14465);
nor U17672 (N_17672,N_10331,N_11157);
xnor U17673 (N_17673,N_10305,N_11930);
and U17674 (N_17674,N_11885,N_12905);
and U17675 (N_17675,N_12125,N_12611);
xor U17676 (N_17676,N_11977,N_11405);
and U17677 (N_17677,N_12693,N_11897);
and U17678 (N_17678,N_12154,N_13652);
nor U17679 (N_17679,N_10917,N_11358);
nand U17680 (N_17680,N_12334,N_13300);
xor U17681 (N_17681,N_12970,N_10300);
xnor U17682 (N_17682,N_10487,N_10044);
nand U17683 (N_17683,N_14000,N_13983);
and U17684 (N_17684,N_11310,N_11188);
and U17685 (N_17685,N_14068,N_12923);
nand U17686 (N_17686,N_10013,N_14423);
nor U17687 (N_17687,N_12378,N_11843);
nand U17688 (N_17688,N_13487,N_10579);
and U17689 (N_17689,N_10081,N_13148);
or U17690 (N_17690,N_11694,N_11130);
nand U17691 (N_17691,N_10166,N_12960);
or U17692 (N_17692,N_12464,N_14560);
or U17693 (N_17693,N_11061,N_14223);
nand U17694 (N_17694,N_10305,N_13422);
nor U17695 (N_17695,N_10833,N_11430);
nand U17696 (N_17696,N_13320,N_11541);
or U17697 (N_17697,N_13762,N_14594);
nor U17698 (N_17698,N_10618,N_13775);
or U17699 (N_17699,N_11493,N_13721);
nor U17700 (N_17700,N_10365,N_10079);
nand U17701 (N_17701,N_13366,N_12942);
nand U17702 (N_17702,N_11265,N_13655);
and U17703 (N_17703,N_12906,N_12492);
and U17704 (N_17704,N_12147,N_14073);
nand U17705 (N_17705,N_11420,N_14678);
nand U17706 (N_17706,N_10518,N_14814);
or U17707 (N_17707,N_10922,N_14222);
nor U17708 (N_17708,N_14288,N_12141);
or U17709 (N_17709,N_13063,N_10530);
or U17710 (N_17710,N_11891,N_11393);
xnor U17711 (N_17711,N_11291,N_13512);
nand U17712 (N_17712,N_14470,N_13022);
nand U17713 (N_17713,N_10028,N_14703);
xnor U17714 (N_17714,N_12008,N_11504);
and U17715 (N_17715,N_12595,N_14956);
nor U17716 (N_17716,N_13170,N_13374);
and U17717 (N_17717,N_14940,N_13884);
or U17718 (N_17718,N_12803,N_14300);
or U17719 (N_17719,N_13003,N_14540);
nor U17720 (N_17720,N_10848,N_14714);
xor U17721 (N_17721,N_14231,N_14453);
nand U17722 (N_17722,N_10827,N_10976);
and U17723 (N_17723,N_13533,N_13789);
xor U17724 (N_17724,N_12688,N_10738);
xor U17725 (N_17725,N_11720,N_12335);
or U17726 (N_17726,N_14281,N_14340);
nand U17727 (N_17727,N_13597,N_14730);
and U17728 (N_17728,N_14314,N_10424);
nor U17729 (N_17729,N_10289,N_14072);
or U17730 (N_17730,N_10378,N_14704);
or U17731 (N_17731,N_10664,N_13141);
or U17732 (N_17732,N_13352,N_13293);
nand U17733 (N_17733,N_13383,N_12633);
nand U17734 (N_17734,N_14700,N_14395);
and U17735 (N_17735,N_14383,N_13659);
or U17736 (N_17736,N_11805,N_13659);
and U17737 (N_17737,N_12050,N_10367);
xnor U17738 (N_17738,N_13704,N_13453);
xnor U17739 (N_17739,N_10940,N_10316);
or U17740 (N_17740,N_12085,N_10764);
xor U17741 (N_17741,N_13273,N_14173);
or U17742 (N_17742,N_10494,N_13494);
and U17743 (N_17743,N_13786,N_14793);
or U17744 (N_17744,N_12995,N_12484);
and U17745 (N_17745,N_12461,N_12837);
nor U17746 (N_17746,N_10816,N_11320);
nor U17747 (N_17747,N_11198,N_14630);
or U17748 (N_17748,N_13113,N_14664);
or U17749 (N_17749,N_11065,N_10039);
or U17750 (N_17750,N_12217,N_12845);
and U17751 (N_17751,N_11299,N_10169);
and U17752 (N_17752,N_10846,N_11814);
or U17753 (N_17753,N_11925,N_14781);
nand U17754 (N_17754,N_14942,N_10485);
or U17755 (N_17755,N_14878,N_11711);
and U17756 (N_17756,N_10900,N_14777);
or U17757 (N_17757,N_12030,N_12876);
nor U17758 (N_17758,N_11349,N_14374);
nand U17759 (N_17759,N_12480,N_14798);
xor U17760 (N_17760,N_10465,N_13353);
nor U17761 (N_17761,N_13410,N_10155);
nor U17762 (N_17762,N_14938,N_10619);
or U17763 (N_17763,N_11832,N_13491);
or U17764 (N_17764,N_12220,N_12676);
nor U17765 (N_17765,N_10121,N_14620);
or U17766 (N_17766,N_11953,N_12068);
nor U17767 (N_17767,N_14665,N_13503);
nor U17768 (N_17768,N_12571,N_12426);
nor U17769 (N_17769,N_13433,N_10585);
and U17770 (N_17770,N_14830,N_13674);
or U17771 (N_17771,N_10830,N_14724);
and U17772 (N_17772,N_11603,N_12307);
and U17773 (N_17773,N_13353,N_14352);
nor U17774 (N_17774,N_12521,N_11374);
or U17775 (N_17775,N_12894,N_10814);
nand U17776 (N_17776,N_14498,N_13967);
or U17777 (N_17777,N_13331,N_12568);
or U17778 (N_17778,N_14815,N_11181);
nor U17779 (N_17779,N_10574,N_14129);
xnor U17780 (N_17780,N_11495,N_10222);
and U17781 (N_17781,N_13374,N_14450);
or U17782 (N_17782,N_10830,N_10477);
xor U17783 (N_17783,N_13737,N_12167);
nor U17784 (N_17784,N_14308,N_11601);
nor U17785 (N_17785,N_13588,N_12706);
and U17786 (N_17786,N_12845,N_12063);
or U17787 (N_17787,N_10387,N_12208);
nand U17788 (N_17788,N_10290,N_12873);
or U17789 (N_17789,N_10064,N_10961);
and U17790 (N_17790,N_10371,N_10368);
nand U17791 (N_17791,N_14726,N_13717);
nor U17792 (N_17792,N_11191,N_10628);
nand U17793 (N_17793,N_12427,N_14254);
nor U17794 (N_17794,N_11305,N_11419);
or U17795 (N_17795,N_12719,N_14618);
nor U17796 (N_17796,N_11117,N_10774);
and U17797 (N_17797,N_12593,N_10445);
nor U17798 (N_17798,N_13026,N_11858);
or U17799 (N_17799,N_12720,N_11908);
xor U17800 (N_17800,N_12855,N_10981);
and U17801 (N_17801,N_10273,N_10693);
nand U17802 (N_17802,N_10757,N_13112);
nor U17803 (N_17803,N_11494,N_12882);
nor U17804 (N_17804,N_12331,N_14856);
or U17805 (N_17805,N_12209,N_10088);
or U17806 (N_17806,N_12048,N_12142);
nand U17807 (N_17807,N_10753,N_13229);
nor U17808 (N_17808,N_12433,N_13443);
nand U17809 (N_17809,N_14695,N_13871);
and U17810 (N_17810,N_12294,N_11583);
nor U17811 (N_17811,N_12373,N_12391);
and U17812 (N_17812,N_11772,N_11532);
and U17813 (N_17813,N_13835,N_10282);
or U17814 (N_17814,N_14065,N_13261);
nand U17815 (N_17815,N_12392,N_14690);
nor U17816 (N_17816,N_10146,N_11155);
or U17817 (N_17817,N_12623,N_10754);
nand U17818 (N_17818,N_13864,N_14563);
nand U17819 (N_17819,N_13571,N_11288);
and U17820 (N_17820,N_13560,N_13827);
or U17821 (N_17821,N_12010,N_12346);
or U17822 (N_17822,N_13484,N_14031);
and U17823 (N_17823,N_11055,N_12331);
and U17824 (N_17824,N_14202,N_13884);
nor U17825 (N_17825,N_14645,N_14599);
xnor U17826 (N_17826,N_11958,N_12544);
and U17827 (N_17827,N_12516,N_10595);
and U17828 (N_17828,N_13331,N_10440);
nor U17829 (N_17829,N_14995,N_13840);
nand U17830 (N_17830,N_11360,N_14679);
and U17831 (N_17831,N_12189,N_14636);
xnor U17832 (N_17832,N_12311,N_11254);
nor U17833 (N_17833,N_11852,N_14142);
nand U17834 (N_17834,N_14449,N_10486);
and U17835 (N_17835,N_14224,N_14169);
nor U17836 (N_17836,N_14000,N_14023);
nand U17837 (N_17837,N_11895,N_12607);
nand U17838 (N_17838,N_12263,N_11007);
nor U17839 (N_17839,N_13976,N_10994);
nor U17840 (N_17840,N_12481,N_10740);
and U17841 (N_17841,N_13790,N_13204);
or U17842 (N_17842,N_10153,N_14289);
and U17843 (N_17843,N_10071,N_11648);
nor U17844 (N_17844,N_13091,N_11375);
nand U17845 (N_17845,N_13807,N_14298);
nor U17846 (N_17846,N_13958,N_14255);
and U17847 (N_17847,N_12461,N_11286);
nor U17848 (N_17848,N_12288,N_13366);
and U17849 (N_17849,N_11244,N_10883);
or U17850 (N_17850,N_14264,N_13264);
nor U17851 (N_17851,N_14615,N_10677);
and U17852 (N_17852,N_13232,N_10451);
or U17853 (N_17853,N_12958,N_12083);
nand U17854 (N_17854,N_14753,N_11869);
and U17855 (N_17855,N_12187,N_13731);
nor U17856 (N_17856,N_10238,N_10862);
nor U17857 (N_17857,N_11493,N_11102);
or U17858 (N_17858,N_13242,N_13869);
nand U17859 (N_17859,N_11357,N_13573);
and U17860 (N_17860,N_12739,N_10043);
and U17861 (N_17861,N_12999,N_12250);
nand U17862 (N_17862,N_12210,N_14895);
xnor U17863 (N_17863,N_11397,N_11527);
nor U17864 (N_17864,N_13015,N_11329);
and U17865 (N_17865,N_13236,N_13785);
nand U17866 (N_17866,N_13221,N_13267);
nand U17867 (N_17867,N_10924,N_14503);
nor U17868 (N_17868,N_13324,N_12317);
nor U17869 (N_17869,N_10406,N_11755);
and U17870 (N_17870,N_11242,N_13051);
and U17871 (N_17871,N_13841,N_14010);
nand U17872 (N_17872,N_10651,N_14321);
and U17873 (N_17873,N_12290,N_13357);
and U17874 (N_17874,N_13271,N_10628);
and U17875 (N_17875,N_12341,N_14425);
nor U17876 (N_17876,N_10285,N_10728);
or U17877 (N_17877,N_14808,N_11613);
or U17878 (N_17878,N_10221,N_13787);
xor U17879 (N_17879,N_12988,N_12120);
or U17880 (N_17880,N_11114,N_10487);
nor U17881 (N_17881,N_13020,N_14620);
nor U17882 (N_17882,N_13422,N_10486);
and U17883 (N_17883,N_11997,N_11628);
nor U17884 (N_17884,N_10285,N_11058);
nor U17885 (N_17885,N_14730,N_12462);
nand U17886 (N_17886,N_10626,N_11550);
or U17887 (N_17887,N_14362,N_12772);
or U17888 (N_17888,N_10306,N_14976);
or U17889 (N_17889,N_11325,N_13365);
and U17890 (N_17890,N_14229,N_13026);
or U17891 (N_17891,N_12409,N_10624);
and U17892 (N_17892,N_14992,N_10505);
nor U17893 (N_17893,N_13198,N_12992);
nor U17894 (N_17894,N_14442,N_10064);
nor U17895 (N_17895,N_13812,N_10159);
nand U17896 (N_17896,N_13099,N_13163);
or U17897 (N_17897,N_13495,N_11409);
and U17898 (N_17898,N_12539,N_13339);
and U17899 (N_17899,N_11858,N_10927);
nor U17900 (N_17900,N_13631,N_12268);
nand U17901 (N_17901,N_10854,N_14991);
or U17902 (N_17902,N_12161,N_14880);
nor U17903 (N_17903,N_12396,N_14551);
nand U17904 (N_17904,N_12817,N_14080);
and U17905 (N_17905,N_10169,N_12166);
or U17906 (N_17906,N_12112,N_13636);
or U17907 (N_17907,N_13625,N_10259);
and U17908 (N_17908,N_11114,N_10823);
nor U17909 (N_17909,N_11422,N_10252);
nor U17910 (N_17910,N_13922,N_12869);
nand U17911 (N_17911,N_12791,N_11344);
nand U17912 (N_17912,N_13942,N_11713);
nand U17913 (N_17913,N_12760,N_10614);
or U17914 (N_17914,N_12826,N_11512);
nand U17915 (N_17915,N_14140,N_12769);
nand U17916 (N_17916,N_10022,N_12929);
nand U17917 (N_17917,N_12687,N_11476);
nand U17918 (N_17918,N_13488,N_12686);
nor U17919 (N_17919,N_13116,N_10838);
nand U17920 (N_17920,N_12124,N_11277);
nor U17921 (N_17921,N_12265,N_14385);
or U17922 (N_17922,N_13773,N_14568);
or U17923 (N_17923,N_11122,N_14703);
nand U17924 (N_17924,N_14962,N_10284);
nor U17925 (N_17925,N_12598,N_13680);
or U17926 (N_17926,N_12472,N_14437);
and U17927 (N_17927,N_10990,N_10643);
xor U17928 (N_17928,N_11450,N_14089);
xor U17929 (N_17929,N_12640,N_12084);
nor U17930 (N_17930,N_14864,N_10401);
nor U17931 (N_17931,N_10076,N_14085);
and U17932 (N_17932,N_13242,N_10692);
nand U17933 (N_17933,N_11132,N_10918);
xor U17934 (N_17934,N_11592,N_11000);
xor U17935 (N_17935,N_12637,N_12686);
and U17936 (N_17936,N_14280,N_11583);
nor U17937 (N_17937,N_12640,N_11446);
nand U17938 (N_17938,N_12007,N_14052);
and U17939 (N_17939,N_12168,N_12247);
nand U17940 (N_17940,N_10437,N_11263);
and U17941 (N_17941,N_12109,N_11080);
nand U17942 (N_17942,N_10955,N_12091);
xnor U17943 (N_17943,N_13307,N_11856);
or U17944 (N_17944,N_11776,N_12310);
and U17945 (N_17945,N_13374,N_11113);
and U17946 (N_17946,N_13100,N_11577);
or U17947 (N_17947,N_11377,N_13648);
nor U17948 (N_17948,N_13974,N_12020);
and U17949 (N_17949,N_11386,N_12294);
or U17950 (N_17950,N_14544,N_14189);
nor U17951 (N_17951,N_10284,N_11696);
nand U17952 (N_17952,N_13189,N_12653);
xor U17953 (N_17953,N_13273,N_10747);
nand U17954 (N_17954,N_11794,N_14920);
nor U17955 (N_17955,N_11197,N_12837);
xor U17956 (N_17956,N_14517,N_12268);
or U17957 (N_17957,N_12253,N_13364);
or U17958 (N_17958,N_12161,N_14821);
and U17959 (N_17959,N_10620,N_13545);
or U17960 (N_17960,N_11123,N_12533);
and U17961 (N_17961,N_12351,N_13520);
nand U17962 (N_17962,N_12436,N_12667);
nor U17963 (N_17963,N_12713,N_14259);
or U17964 (N_17964,N_10859,N_12096);
nand U17965 (N_17965,N_10782,N_11061);
and U17966 (N_17966,N_13588,N_10178);
nor U17967 (N_17967,N_14421,N_11902);
nand U17968 (N_17968,N_12477,N_11284);
and U17969 (N_17969,N_11682,N_11633);
and U17970 (N_17970,N_11572,N_11991);
or U17971 (N_17971,N_12912,N_11648);
nand U17972 (N_17972,N_11620,N_14507);
or U17973 (N_17973,N_13942,N_10540);
and U17974 (N_17974,N_10733,N_13313);
nand U17975 (N_17975,N_10161,N_10568);
and U17976 (N_17976,N_10851,N_11717);
xnor U17977 (N_17977,N_13319,N_14239);
nor U17978 (N_17978,N_11216,N_13756);
nor U17979 (N_17979,N_10151,N_10910);
or U17980 (N_17980,N_11183,N_11522);
nor U17981 (N_17981,N_13370,N_13488);
nand U17982 (N_17982,N_14852,N_11155);
nor U17983 (N_17983,N_11582,N_13324);
and U17984 (N_17984,N_13301,N_11010);
or U17985 (N_17985,N_13296,N_12450);
nand U17986 (N_17986,N_12439,N_13480);
nor U17987 (N_17987,N_13613,N_14079);
and U17988 (N_17988,N_10643,N_13341);
or U17989 (N_17989,N_11379,N_14491);
nand U17990 (N_17990,N_12882,N_14150);
nand U17991 (N_17991,N_12046,N_10462);
xnor U17992 (N_17992,N_10968,N_13781);
or U17993 (N_17993,N_13941,N_10091);
or U17994 (N_17994,N_10684,N_10207);
nand U17995 (N_17995,N_13339,N_12534);
or U17996 (N_17996,N_12391,N_12980);
and U17997 (N_17997,N_13254,N_10385);
or U17998 (N_17998,N_10911,N_10243);
and U17999 (N_17999,N_12644,N_13470);
nand U18000 (N_18000,N_10959,N_10184);
nor U18001 (N_18001,N_11348,N_12377);
xor U18002 (N_18002,N_14950,N_10133);
nor U18003 (N_18003,N_14556,N_11239);
xnor U18004 (N_18004,N_13155,N_10384);
nor U18005 (N_18005,N_12396,N_13910);
and U18006 (N_18006,N_10868,N_14123);
nor U18007 (N_18007,N_14854,N_12479);
or U18008 (N_18008,N_14743,N_13604);
and U18009 (N_18009,N_14463,N_14858);
and U18010 (N_18010,N_11438,N_13623);
or U18011 (N_18011,N_10597,N_14434);
or U18012 (N_18012,N_14766,N_10386);
nand U18013 (N_18013,N_12730,N_10061);
nand U18014 (N_18014,N_10638,N_12747);
nor U18015 (N_18015,N_10380,N_11471);
or U18016 (N_18016,N_10414,N_14094);
nor U18017 (N_18017,N_14369,N_11812);
nor U18018 (N_18018,N_12077,N_10829);
nor U18019 (N_18019,N_14401,N_11135);
nor U18020 (N_18020,N_10098,N_13997);
nor U18021 (N_18021,N_11344,N_12451);
nand U18022 (N_18022,N_11533,N_11545);
nand U18023 (N_18023,N_11569,N_10971);
or U18024 (N_18024,N_10653,N_11483);
and U18025 (N_18025,N_12387,N_13064);
nor U18026 (N_18026,N_12555,N_10991);
and U18027 (N_18027,N_10485,N_11316);
or U18028 (N_18028,N_12993,N_13917);
or U18029 (N_18029,N_12558,N_13346);
nor U18030 (N_18030,N_10117,N_10720);
nand U18031 (N_18031,N_11172,N_11765);
and U18032 (N_18032,N_13094,N_13499);
or U18033 (N_18033,N_13359,N_13954);
or U18034 (N_18034,N_13077,N_10226);
nor U18035 (N_18035,N_13715,N_12580);
or U18036 (N_18036,N_11697,N_14800);
and U18037 (N_18037,N_10279,N_10543);
nand U18038 (N_18038,N_11534,N_14423);
nor U18039 (N_18039,N_11064,N_10433);
and U18040 (N_18040,N_10318,N_13023);
nor U18041 (N_18041,N_11742,N_14646);
or U18042 (N_18042,N_10543,N_12371);
nand U18043 (N_18043,N_13144,N_10101);
or U18044 (N_18044,N_14479,N_11123);
nor U18045 (N_18045,N_11220,N_13315);
xor U18046 (N_18046,N_14918,N_10036);
or U18047 (N_18047,N_13589,N_11255);
xnor U18048 (N_18048,N_11471,N_10840);
and U18049 (N_18049,N_12662,N_12317);
nor U18050 (N_18050,N_11604,N_14376);
nor U18051 (N_18051,N_12921,N_10661);
nand U18052 (N_18052,N_13402,N_14500);
nand U18053 (N_18053,N_12233,N_10868);
nor U18054 (N_18054,N_12344,N_10344);
and U18055 (N_18055,N_11228,N_10139);
and U18056 (N_18056,N_11434,N_11373);
and U18057 (N_18057,N_12399,N_14081);
nand U18058 (N_18058,N_10080,N_11255);
nor U18059 (N_18059,N_11178,N_13137);
and U18060 (N_18060,N_11615,N_14680);
and U18061 (N_18061,N_10714,N_13590);
and U18062 (N_18062,N_10254,N_12007);
xor U18063 (N_18063,N_13177,N_13063);
and U18064 (N_18064,N_11950,N_11296);
xnor U18065 (N_18065,N_12749,N_14782);
nand U18066 (N_18066,N_11421,N_11055);
nor U18067 (N_18067,N_13649,N_12133);
nor U18068 (N_18068,N_12662,N_11163);
or U18069 (N_18069,N_11237,N_13607);
nor U18070 (N_18070,N_12817,N_10390);
and U18071 (N_18071,N_14216,N_13801);
nand U18072 (N_18072,N_13769,N_13094);
and U18073 (N_18073,N_11387,N_10529);
and U18074 (N_18074,N_14053,N_11659);
xnor U18075 (N_18075,N_11031,N_11512);
nand U18076 (N_18076,N_14127,N_13754);
xor U18077 (N_18077,N_10171,N_10999);
nor U18078 (N_18078,N_13909,N_10357);
nor U18079 (N_18079,N_12335,N_10065);
and U18080 (N_18080,N_12781,N_13920);
and U18081 (N_18081,N_11302,N_13802);
nor U18082 (N_18082,N_14211,N_10902);
nand U18083 (N_18083,N_10610,N_12940);
and U18084 (N_18084,N_10069,N_10041);
or U18085 (N_18085,N_13809,N_13911);
and U18086 (N_18086,N_14778,N_10581);
nand U18087 (N_18087,N_10892,N_13909);
nor U18088 (N_18088,N_14493,N_11367);
nor U18089 (N_18089,N_10764,N_11199);
and U18090 (N_18090,N_14724,N_10945);
nor U18091 (N_18091,N_14973,N_14103);
nor U18092 (N_18092,N_10612,N_10793);
or U18093 (N_18093,N_13448,N_12469);
xnor U18094 (N_18094,N_14998,N_11506);
nand U18095 (N_18095,N_13508,N_11107);
or U18096 (N_18096,N_12027,N_13391);
and U18097 (N_18097,N_10595,N_12405);
nor U18098 (N_18098,N_10638,N_13045);
and U18099 (N_18099,N_14621,N_10409);
xnor U18100 (N_18100,N_14058,N_10293);
and U18101 (N_18101,N_10271,N_11660);
or U18102 (N_18102,N_10379,N_10317);
nor U18103 (N_18103,N_10989,N_13673);
and U18104 (N_18104,N_11124,N_14003);
or U18105 (N_18105,N_14142,N_13352);
and U18106 (N_18106,N_13266,N_11375);
and U18107 (N_18107,N_12130,N_13418);
nor U18108 (N_18108,N_14657,N_12674);
xor U18109 (N_18109,N_11844,N_12893);
nand U18110 (N_18110,N_12052,N_13613);
nand U18111 (N_18111,N_12828,N_14670);
or U18112 (N_18112,N_13042,N_12237);
or U18113 (N_18113,N_13672,N_10628);
nor U18114 (N_18114,N_11540,N_14244);
nor U18115 (N_18115,N_14340,N_13143);
nor U18116 (N_18116,N_13264,N_14407);
or U18117 (N_18117,N_13542,N_10347);
nor U18118 (N_18118,N_13212,N_13645);
or U18119 (N_18119,N_10987,N_12385);
nand U18120 (N_18120,N_14962,N_11153);
or U18121 (N_18121,N_13951,N_14310);
nor U18122 (N_18122,N_12944,N_10821);
and U18123 (N_18123,N_14038,N_12630);
nand U18124 (N_18124,N_11075,N_14166);
or U18125 (N_18125,N_12552,N_14680);
nand U18126 (N_18126,N_10237,N_13384);
xnor U18127 (N_18127,N_13936,N_13111);
nand U18128 (N_18128,N_13054,N_10528);
or U18129 (N_18129,N_12080,N_13362);
or U18130 (N_18130,N_10874,N_14362);
and U18131 (N_18131,N_10104,N_14169);
xor U18132 (N_18132,N_14881,N_14969);
xor U18133 (N_18133,N_14392,N_10126);
nor U18134 (N_18134,N_13809,N_12477);
nand U18135 (N_18135,N_12319,N_12286);
nand U18136 (N_18136,N_11799,N_14161);
nand U18137 (N_18137,N_10123,N_12901);
or U18138 (N_18138,N_14639,N_10022);
nor U18139 (N_18139,N_13526,N_12352);
or U18140 (N_18140,N_14637,N_12842);
and U18141 (N_18141,N_10122,N_10761);
nand U18142 (N_18142,N_11184,N_10132);
and U18143 (N_18143,N_13758,N_13389);
xnor U18144 (N_18144,N_12380,N_12641);
or U18145 (N_18145,N_13425,N_14012);
xnor U18146 (N_18146,N_10805,N_14646);
nor U18147 (N_18147,N_11868,N_14581);
nand U18148 (N_18148,N_12813,N_11339);
nor U18149 (N_18149,N_12941,N_13481);
xor U18150 (N_18150,N_10218,N_11838);
nor U18151 (N_18151,N_13938,N_11763);
nand U18152 (N_18152,N_11647,N_13216);
and U18153 (N_18153,N_13301,N_11580);
or U18154 (N_18154,N_10503,N_13700);
and U18155 (N_18155,N_12330,N_11687);
nor U18156 (N_18156,N_12860,N_13476);
and U18157 (N_18157,N_12848,N_12968);
nand U18158 (N_18158,N_14351,N_14263);
nand U18159 (N_18159,N_10791,N_11807);
and U18160 (N_18160,N_12856,N_13716);
or U18161 (N_18161,N_13284,N_13739);
or U18162 (N_18162,N_12482,N_14871);
nor U18163 (N_18163,N_14284,N_12488);
and U18164 (N_18164,N_13059,N_10079);
xnor U18165 (N_18165,N_14658,N_11406);
xnor U18166 (N_18166,N_11471,N_11028);
and U18167 (N_18167,N_12352,N_13556);
nand U18168 (N_18168,N_11436,N_14838);
nor U18169 (N_18169,N_13943,N_14296);
nor U18170 (N_18170,N_11571,N_10249);
or U18171 (N_18171,N_14109,N_10142);
nor U18172 (N_18172,N_12490,N_10398);
or U18173 (N_18173,N_12893,N_10019);
or U18174 (N_18174,N_14228,N_12166);
nor U18175 (N_18175,N_14843,N_11411);
or U18176 (N_18176,N_13232,N_11966);
nand U18177 (N_18177,N_10628,N_11626);
nand U18178 (N_18178,N_11330,N_13546);
nand U18179 (N_18179,N_14789,N_10322);
and U18180 (N_18180,N_12388,N_12532);
or U18181 (N_18181,N_10210,N_14249);
nor U18182 (N_18182,N_11474,N_10703);
nand U18183 (N_18183,N_12632,N_11828);
or U18184 (N_18184,N_11775,N_12371);
nor U18185 (N_18185,N_13164,N_13212);
or U18186 (N_18186,N_14006,N_13623);
or U18187 (N_18187,N_10217,N_13253);
or U18188 (N_18188,N_12381,N_12005);
nand U18189 (N_18189,N_10810,N_12786);
or U18190 (N_18190,N_14376,N_11940);
xnor U18191 (N_18191,N_12557,N_14235);
and U18192 (N_18192,N_10340,N_12827);
nor U18193 (N_18193,N_13755,N_13194);
and U18194 (N_18194,N_10947,N_14265);
nand U18195 (N_18195,N_13516,N_11286);
and U18196 (N_18196,N_11796,N_14519);
or U18197 (N_18197,N_14576,N_14949);
nor U18198 (N_18198,N_10466,N_11878);
nand U18199 (N_18199,N_14849,N_10025);
nand U18200 (N_18200,N_10231,N_13111);
nand U18201 (N_18201,N_10071,N_14665);
or U18202 (N_18202,N_10635,N_14895);
xor U18203 (N_18203,N_11238,N_10150);
xnor U18204 (N_18204,N_14975,N_14967);
xor U18205 (N_18205,N_14224,N_14011);
xnor U18206 (N_18206,N_10549,N_12717);
nor U18207 (N_18207,N_13044,N_11408);
nand U18208 (N_18208,N_11286,N_12880);
xnor U18209 (N_18209,N_13308,N_13598);
nand U18210 (N_18210,N_14759,N_10374);
nor U18211 (N_18211,N_10289,N_12773);
xor U18212 (N_18212,N_12777,N_13942);
nand U18213 (N_18213,N_10078,N_10977);
nor U18214 (N_18214,N_12699,N_11882);
nor U18215 (N_18215,N_12531,N_12980);
nor U18216 (N_18216,N_10522,N_11188);
nor U18217 (N_18217,N_13566,N_14025);
nor U18218 (N_18218,N_12037,N_12086);
nor U18219 (N_18219,N_10404,N_11626);
nand U18220 (N_18220,N_10448,N_10253);
nor U18221 (N_18221,N_14922,N_13075);
nor U18222 (N_18222,N_13114,N_10994);
and U18223 (N_18223,N_14899,N_10580);
nor U18224 (N_18224,N_11787,N_10503);
nor U18225 (N_18225,N_11755,N_10911);
xor U18226 (N_18226,N_14916,N_10387);
nand U18227 (N_18227,N_12961,N_14030);
and U18228 (N_18228,N_11639,N_12157);
nand U18229 (N_18229,N_11710,N_12156);
and U18230 (N_18230,N_13600,N_14020);
and U18231 (N_18231,N_14846,N_11314);
nand U18232 (N_18232,N_12771,N_14311);
and U18233 (N_18233,N_13930,N_11048);
nand U18234 (N_18234,N_12593,N_13193);
nor U18235 (N_18235,N_12082,N_13701);
nand U18236 (N_18236,N_11706,N_10467);
nor U18237 (N_18237,N_12717,N_12819);
nor U18238 (N_18238,N_14801,N_10401);
and U18239 (N_18239,N_10438,N_11209);
nor U18240 (N_18240,N_14348,N_13957);
nand U18241 (N_18241,N_10369,N_11306);
nand U18242 (N_18242,N_13874,N_13229);
and U18243 (N_18243,N_14621,N_13491);
or U18244 (N_18244,N_12726,N_12071);
nor U18245 (N_18245,N_12888,N_11934);
nand U18246 (N_18246,N_12205,N_10287);
nand U18247 (N_18247,N_13376,N_13564);
or U18248 (N_18248,N_12837,N_12029);
nor U18249 (N_18249,N_12265,N_12237);
or U18250 (N_18250,N_10693,N_14978);
or U18251 (N_18251,N_13317,N_11613);
xor U18252 (N_18252,N_12593,N_10425);
xor U18253 (N_18253,N_13677,N_13984);
and U18254 (N_18254,N_13042,N_11075);
or U18255 (N_18255,N_11895,N_10120);
nor U18256 (N_18256,N_13273,N_11279);
nor U18257 (N_18257,N_12908,N_10696);
and U18258 (N_18258,N_14870,N_14544);
and U18259 (N_18259,N_13683,N_11079);
or U18260 (N_18260,N_12365,N_12105);
or U18261 (N_18261,N_11166,N_11061);
and U18262 (N_18262,N_11925,N_11172);
nor U18263 (N_18263,N_14101,N_13597);
nand U18264 (N_18264,N_14037,N_10332);
or U18265 (N_18265,N_13160,N_12113);
and U18266 (N_18266,N_12612,N_10430);
and U18267 (N_18267,N_11372,N_12287);
nand U18268 (N_18268,N_11111,N_10799);
and U18269 (N_18269,N_11863,N_13847);
and U18270 (N_18270,N_14427,N_12253);
nor U18271 (N_18271,N_11966,N_12851);
nand U18272 (N_18272,N_14425,N_12514);
nor U18273 (N_18273,N_12268,N_13362);
xor U18274 (N_18274,N_14159,N_10302);
or U18275 (N_18275,N_13454,N_14295);
xnor U18276 (N_18276,N_12297,N_11081);
nand U18277 (N_18277,N_10507,N_10066);
nand U18278 (N_18278,N_11711,N_10629);
or U18279 (N_18279,N_11158,N_14444);
or U18280 (N_18280,N_12084,N_13542);
nor U18281 (N_18281,N_14245,N_11845);
xor U18282 (N_18282,N_12419,N_11024);
xnor U18283 (N_18283,N_10849,N_13761);
or U18284 (N_18284,N_10356,N_11999);
and U18285 (N_18285,N_12596,N_12087);
nor U18286 (N_18286,N_12260,N_11227);
nor U18287 (N_18287,N_11825,N_11620);
nor U18288 (N_18288,N_12039,N_13804);
xnor U18289 (N_18289,N_13856,N_12912);
or U18290 (N_18290,N_10198,N_11604);
nor U18291 (N_18291,N_11261,N_11779);
and U18292 (N_18292,N_11189,N_14584);
nor U18293 (N_18293,N_12206,N_13026);
xor U18294 (N_18294,N_10101,N_13466);
nand U18295 (N_18295,N_14310,N_13394);
nor U18296 (N_18296,N_14907,N_11357);
and U18297 (N_18297,N_10565,N_10991);
nand U18298 (N_18298,N_11592,N_14501);
or U18299 (N_18299,N_10764,N_12484);
xnor U18300 (N_18300,N_10868,N_10308);
nand U18301 (N_18301,N_10898,N_11727);
nor U18302 (N_18302,N_10672,N_11030);
nor U18303 (N_18303,N_11170,N_12300);
nand U18304 (N_18304,N_10970,N_10866);
xor U18305 (N_18305,N_11112,N_11641);
xor U18306 (N_18306,N_13767,N_12432);
and U18307 (N_18307,N_12740,N_10883);
xnor U18308 (N_18308,N_12976,N_12357);
and U18309 (N_18309,N_13626,N_13650);
nor U18310 (N_18310,N_13350,N_13451);
or U18311 (N_18311,N_14965,N_11656);
or U18312 (N_18312,N_14638,N_12107);
nand U18313 (N_18313,N_10753,N_14982);
or U18314 (N_18314,N_11545,N_14186);
nor U18315 (N_18315,N_13823,N_11986);
nor U18316 (N_18316,N_14263,N_13595);
and U18317 (N_18317,N_10488,N_12545);
or U18318 (N_18318,N_12494,N_11634);
and U18319 (N_18319,N_12631,N_14753);
nor U18320 (N_18320,N_10749,N_13080);
and U18321 (N_18321,N_12060,N_14276);
nand U18322 (N_18322,N_10742,N_11398);
nand U18323 (N_18323,N_12157,N_14806);
nor U18324 (N_18324,N_13157,N_12475);
nand U18325 (N_18325,N_14353,N_11455);
xnor U18326 (N_18326,N_10844,N_13404);
or U18327 (N_18327,N_13787,N_13582);
nor U18328 (N_18328,N_10105,N_10048);
nand U18329 (N_18329,N_13528,N_11524);
or U18330 (N_18330,N_14974,N_12812);
nor U18331 (N_18331,N_10390,N_14413);
and U18332 (N_18332,N_12749,N_13286);
xnor U18333 (N_18333,N_10554,N_10102);
or U18334 (N_18334,N_13850,N_10973);
nor U18335 (N_18335,N_14203,N_14651);
or U18336 (N_18336,N_14647,N_13684);
nand U18337 (N_18337,N_14695,N_12678);
and U18338 (N_18338,N_12615,N_12957);
or U18339 (N_18339,N_14472,N_10698);
or U18340 (N_18340,N_11824,N_10228);
or U18341 (N_18341,N_10068,N_14305);
and U18342 (N_18342,N_14351,N_14819);
nor U18343 (N_18343,N_13313,N_13575);
or U18344 (N_18344,N_14648,N_12248);
nand U18345 (N_18345,N_13125,N_10503);
nand U18346 (N_18346,N_14507,N_13780);
and U18347 (N_18347,N_13841,N_14417);
nor U18348 (N_18348,N_14456,N_12771);
and U18349 (N_18349,N_10214,N_12591);
nor U18350 (N_18350,N_14545,N_11000);
or U18351 (N_18351,N_14148,N_11679);
and U18352 (N_18352,N_13160,N_14338);
and U18353 (N_18353,N_14610,N_14883);
nor U18354 (N_18354,N_11854,N_10461);
xor U18355 (N_18355,N_13295,N_11919);
or U18356 (N_18356,N_13199,N_12697);
nand U18357 (N_18357,N_14835,N_12233);
nand U18358 (N_18358,N_10318,N_14079);
and U18359 (N_18359,N_10909,N_12540);
and U18360 (N_18360,N_10253,N_14675);
and U18361 (N_18361,N_11895,N_12089);
nand U18362 (N_18362,N_12230,N_10296);
and U18363 (N_18363,N_12167,N_13685);
or U18364 (N_18364,N_11427,N_11918);
xnor U18365 (N_18365,N_10907,N_11140);
or U18366 (N_18366,N_10243,N_11336);
nand U18367 (N_18367,N_11297,N_10571);
or U18368 (N_18368,N_10313,N_13917);
and U18369 (N_18369,N_11263,N_10119);
xor U18370 (N_18370,N_13339,N_13909);
nor U18371 (N_18371,N_13315,N_10491);
or U18372 (N_18372,N_14739,N_12149);
or U18373 (N_18373,N_11918,N_10022);
nor U18374 (N_18374,N_12801,N_14043);
and U18375 (N_18375,N_10085,N_13750);
and U18376 (N_18376,N_12974,N_12215);
xor U18377 (N_18377,N_14486,N_10376);
and U18378 (N_18378,N_12840,N_12860);
nand U18379 (N_18379,N_12966,N_10306);
nand U18380 (N_18380,N_11063,N_10612);
or U18381 (N_18381,N_13229,N_14026);
and U18382 (N_18382,N_12841,N_11683);
or U18383 (N_18383,N_13565,N_12022);
or U18384 (N_18384,N_12453,N_12174);
and U18385 (N_18385,N_11104,N_13761);
nor U18386 (N_18386,N_10527,N_14624);
nor U18387 (N_18387,N_14892,N_14799);
or U18388 (N_18388,N_12010,N_11185);
nand U18389 (N_18389,N_13937,N_10432);
nor U18390 (N_18390,N_10794,N_12668);
and U18391 (N_18391,N_11202,N_12776);
nand U18392 (N_18392,N_12189,N_13122);
xnor U18393 (N_18393,N_14532,N_11722);
nand U18394 (N_18394,N_13366,N_14546);
nand U18395 (N_18395,N_11887,N_13102);
nand U18396 (N_18396,N_14988,N_14279);
or U18397 (N_18397,N_12909,N_11128);
nand U18398 (N_18398,N_11074,N_13144);
and U18399 (N_18399,N_11128,N_12607);
and U18400 (N_18400,N_10972,N_13332);
nand U18401 (N_18401,N_12423,N_10984);
nor U18402 (N_18402,N_10096,N_11859);
nand U18403 (N_18403,N_13911,N_12982);
and U18404 (N_18404,N_12193,N_12586);
or U18405 (N_18405,N_11967,N_13282);
and U18406 (N_18406,N_14637,N_11197);
nor U18407 (N_18407,N_13389,N_12576);
nand U18408 (N_18408,N_14982,N_10946);
or U18409 (N_18409,N_13574,N_14133);
nor U18410 (N_18410,N_12752,N_12828);
xor U18411 (N_18411,N_12029,N_13298);
or U18412 (N_18412,N_14835,N_11072);
and U18413 (N_18413,N_10883,N_10691);
or U18414 (N_18414,N_13183,N_14832);
nor U18415 (N_18415,N_14685,N_14842);
nor U18416 (N_18416,N_12773,N_13226);
or U18417 (N_18417,N_12545,N_11294);
nand U18418 (N_18418,N_11732,N_11644);
xor U18419 (N_18419,N_14431,N_11275);
nor U18420 (N_18420,N_13630,N_12391);
xor U18421 (N_18421,N_14041,N_13232);
nand U18422 (N_18422,N_13564,N_12424);
nor U18423 (N_18423,N_14077,N_12699);
and U18424 (N_18424,N_12856,N_11841);
and U18425 (N_18425,N_13600,N_10886);
nand U18426 (N_18426,N_13635,N_11585);
nand U18427 (N_18427,N_10389,N_13466);
nor U18428 (N_18428,N_10381,N_10448);
and U18429 (N_18429,N_13684,N_10946);
nor U18430 (N_18430,N_10249,N_13364);
and U18431 (N_18431,N_12069,N_10845);
xor U18432 (N_18432,N_11256,N_14457);
nor U18433 (N_18433,N_10537,N_10187);
nor U18434 (N_18434,N_14161,N_14609);
and U18435 (N_18435,N_13293,N_12826);
nand U18436 (N_18436,N_12280,N_11931);
or U18437 (N_18437,N_12010,N_11380);
or U18438 (N_18438,N_11446,N_13318);
nand U18439 (N_18439,N_14423,N_13307);
nor U18440 (N_18440,N_10230,N_10572);
nand U18441 (N_18441,N_12069,N_10205);
and U18442 (N_18442,N_10099,N_12224);
or U18443 (N_18443,N_13469,N_14797);
or U18444 (N_18444,N_12757,N_13852);
or U18445 (N_18445,N_10854,N_10216);
and U18446 (N_18446,N_10248,N_13300);
and U18447 (N_18447,N_14969,N_11909);
xnor U18448 (N_18448,N_13518,N_13616);
nand U18449 (N_18449,N_13968,N_14774);
and U18450 (N_18450,N_12151,N_11034);
and U18451 (N_18451,N_10194,N_11388);
and U18452 (N_18452,N_10876,N_13081);
and U18453 (N_18453,N_13984,N_13563);
and U18454 (N_18454,N_13988,N_10734);
nand U18455 (N_18455,N_13074,N_11387);
nand U18456 (N_18456,N_11823,N_10752);
or U18457 (N_18457,N_12214,N_10098);
nor U18458 (N_18458,N_13453,N_11783);
nand U18459 (N_18459,N_12822,N_14434);
nor U18460 (N_18460,N_11283,N_12429);
and U18461 (N_18461,N_13566,N_14266);
xnor U18462 (N_18462,N_12289,N_10171);
nor U18463 (N_18463,N_14546,N_13477);
or U18464 (N_18464,N_14721,N_11448);
or U18465 (N_18465,N_14324,N_13111);
nor U18466 (N_18466,N_13912,N_13311);
and U18467 (N_18467,N_14725,N_14062);
and U18468 (N_18468,N_10871,N_10682);
or U18469 (N_18469,N_13671,N_12864);
nand U18470 (N_18470,N_13680,N_12625);
nand U18471 (N_18471,N_14743,N_13562);
nand U18472 (N_18472,N_12855,N_13001);
and U18473 (N_18473,N_14394,N_12711);
or U18474 (N_18474,N_14113,N_12645);
and U18475 (N_18475,N_10794,N_12335);
and U18476 (N_18476,N_13288,N_11037);
nor U18477 (N_18477,N_12317,N_11755);
and U18478 (N_18478,N_14359,N_14243);
or U18479 (N_18479,N_13967,N_11956);
and U18480 (N_18480,N_10254,N_11947);
nand U18481 (N_18481,N_13754,N_14534);
and U18482 (N_18482,N_11015,N_11518);
or U18483 (N_18483,N_11491,N_10261);
nand U18484 (N_18484,N_12226,N_13354);
nand U18485 (N_18485,N_10759,N_13440);
nor U18486 (N_18486,N_14894,N_12302);
and U18487 (N_18487,N_14741,N_11585);
or U18488 (N_18488,N_10815,N_13891);
or U18489 (N_18489,N_14117,N_14678);
and U18490 (N_18490,N_11164,N_13889);
or U18491 (N_18491,N_11382,N_11862);
xnor U18492 (N_18492,N_10518,N_14186);
or U18493 (N_18493,N_14982,N_13552);
nand U18494 (N_18494,N_13865,N_12882);
nand U18495 (N_18495,N_14055,N_11156);
and U18496 (N_18496,N_10986,N_11252);
xor U18497 (N_18497,N_14217,N_10133);
nor U18498 (N_18498,N_10048,N_14112);
xor U18499 (N_18499,N_14848,N_10407);
and U18500 (N_18500,N_10767,N_14509);
nand U18501 (N_18501,N_13512,N_10325);
nor U18502 (N_18502,N_12965,N_12453);
and U18503 (N_18503,N_13031,N_10536);
or U18504 (N_18504,N_11910,N_10556);
nor U18505 (N_18505,N_11235,N_12413);
nand U18506 (N_18506,N_10427,N_11950);
nand U18507 (N_18507,N_12222,N_11747);
or U18508 (N_18508,N_13591,N_12846);
and U18509 (N_18509,N_10913,N_11242);
or U18510 (N_18510,N_10668,N_11430);
nor U18511 (N_18511,N_13052,N_11688);
or U18512 (N_18512,N_14836,N_10611);
nor U18513 (N_18513,N_10348,N_11677);
and U18514 (N_18514,N_12293,N_14360);
or U18515 (N_18515,N_12641,N_10470);
and U18516 (N_18516,N_10283,N_10094);
nand U18517 (N_18517,N_12939,N_10554);
and U18518 (N_18518,N_12474,N_11144);
nor U18519 (N_18519,N_14849,N_12791);
nor U18520 (N_18520,N_13304,N_12080);
nand U18521 (N_18521,N_11166,N_13939);
xnor U18522 (N_18522,N_10895,N_11269);
nor U18523 (N_18523,N_13394,N_13009);
and U18524 (N_18524,N_10833,N_11701);
or U18525 (N_18525,N_14525,N_12477);
and U18526 (N_18526,N_11629,N_12894);
nand U18527 (N_18527,N_12913,N_13491);
or U18528 (N_18528,N_12431,N_14531);
or U18529 (N_18529,N_12446,N_12824);
and U18530 (N_18530,N_13531,N_11558);
or U18531 (N_18531,N_14465,N_12269);
or U18532 (N_18532,N_13192,N_13413);
and U18533 (N_18533,N_12850,N_12359);
nand U18534 (N_18534,N_12165,N_12560);
nand U18535 (N_18535,N_14934,N_13383);
or U18536 (N_18536,N_12976,N_13394);
or U18537 (N_18537,N_13044,N_11461);
nor U18538 (N_18538,N_12352,N_12340);
nand U18539 (N_18539,N_14756,N_10101);
or U18540 (N_18540,N_12465,N_14504);
or U18541 (N_18541,N_11755,N_11926);
nor U18542 (N_18542,N_10439,N_11344);
nand U18543 (N_18543,N_13944,N_10936);
or U18544 (N_18544,N_10909,N_13529);
nand U18545 (N_18545,N_12784,N_12760);
or U18546 (N_18546,N_10777,N_11204);
nor U18547 (N_18547,N_14813,N_10820);
or U18548 (N_18548,N_12882,N_13022);
nor U18549 (N_18549,N_11976,N_11692);
nor U18550 (N_18550,N_13931,N_12216);
and U18551 (N_18551,N_10298,N_10804);
nand U18552 (N_18552,N_13981,N_12300);
nand U18553 (N_18553,N_12500,N_10673);
nor U18554 (N_18554,N_10432,N_14489);
and U18555 (N_18555,N_12001,N_10272);
or U18556 (N_18556,N_10183,N_14178);
nand U18557 (N_18557,N_11338,N_12144);
or U18558 (N_18558,N_11339,N_11570);
nor U18559 (N_18559,N_10665,N_14348);
or U18560 (N_18560,N_12899,N_12071);
or U18561 (N_18561,N_12421,N_10647);
or U18562 (N_18562,N_10729,N_14851);
nand U18563 (N_18563,N_14560,N_10111);
nand U18564 (N_18564,N_13769,N_12295);
and U18565 (N_18565,N_11247,N_12140);
nor U18566 (N_18566,N_13230,N_10310);
or U18567 (N_18567,N_14196,N_12006);
nand U18568 (N_18568,N_12895,N_10040);
and U18569 (N_18569,N_13713,N_11063);
nor U18570 (N_18570,N_13618,N_10779);
nand U18571 (N_18571,N_11073,N_11596);
nor U18572 (N_18572,N_12520,N_14344);
nand U18573 (N_18573,N_11787,N_10014);
nand U18574 (N_18574,N_12904,N_12004);
xnor U18575 (N_18575,N_13716,N_14278);
nand U18576 (N_18576,N_10263,N_14371);
nor U18577 (N_18577,N_11984,N_10212);
xnor U18578 (N_18578,N_11224,N_14400);
and U18579 (N_18579,N_13647,N_11407);
or U18580 (N_18580,N_14994,N_10308);
nand U18581 (N_18581,N_13313,N_12228);
nand U18582 (N_18582,N_12552,N_10508);
xor U18583 (N_18583,N_12867,N_11884);
nand U18584 (N_18584,N_12303,N_12902);
and U18585 (N_18585,N_13716,N_11700);
and U18586 (N_18586,N_12906,N_12533);
and U18587 (N_18587,N_13291,N_11811);
or U18588 (N_18588,N_10655,N_13446);
or U18589 (N_18589,N_13464,N_10712);
nor U18590 (N_18590,N_13475,N_12766);
and U18591 (N_18591,N_12377,N_11854);
nand U18592 (N_18592,N_11390,N_12718);
nand U18593 (N_18593,N_12339,N_11766);
nor U18594 (N_18594,N_12343,N_14460);
nand U18595 (N_18595,N_10108,N_11406);
nand U18596 (N_18596,N_13026,N_14717);
nor U18597 (N_18597,N_14822,N_13083);
xnor U18598 (N_18598,N_11164,N_10794);
nand U18599 (N_18599,N_12963,N_14168);
nand U18600 (N_18600,N_11427,N_10497);
or U18601 (N_18601,N_12850,N_13371);
nor U18602 (N_18602,N_14905,N_10859);
and U18603 (N_18603,N_11923,N_12414);
xor U18604 (N_18604,N_12851,N_14878);
or U18605 (N_18605,N_10066,N_11778);
or U18606 (N_18606,N_11626,N_12631);
nand U18607 (N_18607,N_10433,N_12340);
and U18608 (N_18608,N_14811,N_14119);
nor U18609 (N_18609,N_11147,N_12329);
nand U18610 (N_18610,N_11951,N_10531);
and U18611 (N_18611,N_12138,N_13955);
xor U18612 (N_18612,N_14880,N_13289);
nor U18613 (N_18613,N_11266,N_14918);
nand U18614 (N_18614,N_14030,N_14390);
xnor U18615 (N_18615,N_14699,N_14275);
or U18616 (N_18616,N_11871,N_13965);
or U18617 (N_18617,N_12415,N_13543);
xnor U18618 (N_18618,N_12318,N_13654);
nand U18619 (N_18619,N_14554,N_13103);
nor U18620 (N_18620,N_11086,N_13005);
xor U18621 (N_18621,N_14460,N_14194);
nand U18622 (N_18622,N_11330,N_10493);
nor U18623 (N_18623,N_13766,N_10793);
and U18624 (N_18624,N_13497,N_13084);
nand U18625 (N_18625,N_14544,N_12698);
or U18626 (N_18626,N_14581,N_13194);
or U18627 (N_18627,N_12866,N_14685);
and U18628 (N_18628,N_10250,N_13092);
nand U18629 (N_18629,N_10433,N_10686);
or U18630 (N_18630,N_13266,N_14515);
or U18631 (N_18631,N_12636,N_12585);
nor U18632 (N_18632,N_12270,N_11378);
and U18633 (N_18633,N_12362,N_14991);
and U18634 (N_18634,N_12940,N_11664);
nor U18635 (N_18635,N_13347,N_14761);
nor U18636 (N_18636,N_12136,N_11907);
and U18637 (N_18637,N_12624,N_11829);
nand U18638 (N_18638,N_11451,N_13168);
xor U18639 (N_18639,N_14894,N_11273);
and U18640 (N_18640,N_10911,N_11416);
xor U18641 (N_18641,N_12271,N_11487);
nor U18642 (N_18642,N_13356,N_10202);
xnor U18643 (N_18643,N_12952,N_10890);
nor U18644 (N_18644,N_12703,N_10841);
nor U18645 (N_18645,N_11788,N_12368);
nand U18646 (N_18646,N_14500,N_10108);
nor U18647 (N_18647,N_12604,N_12727);
or U18648 (N_18648,N_10351,N_12282);
or U18649 (N_18649,N_13040,N_14670);
xnor U18650 (N_18650,N_10730,N_14241);
nand U18651 (N_18651,N_13271,N_10977);
and U18652 (N_18652,N_13638,N_12482);
nand U18653 (N_18653,N_14524,N_12341);
nand U18654 (N_18654,N_13160,N_14894);
and U18655 (N_18655,N_12948,N_11667);
or U18656 (N_18656,N_13802,N_10634);
or U18657 (N_18657,N_13102,N_14342);
and U18658 (N_18658,N_14845,N_13120);
nand U18659 (N_18659,N_10882,N_14358);
or U18660 (N_18660,N_14069,N_14454);
nand U18661 (N_18661,N_12362,N_10633);
and U18662 (N_18662,N_13004,N_11959);
or U18663 (N_18663,N_14399,N_13562);
or U18664 (N_18664,N_14547,N_14898);
xor U18665 (N_18665,N_13280,N_13331);
or U18666 (N_18666,N_14091,N_13209);
or U18667 (N_18667,N_14316,N_13308);
nor U18668 (N_18668,N_10184,N_13504);
and U18669 (N_18669,N_12187,N_12127);
and U18670 (N_18670,N_11852,N_12817);
nor U18671 (N_18671,N_13079,N_12912);
and U18672 (N_18672,N_12604,N_11700);
or U18673 (N_18673,N_14673,N_12187);
and U18674 (N_18674,N_10505,N_12615);
and U18675 (N_18675,N_11430,N_10130);
nor U18676 (N_18676,N_13651,N_12831);
or U18677 (N_18677,N_14157,N_13156);
nor U18678 (N_18678,N_13080,N_12520);
or U18679 (N_18679,N_13004,N_13210);
nand U18680 (N_18680,N_14033,N_11347);
nand U18681 (N_18681,N_11701,N_11346);
nor U18682 (N_18682,N_13020,N_11459);
or U18683 (N_18683,N_14456,N_14152);
and U18684 (N_18684,N_12641,N_14056);
and U18685 (N_18685,N_13212,N_12880);
nor U18686 (N_18686,N_11882,N_13083);
or U18687 (N_18687,N_14834,N_10437);
xnor U18688 (N_18688,N_12666,N_10903);
nor U18689 (N_18689,N_14574,N_10345);
nor U18690 (N_18690,N_14766,N_11839);
xnor U18691 (N_18691,N_10646,N_11916);
and U18692 (N_18692,N_11672,N_10144);
nor U18693 (N_18693,N_14174,N_12780);
nand U18694 (N_18694,N_11224,N_10577);
and U18695 (N_18695,N_14715,N_12530);
and U18696 (N_18696,N_11916,N_10460);
xor U18697 (N_18697,N_12698,N_13223);
and U18698 (N_18698,N_10270,N_13135);
nor U18699 (N_18699,N_13208,N_14650);
and U18700 (N_18700,N_10680,N_14230);
nor U18701 (N_18701,N_12146,N_10473);
or U18702 (N_18702,N_13315,N_11248);
and U18703 (N_18703,N_12466,N_10854);
nand U18704 (N_18704,N_11646,N_13377);
and U18705 (N_18705,N_12214,N_14178);
or U18706 (N_18706,N_14124,N_12093);
xor U18707 (N_18707,N_10236,N_10266);
nor U18708 (N_18708,N_12628,N_12708);
xnor U18709 (N_18709,N_13377,N_11926);
or U18710 (N_18710,N_13796,N_13740);
nand U18711 (N_18711,N_11174,N_12506);
xor U18712 (N_18712,N_10342,N_13719);
and U18713 (N_18713,N_12546,N_11434);
and U18714 (N_18714,N_10034,N_12183);
nor U18715 (N_18715,N_12424,N_14092);
and U18716 (N_18716,N_12972,N_12654);
xnor U18717 (N_18717,N_10447,N_14261);
xnor U18718 (N_18718,N_13825,N_14193);
and U18719 (N_18719,N_12252,N_14525);
nand U18720 (N_18720,N_11751,N_10709);
and U18721 (N_18721,N_13893,N_11727);
nor U18722 (N_18722,N_14406,N_14017);
and U18723 (N_18723,N_12048,N_14155);
or U18724 (N_18724,N_11005,N_14964);
and U18725 (N_18725,N_12145,N_12817);
or U18726 (N_18726,N_13564,N_14551);
xor U18727 (N_18727,N_10833,N_13643);
and U18728 (N_18728,N_12376,N_11649);
nor U18729 (N_18729,N_14948,N_11066);
and U18730 (N_18730,N_12284,N_10462);
nand U18731 (N_18731,N_13601,N_14186);
and U18732 (N_18732,N_14226,N_13695);
nand U18733 (N_18733,N_14514,N_10162);
nor U18734 (N_18734,N_10296,N_13596);
nor U18735 (N_18735,N_13930,N_13744);
or U18736 (N_18736,N_11115,N_14249);
nor U18737 (N_18737,N_10479,N_10931);
nor U18738 (N_18738,N_12682,N_14907);
nor U18739 (N_18739,N_10104,N_10385);
or U18740 (N_18740,N_10557,N_11510);
nor U18741 (N_18741,N_13676,N_14619);
nor U18742 (N_18742,N_10169,N_10009);
nand U18743 (N_18743,N_13800,N_10848);
nand U18744 (N_18744,N_13335,N_14101);
nor U18745 (N_18745,N_13520,N_12877);
and U18746 (N_18746,N_10135,N_12732);
or U18747 (N_18747,N_13497,N_11962);
or U18748 (N_18748,N_14081,N_11928);
nand U18749 (N_18749,N_14811,N_13623);
or U18750 (N_18750,N_13243,N_10636);
nor U18751 (N_18751,N_14267,N_12053);
nor U18752 (N_18752,N_14351,N_14304);
xor U18753 (N_18753,N_11016,N_14256);
nand U18754 (N_18754,N_10681,N_14665);
or U18755 (N_18755,N_12017,N_13638);
nor U18756 (N_18756,N_12339,N_11110);
nor U18757 (N_18757,N_14329,N_14510);
and U18758 (N_18758,N_11844,N_14073);
or U18759 (N_18759,N_13763,N_11115);
or U18760 (N_18760,N_10104,N_10334);
or U18761 (N_18761,N_12275,N_13170);
and U18762 (N_18762,N_14698,N_11369);
xnor U18763 (N_18763,N_10682,N_13501);
or U18764 (N_18764,N_12027,N_13600);
nand U18765 (N_18765,N_12245,N_12262);
and U18766 (N_18766,N_11986,N_14574);
or U18767 (N_18767,N_10034,N_10582);
or U18768 (N_18768,N_11253,N_13727);
nor U18769 (N_18769,N_13485,N_11416);
or U18770 (N_18770,N_14485,N_12123);
or U18771 (N_18771,N_13527,N_13330);
or U18772 (N_18772,N_13916,N_14833);
nand U18773 (N_18773,N_12562,N_14034);
and U18774 (N_18774,N_13655,N_11797);
and U18775 (N_18775,N_14658,N_11138);
or U18776 (N_18776,N_14425,N_11021);
nand U18777 (N_18777,N_12005,N_13670);
nor U18778 (N_18778,N_13224,N_11900);
or U18779 (N_18779,N_10779,N_13155);
and U18780 (N_18780,N_11417,N_13694);
nand U18781 (N_18781,N_14273,N_13439);
and U18782 (N_18782,N_10206,N_10691);
and U18783 (N_18783,N_13919,N_14775);
xnor U18784 (N_18784,N_11495,N_13006);
or U18785 (N_18785,N_14429,N_10192);
nand U18786 (N_18786,N_11806,N_12689);
and U18787 (N_18787,N_13953,N_13613);
nand U18788 (N_18788,N_14483,N_10518);
xor U18789 (N_18789,N_10149,N_11171);
xor U18790 (N_18790,N_14497,N_11703);
nor U18791 (N_18791,N_14535,N_11059);
xor U18792 (N_18792,N_11443,N_14566);
nor U18793 (N_18793,N_12817,N_10385);
nand U18794 (N_18794,N_14695,N_14143);
and U18795 (N_18795,N_13831,N_13850);
or U18796 (N_18796,N_10486,N_12191);
or U18797 (N_18797,N_14597,N_12255);
nand U18798 (N_18798,N_13217,N_11970);
nand U18799 (N_18799,N_12507,N_10014);
or U18800 (N_18800,N_11018,N_11762);
nand U18801 (N_18801,N_14732,N_13202);
nand U18802 (N_18802,N_14318,N_14897);
nor U18803 (N_18803,N_10953,N_13921);
nor U18804 (N_18804,N_13514,N_10811);
or U18805 (N_18805,N_11928,N_10681);
and U18806 (N_18806,N_13426,N_14473);
and U18807 (N_18807,N_12865,N_14223);
or U18808 (N_18808,N_12442,N_14731);
or U18809 (N_18809,N_11678,N_11367);
nor U18810 (N_18810,N_14266,N_14567);
and U18811 (N_18811,N_13583,N_11912);
or U18812 (N_18812,N_10981,N_12064);
or U18813 (N_18813,N_10185,N_11998);
and U18814 (N_18814,N_11954,N_14056);
nand U18815 (N_18815,N_12167,N_13273);
or U18816 (N_18816,N_12544,N_13136);
and U18817 (N_18817,N_12563,N_11537);
or U18818 (N_18818,N_11861,N_12237);
or U18819 (N_18819,N_13783,N_13585);
nor U18820 (N_18820,N_10972,N_14531);
and U18821 (N_18821,N_10159,N_13763);
nand U18822 (N_18822,N_14764,N_11142);
and U18823 (N_18823,N_14297,N_11675);
nand U18824 (N_18824,N_12240,N_12010);
and U18825 (N_18825,N_10085,N_14414);
or U18826 (N_18826,N_12782,N_12164);
nand U18827 (N_18827,N_10257,N_12512);
nand U18828 (N_18828,N_11771,N_10899);
and U18829 (N_18829,N_11619,N_12538);
nand U18830 (N_18830,N_10601,N_12836);
nor U18831 (N_18831,N_10164,N_11176);
and U18832 (N_18832,N_14532,N_11391);
or U18833 (N_18833,N_13726,N_10531);
xnor U18834 (N_18834,N_14195,N_14669);
nor U18835 (N_18835,N_13630,N_11852);
or U18836 (N_18836,N_13733,N_12069);
nand U18837 (N_18837,N_10462,N_11109);
nor U18838 (N_18838,N_10456,N_12094);
and U18839 (N_18839,N_12228,N_12173);
xor U18840 (N_18840,N_13848,N_14564);
nor U18841 (N_18841,N_10180,N_14024);
or U18842 (N_18842,N_14336,N_11648);
or U18843 (N_18843,N_13978,N_10142);
and U18844 (N_18844,N_13708,N_13357);
nor U18845 (N_18845,N_10356,N_13437);
nor U18846 (N_18846,N_13658,N_13198);
nor U18847 (N_18847,N_12515,N_13197);
nand U18848 (N_18848,N_13929,N_10642);
nand U18849 (N_18849,N_14034,N_10599);
nand U18850 (N_18850,N_13449,N_14762);
nor U18851 (N_18851,N_11189,N_11071);
nor U18852 (N_18852,N_10765,N_14159);
or U18853 (N_18853,N_14525,N_12788);
xor U18854 (N_18854,N_10607,N_13692);
or U18855 (N_18855,N_14613,N_13506);
or U18856 (N_18856,N_13004,N_14240);
nand U18857 (N_18857,N_13285,N_14481);
or U18858 (N_18858,N_14550,N_12211);
nor U18859 (N_18859,N_10548,N_13951);
or U18860 (N_18860,N_13805,N_10376);
nor U18861 (N_18861,N_11247,N_10179);
or U18862 (N_18862,N_11932,N_10057);
or U18863 (N_18863,N_10855,N_11752);
nand U18864 (N_18864,N_13233,N_11086);
nor U18865 (N_18865,N_12719,N_10583);
nor U18866 (N_18866,N_11750,N_13123);
or U18867 (N_18867,N_12703,N_10282);
nand U18868 (N_18868,N_12480,N_14941);
nor U18869 (N_18869,N_10609,N_14654);
and U18870 (N_18870,N_12241,N_10533);
nor U18871 (N_18871,N_12436,N_10986);
or U18872 (N_18872,N_10563,N_13500);
nand U18873 (N_18873,N_11686,N_13058);
nor U18874 (N_18874,N_12529,N_11428);
nand U18875 (N_18875,N_12720,N_13726);
nand U18876 (N_18876,N_14180,N_10196);
and U18877 (N_18877,N_14710,N_12395);
nand U18878 (N_18878,N_14616,N_10685);
nand U18879 (N_18879,N_11912,N_13417);
and U18880 (N_18880,N_12367,N_14733);
nor U18881 (N_18881,N_11350,N_14759);
nand U18882 (N_18882,N_14057,N_14826);
or U18883 (N_18883,N_12034,N_10214);
nand U18884 (N_18884,N_11629,N_11576);
or U18885 (N_18885,N_11615,N_13435);
nor U18886 (N_18886,N_10192,N_13021);
nor U18887 (N_18887,N_13963,N_13950);
nor U18888 (N_18888,N_12373,N_10541);
nor U18889 (N_18889,N_14623,N_12088);
nand U18890 (N_18890,N_12390,N_10890);
xor U18891 (N_18891,N_12166,N_11750);
nand U18892 (N_18892,N_14877,N_10288);
nand U18893 (N_18893,N_12314,N_10901);
and U18894 (N_18894,N_11063,N_13057);
xnor U18895 (N_18895,N_10149,N_13647);
and U18896 (N_18896,N_14264,N_12328);
or U18897 (N_18897,N_10399,N_13058);
xor U18898 (N_18898,N_13965,N_10018);
nor U18899 (N_18899,N_12871,N_10095);
nand U18900 (N_18900,N_12757,N_11367);
and U18901 (N_18901,N_11698,N_11000);
nand U18902 (N_18902,N_14177,N_12245);
and U18903 (N_18903,N_11611,N_11501);
nor U18904 (N_18904,N_11839,N_13902);
or U18905 (N_18905,N_11963,N_11618);
nor U18906 (N_18906,N_11616,N_12544);
nand U18907 (N_18907,N_12008,N_13567);
or U18908 (N_18908,N_13426,N_12293);
nand U18909 (N_18909,N_14419,N_12982);
nand U18910 (N_18910,N_11062,N_12967);
xnor U18911 (N_18911,N_11029,N_13000);
and U18912 (N_18912,N_11685,N_10234);
nand U18913 (N_18913,N_12724,N_14423);
or U18914 (N_18914,N_12707,N_13477);
or U18915 (N_18915,N_10014,N_11966);
nand U18916 (N_18916,N_12369,N_12950);
nor U18917 (N_18917,N_12316,N_10380);
or U18918 (N_18918,N_10048,N_11585);
or U18919 (N_18919,N_14969,N_12542);
xnor U18920 (N_18920,N_14072,N_11769);
nand U18921 (N_18921,N_13931,N_14571);
and U18922 (N_18922,N_13850,N_10103);
and U18923 (N_18923,N_14707,N_13015);
and U18924 (N_18924,N_14776,N_11721);
nor U18925 (N_18925,N_13259,N_11992);
and U18926 (N_18926,N_13113,N_10747);
nor U18927 (N_18927,N_13315,N_13991);
nor U18928 (N_18928,N_13841,N_13251);
and U18929 (N_18929,N_13841,N_11898);
nand U18930 (N_18930,N_12782,N_12414);
nand U18931 (N_18931,N_11965,N_14138);
or U18932 (N_18932,N_14240,N_14529);
nor U18933 (N_18933,N_11666,N_10885);
or U18934 (N_18934,N_14202,N_11934);
and U18935 (N_18935,N_14182,N_14884);
and U18936 (N_18936,N_12736,N_11720);
nand U18937 (N_18937,N_11397,N_14564);
or U18938 (N_18938,N_11788,N_12395);
nor U18939 (N_18939,N_14120,N_13455);
nor U18940 (N_18940,N_10248,N_14770);
nand U18941 (N_18941,N_14282,N_12509);
or U18942 (N_18942,N_11948,N_14069);
and U18943 (N_18943,N_12420,N_14177);
nor U18944 (N_18944,N_11268,N_13718);
or U18945 (N_18945,N_11774,N_14727);
and U18946 (N_18946,N_12290,N_11262);
nand U18947 (N_18947,N_13403,N_10332);
xnor U18948 (N_18948,N_14295,N_12746);
nor U18949 (N_18949,N_14104,N_14848);
or U18950 (N_18950,N_10993,N_11598);
or U18951 (N_18951,N_14343,N_11751);
and U18952 (N_18952,N_10046,N_14156);
nand U18953 (N_18953,N_10542,N_13570);
and U18954 (N_18954,N_10318,N_12013);
or U18955 (N_18955,N_11263,N_12523);
xor U18956 (N_18956,N_13593,N_11798);
and U18957 (N_18957,N_11059,N_10757);
nor U18958 (N_18958,N_10547,N_13600);
or U18959 (N_18959,N_11953,N_13867);
or U18960 (N_18960,N_11387,N_11415);
and U18961 (N_18961,N_14028,N_10775);
or U18962 (N_18962,N_12610,N_14539);
and U18963 (N_18963,N_10883,N_12021);
and U18964 (N_18964,N_14734,N_10915);
nor U18965 (N_18965,N_10418,N_13153);
or U18966 (N_18966,N_11021,N_12499);
nand U18967 (N_18967,N_12399,N_12330);
nand U18968 (N_18968,N_11833,N_14495);
nand U18969 (N_18969,N_14574,N_12948);
and U18970 (N_18970,N_14830,N_11081);
or U18971 (N_18971,N_14003,N_13629);
nand U18972 (N_18972,N_14679,N_10484);
or U18973 (N_18973,N_10558,N_10097);
or U18974 (N_18974,N_12891,N_14168);
nand U18975 (N_18975,N_14807,N_14691);
xor U18976 (N_18976,N_12675,N_11379);
xor U18977 (N_18977,N_14468,N_11389);
nor U18978 (N_18978,N_14023,N_10950);
xnor U18979 (N_18979,N_10294,N_14268);
nor U18980 (N_18980,N_10529,N_11264);
and U18981 (N_18981,N_12104,N_11784);
or U18982 (N_18982,N_11043,N_10214);
nand U18983 (N_18983,N_11461,N_13135);
and U18984 (N_18984,N_10135,N_10756);
nor U18985 (N_18985,N_10207,N_14565);
nor U18986 (N_18986,N_13973,N_12405);
nand U18987 (N_18987,N_10502,N_12401);
nand U18988 (N_18988,N_10961,N_13570);
and U18989 (N_18989,N_14251,N_12248);
nand U18990 (N_18990,N_11846,N_10054);
xor U18991 (N_18991,N_12241,N_14562);
nor U18992 (N_18992,N_10317,N_10865);
or U18993 (N_18993,N_11217,N_10743);
and U18994 (N_18994,N_10112,N_14198);
nor U18995 (N_18995,N_11414,N_10835);
nor U18996 (N_18996,N_11914,N_12431);
nand U18997 (N_18997,N_10635,N_11094);
nor U18998 (N_18998,N_12506,N_14085);
and U18999 (N_18999,N_10286,N_11501);
nand U19000 (N_19000,N_14772,N_11363);
xnor U19001 (N_19001,N_14520,N_13257);
nand U19002 (N_19002,N_12286,N_13699);
or U19003 (N_19003,N_12858,N_12148);
nand U19004 (N_19004,N_10395,N_13330);
or U19005 (N_19005,N_10139,N_11353);
and U19006 (N_19006,N_10771,N_10904);
nor U19007 (N_19007,N_10629,N_12244);
or U19008 (N_19008,N_14907,N_10174);
or U19009 (N_19009,N_13097,N_11934);
or U19010 (N_19010,N_12296,N_11684);
or U19011 (N_19011,N_11834,N_12709);
nor U19012 (N_19012,N_10842,N_13756);
and U19013 (N_19013,N_14645,N_12484);
nor U19014 (N_19014,N_12081,N_13947);
nand U19015 (N_19015,N_13802,N_12498);
nor U19016 (N_19016,N_10836,N_11835);
nor U19017 (N_19017,N_13922,N_12582);
or U19018 (N_19018,N_14083,N_11394);
or U19019 (N_19019,N_14858,N_14674);
nand U19020 (N_19020,N_14372,N_14211);
nor U19021 (N_19021,N_13377,N_11940);
and U19022 (N_19022,N_11472,N_14639);
nor U19023 (N_19023,N_11173,N_14077);
or U19024 (N_19024,N_13580,N_12618);
and U19025 (N_19025,N_11817,N_14062);
and U19026 (N_19026,N_11771,N_12283);
and U19027 (N_19027,N_14971,N_11169);
and U19028 (N_19028,N_14720,N_13509);
or U19029 (N_19029,N_14696,N_13583);
or U19030 (N_19030,N_12204,N_13363);
or U19031 (N_19031,N_13966,N_10322);
or U19032 (N_19032,N_14281,N_14291);
nand U19033 (N_19033,N_14070,N_10933);
nor U19034 (N_19034,N_11561,N_13967);
nand U19035 (N_19035,N_10608,N_14203);
and U19036 (N_19036,N_14651,N_11066);
or U19037 (N_19037,N_10835,N_10924);
xor U19038 (N_19038,N_12385,N_11998);
xnor U19039 (N_19039,N_13888,N_13051);
and U19040 (N_19040,N_13277,N_11382);
or U19041 (N_19041,N_14771,N_12373);
or U19042 (N_19042,N_14479,N_14652);
and U19043 (N_19043,N_12088,N_12813);
xnor U19044 (N_19044,N_10574,N_13420);
xor U19045 (N_19045,N_13043,N_14364);
nand U19046 (N_19046,N_13766,N_14358);
nor U19047 (N_19047,N_13534,N_13552);
and U19048 (N_19048,N_14653,N_12994);
nor U19049 (N_19049,N_14599,N_12661);
xor U19050 (N_19050,N_12233,N_14707);
nor U19051 (N_19051,N_12049,N_12716);
and U19052 (N_19052,N_14386,N_11143);
and U19053 (N_19053,N_10791,N_10824);
and U19054 (N_19054,N_10425,N_10559);
nand U19055 (N_19055,N_11564,N_13863);
nand U19056 (N_19056,N_11804,N_13657);
and U19057 (N_19057,N_13419,N_12129);
or U19058 (N_19058,N_11730,N_11338);
nand U19059 (N_19059,N_14004,N_14322);
and U19060 (N_19060,N_14128,N_11146);
nor U19061 (N_19061,N_12236,N_12138);
xor U19062 (N_19062,N_12124,N_10752);
or U19063 (N_19063,N_10905,N_13522);
or U19064 (N_19064,N_11969,N_14039);
or U19065 (N_19065,N_12195,N_10293);
xor U19066 (N_19066,N_13891,N_11900);
and U19067 (N_19067,N_14751,N_13733);
nor U19068 (N_19068,N_13794,N_10609);
or U19069 (N_19069,N_12442,N_10709);
or U19070 (N_19070,N_10338,N_14127);
and U19071 (N_19071,N_12717,N_14420);
nand U19072 (N_19072,N_11379,N_14828);
or U19073 (N_19073,N_10528,N_12240);
nor U19074 (N_19074,N_13671,N_10249);
or U19075 (N_19075,N_10822,N_11259);
nor U19076 (N_19076,N_13602,N_10058);
nor U19077 (N_19077,N_14737,N_13762);
and U19078 (N_19078,N_10544,N_14264);
xnor U19079 (N_19079,N_12751,N_13734);
xnor U19080 (N_19080,N_11954,N_10841);
xor U19081 (N_19081,N_13907,N_12983);
or U19082 (N_19082,N_11245,N_12097);
nor U19083 (N_19083,N_13897,N_10542);
or U19084 (N_19084,N_11318,N_11532);
and U19085 (N_19085,N_11004,N_11821);
or U19086 (N_19086,N_10264,N_11679);
or U19087 (N_19087,N_14773,N_10595);
and U19088 (N_19088,N_11408,N_10928);
or U19089 (N_19089,N_11975,N_10466);
xnor U19090 (N_19090,N_11364,N_10935);
xnor U19091 (N_19091,N_14769,N_14950);
and U19092 (N_19092,N_12715,N_13582);
nand U19093 (N_19093,N_13447,N_13942);
and U19094 (N_19094,N_13833,N_10198);
nand U19095 (N_19095,N_14222,N_11093);
and U19096 (N_19096,N_10459,N_10355);
or U19097 (N_19097,N_10700,N_11065);
nand U19098 (N_19098,N_14134,N_10658);
nor U19099 (N_19099,N_10385,N_10769);
nand U19100 (N_19100,N_11199,N_11113);
or U19101 (N_19101,N_10593,N_12524);
nand U19102 (N_19102,N_14337,N_11991);
nor U19103 (N_19103,N_12420,N_14544);
nand U19104 (N_19104,N_13654,N_11231);
and U19105 (N_19105,N_11861,N_12288);
and U19106 (N_19106,N_10933,N_13634);
and U19107 (N_19107,N_12116,N_14685);
or U19108 (N_19108,N_12967,N_11887);
nor U19109 (N_19109,N_11180,N_14411);
and U19110 (N_19110,N_11683,N_11292);
and U19111 (N_19111,N_14981,N_14398);
nor U19112 (N_19112,N_14269,N_14002);
or U19113 (N_19113,N_13011,N_13900);
nor U19114 (N_19114,N_12225,N_13196);
nand U19115 (N_19115,N_11624,N_10557);
nor U19116 (N_19116,N_12997,N_14291);
nand U19117 (N_19117,N_13917,N_14708);
or U19118 (N_19118,N_13400,N_10882);
nor U19119 (N_19119,N_14510,N_12430);
nor U19120 (N_19120,N_11002,N_14064);
nand U19121 (N_19121,N_11812,N_12994);
and U19122 (N_19122,N_13963,N_14883);
nand U19123 (N_19123,N_12850,N_13052);
nor U19124 (N_19124,N_13568,N_12405);
xor U19125 (N_19125,N_10745,N_14765);
or U19126 (N_19126,N_14868,N_13215);
nand U19127 (N_19127,N_12296,N_11351);
and U19128 (N_19128,N_11016,N_11943);
nand U19129 (N_19129,N_14661,N_14223);
or U19130 (N_19130,N_11808,N_10112);
nor U19131 (N_19131,N_14945,N_11220);
nor U19132 (N_19132,N_11393,N_10103);
and U19133 (N_19133,N_12022,N_10138);
nand U19134 (N_19134,N_11677,N_11688);
or U19135 (N_19135,N_13423,N_11028);
nor U19136 (N_19136,N_12682,N_11735);
nand U19137 (N_19137,N_14520,N_10172);
and U19138 (N_19138,N_10927,N_13093);
nand U19139 (N_19139,N_13577,N_10273);
xnor U19140 (N_19140,N_14071,N_12020);
nor U19141 (N_19141,N_10034,N_12863);
nor U19142 (N_19142,N_11367,N_13530);
or U19143 (N_19143,N_11183,N_11445);
or U19144 (N_19144,N_12384,N_12383);
or U19145 (N_19145,N_12831,N_14062);
nand U19146 (N_19146,N_13866,N_13333);
xnor U19147 (N_19147,N_14302,N_12271);
and U19148 (N_19148,N_13126,N_13183);
and U19149 (N_19149,N_10044,N_10663);
nand U19150 (N_19150,N_12459,N_10482);
nor U19151 (N_19151,N_10714,N_10863);
nor U19152 (N_19152,N_14982,N_14388);
and U19153 (N_19153,N_14485,N_10955);
or U19154 (N_19154,N_12536,N_13277);
nor U19155 (N_19155,N_11150,N_12871);
and U19156 (N_19156,N_12282,N_12651);
nand U19157 (N_19157,N_10933,N_14352);
nor U19158 (N_19158,N_13024,N_12513);
nor U19159 (N_19159,N_14856,N_14927);
or U19160 (N_19160,N_11739,N_12747);
nand U19161 (N_19161,N_10124,N_12406);
nand U19162 (N_19162,N_13587,N_10810);
and U19163 (N_19163,N_10594,N_10206);
or U19164 (N_19164,N_12164,N_12134);
nand U19165 (N_19165,N_10759,N_12639);
and U19166 (N_19166,N_13234,N_12838);
xnor U19167 (N_19167,N_13447,N_13365);
nor U19168 (N_19168,N_13628,N_12990);
nor U19169 (N_19169,N_10866,N_10735);
nand U19170 (N_19170,N_13648,N_11187);
nor U19171 (N_19171,N_13095,N_13115);
and U19172 (N_19172,N_13276,N_11478);
and U19173 (N_19173,N_13837,N_12819);
and U19174 (N_19174,N_11258,N_11585);
or U19175 (N_19175,N_11346,N_14576);
nor U19176 (N_19176,N_14275,N_11169);
and U19177 (N_19177,N_13810,N_13180);
nor U19178 (N_19178,N_13558,N_14692);
nand U19179 (N_19179,N_11789,N_11009);
or U19180 (N_19180,N_12054,N_10590);
xnor U19181 (N_19181,N_12738,N_13982);
nor U19182 (N_19182,N_11849,N_11256);
nand U19183 (N_19183,N_13867,N_14721);
nand U19184 (N_19184,N_14741,N_12011);
and U19185 (N_19185,N_13791,N_10415);
nand U19186 (N_19186,N_13074,N_14808);
nand U19187 (N_19187,N_10160,N_11972);
nor U19188 (N_19188,N_10343,N_13016);
or U19189 (N_19189,N_10267,N_10840);
nand U19190 (N_19190,N_14137,N_12406);
and U19191 (N_19191,N_13891,N_14993);
and U19192 (N_19192,N_11514,N_14360);
or U19193 (N_19193,N_12984,N_10714);
or U19194 (N_19194,N_14312,N_10601);
or U19195 (N_19195,N_14541,N_11965);
and U19196 (N_19196,N_12269,N_12980);
nand U19197 (N_19197,N_14409,N_12133);
xnor U19198 (N_19198,N_10071,N_13434);
nand U19199 (N_19199,N_14176,N_14942);
and U19200 (N_19200,N_10338,N_14318);
and U19201 (N_19201,N_13458,N_13287);
or U19202 (N_19202,N_14620,N_12349);
nand U19203 (N_19203,N_10029,N_12416);
nor U19204 (N_19204,N_11625,N_11904);
nand U19205 (N_19205,N_13893,N_12184);
or U19206 (N_19206,N_10130,N_12822);
or U19207 (N_19207,N_11465,N_14039);
nor U19208 (N_19208,N_10010,N_13514);
nor U19209 (N_19209,N_14207,N_14763);
nor U19210 (N_19210,N_12899,N_13122);
and U19211 (N_19211,N_12871,N_11351);
nand U19212 (N_19212,N_11211,N_14802);
xor U19213 (N_19213,N_11539,N_11556);
or U19214 (N_19214,N_13921,N_13551);
or U19215 (N_19215,N_10880,N_11947);
nor U19216 (N_19216,N_10906,N_11360);
xor U19217 (N_19217,N_14890,N_13688);
or U19218 (N_19218,N_10787,N_12666);
and U19219 (N_19219,N_12471,N_13805);
or U19220 (N_19220,N_10188,N_12420);
xnor U19221 (N_19221,N_14599,N_12810);
and U19222 (N_19222,N_14327,N_13050);
and U19223 (N_19223,N_12325,N_10688);
and U19224 (N_19224,N_14281,N_11381);
or U19225 (N_19225,N_11441,N_14645);
or U19226 (N_19226,N_12134,N_14440);
nand U19227 (N_19227,N_10289,N_14543);
or U19228 (N_19228,N_10558,N_13663);
nor U19229 (N_19229,N_12901,N_10541);
nand U19230 (N_19230,N_11178,N_13190);
xor U19231 (N_19231,N_10133,N_14175);
nor U19232 (N_19232,N_10664,N_13340);
or U19233 (N_19233,N_12244,N_14307);
xor U19234 (N_19234,N_10850,N_11172);
or U19235 (N_19235,N_14844,N_10572);
or U19236 (N_19236,N_10215,N_12200);
or U19237 (N_19237,N_11752,N_14969);
xnor U19238 (N_19238,N_13279,N_10270);
nor U19239 (N_19239,N_11781,N_14407);
xnor U19240 (N_19240,N_14982,N_13187);
and U19241 (N_19241,N_13877,N_13955);
or U19242 (N_19242,N_13069,N_11912);
or U19243 (N_19243,N_11215,N_12229);
or U19244 (N_19244,N_13163,N_12376);
and U19245 (N_19245,N_14545,N_12204);
nand U19246 (N_19246,N_10488,N_11432);
or U19247 (N_19247,N_11267,N_10808);
nand U19248 (N_19248,N_10508,N_13155);
nand U19249 (N_19249,N_11458,N_11109);
or U19250 (N_19250,N_11453,N_11743);
xnor U19251 (N_19251,N_11087,N_10940);
and U19252 (N_19252,N_10165,N_11282);
nand U19253 (N_19253,N_12679,N_11260);
or U19254 (N_19254,N_10178,N_10090);
nor U19255 (N_19255,N_13557,N_13164);
nand U19256 (N_19256,N_14837,N_10464);
or U19257 (N_19257,N_12816,N_11952);
and U19258 (N_19258,N_12196,N_11844);
xnor U19259 (N_19259,N_10309,N_12309);
or U19260 (N_19260,N_11763,N_11092);
nor U19261 (N_19261,N_10544,N_12919);
xnor U19262 (N_19262,N_12371,N_14963);
nand U19263 (N_19263,N_13694,N_10596);
and U19264 (N_19264,N_11319,N_13736);
or U19265 (N_19265,N_12208,N_11463);
nor U19266 (N_19266,N_10830,N_14648);
or U19267 (N_19267,N_11363,N_13576);
or U19268 (N_19268,N_13108,N_12469);
nor U19269 (N_19269,N_10316,N_10542);
nor U19270 (N_19270,N_14268,N_12251);
and U19271 (N_19271,N_11837,N_11625);
and U19272 (N_19272,N_13191,N_10983);
nor U19273 (N_19273,N_13516,N_13915);
or U19274 (N_19274,N_10817,N_13012);
and U19275 (N_19275,N_14981,N_12499);
xor U19276 (N_19276,N_11002,N_14965);
nor U19277 (N_19277,N_13049,N_10857);
or U19278 (N_19278,N_10069,N_12020);
and U19279 (N_19279,N_13038,N_13552);
or U19280 (N_19280,N_10941,N_11493);
and U19281 (N_19281,N_10737,N_11927);
xnor U19282 (N_19282,N_10595,N_13227);
nor U19283 (N_19283,N_10622,N_12650);
nor U19284 (N_19284,N_13474,N_12178);
nand U19285 (N_19285,N_10657,N_11940);
or U19286 (N_19286,N_13410,N_12192);
and U19287 (N_19287,N_12613,N_14133);
nor U19288 (N_19288,N_11195,N_14386);
nor U19289 (N_19289,N_10440,N_14391);
nand U19290 (N_19290,N_14216,N_10923);
nand U19291 (N_19291,N_11539,N_12690);
xor U19292 (N_19292,N_13553,N_12123);
nor U19293 (N_19293,N_11250,N_11963);
nand U19294 (N_19294,N_13809,N_14163);
and U19295 (N_19295,N_14122,N_13684);
xor U19296 (N_19296,N_12663,N_12307);
nor U19297 (N_19297,N_13926,N_12558);
or U19298 (N_19298,N_10393,N_10702);
nand U19299 (N_19299,N_11034,N_13954);
nor U19300 (N_19300,N_10170,N_10885);
and U19301 (N_19301,N_14280,N_13951);
nor U19302 (N_19302,N_11406,N_12661);
xor U19303 (N_19303,N_12765,N_13284);
xor U19304 (N_19304,N_14561,N_11814);
nand U19305 (N_19305,N_11184,N_12909);
or U19306 (N_19306,N_10324,N_10520);
nand U19307 (N_19307,N_12295,N_11999);
and U19308 (N_19308,N_14109,N_10278);
xnor U19309 (N_19309,N_13105,N_11719);
nor U19310 (N_19310,N_12064,N_14337);
nor U19311 (N_19311,N_14616,N_10687);
or U19312 (N_19312,N_10766,N_13474);
nand U19313 (N_19313,N_12816,N_14468);
nand U19314 (N_19314,N_11024,N_12109);
and U19315 (N_19315,N_14300,N_12463);
nor U19316 (N_19316,N_10785,N_10174);
and U19317 (N_19317,N_14827,N_12268);
and U19318 (N_19318,N_10683,N_12179);
nor U19319 (N_19319,N_14408,N_10262);
xor U19320 (N_19320,N_14787,N_10719);
nand U19321 (N_19321,N_10852,N_14718);
nor U19322 (N_19322,N_14098,N_12482);
nand U19323 (N_19323,N_13860,N_11898);
nand U19324 (N_19324,N_13949,N_14365);
nor U19325 (N_19325,N_13476,N_12165);
nand U19326 (N_19326,N_13362,N_10798);
nand U19327 (N_19327,N_14092,N_11159);
nor U19328 (N_19328,N_12488,N_11420);
or U19329 (N_19329,N_12020,N_13237);
nor U19330 (N_19330,N_11462,N_12947);
and U19331 (N_19331,N_14459,N_11075);
and U19332 (N_19332,N_12685,N_14705);
xor U19333 (N_19333,N_13555,N_14437);
or U19334 (N_19334,N_10566,N_11675);
nand U19335 (N_19335,N_11741,N_14749);
nor U19336 (N_19336,N_13775,N_13810);
nor U19337 (N_19337,N_10290,N_14461);
or U19338 (N_19338,N_10981,N_12709);
nand U19339 (N_19339,N_13522,N_14261);
nor U19340 (N_19340,N_12426,N_11218);
and U19341 (N_19341,N_13818,N_12252);
xnor U19342 (N_19342,N_10061,N_10273);
nor U19343 (N_19343,N_11355,N_10007);
or U19344 (N_19344,N_12376,N_10064);
nor U19345 (N_19345,N_13663,N_11446);
or U19346 (N_19346,N_14231,N_11092);
nor U19347 (N_19347,N_12679,N_11728);
nand U19348 (N_19348,N_14155,N_13642);
nand U19349 (N_19349,N_10566,N_12226);
and U19350 (N_19350,N_13326,N_12933);
nor U19351 (N_19351,N_11295,N_12597);
or U19352 (N_19352,N_14864,N_12621);
or U19353 (N_19353,N_11527,N_10058);
xor U19354 (N_19354,N_11456,N_12126);
nor U19355 (N_19355,N_10450,N_10651);
nor U19356 (N_19356,N_13270,N_12174);
nor U19357 (N_19357,N_14722,N_11203);
nor U19358 (N_19358,N_11262,N_12784);
nand U19359 (N_19359,N_13496,N_12891);
nor U19360 (N_19360,N_13669,N_12730);
xnor U19361 (N_19361,N_11719,N_10904);
and U19362 (N_19362,N_13669,N_13543);
and U19363 (N_19363,N_13073,N_13034);
nor U19364 (N_19364,N_12517,N_14945);
or U19365 (N_19365,N_14395,N_13639);
and U19366 (N_19366,N_10109,N_11122);
xnor U19367 (N_19367,N_12062,N_10457);
xnor U19368 (N_19368,N_12920,N_12812);
or U19369 (N_19369,N_14821,N_12076);
and U19370 (N_19370,N_12106,N_12010);
nand U19371 (N_19371,N_12563,N_10515);
and U19372 (N_19372,N_10363,N_13650);
and U19373 (N_19373,N_12142,N_13609);
nor U19374 (N_19374,N_12459,N_13793);
and U19375 (N_19375,N_10314,N_10362);
and U19376 (N_19376,N_10494,N_12370);
nor U19377 (N_19377,N_14557,N_12280);
xor U19378 (N_19378,N_11641,N_11246);
and U19379 (N_19379,N_10389,N_10117);
or U19380 (N_19380,N_14160,N_11624);
and U19381 (N_19381,N_12687,N_11633);
xnor U19382 (N_19382,N_12827,N_12232);
nand U19383 (N_19383,N_11301,N_11549);
or U19384 (N_19384,N_14445,N_10590);
or U19385 (N_19385,N_12466,N_12523);
or U19386 (N_19386,N_14031,N_11273);
or U19387 (N_19387,N_10893,N_14039);
xnor U19388 (N_19388,N_14452,N_13029);
nor U19389 (N_19389,N_10942,N_11130);
or U19390 (N_19390,N_13540,N_12700);
nand U19391 (N_19391,N_13823,N_14169);
nand U19392 (N_19392,N_13417,N_12949);
xor U19393 (N_19393,N_13507,N_10191);
and U19394 (N_19394,N_10704,N_11382);
and U19395 (N_19395,N_11704,N_10532);
or U19396 (N_19396,N_10548,N_13558);
xor U19397 (N_19397,N_14085,N_13314);
nand U19398 (N_19398,N_12885,N_12134);
xor U19399 (N_19399,N_10388,N_14991);
or U19400 (N_19400,N_11943,N_10669);
nand U19401 (N_19401,N_12470,N_14374);
and U19402 (N_19402,N_13232,N_14297);
nand U19403 (N_19403,N_11328,N_13650);
or U19404 (N_19404,N_10093,N_14741);
and U19405 (N_19405,N_11267,N_11298);
nand U19406 (N_19406,N_13363,N_12397);
nand U19407 (N_19407,N_10409,N_13004);
or U19408 (N_19408,N_13560,N_13113);
nor U19409 (N_19409,N_11974,N_12007);
nor U19410 (N_19410,N_12779,N_13173);
nor U19411 (N_19411,N_14177,N_14963);
xor U19412 (N_19412,N_12482,N_11088);
xnor U19413 (N_19413,N_14414,N_10782);
and U19414 (N_19414,N_11605,N_10332);
nor U19415 (N_19415,N_10010,N_11481);
nand U19416 (N_19416,N_11476,N_14424);
or U19417 (N_19417,N_14380,N_10302);
xnor U19418 (N_19418,N_13759,N_12872);
nor U19419 (N_19419,N_12751,N_13436);
or U19420 (N_19420,N_10561,N_11182);
and U19421 (N_19421,N_10798,N_13014);
and U19422 (N_19422,N_13081,N_11245);
or U19423 (N_19423,N_12069,N_14062);
or U19424 (N_19424,N_14312,N_13441);
and U19425 (N_19425,N_12706,N_12105);
nand U19426 (N_19426,N_10419,N_12582);
nand U19427 (N_19427,N_14803,N_14046);
or U19428 (N_19428,N_13468,N_13207);
nor U19429 (N_19429,N_13472,N_14567);
and U19430 (N_19430,N_11320,N_12363);
and U19431 (N_19431,N_13369,N_10609);
nand U19432 (N_19432,N_10012,N_12751);
nand U19433 (N_19433,N_14004,N_11963);
xor U19434 (N_19434,N_11173,N_13884);
and U19435 (N_19435,N_14714,N_13119);
and U19436 (N_19436,N_13922,N_13965);
or U19437 (N_19437,N_12734,N_11339);
or U19438 (N_19438,N_13223,N_12393);
and U19439 (N_19439,N_13643,N_12155);
and U19440 (N_19440,N_11059,N_10990);
nand U19441 (N_19441,N_13663,N_11810);
or U19442 (N_19442,N_10207,N_14045);
and U19443 (N_19443,N_11217,N_10151);
or U19444 (N_19444,N_12741,N_11250);
nand U19445 (N_19445,N_14075,N_13106);
or U19446 (N_19446,N_12486,N_14924);
nand U19447 (N_19447,N_11728,N_11206);
nor U19448 (N_19448,N_12704,N_10110);
and U19449 (N_19449,N_11207,N_10447);
nand U19450 (N_19450,N_10133,N_10311);
and U19451 (N_19451,N_13523,N_13894);
nor U19452 (N_19452,N_12734,N_11431);
and U19453 (N_19453,N_13927,N_14826);
and U19454 (N_19454,N_10165,N_11201);
or U19455 (N_19455,N_12014,N_14723);
nor U19456 (N_19456,N_13666,N_10238);
and U19457 (N_19457,N_12566,N_10601);
nand U19458 (N_19458,N_11577,N_13539);
nand U19459 (N_19459,N_10006,N_14709);
or U19460 (N_19460,N_13996,N_10768);
xnor U19461 (N_19461,N_14564,N_10896);
xor U19462 (N_19462,N_11960,N_11153);
nand U19463 (N_19463,N_12865,N_12197);
nor U19464 (N_19464,N_12536,N_10575);
nand U19465 (N_19465,N_14286,N_12758);
nor U19466 (N_19466,N_13066,N_14883);
nand U19467 (N_19467,N_12902,N_10557);
nor U19468 (N_19468,N_14386,N_12469);
xnor U19469 (N_19469,N_10250,N_13534);
or U19470 (N_19470,N_11329,N_10267);
nor U19471 (N_19471,N_11587,N_10162);
nor U19472 (N_19472,N_11218,N_12436);
nand U19473 (N_19473,N_13941,N_11366);
and U19474 (N_19474,N_11464,N_14280);
xor U19475 (N_19475,N_14380,N_13814);
nor U19476 (N_19476,N_14366,N_13677);
and U19477 (N_19477,N_14482,N_10874);
nor U19478 (N_19478,N_13368,N_12517);
nor U19479 (N_19479,N_14181,N_12434);
and U19480 (N_19480,N_10012,N_11369);
or U19481 (N_19481,N_14832,N_11113);
nand U19482 (N_19482,N_10171,N_10114);
nor U19483 (N_19483,N_14620,N_10788);
nand U19484 (N_19484,N_12454,N_10508);
and U19485 (N_19485,N_13962,N_12289);
or U19486 (N_19486,N_14847,N_10980);
or U19487 (N_19487,N_14081,N_14892);
nand U19488 (N_19488,N_10475,N_14184);
nand U19489 (N_19489,N_12659,N_10029);
nor U19490 (N_19490,N_13273,N_13540);
nand U19491 (N_19491,N_13110,N_13817);
nor U19492 (N_19492,N_14596,N_13672);
or U19493 (N_19493,N_11579,N_10078);
or U19494 (N_19494,N_12020,N_13823);
and U19495 (N_19495,N_11072,N_12117);
nor U19496 (N_19496,N_13014,N_10248);
nor U19497 (N_19497,N_14244,N_10246);
nor U19498 (N_19498,N_12211,N_13522);
and U19499 (N_19499,N_11806,N_13907);
and U19500 (N_19500,N_14152,N_11588);
or U19501 (N_19501,N_10602,N_10801);
nand U19502 (N_19502,N_12139,N_14557);
nor U19503 (N_19503,N_14887,N_12506);
and U19504 (N_19504,N_11899,N_10846);
and U19505 (N_19505,N_14581,N_10745);
nor U19506 (N_19506,N_13307,N_10762);
or U19507 (N_19507,N_10488,N_10582);
nand U19508 (N_19508,N_13314,N_11271);
nor U19509 (N_19509,N_14385,N_14477);
nor U19510 (N_19510,N_13519,N_10630);
or U19511 (N_19511,N_13118,N_10158);
nand U19512 (N_19512,N_13497,N_10341);
xnor U19513 (N_19513,N_13421,N_14043);
or U19514 (N_19514,N_14304,N_10013);
nand U19515 (N_19515,N_10428,N_12722);
and U19516 (N_19516,N_13841,N_10088);
and U19517 (N_19517,N_13193,N_12162);
nand U19518 (N_19518,N_12093,N_10817);
and U19519 (N_19519,N_13022,N_11362);
xor U19520 (N_19520,N_11618,N_14927);
or U19521 (N_19521,N_13033,N_14965);
and U19522 (N_19522,N_10867,N_14413);
xor U19523 (N_19523,N_14047,N_11968);
and U19524 (N_19524,N_11372,N_11201);
or U19525 (N_19525,N_10347,N_11197);
and U19526 (N_19526,N_13392,N_12946);
or U19527 (N_19527,N_14106,N_11525);
and U19528 (N_19528,N_14936,N_10778);
nand U19529 (N_19529,N_11152,N_12425);
or U19530 (N_19530,N_14637,N_10290);
nand U19531 (N_19531,N_11342,N_11452);
nor U19532 (N_19532,N_13483,N_11380);
or U19533 (N_19533,N_11189,N_12322);
nor U19534 (N_19534,N_11892,N_12539);
nor U19535 (N_19535,N_13288,N_10477);
nor U19536 (N_19536,N_14208,N_11498);
nand U19537 (N_19537,N_12240,N_11487);
nand U19538 (N_19538,N_12115,N_12734);
or U19539 (N_19539,N_12187,N_10578);
and U19540 (N_19540,N_13166,N_10765);
nand U19541 (N_19541,N_14594,N_14761);
nor U19542 (N_19542,N_14195,N_10978);
or U19543 (N_19543,N_10988,N_13982);
nor U19544 (N_19544,N_12305,N_14577);
nor U19545 (N_19545,N_10265,N_11344);
or U19546 (N_19546,N_12884,N_12880);
nand U19547 (N_19547,N_14163,N_13133);
and U19548 (N_19548,N_10427,N_14019);
nor U19549 (N_19549,N_14226,N_12124);
and U19550 (N_19550,N_13367,N_14363);
nand U19551 (N_19551,N_14385,N_13123);
nand U19552 (N_19552,N_12970,N_13132);
nand U19553 (N_19553,N_13248,N_13582);
and U19554 (N_19554,N_14179,N_10978);
and U19555 (N_19555,N_11517,N_10308);
and U19556 (N_19556,N_11482,N_10334);
and U19557 (N_19557,N_12844,N_14434);
nor U19558 (N_19558,N_14841,N_11124);
xor U19559 (N_19559,N_11968,N_11270);
or U19560 (N_19560,N_10290,N_10912);
and U19561 (N_19561,N_10018,N_10785);
nor U19562 (N_19562,N_11176,N_13880);
nor U19563 (N_19563,N_10106,N_13810);
or U19564 (N_19564,N_13780,N_13009);
or U19565 (N_19565,N_12741,N_12795);
and U19566 (N_19566,N_13444,N_14846);
nor U19567 (N_19567,N_10085,N_12784);
nor U19568 (N_19568,N_13553,N_10346);
nand U19569 (N_19569,N_10512,N_14661);
nand U19570 (N_19570,N_12067,N_11658);
nand U19571 (N_19571,N_13782,N_11760);
nor U19572 (N_19572,N_10966,N_10911);
nand U19573 (N_19573,N_13215,N_11639);
nand U19574 (N_19574,N_11296,N_13395);
and U19575 (N_19575,N_13593,N_13460);
nand U19576 (N_19576,N_13160,N_10379);
xnor U19577 (N_19577,N_12022,N_11401);
or U19578 (N_19578,N_13628,N_10189);
xnor U19579 (N_19579,N_13408,N_10430);
nand U19580 (N_19580,N_10374,N_10484);
and U19581 (N_19581,N_14560,N_13282);
nor U19582 (N_19582,N_13320,N_11000);
and U19583 (N_19583,N_14486,N_14868);
nor U19584 (N_19584,N_11135,N_11768);
xor U19585 (N_19585,N_11641,N_10619);
xor U19586 (N_19586,N_10442,N_12627);
xnor U19587 (N_19587,N_10920,N_11236);
or U19588 (N_19588,N_14813,N_14111);
or U19589 (N_19589,N_12327,N_13333);
and U19590 (N_19590,N_10619,N_12600);
nor U19591 (N_19591,N_10575,N_11373);
or U19592 (N_19592,N_12509,N_14550);
nand U19593 (N_19593,N_14931,N_13508);
nand U19594 (N_19594,N_11376,N_14626);
nand U19595 (N_19595,N_11792,N_13562);
or U19596 (N_19596,N_12234,N_11693);
or U19597 (N_19597,N_14354,N_13796);
or U19598 (N_19598,N_10502,N_14457);
and U19599 (N_19599,N_12151,N_14714);
nor U19600 (N_19600,N_12254,N_14176);
nor U19601 (N_19601,N_10291,N_12131);
nor U19602 (N_19602,N_12566,N_11155);
or U19603 (N_19603,N_11136,N_14077);
or U19604 (N_19604,N_13426,N_12402);
nand U19605 (N_19605,N_14037,N_11161);
nand U19606 (N_19606,N_14573,N_11808);
nor U19607 (N_19607,N_12348,N_14671);
and U19608 (N_19608,N_10351,N_14714);
nand U19609 (N_19609,N_12946,N_10824);
nor U19610 (N_19610,N_12461,N_10353);
and U19611 (N_19611,N_10879,N_12831);
and U19612 (N_19612,N_13004,N_12101);
xnor U19613 (N_19613,N_14224,N_11310);
and U19614 (N_19614,N_14107,N_12615);
nand U19615 (N_19615,N_14965,N_13924);
nand U19616 (N_19616,N_13057,N_12872);
and U19617 (N_19617,N_10900,N_10491);
nand U19618 (N_19618,N_13527,N_13315);
and U19619 (N_19619,N_10414,N_11614);
xor U19620 (N_19620,N_13285,N_12727);
and U19621 (N_19621,N_11854,N_10763);
or U19622 (N_19622,N_11877,N_11467);
nor U19623 (N_19623,N_11041,N_13971);
nand U19624 (N_19624,N_12710,N_13655);
nor U19625 (N_19625,N_14252,N_11680);
and U19626 (N_19626,N_10092,N_14670);
nand U19627 (N_19627,N_14521,N_10380);
nand U19628 (N_19628,N_12835,N_14715);
and U19629 (N_19629,N_13606,N_10232);
nor U19630 (N_19630,N_14718,N_13276);
nand U19631 (N_19631,N_13167,N_10678);
or U19632 (N_19632,N_10626,N_11956);
or U19633 (N_19633,N_12100,N_13718);
nand U19634 (N_19634,N_14277,N_12620);
nor U19635 (N_19635,N_10914,N_11553);
nor U19636 (N_19636,N_13498,N_13689);
and U19637 (N_19637,N_13747,N_14683);
nand U19638 (N_19638,N_12634,N_10363);
xor U19639 (N_19639,N_13539,N_14683);
xnor U19640 (N_19640,N_10073,N_10356);
nor U19641 (N_19641,N_10569,N_11822);
and U19642 (N_19642,N_11511,N_13135);
nor U19643 (N_19643,N_10413,N_11695);
and U19644 (N_19644,N_10085,N_11793);
nand U19645 (N_19645,N_14508,N_10451);
nor U19646 (N_19646,N_12047,N_13349);
xor U19647 (N_19647,N_10239,N_14139);
xnor U19648 (N_19648,N_11129,N_12679);
or U19649 (N_19649,N_11247,N_14973);
and U19650 (N_19650,N_12079,N_13954);
nor U19651 (N_19651,N_14401,N_14286);
and U19652 (N_19652,N_11936,N_13399);
nor U19653 (N_19653,N_12066,N_14687);
nand U19654 (N_19654,N_10277,N_12900);
nor U19655 (N_19655,N_11489,N_10140);
nand U19656 (N_19656,N_12065,N_12825);
nand U19657 (N_19657,N_14503,N_11469);
or U19658 (N_19658,N_14388,N_14020);
nand U19659 (N_19659,N_11010,N_14288);
xnor U19660 (N_19660,N_10212,N_13896);
xnor U19661 (N_19661,N_13354,N_13852);
and U19662 (N_19662,N_14049,N_11170);
nand U19663 (N_19663,N_11091,N_13831);
nor U19664 (N_19664,N_11531,N_14832);
and U19665 (N_19665,N_12860,N_12330);
nor U19666 (N_19666,N_10801,N_11032);
nand U19667 (N_19667,N_11412,N_11349);
and U19668 (N_19668,N_14862,N_11044);
or U19669 (N_19669,N_14485,N_12623);
or U19670 (N_19670,N_14112,N_11565);
nand U19671 (N_19671,N_10026,N_12643);
nand U19672 (N_19672,N_14209,N_12544);
nand U19673 (N_19673,N_11157,N_11140);
nand U19674 (N_19674,N_13435,N_10948);
nor U19675 (N_19675,N_10474,N_12214);
nor U19676 (N_19676,N_13867,N_14247);
and U19677 (N_19677,N_13051,N_11232);
or U19678 (N_19678,N_11925,N_13931);
nand U19679 (N_19679,N_14938,N_14270);
xnor U19680 (N_19680,N_14361,N_11873);
nor U19681 (N_19681,N_10318,N_14537);
xnor U19682 (N_19682,N_12377,N_11252);
nor U19683 (N_19683,N_11460,N_11484);
or U19684 (N_19684,N_13687,N_13914);
nor U19685 (N_19685,N_12950,N_11889);
and U19686 (N_19686,N_11646,N_11650);
nor U19687 (N_19687,N_14646,N_10916);
nand U19688 (N_19688,N_13758,N_10733);
or U19689 (N_19689,N_12572,N_10399);
or U19690 (N_19690,N_13106,N_14875);
nor U19691 (N_19691,N_13747,N_10525);
nor U19692 (N_19692,N_14793,N_12253);
or U19693 (N_19693,N_13567,N_14143);
and U19694 (N_19694,N_14548,N_13868);
nand U19695 (N_19695,N_10036,N_14259);
or U19696 (N_19696,N_12243,N_11894);
and U19697 (N_19697,N_12862,N_11847);
and U19698 (N_19698,N_12651,N_11676);
and U19699 (N_19699,N_12689,N_13512);
or U19700 (N_19700,N_11702,N_13586);
nor U19701 (N_19701,N_13053,N_12119);
xor U19702 (N_19702,N_10682,N_11776);
nand U19703 (N_19703,N_11056,N_10505);
nor U19704 (N_19704,N_11786,N_12692);
nand U19705 (N_19705,N_14001,N_13905);
nor U19706 (N_19706,N_12590,N_14736);
and U19707 (N_19707,N_12716,N_14111);
xnor U19708 (N_19708,N_11853,N_13995);
or U19709 (N_19709,N_10920,N_14380);
nand U19710 (N_19710,N_10819,N_14860);
or U19711 (N_19711,N_14774,N_14934);
xnor U19712 (N_19712,N_11105,N_10374);
or U19713 (N_19713,N_12428,N_13622);
xnor U19714 (N_19714,N_13047,N_10788);
or U19715 (N_19715,N_14612,N_10831);
and U19716 (N_19716,N_13525,N_10920);
nor U19717 (N_19717,N_12324,N_13070);
nand U19718 (N_19718,N_13595,N_13329);
nor U19719 (N_19719,N_12469,N_14916);
nand U19720 (N_19720,N_10175,N_10118);
and U19721 (N_19721,N_12893,N_13067);
and U19722 (N_19722,N_13532,N_13758);
or U19723 (N_19723,N_11076,N_14882);
nand U19724 (N_19724,N_14465,N_12642);
and U19725 (N_19725,N_12939,N_10085);
or U19726 (N_19726,N_11156,N_12238);
or U19727 (N_19727,N_11605,N_10612);
nor U19728 (N_19728,N_12161,N_10949);
nor U19729 (N_19729,N_10466,N_12673);
nor U19730 (N_19730,N_10844,N_14974);
and U19731 (N_19731,N_13111,N_13327);
nand U19732 (N_19732,N_13481,N_11900);
nor U19733 (N_19733,N_10164,N_10587);
and U19734 (N_19734,N_11136,N_13675);
xor U19735 (N_19735,N_13406,N_12986);
xnor U19736 (N_19736,N_10514,N_11757);
nor U19737 (N_19737,N_11883,N_10855);
or U19738 (N_19738,N_10295,N_14459);
nand U19739 (N_19739,N_14633,N_12006);
nor U19740 (N_19740,N_11752,N_10603);
nor U19741 (N_19741,N_14654,N_11936);
and U19742 (N_19742,N_14346,N_10915);
and U19743 (N_19743,N_11215,N_10212);
and U19744 (N_19744,N_12843,N_13282);
and U19745 (N_19745,N_12242,N_11447);
xnor U19746 (N_19746,N_12126,N_10583);
nor U19747 (N_19747,N_14076,N_14638);
or U19748 (N_19748,N_12144,N_14658);
or U19749 (N_19749,N_11172,N_13880);
nor U19750 (N_19750,N_13518,N_13073);
nor U19751 (N_19751,N_11968,N_13502);
or U19752 (N_19752,N_14991,N_13024);
and U19753 (N_19753,N_11017,N_10648);
or U19754 (N_19754,N_11485,N_11375);
nor U19755 (N_19755,N_13274,N_14578);
or U19756 (N_19756,N_13119,N_12782);
nand U19757 (N_19757,N_11164,N_13096);
nand U19758 (N_19758,N_14233,N_11119);
and U19759 (N_19759,N_12314,N_11731);
xnor U19760 (N_19760,N_12638,N_10076);
xor U19761 (N_19761,N_11800,N_13632);
xor U19762 (N_19762,N_14602,N_14274);
xor U19763 (N_19763,N_14999,N_14913);
or U19764 (N_19764,N_14960,N_13170);
nor U19765 (N_19765,N_12938,N_10915);
or U19766 (N_19766,N_12003,N_13189);
nand U19767 (N_19767,N_10215,N_14157);
nand U19768 (N_19768,N_10659,N_10878);
nor U19769 (N_19769,N_11268,N_11211);
nand U19770 (N_19770,N_11531,N_10050);
nor U19771 (N_19771,N_14624,N_11354);
and U19772 (N_19772,N_10370,N_12293);
xor U19773 (N_19773,N_14607,N_13792);
xnor U19774 (N_19774,N_13996,N_11676);
nand U19775 (N_19775,N_12704,N_11591);
and U19776 (N_19776,N_14981,N_12524);
nor U19777 (N_19777,N_14485,N_13736);
or U19778 (N_19778,N_14149,N_14820);
nand U19779 (N_19779,N_13690,N_11341);
or U19780 (N_19780,N_13270,N_12315);
and U19781 (N_19781,N_13464,N_12219);
or U19782 (N_19782,N_12826,N_10470);
xor U19783 (N_19783,N_14241,N_10163);
and U19784 (N_19784,N_13376,N_10304);
or U19785 (N_19785,N_11114,N_10206);
or U19786 (N_19786,N_10750,N_10289);
or U19787 (N_19787,N_11568,N_12288);
xnor U19788 (N_19788,N_10720,N_14856);
nand U19789 (N_19789,N_12201,N_13664);
and U19790 (N_19790,N_10585,N_11006);
or U19791 (N_19791,N_11686,N_11881);
and U19792 (N_19792,N_14090,N_14022);
nand U19793 (N_19793,N_10837,N_10874);
xor U19794 (N_19794,N_10280,N_14174);
nor U19795 (N_19795,N_13940,N_10286);
nor U19796 (N_19796,N_12593,N_10748);
and U19797 (N_19797,N_12850,N_12954);
xor U19798 (N_19798,N_13153,N_13759);
and U19799 (N_19799,N_14090,N_13172);
nor U19800 (N_19800,N_13339,N_14706);
or U19801 (N_19801,N_12319,N_12808);
and U19802 (N_19802,N_14548,N_10685);
nor U19803 (N_19803,N_11718,N_10762);
nor U19804 (N_19804,N_13342,N_13087);
nand U19805 (N_19805,N_13878,N_11413);
or U19806 (N_19806,N_13672,N_12496);
and U19807 (N_19807,N_11807,N_14795);
nand U19808 (N_19808,N_11168,N_11717);
or U19809 (N_19809,N_10749,N_13937);
xnor U19810 (N_19810,N_12196,N_10205);
and U19811 (N_19811,N_10645,N_12744);
nor U19812 (N_19812,N_10157,N_11003);
or U19813 (N_19813,N_10732,N_10816);
and U19814 (N_19814,N_13415,N_10350);
nand U19815 (N_19815,N_12695,N_13643);
or U19816 (N_19816,N_14346,N_14025);
xor U19817 (N_19817,N_10251,N_13886);
nand U19818 (N_19818,N_13225,N_14130);
nand U19819 (N_19819,N_12436,N_10862);
xor U19820 (N_19820,N_12613,N_10220);
nand U19821 (N_19821,N_11581,N_13707);
nand U19822 (N_19822,N_14432,N_13394);
or U19823 (N_19823,N_12433,N_14940);
and U19824 (N_19824,N_13930,N_11435);
and U19825 (N_19825,N_13261,N_12275);
and U19826 (N_19826,N_10875,N_11459);
nor U19827 (N_19827,N_12935,N_14881);
nand U19828 (N_19828,N_12073,N_14608);
nor U19829 (N_19829,N_13074,N_13223);
or U19830 (N_19830,N_12457,N_12767);
nor U19831 (N_19831,N_12406,N_14773);
or U19832 (N_19832,N_10249,N_14670);
nor U19833 (N_19833,N_14702,N_12865);
nor U19834 (N_19834,N_11226,N_12421);
and U19835 (N_19835,N_11727,N_13158);
nor U19836 (N_19836,N_11953,N_12519);
or U19837 (N_19837,N_12996,N_10028);
xor U19838 (N_19838,N_14679,N_13695);
nor U19839 (N_19839,N_10139,N_14094);
and U19840 (N_19840,N_14061,N_12905);
nand U19841 (N_19841,N_11263,N_14092);
and U19842 (N_19842,N_13483,N_13725);
nor U19843 (N_19843,N_10630,N_14323);
nand U19844 (N_19844,N_14107,N_10391);
or U19845 (N_19845,N_14986,N_10615);
nand U19846 (N_19846,N_13915,N_12316);
xnor U19847 (N_19847,N_11434,N_12566);
and U19848 (N_19848,N_11804,N_12177);
and U19849 (N_19849,N_11167,N_12715);
nor U19850 (N_19850,N_14150,N_14579);
and U19851 (N_19851,N_13281,N_13983);
and U19852 (N_19852,N_12208,N_11475);
and U19853 (N_19853,N_12610,N_11033);
or U19854 (N_19854,N_12740,N_10847);
xnor U19855 (N_19855,N_10764,N_14882);
nor U19856 (N_19856,N_10159,N_12803);
or U19857 (N_19857,N_11701,N_13522);
nor U19858 (N_19858,N_10389,N_14970);
xor U19859 (N_19859,N_12166,N_12729);
and U19860 (N_19860,N_11023,N_14801);
and U19861 (N_19861,N_10089,N_13560);
nand U19862 (N_19862,N_12023,N_14451);
xor U19863 (N_19863,N_11973,N_14446);
nand U19864 (N_19864,N_13561,N_13643);
nor U19865 (N_19865,N_13698,N_14521);
xor U19866 (N_19866,N_11320,N_14932);
nor U19867 (N_19867,N_11235,N_11820);
and U19868 (N_19868,N_12438,N_10079);
nand U19869 (N_19869,N_14613,N_13511);
or U19870 (N_19870,N_12320,N_14243);
nand U19871 (N_19871,N_11691,N_14764);
xor U19872 (N_19872,N_10204,N_13177);
nor U19873 (N_19873,N_10275,N_12099);
or U19874 (N_19874,N_13292,N_13010);
or U19875 (N_19875,N_11621,N_14745);
and U19876 (N_19876,N_11656,N_10014);
nand U19877 (N_19877,N_11988,N_13556);
nor U19878 (N_19878,N_12811,N_11056);
nand U19879 (N_19879,N_13605,N_13114);
xor U19880 (N_19880,N_11005,N_10663);
and U19881 (N_19881,N_11407,N_10121);
xnor U19882 (N_19882,N_13312,N_12870);
and U19883 (N_19883,N_11349,N_10095);
nor U19884 (N_19884,N_10999,N_12935);
nand U19885 (N_19885,N_14986,N_10948);
xor U19886 (N_19886,N_11723,N_13243);
and U19887 (N_19887,N_11753,N_13235);
or U19888 (N_19888,N_11184,N_10163);
and U19889 (N_19889,N_13564,N_11525);
and U19890 (N_19890,N_12798,N_14110);
or U19891 (N_19891,N_12407,N_11097);
nand U19892 (N_19892,N_11145,N_12171);
nand U19893 (N_19893,N_12960,N_11442);
nor U19894 (N_19894,N_12964,N_12725);
and U19895 (N_19895,N_13037,N_12913);
nand U19896 (N_19896,N_10711,N_14787);
and U19897 (N_19897,N_11267,N_14440);
nor U19898 (N_19898,N_10883,N_14855);
or U19899 (N_19899,N_13120,N_13239);
nor U19900 (N_19900,N_14392,N_14365);
xnor U19901 (N_19901,N_11089,N_14630);
and U19902 (N_19902,N_12685,N_11711);
nand U19903 (N_19903,N_11972,N_14395);
and U19904 (N_19904,N_14337,N_11833);
nand U19905 (N_19905,N_13230,N_13602);
nor U19906 (N_19906,N_10471,N_13651);
and U19907 (N_19907,N_13336,N_14801);
nor U19908 (N_19908,N_11940,N_12060);
xnor U19909 (N_19909,N_14913,N_10898);
or U19910 (N_19910,N_12862,N_12854);
xnor U19911 (N_19911,N_11116,N_10665);
nor U19912 (N_19912,N_12683,N_13937);
nand U19913 (N_19913,N_12182,N_11278);
and U19914 (N_19914,N_12620,N_10143);
nand U19915 (N_19915,N_11464,N_13690);
and U19916 (N_19916,N_13455,N_10963);
and U19917 (N_19917,N_13918,N_13884);
nor U19918 (N_19918,N_10398,N_11485);
nor U19919 (N_19919,N_12450,N_13186);
and U19920 (N_19920,N_13098,N_14288);
nand U19921 (N_19921,N_14118,N_13472);
nand U19922 (N_19922,N_14837,N_11797);
or U19923 (N_19923,N_11289,N_10959);
nand U19924 (N_19924,N_14715,N_11527);
or U19925 (N_19925,N_12422,N_14450);
nor U19926 (N_19926,N_11759,N_12958);
and U19927 (N_19927,N_14844,N_14102);
nor U19928 (N_19928,N_11819,N_13417);
nor U19929 (N_19929,N_10203,N_11687);
nand U19930 (N_19930,N_13918,N_12148);
and U19931 (N_19931,N_10808,N_13505);
nor U19932 (N_19932,N_14772,N_11639);
or U19933 (N_19933,N_13572,N_10724);
or U19934 (N_19934,N_12923,N_14385);
and U19935 (N_19935,N_14935,N_13011);
and U19936 (N_19936,N_10142,N_13812);
and U19937 (N_19937,N_13620,N_10856);
nor U19938 (N_19938,N_11683,N_10137);
and U19939 (N_19939,N_11219,N_13653);
or U19940 (N_19940,N_11124,N_11569);
nand U19941 (N_19941,N_10033,N_10272);
nand U19942 (N_19942,N_10242,N_11279);
or U19943 (N_19943,N_12239,N_10759);
xnor U19944 (N_19944,N_10067,N_14272);
or U19945 (N_19945,N_10797,N_13842);
and U19946 (N_19946,N_13082,N_13612);
nand U19947 (N_19947,N_12790,N_12387);
or U19948 (N_19948,N_13052,N_11957);
nor U19949 (N_19949,N_12654,N_10110);
nor U19950 (N_19950,N_11888,N_14660);
and U19951 (N_19951,N_13155,N_10299);
nand U19952 (N_19952,N_10760,N_13282);
or U19953 (N_19953,N_12497,N_10688);
nand U19954 (N_19954,N_13158,N_11182);
nand U19955 (N_19955,N_12035,N_12656);
nand U19956 (N_19956,N_12597,N_14036);
nor U19957 (N_19957,N_10108,N_12257);
or U19958 (N_19958,N_10808,N_10814);
or U19959 (N_19959,N_13451,N_12648);
or U19960 (N_19960,N_11625,N_10037);
or U19961 (N_19961,N_11221,N_11559);
and U19962 (N_19962,N_14622,N_11688);
xor U19963 (N_19963,N_13481,N_10253);
or U19964 (N_19964,N_13554,N_10125);
or U19965 (N_19965,N_13387,N_13993);
nor U19966 (N_19966,N_13291,N_10555);
nand U19967 (N_19967,N_13809,N_13262);
and U19968 (N_19968,N_10354,N_10169);
and U19969 (N_19969,N_12044,N_12086);
and U19970 (N_19970,N_10515,N_10993);
nor U19971 (N_19971,N_14312,N_14716);
and U19972 (N_19972,N_12955,N_10759);
or U19973 (N_19973,N_13352,N_11512);
or U19974 (N_19974,N_12038,N_13407);
or U19975 (N_19975,N_10489,N_10870);
and U19976 (N_19976,N_13737,N_12019);
nor U19977 (N_19977,N_13153,N_13836);
xor U19978 (N_19978,N_13060,N_12860);
or U19979 (N_19979,N_12850,N_10750);
or U19980 (N_19980,N_11009,N_12118);
nor U19981 (N_19981,N_11626,N_10943);
nor U19982 (N_19982,N_12278,N_13382);
nand U19983 (N_19983,N_13456,N_13416);
nand U19984 (N_19984,N_10921,N_13484);
and U19985 (N_19985,N_14100,N_12271);
nand U19986 (N_19986,N_12323,N_13540);
nor U19987 (N_19987,N_14632,N_12971);
and U19988 (N_19988,N_10412,N_12305);
and U19989 (N_19989,N_14819,N_12351);
nand U19990 (N_19990,N_13125,N_12204);
nand U19991 (N_19991,N_10129,N_11200);
nor U19992 (N_19992,N_13759,N_14220);
xnor U19993 (N_19993,N_14168,N_13007);
and U19994 (N_19994,N_13195,N_11286);
and U19995 (N_19995,N_12257,N_14844);
or U19996 (N_19996,N_13834,N_12771);
and U19997 (N_19997,N_10198,N_10086);
or U19998 (N_19998,N_11144,N_14204);
nand U19999 (N_19999,N_10224,N_10220);
nand U20000 (N_20000,N_18266,N_18320);
nand U20001 (N_20001,N_15194,N_15861);
or U20002 (N_20002,N_17461,N_18608);
and U20003 (N_20003,N_19462,N_19415);
nand U20004 (N_20004,N_17655,N_15167);
nor U20005 (N_20005,N_15310,N_15717);
and U20006 (N_20006,N_16505,N_17764);
and U20007 (N_20007,N_15026,N_17545);
nor U20008 (N_20008,N_17557,N_17455);
and U20009 (N_20009,N_16141,N_17847);
and U20010 (N_20010,N_17841,N_17698);
nor U20011 (N_20011,N_15686,N_17578);
nor U20012 (N_20012,N_15363,N_15147);
or U20013 (N_20013,N_17292,N_19589);
nand U20014 (N_20014,N_17616,N_18431);
or U20015 (N_20015,N_18424,N_18255);
nand U20016 (N_20016,N_16076,N_16892);
and U20017 (N_20017,N_19512,N_15777);
and U20018 (N_20018,N_16780,N_19228);
nor U20019 (N_20019,N_19286,N_17444);
and U20020 (N_20020,N_16026,N_17315);
xnor U20021 (N_20021,N_16073,N_16009);
xnor U20022 (N_20022,N_15198,N_15055);
and U20023 (N_20023,N_17185,N_18175);
xor U20024 (N_20024,N_15778,N_15364);
or U20025 (N_20025,N_18218,N_18108);
nor U20026 (N_20026,N_15884,N_18138);
nand U20027 (N_20027,N_19197,N_19143);
or U20028 (N_20028,N_17555,N_19081);
nand U20029 (N_20029,N_15422,N_16305);
nand U20030 (N_20030,N_19435,N_16262);
nor U20031 (N_20031,N_17117,N_15452);
nor U20032 (N_20032,N_17833,N_18500);
or U20033 (N_20033,N_19434,N_15920);
and U20034 (N_20034,N_17222,N_16720);
nor U20035 (N_20035,N_15866,N_16735);
nand U20036 (N_20036,N_16713,N_18678);
or U20037 (N_20037,N_15744,N_18134);
xnor U20038 (N_20038,N_19674,N_19693);
nor U20039 (N_20039,N_18271,N_16559);
or U20040 (N_20040,N_19099,N_16999);
or U20041 (N_20041,N_16702,N_17992);
or U20042 (N_20042,N_18735,N_17425);
or U20043 (N_20043,N_18570,N_17267);
or U20044 (N_20044,N_17167,N_19854);
nand U20045 (N_20045,N_19256,N_17345);
nor U20046 (N_20046,N_19546,N_19118);
and U20047 (N_20047,N_15666,N_19931);
nand U20048 (N_20048,N_18957,N_18044);
or U20049 (N_20049,N_17807,N_18171);
nand U20050 (N_20050,N_19743,N_15405);
nand U20051 (N_20051,N_15819,N_18118);
or U20052 (N_20052,N_17101,N_16056);
nand U20053 (N_20053,N_16164,N_16178);
and U20054 (N_20054,N_17349,N_17361);
nor U20055 (N_20055,N_17058,N_17308);
nand U20056 (N_20056,N_17115,N_17027);
or U20057 (N_20057,N_18600,N_16504);
nor U20058 (N_20058,N_17155,N_18699);
or U20059 (N_20059,N_18212,N_15530);
or U20060 (N_20060,N_15289,N_18144);
xor U20061 (N_20061,N_19588,N_19810);
xnor U20062 (N_20062,N_18596,N_15970);
or U20063 (N_20063,N_18301,N_17376);
nor U20064 (N_20064,N_19889,N_16616);
and U20065 (N_20065,N_15757,N_16240);
and U20066 (N_20066,N_19032,N_18777);
or U20067 (N_20067,N_16339,N_16771);
nor U20068 (N_20068,N_19597,N_17529);
nand U20069 (N_20069,N_17503,N_18952);
nor U20070 (N_20070,N_18421,N_17662);
nor U20071 (N_20071,N_17339,N_19365);
or U20072 (N_20072,N_17424,N_19994);
nor U20073 (N_20073,N_17598,N_17687);
xor U20074 (N_20074,N_17796,N_16923);
xor U20075 (N_20075,N_17596,N_15814);
or U20076 (N_20076,N_19425,N_17776);
xor U20077 (N_20077,N_18286,N_18420);
or U20078 (N_20078,N_15645,N_19928);
xor U20079 (N_20079,N_19431,N_15513);
or U20080 (N_20080,N_16572,N_17128);
and U20081 (N_20081,N_15285,N_18230);
nor U20082 (N_20082,N_17245,N_18644);
nand U20083 (N_20083,N_17443,N_15996);
and U20084 (N_20084,N_16942,N_17287);
and U20085 (N_20085,N_15320,N_15622);
or U20086 (N_20086,N_18261,N_17131);
nor U20087 (N_20087,N_16567,N_16819);
or U20088 (N_20088,N_18358,N_17237);
nor U20089 (N_20089,N_19873,N_15112);
or U20090 (N_20090,N_15114,N_16740);
xor U20091 (N_20091,N_16365,N_18476);
nand U20092 (N_20092,N_16225,N_17886);
or U20093 (N_20093,N_19142,N_15955);
nor U20094 (N_20094,N_16621,N_19257);
nand U20095 (N_20095,N_15252,N_18976);
and U20096 (N_20096,N_19074,N_16871);
or U20097 (N_20097,N_18155,N_16647);
xor U20098 (N_20098,N_19221,N_17572);
or U20099 (N_20099,N_19281,N_19399);
or U20100 (N_20100,N_18438,N_17338);
nand U20101 (N_20101,N_16751,N_15150);
xor U20102 (N_20102,N_17755,N_17613);
nor U20103 (N_20103,N_16238,N_18088);
nor U20104 (N_20104,N_16765,N_15837);
nor U20105 (N_20105,N_15450,N_17102);
or U20106 (N_20106,N_17928,N_17683);
and U20107 (N_20107,N_17576,N_15376);
nor U20108 (N_20108,N_15362,N_16644);
or U20109 (N_20109,N_15346,N_16553);
nor U20110 (N_20110,N_16380,N_17138);
nand U20111 (N_20111,N_18089,N_19944);
or U20112 (N_20112,N_18677,N_16868);
or U20113 (N_20113,N_17047,N_15807);
or U20114 (N_20114,N_18705,N_17408);
nand U20115 (N_20115,N_15143,N_15294);
nor U20116 (N_20116,N_18270,N_18714);
nand U20117 (N_20117,N_16637,N_15343);
nand U20118 (N_20118,N_16784,N_17031);
nor U20119 (N_20119,N_16781,N_17855);
nand U20120 (N_20120,N_15015,N_15742);
or U20121 (N_20121,N_16612,N_16851);
nor U20122 (N_20122,N_17920,N_16040);
nand U20123 (N_20123,N_18321,N_15224);
nand U20124 (N_20124,N_16890,N_16326);
nor U20125 (N_20125,N_18656,N_16375);
nand U20126 (N_20126,N_19710,N_18776);
nor U20127 (N_20127,N_16102,N_19863);
nand U20128 (N_20128,N_19183,N_16261);
or U20129 (N_20129,N_15813,N_19219);
nor U20130 (N_20130,N_19059,N_19877);
or U20131 (N_20131,N_16427,N_19305);
or U20132 (N_20132,N_16506,N_16476);
and U20133 (N_20133,N_16709,N_15284);
xnor U20134 (N_20134,N_19922,N_15020);
and U20135 (N_20135,N_18759,N_18835);
nor U20136 (N_20136,N_16246,N_18703);
nor U20137 (N_20137,N_19622,N_17180);
nor U20138 (N_20138,N_17175,N_17092);
nand U20139 (N_20139,N_17211,N_16747);
and U20140 (N_20140,N_17740,N_17103);
and U20141 (N_20141,N_15215,N_15541);
nand U20142 (N_20142,N_15503,N_16241);
nor U20143 (N_20143,N_18026,N_17984);
or U20144 (N_20144,N_15873,N_19000);
or U20145 (N_20145,N_16194,N_16005);
nor U20146 (N_20146,N_17141,N_17804);
nor U20147 (N_20147,N_19279,N_17696);
nor U20148 (N_20148,N_16383,N_15061);
or U20149 (N_20149,N_16137,N_15738);
nor U20150 (N_20150,N_17769,N_17889);
nor U20151 (N_20151,N_16229,N_16301);
nor U20152 (N_20152,N_18145,N_17643);
and U20153 (N_20153,N_15132,N_17261);
or U20154 (N_20154,N_16158,N_18281);
nand U20155 (N_20155,N_17333,N_15269);
and U20156 (N_20156,N_19720,N_18045);
nand U20157 (N_20157,N_16046,N_17617);
nor U20158 (N_20158,N_16843,N_17157);
nor U20159 (N_20159,N_19429,N_16617);
nor U20160 (N_20160,N_19442,N_16530);
or U20161 (N_20161,N_16988,N_18302);
nor U20162 (N_20162,N_19656,N_15011);
xor U20163 (N_20163,N_15312,N_19215);
or U20164 (N_20164,N_17913,N_17156);
or U20165 (N_20165,N_17232,N_17961);
and U20166 (N_20166,N_15368,N_19995);
nor U20167 (N_20167,N_18824,N_19816);
or U20168 (N_20168,N_17093,N_17347);
and U20169 (N_20169,N_19650,N_15382);
and U20170 (N_20170,N_19340,N_15504);
nand U20171 (N_20171,N_16602,N_15108);
nand U20172 (N_20172,N_17471,N_15766);
or U20173 (N_20173,N_17016,N_19382);
nor U20174 (N_20174,N_17812,N_16521);
nand U20175 (N_20175,N_16269,N_19735);
and U20176 (N_20176,N_17989,N_19213);
and U20177 (N_20177,N_15602,N_16543);
nand U20178 (N_20178,N_16822,N_15942);
nor U20179 (N_20179,N_17709,N_19445);
nor U20180 (N_20180,N_15389,N_18225);
xnor U20181 (N_20181,N_16223,N_17309);
or U20182 (N_20182,N_19273,N_19369);
or U20183 (N_20183,N_17594,N_15037);
nand U20184 (N_20184,N_17149,N_17607);
nor U20185 (N_20185,N_19262,N_16882);
nand U20186 (N_20186,N_17041,N_19869);
nor U20187 (N_20187,N_17561,N_15303);
nor U20188 (N_20188,N_18490,N_16609);
nand U20189 (N_20189,N_18534,N_15505);
and U20190 (N_20190,N_16640,N_19144);
or U20191 (N_20191,N_18662,N_15148);
nand U20192 (N_20192,N_15924,N_18411);
or U20193 (N_20193,N_17351,N_17482);
or U20194 (N_20194,N_15073,N_19677);
or U20195 (N_20195,N_16251,N_18517);
nand U20196 (N_20196,N_19456,N_19130);
nand U20197 (N_20197,N_16214,N_17700);
or U20198 (N_20198,N_15954,N_19073);
or U20199 (N_20199,N_16101,N_17467);
and U20200 (N_20200,N_16408,N_19819);
nor U20201 (N_20201,N_18012,N_18400);
nand U20202 (N_20202,N_18936,N_17303);
nor U20203 (N_20203,N_18993,N_16247);
nor U20204 (N_20204,N_16212,N_17204);
xnor U20205 (N_20205,N_17690,N_18037);
or U20206 (N_20206,N_18780,N_17685);
xnor U20207 (N_20207,N_17898,N_18808);
and U20208 (N_20208,N_19530,N_15975);
or U20209 (N_20209,N_17972,N_16025);
nand U20210 (N_20210,N_19827,N_18602);
and U20211 (N_20211,N_16985,N_16224);
nor U20212 (N_20212,N_15518,N_15542);
nand U20213 (N_20213,N_18278,N_15336);
xnor U20214 (N_20214,N_18629,N_15756);
or U20215 (N_20215,N_18177,N_17669);
or U20216 (N_20216,N_17476,N_16850);
nor U20217 (N_20217,N_19736,N_15980);
nor U20218 (N_20218,N_17739,N_17551);
nor U20219 (N_20219,N_15180,N_18469);
nand U20220 (N_20220,N_19623,N_19439);
nor U20221 (N_20221,N_19111,N_18067);
and U20222 (N_20222,N_15759,N_19586);
nor U20223 (N_20223,N_17895,N_19829);
nor U20224 (N_20224,N_17066,N_17853);
and U20225 (N_20225,N_19420,N_18645);
nor U20226 (N_20226,N_17049,N_17571);
and U20227 (N_20227,N_15072,N_19480);
xnor U20228 (N_20228,N_16179,N_15973);
nand U20229 (N_20229,N_17194,N_18539);
and U20230 (N_20230,N_19204,N_16239);
and U20231 (N_20231,N_17866,N_17534);
nor U20232 (N_20232,N_15120,N_15292);
nor U20233 (N_20233,N_19721,N_17910);
xor U20234 (N_20234,N_16296,N_15893);
nor U20235 (N_20235,N_18484,N_19835);
and U20236 (N_20236,N_16936,N_15386);
and U20237 (N_20237,N_17845,N_16154);
xnor U20238 (N_20238,N_16727,N_16584);
or U20239 (N_20239,N_18744,N_16711);
nand U20240 (N_20240,N_18240,N_17808);
nor U20241 (N_20241,N_15181,N_15403);
or U20242 (N_20242,N_18130,N_16688);
nor U20243 (N_20243,N_16472,N_17635);
nor U20244 (N_20244,N_17137,N_15302);
nand U20245 (N_20245,N_17146,N_18226);
or U20246 (N_20246,N_19632,N_18343);
nand U20247 (N_20247,N_16067,N_18363);
nor U20248 (N_20248,N_17625,N_17849);
nor U20249 (N_20249,N_15624,N_17311);
nand U20250 (N_20250,N_18844,N_18870);
nor U20251 (N_20251,N_19428,N_15628);
nor U20252 (N_20252,N_17198,N_15159);
nor U20253 (N_20253,N_15609,N_18879);
nand U20254 (N_20254,N_19063,N_17404);
nand U20255 (N_20255,N_15959,N_19754);
and U20256 (N_20256,N_15088,N_18625);
nand U20257 (N_20257,N_17507,N_15221);
nor U20258 (N_20258,N_18918,N_17905);
nand U20259 (N_20259,N_18296,N_19903);
or U20260 (N_20260,N_18527,N_16187);
or U20261 (N_20261,N_18196,N_19357);
or U20262 (N_20262,N_16366,N_15111);
nor U20263 (N_20263,N_16719,N_17417);
or U20264 (N_20264,N_16945,N_19795);
or U20265 (N_20265,N_17054,N_17521);
nand U20266 (N_20266,N_15477,N_19946);
or U20267 (N_20267,N_18084,N_18405);
and U20268 (N_20268,N_15634,N_19606);
nor U20269 (N_20269,N_17619,N_18081);
and U20270 (N_20270,N_18273,N_16461);
or U20271 (N_20271,N_15431,N_19745);
nor U20272 (N_20272,N_16157,N_18821);
nor U20273 (N_20273,N_15459,N_19564);
nand U20274 (N_20274,N_19274,N_15806);
or U20275 (N_20275,N_15649,N_15187);
or U20276 (N_20276,N_17336,N_16079);
or U20277 (N_20277,N_15656,N_17178);
nor U20278 (N_20278,N_16113,N_16695);
and U20279 (N_20279,N_16032,N_19297);
nor U20280 (N_20280,N_17676,N_16353);
or U20281 (N_20281,N_17238,N_19731);
nand U20282 (N_20282,N_18298,N_19510);
xor U20283 (N_20283,N_18021,N_19291);
xor U20284 (N_20284,N_19621,N_15056);
and U20285 (N_20285,N_15877,N_18838);
and U20286 (N_20286,N_18640,N_16974);
nor U20287 (N_20287,N_17753,N_16117);
or U20288 (N_20288,N_18519,N_16313);
xnor U20289 (N_20289,N_15435,N_15486);
and U20290 (N_20290,N_15463,N_19545);
nand U20291 (N_20291,N_18324,N_15022);
or U20292 (N_20292,N_16089,N_19595);
nor U20293 (N_20293,N_18943,N_17481);
and U20294 (N_20294,N_16317,N_19051);
and U20295 (N_20295,N_15370,N_19106);
and U20296 (N_20296,N_17565,N_19114);
xor U20297 (N_20297,N_18435,N_19540);
nor U20298 (N_20298,N_18325,N_18911);
and U20299 (N_20299,N_16512,N_17713);
and U20300 (N_20300,N_19767,N_18949);
and U20301 (N_20301,N_16222,N_18079);
or U20302 (N_20302,N_16155,N_16260);
and U20303 (N_20303,N_19568,N_17884);
nand U20304 (N_20304,N_16166,N_15988);
nand U20305 (N_20305,N_15296,N_18720);
nor U20306 (N_20306,N_17968,N_18091);
or U20307 (N_20307,N_16674,N_19047);
nor U20308 (N_20308,N_16038,N_18365);
nor U20309 (N_20309,N_17053,N_18554);
xor U20310 (N_20310,N_17241,N_16970);
nor U20311 (N_20311,N_17527,N_19951);
or U20312 (N_20312,N_15616,N_18001);
xor U20313 (N_20313,N_15745,N_18573);
nand U20314 (N_20314,N_16110,N_19255);
nand U20315 (N_20315,N_19940,N_18087);
and U20316 (N_20316,N_17380,N_17878);
nand U20317 (N_20317,N_19970,N_17078);
nand U20318 (N_20318,N_17597,N_17486);
or U20319 (N_20319,N_15171,N_18074);
or U20320 (N_20320,N_19070,N_18467);
and U20321 (N_20321,N_19925,N_19140);
nor U20322 (N_20322,N_16107,N_15276);
nand U20323 (N_20323,N_18763,N_19726);
nand U20324 (N_20324,N_15694,N_19068);
nor U20325 (N_20325,N_18912,N_18509);
or U20326 (N_20326,N_18470,N_15933);
nand U20327 (N_20327,N_15870,N_17842);
nand U20328 (N_20328,N_19402,N_18101);
and U20329 (N_20329,N_16959,N_16561);
nor U20330 (N_20330,N_18452,N_16714);
nand U20331 (N_20331,N_16129,N_15724);
and U20332 (N_20332,N_15493,N_16675);
nand U20333 (N_20333,N_19179,N_18425);
nor U20334 (N_20334,N_17663,N_19645);
xor U20335 (N_20335,N_19284,N_18129);
xnor U20336 (N_20336,N_15544,N_15981);
and U20337 (N_20337,N_16350,N_16569);
nor U20338 (N_20338,N_15581,N_19129);
and U20339 (N_20339,N_15938,N_19498);
or U20340 (N_20340,N_16918,N_19772);
nand U20341 (N_20341,N_15726,N_15208);
or U20342 (N_20342,N_19108,N_19690);
and U20343 (N_20343,N_19527,N_16642);
nor U20344 (N_20344,N_16883,N_16455);
nand U20345 (N_20345,N_18607,N_18231);
xnor U20346 (N_20346,N_18217,N_17298);
or U20347 (N_20347,N_18981,N_15566);
nor U20348 (N_20348,N_18475,N_16663);
nor U20349 (N_20349,N_18430,N_16968);
or U20350 (N_20350,N_16797,N_18820);
xor U20351 (N_20351,N_18741,N_19804);
xnor U20352 (N_20352,N_16095,N_19594);
xnor U20353 (N_20353,N_16904,N_19796);
nor U20354 (N_20354,N_19160,N_15484);
or U20355 (N_20355,N_18034,N_17327);
nor U20356 (N_20356,N_19296,N_18956);
or U20357 (N_20357,N_15764,N_16285);
nor U20358 (N_20358,N_18288,N_18190);
nand U20359 (N_20359,N_19153,N_19571);
nor U20360 (N_20360,N_15188,N_17415);
and U20361 (N_20361,N_16862,N_15019);
or U20362 (N_20362,N_17391,N_15502);
nor U20363 (N_20363,N_19201,N_16947);
nor U20364 (N_20364,N_19189,N_19393);
nand U20365 (N_20365,N_19906,N_18942);
nor U20366 (N_20366,N_15400,N_17276);
nand U20367 (N_20367,N_17280,N_18841);
or U20368 (N_20368,N_18022,N_17544);
nand U20369 (N_20369,N_19939,N_19843);
nand U20370 (N_20370,N_18622,N_18098);
or U20371 (N_20371,N_19227,N_17464);
and U20372 (N_20372,N_15586,N_16354);
or U20373 (N_20373,N_18536,N_19603);
or U20374 (N_20374,N_16703,N_15990);
nor U20375 (N_20375,N_19737,N_19006);
nand U20376 (N_20376,N_19563,N_16895);
nand U20377 (N_20377,N_17026,N_15474);
nor U20378 (N_20378,N_17290,N_19045);
nor U20379 (N_20379,N_18221,N_17414);
and U20380 (N_20380,N_16308,N_18878);
or U20381 (N_20381,N_15371,N_18392);
and U20382 (N_20382,N_18786,N_16123);
nand U20383 (N_20383,N_16516,N_15106);
nor U20384 (N_20384,N_15115,N_17472);
and U20385 (N_20385,N_16277,N_15149);
nor U20386 (N_20386,N_18888,N_15688);
nand U20387 (N_20387,N_17019,N_17580);
or U20388 (N_20388,N_18069,N_18201);
or U20389 (N_20389,N_18024,N_16048);
nand U20390 (N_20390,N_17973,N_17400);
nand U20391 (N_20391,N_18347,N_17749);
nand U20392 (N_20392,N_17612,N_16293);
xnor U20393 (N_20393,N_17838,N_18446);
and U20394 (N_20394,N_18845,N_17570);
nor U20395 (N_20395,N_16436,N_15632);
or U20396 (N_20396,N_18303,N_19358);
or U20397 (N_20397,N_17939,N_18334);
xnor U20398 (N_20398,N_19131,N_17823);
and U20399 (N_20399,N_18611,N_18974);
nor U20400 (N_20400,N_19789,N_17403);
nand U20401 (N_20401,N_17653,N_18589);
nor U20402 (N_20402,N_15300,N_17517);
nand U20403 (N_20403,N_19018,N_15153);
and U20404 (N_20404,N_18711,N_15126);
nor U20405 (N_20405,N_16651,N_19384);
nor U20406 (N_20406,N_15233,N_19739);
and U20407 (N_20407,N_16481,N_16980);
and U20408 (N_20408,N_18259,N_19790);
and U20409 (N_20409,N_19845,N_18373);
and U20410 (N_20410,N_18983,N_17456);
or U20411 (N_20411,N_16236,N_18252);
and U20412 (N_20412,N_17677,N_16830);
nor U20413 (N_20413,N_15031,N_16940);
nand U20414 (N_20414,N_18901,N_17010);
or U20415 (N_20415,N_17867,N_15944);
or U20416 (N_20416,N_15552,N_18169);
xor U20417 (N_20417,N_18062,N_15982);
nor U20418 (N_20418,N_15608,N_19453);
nand U20419 (N_20419,N_16935,N_18023);
or U20420 (N_20420,N_19011,N_16983);
and U20421 (N_20421,N_17975,N_19562);
xor U20422 (N_20422,N_16925,N_17829);
xnor U20423 (N_20423,N_15962,N_17293);
and U20424 (N_20424,N_15360,N_19014);
nand U20425 (N_20425,N_18823,N_16507);
and U20426 (N_20426,N_18797,N_19681);
nor U20427 (N_20427,N_17985,N_18464);
nor U20428 (N_20428,N_19747,N_16233);
and U20429 (N_20429,N_17600,N_19815);
and U20430 (N_20430,N_16960,N_17152);
nor U20431 (N_20431,N_17286,N_18126);
or U20432 (N_20432,N_18643,N_16244);
nand U20433 (N_20433,N_19141,N_19965);
nor U20434 (N_20434,N_16462,N_19121);
nor U20435 (N_20435,N_15939,N_18771);
and U20436 (N_20436,N_19909,N_19534);
and U20437 (N_20437,N_19526,N_17081);
or U20438 (N_20438,N_17679,N_18616);
or U20439 (N_20439,N_15121,N_17724);
nand U20440 (N_20440,N_17377,N_19338);
or U20441 (N_20441,N_17494,N_19811);
or U20442 (N_20442,N_18992,N_19976);
nand U20443 (N_20443,N_17182,N_15672);
and U20444 (N_20444,N_16515,N_19109);
and U20445 (N_20445,N_15395,N_19318);
and U20446 (N_20446,N_17355,N_16300);
xnor U20447 (N_20447,N_15554,N_17750);
or U20448 (N_20448,N_18465,N_18480);
nor U20449 (N_20449,N_15178,N_18867);
nor U20450 (N_20450,N_17759,N_16404);
nor U20451 (N_20451,N_18852,N_15914);
nand U20452 (N_20452,N_18666,N_19024);
or U20453 (N_20453,N_17289,N_16448);
xor U20454 (N_20454,N_16337,N_15585);
and U20455 (N_20455,N_15263,N_19715);
nand U20456 (N_20456,N_15247,N_17964);
and U20457 (N_20457,N_16428,N_19441);
nand U20458 (N_20458,N_15434,N_15460);
nor U20459 (N_20459,N_15758,N_18399);
xor U20460 (N_20460,N_15855,N_15615);
nor U20461 (N_20461,N_19200,N_18123);
nor U20462 (N_20462,N_15427,N_18238);
nor U20463 (N_20463,N_19330,N_16264);
or U20464 (N_20464,N_15432,N_15872);
and U20465 (N_20465,N_17084,N_19490);
nor U20466 (N_20466,N_18753,N_19805);
nor U20467 (N_20467,N_15130,N_17371);
xor U20468 (N_20468,N_18532,N_19553);
or U20469 (N_20469,N_19549,N_17632);
xnor U20470 (N_20470,N_19465,N_17012);
or U20471 (N_20471,N_17240,N_18158);
xor U20472 (N_20472,N_15021,N_16716);
nand U20473 (N_20473,N_19249,N_17418);
and U20474 (N_20474,N_19208,N_15437);
or U20475 (N_20475,N_19344,N_15625);
nor U20476 (N_20476,N_19506,N_17997);
nor U20477 (N_20477,N_15414,N_18397);
and U20478 (N_20478,N_15937,N_15077);
and U20479 (N_20479,N_17342,N_18968);
nor U20480 (N_20480,N_17639,N_16294);
and U20481 (N_20481,N_17111,N_15638);
nand U20482 (N_20482,N_19437,N_18727);
or U20483 (N_20483,N_19345,N_17949);
nor U20484 (N_20484,N_15323,N_18530);
or U20485 (N_20485,N_17756,N_15089);
and U20486 (N_20486,N_16627,N_19744);
and U20487 (N_20487,N_17420,N_15097);
nand U20488 (N_20488,N_17645,N_19987);
xor U20489 (N_20489,N_17941,N_17840);
and U20490 (N_20490,N_16734,N_16914);
nor U20491 (N_20491,N_18376,N_16570);
and U20492 (N_20492,N_18799,N_16351);
nand U20493 (N_20493,N_16631,N_19091);
and U20494 (N_20494,N_18412,N_19214);
nand U20495 (N_20495,N_16140,N_18377);
nand U20496 (N_20496,N_16963,N_15597);
or U20497 (N_20497,N_15858,N_18227);
or U20498 (N_20498,N_16335,N_16031);
nor U20499 (N_20499,N_19233,N_17320);
nor U20500 (N_20500,N_17250,N_17628);
and U20501 (N_20501,N_16464,N_16343);
nand U20502 (N_20502,N_15157,N_16112);
nand U20503 (N_20503,N_16133,N_18579);
and U20504 (N_20504,N_18831,N_15790);
nor U20505 (N_20505,N_16362,N_18605);
nand U20506 (N_20506,N_19089,N_16450);
nand U20507 (N_20507,N_18576,N_17329);
or U20508 (N_20508,N_18814,N_16479);
nand U20509 (N_20509,N_18423,N_15652);
or U20510 (N_20510,N_18498,N_17697);
xor U20511 (N_20511,N_17497,N_18315);
nand U20512 (N_20512,N_17656,N_18627);
nand U20513 (N_20513,N_15192,N_18894);
and U20514 (N_20514,N_18816,N_17691);
nand U20515 (N_20515,N_17843,N_16730);
or U20516 (N_20516,N_16718,N_15885);
nor U20517 (N_20517,N_17341,N_18842);
or U20518 (N_20518,N_19901,N_16444);
nor U20519 (N_20519,N_15582,N_19020);
nor U20520 (N_20520,N_16770,N_19044);
xor U20521 (N_20521,N_16091,N_19580);
and U20522 (N_20522,N_18210,N_18246);
nand U20523 (N_20523,N_16736,N_16690);
nor U20524 (N_20524,N_15831,N_19640);
or U20525 (N_20525,N_18417,N_17787);
or U20526 (N_20526,N_18219,N_16340);
xor U20527 (N_20527,N_15863,N_19097);
and U20528 (N_20528,N_19759,N_17877);
nand U20529 (N_20529,N_17343,N_18840);
and U20530 (N_20530,N_16106,N_18054);
nand U20531 (N_20531,N_18046,N_16916);
nand U20532 (N_20532,N_18163,N_19707);
xor U20533 (N_20533,N_18116,N_15591);
nand U20534 (N_20534,N_15005,N_15648);
and U20535 (N_20535,N_18745,N_17704);
xnor U20536 (N_20536,N_15596,N_16424);
nor U20537 (N_20537,N_17821,N_15667);
nand U20538 (N_20538,N_17983,N_18548);
nand U20539 (N_20539,N_17470,N_18767);
xnor U20540 (N_20540,N_16619,N_19115);
nor U20541 (N_20541,N_15079,N_18040);
nand U20542 (N_20542,N_16595,N_18989);
nor U20543 (N_20543,N_16327,N_15592);
nor U20544 (N_20544,N_15802,N_19604);
and U20545 (N_20545,N_18587,N_15499);
and U20546 (N_20546,N_18322,N_17991);
and U20547 (N_20547,N_16816,N_18176);
nand U20548 (N_20548,N_16646,N_17370);
and U20549 (N_20549,N_16614,N_19579);
xnor U20550 (N_20550,N_19324,N_16817);
or U20551 (N_20551,N_16182,N_17168);
nand U20552 (N_20552,N_15102,N_18984);
xor U20553 (N_20553,N_16997,N_18331);
nand U20554 (N_20554,N_15352,N_15366);
nand U20555 (N_20555,N_15857,N_18564);
nand U20556 (N_20556,N_16503,N_18404);
nor U20557 (N_20557,N_17661,N_18504);
or U20558 (N_20558,N_15008,N_19126);
nand U20559 (N_20559,N_19786,N_15010);
nand U20560 (N_20560,N_17197,N_17203);
and U20561 (N_20561,N_16807,N_17086);
nand U20562 (N_20562,N_17979,N_18474);
or U20563 (N_20563,N_18768,N_15675);
nor U20564 (N_20564,N_17499,N_18729);
nor U20565 (N_20565,N_19521,N_16352);
nor U20566 (N_20566,N_15304,N_15926);
nand U20567 (N_20567,N_17067,N_17104);
nor U20568 (N_20568,N_15016,N_17732);
nand U20569 (N_20569,N_18466,N_17139);
nor U20570 (N_20570,N_16580,N_18923);
nand U20571 (N_20571,N_19087,N_18390);
and U20572 (N_20572,N_16818,N_19085);
and U20573 (N_20573,N_16951,N_18638);
or U20574 (N_20574,N_15249,N_15109);
and U20575 (N_20575,N_15264,N_19630);
and U20576 (N_20576,N_16087,N_15958);
or U20577 (N_20577,N_17219,N_17301);
nand U20578 (N_20578,N_18567,N_19864);
nand U20579 (N_20579,N_17834,N_16321);
and U20580 (N_20580,N_19315,N_16252);
and U20581 (N_20581,N_17447,N_19569);
nand U20582 (N_20582,N_16589,N_17536);
nor U20583 (N_20583,N_15391,N_19958);
or U20584 (N_20584,N_18810,N_19997);
nor U20585 (N_20585,N_17771,N_18637);
and U20586 (N_20586,N_15448,N_15339);
nand U20587 (N_20587,N_16545,N_17664);
nand U20588 (N_20588,N_16649,N_15827);
or U20589 (N_20589,N_18305,N_17070);
nor U20590 (N_20590,N_18895,N_16219);
nor U20591 (N_20591,N_18332,N_16414);
nor U20592 (N_20592,N_16441,N_16869);
nor U20593 (N_20593,N_17060,N_15138);
xor U20594 (N_20594,N_15177,N_19102);
nand U20595 (N_20595,N_16927,N_17025);
and U20596 (N_20596,N_19250,N_17144);
xnor U20597 (N_20597,N_16355,N_19984);
nand U20598 (N_20598,N_19263,N_18518);
or U20599 (N_20599,N_16967,N_17068);
nand U20600 (N_20600,N_17465,N_19727);
and U20601 (N_20601,N_15963,N_19830);
or U20602 (N_20602,N_19276,N_15415);
xnor U20603 (N_20603,N_19341,N_16976);
and U20604 (N_20604,N_18462,N_19972);
and U20605 (N_20605,N_16650,N_16029);
nand U20606 (N_20606,N_16242,N_17772);
and U20607 (N_20607,N_17080,N_18027);
or U20608 (N_20608,N_17706,N_16286);
nor U20609 (N_20609,N_19698,N_15509);
nor U20610 (N_20610,N_17406,N_16933);
xor U20611 (N_20611,N_19746,N_19508);
or U20612 (N_20612,N_15573,N_16373);
and U20613 (N_20613,N_18529,N_16379);
xnor U20614 (N_20614,N_18429,N_18507);
or U20615 (N_20615,N_17825,N_15306);
nor U20616 (N_20616,N_15214,N_16457);
and U20617 (N_20617,N_16600,N_15250);
nand U20618 (N_20618,N_18619,N_17457);
and U20619 (N_20619,N_17196,N_15711);
or U20620 (N_20620,N_15930,N_17307);
nand U20621 (N_20621,N_16023,N_17252);
or U20622 (N_20622,N_17762,N_18793);
nand U20623 (N_20623,N_19722,N_16524);
or U20624 (N_20624,N_16131,N_17427);
nand U20625 (N_20625,N_18096,N_16952);
nor U20626 (N_20626,N_18005,N_15907);
nor U20627 (N_20627,N_19261,N_18848);
and U20628 (N_20628,N_19252,N_18779);
nor U20629 (N_20629,N_15255,N_15968);
and U20630 (N_20630,N_18892,N_17540);
nand U20631 (N_20631,N_19361,N_15032);
nand U20632 (N_20632,N_17288,N_15222);
or U20633 (N_20633,N_18107,N_17907);
or U20634 (N_20634,N_19868,N_19277);
nor U20635 (N_20635,N_16454,N_17815);
nor U20636 (N_20636,N_19094,N_18545);
or U20637 (N_20637,N_16304,N_18172);
or U20638 (N_20638,N_19448,N_15083);
xnor U20639 (N_20639,N_16813,N_18414);
nor U20640 (N_20640,N_19912,N_19414);
nor U20641 (N_20641,N_18738,N_17248);
nand U20642 (N_20642,N_19801,N_16805);
nor U20643 (N_20643,N_16773,N_16228);
and U20644 (N_20644,N_17262,N_15218);
or U20645 (N_20645,N_19107,N_18834);
or U20646 (N_20646,N_18357,N_15134);
or U20647 (N_20647,N_19348,N_19852);
nor U20648 (N_20648,N_16092,N_15817);
or U20649 (N_20649,N_18066,N_18593);
nand U20650 (N_20650,N_18457,N_19639);
nand U20651 (N_20651,N_18232,N_16659);
xnor U20652 (N_20652,N_18029,N_18864);
nand U20653 (N_20653,N_18401,N_15556);
nand U20654 (N_20654,N_16547,N_18990);
and U20655 (N_20655,N_16180,N_16761);
xor U20656 (N_20656,N_17202,N_17641);
or U20657 (N_20657,N_18599,N_19283);
nor U20658 (N_20658,N_19426,N_15523);
nand U20659 (N_20659,N_16564,N_19803);
and U20660 (N_20660,N_17715,N_15262);
nand U20661 (N_20661,N_15299,N_18247);
nand U20662 (N_20662,N_16386,N_19831);
nor U20663 (N_20663,N_18300,N_18168);
and U20664 (N_20664,N_16203,N_17445);
and U20665 (N_20665,N_19375,N_16656);
and U20666 (N_20666,N_16249,N_19750);
xor U20667 (N_20667,N_17065,N_17348);
nand U20668 (N_20668,N_19779,N_15589);
nor U20669 (N_20669,N_16128,N_16563);
and U20670 (N_20670,N_17610,N_16705);
or U20671 (N_20671,N_19879,N_17802);
nand U20672 (N_20672,N_18198,N_18817);
or U20673 (N_20673,N_17407,N_15101);
nand U20674 (N_20674,N_17751,N_18628);
nor U20675 (N_20675,N_19797,N_19157);
nand U20676 (N_20676,N_17369,N_18000);
nor U20677 (N_20677,N_16655,N_15453);
and U20678 (N_20678,N_16523,N_19923);
nand U20679 (N_20679,N_18053,N_15137);
or U20680 (N_20680,N_18623,N_16715);
and U20681 (N_20681,N_16620,N_17506);
nand U20682 (N_20682,N_15613,N_17806);
or U20683 (N_20683,N_16197,N_17728);
nor U20684 (N_20684,N_17720,N_19757);
nand U20685 (N_20685,N_18085,N_15348);
and U20686 (N_20686,N_15565,N_18565);
nor U20687 (N_20687,N_17748,N_19207);
nand U20688 (N_20688,N_15969,N_15392);
and U20689 (N_20689,N_19777,N_15045);
nor U20690 (N_20690,N_15940,N_18869);
or U20691 (N_20691,N_18119,N_17331);
nand U20692 (N_20692,N_16036,N_16306);
or U20693 (N_20693,N_15239,N_16485);
or U20694 (N_20694,N_18752,N_19637);
or U20695 (N_20695,N_15261,N_18868);
and U20696 (N_20696,N_15859,N_19880);
or U20697 (N_20697,N_18577,N_16012);
nor U20698 (N_20698,N_15800,N_18344);
or U20699 (N_20699,N_19826,N_18133);
or U20700 (N_20700,N_18671,N_17359);
nor U20701 (N_20701,N_16514,N_19396);
or U20702 (N_20702,N_15235,N_18535);
nand U20703 (N_20703,N_15358,N_17729);
or U20704 (N_20704,N_18680,N_18597);
or U20705 (N_20705,N_19738,N_19319);
and U20706 (N_20706,N_16442,N_16865);
or U20707 (N_20707,N_16433,N_16628);
xor U20708 (N_20708,N_15412,N_19851);
or U20709 (N_20709,N_15881,N_17962);
or U20710 (N_20710,N_18179,N_16746);
or U20711 (N_20711,N_18855,N_16061);
or U20712 (N_20712,N_15695,N_18673);
nor U20713 (N_20713,N_17934,N_17957);
nor U20714 (N_20714,N_15878,N_19587);
nor U20715 (N_20715,N_18380,N_18785);
nand U20716 (N_20716,N_17428,N_15612);
or U20717 (N_20717,N_19230,N_19100);
nor U20718 (N_20718,N_17942,N_18603);
xnor U20719 (N_20719,N_16875,N_18257);
and U20720 (N_20720,N_19491,N_15950);
nor U20721 (N_20721,N_19481,N_19775);
nand U20722 (N_20722,N_16593,N_15583);
and U20723 (N_20723,N_18415,N_17705);
nor U20724 (N_20724,N_19494,N_18241);
and U20725 (N_20725,N_16405,N_15576);
xor U20726 (N_20726,N_17169,N_17032);
nand U20727 (N_20727,N_17837,N_19856);
nand U20728 (N_20728,N_19905,N_16522);
nand U20729 (N_20729,N_16437,N_18453);
nor U20730 (N_20730,N_15301,N_19778);
or U20731 (N_20731,N_15080,N_15140);
nand U20732 (N_20732,N_18938,N_17513);
and U20733 (N_20733,N_17183,N_15883);
and U20734 (N_20734,N_17234,N_19380);
or U20735 (N_20735,N_15098,N_18181);
nand U20736 (N_20736,N_16618,N_15816);
or U20737 (N_20737,N_15151,N_19035);
or U20738 (N_20738,N_19828,N_18635);
nand U20739 (N_20739,N_15633,N_16926);
or U20740 (N_20740,N_16911,N_15796);
xor U20741 (N_20741,N_18078,N_15380);
and U20742 (N_20742,N_18506,N_17063);
nor U20743 (N_20743,N_15204,N_18939);
xor U20744 (N_20744,N_16964,N_17229);
or U20745 (N_20745,N_15840,N_15413);
and U20746 (N_20746,N_15527,N_15741);
or U20747 (N_20747,N_19950,N_18445);
nor U20748 (N_20748,N_17963,N_16299);
or U20749 (N_20749,N_15704,N_16151);
xor U20750 (N_20750,N_16738,N_18857);
and U20751 (N_20751,N_16003,N_18148);
nor U20752 (N_20752,N_19765,N_19082);
and U20753 (N_20753,N_19966,N_17487);
and U20754 (N_20754,N_19899,N_15309);
xnor U20755 (N_20755,N_17227,N_16686);
and U20756 (N_20756,N_19194,N_17372);
or U20757 (N_20757,N_17546,N_15620);
or U20758 (N_20758,N_17046,N_16483);
nor U20759 (N_20759,N_15994,N_15760);
nor U20760 (N_20760,N_17368,N_19395);
nand U20761 (N_20761,N_16676,N_19529);
or U20762 (N_20762,N_19374,N_16171);
and U20763 (N_20763,N_18461,N_15546);
xnor U20764 (N_20764,N_15588,N_18909);
nand U20765 (N_20765,N_19664,N_18146);
or U20766 (N_20766,N_19446,N_19942);
and U20767 (N_20767,N_15543,N_19080);
and U20768 (N_20768,N_15657,N_19558);
nand U20769 (N_20769,N_17927,N_17919);
nand U20770 (N_20770,N_16920,N_16216);
and U20771 (N_20771,N_17074,N_16836);
nand U20772 (N_20772,N_16482,N_19933);
or U20773 (N_20773,N_17270,N_17094);
nor U20774 (N_20774,N_15012,N_15248);
nor U20775 (N_20775,N_15929,N_16050);
and U20776 (N_20776,N_19999,N_18349);
or U20777 (N_20777,N_16116,N_17176);
or U20778 (N_20778,N_18812,N_19885);
and U20779 (N_20779,N_19211,N_16546);
nand U20780 (N_20780,N_19180,N_19724);
or U20781 (N_20781,N_19867,N_17142);
nor U20782 (N_20782,N_15844,N_15075);
nor U20783 (N_20783,N_15442,N_18584);
nor U20784 (N_20784,N_18114,N_16028);
or U20785 (N_20785,N_18761,N_19168);
nor U20786 (N_20786,N_15528,N_19444);
or U20787 (N_20787,N_18970,N_18002);
xnor U20788 (N_20788,N_17881,N_17255);
and U20789 (N_20789,N_18790,N_15317);
nor U20790 (N_20790,N_15983,N_16666);
and U20791 (N_20791,N_19537,N_17020);
and U20792 (N_20792,N_18523,N_17668);
or U20793 (N_20793,N_19908,N_15288);
nor U20794 (N_20794,N_15751,N_17966);
nand U20795 (N_20795,N_17514,N_17335);
nand U20796 (N_20796,N_16704,N_19612);
nand U20797 (N_20797,N_15974,N_15809);
nor U20798 (N_20798,N_18604,N_19581);
and U20799 (N_20799,N_16193,N_17218);
and U20800 (N_20800,N_15326,N_19689);
nand U20801 (N_20801,N_17879,N_19733);
xnor U20802 (N_20802,N_19317,N_15076);
or U20803 (N_20803,N_19321,N_18032);
nor U20804 (N_20804,N_18326,N_19075);
or U20805 (N_20805,N_19349,N_15684);
nand U20806 (N_20806,N_18491,N_17044);
nor U20807 (N_20807,N_16673,N_18249);
or U20808 (N_20808,N_16852,N_17816);
and U20809 (N_20809,N_16699,N_18183);
xor U20810 (N_20810,N_15644,N_18811);
nand U20811 (N_20811,N_19613,N_18076);
or U20812 (N_20812,N_15765,N_16877);
nor U20813 (N_20813,N_18162,N_15533);
or U20814 (N_20814,N_15009,N_17108);
nand U20815 (N_20815,N_17993,N_17922);
or U20816 (N_20816,N_16267,N_19019);
xor U20817 (N_20817,N_15833,N_18601);
and U20818 (N_20818,N_17814,N_19583);
nand U20819 (N_20819,N_18493,N_19763);
nor U20820 (N_20820,N_15293,N_19028);
nand U20821 (N_20821,N_17266,N_16722);
and U20822 (N_20822,N_18681,N_18413);
and U20823 (N_20823,N_16030,N_15443);
nor U20824 (N_20824,N_18063,N_15397);
nor U20825 (N_20825,N_18077,N_17794);
and U20826 (N_20826,N_16259,N_18041);
xnor U20827 (N_20827,N_15787,N_15244);
xor U20828 (N_20828,N_18224,N_18382);
nor U20829 (N_20829,N_15964,N_16315);
nor U20830 (N_20830,N_15654,N_15560);
xnor U20831 (N_20831,N_15478,N_16156);
nor U20832 (N_20832,N_15356,N_15774);
nor U20833 (N_20833,N_17667,N_17666);
xnor U20834 (N_20834,N_17689,N_19438);
nand U20835 (N_20835,N_18242,N_19308);
and U20836 (N_20836,N_17217,N_17458);
and U20837 (N_20837,N_16336,N_18856);
nor U20838 (N_20838,N_17468,N_17344);
or U20839 (N_20839,N_19670,N_19531);
and U20840 (N_20840,N_18988,N_19782);
and U20841 (N_20841,N_16471,N_19234);
and U20842 (N_20842,N_17582,N_17797);
nor U20843 (N_20843,N_19626,N_17624);
nor U20844 (N_20844,N_19181,N_17805);
nand U20845 (N_20845,N_17422,N_18265);
nand U20846 (N_20846,N_17518,N_16372);
or U20847 (N_20847,N_18403,N_15709);
nand U20848 (N_20848,N_16377,N_19034);
and U20849 (N_20849,N_15373,N_18388);
and U20850 (N_20850,N_15308,N_18031);
xor U20851 (N_20851,N_17446,N_19193);
or U20852 (N_20852,N_18913,N_17852);
nand U20853 (N_20853,N_18749,N_16831);
or U20854 (N_20854,N_16941,N_16453);
and U20855 (N_20855,N_15674,N_19875);
xor U20856 (N_20856,N_15065,N_18526);
or U20857 (N_20857,N_18586,N_19938);
nand U20858 (N_20858,N_17394,N_15575);
or U20859 (N_20859,N_17875,N_19172);
nand U20860 (N_20860,N_18866,N_17651);
or U20861 (N_20861,N_15776,N_16278);
nor U20862 (N_20862,N_15946,N_19320);
nand U20863 (N_20863,N_16396,N_17466);
nand U20864 (N_20864,N_16000,N_17865);
and U20865 (N_20865,N_16010,N_16525);
or U20866 (N_20866,N_19146,N_18854);
nand U20867 (N_20867,N_19381,N_19247);
or U20868 (N_20868,N_19251,N_16395);
nand U20869 (N_20869,N_17193,N_18755);
or U20870 (N_20870,N_19162,N_19947);
nand U20871 (N_20871,N_16445,N_19892);
nand U20872 (N_20872,N_15421,N_19058);
nor U20873 (N_20873,N_17574,N_18188);
nand U20874 (N_20874,N_19517,N_18289);
and U20875 (N_20875,N_16217,N_17788);
or U20876 (N_20876,N_17120,N_18975);
nand U20877 (N_20877,N_18379,N_17432);
nand U20878 (N_20878,N_18503,N_19977);
nor U20879 (N_20879,N_19388,N_18092);
and U20880 (N_20880,N_17130,N_16645);
or U20881 (N_20881,N_17132,N_19751);
nor U20882 (N_20882,N_16310,N_16748);
nor U20883 (N_20883,N_16901,N_19031);
and U20884 (N_20884,N_18731,N_16266);
and U20885 (N_20885,N_16484,N_17122);
and U20886 (N_20886,N_19489,N_18292);
nand U20887 (N_20887,N_15676,N_19067);
xor U20888 (N_20888,N_16743,N_17314);
nor U20889 (N_20889,N_15334,N_19788);
or U20890 (N_20890,N_15445,N_17909);
nor U20891 (N_20891,N_17354,N_18614);
or U20892 (N_20892,N_18434,N_19149);
nand U20893 (N_20893,N_19061,N_16208);
and U20894 (N_20894,N_15447,N_17431);
nor U20895 (N_20895,N_15074,N_18728);
nand U20896 (N_20896,N_19718,N_16853);
or U20897 (N_20897,N_16276,N_15426);
nand U20898 (N_20898,N_17567,N_17606);
nand U20899 (N_20899,N_18710,N_15361);
or U20900 (N_20900,N_19416,N_15367);
or U20901 (N_20901,N_18511,N_18364);
or U20902 (N_20902,N_15763,N_19217);
xor U20903 (N_20903,N_15567,N_19974);
nor U20904 (N_20904,N_15880,N_15896);
nand U20905 (N_20905,N_18688,N_18047);
nor U20906 (N_20906,N_19117,N_16697);
and U20907 (N_20907,N_19158,N_17817);
nor U20908 (N_20908,N_17897,N_15874);
nand U20909 (N_20909,N_15734,N_17832);
and U20910 (N_20910,N_16623,N_18508);
nor U20911 (N_20911,N_15604,N_18964);
or U20912 (N_20912,N_17680,N_19663);
xnor U20913 (N_20913,N_18541,N_15520);
xor U20914 (N_20914,N_16737,N_15731);
nor U20915 (N_20915,N_18011,N_18234);
nor U20916 (N_20916,N_15211,N_15069);
and U20917 (N_20917,N_19084,N_17035);
nor U20918 (N_20918,N_18633,N_19712);
and U20919 (N_20919,N_16605,N_19443);
or U20920 (N_20920,N_16493,N_17987);
and U20921 (N_20921,N_16161,N_15889);
or U20922 (N_20922,N_18758,N_19672);
nand U20923 (N_20923,N_18685,N_15345);
nor U20924 (N_20924,N_16094,N_15125);
and U20925 (N_20925,N_15913,N_15093);
and U20926 (N_20926,N_19762,N_15618);
nand U20927 (N_20927,N_18202,N_16557);
or U20928 (N_20928,N_16037,N_16792);
xnor U20929 (N_20929,N_16052,N_18304);
nand U20930 (N_20930,N_19316,N_19471);
and U20931 (N_20931,N_17940,N_16809);
and U20932 (N_20932,N_18715,N_16068);
xor U20933 (N_20933,N_18073,N_17831);
nand U20934 (N_20934,N_18687,N_19507);
nor U20935 (N_20935,N_19064,N_17382);
nor U20936 (N_20936,N_15882,N_15918);
and U20937 (N_20937,N_18496,N_18048);
xor U20938 (N_20938,N_15205,N_19222);
or U20939 (N_20939,N_15551,N_15189);
nand U20940 (N_20940,N_17226,N_16124);
and U20941 (N_20941,N_19781,N_19850);
nand U20942 (N_20942,N_17029,N_17900);
or U20943 (N_20943,N_17340,N_15524);
xor U20944 (N_20944,N_18900,N_19732);
nand U20945 (N_20945,N_16088,N_18372);
xor U20946 (N_20946,N_17930,N_19173);
or U20947 (N_20947,N_15538,N_16821);
nand U20948 (N_20948,N_18819,N_19895);
nand U20949 (N_20949,N_17257,N_16192);
or U20950 (N_20950,N_18736,N_16381);
and U20951 (N_20951,N_15278,N_18784);
or U20952 (N_20952,N_16008,N_17017);
and U20953 (N_20953,N_17896,N_19502);
and U20954 (N_20954,N_18036,N_15553);
nor U20955 (N_20955,N_18946,N_17891);
nor U20956 (N_20956,N_17714,N_16406);
nor U20957 (N_20957,N_17502,N_15661);
and U20958 (N_20958,N_18641,N_15681);
nand U20959 (N_20959,N_18582,N_16126);
nand U20960 (N_20960,N_15394,N_18237);
and U20961 (N_20961,N_19910,N_15479);
or U20962 (N_20962,N_15603,N_19147);
nor U20963 (N_20963,N_16376,N_15467);
and U20964 (N_20964,N_16811,N_19333);
xnor U20965 (N_20965,N_17360,N_18860);
nand U20966 (N_20966,N_19567,N_16458);
nor U20967 (N_20967,N_18515,N_16184);
nand U20968 (N_20968,N_15173,N_19948);
and U20969 (N_20969,N_16042,N_15867);
and U20970 (N_20970,N_15852,N_16475);
or U20971 (N_20971,N_17441,N_17857);
nand U20972 (N_20972,N_19287,N_16662);
or U20973 (N_20973,N_16767,N_15512);
nor U20974 (N_20974,N_17478,N_18254);
nand U20975 (N_20975,N_19896,N_15721);
and U20976 (N_20976,N_18284,N_16825);
and U20977 (N_20977,N_16231,N_15476);
nor U20978 (N_20978,N_18293,N_15679);
and U20979 (N_20979,N_18916,N_15408);
nand U20980 (N_20980,N_17819,N_16263);
xnor U20981 (N_20981,N_16913,N_15617);
and U20982 (N_20982,N_18561,N_17284);
nor U20983 (N_20983,N_18951,N_17244);
nand U20984 (N_20984,N_16682,N_18100);
and U20985 (N_20985,N_16210,N_19459);
nand U20986 (N_20986,N_16957,N_19836);
nand U20987 (N_20987,N_18721,N_19684);
and U20988 (N_20988,N_15899,N_16928);
nand U20989 (N_20989,N_16333,N_15662);
and U20990 (N_20990,N_17512,N_18149);
or U20991 (N_20991,N_15772,N_15798);
xnor U20992 (N_20992,N_18850,N_16297);
nor U20993 (N_20993,N_15826,N_17901);
nand U20994 (N_20994,N_15199,N_19969);
and U20995 (N_20995,N_16641,N_18127);
and U20996 (N_20996,N_18664,N_18692);
xor U20997 (N_20997,N_18932,N_15562);
and U20998 (N_20998,N_17039,N_17872);
nor U20999 (N_20999,N_18393,N_18872);
and U21000 (N_21000,N_15152,N_16774);
nor U21001 (N_21001,N_18356,N_18385);
and U21002 (N_21002,N_17893,N_15451);
and U21003 (N_21003,N_18961,N_19990);
and U21004 (N_21004,N_15430,N_19254);
nand U21005 (N_21005,N_16910,N_19855);
nor U21006 (N_21006,N_16790,N_17337);
nand U21007 (N_21007,N_18954,N_17933);
or U21008 (N_21008,N_17099,N_19996);
nor U21009 (N_21009,N_15349,N_15034);
nand U21010 (N_21010,N_18173,N_16874);
nand U21011 (N_21011,N_17501,N_16134);
or U21012 (N_21012,N_19485,N_16949);
xnor U21013 (N_21013,N_19832,N_19464);
and U21014 (N_21014,N_17701,N_15737);
nor U21015 (N_21015,N_19800,N_16345);
nor U21016 (N_21016,N_18520,N_19405);
and U21017 (N_21017,N_15095,N_18544);
or U21018 (N_21018,N_17575,N_18267);
and U21019 (N_21019,N_18004,N_18028);
and U21020 (N_21020,N_17275,N_15381);
nand U21021 (N_21021,N_19136,N_18977);
or U21022 (N_21022,N_15864,N_15514);
and U21023 (N_21023,N_19932,N_19866);
nor U21024 (N_21024,N_19391,N_16271);
and U21025 (N_21025,N_15025,N_18748);
or U21026 (N_21026,N_18667,N_16086);
nor U21027 (N_21027,N_18064,N_17188);
nor U21028 (N_21028,N_19847,N_16226);
and U21029 (N_21029,N_18487,N_19578);
xor U21030 (N_21030,N_19177,N_18948);
nand U21031 (N_21031,N_15338,N_15606);
or U21032 (N_21032,N_15048,N_18479);
and U21033 (N_21033,N_17708,N_15917);
nand U21034 (N_21034,N_17013,N_18141);
or U21035 (N_21035,N_18676,N_19373);
or U21036 (N_21036,N_15329,N_16186);
or U21037 (N_21037,N_19891,N_15702);
or U21038 (N_21038,N_19236,N_19195);
nor U21039 (N_21039,N_18306,N_16749);
xor U21040 (N_21040,N_15082,N_15053);
nand U21041 (N_21041,N_15002,N_18239);
and U21042 (N_21042,N_17516,N_17908);
xnor U21043 (N_21043,N_19343,N_18180);
nand U21044 (N_21044,N_16829,N_17520);
or U21045 (N_21045,N_18341,N_15228);
and U21046 (N_21046,N_15823,N_19394);
or U21047 (N_21047,N_17528,N_18335);
nand U21048 (N_21048,N_16302,N_16728);
and U21049 (N_21049,N_17109,N_19422);
and U21050 (N_21050,N_19857,N_15014);
or U21051 (N_21051,N_19268,N_18375);
xor U21052 (N_21052,N_16590,N_18849);
or U21053 (N_21053,N_17435,N_15860);
and U21054 (N_21054,N_15578,N_17584);
nor U21055 (N_21055,N_18960,N_15838);
or U21056 (N_21056,N_16218,N_19497);
nor U21057 (N_21057,N_19584,N_18533);
and U21058 (N_21058,N_15935,N_17300);
nand U21059 (N_21059,N_19119,N_19675);
xor U21060 (N_21060,N_18875,N_18328);
and U21061 (N_21061,N_18340,N_16881);
nor U21062 (N_21062,N_17703,N_16789);
and U21063 (N_21063,N_17271,N_17224);
and U21064 (N_21064,N_18451,N_16248);
or U21065 (N_21065,N_17537,N_16265);
or U21066 (N_21066,N_17836,N_18440);
or U21067 (N_21067,N_19182,N_17874);
or U21068 (N_21068,N_19980,N_16810);
nand U21069 (N_21069,N_15791,N_19400);
nor U21070 (N_21070,N_15344,N_16799);
or U21071 (N_21071,N_17761,N_17114);
nor U21072 (N_21072,N_19133,N_17069);
or U21073 (N_21073,N_19334,N_15886);
nand U21074 (N_21074,N_18510,N_16407);
and U21075 (N_21075,N_15209,N_18712);
nand U21076 (N_21076,N_17583,N_16984);
nand U21077 (N_21077,N_17774,N_16652);
or U21078 (N_21078,N_18657,N_16429);
nand U21079 (N_21079,N_16332,N_18959);
nor U21080 (N_21080,N_19957,N_19554);
or U21081 (N_21081,N_18747,N_18701);
or U21082 (N_21082,N_19423,N_19823);
and U21083 (N_21083,N_17736,N_16549);
nand U21084 (N_21084,N_16977,N_17599);
nand U21085 (N_21085,N_17030,N_19387);
and U21086 (N_21086,N_15406,N_18314);
and U21087 (N_21087,N_19226,N_15231);
and U21088 (N_21088,N_18547,N_17681);
nand U21089 (N_21089,N_16832,N_15853);
and U21090 (N_21090,N_16213,N_18233);
nor U21091 (N_21091,N_16047,N_15989);
and U21092 (N_21092,N_15232,N_18367);
xnor U21093 (N_21093,N_17064,N_19853);
nor U21094 (N_21094,N_19392,N_15399);
or U21095 (N_21095,N_18277,N_17469);
and U21096 (N_21096,N_19952,N_17129);
nor U21097 (N_21097,N_16191,N_17538);
nor U21098 (N_21098,N_17937,N_16884);
and U21099 (N_21099,N_15119,N_15029);
or U21100 (N_21100,N_18370,N_19487);
and U21101 (N_21101,N_16536,N_15281);
nand U21102 (N_21102,N_17894,N_19466);
nor U21103 (N_21103,N_19555,N_19649);
nand U21104 (N_21104,N_19694,N_19351);
or U21105 (N_21105,N_19043,N_16393);
nor U21106 (N_21106,N_15229,N_17921);
xor U21107 (N_21107,N_19242,N_18630);
nor U21108 (N_21108,N_18528,N_19191);
or U21109 (N_21109,N_17392,N_15275);
nand U21110 (N_21110,N_16848,N_17200);
and U21111 (N_21111,N_18051,N_17186);
nand U21112 (N_21112,N_18502,N_16696);
or U21113 (N_21113,N_19964,N_17281);
nor U21114 (N_21114,N_19883,N_15042);
and U21115 (N_21115,N_16488,N_17725);
xor U21116 (N_21116,N_19524,N_18613);
and U21117 (N_21117,N_16041,N_16409);
or U21118 (N_21118,N_15540,N_18670);
nand U21119 (N_21119,N_17539,N_17970);
or U21120 (N_21120,N_19888,N_16438);
nand U21121 (N_21121,N_16707,N_17792);
or U21122 (N_21122,N_16965,N_15279);
or U21123 (N_21123,N_15832,N_15978);
nor U21124 (N_21124,N_17353,N_18447);
nor U21125 (N_21125,N_19799,N_19295);
nand U21126 (N_21126,N_15411,N_19900);
nand U21127 (N_21127,N_15212,N_15683);
and U21128 (N_21128,N_18965,N_15593);
or U21129 (N_21129,N_19367,N_15267);
and U21130 (N_21130,N_18161,N_16392);
nor U21131 (N_21131,N_19846,N_19914);
nand U21132 (N_21132,N_16019,N_16808);
xor U21133 (N_21133,N_15354,N_19668);
or U21134 (N_21134,N_15060,N_18781);
nor U21135 (N_21135,N_16253,N_16097);
nand U21136 (N_21136,N_16055,N_19450);
nand U21137 (N_21137,N_19551,N_15811);
nor U21138 (N_21138,N_17051,N_19449);
or U21139 (N_21139,N_19918,N_18448);
xnor U21140 (N_21140,N_17665,N_19614);
nand U21141 (N_21141,N_19988,N_15489);
and U21142 (N_21142,N_19807,N_16122);
or U21143 (N_21143,N_19839,N_16534);
and U21144 (N_21144,N_19331,N_19132);
or U21145 (N_21145,N_16661,N_19057);
nor U21146 (N_21146,N_17350,N_16341);
nor U21147 (N_21147,N_16349,N_19608);
nand U21148 (N_21148,N_19412,N_17906);
nand U21149 (N_21149,N_19749,N_15805);
nor U21150 (N_21150,N_19178,N_16919);
nor U21151 (N_21151,N_18734,N_18550);
nand U21152 (N_21152,N_17397,N_18684);
and U21153 (N_21153,N_15993,N_19625);
and U21154 (N_21154,N_19618,N_17022);
nand U21155 (N_21155,N_16494,N_19159);
nand U21156 (N_21156,N_19496,N_19362);
and U21157 (N_21157,N_17633,N_16679);
nor U21158 (N_21158,N_15951,N_19328);
nor U21159 (N_21159,N_19342,N_17357);
nand U21160 (N_21160,N_15815,N_19407);
nand U21161 (N_21161,N_17601,N_15461);
nor U21162 (N_21162,N_18481,N_15641);
xnor U21163 (N_21163,N_17793,N_15465);
xor U21164 (N_21164,N_18998,N_16934);
nand U21165 (N_21165,N_16629,N_15912);
and U21166 (N_21166,N_16518,N_19998);
and U21167 (N_21167,N_16540,N_19610);
or U21168 (N_21168,N_15425,N_19714);
and U21169 (N_21169,N_18213,N_15295);
and U21170 (N_21170,N_16542,N_18473);
and U21171 (N_21171,N_17393,N_17711);
nand U21172 (N_21172,N_18065,N_18581);
nand U21173 (N_21173,N_17967,N_15537);
nor U21174 (N_21174,N_19936,N_18228);
nand U21175 (N_21175,N_19196,N_18941);
nor U21176 (N_21176,N_16939,N_16401);
and U21177 (N_21177,N_17995,N_16207);
nor U21178 (N_21178,N_15277,N_15018);
nor U21179 (N_21179,N_17767,N_15750);
nor U21180 (N_21180,N_19454,N_15468);
nor U21181 (N_21181,N_17923,N_17159);
nor U21182 (N_21182,N_17381,N_17498);
xnor U21183 (N_21183,N_17766,N_19280);
and U21184 (N_21184,N_18972,N_15268);
and U21185 (N_21185,N_17150,N_16130);
or U21186 (N_21186,N_17636,N_16143);
xor U21187 (N_21187,N_19825,N_17614);
and U21188 (N_21188,N_19275,N_16311);
xnor U21189 (N_21189,N_19167,N_15941);
or U21190 (N_21190,N_15900,N_19123);
nand U21191 (N_21191,N_19833,N_15481);
or U21192 (N_21192,N_19771,N_17011);
and U21193 (N_21193,N_17851,N_15017);
nand U21194 (N_21194,N_18258,N_18813);
and U21195 (N_21195,N_17158,N_18985);
nor U21196 (N_21196,N_19654,N_17490);
nand U21197 (N_21197,N_17389,N_15804);
nand U21198 (N_21198,N_15783,N_15482);
nand U21199 (N_21199,N_18620,N_18311);
or U21200 (N_21200,N_16873,N_17009);
nor U21201 (N_21201,N_19760,N_17854);
xnor U21202 (N_21202,N_19575,N_18917);
nand U21203 (N_21203,N_18862,N_15535);
or U21204 (N_21204,N_18514,N_18737);
nand U21205 (N_21205,N_16147,N_19101);
nand U21206 (N_21206,N_17242,N_18934);
nor U21207 (N_21207,N_15398,N_19156);
nor U21208 (N_21208,N_19077,N_17119);
and U21209 (N_21209,N_17777,N_17522);
or U21210 (N_21210,N_15067,N_18789);
or U21211 (N_21211,N_15559,N_16537);
nor U21212 (N_21212,N_19458,N_18386);
nand U21213 (N_21213,N_17483,N_18996);
and U21214 (N_21214,N_15752,N_19154);
and U21215 (N_21215,N_18563,N_17235);
and U21216 (N_21216,N_17014,N_17770);
nand U21217 (N_21217,N_15699,N_19538);
nand U21218 (N_21218,N_17116,N_18222);
or U21219 (N_21219,N_15139,N_15607);
or U21220 (N_21220,N_18394,N_17723);
nand U21221 (N_21221,N_16588,N_16660);
or U21222 (N_21222,N_15984,N_16794);
and U21223 (N_21223,N_18154,N_17413);
or U21224 (N_21224,N_17462,N_17564);
and U21225 (N_21225,N_18014,N_16915);
nand U21226 (N_21226,N_19511,N_16844);
or U21227 (N_21227,N_19038,N_16888);
xor U21228 (N_21228,N_16162,N_19312);
or U21229 (N_21229,N_17100,N_16090);
and U21230 (N_21230,N_19040,N_18588);
nand U21231 (N_21231,N_16969,N_18153);
or U21232 (N_21232,N_18243,N_18410);
nor U21233 (N_21233,N_16344,N_18994);
xnor U21234 (N_21234,N_19216,N_16099);
or U21235 (N_21235,N_18651,N_15639);
or U21236 (N_21236,N_19202,N_17542);
and U21237 (N_21237,N_18800,N_17670);
or U21238 (N_21238,N_16776,N_15162);
nand U21239 (N_21239,N_17316,N_19550);
nor U21240 (N_21240,N_17743,N_15891);
xor U21241 (N_21241,N_18115,N_15332);
or U21242 (N_21242,N_15044,N_15749);
nand U21243 (N_21243,N_18501,N_15496);
and U21244 (N_21244,N_16013,N_16725);
xor U21245 (N_21245,N_17785,N_15631);
xor U21246 (N_21246,N_15905,N_18105);
or U21247 (N_21247,N_18697,N_17085);
nand U21248 (N_21248,N_19418,N_18455);
and U21249 (N_21249,N_19683,N_17225);
and U21250 (N_21250,N_16016,N_18653);
nand U21251 (N_21251,N_15129,N_17548);
nor U21252 (N_21252,N_19169,N_15103);
nand U21253 (N_21253,N_17313,N_17768);
nor U21254 (N_21254,N_19053,N_18804);
nor U21255 (N_21255,N_17390,N_17332);
xor U21256 (N_21256,N_17864,N_18702);
xnor U21257 (N_21257,N_15324,N_19457);
and U21258 (N_21258,N_18890,N_19785);
nand U21259 (N_21259,N_19629,N_19314);
or U21260 (N_21260,N_19350,N_16560);
or U21261 (N_21261,N_15595,N_19874);
or U21262 (N_21262,N_19798,N_17190);
nand U21263 (N_21263,N_17622,N_16465);
xnor U21264 (N_21264,N_16905,N_15651);
nor U21265 (N_21265,N_17754,N_16787);
and U21266 (N_21266,N_15455,N_15160);
and U21267 (N_21267,N_15972,N_18025);
nor U21268 (N_21268,N_18368,N_15668);
xor U21269 (N_21269,N_18186,N_15282);
nor U21270 (N_21270,N_19633,N_15785);
or U21271 (N_21271,N_15911,N_18624);
nor U21272 (N_21272,N_18019,N_18851);
and U21273 (N_21273,N_16636,N_17716);
nand U21274 (N_21274,N_15611,N_19695);
nor U21275 (N_21275,N_16708,N_18336);
nand U21276 (N_21276,N_17786,N_16399);
or U21277 (N_21277,N_16669,N_16996);
nor U21278 (N_21278,N_17640,N_16211);
xnor U21279 (N_21279,N_15161,N_16413);
and U21280 (N_21280,N_15563,N_18197);
nor U21281 (N_21281,N_15068,N_15587);
or U21282 (N_21282,N_15927,N_15729);
or U21283 (N_21283,N_19356,N_16209);
and U21284 (N_21284,N_18060,N_18244);
and U21285 (N_21285,N_15377,N_19267);
and U21286 (N_21286,N_18485,N_15141);
or U21287 (N_21287,N_17126,N_18070);
and U21288 (N_21288,N_15350,N_16795);
nor U21289 (N_21289,N_17166,N_15999);
nand U21290 (N_21290,N_15658,N_19469);
nor U21291 (N_21291,N_18402,N_16363);
nor U21292 (N_21292,N_15601,N_16701);
or U21293 (N_21293,N_16215,N_19886);
nand U21294 (N_21294,N_17734,N_19993);
xor U21295 (N_21295,N_16876,N_17737);
nand U21296 (N_21296,N_15780,N_15291);
xnor U21297 (N_21297,N_17637,N_19005);
or U21298 (N_21298,N_17409,N_15372);
or U21299 (N_21299,N_15767,N_17870);
xor U21300 (N_21300,N_19793,N_15260);
and U21301 (N_21301,N_17170,N_16931);
and U21302 (N_21302,N_16555,N_16854);
xor U21303 (N_21303,N_17718,N_15030);
and U21304 (N_21304,N_16167,N_17056);
nor U21305 (N_21305,N_18159,N_16902);
or U21306 (N_21306,N_18925,N_17523);
nor U21307 (N_21307,N_19773,N_18920);
nor U21308 (N_21308,N_18700,N_15637);
or U21309 (N_21309,N_19669,N_17717);
nor U21310 (N_21310,N_19397,N_17179);
xnor U21311 (N_21311,N_19780,N_18660);
xnor U21312 (N_21312,N_17057,N_18216);
or U21313 (N_21313,N_18686,N_16879);
nand U21314 (N_21314,N_19322,N_16330);
nand U21315 (N_21315,N_17317,N_17780);
nor U21316 (N_21316,N_16397,N_15698);
or U21317 (N_21317,N_19824,N_18672);
nand U21318 (N_21318,N_15843,N_15135);
or U21319 (N_21319,N_15784,N_18009);
nand U21320 (N_21320,N_17605,N_17419);
or U21321 (N_21321,N_15118,N_15471);
xnor U21322 (N_21322,N_16440,N_17189);
xnor U21323 (N_21323,N_18472,N_18513);
or U21324 (N_21324,N_16227,N_19171);
and U21325 (N_21325,N_15472,N_19054);
nor U21326 (N_21326,N_15316,N_16319);
xnor U21327 (N_21327,N_19390,N_17154);
or U21328 (N_21328,N_15013,N_15335);
or U21329 (N_21329,N_16880,N_18449);
nor U21330 (N_21330,N_18963,N_19934);
and U21331 (N_21331,N_15131,N_15754);
or U21332 (N_21332,N_18083,N_19016);
nand U21333 (N_21333,N_19210,N_19174);
and U21334 (N_21334,N_15183,N_18663);
nor U21335 (N_21335,N_16004,N_17902);
or U21336 (N_21336,N_17899,N_17110);
and U21337 (N_21337,N_16533,N_18055);
and U21338 (N_21338,N_18774,N_15605);
or U21339 (N_21339,N_16451,N_17285);
nand U21340 (N_21340,N_18086,N_16739);
nand U21341 (N_21341,N_15646,N_18018);
nand U21342 (N_21342,N_15203,N_15226);
nor U21343 (N_21343,N_16535,N_19598);
and U21344 (N_21344,N_19301,N_19411);
nor U21345 (N_21345,N_18760,N_19651);
nor U21346 (N_21346,N_17647,N_17195);
xor U21347 (N_21347,N_15487,N_18791);
nand U21348 (N_21348,N_15730,N_18250);
or U21349 (N_21349,N_17083,N_19960);
or U21350 (N_21350,N_18058,N_19688);
nand U21351 (N_21351,N_19427,N_15258);
xor U21352 (N_21352,N_19929,N_18291);
and U21353 (N_21353,N_16118,N_19991);
and U21354 (N_21354,N_19953,N_16893);
or U21355 (N_21355,N_16571,N_18756);
nand U21356 (N_21356,N_19915,N_18675);
nand U21357 (N_21357,N_18610,N_17850);
or U21358 (N_21358,N_18442,N_17977);
nand U21359 (N_21359,N_17735,N_16762);
nor U21360 (N_21360,N_18595,N_16415);
and U21361 (N_21361,N_18282,N_15793);
nand U21362 (N_21362,N_18223,N_19323);
xnor U21363 (N_21363,N_17510,N_19244);
and U21364 (N_21364,N_19461,N_19083);
and U21365 (N_21365,N_18454,N_17495);
or U21366 (N_21366,N_16022,N_19535);
xnor U21367 (N_21367,N_16007,N_18329);
nor U21368 (N_21368,N_18068,N_16665);
nor U21369 (N_21369,N_19978,N_15254);
nand U21370 (N_21370,N_15561,N_15094);
nand U21371 (N_21371,N_16800,N_15600);
nand U21372 (N_21372,N_18661,N_17205);
or U21373 (N_21373,N_16820,N_15532);
nand U21374 (N_21374,N_17791,N_19269);
and U21375 (N_21375,N_18632,N_17951);
nor U21376 (N_21376,N_16896,N_19676);
and U21377 (N_21377,N_16754,N_18822);
and U21378 (N_21378,N_15619,N_17965);
nand U21379 (N_21379,N_18263,N_17519);
or U21380 (N_21380,N_15515,N_15185);
xnor U21381 (N_21381,N_15483,N_15473);
nand U21382 (N_21382,N_16500,N_16478);
nor U21383 (N_21383,N_18471,N_19652);
xor U21384 (N_21384,N_19904,N_15895);
nand U21385 (N_21385,N_19659,N_16499);
nor U21386 (N_21386,N_16684,N_18033);
or U21387 (N_21387,N_16150,N_15319);
and U21388 (N_21388,N_19271,N_18378);
and U21389 (N_21389,N_16173,N_15207);
nand U21390 (N_21390,N_16115,N_17699);
nor U21391 (N_21391,N_17760,N_16778);
and U21392 (N_21392,N_16759,N_16237);
nor U21393 (N_21393,N_16074,N_16930);
nand U21394 (N_21394,N_16416,N_17830);
nand U21395 (N_21395,N_15184,N_18764);
nor U21396 (N_21396,N_16601,N_15142);
or U21397 (N_21397,N_15436,N_16189);
xnor U21398 (N_21398,N_17433,N_19278);
nor U21399 (N_21399,N_19865,N_16671);
or U21400 (N_21400,N_19165,N_16532);
or U21401 (N_21401,N_18112,N_17611);
and U21402 (N_21402,N_17978,N_16443);
nor U21403 (N_21403,N_19238,N_17568);
or U21404 (N_21404,N_17945,N_18902);
and U21405 (N_21405,N_18444,N_19660);
nor U21406 (N_21406,N_17493,N_16081);
or U21407 (N_21407,N_19370,N_15869);
nor U21408 (N_21408,N_15307,N_17143);
and U21409 (N_21409,N_18208,N_19542);
nor U21410 (N_21410,N_19306,N_16035);
nand U21411 (N_21411,N_16142,N_15902);
and U21412 (N_21412,N_17820,N_18251);
or U21413 (N_21413,N_17442,N_16014);
or U21414 (N_21414,N_18348,N_16111);
nand U21415 (N_21415,N_19272,N_18099);
or U21416 (N_21416,N_17295,N_16579);
and U21417 (N_21417,N_17588,N_16750);
nand U21418 (N_21418,N_15444,N_15952);
or U21419 (N_21419,N_17379,N_17629);
or U21420 (N_21420,N_17657,N_17868);
nand U21421 (N_21421,N_16257,N_16756);
or U21422 (N_21422,N_18369,N_18826);
nand U21423 (N_21423,N_16085,N_19981);
nand U21424 (N_21424,N_17006,N_16575);
and U21425 (N_21425,N_17004,N_19389);
nand U21426 (N_21426,N_18071,N_17107);
nand U21427 (N_21427,N_16159,N_17304);
and U21428 (N_21428,N_17367,N_15510);
and U21429 (N_21429,N_16658,N_16681);
or U21430 (N_21430,N_17556,N_17395);
xnor U21431 (N_21431,N_18546,N_18121);
or U21432 (N_21432,N_16755,N_15365);
nand U21433 (N_21433,N_17562,N_16948);
xor U21434 (N_21434,N_19424,N_15136);
nor U21435 (N_21435,N_15621,N_19175);
or U21436 (N_21436,N_15176,N_19492);
or U21437 (N_21437,N_15321,N_19368);
nor U21438 (N_21438,N_18896,N_18953);
and U21439 (N_21439,N_19943,N_19577);
and U21440 (N_21440,N_18722,N_16586);
and U21441 (N_21441,N_19814,N_15070);
or U21442 (N_21442,N_16328,N_16806);
or U21443 (N_21443,N_17366,N_16866);
nor U21444 (N_21444,N_18843,N_16152);
nor U21445 (N_21445,N_18409,N_15206);
nor U21446 (N_21446,N_15901,N_16153);
or U21447 (N_21447,N_19447,N_15862);
xnor U21448 (N_21448,N_16955,N_19304);
or U21449 (N_21449,N_19110,N_19919);
and U21450 (N_21450,N_15062,N_15409);
nand U21451 (N_21451,N_18542,N_18236);
nor U21452 (N_21452,N_16566,N_16132);
nand U21453 (N_21453,N_18283,N_17160);
and U21454 (N_21454,N_19152,N_17586);
nand U21455 (N_21455,N_15123,N_17592);
nor U21456 (N_21456,N_15193,N_16254);
and U21457 (N_21457,N_18559,N_18999);
or U21458 (N_21458,N_15024,N_17778);
or U21459 (N_21459,N_18199,N_18669);
and U21460 (N_21460,N_18450,N_18264);
and U21461 (N_21461,N_19026,N_15828);
or U21462 (N_21462,N_17124,N_16498);
nor U21463 (N_21463,N_17828,N_17888);
or U21464 (N_21464,N_19708,N_18307);
nand U21465 (N_21465,N_18272,N_18482);
nor U21466 (N_21466,N_17950,N_17375);
or U21467 (N_21467,N_16105,N_15747);
nor U21468 (N_21468,N_15579,N_15643);
and U21469 (N_21469,N_18463,N_19641);
nor U21470 (N_21470,N_18006,N_17953);
or U21471 (N_21471,N_16772,N_16544);
or U21472 (N_21472,N_16200,N_18733);
or U21473 (N_21473,N_15458,N_16824);
nor U21474 (N_21474,N_18294,N_17021);
nand U21475 (N_21475,N_16638,N_16769);
or U21476 (N_21476,N_18880,N_15703);
and U21477 (N_21477,N_18362,N_19697);
nor U21478 (N_21478,N_17858,N_16786);
and U21479 (N_21479,N_15910,N_19858);
nor U21480 (N_21480,N_17145,N_19260);
xor U21481 (N_21481,N_16034,N_18778);
nand U21482 (N_21482,N_18562,N_17121);
nand U21483 (N_21483,N_17187,N_16900);
and U21484 (N_21484,N_15642,N_18211);
xnor U21485 (N_21485,N_16855,N_16922);
nor U21486 (N_21486,N_15740,N_15979);
or U21487 (N_21487,N_17326,N_15050);
or U21488 (N_21488,N_19590,N_19042);
or U21489 (N_21489,N_15708,N_17810);
nand U21490 (N_21490,N_17862,N_19559);
nand U21491 (N_21491,N_19768,N_16148);
nand U21492 (N_21492,N_18899,N_17648);
and U21493 (N_21493,N_19069,N_18359);
xor U21494 (N_21494,N_17746,N_19353);
or U21495 (N_21495,N_18383,N_16060);
nor U21496 (N_21496,N_17153,N_19209);
and U21497 (N_21497,N_19010,N_18439);
or U21498 (N_21498,N_16470,N_19190);
nor U21499 (N_21499,N_15517,N_18039);
and U21500 (N_21500,N_19025,N_18647);
and U21501 (N_21501,N_15801,N_16496);
xnor U21502 (N_21502,N_16245,N_15217);
nor U21503 (N_21503,N_19138,N_19052);
nand U21504 (N_21504,N_17969,N_18828);
and U21505 (N_21505,N_16420,N_19979);
and U21506 (N_21506,N_19817,N_19332);
or U21507 (N_21507,N_18398,N_18966);
and U21508 (N_21508,N_15710,N_18691);
or U21509 (N_21509,N_15428,N_16577);
nand U21510 (N_21510,N_19232,N_18422);
xnor U21511 (N_21511,N_16135,N_18269);
and U21512 (N_21512,N_17206,N_16100);
or U21513 (N_21513,N_18355,N_15100);
nor U21514 (N_21514,N_19377,N_19699);
or U21515 (N_21515,N_16425,N_18739);
and U21516 (N_21516,N_16342,N_18919);
nand U21517 (N_21517,N_16986,N_16387);
or U21518 (N_21518,N_15508,N_15328);
nand U21519 (N_21519,N_15610,N_18571);
nand U21520 (N_21520,N_17072,N_16760);
nand U21521 (N_21521,N_17533,N_18796);
nor U21522 (N_21522,N_16731,N_15824);
or U21523 (N_21523,N_18538,N_19488);
and U21524 (N_21524,N_17733,N_17509);
xor U21525 (N_21525,N_16723,N_16077);
nand U21526 (N_21526,N_16839,N_15497);
or U21527 (N_21527,N_17043,N_19692);
nor U21528 (N_21528,N_16423,N_18986);
and U21529 (N_21529,N_17671,N_16815);
nor U21530 (N_21530,N_18580,N_19937);
or U21531 (N_21531,N_16389,N_18276);
nand U21532 (N_21532,N_19881,N_16624);
xor U21533 (N_21533,N_19468,N_15998);
nand U21534 (N_21534,N_15713,N_16469);
or U21535 (N_21535,N_17423,N_15227);
nand U21536 (N_21536,N_18787,N_15071);
nand U21537 (N_21537,N_15325,N_17988);
xnor U21538 (N_21538,N_17279,N_16529);
or U21539 (N_21539,N_16753,N_16685);
or U21540 (N_21540,N_18492,N_18353);
and U21541 (N_21541,N_17726,N_15219);
nor U21542 (N_21542,N_18709,N_15063);
nor U21543 (N_21543,N_18740,N_15429);
xnor U21544 (N_21544,N_17822,N_16400);
and U21545 (N_21545,N_16039,N_16598);
nand U21546 (N_21546,N_15337,N_19104);
and U21547 (N_21547,N_18220,N_19364);
nand U21548 (N_21548,N_19605,N_15664);
nor U21549 (N_21549,N_16114,N_15735);
nand U21550 (N_21550,N_17297,N_18094);
or U21551 (N_21551,N_15985,N_19012);
nor U21552 (N_21552,N_18655,N_19379);
nand U21553 (N_21553,N_15822,N_16508);
and U21554 (N_21554,N_15701,N_16006);
nand U21555 (N_21555,N_18782,N_17090);
nand U21556 (N_21556,N_19125,N_15851);
nand U21557 (N_21557,N_15723,N_17453);
or U21558 (N_21558,N_19071,N_15879);
or U21559 (N_21559,N_18516,N_17959);
and U21560 (N_21560,N_17947,N_18468);
nand U21561 (N_21561,N_18809,N_15635);
nor U21562 (N_21562,N_19624,N_19716);
xor U21563 (N_21563,N_16615,N_16729);
xnor U21564 (N_21564,N_16172,N_16398);
and U21565 (N_21565,N_15856,N_15378);
xnor U21566 (N_21566,N_18426,N_19848);
nand U21567 (N_21567,N_16070,N_16840);
nand U21568 (N_21568,N_18436,N_16763);
or U21569 (N_21569,N_18229,N_17485);
xor U21570 (N_21570,N_15976,N_17799);
and U21571 (N_21571,N_17008,N_16284);
and U21572 (N_21572,N_15417,N_18717);
and U21573 (N_21573,N_16049,N_15768);
nand U21574 (N_21574,N_16599,N_15251);
and U21575 (N_21575,N_17491,N_16633);
or U21576 (N_21576,N_17932,N_17136);
nor U21577 (N_21577,N_19299,N_19701);
nand U21578 (N_21578,N_19607,N_17876);
nor U21579 (N_21579,N_17003,N_18770);
xnor U21580 (N_21580,N_15781,N_16606);
nand U21581 (N_21581,N_19231,N_19631);
xnor U21582 (N_21582,N_18762,N_17911);
xor U21583 (N_21583,N_17220,N_18803);
or U21584 (N_21584,N_15992,N_17302);
and U21585 (N_21585,N_17554,N_15947);
xnor U21586 (N_21586,N_15568,N_19235);
xnor U21587 (N_21587,N_17652,N_19678);
or U21588 (N_21588,N_16721,N_18713);
and U21589 (N_21589,N_16144,N_17608);
nor U21590 (N_21590,N_16324,N_19601);
xor U21591 (N_21591,N_15697,N_19473);
nand U21592 (N_21592,N_18167,N_19962);
or U21593 (N_21593,N_15629,N_19655);
nor U21594 (N_21594,N_16018,N_15971);
nor U21595 (N_21595,N_15825,N_18543);
nand U21596 (N_21596,N_19265,N_18626);
nor U21597 (N_21597,N_16288,N_17982);
xnor U21598 (N_21598,N_15059,N_17299);
or U21599 (N_21599,N_17387,N_19383);
nand U21600 (N_21600,N_19347,N_16591);
or U21601 (N_21601,N_17135,N_19009);
and U21602 (N_21602,N_19954,N_17151);
and U21603 (N_21603,N_16410,N_16670);
xor U21604 (N_21604,N_17627,N_19916);
nor U21605 (N_21605,N_18609,N_19658);
nand U21606 (N_21606,N_19566,N_16906);
nand U21607 (N_21607,N_15906,N_19127);
nand U21608 (N_21608,N_15265,N_16519);
and U21609 (N_21609,N_19792,N_19642);
nor U21610 (N_21610,N_17098,N_15803);
xor U21611 (N_21611,N_15987,N_16634);
or U21612 (N_21612,N_18309,N_17532);
or U21613 (N_21613,N_15340,N_18191);
nor U21614 (N_21614,N_17659,N_17541);
or U21615 (N_21615,N_19809,N_19907);
nor U21616 (N_21616,N_19495,N_19520);
and U21617 (N_21617,N_18192,N_19103);
or U21618 (N_21618,N_18551,N_17306);
nor U21619 (N_21619,N_16643,N_15691);
nor U21620 (N_21620,N_18531,N_17405);
xor U21621 (N_21621,N_17230,N_16477);
and U21622 (N_21622,N_16419,N_18945);
nand U21623 (N_21623,N_16538,N_17134);
or U21624 (N_21624,N_19479,N_18182);
or U21625 (N_21625,N_17239,N_15898);
nand U21626 (N_21626,N_18235,N_16513);
nand U21627 (N_21627,N_19514,N_18381);
or U21628 (N_21628,N_18395,N_18969);
or U21629 (N_21629,N_16526,N_18668);
and U21630 (N_21630,N_15812,N_16613);
nor U21631 (N_21631,N_18128,N_16961);
or U21632 (N_21632,N_16183,N_15099);
and U21633 (N_21633,N_15762,N_18958);
nor U21634 (N_21634,N_17383,N_18615);
nand U21635 (N_21635,N_19911,N_16889);
nor U21636 (N_21636,N_17638,N_16290);
and U21637 (N_21637,N_16603,N_15547);
xnor U21638 (N_21638,N_16466,N_19002);
nand U21639 (N_21639,N_18973,N_18732);
nor U21640 (N_21640,N_16826,N_15146);
nand U21641 (N_21641,N_15808,N_19212);
or U21642 (N_21642,N_18955,N_17402);
xor U21643 (N_21643,N_15847,N_17216);
nand U21644 (N_21644,N_15439,N_15677);
nand U21645 (N_21645,N_17192,N_19155);
nand U21646 (N_21646,N_15655,N_17801);
and U21647 (N_21647,N_16958,N_15040);
or U21648 (N_21648,N_18109,N_16668);
or U21649 (N_21649,N_17626,N_16909);
and U21650 (N_21650,N_16700,N_17401);
or U21651 (N_21651,N_15342,N_19812);
xor U21652 (N_21652,N_19463,N_18152);
nor U21653 (N_21653,N_17686,N_16119);
nand U21654 (N_21654,N_15848,N_15519);
xnor U21655 (N_21655,N_17148,N_18887);
nor U21656 (N_21656,N_15494,N_17251);
or U21657 (N_21657,N_16973,N_17604);
or U21658 (N_21658,N_15333,N_16487);
nor U21659 (N_21659,N_15725,N_16539);
nand U21660 (N_21660,N_16744,N_17954);
nand U21661 (N_21661,N_16576,N_18456);
or U21662 (N_21662,N_19404,N_19455);
and U21663 (N_21663,N_17209,N_15539);
or U21664 (N_21664,N_16066,N_19935);
nand U21665 (N_21665,N_18726,N_17091);
nand U21666 (N_21666,N_19992,N_18654);
and U21667 (N_21667,N_15110,N_15771);
nor U21668 (N_21668,N_15480,N_19560);
nand U21669 (N_21669,N_19112,N_18962);
and U21670 (N_21670,N_15165,N_17505);
or U21671 (N_21671,N_17994,N_18908);
nand U21672 (N_21672,N_18926,N_19756);
nand U21673 (N_21673,N_15550,N_17123);
and U21674 (N_21674,N_19062,N_19719);
or U21675 (N_21675,N_15663,N_18583);
and U21676 (N_21676,N_16991,N_17127);
or U21677 (N_21677,N_15836,N_17675);
or U21678 (N_21678,N_16509,N_18944);
nor U21679 (N_21679,N_16782,N_18262);
nor U21680 (N_21680,N_15748,N_15904);
nand U21681 (N_21681,N_17430,N_19619);
and U21682 (N_21682,N_15469,N_15797);
nor U21683 (N_21683,N_17305,N_16630);
nand U21684 (N_21684,N_19258,N_16745);
nand U21685 (N_21685,N_16403,N_19015);
and U21686 (N_21686,N_17184,N_17573);
nor U21687 (N_21687,N_16741,N_16611);
and U21688 (N_21688,N_16798,N_16626);
xor U21689 (N_21689,N_16635,N_17263);
nor U21690 (N_21690,N_16411,N_17352);
and U21691 (N_21691,N_17621,N_19627);
nand U21692 (N_21692,N_16924,N_17118);
nor U21693 (N_21693,N_15081,N_15182);
nor U21694 (N_21694,N_19187,N_15960);
nor U21695 (N_21695,N_18794,N_16104);
and U21696 (N_21696,N_16430,N_17172);
or U21697 (N_21697,N_19547,N_17477);
or U21698 (N_21698,N_18416,N_16490);
or U21699 (N_21699,N_18142,N_17034);
nand U21700 (N_21700,N_19644,N_18718);
xor U21701 (N_21701,N_19783,N_19665);
nand U21702 (N_21702,N_16639,N_17296);
nand U21703 (N_21703,N_17948,N_17374);
or U21704 (N_21704,N_15113,N_16282);
or U21705 (N_21705,N_18194,N_16370);
and U21706 (N_21706,N_18861,N_16903);
or U21707 (N_21707,N_18345,N_15673);
and U21708 (N_21708,N_18807,N_15036);
nor U21709 (N_21709,N_15876,N_17452);
nand U21710 (N_21710,N_19653,N_18203);
and U21711 (N_21711,N_15526,N_18757);
or U21712 (N_21712,N_17484,N_19730);
nor U21713 (N_21713,N_19680,N_17165);
nor U21714 (N_21714,N_18792,N_15388);
or U21715 (N_21715,N_19325,N_15315);
or U21716 (N_21716,N_18783,N_16468);
or U21717 (N_21717,N_18839,N_17265);
nand U21718 (N_21718,N_15511,N_17243);
nand U21719 (N_21719,N_16460,N_18030);
nand U21720 (N_21720,N_15049,N_17783);
and U21721 (N_21721,N_15792,N_15145);
or U21722 (N_21722,N_19769,N_16412);
or U21723 (N_21723,N_15887,N_19041);
nand U21724 (N_21724,N_16946,N_15270);
or U21725 (N_21725,N_16783,N_18387);
xnor U21726 (N_21726,N_15404,N_17587);
nand U21727 (N_21727,N_19398,N_15273);
nor U21728 (N_21728,N_16174,N_16170);
and U21729 (N_21729,N_18950,N_18883);
nor U21730 (N_21730,N_17346,N_19137);
nand U21731 (N_21731,N_17210,N_18592);
and U21732 (N_21732,N_17903,N_15558);
and U21733 (N_21733,N_19336,N_18458);
xnor U21734 (N_21734,N_16680,N_18903);
nor U21735 (N_21735,N_15584,N_19776);
nor U21736 (N_21736,N_18125,N_17463);
nand U21737 (N_21737,N_16103,N_16841);
and U21738 (N_21738,N_18056,N_15023);
nand U21739 (N_21739,N_19556,N_18555);
nand U21740 (N_21740,N_15665,N_19787);
or U21741 (N_21741,N_16827,N_15283);
nand U21742 (N_21742,N_19113,N_15934);
xor U21743 (N_21743,N_18884,N_19122);
nor U21744 (N_21744,N_17018,N_18618);
nand U21745 (N_21745,N_19600,N_19615);
or U21746 (N_21746,N_15495,N_19616);
or U21747 (N_21747,N_19163,N_19065);
or U21748 (N_21748,N_19021,N_18652);
and U21749 (N_21749,N_19941,N_18569);
nor U21750 (N_21750,N_15739,N_18979);
and U21751 (N_21751,N_18374,N_16994);
or U21752 (N_21752,N_15407,N_18103);
xor U21753 (N_21753,N_19717,N_16993);
nand U21754 (N_21754,N_15696,N_19536);
and U21755 (N_21755,N_16497,N_17525);
xnor U21756 (N_21756,N_17781,N_17926);
and U21757 (N_21757,N_19638,N_15379);
nor U21758 (N_21758,N_15921,N_19876);
nand U21759 (N_21759,N_15995,N_16359);
xnor U21760 (N_21760,N_15220,N_16775);
and U21761 (N_21761,N_17125,N_17569);
or U21762 (N_21762,N_15122,N_18187);
and U21763 (N_21763,N_19310,N_18594);
nor U21764 (N_21764,N_19476,N_17744);
nand U21765 (N_21765,N_19573,N_16689);
nand U21766 (N_21766,N_16527,N_17097);
and U21767 (N_21767,N_15571,N_17695);
and U21768 (N_21768,N_17429,N_17113);
nand U21769 (N_21769,N_15234,N_19501);
or U21770 (N_21770,N_15846,N_16139);
nand U21771 (N_21771,N_17660,N_17944);
nand U21772 (N_21772,N_19576,N_17291);
and U21773 (N_21773,N_19893,N_17998);
or U21774 (N_21774,N_15957,N_17826);
or U21775 (N_21775,N_17935,N_15577);
and U21776 (N_21776,N_19647,N_16268);
or U21777 (N_21777,N_17620,N_17956);
or U21778 (N_21778,N_17213,N_16568);
and U21779 (N_21779,N_16384,N_19076);
nand U21780 (N_21780,N_16221,N_17310);
or U21781 (N_21781,N_15245,N_16528);
or U21782 (N_21782,N_17042,N_18907);
xor U21783 (N_21783,N_16796,N_15290);
nand U21784 (N_21784,N_17322,N_18827);
nor U21785 (N_21785,N_16292,N_15769);
nand U21786 (N_21786,N_15190,N_15047);
and U21787 (N_21787,N_18933,N_18719);
nand U21788 (N_21788,N_18560,N_15456);
or U21789 (N_21789,N_18914,N_15107);
nor U21790 (N_21790,N_17650,N_19628);
or U21791 (N_21791,N_19924,N_15225);
xnor U21792 (N_21792,N_18987,N_15163);
or U21793 (N_21793,N_15490,N_19620);
nand U21794 (N_21794,N_15627,N_15498);
or U21795 (N_21795,N_15670,N_15782);
and U21796 (N_21796,N_16001,N_17790);
nor U21797 (N_21797,N_16051,N_15393);
xnor U21798 (N_21798,N_15271,N_17553);
xor U21799 (N_21799,N_19185,N_19460);
or U21800 (N_21800,N_17917,N_17363);
or U21801 (N_21801,N_17249,N_19806);
or U21802 (N_21802,N_16057,N_17365);
and U21803 (N_21803,N_18200,N_15387);
nor U21804 (N_21804,N_16120,N_19266);
nand U21805 (N_21805,N_19878,N_19229);
nand U21806 (N_21806,N_16274,N_17256);
nor U21807 (N_21807,N_18275,N_19975);
nor U21808 (N_21808,N_17330,N_18553);
or U21809 (N_21809,N_17856,N_19770);
and U21810 (N_21810,N_17282,N_19337);
nor U21811 (N_21811,N_18110,N_19700);
and U21812 (N_21812,N_17684,N_15687);
nand U21813 (N_21813,N_19920,N_19702);
nand U21814 (N_21814,N_15090,N_19220);
or U21815 (N_21815,N_16063,N_15313);
or U21816 (N_21816,N_18206,N_15195);
or U21817 (N_21817,N_15678,N_19243);
nand U21818 (N_21818,N_17784,N_19930);
nor U21819 (N_21819,N_16357,N_18922);
xor U21820 (N_21820,N_18342,N_18863);
nor U21821 (N_21821,N_15440,N_17273);
or U21822 (N_21822,N_17844,N_16554);
nand U21823 (N_21823,N_16356,N_16531);
and U21824 (N_21824,N_19725,N_15572);
or U21825 (N_21825,N_15086,N_15928);
nand U21826 (N_21826,N_18082,N_19166);
nand U21827 (N_21827,N_19729,N_16891);
nor U21828 (N_21828,N_19519,N_15314);
nand U21829 (N_21829,N_18505,N_17990);
nor U21830 (N_21830,N_18754,N_19056);
xor U21831 (N_21831,N_16556,N_15521);
or U21832 (N_21832,N_16932,N_17434);
xor U21833 (N_21833,N_17174,N_16683);
and U21834 (N_21834,N_16793,N_16511);
nand U21835 (N_21835,N_15875,N_18818);
nor U21836 (N_21836,N_15569,N_16309);
nor U21837 (N_21837,N_16367,N_17096);
nand U21838 (N_21838,N_17811,N_15051);
and U21839 (N_21839,N_17515,N_16435);
nand U21840 (N_21840,N_16541,N_16431);
nor U21841 (N_21841,N_19532,N_18695);
or U21842 (N_21842,N_17955,N_19748);
nor U21843 (N_21843,N_15598,N_19808);
xnor U21844 (N_21844,N_17312,N_19376);
nor U21845 (N_21845,N_18557,N_17693);
nor U21846 (N_21846,N_17730,N_19989);
and U21847 (N_21847,N_18013,N_18679);
nor U21848 (N_21848,N_16080,N_15850);
xor U21849 (N_21849,N_16585,N_19713);
nor U21850 (N_21850,N_19467,N_15818);
or U21851 (N_21851,N_18617,N_18915);
nor U21852 (N_21852,N_15418,N_19253);
and U21853 (N_21853,N_19758,N_15028);
or U21854 (N_21854,N_18859,N_19366);
xor U21855 (N_21855,N_19066,N_19307);
or U21856 (N_21856,N_18830,N_19329);
nand U21857 (N_21857,N_18881,N_19570);
nor U21858 (N_21858,N_15555,N_17916);
nand U21859 (N_21859,N_17268,N_19433);
or U21860 (N_21860,N_17075,N_17673);
nor U21861 (N_21861,N_18214,N_18906);
and U21862 (N_21862,N_19245,N_17191);
nand U21863 (N_21863,N_19417,N_16495);
and U21864 (N_21864,N_18982,N_18556);
or U21865 (N_21865,N_16757,N_19120);
or U21866 (N_21866,N_15943,N_17089);
nor U21867 (N_21867,N_16692,N_19371);
nand U21868 (N_21868,N_16849,N_19029);
xor U21869 (N_21869,N_17892,N_18773);
and U21870 (N_21870,N_17040,N_19090);
nand U21871 (N_21871,N_19124,N_16587);
or U21872 (N_21872,N_16764,N_19017);
nor U21873 (N_21873,N_16346,N_19949);
nor U21874 (N_21874,N_19523,N_18164);
and U21875 (N_21875,N_18384,N_19860);
or U21876 (N_21876,N_19539,N_16706);
or U21877 (N_21877,N_15253,N_18184);
and U21878 (N_21878,N_16289,N_17827);
or U21879 (N_21879,N_18120,N_15903);
and U21880 (N_21880,N_18137,N_16093);
and U21881 (N_21881,N_19309,N_16447);
nor U21882 (N_21882,N_18007,N_15647);
and U21883 (N_21883,N_18937,N_17779);
or U21884 (N_21884,N_18665,N_16199);
and U21885 (N_21885,N_18441,N_16121);
nor U21886 (N_21886,N_15236,N_19484);
nor U21887 (N_21887,N_15789,N_15213);
and U21888 (N_21888,N_15175,N_17712);
or U21889 (N_21889,N_19030,N_18280);
and U21890 (N_21890,N_15446,N_17095);
or U21891 (N_21891,N_17789,N_15158);
and U21892 (N_21892,N_17033,N_19837);
nand U21893 (N_21893,N_19027,N_16834);
and U21894 (N_21894,N_16058,N_19240);
or U21895 (N_21895,N_16318,N_16320);
xnor U21896 (N_21896,N_15700,N_16912);
nand U21897 (N_21897,N_16250,N_15932);
nor U21898 (N_21898,N_16956,N_19023);
nor U21899 (N_21899,N_19499,N_16917);
nor U21900 (N_21900,N_15197,N_17731);
nand U21901 (N_21901,N_17082,N_16258);
xnor U21902 (N_21902,N_18489,N_15923);
and U21903 (N_21903,N_15347,N_16654);
nand U21904 (N_21904,N_16845,N_18646);
nand U21905 (N_21905,N_18639,N_16021);
and U21906 (N_21906,N_15297,N_18080);
nor U21907 (N_21907,N_19170,N_15038);
nand U21908 (N_21908,N_16205,N_19294);
or U21909 (N_21909,N_15650,N_19834);
and U21910 (N_21910,N_16015,N_19887);
xor U21911 (N_21911,N_16672,N_16175);
xnor U21912 (N_21912,N_16096,N_18585);
and U21913 (N_21913,N_18104,N_18693);
and U21914 (N_21914,N_17278,N_17946);
nor U21915 (N_21915,N_15449,N_17410);
or U21916 (N_21916,N_15728,N_17710);
and U21917 (N_21917,N_15727,N_15680);
nand U21918 (N_21918,N_17399,N_18706);
and U21919 (N_21919,N_15788,N_19794);
and U21920 (N_21920,N_19050,N_15230);
nand U21921 (N_21921,N_15057,N_19223);
nor U21922 (N_21922,N_15004,N_16168);
or U21923 (N_21923,N_16234,N_19116);
nand U21924 (N_21924,N_17318,N_19802);
and U21925 (N_21925,N_19346,N_15223);
nand U21926 (N_21926,N_18650,N_18209);
and U21927 (N_21927,N_18160,N_17426);
or U21928 (N_21928,N_16043,N_16653);
nor U21929 (N_21929,N_15599,N_16368);
nor U21930 (N_21930,N_18407,N_16360);
and U21931 (N_21931,N_17869,N_18351);
nor U21932 (N_21932,N_18419,N_16329);
and U21933 (N_21933,N_19813,N_15755);
nand U21934 (N_21934,N_18935,N_18572);
or U21935 (N_21935,N_18339,N_15419);
or U21936 (N_21936,N_17579,N_19861);
or U21937 (N_21937,N_15256,N_16136);
xor U21938 (N_21938,N_16908,N_17682);
and U21939 (N_21939,N_15925,N_18497);
and U21940 (N_21940,N_18649,N_16492);
and U21941 (N_21941,N_19436,N_19098);
and U21942 (N_21942,N_15842,N_16768);
and U21943 (N_21943,N_19840,N_17496);
nand U21944 (N_21944,N_18093,N_17164);
or U21945 (N_21945,N_17059,N_15359);
and U21946 (N_21946,N_15614,N_17000);
nor U21947 (N_21947,N_16582,N_15475);
or U21948 (N_21948,N_19505,N_19478);
nand U21949 (N_21949,N_18847,N_16551);
nand U21950 (N_21950,N_18333,N_17918);
nand U21951 (N_21951,N_15693,N_17071);
nand U21952 (N_21952,N_17800,N_18591);
and U21953 (N_21953,N_15707,N_17258);
nor U21954 (N_21954,N_18166,N_19884);
or U21955 (N_21955,N_15470,N_19841);
and U21956 (N_21956,N_19259,N_17077);
or U21957 (N_21957,N_15488,N_16954);
nand U21958 (N_21958,N_15549,N_19282);
nor U21959 (N_21959,N_17277,N_16421);
nand U21960 (N_21960,N_19509,N_19859);
and U21961 (N_21961,N_19774,N_17763);
nand U21962 (N_21962,N_19741,N_19818);
and U21963 (N_21963,N_19682,N_18140);
nor U21964 (N_21964,N_19755,N_19335);
nand U21965 (N_21965,N_15243,N_17971);
nor U21966 (N_21966,N_15821,N_16017);
and U21967 (N_21967,N_15286,N_16480);
or U21968 (N_21968,N_18459,N_17915);
and U21969 (N_21969,N_19956,N_15659);
nor U21970 (N_21970,N_18408,N_15685);
nor U21971 (N_21971,N_18350,N_18885);
nand U21972 (N_21972,N_15266,N_18003);
nor U21973 (N_21973,N_18750,N_15201);
and U21974 (N_21974,N_17824,N_17943);
and U21975 (N_21975,N_19148,N_15977);
xnor U21976 (N_21976,N_15272,N_17999);
and U21977 (N_21977,N_15986,N_19451);
and U21978 (N_21978,N_17535,N_19486);
nand U21979 (N_21979,N_18193,N_17719);
or U21980 (N_21980,N_19516,N_15144);
and U21981 (N_21981,N_19533,N_15865);
and U21982 (N_21982,N_18215,N_16712);
and U21983 (N_21983,N_16071,N_18494);
and U21984 (N_21984,N_19599,N_17593);
nor U21985 (N_21985,N_16861,N_16024);
nand U21986 (N_21986,N_17504,N_16929);
nor U21987 (N_21987,N_16987,N_19203);
and U21988 (N_21988,N_19403,N_17861);
or U21989 (N_21989,N_18189,N_17925);
nor U21990 (N_21990,N_17253,N_17264);
or U21991 (N_21991,N_15682,N_16962);
or U21992 (N_21992,N_16054,N_15454);
nor U21993 (N_21993,N_16552,N_16971);
or U21994 (N_21994,N_16127,N_17215);
nand U21995 (N_21995,N_16726,N_17356);
xnor U21996 (N_21996,N_16779,N_18889);
nand U21997 (N_21997,N_19842,N_16181);
nand U21998 (N_21998,N_19897,N_17036);
and U21999 (N_21999,N_15948,N_19004);
or U22000 (N_22000,N_17050,N_18971);
nand U22001 (N_22001,N_16562,N_17052);
and U22002 (N_22002,N_17883,N_17500);
and U22003 (N_22003,N_15997,N_15548);
nand U22004 (N_22004,N_18825,N_16206);
nor U22005 (N_22005,N_16777,N_18433);
and U22006 (N_22006,N_15854,N_18428);
and U22007 (N_22007,N_18927,N_18245);
xnor U22008 (N_22008,N_17105,N_15491);
xor U22009 (N_22009,N_17231,N_15718);
or U22010 (N_22010,N_15916,N_17364);
or U22011 (N_22011,N_18443,N_18928);
nor U22012 (N_22012,N_15841,N_17272);
or U22013 (N_22013,N_18279,N_16664);
nor U22014 (N_22014,N_16190,N_17412);
and U22015 (N_22015,N_16069,N_16108);
or U22016 (N_22016,N_15640,N_15096);
and U22017 (N_22017,N_15154,N_15574);
nor U22018 (N_22018,N_15058,N_18437);
or U22019 (N_22019,N_17758,N_19264);
or U22020 (N_22020,N_15689,N_16272);
nor U22021 (N_22021,N_18704,N_19611);
nor U22022 (N_22022,N_15000,N_16146);
nor U22023 (N_22023,N_15003,N_19483);
nand U22024 (N_22024,N_16710,N_17707);
and U22025 (N_22025,N_19475,N_16693);
nand U22026 (N_22026,N_16632,N_19705);
nor U22027 (N_22027,N_15105,N_19761);
nand U22028 (N_22028,N_17871,N_18967);
or U22029 (N_22029,N_16160,N_16196);
nand U22030 (N_22030,N_15961,N_19105);
or U22031 (N_22031,N_15736,N_15043);
nand U22032 (N_22032,N_15991,N_17782);
or U22033 (N_22033,N_17488,N_15564);
or U22034 (N_22034,N_16291,N_18124);
and U22035 (N_22035,N_18061,N_17448);
nor U22036 (N_22036,N_18097,N_18327);
nand U22037 (N_22037,N_17931,N_15466);
and U22038 (N_22038,N_17848,N_18042);
nor U22039 (N_22039,N_17813,N_19386);
nor U22040 (N_22040,N_19703,N_15623);
and U22041 (N_22041,N_18575,N_18143);
nand U22042 (N_22042,N_16125,N_15035);
nand U22043 (N_22043,N_18742,N_19986);
nand U22044 (N_22044,N_18612,N_18873);
or U22045 (N_22045,N_15536,N_15128);
or U22046 (N_22046,N_15242,N_15839);
nand U22047 (N_22047,N_15945,N_16943);
nand U22048 (N_22048,N_17385,N_17688);
nand U22049 (N_22049,N_19079,N_19410);
nand U22050 (N_22050,N_18248,N_15124);
nor U22051 (N_22051,N_16966,N_18057);
nand U22052 (N_22052,N_19372,N_18802);
or U22053 (N_22053,N_15506,N_18391);
nor U22054 (N_22054,N_18931,N_18117);
nor U22055 (N_22055,N_18260,N_16859);
or U22056 (N_22056,N_17752,N_18788);
nor U22057 (N_22057,N_17474,N_19784);
nand U22058 (N_22058,N_16195,N_18512);
nor U22059 (N_22059,N_19352,N_15500);
nand U22060 (N_22060,N_15357,N_16422);
nor U22061 (N_22061,N_18486,N_19696);
or U22062 (N_22062,N_16907,N_17079);
nor U22063 (N_22063,N_17416,N_19541);
nand U22064 (N_22064,N_17199,N_19477);
nand U22065 (N_22065,N_19528,N_18574);
nor U22066 (N_22066,N_19766,N_15396);
nor U22067 (N_22067,N_15374,N_17436);
and U22068 (N_22068,N_15835,N_19662);
or U22069 (N_22069,N_19033,N_18549);
nor U22070 (N_22070,N_16863,N_15330);
nand U22071 (N_22071,N_17809,N_18725);
or U22072 (N_22072,N_19326,N_17581);
nand U22073 (N_22073,N_19198,N_16953);
nor U22074 (N_22074,N_15257,N_17591);
nor U22075 (N_22075,N_15849,N_18606);
nand U22076 (N_22076,N_19037,N_16550);
nand U22077 (N_22077,N_16075,N_15660);
or U22078 (N_22078,N_19636,N_17885);
or U22079 (N_22079,N_15719,N_19285);
and U22080 (N_22080,N_18389,N_15170);
nand U22081 (N_22081,N_15580,N_15908);
nand U22082 (N_22082,N_17609,N_16995);
nor U22083 (N_22083,N_16062,N_19430);
xnor U22084 (N_22084,N_19862,N_19927);
nand U22085 (N_22085,N_15794,N_18689);
nor U22086 (N_22086,N_15845,N_16255);
nor U22087 (N_22087,N_19968,N_15327);
nor U22088 (N_22088,N_19723,N_16323);
nand U22089 (N_22089,N_16520,N_18330);
nand U22090 (N_22090,N_19515,N_17560);
or U22091 (N_22091,N_18059,N_16364);
nand U22092 (N_22092,N_16177,N_16044);
or U22093 (N_22093,N_18540,N_16979);
nor U22094 (N_22094,N_19482,N_15117);
or U22095 (N_22095,N_18072,N_19055);
and U22096 (N_22096,N_17048,N_19882);
xnor U22097 (N_22097,N_17543,N_15066);
nor U22098 (N_22098,N_17106,N_15240);
and U22099 (N_22099,N_17140,N_19963);
and U22100 (N_22100,N_16388,N_19378);
and U22101 (N_22101,N_17702,N_18876);
nand U22102 (N_22102,N_18113,N_16899);
and U22103 (N_22103,N_16802,N_18552);
nor U22104 (N_22104,N_15529,N_16842);
nand U22105 (N_22105,N_16256,N_15722);
nor U22106 (N_22106,N_15786,N_18205);
and U22107 (N_22107,N_17007,N_18980);
nand U22108 (N_22108,N_18207,N_19921);
and U22109 (N_22109,N_15052,N_15671);
nand U22110 (N_22110,N_17863,N_15690);
or U22111 (N_22111,N_16109,N_16938);
nor U22112 (N_22112,N_16886,N_18483);
or U22113 (N_22113,N_19188,N_18354);
and U22114 (N_22114,N_17321,N_15829);
xor U22115 (N_22115,N_15715,N_16446);
nand U22116 (N_22116,N_17411,N_18035);
or U22117 (N_22117,N_17161,N_18683);
nand U22118 (N_22118,N_16371,N_17328);
and U22119 (N_22119,N_17938,N_17384);
nand U22120 (N_22120,N_17924,N_16950);
nand U22121 (N_22121,N_18634,N_18765);
nor U22122 (N_22122,N_15525,N_15557);
nor U22123 (N_22123,N_16788,N_18102);
nand U22124 (N_22124,N_18524,N_17630);
nor U22125 (N_22125,N_15410,N_15485);
xor U22126 (N_22126,N_19363,N_18139);
or U22127 (N_22127,N_17860,N_16860);
nor U22128 (N_22128,N_17440,N_16594);
nor U22129 (N_22129,N_17958,N_19421);
or U22130 (N_22130,N_18478,N_15156);
nor U22131 (N_22131,N_19176,N_16243);
or U22132 (N_22132,N_17319,N_17171);
or U22133 (N_22133,N_15732,N_17181);
nand U22134 (N_22134,N_15202,N_19917);
nor U22135 (N_22135,N_19327,N_18151);
and U22136 (N_22136,N_15216,N_18522);
nand U22137 (N_22137,N_15462,N_15897);
nand U22138 (N_22138,N_18418,N_16898);
or U22139 (N_22139,N_16648,N_18337);
or U22140 (N_22140,N_18360,N_19300);
nor U22141 (N_22141,N_19289,N_15078);
nand U22142 (N_22142,N_15799,N_17421);
and U22143 (N_22143,N_16678,N_15168);
nand U22144 (N_22144,N_16998,N_16897);
nor U22145 (N_22145,N_16456,N_15438);
nand U22146 (N_22146,N_16581,N_19239);
nor U22147 (N_22147,N_15402,N_18499);
nand U22148 (N_22148,N_19313,N_18075);
nor U22149 (N_22149,N_16439,N_19552);
nor U22150 (N_22150,N_18648,N_16316);
or U22151 (N_22151,N_16165,N_17023);
nor U22152 (N_22152,N_16867,N_19139);
and U22153 (N_22153,N_16283,N_16082);
or U22154 (N_22154,N_16733,N_17163);
and U22155 (N_22155,N_16732,N_18566);
or U22156 (N_22156,N_16622,N_15965);
or U22157 (N_22157,N_15953,N_17912);
or U22158 (N_22158,N_19293,N_16574);
and U22159 (N_22159,N_16220,N_16791);
nor U22160 (N_22160,N_18312,N_16978);
or U22161 (N_22161,N_18295,N_16232);
xor U22162 (N_22162,N_17511,N_15046);
nor U22163 (N_22163,N_15492,N_15457);
nand U22164 (N_22164,N_15516,N_19894);
nand U22165 (N_22165,N_17798,N_17438);
nor U22166 (N_22166,N_16281,N_15423);
nand U22167 (N_22167,N_15746,N_17727);
or U22168 (N_22168,N_18050,N_16072);
nand U22169 (N_22169,N_17960,N_19095);
or U22170 (N_22170,N_18743,N_19409);
nor U22171 (N_22171,N_19302,N_15464);
xor U22172 (N_22172,N_17214,N_18769);
and U22173 (N_22173,N_15922,N_18882);
and U22174 (N_22174,N_16887,N_19128);
nor U22175 (N_22175,N_18043,N_18795);
nand U22176 (N_22176,N_19311,N_16378);
nand U22177 (N_22177,N_17765,N_15892);
and U22178 (N_22178,N_19822,N_19036);
and U22179 (N_22179,N_15116,N_18716);
or U22180 (N_22180,N_18095,N_16273);
or U22181 (N_22181,N_15868,N_17325);
nor U22182 (N_22182,N_16558,N_16990);
xor U22183 (N_22183,N_19821,N_19046);
xor U22184 (N_22184,N_17247,N_19634);
xor U22185 (N_22185,N_15770,N_16287);
nor U22186 (N_22186,N_19493,N_17741);
and U22187 (N_22187,N_15210,N_16625);
or U22188 (N_22188,N_17388,N_17873);
or U22189 (N_22189,N_18772,N_16944);
and U22190 (N_22190,N_19752,N_19643);
nand U22191 (N_22191,N_18897,N_15006);
nor U22192 (N_22192,N_15712,N_15936);
and U22193 (N_22193,N_17839,N_17334);
nand U22194 (N_22194,N_16835,N_17742);
and U22195 (N_22195,N_15351,N_15967);
and U22196 (N_22196,N_17294,N_19355);
and U22197 (N_22197,N_17595,N_17524);
nor U22198 (N_22198,N_16803,N_18558);
and U22199 (N_22199,N_17324,N_19248);
nor U22200 (N_22200,N_19844,N_17323);
xnor U22201 (N_22201,N_19086,N_19648);
or U22202 (N_22202,N_15401,N_16358);
nor U22203 (N_22203,N_15311,N_15705);
and U22204 (N_22204,N_15590,N_15331);
nand U22205 (N_22205,N_18008,N_18156);
nor U22206 (N_22206,N_16610,N_16870);
or U22207 (N_22207,N_18432,N_16937);
or U22208 (N_22208,N_18904,N_19679);
or U22209 (N_22209,N_15355,N_19666);
or U22210 (N_22210,N_15420,N_18352);
nor U22211 (N_22211,N_19186,N_15594);
or U22212 (N_22212,N_19687,N_18308);
or U22213 (N_22213,N_18297,N_15390);
or U22214 (N_22214,N_19401,N_16145);
and U22215 (N_22215,N_17618,N_16502);
or U22216 (N_22216,N_18696,N_15385);
nand U22217 (N_22217,N_19704,N_18730);
and U22218 (N_22218,N_18658,N_19870);
or U22219 (N_22219,N_16856,N_16517);
xnor U22220 (N_22220,N_19513,N_18893);
and U22221 (N_22221,N_17590,N_16202);
or U22222 (N_22222,N_19413,N_18195);
nor U22223 (N_22223,N_19898,N_19596);
xnor U22224 (N_22224,N_16169,N_17386);
or U22225 (N_22225,N_18174,N_17162);
nor U22226 (N_22226,N_17076,N_16592);
nand U22227 (N_22227,N_16742,N_17451);
and U22228 (N_22228,N_19237,N_19983);
or U22229 (N_22229,N_17835,N_16833);
nand U22230 (N_22230,N_19218,N_17259);
xor U22231 (N_22231,N_18299,N_15155);
nor U22232 (N_22232,N_18406,N_19543);
nor U22233 (N_22233,N_19359,N_17236);
or U22234 (N_22234,N_16467,N_16331);
or U22235 (N_22235,N_15087,N_15834);
nor U22236 (N_22236,N_15779,N_17221);
nor U22237 (N_22237,N_16334,N_16814);
and U22238 (N_22238,N_17642,N_19673);
or U22239 (N_22239,N_16275,N_16975);
nand U22240 (N_22240,N_17550,N_17566);
nor U22241 (N_22241,N_16449,N_18724);
and U22242 (N_22242,N_18775,N_15531);
nand U22243 (N_22243,N_18947,N_18924);
nand U22244 (N_22244,N_17358,N_19007);
xnor U22245 (N_22245,N_18940,N_18746);
nand U22246 (N_22246,N_15716,N_18253);
nand U22247 (N_22247,N_15001,N_18150);
nand U22248 (N_22248,N_15890,N_16235);
nor U22249 (N_22249,N_18806,N_15416);
nor U22250 (N_22250,N_19574,N_19135);
and U22251 (N_22251,N_17001,N_17233);
nor U22252 (N_22252,N_17631,N_16604);
nand U22253 (N_22253,N_15172,N_18371);
or U22254 (N_22254,N_18313,N_16270);
nor U22255 (N_22255,N_18135,N_19753);
or U22256 (N_22256,N_17603,N_18132);
or U22257 (N_22257,N_19593,N_15966);
nand U22258 (N_22258,N_19955,N_18858);
nor U22259 (N_22259,N_15305,N_17547);
nand U22260 (N_22260,N_17530,N_15743);
nor U22261 (N_22261,N_19001,N_19048);
nor U22262 (N_22262,N_17005,N_16752);
or U22263 (N_22263,N_15919,N_16694);
or U22264 (N_22264,N_16846,N_16295);
or U22265 (N_22265,N_15956,N_17623);
nand U22266 (N_22266,N_16402,N_19474);
or U22267 (N_22267,N_15636,N_17460);
and U22268 (N_22268,N_17396,N_18090);
nor U22269 (N_22269,N_16185,N_16307);
or U22270 (N_22270,N_17362,N_15888);
or U22271 (N_22271,N_19902,N_18877);
and U22272 (N_22272,N_17646,N_15169);
and U22273 (N_22273,N_19039,N_17062);
and U22274 (N_22274,N_16325,N_16279);
and U22275 (N_22275,N_17549,N_19609);
nand U22276 (N_22276,N_15341,N_16149);
nand U22277 (N_22277,N_18274,N_19288);
xor U22278 (N_22278,N_17914,N_17818);
nor U22279 (N_22279,N_17028,N_16812);
or U22280 (N_22280,N_19472,N_19557);
and U22281 (N_22281,N_17208,N_17038);
or U22282 (N_22282,N_15424,N_19503);
or U22283 (N_22283,N_19151,N_16382);
nand U22284 (N_22284,N_17795,N_18991);
and U22285 (N_22285,N_19973,N_18010);
or U22286 (N_22286,N_18290,N_18708);
or U22287 (N_22287,N_15280,N_18316);
xor U22288 (N_22288,N_19967,N_17745);
nand U22289 (N_22289,N_17585,N_18598);
and U22290 (N_22290,N_16002,N_15041);
nor U22291 (N_22291,N_16698,N_17563);
or U22292 (N_22292,N_19890,N_19872);
and U22293 (N_22293,N_19691,N_15909);
nand U22294 (N_22294,N_19945,N_18317);
nor U22295 (N_22295,N_19072,N_15830);
nand U22296 (N_22296,N_18396,N_19686);
or U22297 (N_22297,N_15298,N_15669);
nand U22298 (N_22298,N_18285,N_15775);
nor U22299 (N_22299,N_19161,N_18460);
and U22300 (N_22300,N_16374,N_17177);
or U22301 (N_22301,N_16878,N_16872);
nor U22302 (N_22302,N_16597,N_18521);
and U22303 (N_22303,N_17088,N_16838);
and U22304 (N_22304,N_15104,N_19224);
nand U22305 (N_22305,N_17283,N_18836);
nand U22306 (N_22306,N_16138,N_18136);
or U22307 (N_22307,N_19192,N_16894);
or U22308 (N_22308,N_19728,N_18578);
nor U22309 (N_22309,N_17439,N_15507);
nand U22310 (N_22310,N_16489,N_18694);
and U22311 (N_22311,N_15007,N_17212);
nor U22312 (N_22312,N_15287,N_16921);
nor U22313 (N_22313,N_16596,N_17112);
xnor U22314 (N_22314,N_17602,N_18256);
xnor U22315 (N_22315,N_17738,N_19764);
nor U22316 (N_22316,N_19406,N_19225);
nor U22317 (N_22317,N_18636,N_18723);
nor U22318 (N_22318,N_15773,N_16432);
nand U22319 (N_22319,N_19706,N_16348);
or U22320 (N_22320,N_17254,N_17489);
nand U22321 (N_22321,N_17615,N_19959);
and U22322 (N_22322,N_19205,N_19709);
or U22323 (N_22323,N_17692,N_18495);
xnor U22324 (N_22324,N_17757,N_19661);
nor U22325 (N_22325,N_18052,N_16473);
nand U22326 (N_22326,N_15501,N_15186);
nand U22327 (N_22327,N_16312,N_18157);
or U22328 (N_22328,N_19740,N_18020);
nand U22329 (N_22329,N_16394,N_19913);
nor U22330 (N_22330,N_19241,N_19657);
or U22331 (N_22331,N_19246,N_18846);
and U22332 (N_22332,N_18707,N_19270);
nor U22333 (N_22333,N_18204,N_18427);
nor U22334 (N_22334,N_19791,N_17492);
and U22335 (N_22335,N_18833,N_18997);
nand U22336 (N_22336,N_18674,N_17437);
nor U22337 (N_22337,N_18537,N_16687);
or U22338 (N_22338,N_19734,N_18015);
and U22339 (N_22339,N_19572,N_16864);
xnor U22340 (N_22340,N_15545,N_18287);
xnor U22341 (N_22341,N_17980,N_19582);
nand U22342 (N_22342,N_18698,N_16198);
or U22343 (N_22343,N_16501,N_16548);
and U22344 (N_22344,N_18659,N_17929);
nor U22345 (N_22345,N_17037,N_17694);
or U22346 (N_22346,N_17147,N_19408);
and U22347 (N_22347,N_16989,N_19961);
nor U22348 (N_22348,N_15570,N_18106);
and U22349 (N_22349,N_19206,N_18930);
nand U22350 (N_22350,N_19088,N_15259);
nand U22351 (N_22351,N_15246,N_16059);
nor U22352 (N_22352,N_19049,N_17015);
or U22353 (N_22353,N_18319,N_19985);
nor U22354 (N_22354,N_18995,N_18886);
nor U22355 (N_22355,N_19646,N_16858);
or U22356 (N_22356,N_15064,N_17133);
nand U22357 (N_22357,N_17246,N_18798);
or U22358 (N_22358,N_16083,N_17986);
nand U22359 (N_22359,N_16280,N_15084);
nor U22360 (N_22360,N_16677,N_19164);
or U22361 (N_22361,N_17996,N_19339);
and U22362 (N_22362,N_15630,N_17674);
or U22363 (N_22363,N_18165,N_16230);
xor U22364 (N_22364,N_16338,N_16391);
nor U22365 (N_22365,N_16607,N_19419);
and U22366 (N_22366,N_19544,N_17207);
and U22367 (N_22367,N_15795,N_18871);
nor U22368 (N_22368,N_17480,N_15322);
nand U22369 (N_22369,N_15534,N_17577);
and U22370 (N_22370,N_16385,N_18905);
nand U22371 (N_22371,N_17658,N_17976);
or U22372 (N_22372,N_16857,N_17952);
nand U22373 (N_22373,N_19290,N_15133);
nor U22374 (N_22374,N_15949,N_16188);
and U22375 (N_22375,N_17087,N_16837);
and U22376 (N_22376,N_15353,N_15237);
or U22377 (N_22377,N_16691,N_16417);
nand U22378 (N_22378,N_16418,N_16065);
nand U22379 (N_22379,N_16766,N_19504);
nand U22380 (N_22380,N_18338,N_19013);
nor U22381 (N_22381,N_18898,N_17508);
xnor U22382 (N_22382,N_17654,N_19470);
xnor U22383 (N_22383,N_16053,N_16463);
nor U22384 (N_22384,N_16992,N_18978);
nor U22385 (N_22385,N_18318,N_16608);
and U22386 (N_22386,N_16657,N_17721);
or U22387 (N_22387,N_18525,N_17974);
and U22388 (N_22388,N_16176,N_16828);
or U22389 (N_22389,N_18131,N_17531);
xor U22390 (N_22390,N_18017,N_17859);
nor U22391 (N_22391,N_16758,N_18921);
nand U22392 (N_22392,N_18488,N_15164);
and U22393 (N_22393,N_15375,N_17803);
or U22394 (N_22394,N_19617,N_15692);
or U22395 (N_22395,N_19303,N_15820);
nand U22396 (N_22396,N_16667,N_17073);
nand U22397 (N_22397,N_16078,N_19298);
or U22398 (N_22398,N_17024,N_16027);
nor U22399 (N_22399,N_16033,N_15166);
or U22400 (N_22400,N_17055,N_16717);
nor U22401 (N_22401,N_16298,N_17644);
nand U22402 (N_22402,N_17880,N_18185);
or U22403 (N_22403,N_16322,N_17201);
or U22404 (N_22404,N_16847,N_16020);
or U22405 (N_22405,N_15127,N_19871);
or U22406 (N_22406,N_18049,N_15274);
or U22407 (N_22407,N_17269,N_19003);
nand U22408 (N_22408,N_19635,N_18766);
or U22409 (N_22409,N_16565,N_18874);
or U22410 (N_22410,N_17473,N_19592);
xnor U22411 (N_22411,N_16369,N_15196);
or U22412 (N_22412,N_15626,N_19184);
or U22413 (N_22413,N_19667,N_17846);
and U22414 (N_22414,N_15369,N_19820);
nor U22415 (N_22415,N_18268,N_18477);
nand U22416 (N_22416,N_15753,N_18910);
nand U22417 (N_22417,N_18590,N_15810);
or U22418 (N_22418,N_17459,N_19432);
nand U22419 (N_22419,N_16303,N_18815);
or U22420 (N_22420,N_18038,N_17454);
and U22421 (N_22421,N_15931,N_15871);
nand U22422 (N_22422,N_15441,N_18805);
nand U22423 (N_22423,N_15915,N_16724);
xor U22424 (N_22424,N_17672,N_18323);
and U22425 (N_22425,N_19971,N_19518);
nand U22426 (N_22426,N_16084,N_16045);
nand U22427 (N_22427,N_16491,N_16583);
or U22428 (N_22428,N_17045,N_19685);
and U22429 (N_22429,N_18366,N_18111);
nor U22430 (N_22430,N_15318,N_16785);
or U22431 (N_22431,N_17773,N_18751);
nor U22432 (N_22432,N_18853,N_19060);
and U22433 (N_22433,N_15027,N_16474);
xor U22434 (N_22434,N_15054,N_17936);
nand U22435 (N_22435,N_19092,N_15039);
xnor U22436 (N_22436,N_17904,N_17649);
nand U22437 (N_22437,N_15761,N_15092);
and U22438 (N_22438,N_18631,N_17526);
nand U22439 (N_22439,N_15174,N_17552);
nand U22440 (N_22440,N_19385,N_17228);
nand U22441 (N_22441,N_19585,N_16578);
nand U22442 (N_22442,N_17450,N_17398);
and U22443 (N_22443,N_18310,N_17589);
nand U22444 (N_22444,N_18929,N_15714);
or U22445 (N_22445,N_19452,N_19199);
and U22446 (N_22446,N_17775,N_19360);
or U22447 (N_22447,N_15191,N_15733);
and U22448 (N_22448,N_19838,N_16011);
nand U22449 (N_22449,N_16972,N_17223);
xor U22450 (N_22450,N_19849,N_17882);
nand U22451 (N_22451,N_16804,N_16390);
nor U22452 (N_22452,N_16823,N_15238);
nand U22453 (N_22453,N_15894,N_16981);
and U22454 (N_22454,N_19602,N_16204);
or U22455 (N_22455,N_19982,N_15720);
and U22456 (N_22456,N_18829,N_18361);
or U22457 (N_22457,N_18147,N_17378);
or U22458 (N_22458,N_18346,N_18865);
and U22459 (N_22459,N_19292,N_16434);
nor U22460 (N_22460,N_19145,N_18690);
nor U22461 (N_22461,N_15433,N_16098);
or U22462 (N_22462,N_17002,N_17173);
or U22463 (N_22463,N_19008,N_15241);
or U22464 (N_22464,N_19561,N_15085);
or U22465 (N_22465,N_19548,N_18801);
or U22466 (N_22466,N_19500,N_15179);
or U22467 (N_22467,N_18837,N_19711);
nor U22468 (N_22468,N_17260,N_16314);
or U22469 (N_22469,N_19134,N_17890);
nor U22470 (N_22470,N_16982,N_16486);
xnor U22471 (N_22471,N_17558,N_17373);
nand U22472 (N_22472,N_16347,N_18178);
or U22473 (N_22473,N_17274,N_18568);
nand U22474 (N_22474,N_15091,N_16201);
nand U22475 (N_22475,N_18016,N_16361);
nand U22476 (N_22476,N_16885,N_17722);
xnor U22477 (N_22477,N_17061,N_16510);
or U22478 (N_22478,N_19671,N_16573);
nand U22479 (N_22479,N_19096,N_17747);
or U22480 (N_22480,N_19093,N_19522);
nor U22481 (N_22481,N_15200,N_15033);
xnor U22482 (N_22482,N_16426,N_19440);
nand U22483 (N_22483,N_17887,N_17559);
nand U22484 (N_22484,N_18170,N_19742);
nand U22485 (N_22485,N_16459,N_16801);
and U22486 (N_22486,N_19150,N_18122);
xnor U22487 (N_22487,N_19525,N_19926);
xor U22488 (N_22488,N_19078,N_19565);
xnor U22489 (N_22489,N_17479,N_17475);
or U22490 (N_22490,N_18621,N_16064);
xor U22491 (N_22491,N_19022,N_17678);
and U22492 (N_22492,N_18642,N_17449);
nand U22493 (N_22493,N_18682,N_17981);
or U22494 (N_22494,N_15653,N_15706);
nand U22495 (N_22495,N_15383,N_18832);
or U22496 (N_22496,N_16452,N_16163);
or U22497 (N_22497,N_17634,N_18891);
nand U22498 (N_22498,N_15384,N_15522);
or U22499 (N_22499,N_19354,N_19591);
nand U22500 (N_22500,N_16992,N_19169);
nor U22501 (N_22501,N_16835,N_15187);
and U22502 (N_22502,N_16192,N_15181);
nand U22503 (N_22503,N_17227,N_16721);
nand U22504 (N_22504,N_18947,N_19734);
and U22505 (N_22505,N_15548,N_15410);
nand U22506 (N_22506,N_19925,N_16464);
nand U22507 (N_22507,N_15217,N_18071);
nor U22508 (N_22508,N_17048,N_16007);
and U22509 (N_22509,N_16648,N_19646);
nand U22510 (N_22510,N_18503,N_16500);
nand U22511 (N_22511,N_15718,N_19094);
or U22512 (N_22512,N_16804,N_18004);
nor U22513 (N_22513,N_18723,N_16758);
nor U22514 (N_22514,N_15623,N_18619);
or U22515 (N_22515,N_19062,N_18347);
nor U22516 (N_22516,N_18809,N_18933);
xnor U22517 (N_22517,N_16855,N_16016);
and U22518 (N_22518,N_18656,N_19259);
xor U22519 (N_22519,N_17567,N_15444);
nand U22520 (N_22520,N_17889,N_17757);
and U22521 (N_22521,N_16305,N_17480);
nor U22522 (N_22522,N_16239,N_17732);
nor U22523 (N_22523,N_15364,N_16693);
or U22524 (N_22524,N_15979,N_15228);
nand U22525 (N_22525,N_16204,N_18892);
and U22526 (N_22526,N_19972,N_19564);
xor U22527 (N_22527,N_17971,N_19390);
and U22528 (N_22528,N_19744,N_16094);
or U22529 (N_22529,N_16803,N_19148);
or U22530 (N_22530,N_18973,N_15941);
nor U22531 (N_22531,N_18131,N_16874);
and U22532 (N_22532,N_15671,N_15097);
and U22533 (N_22533,N_16730,N_18564);
xor U22534 (N_22534,N_15962,N_17851);
nand U22535 (N_22535,N_17463,N_17999);
or U22536 (N_22536,N_15249,N_16072);
nand U22537 (N_22537,N_16361,N_19752);
or U22538 (N_22538,N_18507,N_16470);
nor U22539 (N_22539,N_16141,N_18146);
nand U22540 (N_22540,N_15122,N_19877);
xor U22541 (N_22541,N_17257,N_18939);
nand U22542 (N_22542,N_18631,N_17361);
or U22543 (N_22543,N_16812,N_18108);
xnor U22544 (N_22544,N_15707,N_15588);
nand U22545 (N_22545,N_19933,N_19113);
nand U22546 (N_22546,N_19953,N_16932);
xor U22547 (N_22547,N_15313,N_18221);
nor U22548 (N_22548,N_17338,N_18726);
nor U22549 (N_22549,N_19642,N_19074);
and U22550 (N_22550,N_19442,N_19639);
xnor U22551 (N_22551,N_19832,N_15687);
or U22552 (N_22552,N_15156,N_18059);
and U22553 (N_22553,N_15074,N_15283);
nand U22554 (N_22554,N_19098,N_19819);
nand U22555 (N_22555,N_18886,N_15221);
nor U22556 (N_22556,N_19156,N_17052);
nand U22557 (N_22557,N_16879,N_15019);
and U22558 (N_22558,N_16941,N_16113);
or U22559 (N_22559,N_15147,N_18380);
or U22560 (N_22560,N_16572,N_17204);
or U22561 (N_22561,N_17479,N_19463);
nor U22562 (N_22562,N_19452,N_15735);
or U22563 (N_22563,N_18456,N_18887);
and U22564 (N_22564,N_18137,N_16358);
and U22565 (N_22565,N_19610,N_17175);
nor U22566 (N_22566,N_16496,N_19033);
and U22567 (N_22567,N_17538,N_18020);
xor U22568 (N_22568,N_16912,N_18815);
xor U22569 (N_22569,N_18146,N_18800);
nor U22570 (N_22570,N_17052,N_17394);
or U22571 (N_22571,N_19830,N_19473);
or U22572 (N_22572,N_16857,N_17134);
and U22573 (N_22573,N_15502,N_15724);
and U22574 (N_22574,N_18781,N_16009);
or U22575 (N_22575,N_17791,N_18211);
and U22576 (N_22576,N_19866,N_16988);
nand U22577 (N_22577,N_16938,N_15148);
or U22578 (N_22578,N_15924,N_16641);
nand U22579 (N_22579,N_18544,N_18923);
and U22580 (N_22580,N_16528,N_16831);
nor U22581 (N_22581,N_16504,N_19250);
nor U22582 (N_22582,N_18117,N_15145);
nand U22583 (N_22583,N_15059,N_17955);
and U22584 (N_22584,N_19582,N_17283);
nor U22585 (N_22585,N_15383,N_16090);
or U22586 (N_22586,N_17095,N_17125);
nor U22587 (N_22587,N_15374,N_19639);
nor U22588 (N_22588,N_16985,N_16302);
nand U22589 (N_22589,N_17804,N_19695);
xnor U22590 (N_22590,N_17701,N_17271);
nor U22591 (N_22591,N_17044,N_18022);
and U22592 (N_22592,N_15770,N_16544);
nand U22593 (N_22593,N_15115,N_16816);
nor U22594 (N_22594,N_16213,N_17860);
nand U22595 (N_22595,N_16885,N_15759);
nand U22596 (N_22596,N_19458,N_17265);
or U22597 (N_22597,N_19258,N_16813);
and U22598 (N_22598,N_16811,N_15335);
nor U22599 (N_22599,N_16833,N_15139);
nand U22600 (N_22600,N_15634,N_16189);
and U22601 (N_22601,N_19403,N_17996);
or U22602 (N_22602,N_17730,N_17473);
nand U22603 (N_22603,N_16170,N_15161);
nand U22604 (N_22604,N_18675,N_18185);
xnor U22605 (N_22605,N_15554,N_17365);
nand U22606 (N_22606,N_19094,N_17021);
or U22607 (N_22607,N_16487,N_16631);
and U22608 (N_22608,N_18093,N_19058);
xnor U22609 (N_22609,N_16562,N_15868);
nor U22610 (N_22610,N_15901,N_16820);
or U22611 (N_22611,N_17788,N_15823);
or U22612 (N_22612,N_16234,N_16179);
nor U22613 (N_22613,N_15096,N_18981);
nor U22614 (N_22614,N_16947,N_18744);
nor U22615 (N_22615,N_18886,N_17188);
nor U22616 (N_22616,N_15598,N_19016);
and U22617 (N_22617,N_16669,N_15321);
nand U22618 (N_22618,N_17790,N_17179);
or U22619 (N_22619,N_18271,N_16967);
nor U22620 (N_22620,N_19723,N_17535);
nor U22621 (N_22621,N_15032,N_18347);
nor U22622 (N_22622,N_17610,N_19243);
and U22623 (N_22623,N_15540,N_18621);
xor U22624 (N_22624,N_16775,N_17313);
nor U22625 (N_22625,N_19132,N_16500);
and U22626 (N_22626,N_18141,N_16075);
or U22627 (N_22627,N_15414,N_17861);
or U22628 (N_22628,N_18153,N_19690);
nor U22629 (N_22629,N_16704,N_18988);
and U22630 (N_22630,N_18899,N_16392);
nand U22631 (N_22631,N_19144,N_18206);
and U22632 (N_22632,N_17289,N_16031);
xor U22633 (N_22633,N_19220,N_16263);
nor U22634 (N_22634,N_16061,N_17666);
and U22635 (N_22635,N_17828,N_15938);
or U22636 (N_22636,N_19244,N_19283);
nand U22637 (N_22637,N_16353,N_19557);
xnor U22638 (N_22638,N_15556,N_18505);
and U22639 (N_22639,N_19587,N_19475);
xor U22640 (N_22640,N_18251,N_19948);
nand U22641 (N_22641,N_18642,N_18762);
and U22642 (N_22642,N_15307,N_15704);
or U22643 (N_22643,N_19253,N_18563);
nand U22644 (N_22644,N_18300,N_16884);
or U22645 (N_22645,N_17923,N_16674);
nor U22646 (N_22646,N_19397,N_17315);
or U22647 (N_22647,N_18457,N_19519);
or U22648 (N_22648,N_18334,N_17849);
and U22649 (N_22649,N_18431,N_18088);
nor U22650 (N_22650,N_19982,N_18327);
nand U22651 (N_22651,N_18738,N_15885);
nand U22652 (N_22652,N_17129,N_16386);
nor U22653 (N_22653,N_19577,N_19949);
and U22654 (N_22654,N_19341,N_19116);
and U22655 (N_22655,N_15203,N_18002);
or U22656 (N_22656,N_18459,N_19209);
nand U22657 (N_22657,N_17946,N_16643);
or U22658 (N_22658,N_17446,N_19853);
nand U22659 (N_22659,N_16089,N_17873);
and U22660 (N_22660,N_16788,N_19004);
nor U22661 (N_22661,N_16211,N_17489);
nand U22662 (N_22662,N_18660,N_15436);
nor U22663 (N_22663,N_15022,N_15370);
nand U22664 (N_22664,N_15704,N_15310);
or U22665 (N_22665,N_18965,N_15946);
or U22666 (N_22666,N_19595,N_16811);
or U22667 (N_22667,N_15320,N_16923);
nor U22668 (N_22668,N_18379,N_15128);
and U22669 (N_22669,N_15217,N_17566);
xnor U22670 (N_22670,N_15884,N_15648);
or U22671 (N_22671,N_18536,N_15937);
or U22672 (N_22672,N_17844,N_17914);
nand U22673 (N_22673,N_17952,N_15385);
and U22674 (N_22674,N_16418,N_18560);
nor U22675 (N_22675,N_17840,N_17783);
and U22676 (N_22676,N_17632,N_19986);
and U22677 (N_22677,N_16778,N_17373);
and U22678 (N_22678,N_18612,N_16163);
nand U22679 (N_22679,N_16834,N_15657);
nand U22680 (N_22680,N_18870,N_17847);
and U22681 (N_22681,N_15457,N_19060);
xnor U22682 (N_22682,N_18607,N_15981);
nand U22683 (N_22683,N_19334,N_17463);
and U22684 (N_22684,N_18436,N_16233);
nor U22685 (N_22685,N_15974,N_19259);
nor U22686 (N_22686,N_19627,N_17273);
or U22687 (N_22687,N_17756,N_15722);
nand U22688 (N_22688,N_19712,N_16984);
nor U22689 (N_22689,N_17158,N_18504);
nor U22690 (N_22690,N_17093,N_17866);
and U22691 (N_22691,N_19855,N_15191);
and U22692 (N_22692,N_18844,N_15196);
nor U22693 (N_22693,N_15502,N_17453);
and U22694 (N_22694,N_15468,N_17248);
or U22695 (N_22695,N_17270,N_19629);
nand U22696 (N_22696,N_15316,N_16858);
nand U22697 (N_22697,N_17670,N_18015);
nor U22698 (N_22698,N_17060,N_15861);
nor U22699 (N_22699,N_17165,N_16065);
nand U22700 (N_22700,N_18474,N_15290);
and U22701 (N_22701,N_19701,N_16749);
nand U22702 (N_22702,N_15138,N_16185);
and U22703 (N_22703,N_15262,N_15895);
nand U22704 (N_22704,N_17820,N_16896);
or U22705 (N_22705,N_18895,N_16577);
nor U22706 (N_22706,N_15903,N_16846);
and U22707 (N_22707,N_15124,N_17986);
nand U22708 (N_22708,N_19523,N_19013);
and U22709 (N_22709,N_17145,N_16165);
nor U22710 (N_22710,N_19892,N_19140);
nand U22711 (N_22711,N_19012,N_16374);
or U22712 (N_22712,N_18801,N_18177);
nor U22713 (N_22713,N_19047,N_15276);
nand U22714 (N_22714,N_19752,N_18795);
nor U22715 (N_22715,N_17393,N_15735);
nor U22716 (N_22716,N_16518,N_18699);
nand U22717 (N_22717,N_18377,N_19469);
nor U22718 (N_22718,N_17500,N_19738);
and U22719 (N_22719,N_16933,N_18201);
nor U22720 (N_22720,N_15525,N_19663);
nor U22721 (N_22721,N_17913,N_17898);
nor U22722 (N_22722,N_19098,N_17766);
nand U22723 (N_22723,N_18105,N_18519);
nor U22724 (N_22724,N_15973,N_18380);
nor U22725 (N_22725,N_15053,N_15556);
nand U22726 (N_22726,N_17366,N_15212);
or U22727 (N_22727,N_17089,N_15905);
nor U22728 (N_22728,N_18499,N_19920);
and U22729 (N_22729,N_18983,N_18536);
and U22730 (N_22730,N_15604,N_15515);
and U22731 (N_22731,N_18848,N_17552);
or U22732 (N_22732,N_17512,N_18116);
and U22733 (N_22733,N_17224,N_17787);
or U22734 (N_22734,N_16399,N_17849);
and U22735 (N_22735,N_15050,N_16999);
and U22736 (N_22736,N_16060,N_19863);
xor U22737 (N_22737,N_15630,N_16920);
nand U22738 (N_22738,N_15599,N_19657);
or U22739 (N_22739,N_18175,N_18904);
or U22740 (N_22740,N_18744,N_19081);
nor U22741 (N_22741,N_15735,N_16074);
or U22742 (N_22742,N_19356,N_15373);
nor U22743 (N_22743,N_17289,N_17177);
or U22744 (N_22744,N_15390,N_16178);
nor U22745 (N_22745,N_18988,N_17557);
xor U22746 (N_22746,N_16269,N_17306);
xor U22747 (N_22747,N_15760,N_15965);
or U22748 (N_22748,N_18043,N_19156);
nand U22749 (N_22749,N_17339,N_16801);
and U22750 (N_22750,N_19639,N_19347);
nor U22751 (N_22751,N_19280,N_16774);
nand U22752 (N_22752,N_18192,N_18115);
nor U22753 (N_22753,N_18759,N_15153);
nor U22754 (N_22754,N_15523,N_15374);
nand U22755 (N_22755,N_15444,N_19376);
nor U22756 (N_22756,N_18690,N_19657);
nor U22757 (N_22757,N_15511,N_19295);
or U22758 (N_22758,N_17242,N_16349);
xnor U22759 (N_22759,N_15535,N_16750);
nand U22760 (N_22760,N_19287,N_15901);
xor U22761 (N_22761,N_15089,N_16344);
or U22762 (N_22762,N_18164,N_19916);
or U22763 (N_22763,N_18398,N_17180);
xor U22764 (N_22764,N_18981,N_17278);
nor U22765 (N_22765,N_15760,N_19340);
xor U22766 (N_22766,N_15439,N_18294);
or U22767 (N_22767,N_18771,N_16141);
xnor U22768 (N_22768,N_19540,N_19637);
nor U22769 (N_22769,N_19773,N_15326);
or U22770 (N_22770,N_17892,N_19615);
or U22771 (N_22771,N_18084,N_18952);
nand U22772 (N_22772,N_15939,N_19510);
nor U22773 (N_22773,N_19220,N_19652);
or U22774 (N_22774,N_17828,N_17273);
xnor U22775 (N_22775,N_19413,N_16487);
nor U22776 (N_22776,N_19978,N_15915);
xor U22777 (N_22777,N_16564,N_16178);
nand U22778 (N_22778,N_15234,N_18241);
or U22779 (N_22779,N_18335,N_15882);
nand U22780 (N_22780,N_17633,N_17732);
and U22781 (N_22781,N_18449,N_15487);
nand U22782 (N_22782,N_19025,N_18759);
nor U22783 (N_22783,N_18986,N_18172);
nand U22784 (N_22784,N_17230,N_16424);
or U22785 (N_22785,N_19023,N_19292);
nor U22786 (N_22786,N_18710,N_19501);
or U22787 (N_22787,N_17686,N_18587);
or U22788 (N_22788,N_16302,N_15055);
nor U22789 (N_22789,N_15643,N_19722);
and U22790 (N_22790,N_16562,N_19101);
and U22791 (N_22791,N_16178,N_16452);
nor U22792 (N_22792,N_15049,N_15488);
nor U22793 (N_22793,N_19002,N_18617);
and U22794 (N_22794,N_15697,N_18098);
or U22795 (N_22795,N_19177,N_17360);
and U22796 (N_22796,N_15714,N_18456);
nor U22797 (N_22797,N_17456,N_19465);
xor U22798 (N_22798,N_19199,N_19174);
nand U22799 (N_22799,N_18714,N_16593);
nand U22800 (N_22800,N_16208,N_15671);
nor U22801 (N_22801,N_18795,N_15981);
and U22802 (N_22802,N_19583,N_19809);
nor U22803 (N_22803,N_19212,N_17335);
nand U22804 (N_22804,N_15858,N_15025);
nor U22805 (N_22805,N_17933,N_19472);
and U22806 (N_22806,N_19139,N_17678);
and U22807 (N_22807,N_17479,N_19952);
and U22808 (N_22808,N_19315,N_17367);
and U22809 (N_22809,N_18463,N_18739);
nand U22810 (N_22810,N_15028,N_19515);
or U22811 (N_22811,N_18852,N_15431);
nor U22812 (N_22812,N_19317,N_16500);
xor U22813 (N_22813,N_16153,N_19774);
and U22814 (N_22814,N_15316,N_17807);
and U22815 (N_22815,N_19676,N_15155);
xor U22816 (N_22816,N_16747,N_17775);
nand U22817 (N_22817,N_19451,N_19774);
or U22818 (N_22818,N_18288,N_15201);
or U22819 (N_22819,N_19560,N_18874);
xnor U22820 (N_22820,N_16611,N_17510);
nor U22821 (N_22821,N_16336,N_18654);
and U22822 (N_22822,N_16002,N_16851);
or U22823 (N_22823,N_16835,N_15017);
and U22824 (N_22824,N_19409,N_16301);
nor U22825 (N_22825,N_18030,N_16145);
nand U22826 (N_22826,N_17524,N_18880);
and U22827 (N_22827,N_16169,N_18485);
nor U22828 (N_22828,N_17516,N_16672);
xnor U22829 (N_22829,N_17810,N_18463);
xnor U22830 (N_22830,N_18965,N_15470);
nor U22831 (N_22831,N_18352,N_15373);
xor U22832 (N_22832,N_15840,N_19530);
or U22833 (N_22833,N_15336,N_17627);
nor U22834 (N_22834,N_16039,N_16104);
or U22835 (N_22835,N_16559,N_19344);
nand U22836 (N_22836,N_17022,N_16924);
nand U22837 (N_22837,N_16792,N_15361);
xnor U22838 (N_22838,N_16722,N_17968);
nor U22839 (N_22839,N_15982,N_15260);
or U22840 (N_22840,N_17802,N_16026);
xnor U22841 (N_22841,N_17370,N_17610);
nor U22842 (N_22842,N_18166,N_18599);
nand U22843 (N_22843,N_18559,N_16938);
nand U22844 (N_22844,N_19932,N_17640);
and U22845 (N_22845,N_18980,N_18290);
nor U22846 (N_22846,N_18252,N_19578);
nand U22847 (N_22847,N_15827,N_17789);
nor U22848 (N_22848,N_17373,N_19725);
nor U22849 (N_22849,N_15687,N_17030);
nand U22850 (N_22850,N_17458,N_16190);
or U22851 (N_22851,N_15411,N_15527);
xor U22852 (N_22852,N_19757,N_15778);
nand U22853 (N_22853,N_19679,N_16068);
or U22854 (N_22854,N_19414,N_17377);
and U22855 (N_22855,N_17718,N_17394);
and U22856 (N_22856,N_15921,N_19623);
xor U22857 (N_22857,N_16668,N_17059);
and U22858 (N_22858,N_15326,N_18746);
or U22859 (N_22859,N_19322,N_18802);
xnor U22860 (N_22860,N_15650,N_16876);
nand U22861 (N_22861,N_16430,N_19794);
nand U22862 (N_22862,N_16931,N_18583);
xor U22863 (N_22863,N_19858,N_16728);
xnor U22864 (N_22864,N_17394,N_15823);
nor U22865 (N_22865,N_17061,N_18653);
and U22866 (N_22866,N_18017,N_16656);
xor U22867 (N_22867,N_18468,N_15006);
xor U22868 (N_22868,N_19680,N_17070);
xor U22869 (N_22869,N_15368,N_18182);
xnor U22870 (N_22870,N_17267,N_15583);
nand U22871 (N_22871,N_16602,N_16311);
and U22872 (N_22872,N_18657,N_16001);
nand U22873 (N_22873,N_19352,N_19660);
nor U22874 (N_22874,N_16054,N_19006);
nand U22875 (N_22875,N_17347,N_16930);
or U22876 (N_22876,N_16771,N_19639);
nor U22877 (N_22877,N_19906,N_16016);
nor U22878 (N_22878,N_17980,N_17736);
nand U22879 (N_22879,N_15723,N_16398);
nor U22880 (N_22880,N_18711,N_15352);
nor U22881 (N_22881,N_18747,N_17727);
and U22882 (N_22882,N_19443,N_18936);
and U22883 (N_22883,N_18159,N_17358);
or U22884 (N_22884,N_16311,N_19450);
xnor U22885 (N_22885,N_17968,N_18086);
nand U22886 (N_22886,N_18010,N_16226);
and U22887 (N_22887,N_17643,N_18118);
nor U22888 (N_22888,N_17415,N_19934);
nand U22889 (N_22889,N_16514,N_16280);
and U22890 (N_22890,N_15881,N_16047);
or U22891 (N_22891,N_19992,N_19957);
or U22892 (N_22892,N_19449,N_17429);
xor U22893 (N_22893,N_19753,N_18936);
nor U22894 (N_22894,N_15683,N_16017);
nor U22895 (N_22895,N_18457,N_18204);
or U22896 (N_22896,N_19560,N_15800);
nand U22897 (N_22897,N_19020,N_16440);
nor U22898 (N_22898,N_16518,N_15468);
or U22899 (N_22899,N_15329,N_17843);
xnor U22900 (N_22900,N_18430,N_17730);
xor U22901 (N_22901,N_16017,N_18832);
xnor U22902 (N_22902,N_16466,N_15858);
nand U22903 (N_22903,N_17992,N_16596);
and U22904 (N_22904,N_17355,N_15974);
and U22905 (N_22905,N_15361,N_18093);
nand U22906 (N_22906,N_18336,N_15596);
nor U22907 (N_22907,N_15727,N_19945);
nor U22908 (N_22908,N_17709,N_17476);
nor U22909 (N_22909,N_16993,N_15279);
and U22910 (N_22910,N_17114,N_19816);
nand U22911 (N_22911,N_19683,N_16501);
and U22912 (N_22912,N_19387,N_15824);
and U22913 (N_22913,N_15722,N_15485);
and U22914 (N_22914,N_17005,N_16855);
or U22915 (N_22915,N_16164,N_18451);
nor U22916 (N_22916,N_18419,N_15991);
nor U22917 (N_22917,N_15235,N_19414);
nand U22918 (N_22918,N_17198,N_18726);
and U22919 (N_22919,N_18252,N_19198);
xor U22920 (N_22920,N_19276,N_19178);
or U22921 (N_22921,N_17919,N_15629);
and U22922 (N_22922,N_19526,N_16201);
nor U22923 (N_22923,N_16283,N_16439);
and U22924 (N_22924,N_15731,N_15311);
or U22925 (N_22925,N_15692,N_18834);
or U22926 (N_22926,N_16180,N_17574);
and U22927 (N_22927,N_15815,N_17631);
xor U22928 (N_22928,N_16436,N_15012);
nor U22929 (N_22929,N_18192,N_17254);
nand U22930 (N_22930,N_15445,N_16388);
nand U22931 (N_22931,N_19798,N_18894);
and U22932 (N_22932,N_18952,N_16687);
nand U22933 (N_22933,N_19025,N_15165);
or U22934 (N_22934,N_16390,N_19199);
nor U22935 (N_22935,N_15283,N_19185);
nand U22936 (N_22936,N_16030,N_16039);
and U22937 (N_22937,N_16508,N_18555);
nor U22938 (N_22938,N_17296,N_15410);
nor U22939 (N_22939,N_17154,N_15478);
and U22940 (N_22940,N_19762,N_15010);
and U22941 (N_22941,N_17328,N_17772);
nand U22942 (N_22942,N_18729,N_18546);
or U22943 (N_22943,N_17337,N_19926);
nor U22944 (N_22944,N_15690,N_15146);
and U22945 (N_22945,N_18027,N_16314);
and U22946 (N_22946,N_17461,N_19551);
and U22947 (N_22947,N_18146,N_19576);
and U22948 (N_22948,N_19233,N_15802);
nor U22949 (N_22949,N_16417,N_15709);
nand U22950 (N_22950,N_19152,N_19272);
nor U22951 (N_22951,N_15806,N_17497);
and U22952 (N_22952,N_19672,N_15565);
nor U22953 (N_22953,N_16702,N_19955);
and U22954 (N_22954,N_18702,N_15752);
and U22955 (N_22955,N_16708,N_15050);
nand U22956 (N_22956,N_19177,N_16688);
and U22957 (N_22957,N_19624,N_16655);
nor U22958 (N_22958,N_15885,N_19417);
xnor U22959 (N_22959,N_15990,N_18404);
nand U22960 (N_22960,N_17097,N_19449);
nor U22961 (N_22961,N_16282,N_17746);
or U22962 (N_22962,N_15103,N_17106);
or U22963 (N_22963,N_15590,N_17783);
and U22964 (N_22964,N_19160,N_16024);
and U22965 (N_22965,N_17479,N_17466);
nor U22966 (N_22966,N_19940,N_17423);
nand U22967 (N_22967,N_16317,N_18384);
nand U22968 (N_22968,N_17520,N_16124);
or U22969 (N_22969,N_19160,N_17300);
nor U22970 (N_22970,N_19373,N_18566);
nand U22971 (N_22971,N_16011,N_18696);
nor U22972 (N_22972,N_15772,N_16705);
and U22973 (N_22973,N_17202,N_15990);
nand U22974 (N_22974,N_18965,N_17247);
nor U22975 (N_22975,N_15653,N_19076);
nor U22976 (N_22976,N_19799,N_15591);
xnor U22977 (N_22977,N_18889,N_15316);
or U22978 (N_22978,N_18458,N_17482);
or U22979 (N_22979,N_16033,N_18504);
nor U22980 (N_22980,N_17368,N_16456);
and U22981 (N_22981,N_19224,N_17733);
nand U22982 (N_22982,N_19354,N_15236);
nand U22983 (N_22983,N_16242,N_15872);
or U22984 (N_22984,N_18057,N_16054);
and U22985 (N_22985,N_16419,N_16904);
xor U22986 (N_22986,N_18650,N_17499);
nor U22987 (N_22987,N_18600,N_15395);
xor U22988 (N_22988,N_18486,N_19052);
and U22989 (N_22989,N_16522,N_15542);
xor U22990 (N_22990,N_15541,N_17536);
and U22991 (N_22991,N_15188,N_17167);
and U22992 (N_22992,N_15883,N_17881);
and U22993 (N_22993,N_17408,N_19633);
or U22994 (N_22994,N_19757,N_18394);
nand U22995 (N_22995,N_15053,N_17128);
or U22996 (N_22996,N_18874,N_19205);
nand U22997 (N_22997,N_17621,N_17493);
nor U22998 (N_22998,N_18021,N_16684);
and U22999 (N_22999,N_15211,N_15385);
and U23000 (N_23000,N_19737,N_15679);
nor U23001 (N_23001,N_15570,N_17670);
and U23002 (N_23002,N_15344,N_18966);
nand U23003 (N_23003,N_17828,N_15314);
nand U23004 (N_23004,N_19431,N_17026);
nor U23005 (N_23005,N_19546,N_15107);
nand U23006 (N_23006,N_15347,N_18463);
or U23007 (N_23007,N_16942,N_17676);
and U23008 (N_23008,N_18499,N_15861);
nor U23009 (N_23009,N_17318,N_17242);
or U23010 (N_23010,N_19433,N_18878);
nor U23011 (N_23011,N_15643,N_18930);
nor U23012 (N_23012,N_15901,N_15510);
nor U23013 (N_23013,N_19946,N_16295);
or U23014 (N_23014,N_19522,N_19460);
and U23015 (N_23015,N_17812,N_16016);
nor U23016 (N_23016,N_17272,N_17908);
or U23017 (N_23017,N_19038,N_15516);
and U23018 (N_23018,N_18032,N_18152);
nand U23019 (N_23019,N_19706,N_15385);
and U23020 (N_23020,N_16836,N_16175);
nand U23021 (N_23021,N_17085,N_16462);
nand U23022 (N_23022,N_17857,N_18617);
or U23023 (N_23023,N_15244,N_17686);
nand U23024 (N_23024,N_19148,N_17432);
nor U23025 (N_23025,N_15277,N_16891);
or U23026 (N_23026,N_17355,N_19540);
and U23027 (N_23027,N_18631,N_15866);
or U23028 (N_23028,N_18370,N_17847);
and U23029 (N_23029,N_15007,N_16612);
and U23030 (N_23030,N_16410,N_18704);
or U23031 (N_23031,N_19743,N_18941);
or U23032 (N_23032,N_19520,N_15934);
or U23033 (N_23033,N_15065,N_18592);
nand U23034 (N_23034,N_15790,N_18120);
nand U23035 (N_23035,N_15350,N_17163);
or U23036 (N_23036,N_19667,N_18446);
and U23037 (N_23037,N_16965,N_15657);
nand U23038 (N_23038,N_19242,N_19158);
nor U23039 (N_23039,N_18196,N_18786);
or U23040 (N_23040,N_19291,N_18963);
nor U23041 (N_23041,N_18698,N_19901);
nand U23042 (N_23042,N_17916,N_18013);
nor U23043 (N_23043,N_16653,N_15862);
and U23044 (N_23044,N_18280,N_15401);
or U23045 (N_23045,N_18612,N_17710);
xnor U23046 (N_23046,N_18431,N_18770);
nand U23047 (N_23047,N_16796,N_15542);
and U23048 (N_23048,N_17010,N_18947);
nand U23049 (N_23049,N_18402,N_19906);
nand U23050 (N_23050,N_17281,N_17241);
and U23051 (N_23051,N_17816,N_18732);
xor U23052 (N_23052,N_16743,N_16992);
nor U23053 (N_23053,N_16307,N_17110);
nand U23054 (N_23054,N_18675,N_18552);
and U23055 (N_23055,N_16869,N_16295);
and U23056 (N_23056,N_18683,N_16609);
xnor U23057 (N_23057,N_19352,N_19351);
nand U23058 (N_23058,N_18678,N_16285);
nor U23059 (N_23059,N_16269,N_17090);
or U23060 (N_23060,N_17788,N_15376);
xor U23061 (N_23061,N_18268,N_17151);
and U23062 (N_23062,N_19328,N_15588);
or U23063 (N_23063,N_16450,N_17667);
and U23064 (N_23064,N_15051,N_18305);
nand U23065 (N_23065,N_16708,N_19923);
or U23066 (N_23066,N_19793,N_18894);
and U23067 (N_23067,N_17889,N_16253);
nand U23068 (N_23068,N_18957,N_18490);
nand U23069 (N_23069,N_17935,N_16802);
nand U23070 (N_23070,N_15820,N_19924);
nor U23071 (N_23071,N_17040,N_16127);
and U23072 (N_23072,N_17260,N_17664);
or U23073 (N_23073,N_19496,N_18736);
and U23074 (N_23074,N_19803,N_16099);
or U23075 (N_23075,N_15455,N_19519);
nand U23076 (N_23076,N_16433,N_17727);
and U23077 (N_23077,N_19854,N_19254);
nor U23078 (N_23078,N_18112,N_17095);
or U23079 (N_23079,N_19845,N_16017);
or U23080 (N_23080,N_19553,N_19232);
nor U23081 (N_23081,N_16615,N_18380);
or U23082 (N_23082,N_15416,N_18203);
xnor U23083 (N_23083,N_16318,N_18683);
nor U23084 (N_23084,N_16401,N_18317);
or U23085 (N_23085,N_15878,N_15522);
or U23086 (N_23086,N_16389,N_15283);
xor U23087 (N_23087,N_17615,N_15233);
nor U23088 (N_23088,N_18894,N_17860);
nor U23089 (N_23089,N_16866,N_17860);
or U23090 (N_23090,N_16837,N_17139);
or U23091 (N_23091,N_17160,N_15825);
or U23092 (N_23092,N_18545,N_15805);
nor U23093 (N_23093,N_18770,N_18628);
nor U23094 (N_23094,N_17149,N_19883);
nor U23095 (N_23095,N_18835,N_17717);
nand U23096 (N_23096,N_15182,N_18661);
and U23097 (N_23097,N_18608,N_17299);
and U23098 (N_23098,N_18414,N_19982);
and U23099 (N_23099,N_19912,N_17754);
or U23100 (N_23100,N_19057,N_19115);
nand U23101 (N_23101,N_19534,N_17602);
or U23102 (N_23102,N_16899,N_17209);
nor U23103 (N_23103,N_18401,N_19426);
or U23104 (N_23104,N_18914,N_16455);
nor U23105 (N_23105,N_17740,N_17810);
and U23106 (N_23106,N_19109,N_15476);
and U23107 (N_23107,N_17598,N_15262);
nand U23108 (N_23108,N_19171,N_19858);
or U23109 (N_23109,N_15592,N_19281);
nor U23110 (N_23110,N_19041,N_15989);
nand U23111 (N_23111,N_17393,N_18158);
and U23112 (N_23112,N_16204,N_15454);
and U23113 (N_23113,N_16915,N_17079);
nor U23114 (N_23114,N_16961,N_19710);
nor U23115 (N_23115,N_16589,N_15719);
nor U23116 (N_23116,N_16771,N_15034);
nand U23117 (N_23117,N_19392,N_17513);
and U23118 (N_23118,N_19519,N_16825);
or U23119 (N_23119,N_17338,N_15327);
nand U23120 (N_23120,N_16537,N_18291);
xor U23121 (N_23121,N_19967,N_16467);
xnor U23122 (N_23122,N_19162,N_18408);
and U23123 (N_23123,N_17311,N_15513);
nand U23124 (N_23124,N_19156,N_17329);
or U23125 (N_23125,N_17530,N_18461);
nand U23126 (N_23126,N_19366,N_16987);
or U23127 (N_23127,N_15404,N_18998);
and U23128 (N_23128,N_17906,N_16601);
nand U23129 (N_23129,N_17331,N_15541);
nand U23130 (N_23130,N_16289,N_15558);
nor U23131 (N_23131,N_17786,N_15822);
or U23132 (N_23132,N_16432,N_16376);
and U23133 (N_23133,N_15817,N_17365);
nor U23134 (N_23134,N_19657,N_18642);
or U23135 (N_23135,N_16384,N_15917);
nor U23136 (N_23136,N_19087,N_17640);
xnor U23137 (N_23137,N_18901,N_18971);
nor U23138 (N_23138,N_15533,N_18017);
nand U23139 (N_23139,N_17701,N_15800);
xnor U23140 (N_23140,N_16401,N_16873);
nor U23141 (N_23141,N_17282,N_16315);
and U23142 (N_23142,N_19322,N_18260);
nor U23143 (N_23143,N_15442,N_15466);
and U23144 (N_23144,N_16070,N_19115);
nand U23145 (N_23145,N_19491,N_16455);
nand U23146 (N_23146,N_18460,N_15898);
or U23147 (N_23147,N_15801,N_15471);
and U23148 (N_23148,N_17726,N_16875);
nor U23149 (N_23149,N_18891,N_16559);
nor U23150 (N_23150,N_18761,N_19132);
and U23151 (N_23151,N_16169,N_16382);
nand U23152 (N_23152,N_17810,N_16128);
or U23153 (N_23153,N_19284,N_15210);
nand U23154 (N_23154,N_15126,N_17126);
or U23155 (N_23155,N_18803,N_16354);
xor U23156 (N_23156,N_16812,N_18145);
and U23157 (N_23157,N_17359,N_15330);
nor U23158 (N_23158,N_16761,N_15009);
nor U23159 (N_23159,N_15479,N_19123);
and U23160 (N_23160,N_18662,N_16651);
xnor U23161 (N_23161,N_18804,N_19957);
nor U23162 (N_23162,N_15291,N_17574);
nand U23163 (N_23163,N_16105,N_16513);
and U23164 (N_23164,N_17423,N_19788);
or U23165 (N_23165,N_18372,N_15359);
or U23166 (N_23166,N_19162,N_17734);
and U23167 (N_23167,N_15779,N_19890);
xnor U23168 (N_23168,N_17892,N_17035);
nor U23169 (N_23169,N_17123,N_15351);
xor U23170 (N_23170,N_19804,N_15546);
or U23171 (N_23171,N_17909,N_16601);
or U23172 (N_23172,N_17869,N_16015);
nor U23173 (N_23173,N_18249,N_16392);
nor U23174 (N_23174,N_15113,N_15462);
nand U23175 (N_23175,N_16598,N_16445);
xor U23176 (N_23176,N_17302,N_16805);
or U23177 (N_23177,N_15331,N_17465);
nand U23178 (N_23178,N_16165,N_15014);
or U23179 (N_23179,N_15189,N_18490);
nand U23180 (N_23180,N_17874,N_18914);
and U23181 (N_23181,N_17337,N_19821);
and U23182 (N_23182,N_15196,N_15508);
nand U23183 (N_23183,N_15321,N_19462);
and U23184 (N_23184,N_18455,N_17450);
nor U23185 (N_23185,N_17590,N_16127);
nand U23186 (N_23186,N_15800,N_15278);
and U23187 (N_23187,N_15874,N_15579);
nor U23188 (N_23188,N_17799,N_17123);
nand U23189 (N_23189,N_15205,N_18928);
and U23190 (N_23190,N_17204,N_19303);
nor U23191 (N_23191,N_16496,N_19912);
or U23192 (N_23192,N_16181,N_18263);
and U23193 (N_23193,N_16010,N_16874);
nand U23194 (N_23194,N_16677,N_18058);
or U23195 (N_23195,N_15011,N_18944);
and U23196 (N_23196,N_16828,N_16234);
nor U23197 (N_23197,N_18405,N_16915);
nor U23198 (N_23198,N_15051,N_17606);
xor U23199 (N_23199,N_17505,N_18767);
xnor U23200 (N_23200,N_17203,N_18546);
and U23201 (N_23201,N_19400,N_18593);
nor U23202 (N_23202,N_19495,N_19546);
xor U23203 (N_23203,N_17728,N_16371);
and U23204 (N_23204,N_15217,N_17468);
or U23205 (N_23205,N_19043,N_18745);
nand U23206 (N_23206,N_18026,N_15840);
or U23207 (N_23207,N_18620,N_16830);
xnor U23208 (N_23208,N_16075,N_15547);
nand U23209 (N_23209,N_16935,N_16373);
nand U23210 (N_23210,N_18579,N_19111);
or U23211 (N_23211,N_16478,N_18587);
nor U23212 (N_23212,N_18201,N_17980);
nand U23213 (N_23213,N_15183,N_18908);
and U23214 (N_23214,N_17789,N_19966);
nor U23215 (N_23215,N_17998,N_19063);
or U23216 (N_23216,N_17212,N_17090);
nand U23217 (N_23217,N_15322,N_16346);
or U23218 (N_23218,N_19641,N_15260);
xnor U23219 (N_23219,N_16633,N_15981);
or U23220 (N_23220,N_16764,N_15533);
xor U23221 (N_23221,N_17305,N_18816);
or U23222 (N_23222,N_16827,N_17851);
and U23223 (N_23223,N_18376,N_16827);
and U23224 (N_23224,N_15629,N_17287);
or U23225 (N_23225,N_16285,N_15338);
nor U23226 (N_23226,N_18947,N_15733);
nand U23227 (N_23227,N_19844,N_16798);
and U23228 (N_23228,N_19034,N_16198);
nor U23229 (N_23229,N_19288,N_17612);
xnor U23230 (N_23230,N_16051,N_17192);
nand U23231 (N_23231,N_18802,N_18259);
nand U23232 (N_23232,N_16577,N_17167);
and U23233 (N_23233,N_16780,N_16063);
nand U23234 (N_23234,N_15556,N_16875);
or U23235 (N_23235,N_15712,N_16471);
and U23236 (N_23236,N_15328,N_15976);
nor U23237 (N_23237,N_19410,N_15069);
or U23238 (N_23238,N_19509,N_15844);
nand U23239 (N_23239,N_15720,N_15638);
and U23240 (N_23240,N_15622,N_15123);
and U23241 (N_23241,N_17646,N_15111);
or U23242 (N_23242,N_19954,N_19107);
xor U23243 (N_23243,N_19990,N_19547);
or U23244 (N_23244,N_15269,N_16876);
nor U23245 (N_23245,N_15809,N_15177);
nand U23246 (N_23246,N_17392,N_19652);
or U23247 (N_23247,N_18181,N_15946);
xor U23248 (N_23248,N_18121,N_19273);
and U23249 (N_23249,N_17883,N_16373);
and U23250 (N_23250,N_15603,N_17358);
and U23251 (N_23251,N_17239,N_15849);
and U23252 (N_23252,N_17649,N_19580);
nor U23253 (N_23253,N_15529,N_16465);
and U23254 (N_23254,N_18705,N_15759);
or U23255 (N_23255,N_17467,N_19816);
and U23256 (N_23256,N_18672,N_18125);
nor U23257 (N_23257,N_19598,N_18790);
or U23258 (N_23258,N_16417,N_16650);
nor U23259 (N_23259,N_16320,N_15392);
nor U23260 (N_23260,N_16682,N_17816);
nor U23261 (N_23261,N_18331,N_16572);
and U23262 (N_23262,N_18859,N_18712);
xor U23263 (N_23263,N_16080,N_18081);
nor U23264 (N_23264,N_15596,N_16343);
nor U23265 (N_23265,N_19757,N_18262);
nor U23266 (N_23266,N_17445,N_16789);
xor U23267 (N_23267,N_17717,N_15670);
and U23268 (N_23268,N_17284,N_19487);
and U23269 (N_23269,N_15170,N_19470);
or U23270 (N_23270,N_17628,N_15329);
nand U23271 (N_23271,N_18408,N_19019);
nand U23272 (N_23272,N_16122,N_19578);
nand U23273 (N_23273,N_15295,N_17530);
nor U23274 (N_23274,N_18662,N_16008);
and U23275 (N_23275,N_17605,N_17488);
nand U23276 (N_23276,N_15978,N_17434);
or U23277 (N_23277,N_18988,N_18110);
and U23278 (N_23278,N_15884,N_16564);
nor U23279 (N_23279,N_16032,N_17847);
and U23280 (N_23280,N_16506,N_18828);
and U23281 (N_23281,N_18188,N_16430);
and U23282 (N_23282,N_19907,N_15920);
or U23283 (N_23283,N_17826,N_16031);
nor U23284 (N_23284,N_19157,N_19422);
or U23285 (N_23285,N_18034,N_15602);
xor U23286 (N_23286,N_18878,N_19821);
nand U23287 (N_23287,N_19495,N_19456);
and U23288 (N_23288,N_19109,N_19215);
or U23289 (N_23289,N_17243,N_15205);
nand U23290 (N_23290,N_18616,N_16260);
or U23291 (N_23291,N_17281,N_19994);
or U23292 (N_23292,N_16658,N_17248);
or U23293 (N_23293,N_16159,N_19595);
xnor U23294 (N_23294,N_16635,N_19642);
nor U23295 (N_23295,N_18330,N_17833);
nand U23296 (N_23296,N_18710,N_18950);
xor U23297 (N_23297,N_15013,N_16766);
nor U23298 (N_23298,N_19498,N_16002);
nor U23299 (N_23299,N_15170,N_17242);
nand U23300 (N_23300,N_16862,N_15293);
or U23301 (N_23301,N_15197,N_17177);
and U23302 (N_23302,N_18001,N_17314);
nand U23303 (N_23303,N_18603,N_19660);
nand U23304 (N_23304,N_18774,N_19516);
nand U23305 (N_23305,N_18770,N_16828);
nor U23306 (N_23306,N_19894,N_17774);
or U23307 (N_23307,N_16705,N_16183);
nor U23308 (N_23308,N_18336,N_17850);
xor U23309 (N_23309,N_16098,N_16854);
nor U23310 (N_23310,N_19906,N_17486);
nand U23311 (N_23311,N_17009,N_17568);
nand U23312 (N_23312,N_18512,N_19887);
nand U23313 (N_23313,N_19994,N_15704);
nor U23314 (N_23314,N_19998,N_16869);
nand U23315 (N_23315,N_18296,N_18343);
and U23316 (N_23316,N_16924,N_17274);
or U23317 (N_23317,N_15151,N_19751);
nor U23318 (N_23318,N_19252,N_19707);
nand U23319 (N_23319,N_18686,N_18900);
nor U23320 (N_23320,N_17660,N_18965);
nand U23321 (N_23321,N_17305,N_19920);
nand U23322 (N_23322,N_16721,N_19562);
or U23323 (N_23323,N_16697,N_17715);
and U23324 (N_23324,N_18741,N_19565);
or U23325 (N_23325,N_15626,N_17582);
nand U23326 (N_23326,N_16817,N_15242);
or U23327 (N_23327,N_16821,N_18848);
and U23328 (N_23328,N_16478,N_19166);
nand U23329 (N_23329,N_17881,N_16740);
nor U23330 (N_23330,N_18560,N_15148);
nand U23331 (N_23331,N_15365,N_18309);
nor U23332 (N_23332,N_18371,N_18604);
nand U23333 (N_23333,N_19107,N_15157);
nor U23334 (N_23334,N_19355,N_17183);
or U23335 (N_23335,N_19751,N_16882);
or U23336 (N_23336,N_16409,N_16250);
and U23337 (N_23337,N_16811,N_17278);
xor U23338 (N_23338,N_18207,N_17401);
and U23339 (N_23339,N_18409,N_19257);
nor U23340 (N_23340,N_18019,N_16620);
nor U23341 (N_23341,N_18337,N_19503);
and U23342 (N_23342,N_16651,N_17144);
or U23343 (N_23343,N_16654,N_19056);
nand U23344 (N_23344,N_17126,N_19122);
or U23345 (N_23345,N_15550,N_17159);
or U23346 (N_23346,N_17679,N_18243);
or U23347 (N_23347,N_15511,N_17359);
nor U23348 (N_23348,N_19808,N_19047);
nand U23349 (N_23349,N_15476,N_18962);
or U23350 (N_23350,N_19671,N_19345);
or U23351 (N_23351,N_15157,N_16190);
or U23352 (N_23352,N_17496,N_19918);
nor U23353 (N_23353,N_19029,N_18899);
and U23354 (N_23354,N_16992,N_16340);
and U23355 (N_23355,N_17327,N_19312);
or U23356 (N_23356,N_19257,N_18805);
or U23357 (N_23357,N_19377,N_17196);
xor U23358 (N_23358,N_15456,N_15822);
or U23359 (N_23359,N_15324,N_16272);
xnor U23360 (N_23360,N_15275,N_16327);
and U23361 (N_23361,N_17494,N_16514);
and U23362 (N_23362,N_16611,N_17311);
nand U23363 (N_23363,N_17824,N_17267);
nand U23364 (N_23364,N_17312,N_17192);
nor U23365 (N_23365,N_18166,N_18559);
nand U23366 (N_23366,N_18782,N_18499);
nand U23367 (N_23367,N_18933,N_18456);
or U23368 (N_23368,N_16144,N_15814);
nor U23369 (N_23369,N_19069,N_15630);
and U23370 (N_23370,N_18513,N_17678);
and U23371 (N_23371,N_18360,N_19374);
and U23372 (N_23372,N_16673,N_17012);
or U23373 (N_23373,N_16801,N_15209);
and U23374 (N_23374,N_15644,N_18410);
or U23375 (N_23375,N_17022,N_16977);
and U23376 (N_23376,N_16856,N_15525);
nor U23377 (N_23377,N_15830,N_17679);
nor U23378 (N_23378,N_18782,N_19331);
or U23379 (N_23379,N_16949,N_19834);
nor U23380 (N_23380,N_17188,N_16940);
and U23381 (N_23381,N_16748,N_18314);
nand U23382 (N_23382,N_15864,N_15767);
and U23383 (N_23383,N_18849,N_19977);
nor U23384 (N_23384,N_18919,N_15960);
or U23385 (N_23385,N_17709,N_16002);
or U23386 (N_23386,N_16117,N_16596);
nand U23387 (N_23387,N_17553,N_17458);
or U23388 (N_23388,N_15054,N_16925);
nor U23389 (N_23389,N_15711,N_18280);
xor U23390 (N_23390,N_18440,N_17953);
nand U23391 (N_23391,N_16692,N_17945);
nor U23392 (N_23392,N_17056,N_16526);
xnor U23393 (N_23393,N_18215,N_15060);
or U23394 (N_23394,N_17783,N_18520);
or U23395 (N_23395,N_16257,N_15753);
nor U23396 (N_23396,N_15080,N_18300);
nand U23397 (N_23397,N_19158,N_17677);
and U23398 (N_23398,N_18904,N_19443);
and U23399 (N_23399,N_15976,N_18371);
nor U23400 (N_23400,N_16962,N_15284);
xor U23401 (N_23401,N_18385,N_19499);
nand U23402 (N_23402,N_16505,N_19746);
nand U23403 (N_23403,N_16796,N_19628);
nor U23404 (N_23404,N_17119,N_19144);
and U23405 (N_23405,N_19479,N_17565);
or U23406 (N_23406,N_17703,N_18010);
nor U23407 (N_23407,N_17093,N_17028);
nor U23408 (N_23408,N_16627,N_18150);
nor U23409 (N_23409,N_16822,N_15898);
nand U23410 (N_23410,N_18376,N_18404);
nand U23411 (N_23411,N_17154,N_17387);
or U23412 (N_23412,N_16832,N_15242);
xnor U23413 (N_23413,N_15866,N_17612);
or U23414 (N_23414,N_17709,N_16652);
nand U23415 (N_23415,N_18177,N_16798);
nand U23416 (N_23416,N_16031,N_19005);
nor U23417 (N_23417,N_18150,N_16265);
or U23418 (N_23418,N_17753,N_15321);
or U23419 (N_23419,N_19027,N_19611);
nand U23420 (N_23420,N_15787,N_18548);
or U23421 (N_23421,N_18674,N_16926);
and U23422 (N_23422,N_16006,N_16282);
nand U23423 (N_23423,N_18095,N_17301);
or U23424 (N_23424,N_16360,N_16630);
xor U23425 (N_23425,N_19521,N_15452);
or U23426 (N_23426,N_17690,N_17517);
and U23427 (N_23427,N_18239,N_19646);
and U23428 (N_23428,N_16452,N_15917);
nor U23429 (N_23429,N_16876,N_17031);
or U23430 (N_23430,N_15618,N_18068);
or U23431 (N_23431,N_18777,N_16065);
nor U23432 (N_23432,N_19154,N_18995);
xor U23433 (N_23433,N_15552,N_17639);
nor U23434 (N_23434,N_19560,N_15313);
or U23435 (N_23435,N_17850,N_18182);
and U23436 (N_23436,N_15417,N_16352);
xor U23437 (N_23437,N_17231,N_16873);
or U23438 (N_23438,N_17576,N_19359);
and U23439 (N_23439,N_17939,N_17320);
and U23440 (N_23440,N_17520,N_17571);
xor U23441 (N_23441,N_19219,N_15753);
and U23442 (N_23442,N_15533,N_16966);
nor U23443 (N_23443,N_17046,N_19320);
and U23444 (N_23444,N_18409,N_18603);
and U23445 (N_23445,N_18471,N_16002);
or U23446 (N_23446,N_17396,N_16401);
or U23447 (N_23447,N_17572,N_18399);
nor U23448 (N_23448,N_15301,N_17019);
nor U23449 (N_23449,N_15851,N_17511);
nor U23450 (N_23450,N_15435,N_19876);
nor U23451 (N_23451,N_15067,N_17049);
nor U23452 (N_23452,N_16793,N_16245);
and U23453 (N_23453,N_15085,N_15912);
nand U23454 (N_23454,N_18565,N_17956);
nor U23455 (N_23455,N_19188,N_17900);
or U23456 (N_23456,N_19617,N_18954);
or U23457 (N_23457,N_18656,N_19536);
nor U23458 (N_23458,N_16831,N_17554);
or U23459 (N_23459,N_18594,N_18496);
nor U23460 (N_23460,N_19072,N_15757);
nand U23461 (N_23461,N_17325,N_16091);
and U23462 (N_23462,N_17544,N_16476);
or U23463 (N_23463,N_15271,N_16121);
nor U23464 (N_23464,N_15704,N_15534);
xor U23465 (N_23465,N_17055,N_16745);
nor U23466 (N_23466,N_19649,N_15117);
nand U23467 (N_23467,N_16044,N_18802);
and U23468 (N_23468,N_16781,N_19794);
nor U23469 (N_23469,N_16491,N_17300);
and U23470 (N_23470,N_17531,N_18205);
nand U23471 (N_23471,N_16347,N_17760);
xnor U23472 (N_23472,N_17449,N_16720);
nor U23473 (N_23473,N_17449,N_16471);
and U23474 (N_23474,N_19098,N_18611);
nor U23475 (N_23475,N_15054,N_19589);
nand U23476 (N_23476,N_17242,N_17360);
or U23477 (N_23477,N_17194,N_18477);
or U23478 (N_23478,N_15634,N_19672);
nor U23479 (N_23479,N_16170,N_15785);
nor U23480 (N_23480,N_18081,N_17622);
nor U23481 (N_23481,N_18416,N_15533);
and U23482 (N_23482,N_15270,N_19423);
nand U23483 (N_23483,N_18904,N_19166);
nand U23484 (N_23484,N_15439,N_19288);
nor U23485 (N_23485,N_16890,N_17453);
and U23486 (N_23486,N_16001,N_19729);
nand U23487 (N_23487,N_19967,N_17244);
and U23488 (N_23488,N_19550,N_19882);
nor U23489 (N_23489,N_18181,N_19584);
nor U23490 (N_23490,N_19363,N_17175);
xor U23491 (N_23491,N_15881,N_15460);
nor U23492 (N_23492,N_17483,N_19804);
nand U23493 (N_23493,N_17541,N_16802);
and U23494 (N_23494,N_19329,N_19849);
nand U23495 (N_23495,N_16393,N_15905);
or U23496 (N_23496,N_18170,N_15860);
nand U23497 (N_23497,N_19627,N_18568);
and U23498 (N_23498,N_17644,N_18139);
and U23499 (N_23499,N_18431,N_16813);
nor U23500 (N_23500,N_15053,N_16557);
nor U23501 (N_23501,N_17466,N_18730);
nor U23502 (N_23502,N_17240,N_17449);
nand U23503 (N_23503,N_19352,N_18306);
nand U23504 (N_23504,N_18986,N_18175);
and U23505 (N_23505,N_19235,N_16916);
and U23506 (N_23506,N_19509,N_17722);
nand U23507 (N_23507,N_15741,N_15162);
nand U23508 (N_23508,N_16918,N_16300);
xor U23509 (N_23509,N_16609,N_18676);
nand U23510 (N_23510,N_18203,N_19271);
or U23511 (N_23511,N_17774,N_19959);
and U23512 (N_23512,N_19248,N_19162);
nor U23513 (N_23513,N_18728,N_18245);
or U23514 (N_23514,N_15850,N_17809);
nand U23515 (N_23515,N_15777,N_17244);
or U23516 (N_23516,N_15628,N_15953);
nand U23517 (N_23517,N_18817,N_18916);
and U23518 (N_23518,N_19333,N_16023);
nor U23519 (N_23519,N_16945,N_15577);
or U23520 (N_23520,N_15478,N_16023);
nor U23521 (N_23521,N_19769,N_17097);
nor U23522 (N_23522,N_17586,N_18685);
or U23523 (N_23523,N_17500,N_16012);
and U23524 (N_23524,N_17525,N_16831);
nor U23525 (N_23525,N_19036,N_19817);
nand U23526 (N_23526,N_19252,N_15487);
nor U23527 (N_23527,N_19604,N_17904);
nor U23528 (N_23528,N_16542,N_17599);
and U23529 (N_23529,N_17072,N_15507);
and U23530 (N_23530,N_17052,N_17758);
nand U23531 (N_23531,N_15987,N_17642);
or U23532 (N_23532,N_17873,N_16586);
nor U23533 (N_23533,N_15122,N_16018);
xnor U23534 (N_23534,N_15254,N_17599);
and U23535 (N_23535,N_18279,N_18466);
nor U23536 (N_23536,N_16346,N_15982);
nor U23537 (N_23537,N_19430,N_15753);
and U23538 (N_23538,N_16869,N_17200);
nor U23539 (N_23539,N_16301,N_18868);
or U23540 (N_23540,N_18254,N_19516);
nand U23541 (N_23541,N_19427,N_19883);
and U23542 (N_23542,N_19959,N_19145);
and U23543 (N_23543,N_19204,N_17609);
nor U23544 (N_23544,N_18603,N_15779);
nor U23545 (N_23545,N_17621,N_17102);
and U23546 (N_23546,N_17390,N_19972);
nand U23547 (N_23547,N_15163,N_18797);
nand U23548 (N_23548,N_18564,N_17048);
and U23549 (N_23549,N_15443,N_18021);
nand U23550 (N_23550,N_19548,N_16495);
or U23551 (N_23551,N_19446,N_19089);
nor U23552 (N_23552,N_16754,N_16038);
or U23553 (N_23553,N_15968,N_15527);
or U23554 (N_23554,N_15444,N_16584);
nor U23555 (N_23555,N_18592,N_16416);
nand U23556 (N_23556,N_19011,N_17565);
nand U23557 (N_23557,N_18897,N_17970);
nor U23558 (N_23558,N_19466,N_19200);
nand U23559 (N_23559,N_15450,N_18189);
xor U23560 (N_23560,N_19524,N_17400);
or U23561 (N_23561,N_18764,N_18824);
and U23562 (N_23562,N_19513,N_17476);
and U23563 (N_23563,N_18698,N_18584);
nand U23564 (N_23564,N_15816,N_16261);
and U23565 (N_23565,N_18215,N_15544);
or U23566 (N_23566,N_18945,N_17871);
or U23567 (N_23567,N_19870,N_16724);
or U23568 (N_23568,N_18040,N_19872);
nor U23569 (N_23569,N_16114,N_17403);
nand U23570 (N_23570,N_19294,N_17084);
and U23571 (N_23571,N_18231,N_16093);
nand U23572 (N_23572,N_18434,N_15831);
nand U23573 (N_23573,N_17157,N_15999);
nor U23574 (N_23574,N_18207,N_16512);
nand U23575 (N_23575,N_18471,N_15340);
nor U23576 (N_23576,N_18587,N_19377);
nor U23577 (N_23577,N_17063,N_19839);
or U23578 (N_23578,N_18801,N_16934);
xor U23579 (N_23579,N_15196,N_17241);
nand U23580 (N_23580,N_15520,N_15452);
nand U23581 (N_23581,N_18330,N_18942);
or U23582 (N_23582,N_15814,N_19223);
nor U23583 (N_23583,N_16166,N_19809);
nand U23584 (N_23584,N_18733,N_18950);
or U23585 (N_23585,N_16260,N_19641);
or U23586 (N_23586,N_18876,N_17928);
and U23587 (N_23587,N_19549,N_16859);
or U23588 (N_23588,N_18106,N_18921);
nand U23589 (N_23589,N_18458,N_18505);
or U23590 (N_23590,N_15980,N_15607);
or U23591 (N_23591,N_15151,N_16244);
nor U23592 (N_23592,N_19643,N_18143);
xor U23593 (N_23593,N_16072,N_18919);
nor U23594 (N_23594,N_17543,N_17204);
or U23595 (N_23595,N_16062,N_18741);
or U23596 (N_23596,N_19153,N_18095);
nor U23597 (N_23597,N_16432,N_15500);
nor U23598 (N_23598,N_16949,N_17463);
or U23599 (N_23599,N_16581,N_18300);
or U23600 (N_23600,N_19540,N_15180);
nor U23601 (N_23601,N_17015,N_19642);
or U23602 (N_23602,N_19672,N_19923);
and U23603 (N_23603,N_16061,N_15775);
or U23604 (N_23604,N_18665,N_19561);
and U23605 (N_23605,N_19980,N_18590);
or U23606 (N_23606,N_17465,N_15120);
nor U23607 (N_23607,N_15339,N_19962);
and U23608 (N_23608,N_17498,N_16839);
or U23609 (N_23609,N_17138,N_17990);
nor U23610 (N_23610,N_18077,N_16374);
nor U23611 (N_23611,N_17429,N_18105);
nand U23612 (N_23612,N_19508,N_15884);
nor U23613 (N_23613,N_15060,N_17852);
and U23614 (N_23614,N_17862,N_15512);
or U23615 (N_23615,N_19834,N_19339);
nor U23616 (N_23616,N_15489,N_18358);
or U23617 (N_23617,N_16679,N_19738);
nand U23618 (N_23618,N_15763,N_17536);
or U23619 (N_23619,N_16200,N_17037);
and U23620 (N_23620,N_18211,N_18572);
nand U23621 (N_23621,N_18333,N_19300);
or U23622 (N_23622,N_15934,N_15069);
and U23623 (N_23623,N_16164,N_16634);
or U23624 (N_23624,N_18906,N_15658);
nand U23625 (N_23625,N_15467,N_16244);
xnor U23626 (N_23626,N_15552,N_18959);
or U23627 (N_23627,N_19830,N_16781);
nand U23628 (N_23628,N_17357,N_18497);
and U23629 (N_23629,N_19583,N_19176);
and U23630 (N_23630,N_19447,N_19664);
nor U23631 (N_23631,N_18611,N_17515);
or U23632 (N_23632,N_18196,N_18404);
and U23633 (N_23633,N_16395,N_17490);
xnor U23634 (N_23634,N_15682,N_17916);
or U23635 (N_23635,N_16875,N_15682);
or U23636 (N_23636,N_17674,N_17319);
nor U23637 (N_23637,N_18482,N_19950);
nand U23638 (N_23638,N_18869,N_19489);
or U23639 (N_23639,N_17554,N_19156);
and U23640 (N_23640,N_19180,N_19341);
and U23641 (N_23641,N_17459,N_18852);
and U23642 (N_23642,N_16393,N_18036);
or U23643 (N_23643,N_19334,N_19105);
or U23644 (N_23644,N_18332,N_17210);
nor U23645 (N_23645,N_16568,N_19785);
or U23646 (N_23646,N_17222,N_19018);
and U23647 (N_23647,N_18672,N_16393);
nor U23648 (N_23648,N_15002,N_19090);
nor U23649 (N_23649,N_18823,N_15015);
or U23650 (N_23650,N_15411,N_17329);
or U23651 (N_23651,N_16915,N_19741);
nor U23652 (N_23652,N_18329,N_15246);
and U23653 (N_23653,N_18065,N_19142);
nor U23654 (N_23654,N_15187,N_16988);
xor U23655 (N_23655,N_16247,N_16483);
or U23656 (N_23656,N_17713,N_18750);
and U23657 (N_23657,N_19989,N_17810);
nand U23658 (N_23658,N_19820,N_16726);
xor U23659 (N_23659,N_17338,N_16072);
nor U23660 (N_23660,N_15851,N_15408);
xor U23661 (N_23661,N_18877,N_19616);
nor U23662 (N_23662,N_18735,N_18398);
nor U23663 (N_23663,N_15329,N_17799);
and U23664 (N_23664,N_19347,N_17910);
or U23665 (N_23665,N_17375,N_16261);
or U23666 (N_23666,N_17451,N_19073);
or U23667 (N_23667,N_19293,N_18582);
and U23668 (N_23668,N_17342,N_18874);
nand U23669 (N_23669,N_16943,N_15838);
and U23670 (N_23670,N_18151,N_15882);
and U23671 (N_23671,N_15708,N_16024);
or U23672 (N_23672,N_16101,N_18361);
nand U23673 (N_23673,N_18939,N_18858);
xor U23674 (N_23674,N_19780,N_15321);
and U23675 (N_23675,N_18426,N_17019);
and U23676 (N_23676,N_19328,N_16027);
or U23677 (N_23677,N_16482,N_17275);
nor U23678 (N_23678,N_19707,N_15373);
nor U23679 (N_23679,N_17855,N_15604);
or U23680 (N_23680,N_17114,N_17995);
xor U23681 (N_23681,N_15954,N_19957);
nor U23682 (N_23682,N_17765,N_18247);
or U23683 (N_23683,N_15006,N_18480);
nor U23684 (N_23684,N_15748,N_17565);
nand U23685 (N_23685,N_16268,N_15126);
or U23686 (N_23686,N_16797,N_17894);
xor U23687 (N_23687,N_16848,N_16719);
or U23688 (N_23688,N_15772,N_16699);
nor U23689 (N_23689,N_19163,N_16512);
nor U23690 (N_23690,N_17170,N_19140);
nor U23691 (N_23691,N_19110,N_18974);
nor U23692 (N_23692,N_16581,N_17639);
nor U23693 (N_23693,N_17213,N_19245);
or U23694 (N_23694,N_18851,N_15476);
nor U23695 (N_23695,N_19758,N_19118);
or U23696 (N_23696,N_17189,N_15122);
nand U23697 (N_23697,N_17700,N_18619);
nor U23698 (N_23698,N_18319,N_17270);
or U23699 (N_23699,N_17535,N_15589);
xor U23700 (N_23700,N_16765,N_19090);
and U23701 (N_23701,N_18291,N_17403);
nand U23702 (N_23702,N_18481,N_15148);
nor U23703 (N_23703,N_15961,N_18441);
nor U23704 (N_23704,N_17702,N_15558);
and U23705 (N_23705,N_17817,N_17797);
or U23706 (N_23706,N_18284,N_19600);
nand U23707 (N_23707,N_18794,N_18489);
nand U23708 (N_23708,N_17878,N_16284);
or U23709 (N_23709,N_19961,N_16600);
and U23710 (N_23710,N_17821,N_19861);
nor U23711 (N_23711,N_16659,N_16648);
nand U23712 (N_23712,N_15828,N_16956);
nand U23713 (N_23713,N_16786,N_18031);
and U23714 (N_23714,N_18297,N_18645);
nand U23715 (N_23715,N_16644,N_18344);
nor U23716 (N_23716,N_18536,N_15844);
xor U23717 (N_23717,N_17140,N_16988);
xor U23718 (N_23718,N_17345,N_18349);
and U23719 (N_23719,N_16187,N_18134);
and U23720 (N_23720,N_18202,N_15512);
nor U23721 (N_23721,N_17714,N_17301);
nand U23722 (N_23722,N_18532,N_19839);
and U23723 (N_23723,N_16171,N_17542);
and U23724 (N_23724,N_18550,N_15622);
nand U23725 (N_23725,N_15472,N_17605);
nor U23726 (N_23726,N_18620,N_18410);
and U23727 (N_23727,N_19954,N_16207);
xnor U23728 (N_23728,N_15845,N_15068);
nand U23729 (N_23729,N_18443,N_15948);
nand U23730 (N_23730,N_19792,N_15970);
or U23731 (N_23731,N_17054,N_15259);
xnor U23732 (N_23732,N_16401,N_16138);
xnor U23733 (N_23733,N_17690,N_15545);
or U23734 (N_23734,N_19353,N_19809);
or U23735 (N_23735,N_17819,N_19597);
and U23736 (N_23736,N_17810,N_18680);
nor U23737 (N_23737,N_15511,N_19909);
and U23738 (N_23738,N_16261,N_18151);
nor U23739 (N_23739,N_19513,N_16195);
nor U23740 (N_23740,N_16519,N_16071);
nor U23741 (N_23741,N_16476,N_18253);
nor U23742 (N_23742,N_18432,N_17369);
or U23743 (N_23743,N_17259,N_19297);
nand U23744 (N_23744,N_19303,N_19160);
or U23745 (N_23745,N_19659,N_18868);
nor U23746 (N_23746,N_16476,N_19457);
nand U23747 (N_23747,N_19634,N_15518);
or U23748 (N_23748,N_15830,N_16063);
xor U23749 (N_23749,N_16945,N_15648);
nand U23750 (N_23750,N_18352,N_18766);
and U23751 (N_23751,N_15099,N_18739);
and U23752 (N_23752,N_15436,N_15345);
nor U23753 (N_23753,N_16575,N_17327);
nand U23754 (N_23754,N_18432,N_17472);
and U23755 (N_23755,N_18258,N_18540);
or U23756 (N_23756,N_16389,N_15359);
nand U23757 (N_23757,N_15879,N_19584);
and U23758 (N_23758,N_17410,N_19141);
nor U23759 (N_23759,N_18378,N_18228);
or U23760 (N_23760,N_18376,N_16438);
nand U23761 (N_23761,N_17589,N_16919);
or U23762 (N_23762,N_15939,N_15594);
nor U23763 (N_23763,N_18614,N_16597);
nand U23764 (N_23764,N_19167,N_17613);
nand U23765 (N_23765,N_18379,N_18112);
and U23766 (N_23766,N_17638,N_16118);
nor U23767 (N_23767,N_15551,N_16410);
nand U23768 (N_23768,N_16226,N_17771);
or U23769 (N_23769,N_18048,N_19642);
and U23770 (N_23770,N_18174,N_18640);
or U23771 (N_23771,N_16965,N_16160);
nand U23772 (N_23772,N_17580,N_16348);
nor U23773 (N_23773,N_15497,N_16203);
nand U23774 (N_23774,N_18446,N_15042);
nand U23775 (N_23775,N_18350,N_18895);
and U23776 (N_23776,N_17489,N_17496);
or U23777 (N_23777,N_18898,N_17986);
and U23778 (N_23778,N_16209,N_16093);
and U23779 (N_23779,N_19732,N_16912);
nand U23780 (N_23780,N_15569,N_16663);
xnor U23781 (N_23781,N_19778,N_15667);
or U23782 (N_23782,N_17865,N_17997);
or U23783 (N_23783,N_19423,N_18343);
xnor U23784 (N_23784,N_18500,N_19924);
xnor U23785 (N_23785,N_16400,N_15416);
nor U23786 (N_23786,N_15756,N_17274);
or U23787 (N_23787,N_15693,N_19322);
or U23788 (N_23788,N_15697,N_16773);
or U23789 (N_23789,N_17748,N_15645);
and U23790 (N_23790,N_17174,N_16353);
or U23791 (N_23791,N_18485,N_16376);
nand U23792 (N_23792,N_19079,N_17373);
or U23793 (N_23793,N_18316,N_15410);
nor U23794 (N_23794,N_19112,N_15184);
nor U23795 (N_23795,N_17672,N_18034);
nor U23796 (N_23796,N_18120,N_18285);
and U23797 (N_23797,N_17012,N_16689);
nand U23798 (N_23798,N_19599,N_15408);
nor U23799 (N_23799,N_19597,N_19404);
nand U23800 (N_23800,N_19850,N_19291);
nand U23801 (N_23801,N_18386,N_17979);
nand U23802 (N_23802,N_16206,N_18066);
and U23803 (N_23803,N_16109,N_16531);
nand U23804 (N_23804,N_17335,N_19703);
xor U23805 (N_23805,N_19628,N_19265);
nand U23806 (N_23806,N_15673,N_18806);
or U23807 (N_23807,N_19638,N_15730);
nand U23808 (N_23808,N_19047,N_19909);
or U23809 (N_23809,N_19316,N_15747);
nand U23810 (N_23810,N_16033,N_18136);
nor U23811 (N_23811,N_15162,N_15175);
xor U23812 (N_23812,N_17925,N_18881);
nand U23813 (N_23813,N_19433,N_19924);
xor U23814 (N_23814,N_19816,N_17545);
xnor U23815 (N_23815,N_15882,N_16233);
or U23816 (N_23816,N_15212,N_16770);
nand U23817 (N_23817,N_16207,N_19481);
and U23818 (N_23818,N_18575,N_18408);
nand U23819 (N_23819,N_18058,N_19452);
nand U23820 (N_23820,N_15993,N_17028);
nor U23821 (N_23821,N_15284,N_17227);
nor U23822 (N_23822,N_15968,N_19320);
xnor U23823 (N_23823,N_17814,N_15474);
xnor U23824 (N_23824,N_19300,N_18205);
and U23825 (N_23825,N_16154,N_18555);
xor U23826 (N_23826,N_18759,N_17914);
or U23827 (N_23827,N_17016,N_18902);
xor U23828 (N_23828,N_17328,N_19410);
nor U23829 (N_23829,N_17558,N_15267);
and U23830 (N_23830,N_15848,N_15975);
nor U23831 (N_23831,N_19146,N_18163);
nand U23832 (N_23832,N_18784,N_15591);
nor U23833 (N_23833,N_19153,N_18890);
nand U23834 (N_23834,N_17337,N_17393);
nand U23835 (N_23835,N_16789,N_17901);
or U23836 (N_23836,N_16473,N_19273);
nor U23837 (N_23837,N_15154,N_15881);
xnor U23838 (N_23838,N_18391,N_19541);
nand U23839 (N_23839,N_17019,N_19607);
nor U23840 (N_23840,N_15814,N_18078);
or U23841 (N_23841,N_17277,N_18266);
or U23842 (N_23842,N_19637,N_15352);
and U23843 (N_23843,N_16233,N_15243);
nor U23844 (N_23844,N_15564,N_16268);
and U23845 (N_23845,N_16104,N_19047);
and U23846 (N_23846,N_19593,N_19148);
or U23847 (N_23847,N_19509,N_19950);
nor U23848 (N_23848,N_15972,N_19789);
nor U23849 (N_23849,N_19836,N_18396);
or U23850 (N_23850,N_17033,N_15974);
nand U23851 (N_23851,N_16496,N_15046);
or U23852 (N_23852,N_15364,N_19448);
nand U23853 (N_23853,N_16980,N_19883);
nor U23854 (N_23854,N_19631,N_16716);
and U23855 (N_23855,N_17927,N_19892);
nand U23856 (N_23856,N_19401,N_18624);
nand U23857 (N_23857,N_16804,N_19197);
nand U23858 (N_23858,N_18362,N_17148);
and U23859 (N_23859,N_17133,N_16544);
nand U23860 (N_23860,N_19076,N_18954);
and U23861 (N_23861,N_18020,N_15717);
or U23862 (N_23862,N_15750,N_19387);
or U23863 (N_23863,N_16732,N_15252);
nand U23864 (N_23864,N_19379,N_16297);
or U23865 (N_23865,N_17657,N_16496);
or U23866 (N_23866,N_16081,N_15888);
nand U23867 (N_23867,N_19674,N_17983);
or U23868 (N_23868,N_15979,N_19448);
nand U23869 (N_23869,N_18988,N_18949);
and U23870 (N_23870,N_15474,N_18855);
and U23871 (N_23871,N_15695,N_19551);
or U23872 (N_23872,N_16916,N_17655);
or U23873 (N_23873,N_18057,N_16135);
nor U23874 (N_23874,N_17893,N_18700);
nand U23875 (N_23875,N_15315,N_17076);
or U23876 (N_23876,N_17478,N_19394);
and U23877 (N_23877,N_17578,N_15997);
and U23878 (N_23878,N_16258,N_15084);
and U23879 (N_23879,N_17600,N_18525);
or U23880 (N_23880,N_19229,N_18677);
nand U23881 (N_23881,N_16928,N_19925);
nand U23882 (N_23882,N_16992,N_18561);
xor U23883 (N_23883,N_16097,N_19218);
nand U23884 (N_23884,N_19765,N_15227);
nor U23885 (N_23885,N_19312,N_16791);
nor U23886 (N_23886,N_15110,N_15753);
and U23887 (N_23887,N_17032,N_17630);
and U23888 (N_23888,N_16572,N_19792);
and U23889 (N_23889,N_18352,N_15841);
or U23890 (N_23890,N_16862,N_18292);
nand U23891 (N_23891,N_18392,N_18508);
nand U23892 (N_23892,N_18512,N_17177);
or U23893 (N_23893,N_17305,N_19998);
nand U23894 (N_23894,N_16605,N_19619);
xnor U23895 (N_23895,N_17414,N_17652);
xor U23896 (N_23896,N_17626,N_18569);
nor U23897 (N_23897,N_16106,N_17607);
nand U23898 (N_23898,N_19053,N_18172);
and U23899 (N_23899,N_19882,N_17334);
and U23900 (N_23900,N_19945,N_17644);
nor U23901 (N_23901,N_17768,N_18505);
or U23902 (N_23902,N_17500,N_17512);
xnor U23903 (N_23903,N_18685,N_18792);
or U23904 (N_23904,N_18860,N_18863);
nand U23905 (N_23905,N_19242,N_19085);
nand U23906 (N_23906,N_18882,N_19233);
nand U23907 (N_23907,N_19565,N_17563);
or U23908 (N_23908,N_17883,N_15821);
or U23909 (N_23909,N_15539,N_16329);
and U23910 (N_23910,N_19292,N_18081);
and U23911 (N_23911,N_19424,N_16804);
nand U23912 (N_23912,N_15605,N_19794);
nand U23913 (N_23913,N_18996,N_16767);
nand U23914 (N_23914,N_15133,N_18496);
or U23915 (N_23915,N_16151,N_15855);
nor U23916 (N_23916,N_16191,N_18680);
xnor U23917 (N_23917,N_18845,N_18704);
or U23918 (N_23918,N_19581,N_16689);
and U23919 (N_23919,N_17599,N_16749);
nor U23920 (N_23920,N_18828,N_17392);
nand U23921 (N_23921,N_18139,N_15928);
nor U23922 (N_23922,N_18017,N_19802);
xor U23923 (N_23923,N_16216,N_15922);
and U23924 (N_23924,N_19675,N_18400);
nand U23925 (N_23925,N_16659,N_17958);
or U23926 (N_23926,N_18013,N_19167);
xor U23927 (N_23927,N_15717,N_17750);
or U23928 (N_23928,N_19134,N_15622);
nand U23929 (N_23929,N_18072,N_15851);
nand U23930 (N_23930,N_19947,N_17532);
xnor U23931 (N_23931,N_19102,N_19486);
nand U23932 (N_23932,N_19538,N_18835);
nor U23933 (N_23933,N_17928,N_18905);
nor U23934 (N_23934,N_17206,N_16071);
nand U23935 (N_23935,N_15606,N_18578);
and U23936 (N_23936,N_18276,N_17316);
xor U23937 (N_23937,N_15711,N_19401);
nand U23938 (N_23938,N_18235,N_16639);
or U23939 (N_23939,N_16935,N_18170);
nor U23940 (N_23940,N_18980,N_16723);
and U23941 (N_23941,N_17582,N_16950);
xor U23942 (N_23942,N_15512,N_17297);
or U23943 (N_23943,N_18766,N_15793);
xnor U23944 (N_23944,N_19752,N_17886);
or U23945 (N_23945,N_17991,N_15776);
nor U23946 (N_23946,N_16328,N_16767);
nand U23947 (N_23947,N_17741,N_15294);
nor U23948 (N_23948,N_16366,N_15215);
nand U23949 (N_23949,N_18039,N_16109);
nand U23950 (N_23950,N_16977,N_19317);
nor U23951 (N_23951,N_19699,N_15664);
or U23952 (N_23952,N_18566,N_15424);
and U23953 (N_23953,N_17698,N_19055);
nand U23954 (N_23954,N_15501,N_19145);
and U23955 (N_23955,N_18604,N_15233);
nor U23956 (N_23956,N_18348,N_16599);
nand U23957 (N_23957,N_18181,N_19931);
or U23958 (N_23958,N_16529,N_16312);
nor U23959 (N_23959,N_15160,N_17186);
and U23960 (N_23960,N_18324,N_17462);
nand U23961 (N_23961,N_16317,N_16890);
nor U23962 (N_23962,N_19695,N_18783);
or U23963 (N_23963,N_17034,N_16637);
or U23964 (N_23964,N_17565,N_17959);
xor U23965 (N_23965,N_17018,N_16658);
xor U23966 (N_23966,N_16993,N_19999);
nor U23967 (N_23967,N_17705,N_19075);
nor U23968 (N_23968,N_18318,N_15329);
or U23969 (N_23969,N_15113,N_15751);
and U23970 (N_23970,N_19407,N_18220);
and U23971 (N_23971,N_16173,N_15787);
or U23972 (N_23972,N_19175,N_19883);
nor U23973 (N_23973,N_18205,N_17693);
nor U23974 (N_23974,N_19650,N_16405);
xnor U23975 (N_23975,N_17065,N_16827);
nor U23976 (N_23976,N_19859,N_15673);
xor U23977 (N_23977,N_15890,N_16992);
nor U23978 (N_23978,N_19793,N_15326);
nor U23979 (N_23979,N_15275,N_18113);
or U23980 (N_23980,N_18428,N_17233);
nand U23981 (N_23981,N_17907,N_16814);
and U23982 (N_23982,N_15451,N_17560);
nand U23983 (N_23983,N_15963,N_16479);
nand U23984 (N_23984,N_19967,N_16160);
nor U23985 (N_23985,N_19321,N_18205);
nand U23986 (N_23986,N_17443,N_19103);
and U23987 (N_23987,N_19932,N_16435);
or U23988 (N_23988,N_18768,N_16113);
and U23989 (N_23989,N_15457,N_17928);
nand U23990 (N_23990,N_19115,N_17587);
or U23991 (N_23991,N_16082,N_19712);
xnor U23992 (N_23992,N_17657,N_19452);
and U23993 (N_23993,N_16328,N_17125);
nand U23994 (N_23994,N_15078,N_16518);
or U23995 (N_23995,N_17212,N_15940);
nand U23996 (N_23996,N_18728,N_17614);
nor U23997 (N_23997,N_15293,N_15551);
or U23998 (N_23998,N_16622,N_16277);
nor U23999 (N_23999,N_18225,N_15088);
xnor U24000 (N_24000,N_16920,N_17455);
or U24001 (N_24001,N_17910,N_18092);
or U24002 (N_24002,N_15904,N_19108);
nand U24003 (N_24003,N_15858,N_16730);
or U24004 (N_24004,N_17940,N_19225);
and U24005 (N_24005,N_16987,N_15734);
nor U24006 (N_24006,N_19052,N_17398);
or U24007 (N_24007,N_16699,N_18397);
xnor U24008 (N_24008,N_17623,N_19865);
or U24009 (N_24009,N_18059,N_16355);
xnor U24010 (N_24010,N_15321,N_15316);
and U24011 (N_24011,N_18767,N_16901);
nor U24012 (N_24012,N_19334,N_15278);
and U24013 (N_24013,N_15554,N_15046);
or U24014 (N_24014,N_19641,N_19565);
nand U24015 (N_24015,N_19247,N_19107);
and U24016 (N_24016,N_16261,N_19139);
or U24017 (N_24017,N_17271,N_17666);
nor U24018 (N_24018,N_19637,N_18169);
xor U24019 (N_24019,N_18849,N_19232);
nand U24020 (N_24020,N_16203,N_16524);
or U24021 (N_24021,N_18548,N_19965);
or U24022 (N_24022,N_15315,N_16388);
or U24023 (N_24023,N_15434,N_18889);
nand U24024 (N_24024,N_17108,N_16707);
and U24025 (N_24025,N_19243,N_18242);
nand U24026 (N_24026,N_16990,N_18441);
nor U24027 (N_24027,N_18326,N_19992);
nor U24028 (N_24028,N_17388,N_19472);
and U24029 (N_24029,N_18612,N_18110);
and U24030 (N_24030,N_17231,N_19167);
or U24031 (N_24031,N_19980,N_16557);
nor U24032 (N_24032,N_19883,N_15562);
and U24033 (N_24033,N_16519,N_15820);
nand U24034 (N_24034,N_16273,N_18018);
xor U24035 (N_24035,N_15530,N_18856);
nor U24036 (N_24036,N_16722,N_17154);
nand U24037 (N_24037,N_17409,N_17519);
and U24038 (N_24038,N_18055,N_17374);
and U24039 (N_24039,N_16963,N_15822);
nand U24040 (N_24040,N_15293,N_18503);
nand U24041 (N_24041,N_15538,N_15734);
or U24042 (N_24042,N_19581,N_16092);
xor U24043 (N_24043,N_15251,N_16357);
and U24044 (N_24044,N_18606,N_17574);
xnor U24045 (N_24045,N_15646,N_16052);
nor U24046 (N_24046,N_18910,N_15283);
and U24047 (N_24047,N_15012,N_15410);
nor U24048 (N_24048,N_16974,N_16398);
or U24049 (N_24049,N_17701,N_16119);
nor U24050 (N_24050,N_15127,N_17446);
xor U24051 (N_24051,N_15762,N_19414);
and U24052 (N_24052,N_15625,N_15089);
nor U24053 (N_24053,N_16959,N_19903);
and U24054 (N_24054,N_17402,N_19790);
nor U24055 (N_24055,N_17118,N_15740);
and U24056 (N_24056,N_19007,N_19726);
nand U24057 (N_24057,N_17220,N_19210);
and U24058 (N_24058,N_17826,N_17071);
or U24059 (N_24059,N_19683,N_16393);
or U24060 (N_24060,N_18965,N_17267);
nor U24061 (N_24061,N_17442,N_19440);
nand U24062 (N_24062,N_16290,N_16277);
or U24063 (N_24063,N_17381,N_18924);
nor U24064 (N_24064,N_16473,N_18148);
nor U24065 (N_24065,N_19229,N_19734);
nor U24066 (N_24066,N_16155,N_19734);
nand U24067 (N_24067,N_17325,N_17291);
and U24068 (N_24068,N_17118,N_15206);
nor U24069 (N_24069,N_15021,N_16215);
nand U24070 (N_24070,N_15687,N_16141);
nor U24071 (N_24071,N_18231,N_16987);
or U24072 (N_24072,N_18905,N_16544);
and U24073 (N_24073,N_17995,N_18222);
or U24074 (N_24074,N_15614,N_15180);
xnor U24075 (N_24075,N_15602,N_19923);
or U24076 (N_24076,N_19615,N_18009);
and U24077 (N_24077,N_17352,N_19901);
nand U24078 (N_24078,N_16020,N_15205);
xor U24079 (N_24079,N_19258,N_17053);
and U24080 (N_24080,N_18765,N_17126);
nand U24081 (N_24081,N_18684,N_19402);
xor U24082 (N_24082,N_18169,N_18571);
and U24083 (N_24083,N_15019,N_17598);
xnor U24084 (N_24084,N_17141,N_19047);
nor U24085 (N_24085,N_18915,N_16474);
or U24086 (N_24086,N_17221,N_19717);
or U24087 (N_24087,N_15666,N_19290);
xnor U24088 (N_24088,N_15526,N_19875);
nor U24089 (N_24089,N_19078,N_19322);
nand U24090 (N_24090,N_15529,N_18768);
nor U24091 (N_24091,N_18803,N_19095);
nor U24092 (N_24092,N_15431,N_16969);
nand U24093 (N_24093,N_15141,N_16140);
and U24094 (N_24094,N_18982,N_16482);
or U24095 (N_24095,N_16720,N_15912);
nor U24096 (N_24096,N_16013,N_17427);
and U24097 (N_24097,N_15007,N_15060);
nand U24098 (N_24098,N_16863,N_17891);
nand U24099 (N_24099,N_15419,N_19472);
and U24100 (N_24100,N_18686,N_16290);
xnor U24101 (N_24101,N_15641,N_19169);
nor U24102 (N_24102,N_19363,N_19649);
nor U24103 (N_24103,N_17874,N_18146);
or U24104 (N_24104,N_18007,N_17606);
nor U24105 (N_24105,N_17401,N_17903);
nor U24106 (N_24106,N_19782,N_17134);
or U24107 (N_24107,N_19072,N_19149);
nor U24108 (N_24108,N_18284,N_19791);
xor U24109 (N_24109,N_15952,N_19574);
or U24110 (N_24110,N_19470,N_17964);
or U24111 (N_24111,N_15003,N_16208);
nor U24112 (N_24112,N_16493,N_19317);
nand U24113 (N_24113,N_16358,N_16915);
nor U24114 (N_24114,N_19424,N_18759);
nor U24115 (N_24115,N_19543,N_16057);
nand U24116 (N_24116,N_17542,N_17676);
nor U24117 (N_24117,N_15642,N_18199);
nor U24118 (N_24118,N_18695,N_16005);
nand U24119 (N_24119,N_18259,N_19848);
and U24120 (N_24120,N_17126,N_16486);
and U24121 (N_24121,N_19944,N_15274);
and U24122 (N_24122,N_19732,N_15357);
nand U24123 (N_24123,N_18309,N_18848);
nor U24124 (N_24124,N_18260,N_17991);
nand U24125 (N_24125,N_19058,N_15330);
or U24126 (N_24126,N_17818,N_15425);
nor U24127 (N_24127,N_15408,N_19836);
or U24128 (N_24128,N_18008,N_19998);
and U24129 (N_24129,N_19356,N_18481);
or U24130 (N_24130,N_15831,N_15214);
nor U24131 (N_24131,N_19648,N_15055);
or U24132 (N_24132,N_17793,N_18123);
or U24133 (N_24133,N_18411,N_18587);
nand U24134 (N_24134,N_19923,N_15633);
or U24135 (N_24135,N_17233,N_18741);
and U24136 (N_24136,N_17019,N_19923);
and U24137 (N_24137,N_16433,N_18891);
xor U24138 (N_24138,N_16417,N_18532);
nand U24139 (N_24139,N_15275,N_15727);
and U24140 (N_24140,N_19850,N_15592);
or U24141 (N_24141,N_19271,N_19918);
nor U24142 (N_24142,N_19252,N_19982);
or U24143 (N_24143,N_15427,N_18476);
or U24144 (N_24144,N_15713,N_19497);
and U24145 (N_24145,N_19053,N_15287);
xnor U24146 (N_24146,N_16609,N_15576);
nand U24147 (N_24147,N_15310,N_18504);
nand U24148 (N_24148,N_17596,N_15836);
nand U24149 (N_24149,N_17585,N_16499);
and U24150 (N_24150,N_16568,N_15768);
or U24151 (N_24151,N_15683,N_15241);
nor U24152 (N_24152,N_18879,N_19029);
or U24153 (N_24153,N_15882,N_18553);
and U24154 (N_24154,N_19556,N_19564);
nand U24155 (N_24155,N_15173,N_17812);
nor U24156 (N_24156,N_16488,N_15449);
nand U24157 (N_24157,N_19638,N_16818);
and U24158 (N_24158,N_15550,N_19755);
or U24159 (N_24159,N_15027,N_16728);
xnor U24160 (N_24160,N_18828,N_18714);
and U24161 (N_24161,N_15427,N_15640);
nor U24162 (N_24162,N_16407,N_16027);
nand U24163 (N_24163,N_19243,N_15565);
nor U24164 (N_24164,N_15754,N_16414);
nor U24165 (N_24165,N_18861,N_17821);
xor U24166 (N_24166,N_18674,N_15587);
nor U24167 (N_24167,N_16024,N_16677);
nand U24168 (N_24168,N_18401,N_19732);
xor U24169 (N_24169,N_15711,N_18594);
or U24170 (N_24170,N_15896,N_15135);
and U24171 (N_24171,N_16793,N_19749);
and U24172 (N_24172,N_16503,N_16200);
xnor U24173 (N_24173,N_19426,N_19101);
and U24174 (N_24174,N_16491,N_17661);
nor U24175 (N_24175,N_16040,N_18073);
nand U24176 (N_24176,N_17413,N_16641);
nor U24177 (N_24177,N_16619,N_17533);
nand U24178 (N_24178,N_15749,N_18013);
or U24179 (N_24179,N_19129,N_16987);
nor U24180 (N_24180,N_16090,N_18074);
nand U24181 (N_24181,N_15882,N_18809);
and U24182 (N_24182,N_15327,N_19207);
and U24183 (N_24183,N_17579,N_17171);
or U24184 (N_24184,N_15622,N_18064);
nor U24185 (N_24185,N_16993,N_19814);
nor U24186 (N_24186,N_19642,N_18148);
nand U24187 (N_24187,N_15779,N_19085);
and U24188 (N_24188,N_18039,N_18463);
nand U24189 (N_24189,N_19909,N_19482);
nand U24190 (N_24190,N_19919,N_15096);
and U24191 (N_24191,N_15840,N_15469);
and U24192 (N_24192,N_15720,N_17265);
and U24193 (N_24193,N_18260,N_15525);
and U24194 (N_24194,N_19570,N_15260);
nor U24195 (N_24195,N_19613,N_18018);
or U24196 (N_24196,N_19138,N_17148);
nand U24197 (N_24197,N_18540,N_15008);
or U24198 (N_24198,N_17199,N_15631);
or U24199 (N_24199,N_15510,N_19777);
and U24200 (N_24200,N_16727,N_17035);
nand U24201 (N_24201,N_18019,N_19145);
and U24202 (N_24202,N_16405,N_15661);
nand U24203 (N_24203,N_18333,N_18964);
or U24204 (N_24204,N_17563,N_17204);
nand U24205 (N_24205,N_16952,N_18454);
and U24206 (N_24206,N_18739,N_19890);
or U24207 (N_24207,N_15298,N_19699);
or U24208 (N_24208,N_17895,N_18564);
nand U24209 (N_24209,N_19533,N_19763);
xor U24210 (N_24210,N_18654,N_19209);
nand U24211 (N_24211,N_17719,N_15005);
xnor U24212 (N_24212,N_17372,N_16264);
nand U24213 (N_24213,N_19414,N_18530);
or U24214 (N_24214,N_17114,N_16107);
nor U24215 (N_24215,N_15100,N_19228);
and U24216 (N_24216,N_19678,N_19806);
nand U24217 (N_24217,N_19878,N_16188);
or U24218 (N_24218,N_17447,N_19267);
and U24219 (N_24219,N_17060,N_18593);
and U24220 (N_24220,N_18636,N_19123);
or U24221 (N_24221,N_17670,N_16792);
xnor U24222 (N_24222,N_16411,N_16678);
nand U24223 (N_24223,N_15381,N_16530);
nor U24224 (N_24224,N_15048,N_17547);
or U24225 (N_24225,N_17684,N_17895);
xnor U24226 (N_24226,N_18550,N_15431);
nand U24227 (N_24227,N_19796,N_19876);
nor U24228 (N_24228,N_17115,N_17524);
nor U24229 (N_24229,N_16209,N_16214);
and U24230 (N_24230,N_18514,N_17470);
nand U24231 (N_24231,N_18465,N_15369);
and U24232 (N_24232,N_17642,N_18728);
and U24233 (N_24233,N_19208,N_19710);
and U24234 (N_24234,N_16545,N_16730);
nor U24235 (N_24235,N_16223,N_18565);
nand U24236 (N_24236,N_17621,N_19249);
nand U24237 (N_24237,N_19300,N_17478);
and U24238 (N_24238,N_17884,N_17819);
or U24239 (N_24239,N_17278,N_18594);
nor U24240 (N_24240,N_16038,N_18395);
or U24241 (N_24241,N_17874,N_17728);
nor U24242 (N_24242,N_17343,N_15860);
or U24243 (N_24243,N_18043,N_17816);
nor U24244 (N_24244,N_17266,N_17276);
nor U24245 (N_24245,N_15692,N_16842);
and U24246 (N_24246,N_19911,N_17887);
nand U24247 (N_24247,N_16120,N_19512);
nor U24248 (N_24248,N_15997,N_19791);
nor U24249 (N_24249,N_16472,N_15983);
nor U24250 (N_24250,N_18528,N_19392);
nand U24251 (N_24251,N_17385,N_17222);
or U24252 (N_24252,N_15066,N_16134);
or U24253 (N_24253,N_17003,N_18597);
nor U24254 (N_24254,N_16999,N_18969);
or U24255 (N_24255,N_15245,N_18614);
nand U24256 (N_24256,N_15679,N_17235);
or U24257 (N_24257,N_17677,N_17082);
and U24258 (N_24258,N_16907,N_16327);
and U24259 (N_24259,N_16776,N_16425);
nand U24260 (N_24260,N_16906,N_16945);
nor U24261 (N_24261,N_18407,N_19069);
and U24262 (N_24262,N_18423,N_17058);
nor U24263 (N_24263,N_15892,N_18362);
xnor U24264 (N_24264,N_19171,N_15426);
or U24265 (N_24265,N_16338,N_15897);
xor U24266 (N_24266,N_18933,N_18782);
nor U24267 (N_24267,N_19603,N_16619);
and U24268 (N_24268,N_15720,N_15506);
xnor U24269 (N_24269,N_19420,N_16379);
nand U24270 (N_24270,N_18859,N_18484);
nor U24271 (N_24271,N_15787,N_18493);
nor U24272 (N_24272,N_18594,N_18668);
nor U24273 (N_24273,N_15088,N_19450);
nor U24274 (N_24274,N_16465,N_15951);
nor U24275 (N_24275,N_18481,N_16447);
nor U24276 (N_24276,N_16965,N_17170);
and U24277 (N_24277,N_17394,N_17540);
or U24278 (N_24278,N_19557,N_19868);
nor U24279 (N_24279,N_16106,N_17295);
or U24280 (N_24280,N_18410,N_15424);
and U24281 (N_24281,N_18316,N_17255);
nor U24282 (N_24282,N_16853,N_16659);
nor U24283 (N_24283,N_18956,N_19564);
or U24284 (N_24284,N_18981,N_19146);
nand U24285 (N_24285,N_16935,N_17805);
nand U24286 (N_24286,N_16946,N_15288);
and U24287 (N_24287,N_16401,N_15877);
nor U24288 (N_24288,N_19851,N_18303);
nor U24289 (N_24289,N_15169,N_16085);
nor U24290 (N_24290,N_15340,N_19196);
and U24291 (N_24291,N_16655,N_16245);
or U24292 (N_24292,N_18271,N_16303);
xnor U24293 (N_24293,N_16171,N_15513);
and U24294 (N_24294,N_16251,N_15691);
nand U24295 (N_24295,N_19407,N_15115);
nand U24296 (N_24296,N_16135,N_19725);
nor U24297 (N_24297,N_17559,N_16212);
nor U24298 (N_24298,N_19361,N_18966);
nand U24299 (N_24299,N_15522,N_16724);
nand U24300 (N_24300,N_17438,N_19994);
nor U24301 (N_24301,N_17910,N_19639);
and U24302 (N_24302,N_18331,N_17467);
nand U24303 (N_24303,N_18427,N_19736);
nor U24304 (N_24304,N_15124,N_16768);
or U24305 (N_24305,N_16791,N_19946);
xnor U24306 (N_24306,N_18261,N_17284);
or U24307 (N_24307,N_19003,N_19056);
or U24308 (N_24308,N_18142,N_17236);
nand U24309 (N_24309,N_16130,N_15031);
nor U24310 (N_24310,N_18651,N_15523);
and U24311 (N_24311,N_18468,N_18149);
nand U24312 (N_24312,N_17765,N_16984);
nor U24313 (N_24313,N_17543,N_16382);
or U24314 (N_24314,N_18780,N_17501);
xor U24315 (N_24315,N_18533,N_17503);
nand U24316 (N_24316,N_16090,N_17559);
nand U24317 (N_24317,N_16105,N_15270);
nand U24318 (N_24318,N_17326,N_16029);
xor U24319 (N_24319,N_19020,N_19114);
nor U24320 (N_24320,N_18952,N_17211);
or U24321 (N_24321,N_16935,N_15024);
or U24322 (N_24322,N_19353,N_18038);
and U24323 (N_24323,N_16177,N_18853);
or U24324 (N_24324,N_19068,N_15863);
or U24325 (N_24325,N_19564,N_16829);
xnor U24326 (N_24326,N_15253,N_19155);
or U24327 (N_24327,N_19846,N_16131);
nor U24328 (N_24328,N_15039,N_15278);
or U24329 (N_24329,N_19283,N_17954);
or U24330 (N_24330,N_18097,N_18768);
nand U24331 (N_24331,N_17484,N_19077);
and U24332 (N_24332,N_18035,N_18010);
or U24333 (N_24333,N_18315,N_17707);
nor U24334 (N_24334,N_18984,N_17113);
and U24335 (N_24335,N_19964,N_18715);
or U24336 (N_24336,N_17228,N_18242);
nor U24337 (N_24337,N_16690,N_17100);
or U24338 (N_24338,N_18630,N_18091);
or U24339 (N_24339,N_18481,N_18697);
or U24340 (N_24340,N_17937,N_16316);
and U24341 (N_24341,N_17065,N_15825);
or U24342 (N_24342,N_18044,N_16469);
nor U24343 (N_24343,N_19905,N_16032);
xor U24344 (N_24344,N_16928,N_18160);
nor U24345 (N_24345,N_18827,N_16540);
and U24346 (N_24346,N_15865,N_15923);
and U24347 (N_24347,N_16265,N_16962);
nand U24348 (N_24348,N_19840,N_19464);
and U24349 (N_24349,N_18262,N_19560);
xor U24350 (N_24350,N_17056,N_16619);
nor U24351 (N_24351,N_16089,N_16124);
xor U24352 (N_24352,N_18385,N_16454);
nand U24353 (N_24353,N_15049,N_16740);
nor U24354 (N_24354,N_19210,N_17130);
xnor U24355 (N_24355,N_17761,N_15855);
xnor U24356 (N_24356,N_15853,N_15652);
and U24357 (N_24357,N_16043,N_17212);
and U24358 (N_24358,N_16486,N_15305);
or U24359 (N_24359,N_15367,N_15011);
and U24360 (N_24360,N_18830,N_17342);
nor U24361 (N_24361,N_18691,N_18308);
nor U24362 (N_24362,N_18817,N_16496);
nor U24363 (N_24363,N_16329,N_16359);
xnor U24364 (N_24364,N_19150,N_18201);
or U24365 (N_24365,N_19246,N_16564);
nor U24366 (N_24366,N_15362,N_19870);
or U24367 (N_24367,N_19676,N_19477);
xnor U24368 (N_24368,N_18025,N_17889);
nand U24369 (N_24369,N_15082,N_16992);
nor U24370 (N_24370,N_15521,N_15973);
nor U24371 (N_24371,N_16757,N_18033);
nor U24372 (N_24372,N_19237,N_18456);
or U24373 (N_24373,N_18895,N_16395);
nor U24374 (N_24374,N_16586,N_17761);
or U24375 (N_24375,N_17258,N_16773);
nand U24376 (N_24376,N_15110,N_15095);
and U24377 (N_24377,N_18157,N_15320);
and U24378 (N_24378,N_19124,N_19789);
nor U24379 (N_24379,N_18914,N_16193);
nand U24380 (N_24380,N_18605,N_19836);
xnor U24381 (N_24381,N_18728,N_16073);
nand U24382 (N_24382,N_15995,N_15063);
xor U24383 (N_24383,N_18761,N_19595);
nor U24384 (N_24384,N_17758,N_16816);
nor U24385 (N_24385,N_18351,N_19548);
nor U24386 (N_24386,N_15413,N_17184);
xor U24387 (N_24387,N_17396,N_18750);
nor U24388 (N_24388,N_18721,N_17116);
or U24389 (N_24389,N_18069,N_19179);
nor U24390 (N_24390,N_19171,N_15088);
xnor U24391 (N_24391,N_18668,N_18600);
nor U24392 (N_24392,N_16902,N_18553);
or U24393 (N_24393,N_16647,N_19803);
nand U24394 (N_24394,N_15360,N_15462);
and U24395 (N_24395,N_18499,N_16077);
and U24396 (N_24396,N_16829,N_17861);
and U24397 (N_24397,N_19868,N_15331);
nand U24398 (N_24398,N_16741,N_15732);
and U24399 (N_24399,N_19725,N_17973);
and U24400 (N_24400,N_16563,N_16498);
or U24401 (N_24401,N_17956,N_18668);
nand U24402 (N_24402,N_15561,N_18614);
nor U24403 (N_24403,N_15274,N_19837);
nand U24404 (N_24404,N_19647,N_16966);
nor U24405 (N_24405,N_19633,N_16659);
nor U24406 (N_24406,N_19940,N_18434);
nor U24407 (N_24407,N_16067,N_18065);
and U24408 (N_24408,N_18488,N_19972);
nand U24409 (N_24409,N_15268,N_18941);
nand U24410 (N_24410,N_17648,N_16525);
or U24411 (N_24411,N_18366,N_15819);
and U24412 (N_24412,N_15447,N_16772);
and U24413 (N_24413,N_19651,N_18217);
and U24414 (N_24414,N_19103,N_19137);
xor U24415 (N_24415,N_17718,N_16120);
nand U24416 (N_24416,N_15607,N_18935);
nand U24417 (N_24417,N_17576,N_18263);
and U24418 (N_24418,N_15480,N_16469);
and U24419 (N_24419,N_16255,N_16204);
nor U24420 (N_24420,N_15708,N_17764);
xor U24421 (N_24421,N_17982,N_18603);
or U24422 (N_24422,N_16105,N_15838);
and U24423 (N_24423,N_18983,N_15600);
nor U24424 (N_24424,N_19173,N_15569);
nand U24425 (N_24425,N_18757,N_15229);
nand U24426 (N_24426,N_17325,N_15066);
or U24427 (N_24427,N_15557,N_17389);
nand U24428 (N_24428,N_15242,N_15765);
nand U24429 (N_24429,N_18325,N_19382);
and U24430 (N_24430,N_15429,N_15321);
xnor U24431 (N_24431,N_16418,N_19218);
or U24432 (N_24432,N_15006,N_17972);
and U24433 (N_24433,N_15248,N_17568);
nor U24434 (N_24434,N_18306,N_17600);
and U24435 (N_24435,N_17268,N_19522);
or U24436 (N_24436,N_15728,N_15028);
or U24437 (N_24437,N_19520,N_15886);
or U24438 (N_24438,N_18863,N_17392);
or U24439 (N_24439,N_17770,N_18627);
nor U24440 (N_24440,N_15267,N_18131);
or U24441 (N_24441,N_15804,N_18088);
and U24442 (N_24442,N_19312,N_18398);
xor U24443 (N_24443,N_15093,N_16357);
or U24444 (N_24444,N_17669,N_16930);
nor U24445 (N_24445,N_15734,N_19581);
and U24446 (N_24446,N_16559,N_15074);
or U24447 (N_24447,N_19566,N_16278);
or U24448 (N_24448,N_18381,N_15074);
or U24449 (N_24449,N_18794,N_15850);
nor U24450 (N_24450,N_18352,N_17021);
and U24451 (N_24451,N_15792,N_15670);
nor U24452 (N_24452,N_19014,N_17119);
and U24453 (N_24453,N_18302,N_15103);
or U24454 (N_24454,N_18635,N_16191);
nor U24455 (N_24455,N_17182,N_15239);
or U24456 (N_24456,N_19959,N_18110);
and U24457 (N_24457,N_17411,N_15782);
nand U24458 (N_24458,N_19103,N_15661);
and U24459 (N_24459,N_18658,N_19843);
and U24460 (N_24460,N_19962,N_17106);
or U24461 (N_24461,N_15905,N_16654);
nand U24462 (N_24462,N_19501,N_15014);
and U24463 (N_24463,N_16926,N_19358);
xnor U24464 (N_24464,N_18437,N_18898);
nand U24465 (N_24465,N_15929,N_17906);
nor U24466 (N_24466,N_15706,N_15413);
nor U24467 (N_24467,N_19594,N_17767);
nor U24468 (N_24468,N_16213,N_19162);
nand U24469 (N_24469,N_16074,N_18895);
and U24470 (N_24470,N_15063,N_15752);
and U24471 (N_24471,N_15619,N_15506);
or U24472 (N_24472,N_19808,N_17827);
nand U24473 (N_24473,N_16532,N_15734);
xnor U24474 (N_24474,N_19714,N_16698);
nor U24475 (N_24475,N_17681,N_15958);
and U24476 (N_24476,N_15509,N_15799);
nor U24477 (N_24477,N_18825,N_19628);
or U24478 (N_24478,N_16372,N_18058);
nand U24479 (N_24479,N_18539,N_16646);
and U24480 (N_24480,N_15489,N_17627);
nor U24481 (N_24481,N_15672,N_18773);
nand U24482 (N_24482,N_15411,N_18486);
xor U24483 (N_24483,N_17618,N_19907);
nand U24484 (N_24484,N_19311,N_17294);
nor U24485 (N_24485,N_17622,N_18823);
and U24486 (N_24486,N_17821,N_15416);
nand U24487 (N_24487,N_16971,N_15352);
nand U24488 (N_24488,N_15343,N_16889);
nor U24489 (N_24489,N_16118,N_17684);
nor U24490 (N_24490,N_15277,N_18417);
and U24491 (N_24491,N_17309,N_19196);
and U24492 (N_24492,N_19004,N_16862);
xor U24493 (N_24493,N_18174,N_17067);
xnor U24494 (N_24494,N_19489,N_17380);
and U24495 (N_24495,N_17999,N_17616);
or U24496 (N_24496,N_19903,N_18032);
and U24497 (N_24497,N_15507,N_15823);
xor U24498 (N_24498,N_17481,N_19161);
xor U24499 (N_24499,N_15116,N_19473);
or U24500 (N_24500,N_19176,N_16369);
and U24501 (N_24501,N_18941,N_19016);
nand U24502 (N_24502,N_16681,N_15447);
and U24503 (N_24503,N_15215,N_19533);
or U24504 (N_24504,N_17436,N_16994);
and U24505 (N_24505,N_19862,N_19799);
nand U24506 (N_24506,N_17256,N_17077);
or U24507 (N_24507,N_19254,N_19960);
or U24508 (N_24508,N_17510,N_17604);
or U24509 (N_24509,N_19322,N_16921);
nor U24510 (N_24510,N_17347,N_16370);
nand U24511 (N_24511,N_15890,N_15515);
nand U24512 (N_24512,N_17824,N_15296);
or U24513 (N_24513,N_16532,N_18746);
nor U24514 (N_24514,N_19750,N_18516);
nand U24515 (N_24515,N_17549,N_15013);
nand U24516 (N_24516,N_18090,N_16151);
xnor U24517 (N_24517,N_17866,N_17400);
or U24518 (N_24518,N_18019,N_15588);
nand U24519 (N_24519,N_17629,N_15912);
or U24520 (N_24520,N_18287,N_17594);
nand U24521 (N_24521,N_19796,N_18283);
and U24522 (N_24522,N_17906,N_15641);
nor U24523 (N_24523,N_16007,N_17295);
xor U24524 (N_24524,N_19070,N_18242);
xor U24525 (N_24525,N_16780,N_19603);
nand U24526 (N_24526,N_18653,N_18451);
or U24527 (N_24527,N_19720,N_17980);
or U24528 (N_24528,N_15128,N_15094);
nor U24529 (N_24529,N_17715,N_15616);
or U24530 (N_24530,N_15632,N_18023);
and U24531 (N_24531,N_17372,N_17203);
nand U24532 (N_24532,N_18063,N_17609);
xor U24533 (N_24533,N_19132,N_19582);
and U24534 (N_24534,N_18606,N_15181);
or U24535 (N_24535,N_16494,N_17308);
or U24536 (N_24536,N_19048,N_15427);
and U24537 (N_24537,N_17327,N_19165);
xnor U24538 (N_24538,N_15343,N_17864);
or U24539 (N_24539,N_16653,N_19714);
or U24540 (N_24540,N_15815,N_19252);
and U24541 (N_24541,N_19309,N_15125);
xnor U24542 (N_24542,N_19710,N_18936);
nand U24543 (N_24543,N_16652,N_19072);
nor U24544 (N_24544,N_17588,N_17151);
and U24545 (N_24545,N_16348,N_19988);
and U24546 (N_24546,N_16179,N_16383);
nand U24547 (N_24547,N_18816,N_19016);
or U24548 (N_24548,N_16055,N_15182);
or U24549 (N_24549,N_18918,N_16309);
nand U24550 (N_24550,N_18764,N_15223);
and U24551 (N_24551,N_18207,N_19373);
and U24552 (N_24552,N_17421,N_16512);
or U24553 (N_24553,N_19636,N_18934);
nor U24554 (N_24554,N_16481,N_16776);
nand U24555 (N_24555,N_19881,N_16951);
or U24556 (N_24556,N_15119,N_19711);
nand U24557 (N_24557,N_15962,N_19712);
or U24558 (N_24558,N_19927,N_19504);
nand U24559 (N_24559,N_16419,N_19386);
or U24560 (N_24560,N_18899,N_18569);
nor U24561 (N_24561,N_18227,N_19094);
nand U24562 (N_24562,N_18017,N_15586);
nand U24563 (N_24563,N_16180,N_17240);
nand U24564 (N_24564,N_19655,N_15536);
nor U24565 (N_24565,N_18917,N_18579);
xnor U24566 (N_24566,N_17801,N_18568);
nand U24567 (N_24567,N_16848,N_19845);
nand U24568 (N_24568,N_15325,N_18228);
and U24569 (N_24569,N_19148,N_16739);
or U24570 (N_24570,N_17220,N_18114);
or U24571 (N_24571,N_19342,N_15003);
and U24572 (N_24572,N_15644,N_15456);
nand U24573 (N_24573,N_18134,N_15530);
or U24574 (N_24574,N_17751,N_19274);
nand U24575 (N_24575,N_18894,N_15171);
xor U24576 (N_24576,N_17960,N_18935);
nor U24577 (N_24577,N_15568,N_17271);
or U24578 (N_24578,N_17105,N_19907);
and U24579 (N_24579,N_16578,N_18663);
or U24580 (N_24580,N_19874,N_16723);
nor U24581 (N_24581,N_15778,N_16556);
nor U24582 (N_24582,N_18164,N_18303);
nand U24583 (N_24583,N_18194,N_17866);
nor U24584 (N_24584,N_17693,N_15526);
xor U24585 (N_24585,N_15930,N_15424);
xor U24586 (N_24586,N_15230,N_16403);
nor U24587 (N_24587,N_15631,N_19862);
or U24588 (N_24588,N_16549,N_18852);
nand U24589 (N_24589,N_18536,N_15004);
nor U24590 (N_24590,N_17824,N_18884);
and U24591 (N_24591,N_18651,N_15832);
xor U24592 (N_24592,N_16437,N_16699);
or U24593 (N_24593,N_17693,N_19549);
or U24594 (N_24594,N_15467,N_17883);
or U24595 (N_24595,N_19866,N_18749);
or U24596 (N_24596,N_17577,N_15483);
and U24597 (N_24597,N_19376,N_17800);
xor U24598 (N_24598,N_19095,N_16704);
or U24599 (N_24599,N_18234,N_18272);
and U24600 (N_24600,N_15629,N_15379);
xnor U24601 (N_24601,N_16403,N_18660);
xnor U24602 (N_24602,N_15467,N_19766);
and U24603 (N_24603,N_19244,N_17826);
or U24604 (N_24604,N_18894,N_17598);
nand U24605 (N_24605,N_17919,N_18553);
nand U24606 (N_24606,N_15710,N_19733);
and U24607 (N_24607,N_16303,N_18819);
nand U24608 (N_24608,N_18894,N_19938);
xnor U24609 (N_24609,N_16270,N_15955);
or U24610 (N_24610,N_18287,N_16689);
or U24611 (N_24611,N_16610,N_19654);
or U24612 (N_24612,N_19417,N_17069);
xor U24613 (N_24613,N_15171,N_18282);
nor U24614 (N_24614,N_18084,N_15394);
and U24615 (N_24615,N_17712,N_17946);
nand U24616 (N_24616,N_15565,N_15948);
and U24617 (N_24617,N_19723,N_16259);
nor U24618 (N_24618,N_16785,N_15883);
nand U24619 (N_24619,N_17717,N_17400);
or U24620 (N_24620,N_17080,N_19149);
and U24621 (N_24621,N_15674,N_19096);
or U24622 (N_24622,N_17953,N_16386);
and U24623 (N_24623,N_16841,N_18278);
and U24624 (N_24624,N_15778,N_19180);
or U24625 (N_24625,N_15712,N_19229);
and U24626 (N_24626,N_18357,N_19656);
nor U24627 (N_24627,N_16449,N_17541);
and U24628 (N_24628,N_19308,N_19120);
nand U24629 (N_24629,N_18490,N_17591);
and U24630 (N_24630,N_16814,N_15842);
nor U24631 (N_24631,N_18505,N_19471);
nand U24632 (N_24632,N_17342,N_19053);
nand U24633 (N_24633,N_16258,N_18516);
nor U24634 (N_24634,N_19323,N_19268);
or U24635 (N_24635,N_17411,N_15049);
xnor U24636 (N_24636,N_17251,N_17049);
or U24637 (N_24637,N_19667,N_16396);
and U24638 (N_24638,N_18346,N_18109);
or U24639 (N_24639,N_16386,N_16858);
nor U24640 (N_24640,N_16804,N_18918);
nor U24641 (N_24641,N_15078,N_19429);
or U24642 (N_24642,N_19985,N_16009);
nand U24643 (N_24643,N_17853,N_17905);
or U24644 (N_24644,N_16814,N_17958);
nand U24645 (N_24645,N_16400,N_19282);
nor U24646 (N_24646,N_19875,N_15122);
nand U24647 (N_24647,N_16826,N_18553);
xnor U24648 (N_24648,N_18017,N_18911);
nand U24649 (N_24649,N_15263,N_16151);
nor U24650 (N_24650,N_18918,N_16674);
and U24651 (N_24651,N_19111,N_16988);
and U24652 (N_24652,N_16337,N_19237);
or U24653 (N_24653,N_17828,N_16178);
or U24654 (N_24654,N_16954,N_16767);
and U24655 (N_24655,N_16780,N_16293);
xor U24656 (N_24656,N_16033,N_19842);
and U24657 (N_24657,N_17340,N_19856);
or U24658 (N_24658,N_18097,N_16936);
and U24659 (N_24659,N_18922,N_17844);
or U24660 (N_24660,N_16687,N_16683);
xnor U24661 (N_24661,N_17644,N_18630);
and U24662 (N_24662,N_19918,N_17322);
and U24663 (N_24663,N_19430,N_17429);
or U24664 (N_24664,N_16221,N_19346);
nor U24665 (N_24665,N_18856,N_17592);
xor U24666 (N_24666,N_16073,N_15364);
or U24667 (N_24667,N_16412,N_15082);
and U24668 (N_24668,N_18483,N_19140);
and U24669 (N_24669,N_18397,N_17913);
nor U24670 (N_24670,N_15739,N_15693);
or U24671 (N_24671,N_16674,N_15540);
and U24672 (N_24672,N_19442,N_15467);
xnor U24673 (N_24673,N_15735,N_17827);
nand U24674 (N_24674,N_19578,N_15924);
nor U24675 (N_24675,N_17517,N_15250);
and U24676 (N_24676,N_19578,N_19564);
nor U24677 (N_24677,N_19636,N_16694);
xnor U24678 (N_24678,N_16915,N_17374);
and U24679 (N_24679,N_16982,N_16661);
or U24680 (N_24680,N_19599,N_17398);
nor U24681 (N_24681,N_18081,N_19011);
xor U24682 (N_24682,N_15950,N_15672);
nand U24683 (N_24683,N_18140,N_19673);
nand U24684 (N_24684,N_15217,N_19099);
or U24685 (N_24685,N_17288,N_19044);
or U24686 (N_24686,N_18055,N_19785);
xnor U24687 (N_24687,N_17255,N_18770);
and U24688 (N_24688,N_16250,N_17648);
nor U24689 (N_24689,N_18807,N_17214);
or U24690 (N_24690,N_18746,N_19216);
and U24691 (N_24691,N_17466,N_16885);
nor U24692 (N_24692,N_18179,N_16742);
and U24693 (N_24693,N_16647,N_17137);
and U24694 (N_24694,N_17064,N_19728);
nor U24695 (N_24695,N_15345,N_18470);
xnor U24696 (N_24696,N_17347,N_16856);
nor U24697 (N_24697,N_18839,N_18883);
or U24698 (N_24698,N_16081,N_18986);
xor U24699 (N_24699,N_16018,N_17348);
nand U24700 (N_24700,N_15199,N_19089);
and U24701 (N_24701,N_15403,N_17092);
nor U24702 (N_24702,N_17021,N_15809);
nand U24703 (N_24703,N_17642,N_16476);
or U24704 (N_24704,N_19045,N_15389);
nor U24705 (N_24705,N_19773,N_16815);
nor U24706 (N_24706,N_19163,N_17859);
or U24707 (N_24707,N_19396,N_16350);
or U24708 (N_24708,N_19576,N_16038);
and U24709 (N_24709,N_17157,N_19791);
and U24710 (N_24710,N_18681,N_15986);
nand U24711 (N_24711,N_19496,N_17808);
xor U24712 (N_24712,N_18080,N_19543);
nand U24713 (N_24713,N_15382,N_18594);
nor U24714 (N_24714,N_19832,N_18207);
xnor U24715 (N_24715,N_18427,N_17257);
and U24716 (N_24716,N_18065,N_18485);
and U24717 (N_24717,N_17725,N_16770);
xor U24718 (N_24718,N_16548,N_19378);
or U24719 (N_24719,N_18003,N_18339);
nor U24720 (N_24720,N_19378,N_16180);
nor U24721 (N_24721,N_15739,N_19973);
and U24722 (N_24722,N_16975,N_16870);
or U24723 (N_24723,N_17025,N_17067);
nor U24724 (N_24724,N_19264,N_16927);
and U24725 (N_24725,N_15400,N_15488);
and U24726 (N_24726,N_18475,N_15578);
and U24727 (N_24727,N_19356,N_17045);
xnor U24728 (N_24728,N_16495,N_17199);
and U24729 (N_24729,N_15095,N_16115);
nand U24730 (N_24730,N_16586,N_16710);
and U24731 (N_24731,N_16433,N_15997);
and U24732 (N_24732,N_19698,N_15031);
or U24733 (N_24733,N_15816,N_19365);
nand U24734 (N_24734,N_15996,N_19291);
nor U24735 (N_24735,N_19520,N_17631);
nor U24736 (N_24736,N_17204,N_18406);
and U24737 (N_24737,N_16759,N_18667);
xnor U24738 (N_24738,N_18036,N_16509);
or U24739 (N_24739,N_18835,N_18902);
nand U24740 (N_24740,N_18859,N_19002);
nand U24741 (N_24741,N_17691,N_19291);
or U24742 (N_24742,N_17728,N_18869);
nand U24743 (N_24743,N_17343,N_19132);
nand U24744 (N_24744,N_19782,N_19926);
nand U24745 (N_24745,N_17423,N_15417);
nor U24746 (N_24746,N_15942,N_16451);
or U24747 (N_24747,N_19676,N_17682);
or U24748 (N_24748,N_17561,N_18153);
nor U24749 (N_24749,N_19543,N_15112);
and U24750 (N_24750,N_15372,N_17723);
nor U24751 (N_24751,N_15296,N_18708);
nor U24752 (N_24752,N_18834,N_19031);
xnor U24753 (N_24753,N_18003,N_19486);
nor U24754 (N_24754,N_18989,N_19982);
nor U24755 (N_24755,N_18053,N_16843);
or U24756 (N_24756,N_16251,N_19512);
nor U24757 (N_24757,N_18514,N_16344);
or U24758 (N_24758,N_17790,N_16926);
nor U24759 (N_24759,N_19778,N_18584);
and U24760 (N_24760,N_18639,N_17863);
or U24761 (N_24761,N_15175,N_17077);
nand U24762 (N_24762,N_16692,N_15154);
xnor U24763 (N_24763,N_19215,N_16474);
xor U24764 (N_24764,N_19648,N_18078);
and U24765 (N_24765,N_18404,N_15830);
xnor U24766 (N_24766,N_17203,N_16464);
nor U24767 (N_24767,N_18009,N_15623);
nand U24768 (N_24768,N_15122,N_19987);
and U24769 (N_24769,N_15745,N_19197);
nor U24770 (N_24770,N_15549,N_19492);
nor U24771 (N_24771,N_15487,N_15210);
or U24772 (N_24772,N_19019,N_18461);
or U24773 (N_24773,N_19522,N_17536);
and U24774 (N_24774,N_17652,N_15281);
or U24775 (N_24775,N_17452,N_18940);
nor U24776 (N_24776,N_19933,N_19877);
nand U24777 (N_24777,N_18083,N_16215);
or U24778 (N_24778,N_15230,N_19339);
and U24779 (N_24779,N_15678,N_19827);
or U24780 (N_24780,N_15814,N_16379);
nand U24781 (N_24781,N_15872,N_15328);
nand U24782 (N_24782,N_16160,N_17587);
nor U24783 (N_24783,N_18643,N_16491);
or U24784 (N_24784,N_16614,N_17322);
and U24785 (N_24785,N_17522,N_19032);
and U24786 (N_24786,N_16749,N_18230);
and U24787 (N_24787,N_15837,N_15333);
nor U24788 (N_24788,N_18723,N_17558);
or U24789 (N_24789,N_19012,N_18792);
nand U24790 (N_24790,N_15093,N_18128);
nor U24791 (N_24791,N_17547,N_19580);
nor U24792 (N_24792,N_16683,N_19724);
nand U24793 (N_24793,N_17468,N_19608);
xor U24794 (N_24794,N_18917,N_17691);
xor U24795 (N_24795,N_16213,N_17441);
nand U24796 (N_24796,N_15286,N_19012);
xor U24797 (N_24797,N_17714,N_16667);
or U24798 (N_24798,N_19662,N_15074);
or U24799 (N_24799,N_18595,N_19682);
nor U24800 (N_24800,N_19130,N_17130);
xor U24801 (N_24801,N_18148,N_18732);
or U24802 (N_24802,N_15772,N_18652);
nand U24803 (N_24803,N_19673,N_16714);
nor U24804 (N_24804,N_16929,N_16568);
nor U24805 (N_24805,N_19861,N_16727);
nand U24806 (N_24806,N_16886,N_18738);
nor U24807 (N_24807,N_17688,N_16445);
nor U24808 (N_24808,N_19129,N_19172);
and U24809 (N_24809,N_16426,N_19148);
and U24810 (N_24810,N_18328,N_18825);
nand U24811 (N_24811,N_15604,N_15633);
nor U24812 (N_24812,N_17120,N_15614);
and U24813 (N_24813,N_17256,N_19402);
and U24814 (N_24814,N_19622,N_18589);
nor U24815 (N_24815,N_16337,N_15439);
nand U24816 (N_24816,N_18270,N_17848);
nand U24817 (N_24817,N_18844,N_15386);
or U24818 (N_24818,N_18288,N_15340);
nand U24819 (N_24819,N_19238,N_19283);
or U24820 (N_24820,N_18187,N_16462);
nor U24821 (N_24821,N_19024,N_15683);
and U24822 (N_24822,N_16725,N_16031);
nand U24823 (N_24823,N_18951,N_18003);
nand U24824 (N_24824,N_17288,N_19363);
and U24825 (N_24825,N_16471,N_19747);
nand U24826 (N_24826,N_15170,N_18601);
or U24827 (N_24827,N_19459,N_15537);
or U24828 (N_24828,N_15434,N_17487);
nand U24829 (N_24829,N_19867,N_17783);
and U24830 (N_24830,N_18896,N_16586);
nor U24831 (N_24831,N_16174,N_18584);
and U24832 (N_24832,N_16561,N_19362);
nor U24833 (N_24833,N_16571,N_15728);
or U24834 (N_24834,N_16349,N_15652);
and U24835 (N_24835,N_18364,N_17365);
xor U24836 (N_24836,N_19445,N_18372);
or U24837 (N_24837,N_19619,N_18564);
or U24838 (N_24838,N_15443,N_17252);
nand U24839 (N_24839,N_18528,N_18338);
nand U24840 (N_24840,N_15441,N_15508);
nor U24841 (N_24841,N_17089,N_16361);
and U24842 (N_24842,N_18451,N_15997);
nor U24843 (N_24843,N_18256,N_17260);
nor U24844 (N_24844,N_19910,N_15131);
nor U24845 (N_24845,N_16781,N_17166);
and U24846 (N_24846,N_17786,N_18443);
nor U24847 (N_24847,N_19365,N_17545);
xor U24848 (N_24848,N_15003,N_17559);
xnor U24849 (N_24849,N_17459,N_19583);
nand U24850 (N_24850,N_19283,N_19333);
and U24851 (N_24851,N_19589,N_15826);
or U24852 (N_24852,N_17916,N_19672);
nor U24853 (N_24853,N_19457,N_15465);
nor U24854 (N_24854,N_19167,N_16202);
nand U24855 (N_24855,N_19383,N_19561);
nand U24856 (N_24856,N_15497,N_19461);
nand U24857 (N_24857,N_15814,N_18353);
and U24858 (N_24858,N_16882,N_16195);
or U24859 (N_24859,N_17908,N_16212);
or U24860 (N_24860,N_17240,N_16781);
nand U24861 (N_24861,N_17379,N_18393);
nand U24862 (N_24862,N_16324,N_19025);
or U24863 (N_24863,N_18426,N_19892);
or U24864 (N_24864,N_17772,N_19361);
nor U24865 (N_24865,N_16456,N_17808);
and U24866 (N_24866,N_15318,N_15701);
nor U24867 (N_24867,N_17376,N_17824);
and U24868 (N_24868,N_16151,N_17236);
xor U24869 (N_24869,N_17982,N_15223);
nor U24870 (N_24870,N_17109,N_15994);
or U24871 (N_24871,N_19446,N_19841);
nand U24872 (N_24872,N_17303,N_17789);
nand U24873 (N_24873,N_17912,N_19399);
and U24874 (N_24874,N_18786,N_17247);
and U24875 (N_24875,N_15181,N_18468);
nor U24876 (N_24876,N_17169,N_18543);
or U24877 (N_24877,N_18318,N_18249);
and U24878 (N_24878,N_17293,N_19663);
xor U24879 (N_24879,N_17642,N_18272);
and U24880 (N_24880,N_15225,N_19826);
nor U24881 (N_24881,N_18386,N_17060);
or U24882 (N_24882,N_19414,N_15245);
nand U24883 (N_24883,N_19584,N_16042);
nor U24884 (N_24884,N_18479,N_19388);
or U24885 (N_24885,N_18531,N_18568);
nand U24886 (N_24886,N_19892,N_18170);
or U24887 (N_24887,N_16317,N_16622);
nor U24888 (N_24888,N_15428,N_19280);
xor U24889 (N_24889,N_19129,N_18342);
xnor U24890 (N_24890,N_16612,N_15527);
nand U24891 (N_24891,N_17565,N_18156);
nor U24892 (N_24892,N_17341,N_15611);
nand U24893 (N_24893,N_19638,N_15119);
xor U24894 (N_24894,N_17204,N_15398);
nor U24895 (N_24895,N_18428,N_18800);
or U24896 (N_24896,N_17764,N_16011);
nand U24897 (N_24897,N_17248,N_19522);
or U24898 (N_24898,N_18663,N_15018);
and U24899 (N_24899,N_15715,N_18114);
or U24900 (N_24900,N_18462,N_18243);
xor U24901 (N_24901,N_18101,N_16034);
nor U24902 (N_24902,N_17825,N_16701);
and U24903 (N_24903,N_18175,N_15345);
nor U24904 (N_24904,N_16207,N_15124);
nor U24905 (N_24905,N_19694,N_15944);
or U24906 (N_24906,N_16846,N_15635);
and U24907 (N_24907,N_15741,N_18041);
xnor U24908 (N_24908,N_19543,N_18142);
nor U24909 (N_24909,N_17674,N_16099);
xor U24910 (N_24910,N_17197,N_19029);
nor U24911 (N_24911,N_18342,N_17586);
or U24912 (N_24912,N_17720,N_17263);
nand U24913 (N_24913,N_16241,N_15847);
or U24914 (N_24914,N_16753,N_16081);
nand U24915 (N_24915,N_16725,N_16001);
or U24916 (N_24916,N_15624,N_19944);
and U24917 (N_24917,N_15653,N_19597);
nand U24918 (N_24918,N_18542,N_17013);
and U24919 (N_24919,N_17514,N_17858);
nand U24920 (N_24920,N_18334,N_15104);
and U24921 (N_24921,N_17996,N_15058);
nor U24922 (N_24922,N_15644,N_15223);
or U24923 (N_24923,N_15891,N_18344);
xnor U24924 (N_24924,N_19561,N_19298);
and U24925 (N_24925,N_17411,N_18182);
or U24926 (N_24926,N_19422,N_19929);
and U24927 (N_24927,N_18692,N_18426);
xor U24928 (N_24928,N_18273,N_19805);
or U24929 (N_24929,N_15424,N_16096);
and U24930 (N_24930,N_18983,N_15254);
nand U24931 (N_24931,N_16765,N_19175);
nand U24932 (N_24932,N_18360,N_15273);
nor U24933 (N_24933,N_17004,N_16951);
and U24934 (N_24934,N_19910,N_18247);
or U24935 (N_24935,N_19845,N_18539);
and U24936 (N_24936,N_18807,N_19099);
nand U24937 (N_24937,N_18569,N_15336);
nand U24938 (N_24938,N_16454,N_17809);
nor U24939 (N_24939,N_16536,N_19007);
nor U24940 (N_24940,N_15782,N_16687);
nand U24941 (N_24941,N_19054,N_15664);
or U24942 (N_24942,N_17845,N_19008);
and U24943 (N_24943,N_19666,N_16762);
xor U24944 (N_24944,N_15483,N_18142);
nand U24945 (N_24945,N_15375,N_18434);
or U24946 (N_24946,N_16563,N_15868);
nor U24947 (N_24947,N_17310,N_17209);
nand U24948 (N_24948,N_17735,N_16752);
xnor U24949 (N_24949,N_18195,N_16027);
nor U24950 (N_24950,N_19500,N_19595);
and U24951 (N_24951,N_18897,N_17868);
nand U24952 (N_24952,N_17476,N_16314);
and U24953 (N_24953,N_16956,N_19862);
nor U24954 (N_24954,N_15757,N_16212);
nand U24955 (N_24955,N_17061,N_17320);
and U24956 (N_24956,N_15444,N_18200);
or U24957 (N_24957,N_17521,N_15642);
nor U24958 (N_24958,N_18283,N_15908);
or U24959 (N_24959,N_16270,N_18485);
nor U24960 (N_24960,N_15664,N_18313);
nand U24961 (N_24961,N_15018,N_18179);
or U24962 (N_24962,N_17261,N_16027);
xnor U24963 (N_24963,N_16729,N_19701);
nand U24964 (N_24964,N_19996,N_17612);
nand U24965 (N_24965,N_17465,N_16435);
and U24966 (N_24966,N_16638,N_16644);
nor U24967 (N_24967,N_19398,N_16412);
or U24968 (N_24968,N_18172,N_16223);
and U24969 (N_24969,N_18215,N_17809);
or U24970 (N_24970,N_16923,N_15142);
and U24971 (N_24971,N_18612,N_18576);
nor U24972 (N_24972,N_17198,N_18649);
xnor U24973 (N_24973,N_17945,N_15301);
and U24974 (N_24974,N_19206,N_18531);
and U24975 (N_24975,N_19681,N_19042);
nand U24976 (N_24976,N_19056,N_18279);
and U24977 (N_24977,N_15187,N_15854);
and U24978 (N_24978,N_17532,N_15480);
nand U24979 (N_24979,N_17584,N_17748);
or U24980 (N_24980,N_17777,N_16039);
nor U24981 (N_24981,N_16330,N_16883);
or U24982 (N_24982,N_19719,N_18437);
nor U24983 (N_24983,N_19448,N_16895);
or U24984 (N_24984,N_17691,N_19258);
nand U24985 (N_24985,N_15978,N_17982);
nor U24986 (N_24986,N_15066,N_19150);
or U24987 (N_24987,N_19537,N_18114);
nor U24988 (N_24988,N_15372,N_17054);
and U24989 (N_24989,N_17221,N_17072);
nand U24990 (N_24990,N_16675,N_16805);
or U24991 (N_24991,N_18247,N_17165);
nand U24992 (N_24992,N_18284,N_15129);
nor U24993 (N_24993,N_15787,N_16832);
nand U24994 (N_24994,N_17107,N_15731);
and U24995 (N_24995,N_18915,N_16816);
nand U24996 (N_24996,N_15567,N_18962);
and U24997 (N_24997,N_17552,N_18858);
nand U24998 (N_24998,N_16859,N_18127);
or U24999 (N_24999,N_18824,N_15618);
or UO_0 (O_0,N_23586,N_20997);
and UO_1 (O_1,N_23271,N_24546);
xnor UO_2 (O_2,N_24222,N_21736);
nor UO_3 (O_3,N_23072,N_20840);
and UO_4 (O_4,N_22394,N_20079);
and UO_5 (O_5,N_24143,N_24949);
nor UO_6 (O_6,N_23153,N_22165);
xnor UO_7 (O_7,N_24590,N_22915);
and UO_8 (O_8,N_21885,N_23777);
nand UO_9 (O_9,N_23490,N_21690);
nand UO_10 (O_10,N_23049,N_21727);
nand UO_11 (O_11,N_22121,N_22067);
nor UO_12 (O_12,N_24536,N_20062);
or UO_13 (O_13,N_22535,N_22494);
nand UO_14 (O_14,N_23390,N_24470);
xor UO_15 (O_15,N_23581,N_20090);
and UO_16 (O_16,N_20581,N_22061);
nor UO_17 (O_17,N_21732,N_23065);
and UO_18 (O_18,N_22589,N_20452);
or UO_19 (O_19,N_24390,N_23639);
xnor UO_20 (O_20,N_20702,N_22885);
or UO_21 (O_21,N_24419,N_24057);
nor UO_22 (O_22,N_22795,N_22235);
nor UO_23 (O_23,N_21128,N_22540);
and UO_24 (O_24,N_23740,N_23852);
nand UO_25 (O_25,N_21189,N_23602);
and UO_26 (O_26,N_23019,N_20797);
nand UO_27 (O_27,N_23967,N_20593);
nand UO_28 (O_28,N_20824,N_22723);
and UO_29 (O_29,N_22766,N_23656);
and UO_30 (O_30,N_22192,N_22601);
or UO_31 (O_31,N_21823,N_20028);
or UO_32 (O_32,N_22046,N_23815);
and UO_33 (O_33,N_20891,N_23022);
or UO_34 (O_34,N_20564,N_24811);
nor UO_35 (O_35,N_21996,N_22991);
nand UO_36 (O_36,N_23349,N_23520);
nand UO_37 (O_37,N_20063,N_20269);
and UO_38 (O_38,N_23386,N_23159);
nand UO_39 (O_39,N_22842,N_21509);
nand UO_40 (O_40,N_21891,N_22246);
or UO_41 (O_41,N_20472,N_22947);
nand UO_42 (O_42,N_20537,N_24982);
nor UO_43 (O_43,N_21484,N_24541);
and UO_44 (O_44,N_22602,N_21036);
nor UO_45 (O_45,N_21474,N_22075);
nand UO_46 (O_46,N_22223,N_21227);
nor UO_47 (O_47,N_22533,N_21300);
nor UO_48 (O_48,N_24122,N_23273);
nand UO_49 (O_49,N_22399,N_20332);
xnor UO_50 (O_50,N_24463,N_22379);
and UO_51 (O_51,N_24679,N_22683);
and UO_52 (O_52,N_24499,N_21062);
nor UO_53 (O_53,N_22008,N_22553);
and UO_54 (O_54,N_24738,N_21490);
nand UO_55 (O_55,N_24260,N_22921);
nor UO_56 (O_56,N_21115,N_20083);
nor UO_57 (O_57,N_20590,N_23513);
and UO_58 (O_58,N_20507,N_21763);
and UO_59 (O_59,N_23703,N_23674);
and UO_60 (O_60,N_22346,N_21604);
and UO_61 (O_61,N_23766,N_24598);
nor UO_62 (O_62,N_21129,N_21684);
or UO_63 (O_63,N_22467,N_20831);
nor UO_64 (O_64,N_20397,N_24686);
and UO_65 (O_65,N_20599,N_20610);
nand UO_66 (O_66,N_23610,N_22867);
and UO_67 (O_67,N_23128,N_23201);
and UO_68 (O_68,N_22303,N_20247);
nor UO_69 (O_69,N_23326,N_23872);
nor UO_70 (O_70,N_21724,N_21100);
xor UO_71 (O_71,N_23406,N_20953);
and UO_72 (O_72,N_22083,N_24589);
and UO_73 (O_73,N_24531,N_23700);
xnor UO_74 (O_74,N_20221,N_20485);
and UO_75 (O_75,N_20033,N_22363);
and UO_76 (O_76,N_20329,N_24415);
and UO_77 (O_77,N_21901,N_23214);
xnor UO_78 (O_78,N_21091,N_21913);
or UO_79 (O_79,N_21775,N_21912);
or UO_80 (O_80,N_22471,N_21893);
nand UO_81 (O_81,N_24902,N_23184);
or UO_82 (O_82,N_24066,N_24530);
nand UO_83 (O_83,N_22318,N_21845);
or UO_84 (O_84,N_23257,N_21550);
xnor UO_85 (O_85,N_24860,N_20771);
nand UO_86 (O_86,N_22884,N_23997);
or UO_87 (O_87,N_22018,N_22052);
nand UO_88 (O_88,N_23464,N_21401);
xnor UO_89 (O_89,N_23278,N_22485);
nand UO_90 (O_90,N_23607,N_21756);
nand UO_91 (O_91,N_22116,N_22653);
nor UO_92 (O_92,N_22955,N_23736);
nand UO_93 (O_93,N_20732,N_23532);
and UO_94 (O_94,N_24696,N_21804);
xor UO_95 (O_95,N_24177,N_23922);
nor UO_96 (O_96,N_23626,N_21077);
nand UO_97 (O_97,N_22755,N_20961);
xnor UO_98 (O_98,N_22712,N_21295);
nand UO_99 (O_99,N_21282,N_20100);
nor UO_100 (O_100,N_20143,N_21641);
nor UO_101 (O_101,N_20074,N_23901);
or UO_102 (O_102,N_22605,N_21579);
nand UO_103 (O_103,N_20520,N_20381);
nor UO_104 (O_104,N_23623,N_23794);
and UO_105 (O_105,N_23372,N_23804);
or UO_106 (O_106,N_23891,N_21393);
nand UO_107 (O_107,N_22393,N_20451);
nor UO_108 (O_108,N_21387,N_24987);
or UO_109 (O_109,N_21795,N_22742);
or UO_110 (O_110,N_22942,N_24295);
nand UO_111 (O_111,N_21687,N_24138);
or UO_112 (O_112,N_20570,N_23016);
nor UO_113 (O_113,N_24034,N_21975);
or UO_114 (O_114,N_24911,N_22304);
and UO_115 (O_115,N_23946,N_24535);
and UO_116 (O_116,N_21275,N_20113);
xnor UO_117 (O_117,N_21710,N_20572);
xor UO_118 (O_118,N_22087,N_21962);
and UO_119 (O_119,N_20245,N_21935);
nand UO_120 (O_120,N_22201,N_24141);
and UO_121 (O_121,N_21224,N_24282);
nor UO_122 (O_122,N_20653,N_21750);
or UO_123 (O_123,N_22213,N_23954);
and UO_124 (O_124,N_22846,N_21553);
nand UO_125 (O_125,N_22954,N_24398);
and UO_126 (O_126,N_24191,N_21574);
and UO_127 (O_127,N_22866,N_24578);
nor UO_128 (O_128,N_23751,N_24553);
nand UO_129 (O_129,N_21050,N_20377);
or UO_130 (O_130,N_20528,N_24970);
nor UO_131 (O_131,N_21336,N_24056);
or UO_132 (O_132,N_20493,N_24343);
nand UO_133 (O_133,N_21590,N_23113);
or UO_134 (O_134,N_24897,N_23653);
nor UO_135 (O_135,N_20740,N_20985);
xnor UO_136 (O_136,N_21977,N_24550);
nor UO_137 (O_137,N_21925,N_23523);
and UO_138 (O_138,N_21917,N_23886);
or UO_139 (O_139,N_23732,N_23709);
and UO_140 (O_140,N_24431,N_21086);
nor UO_141 (O_141,N_21456,N_23324);
or UO_142 (O_142,N_20170,N_22319);
nor UO_143 (O_143,N_22076,N_22437);
nor UO_144 (O_144,N_20688,N_23568);
or UO_145 (O_145,N_23043,N_21928);
nand UO_146 (O_146,N_20384,N_23525);
xor UO_147 (O_147,N_23690,N_24663);
nand UO_148 (O_148,N_22349,N_22935);
nor UO_149 (O_149,N_22042,N_23827);
xor UO_150 (O_150,N_23663,N_24921);
nand UO_151 (O_151,N_23236,N_24942);
nor UO_152 (O_152,N_24132,N_21015);
and UO_153 (O_153,N_24196,N_21449);
and UO_154 (O_154,N_22517,N_21647);
or UO_155 (O_155,N_23232,N_24784);
nor UO_156 (O_156,N_21890,N_23823);
nand UO_157 (O_157,N_22300,N_23472);
and UO_158 (O_158,N_23144,N_21668);
nand UO_159 (O_159,N_21476,N_24235);
xnor UO_160 (O_160,N_23512,N_21356);
and UO_161 (O_161,N_20934,N_23105);
nor UO_162 (O_162,N_24330,N_23156);
nand UO_163 (O_163,N_21450,N_20005);
xor UO_164 (O_164,N_24585,N_20408);
or UO_165 (O_165,N_21454,N_24417);
and UO_166 (O_166,N_21184,N_23231);
xor UO_167 (O_167,N_22629,N_21020);
and UO_168 (O_168,N_24665,N_24651);
or UO_169 (O_169,N_20299,N_24610);
and UO_170 (O_170,N_22030,N_23408);
nand UO_171 (O_171,N_21675,N_22093);
or UO_172 (O_172,N_23252,N_24733);
xor UO_173 (O_173,N_20918,N_20061);
nand UO_174 (O_174,N_22004,N_21024);
nor UO_175 (O_175,N_24791,N_22210);
nand UO_176 (O_176,N_23100,N_23391);
nand UO_177 (O_177,N_23389,N_20357);
or UO_178 (O_178,N_24759,N_20678);
nand UO_179 (O_179,N_21370,N_23959);
nand UO_180 (O_180,N_22882,N_24798);
nor UO_181 (O_181,N_22328,N_22176);
and UO_182 (O_182,N_24321,N_24257);
or UO_183 (O_183,N_22356,N_22422);
or UO_184 (O_184,N_20202,N_20322);
nand UO_185 (O_185,N_23861,N_20631);
nor UO_186 (O_186,N_21589,N_21507);
or UO_187 (O_187,N_21742,N_22123);
and UO_188 (O_188,N_22265,N_22445);
nor UO_189 (O_189,N_20066,N_21335);
or UO_190 (O_190,N_21163,N_20255);
nand UO_191 (O_191,N_23333,N_21870);
nor UO_192 (O_192,N_22002,N_22976);
nand UO_193 (O_193,N_22285,N_20624);
nor UO_194 (O_194,N_21943,N_20458);
nor UO_195 (O_195,N_23166,N_20047);
xor UO_196 (O_196,N_23254,N_22894);
nor UO_197 (O_197,N_24605,N_24743);
xnor UO_198 (O_198,N_22207,N_21477);
or UO_199 (O_199,N_23899,N_20746);
or UO_200 (O_200,N_24917,N_21320);
or UO_201 (O_201,N_22660,N_21289);
nand UO_202 (O_202,N_22182,N_20403);
or UO_203 (O_203,N_23315,N_22499);
nand UO_204 (O_204,N_20598,N_24577);
xnor UO_205 (O_205,N_21503,N_22262);
nor UO_206 (O_206,N_21233,N_20502);
or UO_207 (O_207,N_22069,N_20007);
nand UO_208 (O_208,N_20759,N_20883);
and UO_209 (O_209,N_20398,N_24272);
nand UO_210 (O_210,N_23509,N_23483);
and UO_211 (O_211,N_24005,N_24715);
nand UO_212 (O_212,N_24325,N_21805);
nor UO_213 (O_213,N_24139,N_23431);
and UO_214 (O_214,N_24817,N_20549);
nor UO_215 (O_215,N_23423,N_20629);
nand UO_216 (O_216,N_20208,N_22869);
nor UO_217 (O_217,N_24945,N_23527);
nor UO_218 (O_218,N_20849,N_20756);
nor UO_219 (O_219,N_20514,N_24993);
or UO_220 (O_220,N_21759,N_22966);
and UO_221 (O_221,N_23260,N_20527);
or UO_222 (O_222,N_22580,N_21142);
nand UO_223 (O_223,N_21881,N_20944);
nor UO_224 (O_224,N_24616,N_21758);
and UO_225 (O_225,N_22291,N_24753);
and UO_226 (O_226,N_21402,N_20036);
nand UO_227 (O_227,N_23970,N_21243);
and UO_228 (O_228,N_23628,N_22315);
nand UO_229 (O_229,N_24806,N_22106);
nand UO_230 (O_230,N_23162,N_22376);
xor UO_231 (O_231,N_20777,N_21170);
and UO_232 (O_232,N_20547,N_23051);
or UO_233 (O_233,N_23939,N_24347);
nor UO_234 (O_234,N_21960,N_23502);
or UO_235 (O_235,N_21164,N_24304);
or UO_236 (O_236,N_20838,N_23556);
nor UO_237 (O_237,N_23497,N_22470);
nor UO_238 (O_238,N_23651,N_23420);
nand UO_239 (O_239,N_24293,N_22642);
or UO_240 (O_240,N_22927,N_22740);
nand UO_241 (O_241,N_24736,N_22561);
xor UO_242 (O_242,N_23919,N_20966);
or UO_243 (O_243,N_21744,N_21796);
and UO_244 (O_244,N_23036,N_23842);
nand UO_245 (O_245,N_20455,N_22855);
nor UO_246 (O_246,N_24650,N_22902);
nand UO_247 (O_247,N_22980,N_21381);
and UO_248 (O_248,N_21134,N_20766);
xnor UO_249 (O_249,N_22431,N_20737);
nand UO_250 (O_250,N_24825,N_24706);
nor UO_251 (O_251,N_23448,N_22903);
nand UO_252 (O_252,N_23111,N_20981);
nand UO_253 (O_253,N_21284,N_23143);
and UO_254 (O_254,N_23382,N_20866);
and UO_255 (O_255,N_24302,N_23928);
and UO_256 (O_256,N_22989,N_21256);
nor UO_257 (O_257,N_24684,N_24639);
and UO_258 (O_258,N_20665,N_22816);
and UO_259 (O_259,N_23125,N_24277);
nand UO_260 (O_260,N_22148,N_22730);
nand UO_261 (O_261,N_22397,N_20194);
or UO_262 (O_262,N_20155,N_20166);
or UO_263 (O_263,N_20444,N_24493);
nor UO_264 (O_264,N_22586,N_24442);
nor UO_265 (O_265,N_22619,N_22039);
or UO_266 (O_266,N_20248,N_20647);
and UO_267 (O_267,N_24108,N_23476);
and UO_268 (O_268,N_23574,N_21664);
xor UO_269 (O_269,N_20272,N_23742);
nand UO_270 (O_270,N_21333,N_22588);
nand UO_271 (O_271,N_21019,N_20262);
nand UO_272 (O_272,N_21997,N_20752);
and UO_273 (O_273,N_22043,N_20411);
and UO_274 (O_274,N_22336,N_23719);
or UO_275 (O_275,N_21389,N_22697);
xnor UO_276 (O_276,N_22793,N_22143);
and UO_277 (O_277,N_22147,N_24165);
and UO_278 (O_278,N_23799,N_24539);
and UO_279 (O_279,N_21445,N_23417);
or UO_280 (O_280,N_22924,N_20001);
nand UO_281 (O_281,N_23279,N_24007);
xor UO_282 (O_282,N_24259,N_24086);
or UO_283 (O_283,N_20460,N_24412);
xor UO_284 (O_284,N_21220,N_21595);
nor UO_285 (O_285,N_23282,N_22724);
nand UO_286 (O_286,N_20909,N_20817);
or UO_287 (O_287,N_21426,N_21566);
nand UO_288 (O_288,N_22786,N_24595);
or UO_289 (O_289,N_20901,N_23482);
nand UO_290 (O_290,N_24455,N_20121);
or UO_291 (O_291,N_24482,N_20006);
nor UO_292 (O_292,N_21369,N_22216);
nor UO_293 (O_293,N_23754,N_20913);
nor UO_294 (O_294,N_23284,N_24184);
or UO_295 (O_295,N_24351,N_20658);
nor UO_296 (O_296,N_23986,N_23446);
and UO_297 (O_297,N_20104,N_23752);
and UO_298 (O_298,N_24570,N_21978);
and UO_299 (O_299,N_24246,N_24670);
nor UO_300 (O_300,N_22943,N_24730);
nand UO_301 (O_301,N_23761,N_24151);
nand UO_302 (O_302,N_20311,N_21701);
nand UO_303 (O_303,N_22688,N_24904);
nand UO_304 (O_304,N_24331,N_21141);
nor UO_305 (O_305,N_20427,N_24105);
nor UO_306 (O_306,N_23188,N_20153);
nor UO_307 (O_307,N_23864,N_21539);
or UO_308 (O_308,N_24688,N_20701);
nand UO_309 (O_309,N_21153,N_24471);
nor UO_310 (O_310,N_21026,N_20791);
nand UO_311 (O_311,N_23510,N_24354);
and UO_312 (O_312,N_22025,N_23388);
or UO_313 (O_313,N_21860,N_23034);
nand UO_314 (O_314,N_21244,N_24974);
xnor UO_315 (O_315,N_23244,N_21969);
nor UO_316 (O_316,N_20291,N_20636);
or UO_317 (O_317,N_23711,N_24631);
and UO_318 (O_318,N_21521,N_20592);
nand UO_319 (O_319,N_23686,N_23828);
nand UO_320 (O_320,N_22598,N_23149);
or UO_321 (O_321,N_23784,N_23749);
or UO_322 (O_322,N_22154,N_20052);
xnor UO_323 (O_323,N_22965,N_21938);
nor UO_324 (O_324,N_20523,N_22317);
and UO_325 (O_325,N_21957,N_24428);
nor UO_326 (O_326,N_22959,N_24297);
nor UO_327 (O_327,N_20289,N_24461);
nand UO_328 (O_328,N_23035,N_20096);
nor UO_329 (O_329,N_20508,N_24275);
and UO_330 (O_330,N_21570,N_20273);
and UO_331 (O_331,N_20880,N_24374);
or UO_332 (O_332,N_22406,N_21488);
xnor UO_333 (O_333,N_24683,N_21580);
or UO_334 (O_334,N_24283,N_24035);
or UO_335 (O_335,N_22111,N_22405);
nand UO_336 (O_336,N_22142,N_20378);
nor UO_337 (O_337,N_22000,N_23541);
and UO_338 (O_338,N_24816,N_24144);
or UO_339 (O_339,N_24934,N_21993);
and UO_340 (O_340,N_21989,N_24098);
or UO_341 (O_341,N_22878,N_23672);
or UO_342 (O_342,N_21632,N_21785);
nand UO_343 (O_343,N_20591,N_21065);
and UO_344 (O_344,N_24635,N_23121);
or UO_345 (O_345,N_23130,N_22948);
nor UO_346 (O_346,N_20729,N_23381);
nor UO_347 (O_347,N_21048,N_21800);
nand UO_348 (O_348,N_20927,N_23695);
and UO_349 (O_349,N_21752,N_24240);
or UO_350 (O_350,N_24726,N_22362);
nor UO_351 (O_351,N_20167,N_24454);
nor UO_352 (O_352,N_24402,N_24192);
nor UO_353 (O_353,N_23803,N_21657);
or UO_354 (O_354,N_23025,N_24962);
xnor UO_355 (O_355,N_22389,N_23024);
and UO_356 (O_356,N_21191,N_20290);
or UO_357 (O_357,N_23699,N_20580);
xnor UO_358 (O_358,N_20991,N_23538);
nor UO_359 (O_359,N_24608,N_21867);
or UO_360 (O_360,N_20197,N_21360);
or UO_361 (O_361,N_24458,N_20264);
nor UO_362 (O_362,N_20503,N_21847);
nand UO_363 (O_363,N_20780,N_20496);
and UO_364 (O_364,N_21706,N_23898);
or UO_365 (O_365,N_23935,N_22468);
nand UO_366 (O_366,N_24350,N_21693);
nand UO_367 (O_367,N_24219,N_20606);
nor UO_368 (O_368,N_22335,N_22115);
nor UO_369 (O_369,N_22354,N_24317);
nand UO_370 (O_370,N_20727,N_20259);
nand UO_371 (O_371,N_23146,N_21152);
xor UO_372 (O_372,N_20220,N_20163);
and UO_373 (O_373,N_24968,N_21767);
or UO_374 (O_374,N_21303,N_23798);
or UO_375 (O_375,N_21768,N_21691);
nand UO_376 (O_376,N_24563,N_23633);
or UO_377 (O_377,N_21481,N_21738);
xor UO_378 (O_378,N_20526,N_24248);
nand UO_379 (O_379,N_20009,N_22021);
or UO_380 (O_380,N_22525,N_24319);
and UO_381 (O_381,N_20938,N_22624);
and UO_382 (O_382,N_21305,N_24394);
xnor UO_383 (O_383,N_24967,N_23689);
and UO_384 (O_384,N_24055,N_22255);
or UO_385 (O_385,N_20802,N_23664);
nand UO_386 (O_386,N_21955,N_20409);
or UO_387 (O_387,N_23048,N_21246);
nand UO_388 (O_388,N_20789,N_21911);
nor UO_389 (O_389,N_24511,N_22059);
and UO_390 (O_390,N_24393,N_22970);
or UO_391 (O_391,N_22202,N_24886);
or UO_392 (O_392,N_23840,N_22530);
or UO_393 (O_393,N_23988,N_22679);
nor UO_394 (O_394,N_20949,N_23818);
nor UO_395 (O_395,N_22416,N_20360);
nand UO_396 (O_396,N_24781,N_21856);
nor UO_397 (O_397,N_23152,N_20413);
or UO_398 (O_398,N_24498,N_23723);
xnor UO_399 (O_399,N_21995,N_20213);
nand UO_400 (O_400,N_21930,N_22677);
nor UO_401 (O_401,N_21236,N_22352);
and UO_402 (O_402,N_24621,N_23119);
and UO_403 (O_403,N_20931,N_20739);
nand UO_404 (O_404,N_24562,N_24775);
xnor UO_405 (O_405,N_24709,N_21797);
nor UO_406 (O_406,N_24208,N_22957);
nand UO_407 (O_407,N_23114,N_20915);
or UO_408 (O_408,N_23182,N_21672);
nand UO_409 (O_409,N_24205,N_20390);
nand UO_410 (O_410,N_24083,N_21239);
and UO_411 (O_411,N_22434,N_20204);
and UO_412 (O_412,N_24090,N_22556);
nor UO_413 (O_413,N_21296,N_22961);
or UO_414 (O_414,N_22448,N_24912);
and UO_415 (O_415,N_24729,N_24871);
xnor UO_416 (O_416,N_20522,N_24164);
or UO_417 (O_417,N_23501,N_22528);
and UO_418 (O_418,N_24704,N_20280);
and UO_419 (O_419,N_24873,N_23673);
nand UO_420 (O_420,N_24045,N_24113);
nor UO_421 (O_421,N_24660,N_20027);
or UO_422 (O_422,N_24996,N_23097);
nor UO_423 (O_423,N_21215,N_21437);
nand UO_424 (O_424,N_21666,N_24969);
or UO_425 (O_425,N_21394,N_22735);
or UO_426 (O_426,N_23147,N_20900);
and UO_427 (O_427,N_21697,N_20330);
nor UO_428 (O_428,N_21414,N_22355);
or UO_429 (O_429,N_22673,N_23701);
or UO_430 (O_430,N_21452,N_22179);
nor UO_431 (O_431,N_23908,N_21105);
nor UO_432 (O_432,N_22519,N_22790);
nor UO_433 (O_433,N_20882,N_20464);
and UO_434 (O_434,N_24868,N_20353);
nand UO_435 (O_435,N_22627,N_24728);
and UO_436 (O_436,N_22908,N_22791);
xor UO_437 (O_437,N_23013,N_21252);
nand UO_438 (O_438,N_24981,N_20192);
nor UO_439 (O_439,N_24569,N_23942);
nor UO_440 (O_440,N_23876,N_21934);
or UO_441 (O_441,N_23605,N_21415);
xor UO_442 (O_442,N_23191,N_22767);
or UO_443 (O_443,N_20105,N_23615);
xor UO_444 (O_444,N_24664,N_20968);
xnor UO_445 (O_445,N_23210,N_24702);
or UO_446 (O_446,N_24559,N_24014);
nor UO_447 (O_447,N_24274,N_24042);
nor UO_448 (O_448,N_22892,N_23401);
nor UO_449 (O_449,N_24473,N_23211);
nor UO_450 (O_450,N_21051,N_20160);
and UO_451 (O_451,N_20755,N_22709);
or UO_452 (O_452,N_24476,N_21260);
and UO_453 (O_453,N_24346,N_24575);
or UO_454 (O_454,N_24462,N_23580);
nand UO_455 (O_455,N_20559,N_22401);
nand UO_456 (O_456,N_20315,N_23762);
and UO_457 (O_457,N_20187,N_21864);
and UO_458 (O_458,N_24528,N_22898);
or UO_459 (O_459,N_20488,N_22135);
nand UO_460 (O_460,N_21084,N_22806);
xor UO_461 (O_461,N_20386,N_20144);
nand UO_462 (O_462,N_24613,N_20217);
or UO_463 (O_463,N_21221,N_23429);
nor UO_464 (O_464,N_21444,N_24203);
nand UO_465 (O_465,N_24549,N_20969);
nand UO_466 (O_466,N_20453,N_24859);
and UO_467 (O_467,N_21731,N_22275);
nand UO_468 (O_468,N_22051,N_21395);
or UO_469 (O_469,N_22190,N_23577);
nor UO_470 (O_470,N_23241,N_20422);
and UO_471 (O_471,N_22593,N_24667);
nand UO_472 (O_472,N_20491,N_24823);
nand UO_473 (O_473,N_20183,N_23558);
nor UO_474 (O_474,N_23975,N_22321);
nor UO_475 (O_475,N_24285,N_24383);
nor UO_476 (O_476,N_22615,N_23657);
xor UO_477 (O_477,N_24525,N_24800);
and UO_478 (O_478,N_20122,N_24937);
nor UO_479 (O_479,N_21371,N_22747);
xor UO_480 (O_480,N_23503,N_22094);
nor UO_481 (O_481,N_20724,N_22144);
or UO_482 (O_482,N_21597,N_21099);
nor UO_483 (O_483,N_21525,N_23564);
or UO_484 (O_484,N_21311,N_20868);
or UO_485 (O_485,N_24724,N_20268);
and UO_486 (O_486,N_24345,N_23737);
nor UO_487 (O_487,N_21016,N_22364);
nand UO_488 (O_488,N_22849,N_20879);
and UO_489 (O_489,N_23873,N_22780);
xor UO_490 (O_490,N_21603,N_24423);
or UO_491 (O_491,N_23693,N_20649);
or UO_492 (O_492,N_20807,N_23453);
and UO_493 (O_493,N_20596,N_21678);
or UO_494 (O_494,N_22243,N_24384);
xnor UO_495 (O_495,N_24838,N_21774);
or UO_496 (O_496,N_23618,N_24076);
or UO_497 (O_497,N_21910,N_24314);
xnor UO_498 (O_498,N_22875,N_20490);
nand UO_499 (O_499,N_20214,N_23567);
nand UO_500 (O_500,N_23791,N_23594);
nor UO_501 (O_501,N_21276,N_22140);
nor UO_502 (O_502,N_21263,N_23694);
and UO_503 (O_503,N_20484,N_22759);
xnor UO_504 (O_504,N_23212,N_22515);
nor UO_505 (O_505,N_21471,N_24853);
nand UO_506 (O_506,N_21729,N_20054);
and UO_507 (O_507,N_20970,N_23459);
nand UO_508 (O_508,N_21651,N_22783);
xnor UO_509 (O_509,N_21902,N_20858);
and UO_510 (O_510,N_20301,N_23678);
nor UO_511 (O_511,N_22896,N_20787);
and UO_512 (O_512,N_23816,N_24872);
nor UO_513 (O_513,N_21698,N_22563);
xnor UO_514 (O_514,N_23057,N_21347);
nor UO_515 (O_515,N_22023,N_24986);
or UO_516 (O_516,N_22095,N_24755);
or UO_517 (O_517,N_24990,N_20611);
nand UO_518 (O_518,N_20196,N_23219);
or UO_519 (O_519,N_21831,N_21108);
nor UO_520 (O_520,N_20728,N_23320);
nand UO_521 (O_521,N_22294,N_24961);
nand UO_522 (O_522,N_22136,N_21174);
nand UO_523 (O_523,N_24935,N_23397);
nand UO_524 (O_524,N_22203,N_20903);
and UO_525 (O_525,N_20859,N_20768);
or UO_526 (O_526,N_24637,N_24863);
and UO_527 (O_527,N_20243,N_20207);
nor UO_528 (O_528,N_21919,N_20619);
nor UO_529 (O_529,N_21571,N_22256);
or UO_530 (O_530,N_21017,N_24289);
or UO_531 (O_531,N_23115,N_22651);
nor UO_532 (O_532,N_22904,N_22917);
or UO_533 (O_533,N_21114,N_23649);
and UO_534 (O_534,N_24456,N_22944);
nor UO_535 (O_535,N_21704,N_20034);
and UO_536 (O_536,N_24403,N_22891);
nand UO_537 (O_537,N_23078,N_21549);
or UO_538 (O_538,N_20767,N_20260);
nand UO_539 (O_539,N_22539,N_22988);
nand UO_540 (O_540,N_20095,N_24379);
nor UO_541 (O_541,N_24116,N_21915);
nand UO_542 (O_542,N_24880,N_24837);
xor UO_543 (O_543,N_24382,N_23478);
and UO_544 (O_544,N_20664,N_20795);
nand UO_545 (O_545,N_21713,N_24025);
or UO_546 (O_546,N_23213,N_24673);
nand UO_547 (O_547,N_20430,N_20010);
nor UO_548 (O_548,N_20428,N_23867);
and UO_549 (O_549,N_23245,N_23966);
nor UO_550 (O_550,N_23206,N_23859);
or UO_551 (O_551,N_22374,N_22674);
or UO_552 (O_552,N_21846,N_23266);
or UO_553 (O_553,N_24721,N_24410);
nand UO_554 (O_554,N_21548,N_24888);
nand UO_555 (O_555,N_21121,N_20494);
and UO_556 (O_556,N_23780,N_21058);
nor UO_557 (O_557,N_22761,N_20689);
nor UO_558 (O_558,N_24270,N_21607);
or UO_559 (O_559,N_23725,N_22196);
or UO_560 (O_560,N_22611,N_24239);
nor UO_561 (O_561,N_21629,N_21806);
or UO_562 (O_562,N_20278,N_23275);
or UO_563 (O_563,N_24640,N_23735);
nand UO_564 (O_564,N_22269,N_22045);
or UO_565 (O_565,N_24278,N_22809);
or UO_566 (O_566,N_23553,N_21352);
and UO_567 (O_567,N_20011,N_20557);
nand UO_568 (O_568,N_24636,N_21198);
nor UO_569 (O_569,N_23461,N_23611);
and UO_570 (O_570,N_22493,N_22446);
and UO_571 (O_571,N_21979,N_24841);
and UO_572 (O_572,N_24681,N_22146);
nor UO_573 (O_573,N_21653,N_23235);
xnor UO_574 (O_574,N_20026,N_20495);
nor UO_575 (O_575,N_20351,N_22232);
or UO_576 (O_576,N_20854,N_20673);
nand UO_577 (O_577,N_23468,N_23739);
nor UO_578 (O_578,N_24507,N_23305);
nand UO_579 (O_579,N_20227,N_22327);
nand UO_580 (O_580,N_22326,N_21486);
and UO_581 (O_581,N_24612,N_20967);
and UO_582 (O_582,N_20024,N_23764);
or UO_583 (O_583,N_21753,N_21686);
and UO_584 (O_584,N_24944,N_23247);
or UO_585 (O_585,N_21830,N_24842);
nor UO_586 (O_586,N_21781,N_22329);
and UO_587 (O_587,N_21986,N_23248);
and UO_588 (O_588,N_22905,N_20738);
and UO_589 (O_589,N_22931,N_24810);
xnor UO_590 (O_590,N_21081,N_21952);
and UO_591 (O_591,N_21971,N_24867);
nand UO_592 (O_592,N_23486,N_23838);
and UO_593 (O_593,N_24819,N_21309);
nor UO_594 (O_594,N_20801,N_22367);
nor UO_595 (O_595,N_21526,N_21435);
and UO_596 (O_596,N_24503,N_20887);
and UO_597 (O_597,N_24956,N_22837);
or UO_598 (O_598,N_24532,N_22813);
nand UO_599 (O_599,N_21694,N_23142);
and UO_600 (O_600,N_21009,N_22645);
and UO_601 (O_601,N_20424,N_22287);
or UO_602 (O_602,N_23976,N_24429);
and UO_603 (O_603,N_22524,N_21612);
or UO_604 (O_604,N_21783,N_24558);
nor UO_605 (O_605,N_24474,N_23498);
or UO_606 (O_606,N_21208,N_20644);
or UO_607 (O_607,N_23774,N_22286);
xnor UO_608 (O_608,N_21066,N_24071);
nor UO_609 (O_609,N_23234,N_24509);
nand UO_610 (O_610,N_21313,N_24797);
or UO_611 (O_611,N_24112,N_21857);
or UO_612 (O_612,N_24893,N_22879);
nor UO_613 (O_613,N_21118,N_23099);
nor UO_614 (O_614,N_22159,N_24573);
and UO_615 (O_615,N_24305,N_21308);
nor UO_616 (O_616,N_21882,N_23879);
nand UO_617 (O_617,N_23931,N_23327);
nor UO_618 (O_618,N_24407,N_22284);
nor UO_619 (O_619,N_23085,N_21880);
nor UO_620 (O_620,N_23730,N_20661);
nand UO_621 (O_621,N_22534,N_23654);
or UO_622 (O_622,N_24195,N_24228);
nand UO_623 (O_623,N_24763,N_23802);
or UO_624 (O_624,N_24367,N_23352);
or UO_625 (O_625,N_21297,N_23270);
or UO_626 (O_626,N_23038,N_24142);
and UO_627 (O_627,N_23255,N_24154);
or UO_628 (O_628,N_21730,N_20302);
nand UO_629 (O_629,N_20873,N_22247);
and UO_630 (O_630,N_20630,N_22387);
nor UO_631 (O_631,N_22782,N_20154);
or UO_632 (O_632,N_22559,N_24634);
or UO_633 (O_633,N_24168,N_22800);
xnor UO_634 (O_634,N_22827,N_24201);
nand UO_635 (O_635,N_23481,N_21670);
or UO_636 (O_636,N_23083,N_23112);
nand UO_637 (O_637,N_22017,N_24542);
and UO_638 (O_638,N_21074,N_20029);
and UO_639 (O_639,N_20608,N_20088);
or UO_640 (O_640,N_20436,N_24276);
nor UO_641 (O_641,N_20185,N_24421);
nand UO_642 (O_642,N_21457,N_22574);
nand UO_643 (O_643,N_21673,N_20305);
nor UO_644 (O_644,N_24774,N_21104);
nand UO_645 (O_645,N_20479,N_24963);
and UO_646 (O_646,N_22472,N_22035);
and UO_647 (O_647,N_20676,N_24587);
and UO_648 (O_648,N_24218,N_24229);
nor UO_649 (O_649,N_24010,N_20660);
or UO_650 (O_650,N_22488,N_21078);
or UO_651 (O_651,N_22010,N_23168);
or UO_652 (O_652,N_23396,N_24388);
nor UO_653 (O_653,N_23334,N_21585);
nor UO_654 (O_654,N_22040,N_23196);
and UO_655 (O_655,N_21238,N_20441);
or UO_656 (O_656,N_22754,N_23834);
nor UO_657 (O_657,N_20835,N_23341);
and UO_658 (O_658,N_20687,N_23529);
nand UO_659 (O_659,N_23470,N_24727);
and UO_660 (O_660,N_20111,N_23887);
nand UO_661 (O_661,N_23108,N_23795);
xor UO_662 (O_662,N_22330,N_22541);
and UO_663 (O_663,N_22403,N_24475);
and UO_664 (O_664,N_21722,N_20282);
and UO_665 (O_665,N_20806,N_24227);
and UO_666 (O_666,N_23267,N_24149);
and UO_667 (O_667,N_21364,N_23561);
and UO_668 (O_668,N_24049,N_21561);
or UO_669 (O_669,N_20415,N_24692);
nor UO_670 (O_670,N_21937,N_24096);
or UO_671 (O_671,N_24409,N_23309);
nand UO_672 (O_672,N_20733,N_22233);
and UO_673 (O_673,N_24574,N_22655);
nor UO_674 (O_674,N_20861,N_20131);
nand UO_675 (O_675,N_23916,N_24158);
xor UO_676 (O_676,N_23871,N_24459);
and UO_677 (O_677,N_24085,N_24047);
and UO_678 (O_678,N_23949,N_23042);
or UO_679 (O_679,N_20705,N_24984);
nor UO_680 (O_680,N_22695,N_23437);
and UO_681 (O_681,N_20057,N_23398);
or UO_682 (O_682,N_24852,N_24648);
nand UO_683 (O_683,N_21699,N_20819);
nor UO_684 (O_684,N_22504,N_22606);
or UO_685 (O_685,N_21973,N_20750);
or UO_686 (O_686,N_22369,N_21712);
nand UO_687 (O_687,N_21652,N_20829);
and UO_688 (O_688,N_21696,N_24597);
and UO_689 (O_689,N_23753,N_23687);
or UO_690 (O_690,N_24745,N_20847);
xnor UO_691 (O_691,N_23290,N_20857);
nor UO_692 (O_692,N_24839,N_23151);
and UO_693 (O_693,N_20293,N_21267);
nor UO_694 (O_694,N_24803,N_20265);
and UO_695 (O_695,N_22371,N_20341);
nand UO_696 (O_696,N_22368,N_20811);
nor UO_697 (O_697,N_22459,N_24739);
xnor UO_698 (O_698,N_24959,N_24622);
or UO_699 (O_699,N_24754,N_22492);
and UO_700 (O_700,N_21057,N_24002);
nand UO_701 (O_701,N_24628,N_23365);
nor UO_702 (O_702,N_23892,N_21079);
nor UO_703 (O_703,N_21648,N_22543);
nand UO_704 (O_704,N_24487,N_22231);
xnor UO_705 (O_705,N_24882,N_23534);
or UO_706 (O_706,N_20723,N_22312);
nand UO_707 (O_707,N_21137,N_20907);
or UO_708 (O_708,N_21491,N_21624);
and UO_709 (O_709,N_24422,N_24242);
and UO_710 (O_710,N_24765,N_22572);
and UO_711 (O_711,N_20986,N_23009);
xor UO_712 (O_712,N_23030,N_21947);
nand UO_713 (O_713,N_22339,N_23636);
or UO_714 (O_714,N_23089,N_22098);
or UO_715 (O_715,N_23858,N_20579);
nor UO_716 (O_716,N_22267,N_22803);
and UO_717 (O_717,N_24898,N_24520);
nand UO_718 (O_718,N_22388,N_24290);
and UO_719 (O_719,N_20309,N_23311);
and UO_720 (O_720,N_24500,N_23187);
nand UO_721 (O_721,N_24510,N_21475);
nand UO_722 (O_722,N_22373,N_21618);
or UO_723 (O_723,N_22994,N_22462);
or UO_724 (O_724,N_22863,N_22814);
nand UO_725 (O_725,N_20172,N_23463);
and UO_726 (O_726,N_21567,N_23200);
or UO_727 (O_727,N_21338,N_23722);
nand UO_728 (O_728,N_23109,N_22293);
nand UO_729 (O_729,N_24341,N_22604);
nand UO_730 (O_730,N_21615,N_22460);
nor UO_731 (O_731,N_21418,N_24465);
nand UO_732 (O_732,N_20389,N_23945);
nor UO_733 (O_733,N_23854,N_21895);
nor UO_734 (O_734,N_22386,N_22011);
nand UO_735 (O_735,N_20978,N_23878);
and UO_736 (O_736,N_23622,N_24832);
nor UO_737 (O_737,N_22996,N_24666);
or UO_738 (O_738,N_22019,N_22242);
nor UO_739 (O_739,N_23727,N_21194);
or UO_740 (O_740,N_21111,N_24720);
nor UO_741 (O_741,N_20356,N_21351);
xnor UO_742 (O_742,N_24182,N_23821);
and UO_743 (O_743,N_20158,N_24338);
or UO_744 (O_744,N_20108,N_21703);
or UO_745 (O_745,N_22731,N_22852);
xor UO_746 (O_746,N_22254,N_23479);
xor UO_747 (O_747,N_21301,N_22888);
or UO_748 (O_748,N_23371,N_23787);
nor UO_749 (O_749,N_23563,N_23836);
and UO_750 (O_750,N_21813,N_23457);
nor UO_751 (O_751,N_23769,N_23186);
nand UO_752 (O_752,N_24469,N_21131);
and UO_753 (O_753,N_24526,N_23644);
xor UO_754 (O_754,N_22400,N_24938);
nand UO_755 (O_755,N_21985,N_24625);
or UO_756 (O_756,N_22828,N_24019);
or UO_757 (O_757,N_21255,N_22833);
nand UO_758 (O_758,N_21820,N_24329);
or UO_759 (O_759,N_20955,N_24611);
nand UO_760 (O_760,N_23944,N_22271);
or UO_761 (O_761,N_21438,N_21006);
or UO_762 (O_762,N_23906,N_24978);
or UO_763 (O_763,N_21404,N_21413);
or UO_764 (O_764,N_21791,N_21754);
nor UO_765 (O_765,N_20440,N_22811);
nand UO_766 (O_766,N_21950,N_24675);
or UO_767 (O_767,N_21166,N_23075);
nand UO_768 (O_768,N_22920,N_21966);
nand UO_769 (O_769,N_22234,N_20872);
and UO_770 (O_770,N_23124,N_22438);
and UO_771 (O_771,N_22338,N_22359);
nor UO_772 (O_772,N_21872,N_21497);
or UO_773 (O_773,N_22195,N_20270);
and UO_774 (O_774,N_21028,N_22425);
or UO_775 (O_775,N_24626,N_22197);
and UO_776 (O_776,N_22748,N_23455);
and UO_777 (O_777,N_24828,N_20930);
nor UO_778 (O_778,N_22415,N_20878);
nand UO_779 (O_779,N_24323,N_24776);
and UO_780 (O_780,N_22710,N_21746);
and UO_781 (O_781,N_23325,N_22990);
nor UO_782 (O_782,N_21821,N_20731);
nand UO_783 (O_783,N_21839,N_20947);
or UO_784 (O_784,N_23346,N_20335);
and UO_785 (O_785,N_22911,N_22016);
or UO_786 (O_786,N_21366,N_24856);
nor UO_787 (O_787,N_24226,N_22477);
nand UO_788 (O_788,N_21855,N_24807);
nor UO_789 (O_789,N_24711,N_21838);
or UO_790 (O_790,N_23379,N_23971);
and UO_791 (O_791,N_20877,N_20169);
nor UO_792 (O_792,N_23399,N_23885);
and UO_793 (O_793,N_22558,N_21705);
nor UO_794 (O_794,N_23488,N_21799);
nand UO_795 (O_795,N_20889,N_22520);
or UO_796 (O_796,N_23484,N_23023);
nand UO_797 (O_797,N_23883,N_22810);
xnor UO_798 (O_798,N_22169,N_24894);
nand UO_799 (O_799,N_23494,N_24805);
nor UO_800 (O_800,N_20776,N_23306);
and UO_801 (O_801,N_22334,N_22693);
nand UO_802 (O_802,N_24991,N_21959);
nand UO_803 (O_803,N_22139,N_23696);
xnor UO_804 (O_804,N_21522,N_24180);
nor UO_805 (O_805,N_22100,N_20236);
nor UO_806 (O_806,N_23833,N_23449);
and UO_807 (O_807,N_23104,N_23853);
and UO_808 (O_808,N_24915,N_23612);
or UO_809 (O_809,N_24514,N_24834);
xnor UO_810 (O_810,N_21528,N_24363);
nand UO_811 (O_811,N_22776,N_24714);
nand UO_812 (O_812,N_22351,N_23741);
or UO_813 (O_813,N_22797,N_20313);
or UO_814 (O_814,N_24026,N_24740);
nor UO_815 (O_815,N_20827,N_20077);
nor UO_816 (O_816,N_20133,N_23294);
nand UO_817 (O_817,N_24097,N_21453);
or UO_818 (O_818,N_24291,N_24078);
and UO_819 (O_819,N_24821,N_22845);
or UO_820 (O_820,N_24593,N_22897);
xnor UO_821 (O_821,N_22171,N_24854);
nand UO_822 (O_822,N_22983,N_23627);
nand UO_823 (O_823,N_22962,N_24404);
and UO_824 (O_824,N_23027,N_24645);
nor UO_825 (O_825,N_24418,N_21302);
and UO_826 (O_826,N_20355,N_22496);
nand UO_827 (O_827,N_20652,N_21061);
or UO_828 (O_828,N_24923,N_20125);
or UO_829 (O_829,N_20310,N_21489);
and UO_830 (O_830,N_24173,N_24413);
nand UO_831 (O_831,N_22975,N_20863);
nand UO_832 (O_832,N_22546,N_23081);
or UO_833 (O_833,N_23839,N_23050);
or UO_834 (O_834,N_23724,N_22370);
nor UO_835 (O_835,N_20764,N_23982);
or UO_836 (O_836,N_23710,N_23008);
and UO_837 (O_837,N_24375,N_23547);
xor UO_838 (O_838,N_20008,N_22510);
xor UO_839 (O_839,N_21204,N_20246);
nand UO_840 (O_840,N_23958,N_24903);
nor UO_841 (O_841,N_22760,N_23360);
nand UO_842 (O_842,N_24134,N_21588);
nor UO_843 (O_843,N_20613,N_22925);
nor UO_844 (O_844,N_21685,N_22830);
or UO_845 (O_845,N_21682,N_22322);
nor UO_846 (O_846,N_21644,N_21022);
nand UO_847 (O_847,N_24128,N_23268);
and UO_848 (O_848,N_20741,N_20147);
or UO_849 (O_849,N_21376,N_23807);
or UO_850 (O_850,N_23540,N_20140);
or UO_851 (O_851,N_20609,N_20324);
nor UO_852 (O_852,N_22922,N_20211);
nand UO_853 (O_853,N_20218,N_22853);
nor UO_854 (O_854,N_21981,N_23643);
xnor UO_855 (O_855,N_23454,N_23530);
xor UO_856 (O_856,N_21213,N_20816);
or UO_857 (O_857,N_24833,N_21182);
or UO_858 (O_858,N_24533,N_20784);
nor UO_859 (O_859,N_24435,N_23285);
nor UO_860 (O_860,N_21261,N_21951);
nand UO_861 (O_861,N_22175,N_21013);
and UO_862 (O_862,N_22940,N_20045);
nor UO_863 (O_863,N_21802,N_22456);
nand UO_864 (O_864,N_21112,N_23301);
and UO_865 (O_865,N_21034,N_23660);
nor UO_866 (O_866,N_23102,N_23000);
nor UO_867 (O_867,N_20932,N_20684);
and UO_868 (O_868,N_24063,N_22570);
xnor UO_869 (O_869,N_23205,N_23985);
or UO_870 (O_870,N_21633,N_20703);
nor UO_871 (O_871,N_21092,N_21963);
nor UO_872 (O_872,N_20392,N_22483);
xor UO_873 (O_873,N_22726,N_21344);
nand UO_874 (O_874,N_22160,N_23565);
nor UO_875 (O_875,N_20073,N_22129);
nor UO_876 (O_876,N_20833,N_22108);
and UO_877 (O_877,N_23616,N_21259);
or UO_878 (O_878,N_20963,N_20585);
nand UO_879 (O_879,N_22861,N_20896);
and UO_880 (O_880,N_20492,N_21766);
and UO_881 (O_881,N_20736,N_21734);
and UO_882 (O_882,N_21586,N_22705);
nand UO_883 (O_883,N_21596,N_21818);
nand UO_884 (O_884,N_22794,N_24516);
and UO_885 (O_885,N_24999,N_22603);
or UO_886 (O_886,N_21222,N_24178);
nand UO_887 (O_887,N_21844,N_20018);
nor UO_888 (O_888,N_20615,N_20760);
and UO_889 (O_889,N_20876,N_24310);
nand UO_890 (O_890,N_23348,N_24849);
nor UO_891 (O_891,N_24214,N_23177);
and UO_892 (O_892,N_20031,N_22887);
nor UO_893 (O_893,N_21324,N_22029);
and UO_894 (O_894,N_21583,N_24155);
or UO_895 (O_895,N_24719,N_21535);
or UO_896 (O_896,N_21726,N_20085);
or UO_897 (O_897,N_22178,N_21554);
nand UO_898 (O_898,N_24392,N_22872);
and UO_899 (O_899,N_24243,N_21337);
xnor UO_900 (O_900,N_20669,N_22522);
nand UO_901 (O_901,N_20292,N_24439);
xor UO_902 (O_902,N_24448,N_20704);
nand UO_903 (O_903,N_20254,N_23001);
xor UO_904 (O_904,N_23175,N_24145);
and UO_905 (O_905,N_24515,N_21196);
nor UO_906 (O_906,N_20929,N_20911);
nand UO_907 (O_907,N_22419,N_22474);
nand UO_908 (O_908,N_20438,N_20996);
nand UO_909 (O_909,N_21382,N_22873);
nand UO_910 (O_910,N_23227,N_24039);
and UO_911 (O_911,N_22476,N_20641);
and UO_912 (O_912,N_20642,N_22648);
and UO_913 (O_913,N_20770,N_22968);
and UO_914 (O_914,N_23467,N_22802);
nor UO_915 (O_915,N_23261,N_21193);
nand UO_916 (O_916,N_21572,N_23137);
and UO_917 (O_917,N_21887,N_21120);
nor UO_918 (O_918,N_22187,N_23808);
nand UO_919 (O_919,N_22343,N_22238);
nor UO_920 (O_920,N_21920,N_24468);
and UO_921 (O_921,N_20790,N_21605);
or UO_922 (O_922,N_23225,N_24126);
and UO_923 (O_923,N_21610,N_22644);
and UO_924 (O_924,N_22964,N_20992);
nor UO_925 (O_925,N_22820,N_21889);
or UO_926 (O_926,N_22554,N_21984);
xor UO_927 (O_927,N_23058,N_20040);
or UO_928 (O_928,N_22799,N_23974);
or UO_929 (O_929,N_23238,N_20605);
or UO_930 (O_930,N_22858,N_22041);
nor UO_931 (O_931,N_22581,N_21564);
nor UO_932 (O_932,N_21683,N_21098);
or UO_933 (O_933,N_24769,N_22635);
and UO_934 (O_934,N_22220,N_23135);
and UO_935 (O_935,N_21896,N_20718);
nand UO_936 (O_936,N_22676,N_22465);
or UO_937 (O_937,N_20928,N_23650);
or UO_938 (O_938,N_22114,N_22209);
xnor UO_939 (O_939,N_20692,N_23010);
or UO_940 (O_940,N_20134,N_20225);
nor UO_941 (O_941,N_23661,N_21144);
nor UO_942 (O_942,N_23150,N_21770);
or UO_943 (O_943,N_24717,N_23856);
nand UO_944 (O_944,N_21035,N_20917);
xnor UO_945 (O_945,N_20960,N_21067);
and UO_946 (O_946,N_21214,N_20145);
nor UO_947 (O_947,N_23318,N_20534);
and UO_948 (O_948,N_21743,N_21440);
nor UO_949 (O_949,N_24629,N_23702);
nand UO_950 (O_950,N_24555,N_24082);
nand UO_951 (O_951,N_20000,N_21717);
or UO_952 (O_952,N_21832,N_22360);
nand UO_953 (O_953,N_23631,N_23948);
and UO_954 (O_954,N_22999,N_24211);
xor UO_955 (O_955,N_24975,N_22174);
nand UO_956 (O_956,N_24236,N_24910);
xor UO_957 (O_957,N_23179,N_21145);
xnor UO_958 (O_958,N_20201,N_24777);
or UO_959 (O_959,N_23447,N_20112);
or UO_960 (O_960,N_21933,N_21628);
and UO_961 (O_961,N_24932,N_20212);
xnor UO_962 (O_962,N_21323,N_22185);
nor UO_963 (O_963,N_22347,N_20431);
xnor UO_964 (O_964,N_24366,N_21032);
or UO_965 (O_965,N_24538,N_22564);
nand UO_966 (O_966,N_24885,N_22054);
nand UO_967 (O_967,N_24988,N_21349);
and UO_968 (O_968,N_22473,N_21231);
or UO_969 (O_969,N_20097,N_22478);
nor UO_970 (O_970,N_20342,N_23296);
nand UO_971 (O_971,N_22241,N_20657);
or UO_972 (O_972,N_22640,N_23243);
nand UO_973 (O_973,N_24930,N_21298);
or UO_974 (O_974,N_22699,N_21416);
and UO_975 (O_975,N_22261,N_21970);
nand UO_976 (O_976,N_22151,N_23045);
nor UO_977 (O_977,N_22566,N_22844);
nand UO_978 (O_978,N_24440,N_21173);
or UO_979 (O_979,N_20058,N_20382);
nor UO_980 (O_980,N_23677,N_22508);
nand UO_981 (O_981,N_21747,N_20041);
and UO_982 (O_982,N_20602,N_23091);
and UO_983 (O_983,N_23185,N_23157);
nor UO_984 (O_984,N_24215,N_21518);
xor UO_985 (O_985,N_22717,N_22453);
nor UO_986 (O_986,N_20517,N_24883);
nor UO_987 (O_987,N_22597,N_23033);
and UO_988 (O_988,N_20072,N_22715);
and UO_989 (O_989,N_21257,N_21175);
or UO_990 (O_990,N_24490,N_22647);
and UO_991 (O_991,N_20449,N_23844);
nand UO_992 (O_992,N_23830,N_23837);
or UO_993 (O_993,N_20127,N_22649);
and UO_994 (O_994,N_21472,N_22237);
and UO_995 (O_995,N_22283,N_20053);
and UO_996 (O_996,N_20511,N_21278);
xor UO_997 (O_997,N_22153,N_20551);
or UO_998 (O_998,N_23973,N_23106);
nor UO_999 (O_999,N_21419,N_23782);
nor UO_1000 (O_1000,N_21944,N_21230);
or UO_1001 (O_1001,N_24265,N_22280);
or UO_1002 (O_1002,N_20266,N_22050);
xnor UO_1003 (O_1003,N_20751,N_20945);
nor UO_1004 (O_1004,N_22217,N_24387);
nor UO_1005 (O_1005,N_20697,N_24125);
or UO_1006 (O_1006,N_21110,N_22972);
nor UO_1007 (O_1007,N_23473,N_22633);
nand UO_1008 (O_1008,N_22058,N_24013);
nand UO_1009 (O_1009,N_22357,N_24568);
and UO_1010 (O_1010,N_21958,N_24583);
nand UO_1011 (O_1011,N_21190,N_21749);
nor UO_1012 (O_1012,N_24399,N_21926);
nand UO_1013 (O_1013,N_22282,N_24037);
xor UO_1014 (O_1014,N_22092,N_22414);
nand UO_1015 (O_1015,N_20499,N_20181);
xnor UO_1016 (O_1016,N_20685,N_21383);
xnor UO_1017 (O_1017,N_21458,N_20837);
nor UO_1018 (O_1018,N_22411,N_20510);
nor UO_1019 (O_1019,N_20019,N_24518);
nor UO_1020 (O_1020,N_22078,N_22880);
or UO_1021 (O_1021,N_23194,N_23843);
and UO_1022 (O_1022,N_23046,N_23760);
nor UO_1023 (O_1023,N_21334,N_23555);
and UO_1024 (O_1024,N_24649,N_22155);
or UO_1025 (O_1025,N_22253,N_22215);
and UO_1026 (O_1026,N_20078,N_22133);
xnor UO_1027 (O_1027,N_23575,N_24481);
nor UO_1028 (O_1028,N_21075,N_20792);
and UO_1029 (O_1029,N_20707,N_20425);
nand UO_1030 (O_1030,N_20175,N_24831);
nor UO_1031 (O_1031,N_24630,N_21822);
or UO_1032 (O_1032,N_23786,N_21053);
and UO_1033 (O_1033,N_21519,N_24554);
and UO_1034 (O_1034,N_23968,N_22122);
and UO_1035 (O_1035,N_20316,N_20483);
or UO_1036 (O_1036,N_22686,N_22170);
nor UO_1037 (O_1037,N_24093,N_20663);
xor UO_1038 (O_1038,N_20137,N_23117);
xnor UO_1039 (O_1039,N_20796,N_23775);
nor UO_1040 (O_1040,N_24674,N_23566);
nor UO_1041 (O_1041,N_22669,N_24391);
nor UO_1042 (O_1042,N_22479,N_20314);
and UO_1043 (O_1043,N_20060,N_23059);
and UO_1044 (O_1044,N_23291,N_23912);
and UO_1045 (O_1045,N_23474,N_22396);
or UO_1046 (O_1046,N_23685,N_21530);
or UO_1047 (O_1047,N_22744,N_22074);
or UO_1048 (O_1048,N_23913,N_24939);
nand UO_1049 (O_1049,N_22224,N_23317);
or UO_1050 (O_1050,N_21721,N_21751);
and UO_1051 (O_1051,N_22301,N_20401);
or UO_1052 (O_1052,N_22951,N_22992);
xor UO_1053 (O_1053,N_22012,N_24352);
or UO_1054 (O_1054,N_22189,N_20959);
or UO_1055 (O_1055,N_24654,N_23640);
xnor UO_1056 (O_1056,N_24166,N_20414);
nand UO_1057 (O_1057,N_22070,N_23197);
and UO_1058 (O_1058,N_23323,N_20300);
nand UO_1059 (O_1059,N_23920,N_21183);
nor UO_1060 (O_1060,N_20250,N_22173);
nor UO_1061 (O_1061,N_23571,N_24824);
nand UO_1062 (O_1062,N_20588,N_21180);
nand UO_1063 (O_1063,N_20821,N_24947);
nor UO_1064 (O_1064,N_24780,N_21598);
nand UO_1065 (O_1065,N_23286,N_22311);
and UO_1066 (O_1066,N_20312,N_23441);
nand UO_1067 (O_1067,N_21992,N_22770);
nor UO_1068 (O_1068,N_23364,N_23619);
xnor UO_1069 (O_1069,N_20445,N_21343);
nand UO_1070 (O_1070,N_24697,N_24746);
xor UO_1071 (O_1071,N_24813,N_24591);
and UO_1072 (O_1072,N_21942,N_24846);
or UO_1073 (O_1073,N_21562,N_23378);
or UO_1074 (O_1074,N_20237,N_23524);
nand UO_1075 (O_1075,N_22859,N_23570);
or UO_1076 (O_1076,N_21812,N_20933);
or UO_1077 (O_1077,N_22583,N_21842);
or UO_1078 (O_1078,N_24891,N_24433);
or UO_1079 (O_1079,N_23338,N_23133);
and UO_1080 (O_1080,N_20984,N_22569);
and UO_1081 (O_1081,N_20924,N_24353);
nand UO_1082 (O_1082,N_24207,N_20509);
nor UO_1083 (O_1083,N_22077,N_21125);
nor UO_1084 (O_1084,N_24609,N_20800);
nand UO_1085 (O_1085,N_23412,N_21592);
and UO_1086 (O_1086,N_23118,N_23890);
and UO_1087 (O_1087,N_22239,N_24668);
and UO_1088 (O_1088,N_24443,N_23292);
nor UO_1089 (O_1089,N_21327,N_21655);
or UO_1090 (O_1090,N_20690,N_21927);
and UO_1091 (O_1091,N_20867,N_24927);
nand UO_1092 (O_1092,N_20758,N_22720);
xor UO_1093 (O_1093,N_20805,N_23439);
xnor UO_1094 (O_1094,N_24878,N_22031);
xnor UO_1095 (O_1095,N_21412,N_20747);
and UO_1096 (O_1096,N_21976,N_22299);
or UO_1097 (O_1097,N_24460,N_22500);
nand UO_1098 (O_1098,N_20276,N_23923);
xnor UO_1099 (O_1099,N_23981,N_21148);
or UO_1100 (O_1100,N_23433,N_24677);
nand UO_1101 (O_1101,N_20786,N_24427);
nand UO_1102 (O_1102,N_20139,N_24875);
or UO_1103 (O_1103,N_24971,N_24492);
nand UO_1104 (O_1104,N_20554,N_21378);
nor UO_1105 (O_1105,N_22916,N_23770);
nor UO_1106 (O_1106,N_20645,N_21319);
and UO_1107 (O_1107,N_21559,N_24890);
or UO_1108 (O_1108,N_22412,N_20989);
nor UO_1109 (O_1109,N_20612,N_21372);
xnor UO_1110 (O_1110,N_20116,N_21576);
or UO_1111 (O_1111,N_24118,N_23630);
nor UO_1112 (O_1112,N_23123,N_22701);
nor UO_1113 (O_1113,N_24376,N_20107);
nand UO_1114 (O_1114,N_22668,N_22778);
nand UO_1115 (O_1115,N_24284,N_21033);
nand UO_1116 (O_1116,N_20565,N_24693);
nand UO_1117 (O_1117,N_20136,N_23617);
nor UO_1118 (O_1118,N_22973,N_20722);
or UO_1119 (O_1119,N_21465,N_20132);
nand UO_1120 (O_1120,N_20274,N_23545);
or UO_1121 (O_1121,N_22450,N_24919);
nand UO_1122 (O_1122,N_24866,N_21043);
or UO_1123 (O_1123,N_20574,N_21786);
and UO_1124 (O_1124,N_23426,N_20757);
nor UO_1125 (O_1125,N_22125,N_21103);
or UO_1126 (O_1126,N_23139,N_21201);
and UO_1127 (O_1127,N_23728,N_21573);
nand UO_1128 (O_1128,N_23597,N_21689);
and UO_1129 (O_1129,N_21408,N_23380);
and UO_1130 (O_1130,N_24712,N_23178);
nand UO_1131 (O_1131,N_22064,N_24048);
or UO_1132 (O_1132,N_20025,N_21188);
nor UO_1133 (O_1133,N_21626,N_21593);
and UO_1134 (O_1134,N_22969,N_24571);
nand UO_1135 (O_1135,N_22949,N_24908);
nand UO_1136 (O_1136,N_24051,N_21940);
nor UO_1137 (O_1137,N_24337,N_23037);
nor UO_1138 (O_1138,N_20575,N_24848);
or UO_1139 (O_1139,N_20091,N_20973);
and UO_1140 (O_1140,N_22099,N_20720);
nor UO_1141 (O_1141,N_23734,N_21837);
and UO_1142 (O_1142,N_24954,N_21547);
nand UO_1143 (O_1143,N_21714,N_21080);
or UO_1144 (O_1144,N_20568,N_21529);
or UO_1145 (O_1145,N_24031,N_21154);
and UO_1146 (O_1146,N_20337,N_20420);
nand UO_1147 (O_1147,N_22382,N_21322);
or UO_1148 (O_1148,N_21157,N_20012);
and UO_1149 (O_1149,N_24601,N_22798);
and UO_1150 (O_1150,N_24087,N_23265);
nand UO_1151 (O_1151,N_24332,N_23904);
or UO_1152 (O_1152,N_20126,N_22788);
nand UO_1153 (O_1153,N_22501,N_24306);
and UO_1154 (O_1154,N_23706,N_22841);
nand UO_1155 (O_1155,N_23409,N_21793);
and UO_1156 (O_1156,N_24004,N_23755);
xnor UO_1157 (O_1157,N_23165,N_24700);
and UO_1158 (O_1158,N_21373,N_23987);
nor UO_1159 (O_1159,N_23785,N_21312);
and UO_1160 (O_1160,N_22378,N_21353);
or UO_1161 (O_1161,N_21674,N_21527);
nor UO_1162 (O_1162,N_22222,N_23910);
nor UO_1163 (O_1163,N_23938,N_20595);
nor UO_1164 (O_1164,N_21285,N_20843);
nand UO_1165 (O_1165,N_21659,N_22380);
and UO_1166 (O_1166,N_24303,N_24106);
or UO_1167 (O_1167,N_20505,N_24160);
or UO_1168 (O_1168,N_20345,N_24814);
or UO_1169 (O_1169,N_20385,N_24202);
or UO_1170 (O_1170,N_23684,N_22480);
xnor UO_1171 (O_1171,N_24830,N_24193);
or UO_1172 (O_1172,N_23493,N_20646);
and UO_1173 (O_1173,N_22198,N_22081);
and UO_1174 (O_1174,N_22622,N_23535);
nand UO_1175 (O_1175,N_22281,N_22945);
or UO_1176 (O_1176,N_24072,N_20958);
or UO_1177 (O_1177,N_23195,N_23559);
xor UO_1178 (O_1178,N_22974,N_20216);
and UO_1179 (O_1179,N_21854,N_21874);
nor UO_1180 (O_1180,N_22670,N_21932);
or UO_1181 (O_1181,N_22292,N_21304);
or UO_1182 (O_1182,N_21676,N_24602);
or UO_1183 (O_1183,N_24527,N_22537);
nand UO_1184 (O_1184,N_20044,N_20251);
nor UO_1185 (O_1185,N_21249,N_24943);
and UO_1186 (O_1186,N_20391,N_20038);
nand UO_1187 (O_1187,N_21824,N_23811);
or UO_1188 (O_1188,N_21281,N_22096);
or UO_1189 (O_1189,N_20650,N_24936);
nand UO_1190 (O_1190,N_21671,N_23209);
nor UO_1191 (O_1191,N_21126,N_22038);
nor UO_1192 (O_1192,N_23442,N_21482);
and UO_1193 (O_1193,N_20812,N_20783);
nor UO_1194 (O_1194,N_21023,N_23744);
xnor UO_1195 (O_1195,N_24250,N_24931);
nor UO_1196 (O_1196,N_24540,N_24088);
xor UO_1197 (O_1197,N_22487,N_23820);
nand UO_1198 (O_1198,N_23679,N_22481);
or UO_1199 (O_1199,N_22204,N_20988);
or UO_1200 (O_1200,N_22840,N_21317);
and UO_1201 (O_1201,N_22864,N_21386);
nor UO_1202 (O_1202,N_23355,N_24438);
nor UO_1203 (O_1203,N_24135,N_21187);
nand UO_1204 (O_1204,N_24614,N_22551);
and UO_1205 (O_1205,N_21025,N_24676);
and UO_1206 (O_1206,N_21346,N_23688);
and UO_1207 (O_1207,N_23801,N_23300);
xor UO_1208 (O_1208,N_21167,N_21908);
and UO_1209 (O_1209,N_20506,N_20186);
nor UO_1210 (O_1210,N_21424,N_24523);
or UO_1211 (O_1211,N_21608,N_24175);
nor UO_1212 (O_1212,N_24197,N_21631);
and UO_1213 (O_1213,N_23040,N_24682);
nor UO_1214 (O_1214,N_23835,N_24804);
nor UO_1215 (O_1215,N_20515,N_22985);
and UO_1216 (O_1216,N_20119,N_23733);
or UO_1217 (O_1217,N_23593,N_22164);
or UO_1218 (O_1218,N_21341,N_24157);
nand UO_1219 (O_1219,N_24494,N_24922);
and UO_1220 (O_1220,N_22227,N_20864);
and UO_1221 (O_1221,N_20198,N_23810);
and UO_1222 (O_1222,N_24381,N_21946);
nand UO_1223 (O_1223,N_23080,N_20578);
xnor UO_1224 (O_1224,N_21619,N_20529);
nand UO_1225 (O_1225,N_21665,N_23438);
or UO_1226 (O_1226,N_24489,N_24389);
or UO_1227 (O_1227,N_21994,N_22270);
or UO_1228 (O_1228,N_21900,N_24124);
xor UO_1229 (O_1229,N_21362,N_21617);
nand UO_1230 (O_1230,N_21939,N_20683);
nand UO_1231 (O_1231,N_24600,N_23519);
nor UO_1232 (O_1232,N_23164,N_20875);
nor UO_1233 (O_1233,N_20375,N_20446);
nor UO_1234 (O_1234,N_20695,N_24110);
or UO_1235 (O_1235,N_20830,N_22264);
and UO_1236 (O_1236,N_23792,N_23031);
nor UO_1237 (O_1237,N_21679,N_24560);
nand UO_1238 (O_1238,N_22652,N_23435);
nor UO_1239 (O_1239,N_24136,N_20142);
nand UO_1240 (O_1240,N_21464,N_20450);
and UO_1241 (O_1241,N_22607,N_20443);
nand UO_1242 (O_1242,N_23956,N_20084);
or UO_1243 (O_1243,N_21924,N_23458);
or UO_1244 (O_1244,N_21357,N_20836);
nor UO_1245 (O_1245,N_21161,N_24117);
or UO_1246 (O_1246,N_20601,N_23304);
and UO_1247 (O_1247,N_22952,N_20773);
xor UO_1248 (O_1248,N_22618,N_21965);
xor UO_1249 (O_1249,N_23927,N_20895);
nand UO_1250 (O_1250,N_21582,N_23620);
nand UO_1251 (O_1251,N_24464,N_20130);
nor UO_1252 (O_1252,N_22662,N_21649);
and UO_1253 (O_1253,N_24281,N_21314);
nor UO_1254 (O_1254,N_22080,N_22250);
nand UO_1255 (O_1255,N_22441,N_23533);
xnor UO_1256 (O_1256,N_23203,N_22316);
xor UO_1257 (O_1257,N_24296,N_20210);
xnor UO_1258 (O_1258,N_20550,N_22149);
or UO_1259 (O_1259,N_20275,N_23675);
nand UO_1260 (O_1260,N_21350,N_22079);
nand UO_1261 (O_1261,N_21030,N_23462);
or UO_1262 (O_1262,N_20497,N_24359);
xnor UO_1263 (O_1263,N_21082,N_24644);
nor UO_1264 (O_1264,N_24220,N_21374);
nor UO_1265 (O_1265,N_21038,N_24365);
nor UO_1266 (O_1266,N_22823,N_24267);
and UO_1267 (O_1267,N_22591,N_24623);
nor UO_1268 (O_1268,N_23171,N_23303);
xnor UO_1269 (O_1269,N_24657,N_24263);
and UO_1270 (O_1270,N_22308,N_20059);
and UO_1271 (O_1271,N_21375,N_20546);
or UO_1272 (O_1272,N_24163,N_22856);
and UO_1273 (O_1273,N_24029,N_21833);
nand UO_1274 (O_1274,N_20152,N_23103);
xnor UO_1275 (O_1275,N_24820,N_24204);
nand UO_1276 (O_1276,N_22340,N_23508);
nand UO_1277 (O_1277,N_23425,N_20219);
nor UO_1278 (O_1278,N_22919,N_22248);
nor UO_1279 (O_1279,N_21294,N_23246);
and UO_1280 (O_1280,N_21398,N_20745);
nand UO_1281 (O_1281,N_20846,N_24269);
nor UO_1282 (O_1282,N_23712,N_21851);
nand UO_1283 (O_1283,N_21663,N_22834);
and UO_1284 (O_1284,N_21899,N_20809);
and UO_1285 (O_1285,N_21803,N_24513);
or UO_1286 (O_1286,N_20761,N_21124);
or UO_1287 (O_1287,N_24735,N_23233);
or UO_1288 (O_1288,N_22200,N_20717);
or UO_1289 (O_1289,N_21849,N_20628);
nand UO_1290 (O_1290,N_21447,N_21109);
xnor UO_1291 (O_1291,N_23250,N_22342);
and UO_1292 (O_1292,N_22053,N_24333);
or UO_1293 (O_1293,N_23277,N_23697);
nand UO_1294 (O_1294,N_23926,N_24483);
or UO_1295 (O_1295,N_22225,N_23569);
or UO_1296 (O_1296,N_23831,N_21431);
nor UO_1297 (O_1297,N_24844,N_23983);
xnor UO_1298 (O_1298,N_23905,N_23805);
or UO_1299 (O_1299,N_20748,N_23357);
nor UO_1300 (O_1300,N_21485,N_23082);
and UO_1301 (O_1301,N_24121,N_24406);
xor UO_1302 (O_1302,N_24565,N_24444);
xnor UO_1303 (O_1303,N_22062,N_22718);
nor UO_1304 (O_1304,N_24864,N_21948);
or UO_1305 (O_1305,N_23726,N_22758);
nand UO_1306 (O_1306,N_20240,N_20638);
nand UO_1307 (O_1307,N_24851,N_21270);
or UO_1308 (O_1308,N_22503,N_22348);
nor UO_1309 (O_1309,N_20576,N_22245);
xor UO_1310 (O_1310,N_20696,N_24339);
nor UO_1311 (O_1311,N_23601,N_21367);
xor UO_1312 (O_1312,N_22523,N_24501);
nor UO_1313 (O_1313,N_24119,N_23642);
and UO_1314 (O_1314,N_24225,N_21266);
nor UO_1315 (O_1315,N_22168,N_24199);
and UO_1316 (O_1316,N_21591,N_22703);
nand UO_1317 (O_1317,N_23647,N_23896);
and UO_1318 (O_1318,N_24294,N_20832);
xor UO_1319 (O_1319,N_24506,N_21326);
xor UO_1320 (O_1320,N_21523,N_23729);
nand UO_1321 (O_1321,N_23062,N_22937);
or UO_1322 (O_1322,N_23897,N_21094);
nand UO_1323 (O_1323,N_22984,N_22933);
nor UO_1324 (O_1324,N_20365,N_24773);
nand UO_1325 (O_1325,N_23592,N_20536);
nor UO_1326 (O_1326,N_24094,N_22579);
and UO_1327 (O_1327,N_21581,N_20941);
nand UO_1328 (O_1328,N_21493,N_20856);
nand UO_1329 (O_1329,N_20002,N_20993);
nor UO_1330 (O_1330,N_24543,N_24976);
nor UO_1331 (O_1331,N_20416,N_20533);
or UO_1332 (O_1332,N_24472,N_22678);
nor UO_1333 (O_1333,N_21209,N_21253);
and UO_1334 (O_1334,N_22641,N_21479);
nand UO_1335 (O_1335,N_23943,N_22532);
nor UO_1336 (O_1336,N_23721,N_22194);
xnor UO_1337 (O_1337,N_22821,N_21171);
or UO_1338 (O_1338,N_20825,N_23405);
nand UO_1339 (O_1339,N_22753,N_24364);
xnor UO_1340 (O_1340,N_22621,N_23460);
or UO_1341 (O_1341,N_22439,N_22713);
or UO_1342 (O_1342,N_22228,N_23430);
or UO_1343 (O_1343,N_20513,N_24373);
nor UO_1344 (O_1344,N_23667,N_21331);
nand UO_1345 (O_1345,N_23718,N_20749);
nand UO_1346 (O_1346,N_21041,N_22576);
or UO_1347 (O_1347,N_24405,N_20184);
and UO_1348 (O_1348,N_21480,N_23351);
xnor UO_1349 (O_1349,N_20482,N_22682);
or UO_1350 (O_1350,N_20977,N_22193);
nor UO_1351 (O_1351,N_20388,N_24985);
and UO_1352 (O_1352,N_20297,N_22733);
nor UO_1353 (O_1353,N_21843,N_22218);
and UO_1354 (O_1354,N_23032,N_23259);
or UO_1355 (O_1355,N_22134,N_24017);
nand UO_1356 (O_1356,N_23126,N_23977);
nor UO_1357 (O_1357,N_22272,N_23189);
and UO_1358 (O_1358,N_23087,N_20364);
nand UO_1359 (O_1359,N_23264,N_23507);
or UO_1360 (O_1360,N_21247,N_20808);
and UO_1361 (O_1361,N_21143,N_23557);
xnor UO_1362 (O_1362,N_22739,N_24638);
or UO_1363 (O_1363,N_21557,N_23763);
or UO_1364 (O_1364,N_20699,N_24152);
and UO_1365 (O_1365,N_20379,N_20594);
or UO_1366 (O_1366,N_23953,N_20150);
or UO_1367 (O_1367,N_20845,N_23394);
and UO_1368 (O_1368,N_20165,N_24411);
or UO_1369 (O_1369,N_20093,N_20099);
xor UO_1370 (O_1370,N_23020,N_20541);
nor UO_1371 (O_1371,N_20552,N_22113);
nand UO_1372 (O_1372,N_24529,N_22451);
and UO_1373 (O_1373,N_23129,N_20174);
or UO_1374 (O_1374,N_24104,N_21122);
nor UO_1375 (O_1375,N_23964,N_21072);
or UO_1376 (O_1376,N_22594,N_23800);
and UO_1377 (O_1377,N_24603,N_20713);
nand UO_1378 (O_1378,N_24958,N_21762);
nor UO_1379 (O_1379,N_21906,N_21439);
nand UO_1380 (O_1380,N_20319,N_22314);
and UO_1381 (O_1381,N_24544,N_23866);
nand UO_1382 (O_1382,N_22946,N_24918);
or UO_1383 (O_1383,N_24022,N_24238);
nand UO_1384 (O_1384,N_20021,N_20623);
xor UO_1385 (O_1385,N_23608,N_20318);
or UO_1386 (O_1386,N_20320,N_23796);
nand UO_1387 (O_1387,N_24870,N_21953);
and UO_1388 (O_1388,N_21620,N_21403);
xor UO_1389 (O_1389,N_23918,N_21883);
or UO_1390 (O_1390,N_21014,N_22719);
xor UO_1391 (O_1391,N_23208,N_22764);
nand UO_1392 (O_1392,N_22402,N_22585);
and UO_1393 (O_1393,N_20839,N_21868);
and UO_1394 (O_1394,N_23095,N_20983);
nand UO_1395 (O_1395,N_23537,N_20998);
and UO_1396 (O_1396,N_21460,N_21511);
nand UO_1397 (O_1397,N_22409,N_24059);
or UO_1398 (O_1398,N_21740,N_20763);
or UO_1399 (O_1399,N_20540,N_23793);
xnor UO_1400 (O_1400,N_21315,N_24488);
nor UO_1401 (O_1401,N_21052,N_21292);
nand UO_1402 (O_1402,N_23708,N_22721);
nand UO_1403 (O_1403,N_21254,N_21342);
nand UO_1404 (O_1404,N_22936,N_23952);
nand UO_1405 (O_1405,N_22433,N_22926);
nor UO_1406 (O_1406,N_23576,N_20263);
nand UO_1407 (O_1407,N_20965,N_23877);
nand UO_1408 (O_1408,N_23155,N_24186);
and UO_1409 (O_1409,N_24452,N_24653);
nor UO_1410 (O_1410,N_24183,N_21093);
xnor UO_1411 (O_1411,N_23312,N_20979);
xor UO_1412 (O_1412,N_20229,N_22900);
or UO_1413 (O_1413,N_23600,N_23937);
nor UO_1414 (O_1414,N_24016,N_22658);
and UO_1415 (O_1415,N_21008,N_21071);
and UO_1416 (O_1416,N_24368,N_22956);
nand UO_1417 (O_1417,N_23280,N_21876);
or UO_1418 (O_1418,N_24033,N_20106);
or UO_1419 (O_1419,N_20753,N_23941);
and UO_1420 (O_1420,N_20544,N_21088);
and UO_1421 (O_1421,N_21291,N_24497);
nor UO_1422 (O_1422,N_20532,N_23542);
xnor UO_1423 (O_1423,N_23076,N_21929);
and UO_1424 (O_1424,N_22305,N_24140);
xnor UO_1425 (O_1425,N_23745,N_23283);
or UO_1426 (O_1426,N_24252,N_22206);
nand UO_1427 (O_1427,N_24671,N_23181);
and UO_1428 (O_1428,N_23846,N_20834);
or UO_1429 (O_1429,N_21863,N_22107);
nor UO_1430 (O_1430,N_20881,N_20719);
nor UO_1431 (O_1431,N_21411,N_20951);
or UO_1432 (O_1432,N_22390,N_24217);
and UO_1433 (O_1433,N_20521,N_22865);
nor UO_1434 (O_1434,N_23680,N_23950);
nor UO_1435 (O_1435,N_23572,N_24519);
nand UO_1436 (O_1436,N_22404,N_21045);
nand UO_1437 (O_1437,N_23006,N_24751);
or UO_1438 (O_1438,N_22839,N_21197);
xor UO_1439 (O_1439,N_22741,N_21106);
or UO_1440 (O_1440,N_23154,N_22729);
nor UO_1441 (O_1441,N_22550,N_21584);
nand UO_1442 (O_1442,N_20222,N_23160);
nand UO_1443 (O_1443,N_23204,N_22413);
or UO_1444 (O_1444,N_21021,N_21068);
or UO_1445 (O_1445,N_23848,N_22599);
nor UO_1446 (O_1446,N_21089,N_20667);
and UO_1447 (O_1447,N_22663,N_20205);
xnor UO_1448 (O_1448,N_20804,N_22526);
or UO_1449 (O_1449,N_24809,N_21545);
and UO_1450 (O_1450,N_20936,N_21532);
or UO_1451 (O_1451,N_21898,N_24502);
nand UO_1452 (O_1452,N_23240,N_20457);
and UO_1453 (O_1453,N_21622,N_23996);
and UO_1454 (O_1454,N_23070,N_21825);
or UO_1455 (O_1455,N_20487,N_23288);
or UO_1456 (O_1456,N_22596,N_21436);
xnor UO_1457 (O_1457,N_20614,N_24477);
nand UO_1458 (O_1458,N_24998,N_21537);
xor UO_1459 (O_1459,N_21873,N_20946);
or UO_1460 (O_1460,N_23598,N_21956);
nor UO_1461 (O_1461,N_23924,N_23060);
nor UO_1462 (O_1462,N_20616,N_21459);
nand UO_1463 (O_1463,N_22138,N_21186);
nand UO_1464 (O_1464,N_22452,N_21542);
and UO_1465 (O_1465,N_23851,N_22906);
nand UO_1466 (O_1466,N_21432,N_23665);
nor UO_1467 (O_1467,N_22613,N_24231);
nand UO_1468 (O_1468,N_22365,N_22822);
nand UO_1469 (O_1469,N_24247,N_22637);
xor UO_1470 (O_1470,N_23850,N_21556);
or UO_1471 (O_1471,N_23979,N_21980);
nand UO_1472 (O_1472,N_20620,N_22868);
and UO_1473 (O_1473,N_20046,N_20640);
nand UO_1474 (O_1474,N_24241,N_21987);
or UO_1475 (O_1475,N_21172,N_24268);
nand UO_1476 (O_1476,N_21390,N_24997);
nor UO_1477 (O_1477,N_23223,N_23789);
and UO_1478 (O_1478,N_22145,N_24170);
nor UO_1479 (O_1479,N_20769,N_21923);
or UO_1480 (O_1480,N_20015,N_20618);
or UO_1481 (O_1481,N_20956,N_22818);
nor UO_1482 (O_1482,N_23229,N_23992);
xor UO_1483 (O_1483,N_21240,N_22614);
or UO_1484 (O_1484,N_21127,N_23646);
nor UO_1485 (O_1485,N_23375,N_21055);
nand UO_1486 (O_1486,N_20603,N_22297);
nand UO_1487 (O_1487,N_22584,N_24989);
nand UO_1488 (O_1488,N_22610,N_24064);
nand UO_1489 (O_1489,N_24044,N_23504);
and UO_1490 (O_1490,N_20693,N_21569);
and UO_1491 (O_1491,N_22068,N_21496);
nor UO_1492 (O_1492,N_24187,N_21988);
and UO_1493 (O_1493,N_20101,N_22323);
nor UO_1494 (O_1494,N_24887,N_20675);
nor UO_1495 (O_1495,N_23456,N_21999);
nor UO_1496 (O_1496,N_23376,N_23984);
or UO_1497 (O_1497,N_23469,N_23258);
nor UO_1498 (O_1498,N_21469,N_23863);
or UO_1499 (O_1499,N_24299,N_20726);
nand UO_1500 (O_1500,N_23041,N_20583);
and UO_1501 (O_1501,N_21004,N_22398);
nand UO_1502 (O_1502,N_24065,N_22102);
nor UO_1503 (O_1503,N_21991,N_23961);
nand UO_1504 (O_1504,N_22848,N_24678);
and UO_1505 (O_1505,N_24960,N_23638);
nor UO_1506 (O_1506,N_21160,N_20049);
nor UO_1507 (O_1507,N_20885,N_23522);
or UO_1508 (O_1508,N_23480,N_24829);
and UO_1509 (O_1509,N_23582,N_23999);
nor UO_1510 (O_1510,N_24340,N_23652);
nand UO_1511 (O_1511,N_21135,N_20284);
or UO_1512 (O_1512,N_21888,N_22013);
and UO_1513 (O_1513,N_24362,N_22890);
nor UO_1514 (O_1514,N_23061,N_21757);
or UO_1515 (O_1515,N_21780,N_22457);
nand UO_1516 (O_1516,N_22131,N_22918);
nand UO_1517 (O_1517,N_24790,N_21113);
or UO_1518 (O_1518,N_20888,N_22860);
nand UO_1519 (O_1519,N_22259,N_21961);
or UO_1520 (O_1520,N_22333,N_20114);
or UO_1521 (O_1521,N_24130,N_23336);
nand UO_1522 (O_1522,N_20234,N_24318);
nand UO_1523 (O_1523,N_20468,N_22117);
or UO_1524 (O_1524,N_22781,N_23562);
or UO_1525 (O_1525,N_24580,N_21392);
xnor UO_1526 (O_1526,N_23771,N_24778);
nand UO_1527 (O_1527,N_24054,N_21669);
and UO_1528 (O_1528,N_22568,N_20344);
nor UO_1529 (O_1529,N_22313,N_24342);
and UO_1530 (O_1530,N_23543,N_24213);
nor UO_1531 (O_1531,N_20617,N_22172);
and UO_1532 (O_1532,N_21064,N_23496);
or UO_1533 (O_1533,N_20209,N_21425);
xnor UO_1534 (O_1534,N_22847,N_21723);
or UO_1535 (O_1535,N_23067,N_20432);
xor UO_1536 (O_1536,N_22188,N_24335);
and UO_1537 (O_1537,N_24162,N_22072);
or UO_1538 (O_1538,N_24479,N_22001);
nand UO_1539 (O_1539,N_24596,N_23881);
or UO_1540 (O_1540,N_22617,N_20238);
nor UO_1541 (O_1541,N_24006,N_23199);
or UO_1542 (O_1542,N_20584,N_24869);
or UO_1543 (O_1543,N_20016,N_22907);
nor UO_1544 (O_1544,N_22498,N_20625);
or UO_1545 (O_1545,N_20714,N_22443);
xor UO_1546 (O_1546,N_21169,N_21524);
or UO_1547 (O_1547,N_24349,N_22531);
nand UO_1548 (O_1548,N_23377,N_24131);
or UO_1549 (O_1549,N_24309,N_21809);
or UO_1550 (O_1550,N_21777,N_21430);
and UO_1551 (O_1551,N_21878,N_24397);
or UO_1552 (O_1552,N_22063,N_21536);
nand UO_1553 (O_1553,N_21423,N_24703);
nor UO_1554 (O_1554,N_23385,N_21299);
or UO_1555 (O_1555,N_22930,N_23444);
nand UO_1556 (O_1556,N_20086,N_20032);
or UO_1557 (O_1557,N_23015,N_23237);
or UO_1558 (O_1558,N_21226,N_21420);
nand UO_1559 (O_1559,N_22851,N_22156);
nand UO_1560 (O_1560,N_20923,N_22306);
or UO_1561 (O_1561,N_20406,N_21702);
and UO_1562 (O_1562,N_22130,N_24786);
and UO_1563 (O_1563,N_20261,N_24995);
and UO_1564 (O_1564,N_23868,N_22685);
nand UO_1565 (O_1565,N_21087,N_23071);
and UO_1566 (O_1566,N_21130,N_20358);
nor UO_1567 (O_1567,N_21789,N_20476);
and UO_1568 (O_1568,N_22375,N_23445);
nand UO_1569 (O_1569,N_20823,N_21293);
and UO_1570 (O_1570,N_24757,N_24198);
nand UO_1571 (O_1571,N_20069,N_20129);
or UO_1572 (O_1572,N_22034,N_23068);
and UO_1573 (O_1573,N_24190,N_24380);
or UO_1574 (O_1574,N_21399,N_23829);
nand UO_1575 (O_1575,N_21716,N_20524);
or UO_1576 (O_1576,N_22557,N_20419);
nand UO_1577 (O_1577,N_20815,N_23874);
nand UO_1578 (O_1578,N_22595,N_21049);
nor UO_1579 (O_1579,N_24023,N_23757);
and UO_1580 (O_1580,N_23198,N_22044);
xnor UO_1581 (O_1581,N_20489,N_23783);
nor UO_1582 (O_1582,N_20231,N_23515);
xnor UO_1583 (O_1583,N_20267,N_21310);
nand UO_1584 (O_1584,N_20535,N_20950);
or UO_1585 (O_1585,N_24705,N_20920);
and UO_1586 (O_1586,N_21433,N_21001);
nor UO_1587 (O_1587,N_20109,N_21339);
or UO_1588 (O_1588,N_23914,N_24313);
nor UO_1589 (O_1589,N_23641,N_20622);
nor UO_1590 (O_1590,N_23990,N_21316);
or UO_1591 (O_1591,N_21640,N_20715);
xor UO_1592 (O_1592,N_20922,N_20287);
or UO_1593 (O_1593,N_24446,N_21073);
and UO_1594 (O_1594,N_20051,N_20370);
nor UO_1595 (O_1595,N_22199,N_20682);
nand UO_1596 (O_1596,N_20474,N_20461);
or UO_1597 (O_1597,N_24273,N_22410);
xor UO_1598 (O_1598,N_21000,N_23098);
nor UO_1599 (O_1599,N_20075,N_22118);
and UO_1600 (O_1600,N_24062,N_21235);
and UO_1601 (O_1601,N_23902,N_23403);
or UO_1602 (O_1602,N_20952,N_24557);
or UO_1603 (O_1603,N_24742,N_21639);
nand UO_1604 (O_1604,N_24761,N_23965);
or UO_1605 (O_1605,N_22680,N_20994);
or UO_1606 (O_1606,N_21442,N_21462);
and UO_1607 (O_1607,N_20607,N_23217);
or UO_1608 (O_1608,N_21328,N_23302);
and UO_1609 (O_1609,N_24437,N_20233);
nand UO_1610 (O_1610,N_22128,N_24695);
xnor UO_1611 (O_1611,N_20141,N_24764);
xnor UO_1612 (O_1612,N_21205,N_20235);
xor UO_1613 (O_1613,N_21968,N_24244);
or UO_1614 (O_1614,N_22407,N_22843);
xnor UO_1615 (O_1615,N_22745,N_24718);
nand UO_1616 (O_1616,N_23998,N_23884);
nor UO_1617 (O_1617,N_23506,N_22162);
or UO_1618 (O_1618,N_24298,N_20394);
and UO_1619 (O_1619,N_22609,N_24053);
nand UO_1620 (O_1620,N_24052,N_22502);
nor UO_1621 (O_1621,N_21397,N_23056);
nor UO_1622 (O_1622,N_22490,N_21400);
or UO_1623 (O_1623,N_21391,N_23817);
nor UO_1624 (O_1624,N_21181,N_23363);
nand UO_1625 (O_1625,N_24586,N_23367);
or UO_1626 (O_1626,N_21421,N_22475);
nor UO_1627 (O_1627,N_20635,N_23387);
and UO_1628 (O_1628,N_23511,N_21159);
nand UO_1629 (O_1629,N_20366,N_20906);
nor UO_1630 (O_1630,N_21150,N_20480);
xor UO_1631 (O_1631,N_23492,N_24691);
or UO_1632 (O_1632,N_24537,N_20679);
nor UO_1633 (O_1633,N_23485,N_24038);
or UO_1634 (O_1634,N_24355,N_21044);
nor UO_1635 (O_1635,N_20135,N_24933);
nor UO_1636 (O_1636,N_23554,N_21658);
and UO_1637 (O_1637,N_20448,N_23546);
or UO_1638 (O_1638,N_20421,N_24606);
nand UO_1639 (O_1639,N_24618,N_20855);
nand UO_1640 (O_1640,N_21102,N_21499);
nor UO_1641 (O_1641,N_21422,N_22850);
nor UO_1642 (O_1642,N_20542,N_20975);
nor UO_1643 (O_1643,N_23614,N_22979);
nor UO_1644 (O_1644,N_21840,N_21614);
and UO_1645 (O_1645,N_23276,N_20957);
and UO_1646 (O_1646,N_24020,N_21852);
nor UO_1647 (O_1647,N_22240,N_20711);
nand UO_1648 (O_1648,N_22608,N_20651);
xor UO_1649 (O_1649,N_20371,N_21040);
nor UO_1650 (O_1650,N_22082,N_20178);
xor UO_1651 (O_1651,N_20921,N_21516);
nand UO_1652 (O_1652,N_22804,N_23637);
or UO_1653 (O_1653,N_22912,N_21417);
and UO_1654 (O_1654,N_22005,N_23748);
or UO_1655 (O_1655,N_21095,N_22706);
and UO_1656 (O_1656,N_24701,N_23183);
and UO_1657 (O_1657,N_22181,N_23400);
nand UO_1658 (O_1658,N_23536,N_24344);
nor UO_1659 (O_1659,N_23635,N_21012);
nor UO_1660 (O_1660,N_22022,N_21097);
nand UO_1661 (O_1661,N_20633,N_23705);
and UO_1662 (O_1662,N_21117,N_20826);
xor UO_1663 (O_1663,N_23052,N_22913);
and UO_1664 (O_1664,N_24147,N_22817);
and UO_1665 (O_1665,N_23549,N_24508);
nor UO_1666 (O_1666,N_23101,N_21866);
or UO_1667 (O_1667,N_22258,N_20224);
nand UO_1668 (O_1668,N_24255,N_20735);
xnor UO_1669 (O_1669,N_21268,N_24551);
or UO_1670 (O_1670,N_24687,N_21162);
nor UO_1671 (O_1671,N_22212,N_21396);
nand UO_1672 (O_1672,N_20256,N_20117);
or UO_1673 (O_1673,N_23413,N_21365);
and UO_1674 (O_1674,N_22177,N_23404);
nand UO_1675 (O_1675,N_21332,N_21107);
and UO_1676 (O_1676,N_23310,N_23256);
or UO_1677 (O_1677,N_23776,N_22716);
and UO_1678 (O_1678,N_21330,N_23765);
xnor UO_1679 (O_1679,N_24766,N_24189);
nor UO_1680 (O_1680,N_22700,N_20103);
nor UO_1681 (O_1681,N_24505,N_24913);
and UO_1682 (O_1682,N_23414,N_20582);
nand UO_1683 (O_1683,N_20304,N_22707);
or UO_1684 (O_1684,N_22505,N_23224);
and UO_1685 (O_1685,N_21737,N_24107);
xnor UO_1686 (O_1686,N_22236,N_24050);
or UO_1687 (O_1687,N_23993,N_22928);
nand UO_1688 (O_1688,N_22320,N_24425);
nor UO_1689 (O_1689,N_22447,N_21039);
nand UO_1690 (O_1690,N_21200,N_21101);
or UO_1691 (O_1691,N_22421,N_24430);
xor UO_1692 (O_1692,N_21848,N_21560);
nand UO_1693 (O_1693,N_20662,N_24249);
nand UO_1694 (O_1694,N_21841,N_20387);
or UO_1695 (O_1695,N_21616,N_22444);
nand UO_1696 (O_1696,N_24077,N_22221);
nor UO_1697 (O_1697,N_23215,N_22290);
and UO_1698 (O_1698,N_24245,N_24060);
nor UO_1699 (O_1699,N_24146,N_21558);
or UO_1700 (O_1700,N_23613,N_22625);
nand UO_1701 (O_1701,N_23682,N_20242);
or UO_1702 (O_1702,N_21862,N_20022);
nand UO_1703 (O_1703,N_20159,N_23666);
nor UO_1704 (O_1704,N_21046,N_20372);
nand UO_1705 (O_1705,N_21363,N_20285);
xnor UO_1706 (O_1706,N_24689,N_21745);
nand UO_1707 (O_1707,N_20561,N_24892);
nand UO_1708 (O_1708,N_20030,N_20232);
nor UO_1709 (O_1709,N_23230,N_20190);
xor UO_1710 (O_1710,N_21434,N_22824);
and UO_1711 (O_1711,N_22774,N_20087);
and UO_1712 (O_1712,N_24091,N_24271);
xnor UO_1713 (O_1713,N_23475,N_22711);
nand UO_1714 (O_1714,N_24884,N_20399);
xnor UO_1715 (O_1715,N_21601,N_22091);
nand UO_1716 (O_1716,N_24983,N_22886);
xnor UO_1717 (O_1717,N_20639,N_21718);
nor UO_1718 (O_1718,N_22229,N_22086);
and UO_1719 (O_1719,N_24524,N_22381);
nand UO_1720 (O_1720,N_21168,N_20475);
or UO_1721 (O_1721,N_23779,N_21241);
nor UO_1722 (O_1722,N_24879,N_22636);
nand UO_1723 (O_1723,N_24946,N_20470);
nor UO_1724 (O_1724,N_22110,N_20948);
nor UO_1725 (O_1725,N_24707,N_20567);
nor UO_1726 (O_1726,N_20940,N_22545);
nor UO_1727 (O_1727,N_23356,N_23917);
nand UO_1728 (O_1728,N_24080,N_21667);
and UO_1729 (O_1729,N_24789,N_24369);
nor UO_1730 (O_1730,N_20571,N_21695);
nand UO_1731 (O_1731,N_24467,N_22862);
nand UO_1732 (O_1732,N_20395,N_23692);
and UO_1733 (O_1733,N_20539,N_23383);
nor UO_1734 (O_1734,N_20226,N_23321);
nand UO_1735 (O_1735,N_22582,N_21645);
or UO_1736 (O_1736,N_20288,N_20668);
and UO_1737 (O_1737,N_23077,N_22205);
xnor UO_1738 (O_1738,N_21739,N_21660);
xnor UO_1739 (O_1739,N_20081,N_24845);
nand UO_1740 (O_1740,N_20677,N_22932);
nand UO_1741 (O_1741,N_23316,N_20042);
nor UO_1742 (O_1742,N_24447,N_21237);
or UO_1743 (O_1743,N_20043,N_24992);
nand UO_1744 (O_1744,N_23781,N_24521);
or UO_1745 (O_1745,N_21288,N_24652);
and UO_1746 (O_1746,N_24316,N_24522);
nor UO_1747 (O_1747,N_20730,N_20252);
and UO_1748 (O_1748,N_24073,N_23933);
nor UO_1749 (O_1749,N_23093,N_22366);
nor UO_1750 (O_1750,N_23947,N_21203);
nor UO_1751 (O_1751,N_23249,N_20380);
nand UO_1752 (O_1752,N_24015,N_23173);
nand UO_1753 (O_1753,N_20548,N_20410);
and UO_1754 (O_1754,N_24233,N_20525);
and UO_1755 (O_1755,N_21627,N_24785);
xor UO_1756 (O_1756,N_22065,N_22681);
or UO_1757 (O_1757,N_20437,N_23345);
and UO_1758 (O_1758,N_23411,N_24426);
nor UO_1759 (O_1759,N_24641,N_22751);
nor UO_1760 (O_1760,N_24070,N_23849);
nand UO_1761 (O_1761,N_20666,N_22047);
or UO_1762 (O_1762,N_24496,N_20518);
or UO_1763 (O_1763,N_21613,N_20343);
xor UO_1764 (O_1764,N_20774,N_24788);
nor UO_1765 (O_1765,N_21090,N_20149);
or UO_1766 (O_1766,N_21069,N_20530);
or UO_1767 (O_1767,N_23343,N_21467);
or UO_1768 (O_1768,N_23921,N_23328);
nand UO_1769 (O_1769,N_20504,N_21871);
and UO_1770 (O_1770,N_21318,N_24545);
nand UO_1771 (O_1771,N_23308,N_21149);
or UO_1772 (O_1772,N_23790,N_21865);
xor UO_1773 (O_1773,N_21031,N_22536);
xnor UO_1774 (O_1774,N_20897,N_24627);
xor UO_1775 (O_1775,N_21429,N_22592);
or UO_1776 (O_1776,N_23017,N_22009);
or UO_1777 (O_1777,N_24075,N_22103);
nor UO_1778 (O_1778,N_24092,N_22455);
xnor UO_1779 (O_1779,N_20820,N_22180);
and UO_1780 (O_1780,N_23746,N_21512);
and UO_1781 (O_1781,N_20793,N_20110);
or UO_1782 (O_1782,N_21794,N_22646);
nand UO_1783 (O_1783,N_21123,N_22838);
or UO_1784 (O_1784,N_23658,N_21715);
and UO_1785 (O_1785,N_20538,N_23428);
nand UO_1786 (O_1786,N_21218,N_24907);
or UO_1787 (O_1787,N_22277,N_21931);
xnor UO_1788 (O_1788,N_22491,N_21007);
nand UO_1789 (O_1789,N_24232,N_22049);
nor UO_1790 (O_1790,N_21552,N_24914);
and UO_1791 (O_1791,N_23466,N_21982);
nor UO_1792 (O_1792,N_23865,N_21760);
xor UO_1793 (O_1793,N_22420,N_24862);
or UO_1794 (O_1794,N_22769,N_20659);
nand UO_1795 (O_1795,N_22792,N_22244);
nand UO_1796 (O_1796,N_22372,N_23148);
nor UO_1797 (O_1797,N_20919,N_20893);
xor UO_1798 (O_1798,N_20942,N_24710);
and UO_1799 (O_1799,N_24495,N_20020);
nor UO_1800 (O_1800,N_23359,N_21808);
or UO_1801 (O_1801,N_21990,N_24950);
or UO_1802 (O_1802,N_23003,N_20577);
xnor UO_1803 (O_1803,N_20926,N_20064);
and UO_1804 (O_1804,N_24449,N_24061);
xor UO_1805 (O_1805,N_21076,N_24615);
nor UO_1806 (O_1806,N_22484,N_22028);
nor UO_1807 (O_1807,N_22385,N_20779);
nand UO_1808 (O_1808,N_23671,N_23170);
and UO_1809 (O_1809,N_21002,N_24261);
and UO_1810 (O_1810,N_20067,N_20334);
or UO_1811 (O_1811,N_20516,N_21379);
nand UO_1812 (O_1812,N_20070,N_20161);
nor UO_1813 (O_1813,N_22288,N_20566);
or UO_1814 (O_1814,N_20467,N_21983);
xor UO_1815 (O_1815,N_20935,N_22987);
or UO_1816 (O_1816,N_21037,N_20303);
nand UO_1817 (O_1817,N_21661,N_23122);
nand UO_1818 (O_1818,N_21470,N_20902);
nor UO_1819 (O_1819,N_21711,N_20376);
and UO_1820 (O_1820,N_22667,N_22939);
nand UO_1821 (O_1821,N_24572,N_22020);
nor UO_1822 (O_1822,N_21720,N_21210);
or UO_1823 (O_1823,N_21199,N_24484);
nor UO_1824 (O_1824,N_23169,N_23517);
nand UO_1825 (O_1825,N_21277,N_21541);
nor UO_1826 (O_1826,N_21909,N_24043);
nand UO_1827 (O_1827,N_22105,N_23330);
and UO_1828 (O_1828,N_23814,N_22986);
xnor UO_1829 (O_1829,N_22007,N_24021);
and UO_1830 (O_1830,N_23862,N_22881);
or UO_1831 (O_1831,N_20193,N_20862);
and UO_1832 (O_1832,N_24699,N_23281);
nor UO_1833 (O_1833,N_22060,N_24793);
xnor UO_1834 (O_1834,N_23014,N_21861);
nand UO_1835 (O_1835,N_23427,N_23088);
nor UO_1836 (O_1836,N_21274,N_23161);
nor UO_1837 (O_1837,N_21085,N_20982);
nor UO_1838 (O_1838,N_21359,N_21140);
or UO_1839 (O_1839,N_24466,N_20654);
and UO_1840 (O_1840,N_22377,N_20560);
and UO_1841 (O_1841,N_22418,N_21563);
nor UO_1842 (O_1842,N_23226,N_22084);
and UO_1843 (O_1843,N_24103,N_21728);
nor UO_1844 (O_1844,N_20094,N_22085);
or UO_1845 (O_1845,N_22575,N_22600);
and UO_1846 (O_1846,N_24262,N_23589);
xor UO_1847 (O_1847,N_22555,N_24001);
xor UO_1848 (O_1848,N_24079,N_22249);
nor UO_1849 (O_1849,N_20426,N_21005);
and UO_1850 (O_1850,N_20478,N_24137);
nand UO_1851 (O_1851,N_22958,N_22612);
and UO_1852 (O_1852,N_20283,N_23585);
or UO_1853 (O_1853,N_20974,N_24445);
and UO_1854 (O_1854,N_23272,N_24767);
nand UO_1855 (O_1855,N_22560,N_23632);
nor UO_1856 (O_1856,N_22971,N_24799);
nor UO_1857 (O_1857,N_23659,N_22427);
nor UO_1858 (O_1858,N_22073,N_20627);
nand UO_1859 (O_1859,N_23145,N_20168);
nand UO_1860 (O_1860,N_20286,N_24000);
nor UO_1861 (O_1861,N_21345,N_23337);
or UO_1862 (O_1862,N_23407,N_22626);
nand UO_1863 (O_1863,N_21178,N_21630);
or UO_1864 (O_1864,N_23624,N_24258);
nand UO_1865 (O_1865,N_20772,N_21894);
or UO_1866 (O_1866,N_22458,N_21850);
nor UO_1867 (O_1867,N_21513,N_23758);
nand UO_1868 (O_1868,N_23991,N_22910);
and UO_1869 (O_1869,N_21207,N_22934);
or UO_1870 (O_1870,N_24876,N_21368);
or UO_1871 (O_1871,N_21945,N_20905);
nand UO_1872 (O_1872,N_21918,N_21904);
nand UO_1873 (O_1873,N_21587,N_20775);
or UO_1874 (O_1874,N_24089,N_20637);
and UO_1875 (O_1875,N_21531,N_24835);
and UO_1876 (O_1876,N_23903,N_24926);
nand UO_1877 (O_1877,N_22463,N_22763);
nand UO_1878 (O_1878,N_23860,N_22874);
nand UO_1879 (O_1879,N_22914,N_21510);
xor UO_1880 (O_1880,N_20241,N_20393);
and UO_1881 (O_1881,N_23207,N_22738);
nand UO_1882 (O_1882,N_24840,N_24646);
nand UO_1883 (O_1883,N_20369,N_21063);
and UO_1884 (O_1884,N_22773,N_23599);
nand UO_1885 (O_1885,N_21761,N_23361);
nand UO_1886 (O_1886,N_23443,N_20634);
xor UO_1887 (O_1887,N_24581,N_20563);
or UO_1888 (O_1888,N_23402,N_22728);
nor UO_1889 (O_1889,N_24095,N_24074);
nor UO_1890 (O_1890,N_24647,N_23084);
or UO_1891 (O_1891,N_24133,N_24979);
or UO_1892 (O_1892,N_20971,N_24752);
nor UO_1893 (O_1893,N_23528,N_23994);
and UO_1894 (O_1894,N_20433,N_22661);
and UO_1895 (O_1895,N_22630,N_20655);
nor UO_1896 (O_1896,N_24266,N_23889);
and UO_1897 (O_1897,N_20400,N_22157);
and UO_1898 (O_1898,N_23299,N_20014);
or UO_1899 (O_1899,N_22675,N_23683);
and UO_1900 (O_1900,N_22941,N_24450);
xnor UO_1901 (O_1901,N_22127,N_21495);
and UO_1902 (O_1902,N_22929,N_20810);
and UO_1903 (O_1903,N_24812,N_20462);
nor UO_1904 (O_1904,N_21502,N_21156);
and UO_1905 (O_1905,N_21271,N_24280);
nand UO_1906 (O_1906,N_24420,N_24802);
or UO_1907 (O_1907,N_20725,N_23432);
and UO_1908 (O_1908,N_22055,N_20325);
or UO_1909 (O_1909,N_22656,N_20333);
nand UO_1910 (O_1910,N_22779,N_20279);
and UO_1911 (O_1911,N_22518,N_22104);
and UO_1912 (O_1912,N_23662,N_24685);
nand UO_1913 (O_1913,N_21650,N_24179);
nor UO_1914 (O_1914,N_23028,N_21155);
and UO_1915 (O_1915,N_21202,N_20244);
and UO_1916 (O_1916,N_24336,N_21599);
nand UO_1917 (O_1917,N_22620,N_20206);
nor UO_1918 (O_1918,N_22771,N_22805);
nor UO_1919 (O_1919,N_24582,N_21219);
nor UO_1920 (O_1920,N_22963,N_23857);
nor UO_1921 (O_1921,N_23925,N_24925);
xnor UO_1922 (O_1922,N_20698,N_24980);
and UO_1923 (O_1923,N_22756,N_23066);
or UO_1924 (O_1924,N_20555,N_22737);
nand UO_1925 (O_1925,N_22529,N_20562);
xnor UO_1926 (O_1926,N_22252,N_22967);
and UO_1927 (O_1927,N_22033,N_22982);
nor UO_1928 (O_1928,N_20013,N_20230);
nor UO_1929 (O_1929,N_24485,N_20362);
nand UO_1930 (O_1930,N_23007,N_23629);
nor UO_1931 (O_1931,N_23221,N_22857);
nor UO_1932 (O_1932,N_24966,N_24230);
nor UO_1933 (O_1933,N_24171,N_21634);
nor UO_1934 (O_1934,N_22757,N_20486);
nand UO_1935 (O_1935,N_24036,N_24617);
and UO_1936 (O_1936,N_24129,N_21264);
or UO_1937 (O_1937,N_24827,N_22408);
xnor UO_1938 (O_1938,N_21279,N_21914);
nor UO_1939 (O_1939,N_23989,N_20589);
nor UO_1940 (O_1940,N_21778,N_21819);
and UO_1941 (O_1941,N_24865,N_20818);
nand UO_1942 (O_1942,N_21242,N_22722);
nand UO_1943 (O_1943,N_22424,N_22765);
xor UO_1944 (O_1944,N_23772,N_24478);
nand UO_1945 (O_1945,N_21265,N_20828);
nor UO_1946 (O_1946,N_22650,N_23962);
nand UO_1947 (O_1947,N_20708,N_23293);
or UO_1948 (O_1948,N_20742,N_21059);
or UO_1949 (O_1949,N_23313,N_24030);
and UO_1950 (O_1950,N_24588,N_24579);
nand UO_1951 (O_1951,N_22090,N_22056);
or UO_1952 (O_1952,N_21733,N_20884);
nor UO_1953 (O_1953,N_20182,N_22807);
nand UO_1954 (O_1954,N_23621,N_21283);
nor UO_1955 (O_1955,N_20980,N_22150);
and UO_1956 (O_1956,N_20454,N_20943);
or UO_1957 (O_1957,N_21534,N_24312);
nand UO_1958 (O_1958,N_20712,N_23560);
xnor UO_1959 (O_1959,N_21176,N_24328);
nor UO_1960 (O_1960,N_22027,N_24194);
and UO_1961 (O_1961,N_21884,N_24357);
or UO_1962 (O_1962,N_22628,N_22883);
or UO_1963 (O_1963,N_22734,N_24905);
nor UO_1964 (O_1964,N_23670,N_21461);
nor UO_1965 (O_1965,N_22152,N_21755);
and UO_1966 (O_1966,N_22066,N_24566);
xnor UO_1967 (O_1967,N_21042,N_23768);
or UO_1968 (O_1968,N_21478,N_22750);
xor UO_1969 (O_1969,N_21096,N_22324);
or UO_1970 (O_1970,N_20586,N_22392);
and UO_1971 (O_1971,N_23368,N_21262);
and UO_1972 (O_1972,N_20465,N_21829);
nor UO_1973 (O_1973,N_22752,N_23797);
nand UO_1974 (O_1974,N_21406,N_23410);
nand UO_1975 (O_1975,N_21269,N_22698);
nand UO_1976 (O_1976,N_20656,N_23262);
or UO_1977 (O_1977,N_23086,N_24661);
and UO_1978 (O_1978,N_23004,N_23487);
and UO_1979 (O_1979,N_23698,N_23079);
and UO_1980 (O_1980,N_21810,N_23140);
and UO_1981 (O_1981,N_22950,N_24377);
or UO_1982 (O_1982,N_20200,N_20851);
nor UO_1983 (O_1983,N_23813,N_20716);
or UO_1984 (O_1984,N_24111,N_21290);
or UO_1985 (O_1985,N_20162,N_23220);
and UO_1986 (O_1986,N_24221,N_20039);
nor UO_1987 (O_1987,N_23911,N_20157);
and UO_1988 (O_1988,N_20071,N_21643);
xor UO_1989 (O_1989,N_24818,N_20338);
nor UO_1990 (O_1990,N_21972,N_20870);
xor UO_1991 (O_1991,N_23366,N_24795);
nor UO_1992 (O_1992,N_24896,N_20156);
and UO_1993 (O_1993,N_22469,N_24732);
or UO_1994 (O_1994,N_21784,N_22671);
and UO_1995 (O_1995,N_23743,N_22024);
nand UO_1996 (O_1996,N_21681,N_20621);
nand UO_1997 (O_1997,N_24251,N_23218);
nor UO_1998 (O_1998,N_20643,N_21010);
and UO_1999 (O_1999,N_23806,N_21941);
and UO_2000 (O_2000,N_23069,N_21764);
and UO_2001 (O_2001,N_22995,N_24436);
and UO_2002 (O_2002,N_20754,N_20294);
or UO_2003 (O_2003,N_23655,N_22938);
or UO_2004 (O_2004,N_20910,N_20188);
nand UO_2005 (O_2005,N_23107,N_24237);
xnor UO_2006 (O_2006,N_22923,N_20744);
or UO_2007 (O_2007,N_23720,N_20937);
or UO_2008 (O_2008,N_22704,N_24964);
or UO_2009 (O_2009,N_22812,N_23778);
nand UO_2010 (O_2010,N_22226,N_23596);
or UO_2011 (O_2011,N_21638,N_21551);
and UO_2012 (O_2012,N_24855,N_21772);
xor UO_2013 (O_2013,N_22587,N_24174);
or UO_2014 (O_2014,N_24672,N_20405);
nand UO_2015 (O_2015,N_24212,N_23603);
nand UO_2016 (O_2016,N_20317,N_22230);
xnor UO_2017 (O_2017,N_20363,N_20429);
and UO_2018 (O_2018,N_20648,N_20842);
nor UO_2019 (O_2019,N_23172,N_21707);
xor UO_2020 (O_2020,N_24167,N_21451);
nor UO_2021 (O_2021,N_23759,N_20151);
and UO_2022 (O_2022,N_20098,N_21635);
xnor UO_2023 (O_2023,N_22266,N_24120);
and UO_2024 (O_2024,N_20128,N_24223);
and UO_2025 (O_2025,N_21636,N_20089);
and UO_2026 (O_2026,N_21877,N_20569);
or UO_2027 (O_2027,N_24850,N_23047);
or UO_2028 (O_2028,N_24287,N_21258);
nand UO_2029 (O_2029,N_21192,N_23888);
nand UO_2030 (O_2030,N_23422,N_22464);
xnor UO_2031 (O_2031,N_20050,N_23174);
nor UO_2032 (O_2032,N_23590,N_24161);
xnor UO_2033 (O_2033,N_22466,N_24900);
nor UO_2034 (O_2034,N_20874,N_24948);
or UO_2035 (O_2035,N_21578,N_23332);
nand UO_2036 (O_2036,N_22126,N_21835);
nor UO_2037 (O_2037,N_24027,N_23063);
and UO_2038 (O_2038,N_20418,N_23750);
or UO_2039 (O_2039,N_21212,N_24576);
nor UO_2040 (O_2040,N_22899,N_24491);
or UO_2041 (O_2041,N_22057,N_23951);
and UO_2042 (O_2042,N_21974,N_21646);
nand UO_2043 (O_2043,N_21748,N_20023);
nand UO_2044 (O_2044,N_24941,N_20148);
nand UO_2045 (O_2045,N_20671,N_24619);
or UO_2046 (O_2046,N_23552,N_22829);
xor UO_2047 (O_2047,N_23909,N_24768);
nor UO_2048 (O_2048,N_24308,N_20999);
and UO_2049 (O_2049,N_20471,N_22654);
or UO_2050 (O_2050,N_21029,N_22643);
nor UO_2051 (O_2051,N_24360,N_24556);
nand UO_2052 (O_2052,N_21807,N_24874);
nor UO_2053 (O_2053,N_21177,N_20402);
and UO_2054 (O_2054,N_20531,N_21538);
or UO_2055 (O_2055,N_23415,N_21325);
or UO_2056 (O_2056,N_23676,N_22071);
nor UO_2057 (O_2057,N_22960,N_21228);
nor UO_2058 (O_2058,N_24327,N_22749);
and UO_2059 (O_2059,N_24698,N_22694);
or UO_2060 (O_2060,N_23756,N_24749);
or UO_2061 (O_2061,N_20203,N_24889);
and UO_2062 (O_2062,N_21340,N_23940);
and UO_2063 (O_2063,N_21018,N_22495);
and UO_2064 (O_2064,N_20307,N_21828);
nand UO_2065 (O_2065,N_20055,N_22341);
and UO_2066 (O_2066,N_23915,N_20597);
nand UO_2067 (O_2067,N_20604,N_21609);
xor UO_2068 (O_2068,N_20674,N_22998);
nand UO_2069 (O_2069,N_23832,N_22895);
or UO_2070 (O_2070,N_21487,N_24370);
nor UO_2071 (O_2071,N_23298,N_22278);
xnor UO_2072 (O_2072,N_24099,N_20706);
nor UO_2073 (O_2073,N_22353,N_23228);
xor UO_2074 (O_2074,N_22263,N_20295);
nand UO_2075 (O_2075,N_24658,N_22567);
xor UO_2076 (O_2076,N_23120,N_20146);
nand UO_2077 (O_2077,N_20102,N_24024);
or UO_2078 (O_2078,N_23489,N_23505);
and UO_2079 (O_2079,N_24723,N_21060);
and UO_2080 (O_2080,N_22819,N_22279);
nor UO_2081 (O_2081,N_20672,N_20253);
nand UO_2082 (O_2082,N_22808,N_22208);
or UO_2083 (O_2083,N_21428,N_20056);
or UO_2084 (O_2084,N_21967,N_24643);
nor UO_2085 (O_2085,N_21500,N_22191);
and UO_2086 (O_2086,N_22036,N_22893);
and UO_2087 (O_2087,N_21492,N_23074);
nand UO_2088 (O_2088,N_20349,N_20177);
nor UO_2089 (O_2089,N_22997,N_24895);
nand UO_2090 (O_2090,N_24256,N_22361);
nand UO_2091 (O_2091,N_22623,N_21146);
nand UO_2092 (O_2092,N_23342,N_24480);
or UO_2093 (O_2093,N_22777,N_20473);
nand UO_2094 (O_2094,N_23344,N_23239);
or UO_2095 (O_2095,N_24003,N_20065);
and UO_2096 (O_2096,N_23314,N_23625);
and UO_2097 (O_2097,N_24787,N_23972);
nor UO_2098 (O_2098,N_22692,N_20118);
nor UO_2099 (O_2099,N_20573,N_22527);
nor UO_2100 (O_2100,N_23606,N_21251);
and UO_2101 (O_2101,N_24315,N_20180);
nor UO_2102 (O_2102,N_20179,N_23882);
nand UO_2103 (O_2103,N_23773,N_23373);
nand UO_2104 (O_2104,N_21834,N_20781);
nand UO_2105 (O_2105,N_21921,N_23354);
nand UO_2106 (O_2106,N_20368,N_20670);
nand UO_2107 (O_2107,N_21543,N_21623);
nor UO_2108 (O_2108,N_24011,N_20477);
and UO_2109 (O_2109,N_20691,N_24722);
nand UO_2110 (O_2110,N_20778,N_21011);
and UO_2111 (O_2111,N_21735,N_20296);
nand UO_2112 (O_2112,N_23491,N_23090);
nand UO_2113 (O_2113,N_23929,N_21441);
nand UO_2114 (O_2114,N_23518,N_22331);
and UO_2115 (O_2115,N_24656,N_21329);
nor UO_2116 (O_2116,N_22762,N_21463);
and UO_2117 (O_2117,N_24009,N_24877);
nor UO_2118 (O_2118,N_23138,N_23419);
and UO_2119 (O_2119,N_20076,N_21306);
xnor UO_2120 (O_2120,N_21468,N_20886);
nand UO_2121 (O_2121,N_20600,N_22032);
nor UO_2122 (O_2122,N_22815,N_23957);
or UO_2123 (O_2123,N_23907,N_21473);
nand UO_2124 (O_2124,N_24632,N_22889);
nand UO_2125 (O_2125,N_22428,N_24940);
or UO_2126 (O_2126,N_21811,N_23767);
nor UO_2127 (O_2127,N_24286,N_22562);
nand UO_2128 (O_2128,N_24552,N_21027);
or UO_2129 (O_2129,N_21501,N_20257);
nand UO_2130 (O_2130,N_23263,N_23269);
and UO_2131 (O_2131,N_22548,N_21853);
nand UO_2132 (O_2132,N_24040,N_23645);
and UO_2133 (O_2133,N_24952,N_23073);
and UO_2134 (O_2134,N_21798,N_21814);
and UO_2135 (O_2135,N_23339,N_23242);
nand UO_2136 (O_2136,N_23731,N_22571);
nand UO_2137 (O_2137,N_24102,N_21223);
or UO_2138 (O_2138,N_20899,N_22953);
and UO_2139 (O_2139,N_23029,N_22435);
or UO_2140 (O_2140,N_24209,N_24708);
or UO_2141 (O_2141,N_21611,N_22785);
or UO_2142 (O_2142,N_23297,N_21217);
xnor UO_2143 (O_2143,N_22186,N_22978);
nand UO_2144 (O_2144,N_23192,N_22547);
xnor UO_2145 (O_2145,N_21377,N_23825);
nand UO_2146 (O_2146,N_22732,N_20721);
nor UO_2147 (O_2147,N_21903,N_23609);
nand UO_2148 (O_2148,N_21792,N_20373);
and UO_2149 (O_2149,N_20814,N_24534);
xnor UO_2150 (O_2150,N_20892,N_21307);
and UO_2151 (O_2151,N_21229,N_21158);
nor UO_2152 (O_2152,N_21250,N_23216);
and UO_2153 (O_2153,N_20813,N_21056);
or UO_2154 (O_2154,N_24400,N_21354);
and UO_2155 (O_2155,N_23434,N_22449);
nand UO_2156 (O_2156,N_24028,N_23026);
xnor UO_2157 (O_2157,N_20004,N_24114);
or UO_2158 (O_2158,N_23421,N_21827);
and UO_2159 (O_2159,N_24159,N_23588);
or UO_2160 (O_2160,N_20115,N_22775);
nand UO_2161 (O_2161,N_20853,N_20694);
and UO_2162 (O_2162,N_22015,N_20348);
or UO_2163 (O_2163,N_24385,N_24747);
and UO_2164 (O_2164,N_24642,N_21568);
and UO_2165 (O_2165,N_23551,N_20976);
or UO_2166 (O_2166,N_22006,N_24067);
or UO_2167 (O_2167,N_20249,N_24801);
or UO_2168 (O_2168,N_20339,N_20340);
and UO_2169 (O_2169,N_24185,N_23163);
nor UO_2170 (O_2170,N_20939,N_23634);
nand UO_2171 (O_2171,N_21546,N_24046);
and UO_2172 (O_2172,N_22440,N_21905);
nor UO_2173 (O_2173,N_24906,N_24386);
or UO_2174 (O_2174,N_22391,N_23251);
and UO_2175 (O_2175,N_24584,N_24408);
xnor UO_2176 (O_2176,N_21700,N_22307);
or UO_2177 (O_2177,N_24770,N_23370);
or UO_2178 (O_2178,N_20003,N_20558);
nand UO_2179 (O_2179,N_20306,N_20916);
xor UO_2180 (O_2180,N_20964,N_23875);
xnor UO_2181 (O_2181,N_24994,N_20336);
nand UO_2182 (O_2182,N_24599,N_21054);
and UO_2183 (O_2183,N_24081,N_22538);
nor UO_2184 (O_2184,N_24041,N_23132);
nor UO_2185 (O_2185,N_22666,N_24101);
nor UO_2186 (O_2186,N_20326,N_22736);
nor UO_2187 (O_2187,N_20367,N_22436);
nand UO_2188 (O_2188,N_24008,N_22423);
or UO_2189 (O_2189,N_20908,N_23514);
nand UO_2190 (O_2190,N_23424,N_23418);
or UO_2191 (O_2191,N_23969,N_20822);
and UO_2192 (O_2192,N_22639,N_24957);
and UO_2193 (O_2193,N_23384,N_23544);
nor UO_2194 (O_2194,N_24771,N_23573);
xor UO_2195 (O_2195,N_20762,N_24744);
nand UO_2196 (O_2196,N_21677,N_20080);
and UO_2197 (O_2197,N_24783,N_21709);
nand UO_2198 (O_2198,N_20176,N_23176);
nand UO_2199 (O_2199,N_24741,N_21273);
xor UO_2200 (O_2200,N_20396,N_23340);
nor UO_2201 (O_2201,N_24441,N_23393);
nand UO_2202 (O_2202,N_21070,N_22383);
nor UO_2203 (O_2203,N_21637,N_23499);
xnor UO_2204 (O_2204,N_22430,N_24953);
xnor UO_2205 (O_2205,N_24288,N_20848);
nor UO_2206 (O_2206,N_24307,N_22289);
nor UO_2207 (O_2207,N_21388,N_23451);
nand UO_2208 (O_2208,N_23044,N_24633);
nand UO_2209 (O_2209,N_23353,N_22672);
nor UO_2210 (O_2210,N_20995,N_23329);
or UO_2211 (O_2211,N_22702,N_22787);
nor UO_2212 (O_2212,N_20228,N_24659);
or UO_2213 (O_2213,N_23980,N_21769);
nand UO_2214 (O_2214,N_22725,N_22870);
or UO_2215 (O_2215,N_21136,N_24929);
xnor UO_2216 (O_2216,N_23287,N_20347);
nor UO_2217 (O_2217,N_21132,N_21165);
and UO_2218 (O_2218,N_23717,N_20374);
or UO_2219 (O_2219,N_24826,N_24762);
and UO_2220 (O_2220,N_21916,N_21380);
or UO_2221 (O_2221,N_22511,N_20308);
or UO_2222 (O_2222,N_24115,N_22772);
xnor UO_2223 (O_2223,N_21816,N_24782);
xnor UO_2224 (O_2224,N_24356,N_22659);
nand UO_2225 (O_2225,N_23826,N_23738);
and UO_2226 (O_2226,N_20298,N_20794);
or UO_2227 (O_2227,N_23788,N_23960);
nand UO_2228 (O_2228,N_22219,N_22909);
nand UO_2229 (O_2229,N_23274,N_20434);
nand UO_2230 (O_2230,N_23934,N_20962);
nand UO_2231 (O_2231,N_23011,N_22211);
or UO_2232 (O_2232,N_20215,N_20164);
or UO_2233 (O_2233,N_20626,N_24607);
and UO_2234 (O_2234,N_20037,N_22689);
or UO_2235 (O_2235,N_24216,N_20331);
and UO_2236 (O_2236,N_23715,N_24690);
or UO_2237 (O_2237,N_20987,N_23039);
or UO_2238 (O_2238,N_21147,N_23350);
and UO_2239 (O_2239,N_21922,N_24058);
or UO_2240 (O_2240,N_22871,N_20258);
nand UO_2241 (O_2241,N_22516,N_21936);
and UO_2242 (O_2242,N_20346,N_22691);
nor UO_2243 (O_2243,N_24564,N_21133);
or UO_2244 (O_2244,N_20686,N_24127);
nand UO_2245 (O_2245,N_24084,N_22513);
or UO_2246 (O_2246,N_22132,N_22337);
or UO_2247 (O_2247,N_22119,N_22432);
nand UO_2248 (O_2248,N_24200,N_23018);
nor UO_2249 (O_2249,N_22310,N_24123);
nor UO_2250 (O_2250,N_23116,N_21321);
and UO_2251 (O_2251,N_21211,N_21506);
or UO_2252 (O_2252,N_24620,N_22727);
and UO_2253 (O_2253,N_24734,N_22395);
nand UO_2254 (O_2254,N_20412,N_21688);
xor UO_2255 (O_2255,N_21680,N_22507);
nand UO_2256 (O_2256,N_21625,N_22101);
or UO_2257 (O_2257,N_23167,N_21817);
nor UO_2258 (O_2258,N_21466,N_24378);
nor UO_2259 (O_2259,N_22993,N_24100);
nor UO_2260 (O_2260,N_20681,N_21621);
nor UO_2261 (O_2261,N_22901,N_20352);
and UO_2262 (O_2262,N_20404,N_24604);
nor UO_2263 (O_2263,N_20890,N_22552);
nor UO_2264 (O_2264,N_22384,N_23894);
or UO_2265 (O_2265,N_21446,N_21954);
and UO_2266 (O_2266,N_22836,N_23295);
nand UO_2267 (O_2267,N_22665,N_22251);
nand UO_2268 (O_2268,N_20865,N_20803);
and UO_2269 (O_2269,N_24680,N_20035);
or UO_2270 (O_2270,N_22345,N_23930);
xor UO_2271 (O_2271,N_24334,N_24547);
nor UO_2272 (O_2272,N_21225,N_23669);
nand UO_2273 (O_2273,N_23963,N_22690);
nor UO_2274 (O_2274,N_20447,N_22273);
nand UO_2275 (O_2275,N_24188,N_23358);
nor UO_2276 (O_2276,N_22426,N_22268);
nand UO_2277 (O_2277,N_21642,N_20914);
xnor UO_2278 (O_2278,N_24920,N_21448);
and UO_2279 (O_2279,N_24916,N_22089);
nand UO_2280 (O_2280,N_22167,N_24624);
and UO_2281 (O_2281,N_23002,N_21875);
or UO_2282 (O_2282,N_22831,N_21483);
nand UO_2283 (O_2283,N_23880,N_22743);
and UO_2284 (O_2284,N_21869,N_22634);
nor UO_2285 (O_2285,N_22461,N_21287);
or UO_2286 (O_2286,N_23936,N_23516);
and UO_2287 (O_2287,N_20852,N_23471);
nor UO_2288 (O_2288,N_22097,N_21179);
or UO_2289 (O_2289,N_24432,N_23713);
nor UO_2290 (O_2290,N_24068,N_22877);
or UO_2291 (O_2291,N_24977,N_22429);
nand UO_2292 (O_2292,N_24264,N_21741);
nor UO_2293 (O_2293,N_21455,N_22544);
nand UO_2294 (O_2294,N_21907,N_22565);
and UO_2295 (O_2295,N_20082,N_21773);
xnor UO_2296 (O_2296,N_24808,N_24861);
or UO_2297 (O_2297,N_23841,N_23707);
xor UO_2298 (O_2298,N_21151,N_20239);
nor UO_2299 (O_2299,N_21782,N_24713);
nor UO_2300 (O_2300,N_20512,N_20354);
and UO_2301 (O_2301,N_21859,N_23395);
nand UO_2302 (O_2302,N_21964,N_24414);
nor UO_2303 (O_2303,N_22825,N_22417);
or UO_2304 (O_2304,N_20123,N_24881);
nor UO_2305 (O_2305,N_23521,N_24311);
or UO_2306 (O_2306,N_21886,N_23824);
or UO_2307 (O_2307,N_21836,N_20925);
nor UO_2308 (O_2308,N_23595,N_21508);
or UO_2309 (O_2309,N_24451,N_21407);
nand UO_2310 (O_2310,N_24424,N_20189);
and UO_2311 (O_2311,N_20463,N_20481);
or UO_2312 (O_2312,N_24206,N_23374);
nand UO_2313 (O_2313,N_21879,N_20361);
or UO_2314 (O_2314,N_21788,N_23714);
nand UO_2315 (O_2315,N_23141,N_21654);
and UO_2316 (O_2316,N_23465,N_21494);
nand UO_2317 (O_2317,N_21514,N_24234);
and UO_2318 (O_2318,N_24372,N_22854);
nand UO_2319 (O_2319,N_22158,N_24396);
nor UO_2320 (O_2320,N_22137,N_24032);
or UO_2321 (O_2321,N_21138,N_23012);
nor UO_2322 (O_2322,N_22638,N_23319);
and UO_2323 (O_2323,N_24592,N_21216);
nor UO_2324 (O_2324,N_23893,N_20423);
and UO_2325 (O_2325,N_22835,N_22120);
nor UO_2326 (O_2326,N_20788,N_23131);
nand UO_2327 (O_2327,N_21708,N_20894);
or UO_2328 (O_2328,N_24772,N_21427);
and UO_2329 (O_2329,N_20456,N_20017);
or UO_2330 (O_2330,N_23158,N_20417);
nand UO_2331 (O_2331,N_23392,N_23322);
and UO_2332 (O_2332,N_24326,N_23668);
nor UO_2333 (O_2333,N_22506,N_21358);
nor UO_2334 (O_2334,N_20519,N_23005);
nand UO_2335 (O_2335,N_23681,N_22026);
nand UO_2336 (O_2336,N_24909,N_22037);
nor UO_2337 (O_2337,N_24150,N_22549);
nor UO_2338 (O_2338,N_22295,N_24176);
or UO_2339 (O_2339,N_23021,N_22577);
or UO_2340 (O_2340,N_22826,N_22497);
and UO_2341 (O_2341,N_21272,N_20860);
or UO_2342 (O_2342,N_24794,N_22514);
and UO_2343 (O_2343,N_20734,N_20323);
nand UO_2344 (O_2344,N_22124,N_20277);
or UO_2345 (O_2345,N_24899,N_21185);
or UO_2346 (O_2346,N_22632,N_21555);
xnor UO_2347 (O_2347,N_20841,N_21195);
nor UO_2348 (O_2348,N_24750,N_22014);
and UO_2349 (O_2349,N_20439,N_22003);
and UO_2350 (O_2350,N_23584,N_22832);
and UO_2351 (O_2351,N_24731,N_21409);
xnor UO_2352 (O_2352,N_24358,N_23819);
and UO_2353 (O_2353,N_20743,N_21776);
nor UO_2354 (O_2354,N_24109,N_21787);
and UO_2355 (O_2355,N_20407,N_23500);
and UO_2356 (O_2356,N_20850,N_24300);
xor UO_2357 (O_2357,N_22332,N_21565);
and UO_2358 (O_2358,N_24822,N_21600);
and UO_2359 (O_2359,N_23127,N_23450);
or UO_2360 (O_2360,N_22542,N_21245);
and UO_2361 (O_2361,N_20383,N_22048);
nand UO_2362 (O_2362,N_24836,N_21801);
nor UO_2363 (O_2363,N_23134,N_24324);
xnor UO_2364 (O_2364,N_24322,N_22977);
nand UO_2365 (O_2365,N_20587,N_22616);
or UO_2366 (O_2366,N_20092,N_24361);
and UO_2367 (O_2367,N_24796,N_20912);
or UO_2368 (O_2368,N_20199,N_23591);
nor UO_2369 (O_2369,N_20048,N_20191);
nand UO_2370 (O_2370,N_24395,N_20500);
nor UO_2371 (O_2371,N_21003,N_23704);
xnor UO_2372 (O_2372,N_23495,N_24669);
nand UO_2373 (O_2373,N_23648,N_23869);
or UO_2374 (O_2374,N_24951,N_22768);
and UO_2375 (O_2375,N_20068,N_22664);
and UO_2376 (O_2376,N_23180,N_24153);
xor UO_2377 (O_2377,N_21725,N_24725);
or UO_2378 (O_2378,N_24694,N_24548);
nor UO_2379 (O_2379,N_22260,N_23531);
nand UO_2380 (O_2380,N_21384,N_23995);
nor UO_2381 (O_2381,N_21498,N_23845);
nor UO_2382 (O_2382,N_22141,N_23539);
or UO_2383 (O_2383,N_22521,N_22344);
nand UO_2384 (O_2384,N_22482,N_21575);
xor UO_2385 (O_2385,N_20321,N_24453);
and UO_2386 (O_2386,N_20498,N_20782);
nor UO_2387 (O_2387,N_23747,N_24857);
or UO_2388 (O_2388,N_24924,N_24972);
xnor UO_2389 (O_2389,N_20350,N_21771);
or UO_2390 (O_2390,N_20954,N_22486);
nor UO_2391 (O_2391,N_22784,N_20281);
and UO_2392 (O_2392,N_22684,N_23053);
nor UO_2393 (O_2393,N_22302,N_23578);
or UO_2394 (O_2394,N_24901,N_24561);
nand UO_2395 (O_2395,N_24973,N_24301);
and UO_2396 (O_2396,N_20972,N_20680);
and UO_2397 (O_2397,N_24655,N_22489);
nand UO_2398 (O_2398,N_23691,N_24716);
and UO_2399 (O_2399,N_24843,N_21505);
and UO_2400 (O_2400,N_23436,N_22509);
and UO_2401 (O_2401,N_24279,N_23604);
xor UO_2402 (O_2402,N_24224,N_21606);
and UO_2403 (O_2403,N_23289,N_22796);
nor UO_2404 (O_2404,N_23900,N_23847);
xnor UO_2405 (O_2405,N_22512,N_23347);
nand UO_2406 (O_2406,N_23110,N_23452);
nand UO_2407 (O_2407,N_24012,N_23222);
nor UO_2408 (O_2408,N_22274,N_23716);
or UO_2409 (O_2409,N_24371,N_21602);
or UO_2410 (O_2410,N_22789,N_23094);
nor UO_2411 (O_2411,N_22112,N_24169);
or UO_2412 (O_2412,N_23307,N_20904);
nor UO_2413 (O_2413,N_20328,N_24662);
nand UO_2414 (O_2414,N_22590,N_21897);
nor UO_2415 (O_2415,N_23253,N_22708);
and UO_2416 (O_2416,N_22109,N_24181);
and UO_2417 (O_2417,N_24815,N_21234);
xor UO_2418 (O_2418,N_21765,N_20124);
nor UO_2419 (O_2419,N_20271,N_20990);
or UO_2420 (O_2420,N_24955,N_21504);
or UO_2421 (O_2421,N_22309,N_20798);
and UO_2422 (O_2422,N_22714,N_20173);
nor UO_2423 (O_2423,N_21232,N_20844);
and UO_2424 (O_2424,N_22631,N_23955);
nand UO_2425 (O_2425,N_20171,N_24594);
nor UO_2426 (O_2426,N_20545,N_21139);
nand UO_2427 (O_2427,N_20799,N_20871);
nor UO_2428 (O_2428,N_20466,N_21361);
nand UO_2429 (O_2429,N_21385,N_21577);
and UO_2430 (O_2430,N_22350,N_21533);
or UO_2431 (O_2431,N_24254,N_21594);
xor UO_2432 (O_2432,N_23335,N_21540);
nor UO_2433 (O_2433,N_24348,N_20120);
nor UO_2434 (O_2434,N_23809,N_21892);
and UO_2435 (O_2435,N_24758,N_23477);
or UO_2436 (O_2436,N_20632,N_23193);
nand UO_2437 (O_2437,N_23054,N_21656);
and UO_2438 (O_2438,N_20543,N_23096);
or UO_2439 (O_2439,N_24292,N_22801);
nand UO_2440 (O_2440,N_24748,N_20785);
or UO_2441 (O_2441,N_23416,N_21280);
and UO_2442 (O_2442,N_23331,N_24434);
nor UO_2443 (O_2443,N_22876,N_24457);
nand UO_2444 (O_2444,N_21998,N_23369);
nor UO_2445 (O_2445,N_24517,N_20898);
nand UO_2446 (O_2446,N_22578,N_24018);
or UO_2447 (O_2447,N_24965,N_23812);
nand UO_2448 (O_2448,N_23579,N_24928);
or UO_2449 (O_2449,N_21815,N_23895);
xnor UO_2450 (O_2450,N_20709,N_21248);
nor UO_2451 (O_2451,N_21119,N_21410);
xor UO_2452 (O_2452,N_20710,N_21405);
nand UO_2453 (O_2453,N_23855,N_24486);
nand UO_2454 (O_2454,N_24148,N_22696);
or UO_2455 (O_2455,N_20435,N_22687);
nor UO_2456 (O_2456,N_22981,N_21515);
and UO_2457 (O_2457,N_24401,N_23362);
nor UO_2458 (O_2458,N_23978,N_21779);
nor UO_2459 (O_2459,N_21949,N_20553);
xnor UO_2460 (O_2460,N_23440,N_21116);
nand UO_2461 (O_2461,N_20469,N_21047);
nor UO_2462 (O_2462,N_23870,N_22454);
and UO_2463 (O_2463,N_21348,N_24792);
or UO_2464 (O_2464,N_22296,N_20765);
and UO_2465 (O_2465,N_22746,N_22358);
nand UO_2466 (O_2466,N_23136,N_21544);
nand UO_2467 (O_2467,N_22442,N_22298);
and UO_2468 (O_2468,N_20556,N_20442);
nor UO_2469 (O_2469,N_23064,N_24756);
and UO_2470 (O_2470,N_20459,N_23932);
or UO_2471 (O_2471,N_22257,N_22184);
nor UO_2472 (O_2472,N_22166,N_22276);
or UO_2473 (O_2473,N_21206,N_20138);
and UO_2474 (O_2474,N_22573,N_22183);
and UO_2475 (O_2475,N_20223,N_23583);
and UO_2476 (O_2476,N_21662,N_24416);
and UO_2477 (O_2477,N_22325,N_21517);
nor UO_2478 (O_2478,N_24069,N_24779);
nand UO_2479 (O_2479,N_24156,N_24847);
or UO_2480 (O_2480,N_21692,N_24210);
and UO_2481 (O_2481,N_20501,N_24760);
and UO_2482 (O_2482,N_23190,N_24172);
or UO_2483 (O_2483,N_23526,N_22657);
or UO_2484 (O_2484,N_20869,N_24320);
and UO_2485 (O_2485,N_21443,N_23587);
xor UO_2486 (O_2486,N_22088,N_21355);
or UO_2487 (O_2487,N_24504,N_24253);
nand UO_2488 (O_2488,N_23822,N_23202);
or UO_2489 (O_2489,N_23092,N_21790);
and UO_2490 (O_2490,N_24567,N_22163);
and UO_2491 (O_2491,N_22161,N_24512);
nor UO_2492 (O_2492,N_23548,N_23550);
nor UO_2493 (O_2493,N_21083,N_21520);
and UO_2494 (O_2494,N_20359,N_20327);
or UO_2495 (O_2495,N_20700,N_24858);
and UO_2496 (O_2496,N_21858,N_24737);
or UO_2497 (O_2497,N_22214,N_21719);
xor UO_2498 (O_2498,N_23055,N_21286);
and UO_2499 (O_2499,N_21826,N_20195);
nor UO_2500 (O_2500,N_20996,N_22186);
and UO_2501 (O_2501,N_22475,N_22875);
or UO_2502 (O_2502,N_23686,N_24088);
nor UO_2503 (O_2503,N_22354,N_22562);
and UO_2504 (O_2504,N_24252,N_21598);
and UO_2505 (O_2505,N_22276,N_24008);
or UO_2506 (O_2506,N_24867,N_21252);
nand UO_2507 (O_2507,N_20141,N_23831);
and UO_2508 (O_2508,N_20738,N_21467);
or UO_2509 (O_2509,N_24138,N_22518);
or UO_2510 (O_2510,N_24890,N_22710);
nand UO_2511 (O_2511,N_20403,N_22738);
xor UO_2512 (O_2512,N_22203,N_21002);
nand UO_2513 (O_2513,N_20156,N_20608);
and UO_2514 (O_2514,N_22649,N_23660);
or UO_2515 (O_2515,N_20973,N_22659);
and UO_2516 (O_2516,N_23603,N_23057);
nand UO_2517 (O_2517,N_22566,N_20509);
and UO_2518 (O_2518,N_23522,N_23494);
xnor UO_2519 (O_2519,N_21813,N_24021);
xor UO_2520 (O_2520,N_22386,N_21701);
or UO_2521 (O_2521,N_22341,N_21081);
or UO_2522 (O_2522,N_24747,N_20855);
nor UO_2523 (O_2523,N_22422,N_20711);
xnor UO_2524 (O_2524,N_21789,N_20152);
or UO_2525 (O_2525,N_22991,N_21244);
or UO_2526 (O_2526,N_23992,N_20224);
or UO_2527 (O_2527,N_23525,N_21866);
or UO_2528 (O_2528,N_23645,N_22943);
nand UO_2529 (O_2529,N_20190,N_20611);
or UO_2530 (O_2530,N_22312,N_20483);
or UO_2531 (O_2531,N_22098,N_23137);
or UO_2532 (O_2532,N_20380,N_20460);
xnor UO_2533 (O_2533,N_24298,N_24854);
and UO_2534 (O_2534,N_23355,N_22917);
or UO_2535 (O_2535,N_22058,N_23707);
and UO_2536 (O_2536,N_24908,N_20500);
nand UO_2537 (O_2537,N_20230,N_23144);
nor UO_2538 (O_2538,N_22244,N_21275);
or UO_2539 (O_2539,N_21242,N_22827);
xnor UO_2540 (O_2540,N_23351,N_20924);
nor UO_2541 (O_2541,N_22755,N_22722);
nor UO_2542 (O_2542,N_23647,N_21896);
nand UO_2543 (O_2543,N_24708,N_24156);
or UO_2544 (O_2544,N_22456,N_24861);
nor UO_2545 (O_2545,N_24119,N_21914);
nor UO_2546 (O_2546,N_21384,N_24328);
nand UO_2547 (O_2547,N_21007,N_22589);
xnor UO_2548 (O_2548,N_23995,N_24486);
nand UO_2549 (O_2549,N_20387,N_24539);
nand UO_2550 (O_2550,N_24979,N_21199);
and UO_2551 (O_2551,N_24337,N_21711);
nand UO_2552 (O_2552,N_22552,N_24152);
nand UO_2553 (O_2553,N_23533,N_23050);
and UO_2554 (O_2554,N_23425,N_22336);
nand UO_2555 (O_2555,N_24131,N_20686);
or UO_2556 (O_2556,N_20386,N_24742);
nor UO_2557 (O_2557,N_23694,N_21739);
or UO_2558 (O_2558,N_22527,N_24416);
and UO_2559 (O_2559,N_23893,N_23138);
nor UO_2560 (O_2560,N_23599,N_20416);
nor UO_2561 (O_2561,N_21961,N_24086);
nor UO_2562 (O_2562,N_22526,N_21367);
and UO_2563 (O_2563,N_21076,N_22582);
nand UO_2564 (O_2564,N_20597,N_22407);
and UO_2565 (O_2565,N_23583,N_21798);
or UO_2566 (O_2566,N_23898,N_23144);
or UO_2567 (O_2567,N_23757,N_24234);
or UO_2568 (O_2568,N_22597,N_20116);
and UO_2569 (O_2569,N_20376,N_22897);
nor UO_2570 (O_2570,N_22420,N_20227);
or UO_2571 (O_2571,N_23126,N_21298);
nor UO_2572 (O_2572,N_21882,N_22531);
or UO_2573 (O_2573,N_24071,N_21633);
nor UO_2574 (O_2574,N_22696,N_22307);
or UO_2575 (O_2575,N_20174,N_20999);
or UO_2576 (O_2576,N_21109,N_22265);
or UO_2577 (O_2577,N_23011,N_24727);
nand UO_2578 (O_2578,N_20604,N_22236);
or UO_2579 (O_2579,N_22931,N_20740);
nand UO_2580 (O_2580,N_20082,N_24688);
nand UO_2581 (O_2581,N_22503,N_20681);
or UO_2582 (O_2582,N_23792,N_22709);
or UO_2583 (O_2583,N_23734,N_20100);
nand UO_2584 (O_2584,N_21047,N_23160);
or UO_2585 (O_2585,N_22859,N_24227);
and UO_2586 (O_2586,N_21117,N_20896);
nand UO_2587 (O_2587,N_24041,N_23500);
nor UO_2588 (O_2588,N_20191,N_20431);
and UO_2589 (O_2589,N_22668,N_22051);
xnor UO_2590 (O_2590,N_24147,N_21902);
nor UO_2591 (O_2591,N_21653,N_22358);
nor UO_2592 (O_2592,N_22988,N_21951);
xnor UO_2593 (O_2593,N_24251,N_24357);
and UO_2594 (O_2594,N_22045,N_21502);
nor UO_2595 (O_2595,N_21350,N_24025);
nor UO_2596 (O_2596,N_21910,N_21192);
or UO_2597 (O_2597,N_20425,N_23478);
nor UO_2598 (O_2598,N_21657,N_23762);
or UO_2599 (O_2599,N_21703,N_22772);
and UO_2600 (O_2600,N_21879,N_22934);
nor UO_2601 (O_2601,N_21536,N_21596);
nand UO_2602 (O_2602,N_20395,N_21007);
and UO_2603 (O_2603,N_20150,N_22576);
xnor UO_2604 (O_2604,N_22152,N_20228);
or UO_2605 (O_2605,N_20644,N_20060);
nor UO_2606 (O_2606,N_23189,N_24666);
or UO_2607 (O_2607,N_20623,N_22767);
or UO_2608 (O_2608,N_20915,N_22443);
and UO_2609 (O_2609,N_24532,N_24298);
and UO_2610 (O_2610,N_23702,N_24318);
nand UO_2611 (O_2611,N_21786,N_21355);
or UO_2612 (O_2612,N_23156,N_23775);
nand UO_2613 (O_2613,N_22834,N_23964);
or UO_2614 (O_2614,N_21473,N_20519);
or UO_2615 (O_2615,N_21372,N_24005);
and UO_2616 (O_2616,N_23890,N_23094);
nor UO_2617 (O_2617,N_21654,N_22928);
xnor UO_2618 (O_2618,N_23013,N_23125);
nand UO_2619 (O_2619,N_24943,N_24085);
xnor UO_2620 (O_2620,N_20208,N_22062);
or UO_2621 (O_2621,N_22542,N_20023);
nor UO_2622 (O_2622,N_24143,N_21014);
nor UO_2623 (O_2623,N_23148,N_21939);
and UO_2624 (O_2624,N_23399,N_24388);
nand UO_2625 (O_2625,N_24351,N_20105);
or UO_2626 (O_2626,N_21508,N_22951);
xor UO_2627 (O_2627,N_23366,N_20775);
or UO_2628 (O_2628,N_22523,N_22765);
and UO_2629 (O_2629,N_22837,N_23819);
and UO_2630 (O_2630,N_21089,N_23876);
or UO_2631 (O_2631,N_20104,N_24418);
or UO_2632 (O_2632,N_22466,N_20657);
xnor UO_2633 (O_2633,N_23344,N_24586);
or UO_2634 (O_2634,N_20099,N_21100);
nor UO_2635 (O_2635,N_24246,N_24933);
nor UO_2636 (O_2636,N_20191,N_22719);
and UO_2637 (O_2637,N_22528,N_21660);
or UO_2638 (O_2638,N_22641,N_24839);
nor UO_2639 (O_2639,N_23293,N_20248);
and UO_2640 (O_2640,N_20727,N_20610);
nor UO_2641 (O_2641,N_20020,N_20813);
nor UO_2642 (O_2642,N_24418,N_20026);
or UO_2643 (O_2643,N_24134,N_22102);
or UO_2644 (O_2644,N_23897,N_24133);
nand UO_2645 (O_2645,N_23441,N_23175);
nor UO_2646 (O_2646,N_24304,N_20322);
and UO_2647 (O_2647,N_23710,N_20542);
and UO_2648 (O_2648,N_24600,N_20067);
nand UO_2649 (O_2649,N_20345,N_20581);
and UO_2650 (O_2650,N_20674,N_21655);
nor UO_2651 (O_2651,N_20591,N_22349);
and UO_2652 (O_2652,N_20942,N_20346);
nor UO_2653 (O_2653,N_23247,N_23898);
and UO_2654 (O_2654,N_21924,N_22870);
nor UO_2655 (O_2655,N_20760,N_23281);
nor UO_2656 (O_2656,N_22914,N_22620);
nand UO_2657 (O_2657,N_24364,N_23454);
nor UO_2658 (O_2658,N_23800,N_21513);
nor UO_2659 (O_2659,N_24813,N_20434);
and UO_2660 (O_2660,N_22745,N_22446);
nor UO_2661 (O_2661,N_23793,N_21337);
nor UO_2662 (O_2662,N_22275,N_20971);
nand UO_2663 (O_2663,N_20365,N_23006);
nand UO_2664 (O_2664,N_21032,N_21894);
and UO_2665 (O_2665,N_22889,N_22270);
nand UO_2666 (O_2666,N_23151,N_24002);
nor UO_2667 (O_2667,N_24076,N_23275);
nor UO_2668 (O_2668,N_24577,N_20529);
xnor UO_2669 (O_2669,N_24939,N_24964);
nor UO_2670 (O_2670,N_21248,N_24342);
or UO_2671 (O_2671,N_20081,N_23146);
and UO_2672 (O_2672,N_24623,N_21064);
or UO_2673 (O_2673,N_20505,N_22017);
nor UO_2674 (O_2674,N_24675,N_24410);
nor UO_2675 (O_2675,N_22096,N_24514);
or UO_2676 (O_2676,N_21704,N_23455);
nor UO_2677 (O_2677,N_22414,N_21739);
nand UO_2678 (O_2678,N_23423,N_21314);
or UO_2679 (O_2679,N_21428,N_20799);
and UO_2680 (O_2680,N_23133,N_22846);
and UO_2681 (O_2681,N_24162,N_23298);
nor UO_2682 (O_2682,N_21211,N_23210);
nand UO_2683 (O_2683,N_22794,N_23815);
nand UO_2684 (O_2684,N_21887,N_22698);
nor UO_2685 (O_2685,N_23735,N_24469);
nor UO_2686 (O_2686,N_20440,N_22860);
and UO_2687 (O_2687,N_22430,N_24571);
xor UO_2688 (O_2688,N_21246,N_20807);
nor UO_2689 (O_2689,N_22032,N_22919);
nand UO_2690 (O_2690,N_20659,N_23643);
nor UO_2691 (O_2691,N_22992,N_20522);
xnor UO_2692 (O_2692,N_24312,N_22525);
nor UO_2693 (O_2693,N_23472,N_24217);
and UO_2694 (O_2694,N_21262,N_20395);
nor UO_2695 (O_2695,N_22261,N_20099);
xnor UO_2696 (O_2696,N_22808,N_24495);
nand UO_2697 (O_2697,N_21262,N_23683);
or UO_2698 (O_2698,N_22314,N_21066);
and UO_2699 (O_2699,N_22529,N_20733);
and UO_2700 (O_2700,N_23560,N_22078);
or UO_2701 (O_2701,N_23151,N_20464);
or UO_2702 (O_2702,N_23935,N_23590);
nor UO_2703 (O_2703,N_24241,N_21501);
nand UO_2704 (O_2704,N_20915,N_21524);
or UO_2705 (O_2705,N_23176,N_20095);
nor UO_2706 (O_2706,N_20180,N_21133);
nor UO_2707 (O_2707,N_24899,N_20741);
or UO_2708 (O_2708,N_22771,N_24106);
or UO_2709 (O_2709,N_22270,N_22365);
nor UO_2710 (O_2710,N_22992,N_20576);
nand UO_2711 (O_2711,N_22086,N_23025);
nand UO_2712 (O_2712,N_24859,N_23622);
and UO_2713 (O_2713,N_24287,N_23574);
and UO_2714 (O_2714,N_20674,N_24316);
nor UO_2715 (O_2715,N_22557,N_20547);
and UO_2716 (O_2716,N_24533,N_21873);
nand UO_2717 (O_2717,N_22807,N_23282);
and UO_2718 (O_2718,N_21035,N_24660);
nor UO_2719 (O_2719,N_22897,N_22738);
nor UO_2720 (O_2720,N_21185,N_21385);
nand UO_2721 (O_2721,N_23688,N_24808);
xnor UO_2722 (O_2722,N_20182,N_21044);
xnor UO_2723 (O_2723,N_23350,N_21644);
or UO_2724 (O_2724,N_22442,N_21432);
xnor UO_2725 (O_2725,N_22808,N_21432);
nor UO_2726 (O_2726,N_23336,N_21155);
nand UO_2727 (O_2727,N_24003,N_22665);
nor UO_2728 (O_2728,N_24153,N_22808);
and UO_2729 (O_2729,N_21918,N_24937);
and UO_2730 (O_2730,N_24184,N_20708);
nand UO_2731 (O_2731,N_24598,N_21365);
xnor UO_2732 (O_2732,N_21968,N_20428);
or UO_2733 (O_2733,N_20402,N_22815);
and UO_2734 (O_2734,N_23520,N_22710);
nand UO_2735 (O_2735,N_22279,N_24314);
nor UO_2736 (O_2736,N_20322,N_21069);
nand UO_2737 (O_2737,N_21717,N_20437);
and UO_2738 (O_2738,N_22287,N_22509);
or UO_2739 (O_2739,N_21778,N_23224);
and UO_2740 (O_2740,N_20137,N_20314);
and UO_2741 (O_2741,N_24668,N_24388);
nand UO_2742 (O_2742,N_22255,N_21760);
and UO_2743 (O_2743,N_22590,N_20372);
nand UO_2744 (O_2744,N_21549,N_24012);
nand UO_2745 (O_2745,N_22559,N_24758);
nand UO_2746 (O_2746,N_24077,N_20052);
nand UO_2747 (O_2747,N_22731,N_21782);
or UO_2748 (O_2748,N_24520,N_23259);
nor UO_2749 (O_2749,N_23341,N_23679);
and UO_2750 (O_2750,N_23785,N_21468);
and UO_2751 (O_2751,N_21352,N_24350);
or UO_2752 (O_2752,N_21703,N_20699);
nand UO_2753 (O_2753,N_23108,N_23730);
xnor UO_2754 (O_2754,N_21695,N_23733);
and UO_2755 (O_2755,N_20976,N_20629);
nand UO_2756 (O_2756,N_24422,N_20948);
or UO_2757 (O_2757,N_22053,N_24917);
and UO_2758 (O_2758,N_23916,N_21065);
or UO_2759 (O_2759,N_24135,N_21742);
nand UO_2760 (O_2760,N_23988,N_24625);
or UO_2761 (O_2761,N_24425,N_20309);
nand UO_2762 (O_2762,N_21276,N_24143);
nor UO_2763 (O_2763,N_20165,N_22963);
nand UO_2764 (O_2764,N_21727,N_22851);
and UO_2765 (O_2765,N_20312,N_20398);
and UO_2766 (O_2766,N_24847,N_22960);
and UO_2767 (O_2767,N_22367,N_21788);
xnor UO_2768 (O_2768,N_24036,N_21456);
nand UO_2769 (O_2769,N_22567,N_21998);
nand UO_2770 (O_2770,N_23291,N_23285);
nand UO_2771 (O_2771,N_24974,N_23556);
or UO_2772 (O_2772,N_21347,N_20184);
and UO_2773 (O_2773,N_23078,N_24697);
nor UO_2774 (O_2774,N_21256,N_22876);
or UO_2775 (O_2775,N_21224,N_23144);
or UO_2776 (O_2776,N_22926,N_22937);
or UO_2777 (O_2777,N_24629,N_22395);
nand UO_2778 (O_2778,N_20626,N_22899);
nand UO_2779 (O_2779,N_20406,N_21421);
and UO_2780 (O_2780,N_21305,N_24614);
nand UO_2781 (O_2781,N_22304,N_23069);
nor UO_2782 (O_2782,N_21685,N_22368);
and UO_2783 (O_2783,N_23674,N_24829);
or UO_2784 (O_2784,N_20837,N_24474);
nand UO_2785 (O_2785,N_22434,N_20382);
or UO_2786 (O_2786,N_22255,N_24364);
and UO_2787 (O_2787,N_24641,N_22699);
nor UO_2788 (O_2788,N_24968,N_22895);
nand UO_2789 (O_2789,N_20360,N_20443);
and UO_2790 (O_2790,N_23212,N_24780);
and UO_2791 (O_2791,N_24726,N_24982);
or UO_2792 (O_2792,N_24663,N_20111);
and UO_2793 (O_2793,N_24419,N_22119);
nor UO_2794 (O_2794,N_24376,N_21274);
and UO_2795 (O_2795,N_21325,N_23114);
nand UO_2796 (O_2796,N_21060,N_23657);
xnor UO_2797 (O_2797,N_24990,N_23131);
nand UO_2798 (O_2798,N_20380,N_20526);
or UO_2799 (O_2799,N_21973,N_22691);
nor UO_2800 (O_2800,N_22109,N_22291);
and UO_2801 (O_2801,N_24285,N_21637);
nand UO_2802 (O_2802,N_21823,N_24098);
or UO_2803 (O_2803,N_23011,N_23211);
nor UO_2804 (O_2804,N_24035,N_20633);
nand UO_2805 (O_2805,N_24969,N_20823);
nand UO_2806 (O_2806,N_22120,N_20296);
nand UO_2807 (O_2807,N_21744,N_20848);
and UO_2808 (O_2808,N_23995,N_21548);
nor UO_2809 (O_2809,N_21389,N_24631);
and UO_2810 (O_2810,N_21160,N_22341);
or UO_2811 (O_2811,N_21804,N_22692);
or UO_2812 (O_2812,N_21511,N_20026);
nand UO_2813 (O_2813,N_21316,N_20116);
xnor UO_2814 (O_2814,N_22991,N_24594);
nand UO_2815 (O_2815,N_22696,N_20082);
nand UO_2816 (O_2816,N_23709,N_23392);
and UO_2817 (O_2817,N_24235,N_22521);
and UO_2818 (O_2818,N_21919,N_20557);
nor UO_2819 (O_2819,N_23610,N_20968);
nor UO_2820 (O_2820,N_23668,N_23577);
xnor UO_2821 (O_2821,N_20543,N_21410);
and UO_2822 (O_2822,N_24402,N_23041);
nor UO_2823 (O_2823,N_20009,N_20761);
nor UO_2824 (O_2824,N_21941,N_22377);
or UO_2825 (O_2825,N_22949,N_21926);
or UO_2826 (O_2826,N_24622,N_22866);
nand UO_2827 (O_2827,N_23499,N_21216);
nor UO_2828 (O_2828,N_21466,N_21042);
or UO_2829 (O_2829,N_21846,N_24290);
nand UO_2830 (O_2830,N_24441,N_22810);
nor UO_2831 (O_2831,N_23610,N_23177);
or UO_2832 (O_2832,N_21833,N_21035);
nand UO_2833 (O_2833,N_23679,N_22986);
and UO_2834 (O_2834,N_22973,N_21291);
or UO_2835 (O_2835,N_21764,N_21674);
nand UO_2836 (O_2836,N_20014,N_23273);
and UO_2837 (O_2837,N_24461,N_20638);
nor UO_2838 (O_2838,N_22202,N_21946);
or UO_2839 (O_2839,N_21129,N_24942);
nand UO_2840 (O_2840,N_23844,N_23399);
nor UO_2841 (O_2841,N_23506,N_23518);
and UO_2842 (O_2842,N_21939,N_23070);
or UO_2843 (O_2843,N_21546,N_21394);
and UO_2844 (O_2844,N_24783,N_24955);
or UO_2845 (O_2845,N_21861,N_23891);
and UO_2846 (O_2846,N_21446,N_20347);
and UO_2847 (O_2847,N_21576,N_22741);
nor UO_2848 (O_2848,N_20891,N_23863);
and UO_2849 (O_2849,N_24325,N_23192);
nand UO_2850 (O_2850,N_21806,N_23373);
or UO_2851 (O_2851,N_23434,N_21841);
xnor UO_2852 (O_2852,N_21762,N_20603);
nor UO_2853 (O_2853,N_21349,N_22151);
xnor UO_2854 (O_2854,N_20265,N_22828);
and UO_2855 (O_2855,N_22608,N_24972);
xor UO_2856 (O_2856,N_24449,N_20569);
nor UO_2857 (O_2857,N_22902,N_23318);
nor UO_2858 (O_2858,N_22595,N_20249);
nand UO_2859 (O_2859,N_24666,N_21944);
nand UO_2860 (O_2860,N_20914,N_22169);
nor UO_2861 (O_2861,N_24145,N_22298);
or UO_2862 (O_2862,N_21911,N_20815);
xnor UO_2863 (O_2863,N_22636,N_24890);
nor UO_2864 (O_2864,N_23476,N_22263);
and UO_2865 (O_2865,N_21552,N_20253);
nand UO_2866 (O_2866,N_24388,N_21736);
nand UO_2867 (O_2867,N_21779,N_20444);
or UO_2868 (O_2868,N_21842,N_21284);
nor UO_2869 (O_2869,N_23845,N_24288);
nand UO_2870 (O_2870,N_23092,N_24236);
nor UO_2871 (O_2871,N_20986,N_22808);
nand UO_2872 (O_2872,N_24189,N_24954);
nand UO_2873 (O_2873,N_23445,N_21525);
nor UO_2874 (O_2874,N_23101,N_23664);
nor UO_2875 (O_2875,N_24456,N_21263);
nand UO_2876 (O_2876,N_20523,N_20283);
or UO_2877 (O_2877,N_22793,N_22459);
or UO_2878 (O_2878,N_21672,N_24378);
nand UO_2879 (O_2879,N_22011,N_24990);
nor UO_2880 (O_2880,N_21325,N_22010);
and UO_2881 (O_2881,N_24809,N_20800);
and UO_2882 (O_2882,N_20319,N_21020);
and UO_2883 (O_2883,N_23791,N_24094);
nor UO_2884 (O_2884,N_22247,N_22278);
and UO_2885 (O_2885,N_21419,N_21996);
and UO_2886 (O_2886,N_22338,N_22762);
or UO_2887 (O_2887,N_23456,N_23244);
xnor UO_2888 (O_2888,N_20932,N_22260);
nor UO_2889 (O_2889,N_23373,N_20498);
and UO_2890 (O_2890,N_23006,N_20183);
and UO_2891 (O_2891,N_24150,N_23056);
nand UO_2892 (O_2892,N_21255,N_20655);
nor UO_2893 (O_2893,N_21677,N_22277);
or UO_2894 (O_2894,N_20432,N_21368);
and UO_2895 (O_2895,N_24341,N_23765);
or UO_2896 (O_2896,N_23779,N_22768);
and UO_2897 (O_2897,N_21706,N_24311);
nand UO_2898 (O_2898,N_21550,N_24389);
and UO_2899 (O_2899,N_20022,N_23153);
and UO_2900 (O_2900,N_20592,N_24385);
and UO_2901 (O_2901,N_21371,N_23230);
nor UO_2902 (O_2902,N_21323,N_22471);
xor UO_2903 (O_2903,N_21832,N_22279);
nor UO_2904 (O_2904,N_22868,N_20441);
and UO_2905 (O_2905,N_21597,N_24502);
and UO_2906 (O_2906,N_20525,N_23137);
nor UO_2907 (O_2907,N_23261,N_22522);
xnor UO_2908 (O_2908,N_23181,N_24659);
nor UO_2909 (O_2909,N_22727,N_23863);
nor UO_2910 (O_2910,N_23589,N_21236);
and UO_2911 (O_2911,N_23297,N_20327);
and UO_2912 (O_2912,N_22975,N_22200);
nor UO_2913 (O_2913,N_24192,N_23712);
and UO_2914 (O_2914,N_23539,N_23583);
or UO_2915 (O_2915,N_20389,N_23929);
and UO_2916 (O_2916,N_23701,N_21866);
nand UO_2917 (O_2917,N_21705,N_22335);
and UO_2918 (O_2918,N_21112,N_24953);
and UO_2919 (O_2919,N_21307,N_21984);
nor UO_2920 (O_2920,N_24218,N_21830);
and UO_2921 (O_2921,N_24597,N_20482);
nor UO_2922 (O_2922,N_24443,N_22435);
and UO_2923 (O_2923,N_20552,N_22981);
nor UO_2924 (O_2924,N_23811,N_21867);
nand UO_2925 (O_2925,N_22751,N_22266);
nor UO_2926 (O_2926,N_24762,N_24507);
nor UO_2927 (O_2927,N_23820,N_20237);
xor UO_2928 (O_2928,N_21041,N_21163);
nor UO_2929 (O_2929,N_21467,N_23144);
nand UO_2930 (O_2930,N_24639,N_21163);
nor UO_2931 (O_2931,N_23268,N_21791);
nor UO_2932 (O_2932,N_20711,N_20330);
and UO_2933 (O_2933,N_23444,N_20598);
xnor UO_2934 (O_2934,N_22218,N_22748);
nor UO_2935 (O_2935,N_20775,N_21184);
nor UO_2936 (O_2936,N_21782,N_23298);
nor UO_2937 (O_2937,N_20147,N_21750);
nor UO_2938 (O_2938,N_20230,N_22079);
or UO_2939 (O_2939,N_21415,N_24730);
or UO_2940 (O_2940,N_20117,N_20933);
nor UO_2941 (O_2941,N_24368,N_22405);
and UO_2942 (O_2942,N_24967,N_22739);
and UO_2943 (O_2943,N_24850,N_21773);
or UO_2944 (O_2944,N_24337,N_23633);
and UO_2945 (O_2945,N_22275,N_24493);
nand UO_2946 (O_2946,N_24317,N_22041);
nand UO_2947 (O_2947,N_23272,N_24017);
and UO_2948 (O_2948,N_24445,N_22714);
or UO_2949 (O_2949,N_22927,N_21044);
nor UO_2950 (O_2950,N_24765,N_22750);
or UO_2951 (O_2951,N_21263,N_23648);
and UO_2952 (O_2952,N_23511,N_22096);
and UO_2953 (O_2953,N_21545,N_23954);
or UO_2954 (O_2954,N_20302,N_23501);
or UO_2955 (O_2955,N_24565,N_20636);
nand UO_2956 (O_2956,N_22497,N_22477);
and UO_2957 (O_2957,N_21731,N_20411);
nand UO_2958 (O_2958,N_22224,N_20073);
and UO_2959 (O_2959,N_23958,N_22133);
and UO_2960 (O_2960,N_20655,N_23238);
and UO_2961 (O_2961,N_20057,N_20452);
or UO_2962 (O_2962,N_24924,N_23880);
and UO_2963 (O_2963,N_20883,N_24931);
or UO_2964 (O_2964,N_24686,N_24604);
nor UO_2965 (O_2965,N_24257,N_24863);
or UO_2966 (O_2966,N_23627,N_21220);
or UO_2967 (O_2967,N_22559,N_21939);
nor UO_2968 (O_2968,N_24500,N_22564);
and UO_2969 (O_2969,N_23810,N_20905);
xnor UO_2970 (O_2970,N_24765,N_22784);
nor UO_2971 (O_2971,N_24060,N_22957);
nand UO_2972 (O_2972,N_22155,N_22245);
nand UO_2973 (O_2973,N_22280,N_24554);
nand UO_2974 (O_2974,N_20892,N_23080);
or UO_2975 (O_2975,N_22128,N_20776);
and UO_2976 (O_2976,N_21986,N_22306);
or UO_2977 (O_2977,N_22101,N_23577);
and UO_2978 (O_2978,N_24070,N_22500);
nor UO_2979 (O_2979,N_22795,N_21332);
xor UO_2980 (O_2980,N_20042,N_22456);
nand UO_2981 (O_2981,N_21203,N_24363);
and UO_2982 (O_2982,N_24708,N_24599);
nand UO_2983 (O_2983,N_20697,N_20445);
or UO_2984 (O_2984,N_24604,N_21939);
and UO_2985 (O_2985,N_23241,N_22531);
nor UO_2986 (O_2986,N_24715,N_22468);
nand UO_2987 (O_2987,N_20358,N_21354);
xor UO_2988 (O_2988,N_22545,N_24428);
nand UO_2989 (O_2989,N_21172,N_24638);
or UO_2990 (O_2990,N_24331,N_22042);
or UO_2991 (O_2991,N_22251,N_23117);
and UO_2992 (O_2992,N_22615,N_22535);
nand UO_2993 (O_2993,N_24446,N_22492);
nor UO_2994 (O_2994,N_20116,N_24161);
nand UO_2995 (O_2995,N_22333,N_21401);
or UO_2996 (O_2996,N_24684,N_23158);
or UO_2997 (O_2997,N_24058,N_22629);
or UO_2998 (O_2998,N_21547,N_24529);
xnor UO_2999 (O_2999,N_20146,N_22147);
endmodule