module basic_1000_10000_1500_2_levels_1xor_7(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5002,N_5003,N_5004,N_5007,N_5008,N_5011,N_5012,N_5013,N_5015,N_5016,N_5017,N_5018,N_5021,N_5022,N_5025,N_5027,N_5028,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5038,N_5039,N_5043,N_5044,N_5045,N_5046,N_5047,N_5049,N_5050,N_5052,N_5053,N_5054,N_5055,N_5059,N_5063,N_5065,N_5067,N_5068,N_5069,N_5071,N_5073,N_5074,N_5075,N_5076,N_5077,N_5080,N_5084,N_5085,N_5089,N_5090,N_5091,N_5093,N_5094,N_5096,N_5097,N_5099,N_5100,N_5102,N_5104,N_5105,N_5106,N_5108,N_5110,N_5112,N_5114,N_5115,N_5116,N_5117,N_5118,N_5123,N_5124,N_5126,N_5127,N_5128,N_5130,N_5131,N_5133,N_5135,N_5137,N_5138,N_5140,N_5141,N_5145,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5159,N_5162,N_5163,N_5164,N_5166,N_5169,N_5170,N_5171,N_5173,N_5175,N_5176,N_5177,N_5178,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5191,N_5192,N_5194,N_5197,N_5199,N_5200,N_5203,N_5204,N_5205,N_5206,N_5208,N_5209,N_5210,N_5211,N_5214,N_5215,N_5216,N_5217,N_5219,N_5220,N_5221,N_5222,N_5225,N_5226,N_5227,N_5228,N_5230,N_5231,N_5232,N_5236,N_5237,N_5238,N_5239,N_5240,N_5243,N_5244,N_5247,N_5248,N_5249,N_5250,N_5251,N_5253,N_5255,N_5259,N_5263,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5276,N_5278,N_5279,N_5280,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5290,N_5292,N_5293,N_5295,N_5296,N_5298,N_5299,N_5300,N_5301,N_5303,N_5306,N_5309,N_5312,N_5314,N_5315,N_5316,N_5318,N_5320,N_5321,N_5322,N_5324,N_5328,N_5329,N_5332,N_5334,N_5335,N_5337,N_5338,N_5339,N_5340,N_5342,N_5343,N_5344,N_5347,N_5348,N_5351,N_5354,N_5356,N_5357,N_5358,N_5361,N_5363,N_5364,N_5366,N_5368,N_5373,N_5375,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5391,N_5394,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5405,N_5407,N_5409,N_5410,N_5411,N_5412,N_5413,N_5415,N_5417,N_5422,N_5423,N_5424,N_5425,N_5430,N_5432,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5441,N_5442,N_5443,N_5446,N_5447,N_5448,N_5451,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5461,N_5463,N_5466,N_5469,N_5471,N_5473,N_5474,N_5475,N_5480,N_5481,N_5483,N_5484,N_5485,N_5486,N_5487,N_5489,N_5490,N_5493,N_5497,N_5498,N_5499,N_5500,N_5504,N_5507,N_5508,N_5509,N_5510,N_5515,N_5516,N_5517,N_5519,N_5521,N_5522,N_5523,N_5525,N_5526,N_5529,N_5532,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5552,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5562,N_5564,N_5565,N_5566,N_5567,N_5569,N_5571,N_5572,N_5573,N_5576,N_5577,N_5578,N_5579,N_5581,N_5582,N_5583,N_5585,N_5590,N_5595,N_5596,N_5598,N_5599,N_5602,N_5603,N_5608,N_5609,N_5610,N_5612,N_5614,N_5615,N_5616,N_5618,N_5622,N_5623,N_5627,N_5628,N_5629,N_5631,N_5632,N_5636,N_5638,N_5639,N_5640,N_5641,N_5644,N_5646,N_5647,N_5651,N_5654,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5665,N_5666,N_5668,N_5670,N_5671,N_5673,N_5674,N_5675,N_5676,N_5677,N_5679,N_5680,N_5681,N_5682,N_5686,N_5687,N_5688,N_5689,N_5692,N_5693,N_5694,N_5697,N_5698,N_5699,N_5703,N_5704,N_5705,N_5708,N_5709,N_5711,N_5712,N_5716,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5727,N_5728,N_5729,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5743,N_5745,N_5747,N_5749,N_5751,N_5752,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5761,N_5762,N_5763,N_5764,N_5766,N_5767,N_5769,N_5770,N_5772,N_5776,N_5777,N_5778,N_5779,N_5781,N_5782,N_5784,N_5786,N_5790,N_5792,N_5794,N_5795,N_5798,N_5799,N_5800,N_5801,N_5803,N_5804,N_5805,N_5807,N_5808,N_5809,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5823,N_5824,N_5825,N_5826,N_5828,N_5829,N_5834,N_5835,N_5837,N_5838,N_5839,N_5841,N_5842,N_5843,N_5844,N_5849,N_5851,N_5852,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5871,N_5872,N_5874,N_5875,N_5876,N_5879,N_5881,N_5882,N_5887,N_5889,N_5890,N_5892,N_5895,N_5896,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5910,N_5914,N_5918,N_5920,N_5921,N_5924,N_5925,N_5926,N_5927,N_5932,N_5933,N_5934,N_5936,N_5939,N_5940,N_5941,N_5946,N_5947,N_5948,N_5949,N_5951,N_5952,N_5954,N_5956,N_5957,N_5958,N_5959,N_5960,N_5962,N_5963,N_5964,N_5965,N_5966,N_5969,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5980,N_5981,N_5985,N_5986,N_5989,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6005,N_6006,N_6007,N_6009,N_6010,N_6011,N_6013,N_6014,N_6015,N_6017,N_6019,N_6021,N_6022,N_6023,N_6025,N_6027,N_6032,N_6033,N_6035,N_6037,N_6038,N_6041,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6053,N_6054,N_6056,N_6057,N_6059,N_6061,N_6062,N_6063,N_6064,N_6066,N_6067,N_6068,N_6070,N_6071,N_6072,N_6073,N_6077,N_6078,N_6079,N_6080,N_6083,N_6084,N_6086,N_6087,N_6089,N_6090,N_6091,N_6094,N_6096,N_6098,N_6099,N_6101,N_6102,N_6105,N_6107,N_6109,N_6110,N_6112,N_6114,N_6118,N_6120,N_6121,N_6122,N_6124,N_6125,N_6126,N_6127,N_6130,N_6131,N_6132,N_6134,N_6139,N_6140,N_6141,N_6143,N_6149,N_6150,N_6152,N_6153,N_6154,N_6155,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6165,N_6166,N_6167,N_6169,N_6170,N_6171,N_6172,N_6173,N_6175,N_6177,N_6178,N_6179,N_6181,N_6182,N_6183,N_6185,N_6186,N_6191,N_6192,N_6193,N_6195,N_6198,N_6200,N_6204,N_6205,N_6206,N_6208,N_6210,N_6211,N_6212,N_6216,N_6217,N_6218,N_6219,N_6220,N_6223,N_6224,N_6225,N_6226,N_6228,N_6229,N_6232,N_6234,N_6237,N_6238,N_6239,N_6240,N_6241,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6253,N_6254,N_6255,N_6256,N_6257,N_6259,N_6261,N_6262,N_6263,N_6266,N_6269,N_6270,N_6271,N_6272,N_6275,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6291,N_6292,N_6293,N_6295,N_6297,N_6298,N_6299,N_6304,N_6306,N_6308,N_6309,N_6310,N_6313,N_6315,N_6316,N_6318,N_6319,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6343,N_6344,N_6347,N_6348,N_6350,N_6353,N_6354,N_6355,N_6362,N_6363,N_6364,N_6367,N_6368,N_6369,N_6373,N_6375,N_6376,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6390,N_6391,N_6393,N_6397,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6406,N_6409,N_6410,N_6412,N_6413,N_6414,N_6415,N_6419,N_6420,N_6422,N_6423,N_6424,N_6426,N_6427,N_6428,N_6429,N_6431,N_6432,N_6433,N_6434,N_6435,N_6437,N_6438,N_6439,N_6442,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6454,N_6455,N_6458,N_6459,N_6460,N_6465,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6480,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6492,N_6494,N_6495,N_6496,N_6498,N_6499,N_6500,N_6503,N_6505,N_6509,N_6510,N_6511,N_6512,N_6514,N_6518,N_6519,N_6521,N_6522,N_6523,N_6524,N_6525,N_6528,N_6534,N_6535,N_6536,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6547,N_6552,N_6554,N_6558,N_6559,N_6560,N_6561,N_6564,N_6566,N_6568,N_6569,N_6570,N_6572,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6582,N_6584,N_6585,N_6586,N_6589,N_6595,N_6598,N_6599,N_6601,N_6602,N_6605,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6620,N_6621,N_6623,N_6624,N_6628,N_6629,N_6630,N_6632,N_6634,N_6635,N_6636,N_6638,N_6639,N_6640,N_6644,N_6645,N_6648,N_6653,N_6654,N_6655,N_6657,N_6658,N_6661,N_6662,N_6664,N_6668,N_6671,N_6673,N_6674,N_6676,N_6677,N_6678,N_6679,N_6683,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6703,N_6704,N_6706,N_6707,N_6708,N_6709,N_6710,N_6712,N_6713,N_6714,N_6715,N_6717,N_6718,N_6719,N_6720,N_6722,N_6723,N_6725,N_6726,N_6727,N_6730,N_6732,N_6734,N_6737,N_6738,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6749,N_6751,N_6752,N_6753,N_6755,N_6756,N_6759,N_6760,N_6762,N_6763,N_6764,N_6767,N_6769,N_6771,N_6774,N_6775,N_6776,N_6779,N_6783,N_6784,N_6788,N_6789,N_6790,N_6794,N_6795,N_6797,N_6798,N_6799,N_6801,N_6802,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6812,N_6813,N_6814,N_6817,N_6818,N_6819,N_6820,N_6821,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6846,N_6847,N_6849,N_6852,N_6853,N_6855,N_6856,N_6858,N_6859,N_6862,N_6863,N_6864,N_6865,N_6866,N_6868,N_6870,N_6871,N_6872,N_6873,N_6874,N_6876,N_6878,N_6879,N_6880,N_6882,N_6883,N_6884,N_6885,N_6887,N_6890,N_6891,N_6892,N_6895,N_6896,N_6897,N_6898,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6909,N_6912,N_6913,N_6914,N_6915,N_6918,N_6919,N_6920,N_6922,N_6925,N_6927,N_6930,N_6931,N_6932,N_6934,N_6935,N_6936,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6946,N_6948,N_6950,N_6951,N_6952,N_6956,N_6957,N_6958,N_6959,N_6962,N_6963,N_6964,N_6965,N_6966,N_6971,N_6973,N_6975,N_6977,N_6978,N_6980,N_6981,N_6982,N_6985,N_6989,N_6990,N_6994,N_6996,N_6998,N_6999,N_7001,N_7002,N_7006,N_7007,N_7009,N_7010,N_7011,N_7015,N_7016,N_7017,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7030,N_7031,N_7032,N_7037,N_7038,N_7041,N_7043,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7063,N_7064,N_7065,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7078,N_7083,N_7085,N_7086,N_7088,N_7090,N_7091,N_7093,N_7094,N_7097,N_7098,N_7100,N_7104,N_7106,N_7109,N_7111,N_7114,N_7115,N_7117,N_7118,N_7119,N_7120,N_7125,N_7127,N_7130,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7142,N_7144,N_7145,N_7146,N_7148,N_7152,N_7158,N_7159,N_7161,N_7164,N_7165,N_7168,N_7170,N_7171,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7180,N_7181,N_7182,N_7186,N_7187,N_7189,N_7194,N_7195,N_7198,N_7199,N_7200,N_7202,N_7203,N_7205,N_7210,N_7214,N_7216,N_7218,N_7221,N_7222,N_7223,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7232,N_7233,N_7234,N_7235,N_7238,N_7240,N_7241,N_7244,N_7245,N_7247,N_7248,N_7249,N_7250,N_7252,N_7254,N_7255,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7264,N_7266,N_7268,N_7269,N_7270,N_7271,N_7273,N_7274,N_7275,N_7277,N_7279,N_7283,N_7284,N_7285,N_7289,N_7290,N_7294,N_7295,N_7296,N_7297,N_7299,N_7301,N_7302,N_7304,N_7305,N_7306,N_7307,N_7309,N_7312,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7334,N_7335,N_7336,N_7338,N_7339,N_7344,N_7345,N_7349,N_7350,N_7352,N_7353,N_7355,N_7358,N_7360,N_7362,N_7363,N_7365,N_7366,N_7368,N_7369,N_7372,N_7373,N_7374,N_7376,N_7377,N_7378,N_7379,N_7380,N_7384,N_7385,N_7387,N_7389,N_7391,N_7392,N_7393,N_7394,N_7396,N_7400,N_7403,N_7404,N_7406,N_7407,N_7408,N_7409,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7421,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7433,N_7434,N_7436,N_7438,N_7439,N_7441,N_7442,N_7443,N_7446,N_7447,N_7448,N_7450,N_7451,N_7455,N_7457,N_7458,N_7459,N_7463,N_7464,N_7465,N_7467,N_7468,N_7470,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7488,N_7491,N_7493,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7503,N_7505,N_7507,N_7508,N_7509,N_7511,N_7513,N_7514,N_7520,N_7521,N_7522,N_7523,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7541,N_7542,N_7544,N_7546,N_7550,N_7551,N_7553,N_7554,N_7555,N_7556,N_7558,N_7560,N_7563,N_7566,N_7567,N_7569,N_7572,N_7573,N_7574,N_7579,N_7580,N_7582,N_7584,N_7587,N_7588,N_7589,N_7591,N_7592,N_7593,N_7594,N_7596,N_7597,N_7598,N_7599,N_7601,N_7603,N_7604,N_7607,N_7608,N_7611,N_7612,N_7613,N_7614,N_7616,N_7617,N_7618,N_7620,N_7622,N_7623,N_7625,N_7627,N_7629,N_7630,N_7631,N_7634,N_7635,N_7636,N_7640,N_7641,N_7642,N_7643,N_7645,N_7646,N_7651,N_7652,N_7654,N_7656,N_7659,N_7661,N_7663,N_7664,N_7665,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7677,N_7678,N_7679,N_7681,N_7682,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7691,N_7692,N_7694,N_7695,N_7696,N_7700,N_7701,N_7703,N_7704,N_7706,N_7707,N_7711,N_7714,N_7715,N_7716,N_7718,N_7719,N_7720,N_7722,N_7725,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7736,N_7737,N_7741,N_7743,N_7746,N_7747,N_7750,N_7751,N_7752,N_7754,N_7755,N_7757,N_7761,N_7763,N_7764,N_7765,N_7769,N_7770,N_7774,N_7776,N_7777,N_7778,N_7780,N_7784,N_7785,N_7786,N_7787,N_7789,N_7790,N_7792,N_7793,N_7794,N_7797,N_7798,N_7799,N_7802,N_7803,N_7804,N_7805,N_7807,N_7808,N_7809,N_7810,N_7812,N_7813,N_7814,N_7815,N_7817,N_7819,N_7821,N_7823,N_7830,N_7831,N_7832,N_7834,N_7837,N_7838,N_7839,N_7841,N_7842,N_7843,N_7845,N_7846,N_7847,N_7850,N_7851,N_7857,N_7858,N_7862,N_7863,N_7867,N_7868,N_7869,N_7871,N_7872,N_7873,N_7877,N_7878,N_7882,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7893,N_7895,N_7896,N_7897,N_7899,N_7900,N_7902,N_7903,N_7905,N_7906,N_7907,N_7909,N_7912,N_7914,N_7915,N_7916,N_7918,N_7920,N_7921,N_7924,N_7925,N_7926,N_7927,N_7928,N_7930,N_7931,N_7933,N_7934,N_7936,N_7937,N_7939,N_7940,N_7942,N_7944,N_7945,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7968,N_7970,N_7971,N_7973,N_7974,N_7975,N_7976,N_7981,N_7982,N_7984,N_7985,N_7987,N_7988,N_7989,N_7990,N_7995,N_7996,N_7998,N_8001,N_8003,N_8006,N_8008,N_8010,N_8012,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8026,N_8027,N_8028,N_8029,N_8031,N_8032,N_8034,N_8035,N_8036,N_8040,N_8041,N_8045,N_8047,N_8048,N_8049,N_8050,N_8051,N_8053,N_8054,N_8055,N_8058,N_8059,N_8065,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8078,N_8080,N_8081,N_8083,N_8084,N_8086,N_8087,N_8092,N_8095,N_8097,N_8099,N_8100,N_8101,N_8103,N_8104,N_8105,N_8109,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8124,N_8127,N_8129,N_8130,N_8131,N_8132,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8143,N_8149,N_8150,N_8151,N_8153,N_8154,N_8156,N_8159,N_8162,N_8163,N_8165,N_8167,N_8169,N_8170,N_8171,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8181,N_8183,N_8184,N_8185,N_8187,N_8191,N_8194,N_8196,N_8197,N_8198,N_8200,N_8201,N_8205,N_8207,N_8208,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8219,N_8220,N_8221,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8230,N_8231,N_8234,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8264,N_8268,N_8269,N_8270,N_8274,N_8275,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8284,N_8285,N_8286,N_8289,N_8291,N_8292,N_8293,N_8295,N_8296,N_8297,N_8300,N_8302,N_8303,N_8306,N_8307,N_8309,N_8311,N_8312,N_8313,N_8316,N_8318,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8331,N_8332,N_8333,N_8336,N_8337,N_8339,N_8340,N_8342,N_8343,N_8344,N_8345,N_8348,N_8349,N_8350,N_8352,N_8353,N_8356,N_8358,N_8359,N_8362,N_8363,N_8365,N_8366,N_8371,N_8372,N_8374,N_8375,N_8376,N_8377,N_8379,N_8381,N_8382,N_8383,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8395,N_8397,N_8398,N_8399,N_8401,N_8402,N_8405,N_8406,N_8408,N_8410,N_8412,N_8415,N_8417,N_8418,N_8420,N_8422,N_8423,N_8424,N_8427,N_8428,N_8431,N_8433,N_8435,N_8437,N_8438,N_8439,N_8442,N_8445,N_8447,N_8448,N_8449,N_8450,N_8452,N_8453,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8462,N_8463,N_8464,N_8466,N_8467,N_8469,N_8470,N_8471,N_8473,N_8474,N_8477,N_8479,N_8484,N_8485,N_8486,N_8491,N_8494,N_8495,N_8496,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8505,N_8506,N_8511,N_8513,N_8514,N_8517,N_8519,N_8520,N_8522,N_8523,N_8524,N_8525,N_8527,N_8528,N_8529,N_8533,N_8534,N_8535,N_8537,N_8538,N_8539,N_8540,N_8542,N_8543,N_8544,N_8545,N_8547,N_8549,N_8552,N_8553,N_8554,N_8555,N_8557,N_8558,N_8562,N_8563,N_8566,N_8568,N_8569,N_8570,N_8574,N_8577,N_8578,N_8582,N_8583,N_8585,N_8586,N_8588,N_8590,N_8591,N_8592,N_8593,N_8595,N_8596,N_8597,N_8600,N_8603,N_8605,N_8606,N_8608,N_8609,N_8610,N_8612,N_8613,N_8614,N_8616,N_8617,N_8619,N_8620,N_8622,N_8623,N_8624,N_8625,N_8627,N_8632,N_8634,N_8635,N_8639,N_8641,N_8643,N_8647,N_8648,N_8649,N_8650,N_8652,N_8654,N_8656,N_8657,N_8659,N_8660,N_8661,N_8663,N_8664,N_8665,N_8667,N_8668,N_8670,N_8671,N_8674,N_8675,N_8677,N_8678,N_8680,N_8681,N_8682,N_8683,N_8687,N_8688,N_8689,N_8690,N_8691,N_8693,N_8695,N_8696,N_8698,N_8699,N_8701,N_8703,N_8705,N_8706,N_8707,N_8713,N_8715,N_8716,N_8717,N_8719,N_8720,N_8721,N_8722,N_8723,N_8727,N_8728,N_8730,N_8731,N_8735,N_8736,N_8738,N_8739,N_8741,N_8743,N_8748,N_8749,N_8751,N_8754,N_8755,N_8756,N_8761,N_8762,N_8763,N_8766,N_8767,N_8768,N_8771,N_8772,N_8773,N_8774,N_8777,N_8779,N_8780,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8801,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8810,N_8811,N_8812,N_8813,N_8815,N_8819,N_8820,N_8823,N_8824,N_8828,N_8830,N_8833,N_8834,N_8835,N_8836,N_8837,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8847,N_8848,N_8852,N_8853,N_8854,N_8855,N_8858,N_8859,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8876,N_8877,N_8878,N_8879,N_8883,N_8884,N_8885,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8894,N_8896,N_8899,N_8900,N_8902,N_8903,N_8904,N_8906,N_8907,N_8910,N_8911,N_8913,N_8916,N_8918,N_8919,N_8922,N_8923,N_8924,N_8925,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8936,N_8937,N_8938,N_8939,N_8940,N_8942,N_8943,N_8945,N_8946,N_8948,N_8950,N_8951,N_8952,N_8953,N_8955,N_8957,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8978,N_8979,N_8982,N_8983,N_8984,N_8986,N_8988,N_8993,N_8994,N_8995,N_8997,N_9003,N_9004,N_9005,N_9006,N_9007,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9017,N_9019,N_9020,N_9023,N_9025,N_9026,N_9029,N_9030,N_9034,N_9035,N_9036,N_9038,N_9039,N_9040,N_9041,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9051,N_9053,N_9054,N_9056,N_9059,N_9060,N_9062,N_9063,N_9065,N_9067,N_9068,N_9070,N_9071,N_9072,N_9073,N_9074,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9089,N_9090,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9102,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9111,N_9112,N_9113,N_9115,N_9118,N_9120,N_9121,N_9123,N_9124,N_9125,N_9126,N_9128,N_9130,N_9132,N_9133,N_9134,N_9135,N_9137,N_9138,N_9139,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9149,N_9150,N_9151,N_9153,N_9154,N_9158,N_9159,N_9160,N_9161,N_9164,N_9165,N_9167,N_9168,N_9169,N_9171,N_9173,N_9174,N_9175,N_9176,N_9180,N_9181,N_9182,N_9189,N_9190,N_9191,N_9193,N_9194,N_9197,N_9198,N_9200,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9210,N_9212,N_9213,N_9216,N_9217,N_9218,N_9219,N_9220,N_9222,N_9223,N_9229,N_9231,N_9233,N_9234,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9246,N_9248,N_9249,N_9250,N_9251,N_9252,N_9258,N_9259,N_9260,N_9264,N_9265,N_9266,N_9268,N_9269,N_9270,N_9271,N_9272,N_9274,N_9275,N_9277,N_9279,N_9280,N_9281,N_9284,N_9285,N_9287,N_9289,N_9291,N_9293,N_9294,N_9297,N_9300,N_9301,N_9303,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9312,N_9314,N_9315,N_9319,N_9321,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9335,N_9337,N_9340,N_9342,N_9343,N_9346,N_9347,N_9348,N_9351,N_9352,N_9357,N_9358,N_9359,N_9360,N_9361,N_9363,N_9365,N_9366,N_9368,N_9369,N_9373,N_9374,N_9375,N_9376,N_9378,N_9379,N_9380,N_9383,N_9385,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9400,N_9403,N_9406,N_9409,N_9410,N_9412,N_9415,N_9416,N_9417,N_9419,N_9423,N_9424,N_9426,N_9433,N_9434,N_9436,N_9438,N_9439,N_9441,N_9442,N_9443,N_9444,N_9446,N_9449,N_9450,N_9453,N_9455,N_9460,N_9461,N_9463,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9472,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9495,N_9496,N_9499,N_9503,N_9504,N_9508,N_9509,N_9511,N_9512,N_9513,N_9515,N_9516,N_9518,N_9519,N_9520,N_9521,N_9522,N_9527,N_9532,N_9533,N_9535,N_9538,N_9539,N_9542,N_9543,N_9544,N_9549,N_9550,N_9553,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9564,N_9565,N_9567,N_9569,N_9572,N_9573,N_9574,N_9578,N_9581,N_9582,N_9583,N_9585,N_9586,N_9588,N_9589,N_9590,N_9596,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9607,N_9608,N_9609,N_9611,N_9612,N_9613,N_9614,N_9617,N_9618,N_9619,N_9621,N_9622,N_9623,N_9627,N_9628,N_9632,N_9633,N_9634,N_9635,N_9636,N_9638,N_9640,N_9641,N_9646,N_9649,N_9650,N_9654,N_9655,N_9656,N_9658,N_9659,N_9661,N_9662,N_9664,N_9665,N_9666,N_9667,N_9668,N_9670,N_9672,N_9673,N_9676,N_9677,N_9678,N_9679,N_9681,N_9683,N_9684,N_9686,N_9689,N_9690,N_9691,N_9692,N_9694,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9710,N_9711,N_9713,N_9714,N_9718,N_9726,N_9728,N_9733,N_9738,N_9739,N_9744,N_9746,N_9750,N_9752,N_9753,N_9754,N_9755,N_9757,N_9758,N_9761,N_9762,N_9763,N_9766,N_9767,N_9768,N_9769,N_9770,N_9773,N_9774,N_9775,N_9778,N_9779,N_9781,N_9782,N_9783,N_9784,N_9788,N_9790,N_9791,N_9792,N_9793,N_9796,N_9798,N_9801,N_9803,N_9804,N_9811,N_9812,N_9816,N_9817,N_9820,N_9823,N_9825,N_9828,N_9829,N_9831,N_9835,N_9836,N_9838,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9850,N_9851,N_9853,N_9856,N_9860,N_9862,N_9864,N_9865,N_9866,N_9867,N_9869,N_9871,N_9873,N_9874,N_9875,N_9876,N_9878,N_9883,N_9886,N_9888,N_9889,N_9890,N_9891,N_9893,N_9894,N_9895,N_9896,N_9899,N_9901,N_9902,N_9904,N_9905,N_9906,N_9908,N_9909,N_9911,N_9912,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9929,N_9931,N_9932,N_9933,N_9934,N_9936,N_9937,N_9939,N_9941,N_9942,N_9945,N_9946,N_9948,N_9949,N_9951,N_9952,N_9953,N_9955,N_9957,N_9960,N_9961,N_9962,N_9964,N_9965,N_9966,N_9967,N_9970,N_9971,N_9974,N_9975,N_9977,N_9978,N_9981,N_9982,N_9986,N_9988,N_9990,N_9992,N_9994,N_9995,N_9996,N_9998;
or U0 (N_0,In_62,In_379);
and U1 (N_1,In_866,In_954);
or U2 (N_2,In_128,In_160);
nand U3 (N_3,In_692,In_33);
and U4 (N_4,In_514,In_275);
nor U5 (N_5,In_237,In_783);
nor U6 (N_6,In_52,In_676);
or U7 (N_7,In_206,In_962);
nand U8 (N_8,In_842,In_386);
nor U9 (N_9,In_926,In_607);
and U10 (N_10,In_3,In_63);
nor U11 (N_11,In_891,In_222);
and U12 (N_12,In_967,In_277);
nand U13 (N_13,In_307,In_689);
and U14 (N_14,In_117,In_507);
nor U15 (N_15,In_677,In_569);
nand U16 (N_16,In_558,In_321);
and U17 (N_17,In_825,In_953);
and U18 (N_18,In_606,In_356);
and U19 (N_19,In_452,In_134);
nor U20 (N_20,In_732,In_887);
nor U21 (N_21,In_309,In_55);
or U22 (N_22,In_451,In_862);
nand U23 (N_23,In_700,In_845);
nor U24 (N_24,In_227,In_194);
nand U25 (N_25,In_699,In_369);
nor U26 (N_26,In_748,In_588);
or U27 (N_27,In_909,In_658);
nor U28 (N_28,In_453,In_805);
or U29 (N_29,In_879,In_565);
and U30 (N_30,In_491,In_621);
nand U31 (N_31,In_428,In_619);
and U32 (N_32,In_290,In_794);
or U33 (N_33,In_838,In_121);
nand U34 (N_34,In_422,In_200);
or U35 (N_35,In_168,In_178);
nand U36 (N_36,In_276,In_426);
nand U37 (N_37,In_1,In_877);
or U38 (N_38,In_934,In_939);
and U39 (N_39,In_305,In_482);
or U40 (N_40,In_601,In_343);
nand U41 (N_41,In_557,In_511);
nand U42 (N_42,In_720,In_522);
and U43 (N_43,In_424,In_314);
or U44 (N_44,In_9,In_544);
xor U45 (N_45,In_861,In_261);
and U46 (N_46,In_463,In_266);
nand U47 (N_47,In_418,In_553);
nor U48 (N_48,In_585,In_888);
nor U49 (N_49,In_533,In_211);
nor U50 (N_50,In_567,In_716);
and U51 (N_51,In_208,In_415);
or U52 (N_52,In_802,In_254);
or U53 (N_53,In_552,In_516);
xnor U54 (N_54,In_102,In_738);
and U55 (N_55,In_224,In_319);
and U56 (N_56,In_219,In_251);
or U57 (N_57,In_824,In_366);
and U58 (N_58,In_855,In_368);
or U59 (N_59,In_731,In_804);
nor U60 (N_60,In_527,In_594);
and U61 (N_61,In_365,In_332);
nand U62 (N_62,In_893,In_958);
and U63 (N_63,In_611,In_929);
or U64 (N_64,In_859,In_23);
and U65 (N_65,In_543,In_395);
or U66 (N_66,In_18,In_79);
or U67 (N_67,In_73,In_221);
and U68 (N_68,In_743,In_556);
nand U69 (N_69,In_617,In_708);
or U70 (N_70,In_581,In_727);
nand U71 (N_71,In_671,In_678);
nor U72 (N_72,In_806,In_480);
or U73 (N_73,In_414,In_59);
nand U74 (N_74,In_749,In_74);
or U75 (N_75,In_84,In_597);
or U76 (N_76,In_477,In_40);
or U77 (N_77,In_50,In_791);
nand U78 (N_78,In_287,In_538);
or U79 (N_79,In_184,In_260);
nor U80 (N_80,In_897,In_564);
nand U81 (N_81,In_448,In_603);
nand U82 (N_82,In_333,In_620);
nand U83 (N_83,In_111,In_163);
nor U84 (N_84,In_471,In_975);
nand U85 (N_85,In_93,In_881);
nor U86 (N_86,In_735,In_679);
nor U87 (N_87,In_705,In_863);
and U88 (N_88,In_807,In_230);
and U89 (N_89,In_255,In_622);
nand U90 (N_90,In_0,In_2);
and U91 (N_91,In_823,In_34);
nand U92 (N_92,In_346,In_615);
or U93 (N_93,In_762,In_940);
and U94 (N_94,In_944,In_412);
nand U95 (N_95,In_231,In_515);
nand U96 (N_96,In_288,In_793);
or U97 (N_97,In_675,In_752);
nor U98 (N_98,In_795,In_798);
and U99 (N_99,In_374,In_834);
or U100 (N_100,In_481,In_833);
nor U101 (N_101,In_417,In_542);
nor U102 (N_102,In_618,In_956);
and U103 (N_103,In_596,In_870);
and U104 (N_104,In_638,In_867);
nand U105 (N_105,In_754,In_430);
nand U106 (N_106,In_454,In_15);
and U107 (N_107,In_22,In_460);
or U108 (N_108,In_691,In_822);
nand U109 (N_109,In_755,In_548);
and U110 (N_110,In_587,In_892);
or U111 (N_111,In_391,In_46);
nand U112 (N_112,In_229,In_433);
and U113 (N_113,In_693,In_397);
nor U114 (N_114,In_715,In_610);
nor U115 (N_115,In_498,In_924);
nand U116 (N_116,In_598,In_936);
nor U117 (N_117,In_92,In_264);
nand U118 (N_118,In_279,In_961);
or U119 (N_119,In_812,In_817);
and U120 (N_120,In_786,In_774);
and U121 (N_121,In_392,In_189);
or U122 (N_122,In_435,In_164);
and U123 (N_123,In_509,In_563);
and U124 (N_124,In_972,In_31);
nand U125 (N_125,In_697,In_803);
nor U126 (N_126,In_898,In_354);
xnor U127 (N_127,In_513,In_416);
nand U128 (N_128,In_681,In_797);
nand U129 (N_129,In_730,In_476);
nand U130 (N_130,In_937,In_64);
nand U131 (N_131,In_196,In_760);
or U132 (N_132,In_289,In_351);
and U133 (N_133,In_497,In_580);
nand U134 (N_134,In_555,In_966);
nor U135 (N_135,In_151,In_65);
nand U136 (N_136,In_641,In_869);
xnor U137 (N_137,In_880,In_85);
and U138 (N_138,In_914,In_437);
and U139 (N_139,In_896,In_571);
nor U140 (N_140,In_714,In_69);
or U141 (N_141,In_525,In_987);
nand U142 (N_142,In_505,In_129);
nand U143 (N_143,In_328,In_792);
or U144 (N_144,In_209,In_135);
and U145 (N_145,In_474,In_42);
or U146 (N_146,In_917,In_665);
or U147 (N_147,In_378,In_876);
nor U148 (N_148,In_205,In_335);
nand U149 (N_149,In_218,In_413);
or U150 (N_150,In_996,In_244);
or U151 (N_151,In_889,In_48);
nand U152 (N_152,In_763,In_44);
nor U153 (N_153,In_5,In_600);
or U154 (N_154,In_348,In_370);
nand U155 (N_155,In_971,In_311);
nand U156 (N_156,In_297,In_796);
nor U157 (N_157,In_267,In_947);
nand U158 (N_158,In_80,In_964);
nor U159 (N_159,In_901,In_979);
nor U160 (N_160,In_994,In_165);
nand U161 (N_161,In_490,In_713);
or U162 (N_162,In_106,In_560);
or U163 (N_163,In_801,In_166);
or U164 (N_164,In_589,In_965);
or U165 (N_165,In_91,In_295);
and U166 (N_166,In_313,In_225);
nor U167 (N_167,In_158,In_988);
or U168 (N_168,In_811,In_161);
and U169 (N_169,In_293,In_153);
and U170 (N_170,In_90,In_843);
nand U171 (N_171,In_359,In_247);
nand U172 (N_172,In_920,In_182);
or U173 (N_173,In_957,In_103);
nor U174 (N_174,In_724,In_449);
nand U175 (N_175,In_739,In_464);
nand U176 (N_176,In_86,In_900);
nor U177 (N_177,In_946,In_942);
nor U178 (N_178,In_711,In_499);
xor U179 (N_179,In_761,In_857);
nand U180 (N_180,In_656,In_292);
xnor U181 (N_181,In_787,In_4);
nand U182 (N_182,In_922,In_701);
nor U183 (N_183,In_586,In_660);
nand U184 (N_184,In_253,In_546);
and U185 (N_185,In_410,In_210);
nor U186 (N_186,In_409,In_506);
nand U187 (N_187,In_959,In_466);
and U188 (N_188,In_853,In_672);
and U189 (N_189,In_736,In_604);
or U190 (N_190,In_142,In_127);
nor U191 (N_191,In_30,In_104);
or U192 (N_192,In_841,In_578);
or U193 (N_193,In_240,In_149);
and U194 (N_194,In_223,In_646);
nor U195 (N_195,In_173,In_338);
and U196 (N_196,In_951,In_123);
nor U197 (N_197,In_758,In_751);
or U198 (N_198,In_457,In_561);
nand U199 (N_199,In_518,In_281);
nand U200 (N_200,In_388,In_118);
and U201 (N_201,In_753,In_20);
nor U202 (N_202,In_57,In_503);
nor U203 (N_203,In_180,In_14);
nand U204 (N_204,In_875,In_915);
or U205 (N_205,In_155,In_584);
and U206 (N_206,In_306,In_634);
and U207 (N_207,In_698,In_312);
and U208 (N_208,In_54,In_745);
xnor U209 (N_209,In_726,In_851);
and U210 (N_210,In_334,In_285);
nand U211 (N_211,In_318,In_636);
nand U212 (N_212,In_568,In_327);
nand U213 (N_213,In_496,In_349);
or U214 (N_214,In_818,In_242);
or U215 (N_215,In_950,In_355);
nor U216 (N_216,In_902,In_24);
nand U217 (N_217,In_616,In_912);
and U218 (N_218,In_26,In_539);
and U219 (N_219,In_188,In_226);
or U220 (N_220,In_262,In_228);
nand U221 (N_221,In_592,In_114);
nor U222 (N_222,In_258,In_702);
nor U223 (N_223,In_444,In_868);
nor U224 (N_224,In_765,In_904);
nand U225 (N_225,In_394,In_411);
nor U226 (N_226,In_704,In_268);
or U227 (N_227,In_955,In_174);
nor U228 (N_228,In_233,In_286);
or U229 (N_229,In_150,In_559);
and U230 (N_230,In_642,In_878);
nor U231 (N_231,In_528,In_245);
nor U232 (N_232,In_582,In_94);
nand U233 (N_233,In_81,In_814);
and U234 (N_234,In_913,In_908);
and U235 (N_235,In_991,In_742);
nand U236 (N_236,In_146,In_510);
xor U237 (N_237,In_58,In_393);
nor U238 (N_238,In_329,In_381);
nand U239 (N_239,In_300,In_298);
nor U240 (N_240,In_750,In_273);
nand U241 (N_241,In_99,In_952);
or U242 (N_242,In_570,In_487);
nand U243 (N_243,In_256,In_687);
nor U244 (N_244,In_199,In_140);
nor U245 (N_245,In_154,In_272);
nor U246 (N_246,In_989,In_183);
nand U247 (N_247,In_484,In_640);
and U248 (N_248,In_246,In_217);
and U249 (N_249,In_116,In_204);
nor U250 (N_250,In_326,In_643);
xor U251 (N_251,In_45,In_688);
nor U252 (N_252,In_984,In_769);
nor U253 (N_253,In_402,In_839);
nand U254 (N_254,In_88,In_718);
or U255 (N_255,In_363,In_921);
and U256 (N_256,In_446,In_631);
or U257 (N_257,In_894,In_171);
nor U258 (N_258,In_108,In_832);
and U259 (N_259,In_554,In_494);
and U260 (N_260,In_593,In_722);
or U261 (N_261,In_635,In_197);
and U262 (N_262,In_847,In_304);
and U263 (N_263,In_690,In_632);
nand U264 (N_264,In_998,In_16);
nand U265 (N_265,In_982,In_213);
nor U266 (N_266,In_458,In_707);
nand U267 (N_267,In_485,In_37);
nand U268 (N_268,In_540,In_170);
and U269 (N_269,In_933,In_263);
nand U270 (N_270,In_980,In_865);
nand U271 (N_271,In_895,In_777);
nor U272 (N_272,In_265,In_408);
nand U273 (N_273,In_575,In_17);
nor U274 (N_274,In_639,In_339);
nand U275 (N_275,In_113,In_993);
nand U276 (N_276,In_932,In_82);
or U277 (N_277,In_456,In_323);
nor U278 (N_278,In_523,In_19);
or U279 (N_279,In_423,In_479);
nor U280 (N_280,In_455,In_668);
and U281 (N_281,In_269,In_931);
nand U282 (N_282,In_978,In_280);
nand U283 (N_283,In_800,In_759);
or U284 (N_284,In_187,In_907);
and U285 (N_285,In_500,In_923);
nand U286 (N_286,In_808,In_77);
nand U287 (N_287,In_181,In_473);
nand U288 (N_288,In_949,In_345);
nand U289 (N_289,In_826,In_562);
nor U290 (N_290,In_438,In_203);
nor U291 (N_291,In_566,In_100);
nand U292 (N_292,In_885,In_72);
or U293 (N_293,In_470,In_459);
nor U294 (N_294,In_502,In_41);
xor U295 (N_295,In_819,In_630);
and U296 (N_296,In_176,In_11);
or U297 (N_297,In_999,In_440);
nor U298 (N_298,In_519,In_551);
or U299 (N_299,In_399,In_633);
and U300 (N_300,In_919,In_78);
nand U301 (N_301,In_212,In_274);
or U302 (N_302,In_465,In_706);
and U303 (N_303,In_145,In_771);
and U304 (N_304,In_756,In_325);
or U305 (N_305,In_126,In_935);
or U306 (N_306,In_770,In_725);
and U307 (N_307,In_28,In_846);
or U308 (N_308,In_372,In_89);
or U309 (N_309,In_776,In_766);
nor U310 (N_310,In_501,In_772);
and U311 (N_311,In_827,In_864);
or U312 (N_312,In_493,In_719);
nor U313 (N_313,In_652,In_330);
xnor U314 (N_314,In_873,In_721);
nand U315 (N_315,In_669,In_547);
and U316 (N_316,In_775,In_741);
nand U317 (N_317,In_821,In_340);
nor U318 (N_318,In_162,In_76);
nor U319 (N_319,In_122,In_773);
and U320 (N_320,In_96,In_429);
nor U321 (N_321,In_524,In_884);
nand U322 (N_322,In_530,In_406);
nand U323 (N_323,In_469,In_653);
nand U324 (N_324,In_960,In_572);
or U325 (N_325,In_696,In_709);
and U326 (N_326,In_216,In_790);
nand U327 (N_327,In_605,In_549);
nand U328 (N_328,In_673,In_647);
nor U329 (N_329,In_109,In_717);
nor U330 (N_330,In_70,In_201);
and U331 (N_331,In_341,In_781);
nand U332 (N_332,In_905,In_789);
nand U333 (N_333,In_71,In_405);
nor U334 (N_334,In_39,In_746);
nand U335 (N_335,In_331,In_357);
nand U336 (N_336,In_152,In_627);
and U337 (N_337,In_238,In_29);
or U338 (N_338,In_443,In_852);
nand U339 (N_339,In_710,In_358);
and U340 (N_340,In_764,In_157);
and U341 (N_341,In_813,In_963);
or U342 (N_342,In_550,In_504);
or U343 (N_343,In_175,In_899);
nor U344 (N_344,In_712,In_360);
nor U345 (N_345,In_10,In_347);
and U346 (N_346,In_32,In_747);
or U347 (N_347,In_8,In_95);
or U348 (N_348,In_371,In_384);
and U349 (N_349,In_910,In_667);
nor U350 (N_350,In_650,In_396);
nand U351 (N_351,In_930,In_436);
or U352 (N_352,In_419,In_684);
nor U353 (N_353,In_661,In_387);
nand U354 (N_354,In_737,In_535);
nand U355 (N_355,In_829,In_202);
or U356 (N_356,In_545,In_651);
nand U357 (N_357,In_220,In_434);
nand U358 (N_358,In_427,In_788);
or U359 (N_359,In_119,In_682);
and U360 (N_360,In_740,In_657);
nand U361 (N_361,In_124,In_373);
nand U362 (N_362,In_591,In_239);
nor U363 (N_363,In_782,In_850);
or U364 (N_364,In_467,In_249);
nand U365 (N_365,In_301,In_21);
nor U366 (N_366,In_649,In_837);
and U367 (N_367,In_299,In_315);
and U368 (N_368,In_830,In_531);
xnor U369 (N_369,In_574,In_733);
or U370 (N_370,In_400,In_190);
nor U371 (N_371,In_780,In_324);
nor U372 (N_372,In_489,In_871);
or U373 (N_373,In_398,In_385);
nor U374 (N_374,In_541,In_43);
or U375 (N_375,In_602,In_337);
nand U376 (N_376,In_51,In_906);
or U377 (N_377,In_259,In_310);
xor U378 (N_378,In_840,In_447);
and U379 (N_379,In_317,In_67);
or U380 (N_380,In_167,In_138);
nand U381 (N_381,In_976,In_623);
or U382 (N_382,In_744,In_445);
and U383 (N_383,In_512,In_407);
nor U384 (N_384,In_53,In_87);
nand U385 (N_385,In_608,In_526);
nand U386 (N_386,In_590,In_488);
nor U387 (N_387,In_757,In_799);
or U388 (N_388,In_35,In_257);
or U389 (N_389,In_132,In_60);
nor U390 (N_390,In_7,In_831);
nand U391 (N_391,In_107,In_844);
or U392 (N_392,In_291,In_810);
or U393 (N_393,In_441,In_316);
nand U394 (N_394,In_674,In_13);
and U395 (N_395,In_784,In_537);
or U396 (N_396,In_520,In_320);
nor U397 (N_397,In_101,In_362);
and U398 (N_398,In_144,In_115);
or U399 (N_399,In_141,In_886);
nor U400 (N_400,In_336,In_663);
or U401 (N_401,In_364,In_179);
nor U402 (N_402,In_626,In_296);
nand U403 (N_403,In_49,In_483);
and U404 (N_404,In_284,In_612);
nor U405 (N_405,In_270,In_38);
or U406 (N_406,In_376,In_854);
or U407 (N_407,In_918,In_353);
nor U408 (N_408,In_521,In_990);
nor U409 (N_409,In_628,In_637);
nand U410 (N_410,In_685,In_856);
and U411 (N_411,In_125,In_985);
nor U412 (N_412,In_97,In_986);
and U413 (N_413,In_403,In_431);
nand U414 (N_414,In_768,In_883);
nor U415 (N_415,In_380,In_198);
and U416 (N_416,In_517,In_629);
nor U417 (N_417,In_664,In_579);
nor U418 (N_418,In_302,In_599);
or U419 (N_419,In_83,In_172);
and U420 (N_420,In_450,In_243);
nand U421 (N_421,In_835,In_420);
or U422 (N_422,In_723,In_820);
nand U423 (N_423,In_858,In_252);
nor U424 (N_424,In_683,In_981);
or U425 (N_425,In_432,In_421);
nor U426 (N_426,In_992,In_468);
or U427 (N_427,In_595,In_105);
or U428 (N_428,In_214,In_995);
or U429 (N_429,In_271,In_66);
nand U430 (N_430,In_734,In_472);
nand U431 (N_431,In_508,In_112);
or U432 (N_432,In_352,In_344);
nand U433 (N_433,In_968,In_282);
nand U434 (N_434,In_404,In_767);
nand U435 (N_435,In_577,In_241);
or U436 (N_436,In_156,In_903);
nor U437 (N_437,In_215,In_342);
nand U438 (N_438,In_928,In_177);
or U439 (N_439,In_322,In_495);
nor U440 (N_440,In_614,In_25);
nand U441 (N_441,In_695,In_872);
or U442 (N_442,In_439,In_644);
nor U443 (N_443,In_882,In_350);
and U444 (N_444,In_442,In_655);
nand U445 (N_445,In_475,In_534);
nand U446 (N_446,In_778,In_848);
nor U447 (N_447,In_207,In_461);
nand U448 (N_448,In_694,In_12);
and U449 (N_449,In_927,In_159);
nor U450 (N_450,In_390,In_308);
nand U451 (N_451,In_492,In_779);
nor U452 (N_452,In_478,In_816);
nor U453 (N_453,In_785,In_193);
nand U454 (N_454,In_248,In_662);
nor U455 (N_455,In_997,In_573);
nor U456 (N_456,In_120,In_462);
xnor U457 (N_457,In_576,In_139);
nor U458 (N_458,In_874,In_147);
nand U459 (N_459,In_624,In_130);
and U460 (N_460,In_136,In_536);
nor U461 (N_461,In_729,In_703);
and U462 (N_462,In_294,In_186);
and U463 (N_463,In_583,In_983);
or U464 (N_464,In_728,In_659);
nor U465 (N_465,In_860,In_283);
nor U466 (N_466,In_185,In_836);
and U467 (N_467,In_969,In_133);
or U468 (N_468,In_815,In_137);
or U469 (N_469,In_47,In_973);
or U470 (N_470,In_235,In_849);
and U471 (N_471,In_911,In_303);
nor U472 (N_472,In_828,In_532);
nor U473 (N_473,In_890,In_367);
nand U474 (N_474,In_169,In_686);
xnor U475 (N_475,In_941,In_645);
nand U476 (N_476,In_36,In_648);
nor U477 (N_477,In_110,In_389);
and U478 (N_478,In_27,In_75);
nand U479 (N_479,In_529,In_191);
or U480 (N_480,In_56,In_925);
or U481 (N_481,In_613,In_131);
nand U482 (N_482,In_232,In_486);
nor U483 (N_483,In_98,In_382);
nor U484 (N_484,In_670,In_680);
nand U485 (N_485,In_916,In_948);
xor U486 (N_486,In_61,In_68);
or U487 (N_487,In_809,In_148);
and U488 (N_488,In_977,In_974);
and U489 (N_489,In_943,In_970);
nand U490 (N_490,In_401,In_375);
nand U491 (N_491,In_625,In_236);
and U492 (N_492,In_278,In_654);
nor U493 (N_493,In_250,In_143);
and U494 (N_494,In_234,In_195);
nand U495 (N_495,In_361,In_383);
or U496 (N_496,In_609,In_192);
or U497 (N_497,In_666,In_945);
nor U498 (N_498,In_377,In_425);
nand U499 (N_499,In_6,In_938);
and U500 (N_500,In_459,In_47);
nor U501 (N_501,In_154,In_114);
nand U502 (N_502,In_839,In_834);
or U503 (N_503,In_963,In_907);
or U504 (N_504,In_980,In_341);
nand U505 (N_505,In_491,In_663);
and U506 (N_506,In_872,In_647);
nor U507 (N_507,In_69,In_163);
and U508 (N_508,In_307,In_138);
nor U509 (N_509,In_995,In_649);
or U510 (N_510,In_725,In_704);
nand U511 (N_511,In_696,In_214);
nand U512 (N_512,In_639,In_99);
nand U513 (N_513,In_260,In_673);
or U514 (N_514,In_128,In_189);
and U515 (N_515,In_502,In_609);
nand U516 (N_516,In_992,In_78);
and U517 (N_517,In_508,In_501);
and U518 (N_518,In_75,In_451);
or U519 (N_519,In_237,In_612);
and U520 (N_520,In_584,In_303);
nor U521 (N_521,In_599,In_936);
and U522 (N_522,In_899,In_433);
nor U523 (N_523,In_909,In_536);
or U524 (N_524,In_543,In_758);
or U525 (N_525,In_730,In_872);
or U526 (N_526,In_275,In_906);
nand U527 (N_527,In_885,In_237);
or U528 (N_528,In_177,In_111);
nor U529 (N_529,In_773,In_755);
and U530 (N_530,In_407,In_215);
nor U531 (N_531,In_474,In_812);
and U532 (N_532,In_657,In_15);
nor U533 (N_533,In_259,In_600);
nand U534 (N_534,In_352,In_615);
or U535 (N_535,In_975,In_428);
nand U536 (N_536,In_734,In_271);
nand U537 (N_537,In_214,In_177);
and U538 (N_538,In_411,In_634);
and U539 (N_539,In_478,In_170);
and U540 (N_540,In_655,In_276);
nor U541 (N_541,In_769,In_189);
and U542 (N_542,In_839,In_435);
or U543 (N_543,In_352,In_508);
or U544 (N_544,In_873,In_681);
and U545 (N_545,In_131,In_72);
or U546 (N_546,In_715,In_342);
nor U547 (N_547,In_234,In_917);
and U548 (N_548,In_167,In_68);
nor U549 (N_549,In_30,In_374);
nand U550 (N_550,In_584,In_341);
nor U551 (N_551,In_852,In_111);
or U552 (N_552,In_846,In_400);
nor U553 (N_553,In_791,In_249);
nor U554 (N_554,In_896,In_838);
and U555 (N_555,In_27,In_386);
nand U556 (N_556,In_5,In_404);
and U557 (N_557,In_634,In_958);
nor U558 (N_558,In_328,In_734);
nand U559 (N_559,In_731,In_137);
or U560 (N_560,In_413,In_873);
and U561 (N_561,In_9,In_637);
nand U562 (N_562,In_393,In_713);
nor U563 (N_563,In_986,In_985);
nand U564 (N_564,In_535,In_179);
and U565 (N_565,In_132,In_81);
and U566 (N_566,In_222,In_949);
nor U567 (N_567,In_609,In_151);
nand U568 (N_568,In_190,In_9);
nand U569 (N_569,In_801,In_321);
nor U570 (N_570,In_791,In_459);
or U571 (N_571,In_586,In_37);
and U572 (N_572,In_899,In_851);
nand U573 (N_573,In_64,In_52);
nand U574 (N_574,In_641,In_944);
or U575 (N_575,In_255,In_594);
nand U576 (N_576,In_121,In_53);
and U577 (N_577,In_51,In_552);
nor U578 (N_578,In_530,In_169);
nand U579 (N_579,In_918,In_334);
and U580 (N_580,In_952,In_325);
and U581 (N_581,In_878,In_621);
nor U582 (N_582,In_469,In_348);
and U583 (N_583,In_223,In_300);
nand U584 (N_584,In_930,In_686);
and U585 (N_585,In_982,In_825);
or U586 (N_586,In_404,In_667);
or U587 (N_587,In_923,In_72);
nor U588 (N_588,In_168,In_537);
or U589 (N_589,In_521,In_34);
nor U590 (N_590,In_628,In_662);
or U591 (N_591,In_477,In_20);
nor U592 (N_592,In_747,In_708);
or U593 (N_593,In_616,In_208);
and U594 (N_594,In_953,In_580);
or U595 (N_595,In_949,In_61);
nand U596 (N_596,In_982,In_631);
nand U597 (N_597,In_923,In_650);
and U598 (N_598,In_746,In_547);
or U599 (N_599,In_179,In_173);
nand U600 (N_600,In_187,In_500);
nor U601 (N_601,In_513,In_407);
nand U602 (N_602,In_434,In_450);
or U603 (N_603,In_446,In_86);
xnor U604 (N_604,In_361,In_437);
and U605 (N_605,In_275,In_60);
and U606 (N_606,In_523,In_839);
and U607 (N_607,In_236,In_849);
nor U608 (N_608,In_353,In_435);
and U609 (N_609,In_941,In_923);
nor U610 (N_610,In_596,In_937);
and U611 (N_611,In_609,In_714);
and U612 (N_612,In_726,In_410);
or U613 (N_613,In_865,In_618);
or U614 (N_614,In_491,In_969);
and U615 (N_615,In_661,In_116);
and U616 (N_616,In_272,In_373);
nor U617 (N_617,In_598,In_96);
or U618 (N_618,In_913,In_866);
or U619 (N_619,In_867,In_864);
and U620 (N_620,In_405,In_636);
nor U621 (N_621,In_946,In_294);
nor U622 (N_622,In_139,In_523);
nand U623 (N_623,In_848,In_158);
or U624 (N_624,In_80,In_114);
nand U625 (N_625,In_739,In_10);
and U626 (N_626,In_964,In_965);
or U627 (N_627,In_767,In_492);
and U628 (N_628,In_899,In_44);
or U629 (N_629,In_199,In_485);
or U630 (N_630,In_88,In_776);
and U631 (N_631,In_61,In_529);
nor U632 (N_632,In_808,In_7);
nor U633 (N_633,In_925,In_112);
nor U634 (N_634,In_943,In_738);
nand U635 (N_635,In_802,In_902);
and U636 (N_636,In_933,In_299);
or U637 (N_637,In_734,In_90);
or U638 (N_638,In_858,In_141);
nor U639 (N_639,In_144,In_459);
nor U640 (N_640,In_553,In_589);
nor U641 (N_641,In_204,In_945);
xor U642 (N_642,In_159,In_26);
nand U643 (N_643,In_14,In_419);
nand U644 (N_644,In_370,In_520);
or U645 (N_645,In_540,In_628);
and U646 (N_646,In_5,In_818);
nand U647 (N_647,In_372,In_234);
and U648 (N_648,In_304,In_610);
and U649 (N_649,In_57,In_579);
or U650 (N_650,In_968,In_127);
or U651 (N_651,In_768,In_20);
or U652 (N_652,In_536,In_273);
nand U653 (N_653,In_463,In_219);
and U654 (N_654,In_705,In_134);
nor U655 (N_655,In_754,In_520);
nand U656 (N_656,In_454,In_645);
nor U657 (N_657,In_450,In_940);
nor U658 (N_658,In_344,In_911);
or U659 (N_659,In_920,In_939);
and U660 (N_660,In_763,In_995);
or U661 (N_661,In_90,In_760);
nor U662 (N_662,In_968,In_818);
nor U663 (N_663,In_858,In_293);
nand U664 (N_664,In_63,In_48);
or U665 (N_665,In_561,In_918);
and U666 (N_666,In_518,In_728);
nor U667 (N_667,In_900,In_443);
and U668 (N_668,In_313,In_211);
and U669 (N_669,In_490,In_416);
or U670 (N_670,In_273,In_421);
nand U671 (N_671,In_103,In_890);
and U672 (N_672,In_504,In_334);
nand U673 (N_673,In_920,In_306);
and U674 (N_674,In_808,In_938);
nand U675 (N_675,In_541,In_928);
nor U676 (N_676,In_152,In_380);
and U677 (N_677,In_263,In_5);
or U678 (N_678,In_452,In_434);
or U679 (N_679,In_749,In_989);
xor U680 (N_680,In_387,In_551);
nand U681 (N_681,In_429,In_22);
or U682 (N_682,In_453,In_310);
and U683 (N_683,In_12,In_526);
nor U684 (N_684,In_647,In_490);
nand U685 (N_685,In_958,In_33);
nor U686 (N_686,In_553,In_327);
nand U687 (N_687,In_914,In_1);
or U688 (N_688,In_812,In_18);
nor U689 (N_689,In_90,In_459);
and U690 (N_690,In_399,In_250);
nor U691 (N_691,In_847,In_456);
nor U692 (N_692,In_209,In_935);
nor U693 (N_693,In_747,In_166);
and U694 (N_694,In_136,In_241);
and U695 (N_695,In_781,In_29);
nor U696 (N_696,In_519,In_440);
nand U697 (N_697,In_26,In_773);
nand U698 (N_698,In_816,In_228);
nor U699 (N_699,In_663,In_138);
nand U700 (N_700,In_660,In_88);
or U701 (N_701,In_5,In_357);
or U702 (N_702,In_612,In_887);
and U703 (N_703,In_218,In_124);
xnor U704 (N_704,In_133,In_587);
nor U705 (N_705,In_695,In_63);
nand U706 (N_706,In_366,In_220);
nor U707 (N_707,In_546,In_12);
nor U708 (N_708,In_786,In_346);
nor U709 (N_709,In_368,In_802);
nand U710 (N_710,In_738,In_882);
nand U711 (N_711,In_945,In_671);
or U712 (N_712,In_159,In_779);
nand U713 (N_713,In_157,In_797);
nor U714 (N_714,In_207,In_264);
or U715 (N_715,In_991,In_586);
and U716 (N_716,In_739,In_22);
nor U717 (N_717,In_432,In_346);
and U718 (N_718,In_630,In_948);
nor U719 (N_719,In_896,In_931);
and U720 (N_720,In_815,In_656);
and U721 (N_721,In_917,In_278);
nor U722 (N_722,In_998,In_753);
nand U723 (N_723,In_304,In_33);
and U724 (N_724,In_963,In_339);
or U725 (N_725,In_757,In_811);
and U726 (N_726,In_59,In_943);
nand U727 (N_727,In_659,In_158);
or U728 (N_728,In_711,In_291);
nor U729 (N_729,In_569,In_407);
and U730 (N_730,In_73,In_754);
nand U731 (N_731,In_572,In_295);
and U732 (N_732,In_901,In_9);
or U733 (N_733,In_890,In_898);
nand U734 (N_734,In_740,In_618);
and U735 (N_735,In_139,In_934);
or U736 (N_736,In_916,In_295);
or U737 (N_737,In_234,In_491);
nor U738 (N_738,In_184,In_160);
nor U739 (N_739,In_666,In_53);
nand U740 (N_740,In_61,In_996);
or U741 (N_741,In_445,In_599);
nor U742 (N_742,In_153,In_85);
and U743 (N_743,In_862,In_456);
nand U744 (N_744,In_871,In_71);
nand U745 (N_745,In_965,In_257);
nor U746 (N_746,In_570,In_843);
nor U747 (N_747,In_460,In_329);
nand U748 (N_748,In_642,In_746);
or U749 (N_749,In_514,In_576);
or U750 (N_750,In_381,In_341);
and U751 (N_751,In_35,In_641);
and U752 (N_752,In_277,In_1);
nand U753 (N_753,In_510,In_145);
and U754 (N_754,In_953,In_438);
nor U755 (N_755,In_959,In_747);
nand U756 (N_756,In_923,In_75);
nand U757 (N_757,In_996,In_960);
nand U758 (N_758,In_26,In_847);
and U759 (N_759,In_164,In_361);
nand U760 (N_760,In_157,In_99);
and U761 (N_761,In_506,In_970);
or U762 (N_762,In_468,In_639);
nor U763 (N_763,In_959,In_207);
nand U764 (N_764,In_989,In_401);
and U765 (N_765,In_273,In_610);
nor U766 (N_766,In_485,In_656);
or U767 (N_767,In_486,In_789);
or U768 (N_768,In_317,In_673);
nor U769 (N_769,In_27,In_467);
nand U770 (N_770,In_567,In_601);
nor U771 (N_771,In_598,In_819);
nor U772 (N_772,In_841,In_41);
and U773 (N_773,In_500,In_713);
nor U774 (N_774,In_626,In_56);
nand U775 (N_775,In_280,In_517);
or U776 (N_776,In_138,In_647);
or U777 (N_777,In_179,In_222);
nor U778 (N_778,In_55,In_152);
or U779 (N_779,In_909,In_292);
or U780 (N_780,In_542,In_309);
nor U781 (N_781,In_680,In_84);
nor U782 (N_782,In_955,In_801);
nand U783 (N_783,In_308,In_171);
nor U784 (N_784,In_54,In_506);
or U785 (N_785,In_396,In_643);
or U786 (N_786,In_766,In_704);
nor U787 (N_787,In_451,In_486);
nor U788 (N_788,In_147,In_986);
or U789 (N_789,In_101,In_79);
and U790 (N_790,In_772,In_742);
nand U791 (N_791,In_940,In_769);
nand U792 (N_792,In_493,In_964);
and U793 (N_793,In_314,In_330);
and U794 (N_794,In_690,In_628);
and U795 (N_795,In_121,In_598);
nand U796 (N_796,In_514,In_78);
and U797 (N_797,In_118,In_943);
xnor U798 (N_798,In_622,In_653);
nand U799 (N_799,In_198,In_118);
nor U800 (N_800,In_925,In_663);
and U801 (N_801,In_403,In_577);
nand U802 (N_802,In_841,In_759);
nand U803 (N_803,In_211,In_406);
and U804 (N_804,In_545,In_566);
or U805 (N_805,In_172,In_549);
and U806 (N_806,In_884,In_89);
nand U807 (N_807,In_71,In_767);
or U808 (N_808,In_775,In_215);
nand U809 (N_809,In_837,In_620);
and U810 (N_810,In_353,In_436);
nor U811 (N_811,In_688,In_189);
nor U812 (N_812,In_420,In_793);
or U813 (N_813,In_664,In_269);
xnor U814 (N_814,In_197,In_17);
nand U815 (N_815,In_46,In_217);
or U816 (N_816,In_980,In_302);
nand U817 (N_817,In_866,In_472);
nand U818 (N_818,In_205,In_29);
nor U819 (N_819,In_901,In_548);
nor U820 (N_820,In_697,In_646);
and U821 (N_821,In_561,In_84);
nand U822 (N_822,In_910,In_480);
nand U823 (N_823,In_438,In_397);
and U824 (N_824,In_929,In_340);
nor U825 (N_825,In_179,In_709);
nor U826 (N_826,In_358,In_820);
and U827 (N_827,In_359,In_169);
nor U828 (N_828,In_48,In_600);
and U829 (N_829,In_800,In_947);
and U830 (N_830,In_665,In_72);
nor U831 (N_831,In_150,In_852);
and U832 (N_832,In_761,In_70);
nand U833 (N_833,In_428,In_323);
or U834 (N_834,In_501,In_339);
and U835 (N_835,In_524,In_151);
nand U836 (N_836,In_730,In_204);
nand U837 (N_837,In_935,In_771);
and U838 (N_838,In_209,In_775);
or U839 (N_839,In_258,In_733);
nand U840 (N_840,In_949,In_834);
xnor U841 (N_841,In_141,In_372);
nand U842 (N_842,In_615,In_577);
nand U843 (N_843,In_303,In_73);
or U844 (N_844,In_238,In_455);
nand U845 (N_845,In_857,In_111);
nor U846 (N_846,In_946,In_517);
or U847 (N_847,In_297,In_267);
or U848 (N_848,In_850,In_112);
nand U849 (N_849,In_255,In_773);
or U850 (N_850,In_268,In_590);
nand U851 (N_851,In_418,In_978);
nor U852 (N_852,In_603,In_863);
nand U853 (N_853,In_56,In_698);
or U854 (N_854,In_815,In_771);
and U855 (N_855,In_70,In_558);
or U856 (N_856,In_944,In_982);
nand U857 (N_857,In_400,In_553);
and U858 (N_858,In_23,In_376);
nor U859 (N_859,In_169,In_923);
or U860 (N_860,In_781,In_953);
and U861 (N_861,In_900,In_742);
nand U862 (N_862,In_210,In_842);
and U863 (N_863,In_693,In_140);
nor U864 (N_864,In_906,In_119);
nand U865 (N_865,In_869,In_205);
nand U866 (N_866,In_256,In_924);
nor U867 (N_867,In_373,In_46);
nor U868 (N_868,In_479,In_292);
nand U869 (N_869,In_341,In_99);
or U870 (N_870,In_692,In_494);
nand U871 (N_871,In_976,In_109);
nand U872 (N_872,In_584,In_788);
and U873 (N_873,In_566,In_548);
and U874 (N_874,In_827,In_606);
or U875 (N_875,In_742,In_447);
or U876 (N_876,In_995,In_629);
nand U877 (N_877,In_763,In_141);
and U878 (N_878,In_122,In_426);
or U879 (N_879,In_578,In_242);
or U880 (N_880,In_825,In_452);
nor U881 (N_881,In_654,In_515);
and U882 (N_882,In_874,In_422);
or U883 (N_883,In_204,In_421);
or U884 (N_884,In_450,In_882);
or U885 (N_885,In_664,In_860);
nand U886 (N_886,In_355,In_204);
or U887 (N_887,In_492,In_65);
and U888 (N_888,In_996,In_148);
or U889 (N_889,In_920,In_898);
or U890 (N_890,In_818,In_47);
and U891 (N_891,In_681,In_168);
nor U892 (N_892,In_89,In_687);
and U893 (N_893,In_387,In_353);
and U894 (N_894,In_789,In_857);
nand U895 (N_895,In_140,In_700);
nand U896 (N_896,In_509,In_341);
xor U897 (N_897,In_225,In_567);
and U898 (N_898,In_243,In_737);
nor U899 (N_899,In_609,In_431);
nor U900 (N_900,In_659,In_95);
or U901 (N_901,In_697,In_85);
nand U902 (N_902,In_992,In_209);
or U903 (N_903,In_532,In_547);
nand U904 (N_904,In_526,In_674);
or U905 (N_905,In_638,In_349);
or U906 (N_906,In_424,In_516);
nand U907 (N_907,In_480,In_265);
nand U908 (N_908,In_581,In_32);
nor U909 (N_909,In_847,In_389);
and U910 (N_910,In_925,In_155);
nand U911 (N_911,In_343,In_452);
nand U912 (N_912,In_275,In_167);
nor U913 (N_913,In_496,In_390);
and U914 (N_914,In_69,In_683);
and U915 (N_915,In_851,In_580);
and U916 (N_916,In_880,In_275);
or U917 (N_917,In_849,In_997);
or U918 (N_918,In_464,In_126);
and U919 (N_919,In_559,In_88);
nand U920 (N_920,In_737,In_398);
and U921 (N_921,In_282,In_838);
nor U922 (N_922,In_980,In_596);
nor U923 (N_923,In_787,In_466);
nand U924 (N_924,In_422,In_750);
or U925 (N_925,In_397,In_798);
nand U926 (N_926,In_268,In_908);
or U927 (N_927,In_63,In_185);
or U928 (N_928,In_236,In_624);
or U929 (N_929,In_412,In_544);
and U930 (N_930,In_470,In_252);
nand U931 (N_931,In_367,In_972);
nand U932 (N_932,In_756,In_191);
nor U933 (N_933,In_219,In_268);
and U934 (N_934,In_710,In_206);
nor U935 (N_935,In_73,In_968);
and U936 (N_936,In_159,In_511);
and U937 (N_937,In_101,In_460);
or U938 (N_938,In_912,In_51);
or U939 (N_939,In_917,In_126);
nor U940 (N_940,In_811,In_24);
or U941 (N_941,In_560,In_352);
and U942 (N_942,In_721,In_748);
or U943 (N_943,In_113,In_428);
and U944 (N_944,In_504,In_255);
nand U945 (N_945,In_239,In_402);
nor U946 (N_946,In_283,In_67);
and U947 (N_947,In_268,In_650);
nor U948 (N_948,In_659,In_78);
or U949 (N_949,In_552,In_856);
and U950 (N_950,In_930,In_699);
nor U951 (N_951,In_394,In_732);
and U952 (N_952,In_199,In_562);
nor U953 (N_953,In_888,In_221);
nor U954 (N_954,In_42,In_863);
nand U955 (N_955,In_832,In_187);
or U956 (N_956,In_234,In_664);
and U957 (N_957,In_639,In_841);
and U958 (N_958,In_453,In_345);
nor U959 (N_959,In_910,In_112);
and U960 (N_960,In_526,In_346);
nand U961 (N_961,In_314,In_16);
or U962 (N_962,In_849,In_791);
nor U963 (N_963,In_687,In_799);
nand U964 (N_964,In_112,In_761);
nor U965 (N_965,In_511,In_508);
nor U966 (N_966,In_519,In_888);
nand U967 (N_967,In_199,In_877);
or U968 (N_968,In_221,In_532);
and U969 (N_969,In_513,In_633);
nand U970 (N_970,In_853,In_173);
xor U971 (N_971,In_187,In_29);
nand U972 (N_972,In_806,In_574);
nor U973 (N_973,In_283,In_322);
nor U974 (N_974,In_448,In_476);
nand U975 (N_975,In_426,In_215);
nor U976 (N_976,In_427,In_666);
or U977 (N_977,In_234,In_270);
or U978 (N_978,In_22,In_256);
nor U979 (N_979,In_302,In_508);
or U980 (N_980,In_642,In_838);
and U981 (N_981,In_987,In_721);
or U982 (N_982,In_581,In_946);
and U983 (N_983,In_552,In_536);
or U984 (N_984,In_842,In_116);
and U985 (N_985,In_604,In_130);
nand U986 (N_986,In_850,In_957);
nor U987 (N_987,In_251,In_406);
nor U988 (N_988,In_840,In_34);
and U989 (N_989,In_710,In_802);
and U990 (N_990,In_922,In_652);
xor U991 (N_991,In_962,In_202);
nand U992 (N_992,In_31,In_976);
nand U993 (N_993,In_182,In_133);
and U994 (N_994,In_293,In_974);
nand U995 (N_995,In_875,In_777);
or U996 (N_996,In_625,In_492);
or U997 (N_997,In_32,In_320);
nand U998 (N_998,In_714,In_936);
nor U999 (N_999,In_625,In_580);
or U1000 (N_1000,In_358,In_533);
and U1001 (N_1001,In_478,In_330);
and U1002 (N_1002,In_441,In_634);
nand U1003 (N_1003,In_520,In_140);
or U1004 (N_1004,In_206,In_979);
nor U1005 (N_1005,In_673,In_142);
nor U1006 (N_1006,In_921,In_839);
and U1007 (N_1007,In_373,In_337);
nor U1008 (N_1008,In_217,In_845);
or U1009 (N_1009,In_999,In_862);
nand U1010 (N_1010,In_339,In_265);
nand U1011 (N_1011,In_152,In_491);
and U1012 (N_1012,In_654,In_78);
and U1013 (N_1013,In_500,In_410);
nor U1014 (N_1014,In_928,In_874);
or U1015 (N_1015,In_661,In_375);
nor U1016 (N_1016,In_923,In_604);
and U1017 (N_1017,In_638,In_514);
or U1018 (N_1018,In_184,In_670);
and U1019 (N_1019,In_551,In_776);
nand U1020 (N_1020,In_106,In_469);
and U1021 (N_1021,In_542,In_383);
nand U1022 (N_1022,In_503,In_790);
or U1023 (N_1023,In_505,In_398);
nor U1024 (N_1024,In_502,In_993);
nand U1025 (N_1025,In_271,In_394);
nor U1026 (N_1026,In_453,In_516);
and U1027 (N_1027,In_459,In_190);
or U1028 (N_1028,In_389,In_162);
nand U1029 (N_1029,In_233,In_845);
nand U1030 (N_1030,In_611,In_843);
or U1031 (N_1031,In_164,In_687);
nor U1032 (N_1032,In_929,In_783);
nand U1033 (N_1033,In_854,In_631);
and U1034 (N_1034,In_987,In_776);
nor U1035 (N_1035,In_877,In_404);
nand U1036 (N_1036,In_320,In_729);
nand U1037 (N_1037,In_588,In_871);
or U1038 (N_1038,In_600,In_152);
and U1039 (N_1039,In_479,In_429);
or U1040 (N_1040,In_42,In_475);
nor U1041 (N_1041,In_583,In_986);
or U1042 (N_1042,In_570,In_424);
xnor U1043 (N_1043,In_824,In_368);
nand U1044 (N_1044,In_139,In_663);
or U1045 (N_1045,In_325,In_620);
and U1046 (N_1046,In_710,In_291);
nand U1047 (N_1047,In_689,In_939);
xor U1048 (N_1048,In_683,In_667);
and U1049 (N_1049,In_358,In_142);
or U1050 (N_1050,In_545,In_797);
or U1051 (N_1051,In_270,In_112);
nand U1052 (N_1052,In_39,In_604);
nor U1053 (N_1053,In_829,In_98);
nor U1054 (N_1054,In_82,In_449);
or U1055 (N_1055,In_637,In_689);
nor U1056 (N_1056,In_931,In_908);
nor U1057 (N_1057,In_550,In_145);
nor U1058 (N_1058,In_361,In_600);
or U1059 (N_1059,In_161,In_75);
nand U1060 (N_1060,In_500,In_85);
or U1061 (N_1061,In_431,In_61);
and U1062 (N_1062,In_628,In_671);
nand U1063 (N_1063,In_211,In_972);
and U1064 (N_1064,In_350,In_443);
nor U1065 (N_1065,In_594,In_419);
nand U1066 (N_1066,In_982,In_105);
nand U1067 (N_1067,In_850,In_587);
nand U1068 (N_1068,In_322,In_608);
or U1069 (N_1069,In_81,In_98);
and U1070 (N_1070,In_481,In_811);
and U1071 (N_1071,In_733,In_57);
nand U1072 (N_1072,In_745,In_257);
nand U1073 (N_1073,In_589,In_112);
and U1074 (N_1074,In_857,In_383);
nand U1075 (N_1075,In_307,In_934);
or U1076 (N_1076,In_545,In_658);
nor U1077 (N_1077,In_820,In_686);
and U1078 (N_1078,In_224,In_551);
nand U1079 (N_1079,In_795,In_550);
and U1080 (N_1080,In_858,In_789);
nand U1081 (N_1081,In_684,In_415);
nor U1082 (N_1082,In_875,In_618);
or U1083 (N_1083,In_551,In_825);
nor U1084 (N_1084,In_623,In_7);
nor U1085 (N_1085,In_63,In_801);
nor U1086 (N_1086,In_352,In_898);
nor U1087 (N_1087,In_183,In_80);
and U1088 (N_1088,In_964,In_890);
or U1089 (N_1089,In_656,In_653);
and U1090 (N_1090,In_412,In_171);
and U1091 (N_1091,In_671,In_717);
and U1092 (N_1092,In_498,In_394);
nand U1093 (N_1093,In_982,In_743);
nand U1094 (N_1094,In_120,In_371);
nand U1095 (N_1095,In_304,In_700);
and U1096 (N_1096,In_716,In_886);
nand U1097 (N_1097,In_825,In_745);
xor U1098 (N_1098,In_501,In_272);
or U1099 (N_1099,In_740,In_429);
nor U1100 (N_1100,In_56,In_640);
nor U1101 (N_1101,In_779,In_870);
and U1102 (N_1102,In_331,In_561);
or U1103 (N_1103,In_369,In_475);
nor U1104 (N_1104,In_968,In_641);
and U1105 (N_1105,In_593,In_224);
or U1106 (N_1106,In_830,In_457);
nand U1107 (N_1107,In_256,In_159);
or U1108 (N_1108,In_959,In_757);
nand U1109 (N_1109,In_464,In_696);
nand U1110 (N_1110,In_77,In_177);
nor U1111 (N_1111,In_531,In_960);
nor U1112 (N_1112,In_839,In_808);
and U1113 (N_1113,In_160,In_57);
nand U1114 (N_1114,In_366,In_610);
nand U1115 (N_1115,In_430,In_384);
or U1116 (N_1116,In_134,In_689);
nor U1117 (N_1117,In_338,In_157);
nand U1118 (N_1118,In_465,In_179);
nand U1119 (N_1119,In_862,In_444);
nand U1120 (N_1120,In_430,In_132);
nand U1121 (N_1121,In_942,In_271);
or U1122 (N_1122,In_956,In_204);
or U1123 (N_1123,In_922,In_486);
nor U1124 (N_1124,In_79,In_514);
nor U1125 (N_1125,In_4,In_256);
nor U1126 (N_1126,In_182,In_836);
or U1127 (N_1127,In_259,In_502);
or U1128 (N_1128,In_677,In_77);
nand U1129 (N_1129,In_153,In_934);
nor U1130 (N_1130,In_388,In_827);
or U1131 (N_1131,In_782,In_649);
or U1132 (N_1132,In_178,In_119);
or U1133 (N_1133,In_58,In_833);
and U1134 (N_1134,In_670,In_395);
and U1135 (N_1135,In_405,In_312);
nand U1136 (N_1136,In_21,In_921);
nand U1137 (N_1137,In_779,In_831);
or U1138 (N_1138,In_961,In_875);
or U1139 (N_1139,In_310,In_77);
nor U1140 (N_1140,In_464,In_474);
or U1141 (N_1141,In_490,In_94);
and U1142 (N_1142,In_222,In_157);
nand U1143 (N_1143,In_861,In_395);
or U1144 (N_1144,In_214,In_979);
or U1145 (N_1145,In_935,In_644);
nor U1146 (N_1146,In_369,In_929);
or U1147 (N_1147,In_986,In_293);
nand U1148 (N_1148,In_7,In_874);
xnor U1149 (N_1149,In_206,In_349);
and U1150 (N_1150,In_192,In_869);
or U1151 (N_1151,In_257,In_170);
or U1152 (N_1152,In_944,In_81);
or U1153 (N_1153,In_615,In_714);
nor U1154 (N_1154,In_759,In_812);
or U1155 (N_1155,In_12,In_818);
or U1156 (N_1156,In_988,In_930);
or U1157 (N_1157,In_571,In_244);
nand U1158 (N_1158,In_665,In_927);
or U1159 (N_1159,In_719,In_57);
and U1160 (N_1160,In_528,In_227);
nor U1161 (N_1161,In_179,In_166);
nand U1162 (N_1162,In_176,In_808);
and U1163 (N_1163,In_177,In_347);
nand U1164 (N_1164,In_803,In_449);
and U1165 (N_1165,In_229,In_497);
nor U1166 (N_1166,In_721,In_459);
or U1167 (N_1167,In_792,In_230);
nor U1168 (N_1168,In_65,In_585);
xor U1169 (N_1169,In_775,In_587);
and U1170 (N_1170,In_872,In_569);
and U1171 (N_1171,In_568,In_178);
nor U1172 (N_1172,In_353,In_860);
or U1173 (N_1173,In_904,In_331);
or U1174 (N_1174,In_158,In_755);
nor U1175 (N_1175,In_183,In_765);
or U1176 (N_1176,In_120,In_932);
xnor U1177 (N_1177,In_448,In_355);
nor U1178 (N_1178,In_614,In_430);
and U1179 (N_1179,In_897,In_185);
nand U1180 (N_1180,In_140,In_371);
nor U1181 (N_1181,In_202,In_838);
or U1182 (N_1182,In_894,In_667);
nand U1183 (N_1183,In_0,In_530);
and U1184 (N_1184,In_783,In_920);
and U1185 (N_1185,In_522,In_277);
nand U1186 (N_1186,In_617,In_502);
or U1187 (N_1187,In_667,In_709);
and U1188 (N_1188,In_56,In_736);
nand U1189 (N_1189,In_63,In_275);
nand U1190 (N_1190,In_19,In_390);
or U1191 (N_1191,In_812,In_365);
nor U1192 (N_1192,In_373,In_93);
and U1193 (N_1193,In_296,In_946);
or U1194 (N_1194,In_479,In_409);
nand U1195 (N_1195,In_402,In_865);
or U1196 (N_1196,In_252,In_856);
or U1197 (N_1197,In_410,In_260);
nor U1198 (N_1198,In_348,In_579);
and U1199 (N_1199,In_863,In_124);
nand U1200 (N_1200,In_16,In_199);
nor U1201 (N_1201,In_810,In_751);
or U1202 (N_1202,In_312,In_354);
or U1203 (N_1203,In_515,In_445);
or U1204 (N_1204,In_474,In_855);
and U1205 (N_1205,In_553,In_41);
or U1206 (N_1206,In_364,In_953);
nand U1207 (N_1207,In_765,In_172);
and U1208 (N_1208,In_8,In_632);
nor U1209 (N_1209,In_250,In_483);
or U1210 (N_1210,In_864,In_229);
nand U1211 (N_1211,In_989,In_543);
and U1212 (N_1212,In_606,In_644);
nand U1213 (N_1213,In_839,In_352);
nand U1214 (N_1214,In_330,In_822);
and U1215 (N_1215,In_701,In_291);
nor U1216 (N_1216,In_846,In_786);
nand U1217 (N_1217,In_708,In_677);
nor U1218 (N_1218,In_617,In_550);
nor U1219 (N_1219,In_970,In_638);
nor U1220 (N_1220,In_768,In_95);
and U1221 (N_1221,In_986,In_513);
nand U1222 (N_1222,In_652,In_499);
and U1223 (N_1223,In_668,In_236);
nor U1224 (N_1224,In_247,In_449);
or U1225 (N_1225,In_80,In_694);
nor U1226 (N_1226,In_541,In_527);
and U1227 (N_1227,In_3,In_917);
nor U1228 (N_1228,In_909,In_459);
and U1229 (N_1229,In_755,In_737);
and U1230 (N_1230,In_450,In_963);
nor U1231 (N_1231,In_654,In_722);
and U1232 (N_1232,In_377,In_688);
nor U1233 (N_1233,In_261,In_829);
and U1234 (N_1234,In_958,In_257);
nand U1235 (N_1235,In_544,In_970);
or U1236 (N_1236,In_354,In_338);
nand U1237 (N_1237,In_22,In_955);
or U1238 (N_1238,In_144,In_428);
nor U1239 (N_1239,In_374,In_15);
and U1240 (N_1240,In_399,In_569);
or U1241 (N_1241,In_62,In_927);
nand U1242 (N_1242,In_415,In_876);
nand U1243 (N_1243,In_369,In_0);
nand U1244 (N_1244,In_125,In_956);
nor U1245 (N_1245,In_169,In_145);
or U1246 (N_1246,In_886,In_197);
nand U1247 (N_1247,In_885,In_697);
nand U1248 (N_1248,In_290,In_328);
or U1249 (N_1249,In_636,In_117);
nand U1250 (N_1250,In_194,In_108);
or U1251 (N_1251,In_420,In_126);
and U1252 (N_1252,In_136,In_394);
or U1253 (N_1253,In_565,In_69);
nor U1254 (N_1254,In_252,In_757);
or U1255 (N_1255,In_205,In_128);
and U1256 (N_1256,In_367,In_362);
nor U1257 (N_1257,In_480,In_451);
and U1258 (N_1258,In_301,In_611);
and U1259 (N_1259,In_870,In_727);
nand U1260 (N_1260,In_737,In_624);
or U1261 (N_1261,In_599,In_316);
nand U1262 (N_1262,In_631,In_494);
or U1263 (N_1263,In_195,In_423);
and U1264 (N_1264,In_769,In_576);
and U1265 (N_1265,In_591,In_657);
nand U1266 (N_1266,In_644,In_512);
nor U1267 (N_1267,In_543,In_762);
and U1268 (N_1268,In_785,In_714);
or U1269 (N_1269,In_609,In_85);
and U1270 (N_1270,In_90,In_447);
nand U1271 (N_1271,In_574,In_658);
nor U1272 (N_1272,In_816,In_539);
nor U1273 (N_1273,In_356,In_149);
nor U1274 (N_1274,In_965,In_521);
and U1275 (N_1275,In_806,In_887);
or U1276 (N_1276,In_26,In_954);
nor U1277 (N_1277,In_187,In_86);
nor U1278 (N_1278,In_517,In_738);
nor U1279 (N_1279,In_60,In_834);
and U1280 (N_1280,In_793,In_568);
or U1281 (N_1281,In_283,In_187);
or U1282 (N_1282,In_524,In_292);
nand U1283 (N_1283,In_108,In_861);
nor U1284 (N_1284,In_486,In_359);
and U1285 (N_1285,In_367,In_500);
and U1286 (N_1286,In_656,In_25);
or U1287 (N_1287,In_68,In_768);
or U1288 (N_1288,In_130,In_757);
nor U1289 (N_1289,In_844,In_683);
nand U1290 (N_1290,In_583,In_19);
nor U1291 (N_1291,In_321,In_956);
nand U1292 (N_1292,In_45,In_523);
or U1293 (N_1293,In_758,In_403);
or U1294 (N_1294,In_381,In_35);
or U1295 (N_1295,In_611,In_25);
and U1296 (N_1296,In_636,In_559);
and U1297 (N_1297,In_867,In_366);
or U1298 (N_1298,In_619,In_70);
or U1299 (N_1299,In_688,In_781);
nand U1300 (N_1300,In_554,In_435);
nor U1301 (N_1301,In_586,In_885);
nor U1302 (N_1302,In_494,In_922);
and U1303 (N_1303,In_600,In_203);
nand U1304 (N_1304,In_932,In_474);
and U1305 (N_1305,In_115,In_754);
nand U1306 (N_1306,In_132,In_915);
nor U1307 (N_1307,In_300,In_72);
nand U1308 (N_1308,In_381,In_945);
or U1309 (N_1309,In_710,In_848);
and U1310 (N_1310,In_818,In_962);
nand U1311 (N_1311,In_951,In_315);
nand U1312 (N_1312,In_896,In_774);
and U1313 (N_1313,In_493,In_206);
nor U1314 (N_1314,In_917,In_849);
or U1315 (N_1315,In_234,In_488);
and U1316 (N_1316,In_818,In_491);
nand U1317 (N_1317,In_428,In_971);
nand U1318 (N_1318,In_677,In_69);
or U1319 (N_1319,In_635,In_659);
nand U1320 (N_1320,In_108,In_246);
nor U1321 (N_1321,In_622,In_44);
and U1322 (N_1322,In_165,In_177);
nand U1323 (N_1323,In_928,In_276);
xor U1324 (N_1324,In_246,In_411);
nor U1325 (N_1325,In_166,In_79);
nor U1326 (N_1326,In_748,In_960);
nor U1327 (N_1327,In_594,In_829);
nor U1328 (N_1328,In_131,In_493);
nor U1329 (N_1329,In_208,In_222);
and U1330 (N_1330,In_345,In_381);
and U1331 (N_1331,In_666,In_925);
or U1332 (N_1332,In_955,In_36);
nor U1333 (N_1333,In_258,In_549);
nand U1334 (N_1334,In_765,In_252);
nor U1335 (N_1335,In_496,In_703);
nand U1336 (N_1336,In_174,In_489);
nor U1337 (N_1337,In_632,In_833);
and U1338 (N_1338,In_592,In_754);
nand U1339 (N_1339,In_563,In_811);
and U1340 (N_1340,In_91,In_426);
nand U1341 (N_1341,In_671,In_818);
or U1342 (N_1342,In_493,In_290);
nor U1343 (N_1343,In_335,In_680);
and U1344 (N_1344,In_370,In_151);
nand U1345 (N_1345,In_969,In_701);
nand U1346 (N_1346,In_345,In_336);
or U1347 (N_1347,In_752,In_586);
or U1348 (N_1348,In_798,In_482);
or U1349 (N_1349,In_513,In_847);
nor U1350 (N_1350,In_76,In_33);
and U1351 (N_1351,In_478,In_574);
nor U1352 (N_1352,In_223,In_804);
or U1353 (N_1353,In_234,In_94);
nor U1354 (N_1354,In_777,In_95);
and U1355 (N_1355,In_430,In_403);
nor U1356 (N_1356,In_546,In_919);
nor U1357 (N_1357,In_270,In_995);
and U1358 (N_1358,In_303,In_681);
and U1359 (N_1359,In_681,In_882);
and U1360 (N_1360,In_453,In_712);
nor U1361 (N_1361,In_97,In_782);
and U1362 (N_1362,In_491,In_328);
and U1363 (N_1363,In_467,In_429);
or U1364 (N_1364,In_508,In_5);
or U1365 (N_1365,In_522,In_540);
nand U1366 (N_1366,In_789,In_705);
nand U1367 (N_1367,In_846,In_501);
and U1368 (N_1368,In_386,In_134);
and U1369 (N_1369,In_869,In_918);
nor U1370 (N_1370,In_882,In_741);
and U1371 (N_1371,In_390,In_386);
nor U1372 (N_1372,In_578,In_298);
or U1373 (N_1373,In_75,In_800);
or U1374 (N_1374,In_800,In_904);
nor U1375 (N_1375,In_436,In_545);
nor U1376 (N_1376,In_288,In_951);
or U1377 (N_1377,In_136,In_852);
and U1378 (N_1378,In_232,In_639);
or U1379 (N_1379,In_759,In_774);
and U1380 (N_1380,In_100,In_182);
xnor U1381 (N_1381,In_544,In_360);
and U1382 (N_1382,In_969,In_820);
nor U1383 (N_1383,In_695,In_117);
and U1384 (N_1384,In_43,In_427);
nand U1385 (N_1385,In_730,In_848);
nor U1386 (N_1386,In_356,In_536);
nand U1387 (N_1387,In_69,In_168);
and U1388 (N_1388,In_787,In_441);
nand U1389 (N_1389,In_410,In_829);
nand U1390 (N_1390,In_417,In_864);
and U1391 (N_1391,In_321,In_25);
and U1392 (N_1392,In_239,In_484);
or U1393 (N_1393,In_2,In_966);
or U1394 (N_1394,In_186,In_652);
nand U1395 (N_1395,In_950,In_515);
nand U1396 (N_1396,In_23,In_200);
and U1397 (N_1397,In_901,In_475);
and U1398 (N_1398,In_861,In_539);
or U1399 (N_1399,In_853,In_357);
nand U1400 (N_1400,In_360,In_9);
or U1401 (N_1401,In_5,In_673);
and U1402 (N_1402,In_331,In_338);
nor U1403 (N_1403,In_449,In_273);
or U1404 (N_1404,In_323,In_553);
or U1405 (N_1405,In_480,In_351);
nor U1406 (N_1406,In_214,In_565);
nand U1407 (N_1407,In_903,In_714);
nor U1408 (N_1408,In_565,In_258);
nor U1409 (N_1409,In_416,In_3);
and U1410 (N_1410,In_155,In_243);
nand U1411 (N_1411,In_202,In_67);
and U1412 (N_1412,In_700,In_525);
nand U1413 (N_1413,In_501,In_316);
nor U1414 (N_1414,In_503,In_650);
nand U1415 (N_1415,In_311,In_628);
and U1416 (N_1416,In_269,In_48);
and U1417 (N_1417,In_898,In_295);
or U1418 (N_1418,In_960,In_650);
nand U1419 (N_1419,In_144,In_479);
nand U1420 (N_1420,In_276,In_704);
and U1421 (N_1421,In_294,In_150);
nand U1422 (N_1422,In_31,In_775);
and U1423 (N_1423,In_499,In_385);
nor U1424 (N_1424,In_845,In_343);
or U1425 (N_1425,In_891,In_351);
nand U1426 (N_1426,In_730,In_54);
or U1427 (N_1427,In_297,In_949);
xnor U1428 (N_1428,In_198,In_596);
nor U1429 (N_1429,In_864,In_651);
nor U1430 (N_1430,In_444,In_323);
nand U1431 (N_1431,In_53,In_725);
and U1432 (N_1432,In_734,In_119);
nor U1433 (N_1433,In_398,In_919);
nor U1434 (N_1434,In_229,In_761);
or U1435 (N_1435,In_126,In_684);
and U1436 (N_1436,In_445,In_497);
nor U1437 (N_1437,In_854,In_323);
or U1438 (N_1438,In_818,In_111);
and U1439 (N_1439,In_693,In_162);
nor U1440 (N_1440,In_465,In_607);
nor U1441 (N_1441,In_441,In_708);
and U1442 (N_1442,In_418,In_543);
or U1443 (N_1443,In_545,In_467);
nor U1444 (N_1444,In_181,In_392);
and U1445 (N_1445,In_354,In_31);
or U1446 (N_1446,In_105,In_108);
or U1447 (N_1447,In_18,In_870);
and U1448 (N_1448,In_553,In_741);
and U1449 (N_1449,In_733,In_899);
nand U1450 (N_1450,In_511,In_417);
nand U1451 (N_1451,In_414,In_647);
nor U1452 (N_1452,In_657,In_772);
and U1453 (N_1453,In_784,In_148);
and U1454 (N_1454,In_483,In_947);
nand U1455 (N_1455,In_551,In_982);
nor U1456 (N_1456,In_666,In_757);
and U1457 (N_1457,In_140,In_565);
or U1458 (N_1458,In_298,In_521);
nand U1459 (N_1459,In_846,In_852);
and U1460 (N_1460,In_799,In_60);
nand U1461 (N_1461,In_255,In_793);
nor U1462 (N_1462,In_420,In_598);
or U1463 (N_1463,In_197,In_350);
or U1464 (N_1464,In_639,In_870);
nor U1465 (N_1465,In_136,In_109);
or U1466 (N_1466,In_204,In_139);
or U1467 (N_1467,In_31,In_759);
nor U1468 (N_1468,In_933,In_19);
and U1469 (N_1469,In_391,In_599);
nand U1470 (N_1470,In_96,In_79);
nand U1471 (N_1471,In_202,In_753);
nand U1472 (N_1472,In_584,In_508);
nand U1473 (N_1473,In_840,In_956);
and U1474 (N_1474,In_391,In_753);
nand U1475 (N_1475,In_49,In_579);
and U1476 (N_1476,In_118,In_871);
and U1477 (N_1477,In_605,In_858);
or U1478 (N_1478,In_852,In_79);
nand U1479 (N_1479,In_255,In_420);
or U1480 (N_1480,In_822,In_41);
xor U1481 (N_1481,In_726,In_187);
or U1482 (N_1482,In_607,In_551);
nand U1483 (N_1483,In_66,In_247);
nor U1484 (N_1484,In_151,In_855);
nand U1485 (N_1485,In_337,In_83);
nand U1486 (N_1486,In_626,In_661);
or U1487 (N_1487,In_797,In_240);
and U1488 (N_1488,In_616,In_889);
and U1489 (N_1489,In_403,In_57);
nand U1490 (N_1490,In_656,In_922);
and U1491 (N_1491,In_170,In_178);
nor U1492 (N_1492,In_505,In_0);
and U1493 (N_1493,In_484,In_447);
and U1494 (N_1494,In_940,In_565);
or U1495 (N_1495,In_829,In_613);
or U1496 (N_1496,In_553,In_396);
or U1497 (N_1497,In_603,In_67);
nand U1498 (N_1498,In_443,In_832);
or U1499 (N_1499,In_11,In_246);
nand U1500 (N_1500,In_373,In_513);
nor U1501 (N_1501,In_530,In_316);
nor U1502 (N_1502,In_62,In_315);
or U1503 (N_1503,In_762,In_676);
nand U1504 (N_1504,In_90,In_421);
nand U1505 (N_1505,In_961,In_365);
nand U1506 (N_1506,In_229,In_716);
nor U1507 (N_1507,In_187,In_768);
nand U1508 (N_1508,In_310,In_729);
or U1509 (N_1509,In_162,In_184);
nor U1510 (N_1510,In_278,In_203);
nand U1511 (N_1511,In_175,In_766);
nand U1512 (N_1512,In_967,In_540);
or U1513 (N_1513,In_995,In_943);
xnor U1514 (N_1514,In_959,In_294);
nor U1515 (N_1515,In_897,In_672);
nand U1516 (N_1516,In_77,In_391);
nor U1517 (N_1517,In_14,In_413);
xor U1518 (N_1518,In_122,In_761);
nand U1519 (N_1519,In_865,In_357);
xnor U1520 (N_1520,In_866,In_44);
nand U1521 (N_1521,In_352,In_263);
or U1522 (N_1522,In_832,In_587);
nand U1523 (N_1523,In_598,In_419);
or U1524 (N_1524,In_149,In_173);
and U1525 (N_1525,In_140,In_870);
nand U1526 (N_1526,In_977,In_207);
or U1527 (N_1527,In_942,In_857);
nand U1528 (N_1528,In_600,In_776);
and U1529 (N_1529,In_504,In_945);
and U1530 (N_1530,In_359,In_643);
and U1531 (N_1531,In_567,In_864);
nand U1532 (N_1532,In_11,In_433);
and U1533 (N_1533,In_359,In_654);
and U1534 (N_1534,In_943,In_529);
or U1535 (N_1535,In_254,In_565);
or U1536 (N_1536,In_477,In_884);
nand U1537 (N_1537,In_976,In_555);
nor U1538 (N_1538,In_677,In_859);
or U1539 (N_1539,In_113,In_37);
and U1540 (N_1540,In_513,In_169);
nand U1541 (N_1541,In_517,In_475);
and U1542 (N_1542,In_634,In_120);
and U1543 (N_1543,In_873,In_86);
or U1544 (N_1544,In_850,In_655);
or U1545 (N_1545,In_98,In_992);
nor U1546 (N_1546,In_771,In_830);
or U1547 (N_1547,In_276,In_438);
nor U1548 (N_1548,In_171,In_814);
and U1549 (N_1549,In_195,In_624);
and U1550 (N_1550,In_812,In_423);
and U1551 (N_1551,In_743,In_500);
and U1552 (N_1552,In_611,In_139);
or U1553 (N_1553,In_619,In_840);
nand U1554 (N_1554,In_952,In_835);
and U1555 (N_1555,In_670,In_1);
nor U1556 (N_1556,In_161,In_73);
and U1557 (N_1557,In_99,In_610);
and U1558 (N_1558,In_471,In_462);
or U1559 (N_1559,In_296,In_475);
and U1560 (N_1560,In_335,In_442);
nor U1561 (N_1561,In_436,In_603);
and U1562 (N_1562,In_384,In_122);
and U1563 (N_1563,In_887,In_58);
or U1564 (N_1564,In_136,In_837);
or U1565 (N_1565,In_422,In_720);
or U1566 (N_1566,In_485,In_962);
nor U1567 (N_1567,In_32,In_88);
and U1568 (N_1568,In_622,In_972);
and U1569 (N_1569,In_555,In_560);
and U1570 (N_1570,In_887,In_331);
nor U1571 (N_1571,In_873,In_821);
nand U1572 (N_1572,In_67,In_796);
or U1573 (N_1573,In_577,In_329);
and U1574 (N_1574,In_752,In_358);
or U1575 (N_1575,In_10,In_559);
xor U1576 (N_1576,In_181,In_502);
nor U1577 (N_1577,In_3,In_779);
or U1578 (N_1578,In_119,In_401);
nand U1579 (N_1579,In_307,In_993);
or U1580 (N_1580,In_846,In_990);
nor U1581 (N_1581,In_612,In_675);
or U1582 (N_1582,In_576,In_208);
nand U1583 (N_1583,In_710,In_840);
or U1584 (N_1584,In_22,In_212);
and U1585 (N_1585,In_63,In_682);
and U1586 (N_1586,In_361,In_671);
and U1587 (N_1587,In_566,In_533);
or U1588 (N_1588,In_648,In_630);
nor U1589 (N_1589,In_58,In_440);
nor U1590 (N_1590,In_987,In_337);
or U1591 (N_1591,In_847,In_471);
nor U1592 (N_1592,In_451,In_700);
and U1593 (N_1593,In_791,In_373);
or U1594 (N_1594,In_316,In_866);
and U1595 (N_1595,In_970,In_50);
or U1596 (N_1596,In_254,In_175);
and U1597 (N_1597,In_838,In_6);
nor U1598 (N_1598,In_303,In_989);
or U1599 (N_1599,In_860,In_358);
nand U1600 (N_1600,In_504,In_186);
nand U1601 (N_1601,In_897,In_3);
and U1602 (N_1602,In_737,In_642);
nor U1603 (N_1603,In_677,In_664);
or U1604 (N_1604,In_429,In_857);
nor U1605 (N_1605,In_427,In_814);
or U1606 (N_1606,In_23,In_444);
nor U1607 (N_1607,In_748,In_819);
nor U1608 (N_1608,In_425,In_253);
or U1609 (N_1609,In_897,In_121);
nand U1610 (N_1610,In_696,In_726);
nor U1611 (N_1611,In_919,In_125);
nand U1612 (N_1612,In_745,In_516);
nor U1613 (N_1613,In_262,In_841);
and U1614 (N_1614,In_908,In_387);
nor U1615 (N_1615,In_494,In_676);
nor U1616 (N_1616,In_323,In_908);
nand U1617 (N_1617,In_597,In_762);
nand U1618 (N_1618,In_983,In_484);
nor U1619 (N_1619,In_232,In_184);
or U1620 (N_1620,In_698,In_867);
or U1621 (N_1621,In_675,In_580);
nand U1622 (N_1622,In_233,In_788);
and U1623 (N_1623,In_926,In_216);
nor U1624 (N_1624,In_55,In_185);
nor U1625 (N_1625,In_600,In_526);
and U1626 (N_1626,In_696,In_642);
nor U1627 (N_1627,In_751,In_617);
and U1628 (N_1628,In_551,In_459);
and U1629 (N_1629,In_810,In_134);
and U1630 (N_1630,In_635,In_248);
or U1631 (N_1631,In_364,In_91);
nand U1632 (N_1632,In_313,In_618);
and U1633 (N_1633,In_343,In_66);
and U1634 (N_1634,In_325,In_578);
or U1635 (N_1635,In_294,In_996);
and U1636 (N_1636,In_687,In_314);
and U1637 (N_1637,In_752,In_664);
nand U1638 (N_1638,In_752,In_719);
nor U1639 (N_1639,In_94,In_256);
nand U1640 (N_1640,In_838,In_667);
nor U1641 (N_1641,In_888,In_264);
nand U1642 (N_1642,In_732,In_981);
and U1643 (N_1643,In_172,In_41);
and U1644 (N_1644,In_926,In_309);
or U1645 (N_1645,In_697,In_38);
and U1646 (N_1646,In_886,In_704);
or U1647 (N_1647,In_138,In_322);
nand U1648 (N_1648,In_53,In_466);
nand U1649 (N_1649,In_686,In_740);
nand U1650 (N_1650,In_292,In_407);
nor U1651 (N_1651,In_976,In_843);
nand U1652 (N_1652,In_544,In_747);
nor U1653 (N_1653,In_595,In_396);
nor U1654 (N_1654,In_58,In_231);
nor U1655 (N_1655,In_521,In_425);
and U1656 (N_1656,In_273,In_454);
nand U1657 (N_1657,In_936,In_35);
nand U1658 (N_1658,In_148,In_860);
or U1659 (N_1659,In_772,In_873);
nor U1660 (N_1660,In_278,In_364);
nand U1661 (N_1661,In_503,In_113);
nand U1662 (N_1662,In_362,In_396);
nor U1663 (N_1663,In_287,In_351);
nand U1664 (N_1664,In_139,In_127);
and U1665 (N_1665,In_816,In_50);
nor U1666 (N_1666,In_728,In_991);
nor U1667 (N_1667,In_365,In_444);
or U1668 (N_1668,In_43,In_461);
nand U1669 (N_1669,In_790,In_563);
and U1670 (N_1670,In_843,In_477);
and U1671 (N_1671,In_240,In_50);
nor U1672 (N_1672,In_108,In_112);
or U1673 (N_1673,In_602,In_469);
nor U1674 (N_1674,In_740,In_960);
nor U1675 (N_1675,In_596,In_471);
nand U1676 (N_1676,In_582,In_807);
nand U1677 (N_1677,In_501,In_951);
and U1678 (N_1678,In_646,In_618);
nor U1679 (N_1679,In_80,In_578);
nor U1680 (N_1680,In_709,In_729);
or U1681 (N_1681,In_164,In_292);
or U1682 (N_1682,In_925,In_852);
nor U1683 (N_1683,In_384,In_965);
nor U1684 (N_1684,In_679,In_629);
nor U1685 (N_1685,In_38,In_987);
nor U1686 (N_1686,In_262,In_534);
and U1687 (N_1687,In_981,In_33);
nand U1688 (N_1688,In_743,In_251);
and U1689 (N_1689,In_3,In_438);
nor U1690 (N_1690,In_877,In_833);
or U1691 (N_1691,In_447,In_322);
nor U1692 (N_1692,In_271,In_304);
nor U1693 (N_1693,In_4,In_7);
nand U1694 (N_1694,In_544,In_186);
nor U1695 (N_1695,In_365,In_120);
or U1696 (N_1696,In_486,In_234);
and U1697 (N_1697,In_10,In_704);
and U1698 (N_1698,In_373,In_275);
nor U1699 (N_1699,In_49,In_306);
and U1700 (N_1700,In_116,In_704);
and U1701 (N_1701,In_902,In_166);
nand U1702 (N_1702,In_717,In_268);
and U1703 (N_1703,In_757,In_312);
nor U1704 (N_1704,In_723,In_898);
and U1705 (N_1705,In_986,In_887);
nand U1706 (N_1706,In_88,In_637);
and U1707 (N_1707,In_848,In_50);
nor U1708 (N_1708,In_221,In_421);
nand U1709 (N_1709,In_34,In_854);
nor U1710 (N_1710,In_115,In_128);
and U1711 (N_1711,In_345,In_331);
nor U1712 (N_1712,In_44,In_871);
nor U1713 (N_1713,In_436,In_502);
and U1714 (N_1714,In_630,In_201);
nand U1715 (N_1715,In_210,In_469);
or U1716 (N_1716,In_748,In_44);
nor U1717 (N_1717,In_856,In_861);
nor U1718 (N_1718,In_206,In_513);
nand U1719 (N_1719,In_272,In_525);
and U1720 (N_1720,In_43,In_265);
and U1721 (N_1721,In_662,In_582);
or U1722 (N_1722,In_692,In_547);
or U1723 (N_1723,In_849,In_5);
and U1724 (N_1724,In_876,In_996);
nor U1725 (N_1725,In_152,In_595);
nand U1726 (N_1726,In_54,In_69);
nor U1727 (N_1727,In_405,In_693);
nand U1728 (N_1728,In_928,In_381);
and U1729 (N_1729,In_86,In_196);
nor U1730 (N_1730,In_972,In_957);
nor U1731 (N_1731,In_596,In_341);
nor U1732 (N_1732,In_906,In_48);
or U1733 (N_1733,In_902,In_754);
and U1734 (N_1734,In_871,In_92);
nor U1735 (N_1735,In_272,In_725);
and U1736 (N_1736,In_158,In_727);
nand U1737 (N_1737,In_282,In_637);
or U1738 (N_1738,In_879,In_749);
or U1739 (N_1739,In_288,In_836);
nor U1740 (N_1740,In_784,In_17);
and U1741 (N_1741,In_463,In_183);
nand U1742 (N_1742,In_451,In_915);
nor U1743 (N_1743,In_509,In_198);
or U1744 (N_1744,In_512,In_273);
and U1745 (N_1745,In_663,In_866);
nor U1746 (N_1746,In_262,In_636);
nand U1747 (N_1747,In_717,In_10);
nor U1748 (N_1748,In_631,In_521);
nor U1749 (N_1749,In_45,In_32);
and U1750 (N_1750,In_272,In_710);
nor U1751 (N_1751,In_911,In_42);
nand U1752 (N_1752,In_6,In_27);
nor U1753 (N_1753,In_88,In_535);
nand U1754 (N_1754,In_438,In_590);
and U1755 (N_1755,In_272,In_875);
nand U1756 (N_1756,In_670,In_955);
nand U1757 (N_1757,In_417,In_976);
xor U1758 (N_1758,In_143,In_921);
or U1759 (N_1759,In_515,In_778);
nor U1760 (N_1760,In_431,In_957);
nand U1761 (N_1761,In_98,In_243);
nand U1762 (N_1762,In_87,In_633);
nor U1763 (N_1763,In_558,In_601);
nand U1764 (N_1764,In_893,In_492);
or U1765 (N_1765,In_152,In_719);
or U1766 (N_1766,In_578,In_205);
and U1767 (N_1767,In_168,In_323);
nor U1768 (N_1768,In_799,In_862);
or U1769 (N_1769,In_612,In_664);
or U1770 (N_1770,In_341,In_879);
nor U1771 (N_1771,In_131,In_434);
nand U1772 (N_1772,In_928,In_270);
or U1773 (N_1773,In_179,In_395);
or U1774 (N_1774,In_126,In_607);
nand U1775 (N_1775,In_748,In_755);
or U1776 (N_1776,In_483,In_71);
nor U1777 (N_1777,In_190,In_266);
or U1778 (N_1778,In_575,In_531);
and U1779 (N_1779,In_743,In_692);
nand U1780 (N_1780,In_395,In_798);
nor U1781 (N_1781,In_113,In_450);
or U1782 (N_1782,In_52,In_829);
nand U1783 (N_1783,In_888,In_366);
nand U1784 (N_1784,In_447,In_940);
or U1785 (N_1785,In_751,In_894);
or U1786 (N_1786,In_409,In_180);
nand U1787 (N_1787,In_93,In_8);
nor U1788 (N_1788,In_155,In_558);
or U1789 (N_1789,In_601,In_807);
and U1790 (N_1790,In_482,In_182);
or U1791 (N_1791,In_545,In_496);
xnor U1792 (N_1792,In_88,In_542);
and U1793 (N_1793,In_627,In_785);
nand U1794 (N_1794,In_6,In_530);
nand U1795 (N_1795,In_27,In_0);
and U1796 (N_1796,In_41,In_163);
nor U1797 (N_1797,In_142,In_366);
and U1798 (N_1798,In_441,In_568);
and U1799 (N_1799,In_270,In_522);
or U1800 (N_1800,In_709,In_56);
or U1801 (N_1801,In_839,In_84);
nand U1802 (N_1802,In_381,In_623);
or U1803 (N_1803,In_292,In_619);
or U1804 (N_1804,In_246,In_681);
and U1805 (N_1805,In_852,In_8);
nand U1806 (N_1806,In_812,In_799);
xor U1807 (N_1807,In_509,In_479);
nor U1808 (N_1808,In_724,In_719);
nand U1809 (N_1809,In_836,In_214);
nand U1810 (N_1810,In_637,In_552);
and U1811 (N_1811,In_423,In_252);
or U1812 (N_1812,In_268,In_889);
and U1813 (N_1813,In_315,In_836);
nor U1814 (N_1814,In_759,In_189);
or U1815 (N_1815,In_503,In_609);
or U1816 (N_1816,In_982,In_37);
nor U1817 (N_1817,In_174,In_380);
and U1818 (N_1818,In_15,In_153);
nand U1819 (N_1819,In_833,In_972);
or U1820 (N_1820,In_316,In_40);
nor U1821 (N_1821,In_481,In_764);
nand U1822 (N_1822,In_267,In_93);
and U1823 (N_1823,In_126,In_800);
nor U1824 (N_1824,In_632,In_856);
nor U1825 (N_1825,In_61,In_273);
nand U1826 (N_1826,In_255,In_953);
and U1827 (N_1827,In_93,In_209);
nor U1828 (N_1828,In_45,In_433);
nand U1829 (N_1829,In_53,In_52);
and U1830 (N_1830,In_599,In_154);
nor U1831 (N_1831,In_775,In_71);
nor U1832 (N_1832,In_925,In_953);
nand U1833 (N_1833,In_926,In_880);
or U1834 (N_1834,In_309,In_544);
nor U1835 (N_1835,In_746,In_336);
nand U1836 (N_1836,In_478,In_594);
nor U1837 (N_1837,In_797,In_525);
nor U1838 (N_1838,In_230,In_770);
or U1839 (N_1839,In_806,In_261);
and U1840 (N_1840,In_855,In_630);
and U1841 (N_1841,In_205,In_892);
or U1842 (N_1842,In_966,In_337);
nand U1843 (N_1843,In_50,In_554);
nor U1844 (N_1844,In_200,In_665);
nor U1845 (N_1845,In_686,In_20);
nand U1846 (N_1846,In_218,In_408);
or U1847 (N_1847,In_93,In_551);
nor U1848 (N_1848,In_482,In_752);
and U1849 (N_1849,In_99,In_778);
or U1850 (N_1850,In_363,In_270);
and U1851 (N_1851,In_862,In_943);
or U1852 (N_1852,In_623,In_308);
nand U1853 (N_1853,In_109,In_764);
nand U1854 (N_1854,In_828,In_669);
xor U1855 (N_1855,In_433,In_333);
nand U1856 (N_1856,In_780,In_45);
or U1857 (N_1857,In_75,In_232);
and U1858 (N_1858,In_12,In_841);
nor U1859 (N_1859,In_554,In_152);
or U1860 (N_1860,In_373,In_190);
nor U1861 (N_1861,In_593,In_457);
nand U1862 (N_1862,In_798,In_827);
or U1863 (N_1863,In_975,In_292);
nand U1864 (N_1864,In_448,In_305);
or U1865 (N_1865,In_399,In_923);
nor U1866 (N_1866,In_916,In_94);
or U1867 (N_1867,In_4,In_292);
or U1868 (N_1868,In_923,In_49);
or U1869 (N_1869,In_846,In_36);
nand U1870 (N_1870,In_122,In_841);
and U1871 (N_1871,In_403,In_735);
nand U1872 (N_1872,In_903,In_159);
or U1873 (N_1873,In_230,In_835);
or U1874 (N_1874,In_358,In_376);
or U1875 (N_1875,In_445,In_135);
nand U1876 (N_1876,In_799,In_195);
nor U1877 (N_1877,In_560,In_658);
nor U1878 (N_1878,In_343,In_3);
and U1879 (N_1879,In_518,In_649);
nor U1880 (N_1880,In_588,In_170);
or U1881 (N_1881,In_142,In_356);
and U1882 (N_1882,In_61,In_97);
nor U1883 (N_1883,In_572,In_485);
nor U1884 (N_1884,In_47,In_406);
nor U1885 (N_1885,In_669,In_689);
nor U1886 (N_1886,In_682,In_625);
or U1887 (N_1887,In_639,In_323);
nand U1888 (N_1888,In_623,In_732);
and U1889 (N_1889,In_419,In_635);
nand U1890 (N_1890,In_993,In_627);
and U1891 (N_1891,In_274,In_278);
and U1892 (N_1892,In_430,In_815);
and U1893 (N_1893,In_253,In_671);
nor U1894 (N_1894,In_194,In_904);
and U1895 (N_1895,In_692,In_79);
nand U1896 (N_1896,In_370,In_144);
nand U1897 (N_1897,In_189,In_597);
or U1898 (N_1898,In_394,In_114);
nor U1899 (N_1899,In_721,In_276);
or U1900 (N_1900,In_782,In_98);
nand U1901 (N_1901,In_422,In_428);
or U1902 (N_1902,In_913,In_32);
nor U1903 (N_1903,In_94,In_226);
or U1904 (N_1904,In_583,In_887);
and U1905 (N_1905,In_661,In_465);
or U1906 (N_1906,In_254,In_355);
and U1907 (N_1907,In_258,In_983);
nand U1908 (N_1908,In_278,In_999);
nand U1909 (N_1909,In_976,In_913);
nand U1910 (N_1910,In_903,In_166);
or U1911 (N_1911,In_639,In_609);
nand U1912 (N_1912,In_865,In_682);
nand U1913 (N_1913,In_549,In_722);
nor U1914 (N_1914,In_699,In_635);
and U1915 (N_1915,In_769,In_733);
and U1916 (N_1916,In_937,In_86);
nor U1917 (N_1917,In_584,In_225);
or U1918 (N_1918,In_705,In_861);
nor U1919 (N_1919,In_246,In_316);
xnor U1920 (N_1920,In_789,In_605);
nor U1921 (N_1921,In_818,In_123);
nor U1922 (N_1922,In_976,In_152);
or U1923 (N_1923,In_942,In_887);
and U1924 (N_1924,In_158,In_399);
nand U1925 (N_1925,In_544,In_19);
and U1926 (N_1926,In_972,In_234);
nor U1927 (N_1927,In_215,In_385);
nand U1928 (N_1928,In_298,In_881);
and U1929 (N_1929,In_707,In_709);
nor U1930 (N_1930,In_501,In_297);
nor U1931 (N_1931,In_454,In_905);
or U1932 (N_1932,In_75,In_558);
nor U1933 (N_1933,In_577,In_785);
nor U1934 (N_1934,In_694,In_618);
or U1935 (N_1935,In_343,In_897);
nor U1936 (N_1936,In_695,In_795);
or U1937 (N_1937,In_982,In_720);
nand U1938 (N_1938,In_324,In_77);
and U1939 (N_1939,In_450,In_529);
or U1940 (N_1940,In_199,In_603);
nor U1941 (N_1941,In_497,In_442);
and U1942 (N_1942,In_413,In_498);
or U1943 (N_1943,In_907,In_337);
nor U1944 (N_1944,In_579,In_98);
or U1945 (N_1945,In_108,In_500);
or U1946 (N_1946,In_202,In_607);
nand U1947 (N_1947,In_70,In_352);
or U1948 (N_1948,In_778,In_59);
or U1949 (N_1949,In_505,In_296);
or U1950 (N_1950,In_969,In_905);
nand U1951 (N_1951,In_923,In_993);
and U1952 (N_1952,In_865,In_37);
nor U1953 (N_1953,In_916,In_754);
nor U1954 (N_1954,In_640,In_754);
nor U1955 (N_1955,In_462,In_508);
and U1956 (N_1956,In_298,In_204);
and U1957 (N_1957,In_811,In_281);
and U1958 (N_1958,In_432,In_473);
nand U1959 (N_1959,In_192,In_329);
and U1960 (N_1960,In_731,In_849);
nor U1961 (N_1961,In_356,In_505);
nor U1962 (N_1962,In_853,In_698);
and U1963 (N_1963,In_597,In_115);
nor U1964 (N_1964,In_933,In_150);
nor U1965 (N_1965,In_318,In_366);
nor U1966 (N_1966,In_313,In_833);
and U1967 (N_1967,In_294,In_818);
nor U1968 (N_1968,In_491,In_635);
nor U1969 (N_1969,In_464,In_270);
nand U1970 (N_1970,In_110,In_335);
nand U1971 (N_1971,In_920,In_722);
nand U1972 (N_1972,In_407,In_846);
nand U1973 (N_1973,In_297,In_47);
or U1974 (N_1974,In_744,In_630);
nand U1975 (N_1975,In_517,In_813);
nor U1976 (N_1976,In_876,In_338);
and U1977 (N_1977,In_786,In_182);
or U1978 (N_1978,In_859,In_99);
or U1979 (N_1979,In_792,In_885);
nand U1980 (N_1980,In_708,In_13);
nand U1981 (N_1981,In_873,In_101);
and U1982 (N_1982,In_643,In_869);
nand U1983 (N_1983,In_916,In_398);
nand U1984 (N_1984,In_702,In_824);
and U1985 (N_1985,In_498,In_975);
nand U1986 (N_1986,In_65,In_722);
nand U1987 (N_1987,In_571,In_449);
and U1988 (N_1988,In_821,In_908);
and U1989 (N_1989,In_58,In_453);
nor U1990 (N_1990,In_945,In_355);
and U1991 (N_1991,In_93,In_934);
or U1992 (N_1992,In_902,In_375);
nor U1993 (N_1993,In_666,In_306);
and U1994 (N_1994,In_4,In_558);
or U1995 (N_1995,In_450,In_38);
and U1996 (N_1996,In_227,In_505);
or U1997 (N_1997,In_238,In_315);
and U1998 (N_1998,In_227,In_770);
and U1999 (N_1999,In_828,In_501);
and U2000 (N_2000,In_578,In_194);
nand U2001 (N_2001,In_569,In_649);
nand U2002 (N_2002,In_388,In_713);
nand U2003 (N_2003,In_974,In_534);
or U2004 (N_2004,In_836,In_356);
nand U2005 (N_2005,In_475,In_485);
nand U2006 (N_2006,In_376,In_981);
nor U2007 (N_2007,In_508,In_992);
nor U2008 (N_2008,In_348,In_78);
nand U2009 (N_2009,In_104,In_841);
nand U2010 (N_2010,In_418,In_886);
nor U2011 (N_2011,In_515,In_843);
nand U2012 (N_2012,In_374,In_620);
nand U2013 (N_2013,In_172,In_378);
and U2014 (N_2014,In_588,In_186);
nand U2015 (N_2015,In_548,In_612);
nand U2016 (N_2016,In_915,In_208);
or U2017 (N_2017,In_822,In_789);
or U2018 (N_2018,In_202,In_786);
nor U2019 (N_2019,In_694,In_560);
or U2020 (N_2020,In_958,In_422);
nand U2021 (N_2021,In_846,In_55);
nor U2022 (N_2022,In_722,In_256);
or U2023 (N_2023,In_164,In_416);
nand U2024 (N_2024,In_89,In_92);
nor U2025 (N_2025,In_364,In_909);
nand U2026 (N_2026,In_166,In_770);
and U2027 (N_2027,In_286,In_93);
nand U2028 (N_2028,In_488,In_301);
nor U2029 (N_2029,In_764,In_635);
nor U2030 (N_2030,In_107,In_552);
or U2031 (N_2031,In_937,In_673);
or U2032 (N_2032,In_367,In_414);
and U2033 (N_2033,In_202,In_836);
nand U2034 (N_2034,In_590,In_310);
nor U2035 (N_2035,In_772,In_397);
nand U2036 (N_2036,In_596,In_466);
nor U2037 (N_2037,In_714,In_33);
and U2038 (N_2038,In_610,In_880);
and U2039 (N_2039,In_500,In_136);
nand U2040 (N_2040,In_647,In_713);
or U2041 (N_2041,In_454,In_732);
nor U2042 (N_2042,In_888,In_328);
nand U2043 (N_2043,In_98,In_551);
or U2044 (N_2044,In_609,In_430);
nor U2045 (N_2045,In_763,In_605);
nor U2046 (N_2046,In_954,In_932);
nor U2047 (N_2047,In_639,In_930);
and U2048 (N_2048,In_633,In_624);
nor U2049 (N_2049,In_185,In_166);
or U2050 (N_2050,In_513,In_749);
or U2051 (N_2051,In_297,In_953);
and U2052 (N_2052,In_121,In_788);
nor U2053 (N_2053,In_645,In_398);
or U2054 (N_2054,In_656,In_731);
and U2055 (N_2055,In_236,In_706);
or U2056 (N_2056,In_511,In_965);
nor U2057 (N_2057,In_172,In_836);
nor U2058 (N_2058,In_159,In_346);
and U2059 (N_2059,In_51,In_218);
and U2060 (N_2060,In_380,In_528);
or U2061 (N_2061,In_631,In_688);
nand U2062 (N_2062,In_332,In_434);
and U2063 (N_2063,In_847,In_370);
nor U2064 (N_2064,In_99,In_352);
and U2065 (N_2065,In_337,In_466);
nor U2066 (N_2066,In_882,In_256);
nor U2067 (N_2067,In_485,In_675);
or U2068 (N_2068,In_571,In_405);
or U2069 (N_2069,In_681,In_725);
nor U2070 (N_2070,In_868,In_161);
or U2071 (N_2071,In_383,In_385);
and U2072 (N_2072,In_22,In_248);
or U2073 (N_2073,In_715,In_325);
and U2074 (N_2074,In_470,In_364);
and U2075 (N_2075,In_888,In_294);
nor U2076 (N_2076,In_529,In_707);
nand U2077 (N_2077,In_913,In_743);
and U2078 (N_2078,In_823,In_62);
nor U2079 (N_2079,In_772,In_202);
or U2080 (N_2080,In_953,In_643);
or U2081 (N_2081,In_665,In_746);
nand U2082 (N_2082,In_193,In_676);
or U2083 (N_2083,In_796,In_300);
or U2084 (N_2084,In_378,In_919);
nand U2085 (N_2085,In_771,In_976);
and U2086 (N_2086,In_711,In_69);
xor U2087 (N_2087,In_479,In_543);
or U2088 (N_2088,In_668,In_706);
nor U2089 (N_2089,In_838,In_699);
nand U2090 (N_2090,In_994,In_102);
nor U2091 (N_2091,In_819,In_906);
nor U2092 (N_2092,In_54,In_861);
and U2093 (N_2093,In_149,In_634);
and U2094 (N_2094,In_242,In_934);
nand U2095 (N_2095,In_74,In_608);
and U2096 (N_2096,In_497,In_100);
nor U2097 (N_2097,In_470,In_967);
or U2098 (N_2098,In_491,In_528);
nor U2099 (N_2099,In_876,In_578);
and U2100 (N_2100,In_324,In_166);
and U2101 (N_2101,In_340,In_383);
nand U2102 (N_2102,In_559,In_113);
and U2103 (N_2103,In_316,In_678);
nor U2104 (N_2104,In_872,In_354);
and U2105 (N_2105,In_283,In_993);
or U2106 (N_2106,In_522,In_680);
or U2107 (N_2107,In_289,In_146);
or U2108 (N_2108,In_371,In_849);
nand U2109 (N_2109,In_505,In_117);
nor U2110 (N_2110,In_142,In_229);
and U2111 (N_2111,In_102,In_192);
and U2112 (N_2112,In_33,In_106);
nand U2113 (N_2113,In_739,In_771);
nor U2114 (N_2114,In_659,In_471);
and U2115 (N_2115,In_419,In_37);
nor U2116 (N_2116,In_650,In_385);
or U2117 (N_2117,In_76,In_208);
nand U2118 (N_2118,In_318,In_957);
nor U2119 (N_2119,In_336,In_431);
nor U2120 (N_2120,In_518,In_678);
nor U2121 (N_2121,In_873,In_246);
and U2122 (N_2122,In_212,In_937);
nand U2123 (N_2123,In_468,In_310);
nor U2124 (N_2124,In_924,In_554);
or U2125 (N_2125,In_763,In_143);
nand U2126 (N_2126,In_85,In_215);
or U2127 (N_2127,In_933,In_351);
or U2128 (N_2128,In_209,In_543);
and U2129 (N_2129,In_57,In_689);
or U2130 (N_2130,In_589,In_574);
nor U2131 (N_2131,In_947,In_972);
nand U2132 (N_2132,In_784,In_331);
and U2133 (N_2133,In_405,In_374);
or U2134 (N_2134,In_780,In_640);
and U2135 (N_2135,In_717,In_537);
xnor U2136 (N_2136,In_408,In_392);
nor U2137 (N_2137,In_235,In_940);
and U2138 (N_2138,In_60,In_853);
and U2139 (N_2139,In_991,In_614);
and U2140 (N_2140,In_521,In_964);
nor U2141 (N_2141,In_810,In_749);
and U2142 (N_2142,In_800,In_150);
nand U2143 (N_2143,In_941,In_879);
nand U2144 (N_2144,In_138,In_118);
and U2145 (N_2145,In_710,In_104);
and U2146 (N_2146,In_333,In_70);
nand U2147 (N_2147,In_446,In_769);
nor U2148 (N_2148,In_942,In_971);
and U2149 (N_2149,In_168,In_216);
or U2150 (N_2150,In_190,In_380);
nor U2151 (N_2151,In_429,In_84);
and U2152 (N_2152,In_651,In_257);
nor U2153 (N_2153,In_46,In_265);
or U2154 (N_2154,In_714,In_377);
or U2155 (N_2155,In_860,In_8);
and U2156 (N_2156,In_698,In_27);
or U2157 (N_2157,In_259,In_122);
or U2158 (N_2158,In_280,In_384);
nor U2159 (N_2159,In_576,In_251);
xor U2160 (N_2160,In_423,In_373);
and U2161 (N_2161,In_184,In_973);
nand U2162 (N_2162,In_900,In_424);
and U2163 (N_2163,In_629,In_838);
nor U2164 (N_2164,In_51,In_161);
nand U2165 (N_2165,In_366,In_853);
nor U2166 (N_2166,In_529,In_122);
xnor U2167 (N_2167,In_335,In_112);
nor U2168 (N_2168,In_55,In_53);
and U2169 (N_2169,In_453,In_925);
and U2170 (N_2170,In_312,In_781);
nor U2171 (N_2171,In_123,In_187);
or U2172 (N_2172,In_811,In_33);
and U2173 (N_2173,In_337,In_363);
or U2174 (N_2174,In_553,In_501);
nor U2175 (N_2175,In_667,In_581);
nand U2176 (N_2176,In_786,In_603);
nand U2177 (N_2177,In_861,In_801);
or U2178 (N_2178,In_913,In_853);
nor U2179 (N_2179,In_314,In_703);
or U2180 (N_2180,In_795,In_277);
nand U2181 (N_2181,In_211,In_371);
or U2182 (N_2182,In_699,In_674);
nor U2183 (N_2183,In_271,In_773);
nor U2184 (N_2184,In_536,In_571);
nand U2185 (N_2185,In_856,In_931);
nand U2186 (N_2186,In_766,In_632);
or U2187 (N_2187,In_738,In_387);
nor U2188 (N_2188,In_245,In_998);
and U2189 (N_2189,In_411,In_13);
nor U2190 (N_2190,In_658,In_590);
or U2191 (N_2191,In_981,In_888);
nand U2192 (N_2192,In_571,In_390);
and U2193 (N_2193,In_993,In_468);
or U2194 (N_2194,In_523,In_736);
or U2195 (N_2195,In_860,In_144);
and U2196 (N_2196,In_751,In_815);
nand U2197 (N_2197,In_620,In_360);
nand U2198 (N_2198,In_47,In_251);
nand U2199 (N_2199,In_665,In_530);
nor U2200 (N_2200,In_175,In_360);
nor U2201 (N_2201,In_304,In_350);
nor U2202 (N_2202,In_373,In_146);
and U2203 (N_2203,In_303,In_362);
or U2204 (N_2204,In_817,In_90);
and U2205 (N_2205,In_830,In_645);
and U2206 (N_2206,In_619,In_171);
or U2207 (N_2207,In_413,In_692);
nand U2208 (N_2208,In_240,In_25);
or U2209 (N_2209,In_178,In_350);
nand U2210 (N_2210,In_87,In_290);
and U2211 (N_2211,In_223,In_629);
and U2212 (N_2212,In_219,In_127);
nand U2213 (N_2213,In_353,In_95);
nand U2214 (N_2214,In_711,In_817);
nor U2215 (N_2215,In_284,In_453);
and U2216 (N_2216,In_391,In_479);
nor U2217 (N_2217,In_799,In_216);
and U2218 (N_2218,In_382,In_518);
nor U2219 (N_2219,In_514,In_87);
and U2220 (N_2220,In_381,In_484);
or U2221 (N_2221,In_437,In_72);
or U2222 (N_2222,In_123,In_642);
and U2223 (N_2223,In_409,In_890);
nor U2224 (N_2224,In_889,In_831);
nor U2225 (N_2225,In_411,In_320);
nor U2226 (N_2226,In_571,In_854);
and U2227 (N_2227,In_7,In_219);
nor U2228 (N_2228,In_934,In_920);
or U2229 (N_2229,In_477,In_743);
nand U2230 (N_2230,In_709,In_16);
nand U2231 (N_2231,In_75,In_471);
or U2232 (N_2232,In_579,In_209);
nand U2233 (N_2233,In_169,In_554);
and U2234 (N_2234,In_49,In_340);
or U2235 (N_2235,In_144,In_170);
nor U2236 (N_2236,In_941,In_755);
or U2237 (N_2237,In_467,In_267);
nor U2238 (N_2238,In_96,In_118);
nor U2239 (N_2239,In_206,In_267);
nand U2240 (N_2240,In_717,In_145);
or U2241 (N_2241,In_291,In_676);
nand U2242 (N_2242,In_661,In_56);
nor U2243 (N_2243,In_847,In_200);
or U2244 (N_2244,In_599,In_728);
or U2245 (N_2245,In_458,In_622);
nand U2246 (N_2246,In_366,In_481);
nor U2247 (N_2247,In_878,In_627);
or U2248 (N_2248,In_275,In_770);
nor U2249 (N_2249,In_304,In_532);
nor U2250 (N_2250,In_91,In_425);
or U2251 (N_2251,In_256,In_254);
nand U2252 (N_2252,In_440,In_73);
nand U2253 (N_2253,In_674,In_499);
nor U2254 (N_2254,In_802,In_652);
or U2255 (N_2255,In_206,In_116);
xnor U2256 (N_2256,In_223,In_343);
or U2257 (N_2257,In_900,In_624);
or U2258 (N_2258,In_1,In_88);
and U2259 (N_2259,In_852,In_244);
nand U2260 (N_2260,In_311,In_532);
nor U2261 (N_2261,In_719,In_571);
nand U2262 (N_2262,In_747,In_259);
and U2263 (N_2263,In_801,In_446);
or U2264 (N_2264,In_251,In_162);
nand U2265 (N_2265,In_336,In_527);
or U2266 (N_2266,In_151,In_360);
and U2267 (N_2267,In_938,In_94);
and U2268 (N_2268,In_428,In_1);
or U2269 (N_2269,In_519,In_635);
or U2270 (N_2270,In_209,In_354);
nor U2271 (N_2271,In_642,In_558);
nand U2272 (N_2272,In_743,In_734);
nand U2273 (N_2273,In_856,In_201);
or U2274 (N_2274,In_42,In_255);
and U2275 (N_2275,In_191,In_25);
nor U2276 (N_2276,In_382,In_556);
or U2277 (N_2277,In_108,In_101);
and U2278 (N_2278,In_988,In_107);
or U2279 (N_2279,In_644,In_605);
nor U2280 (N_2280,In_361,In_317);
nand U2281 (N_2281,In_128,In_525);
and U2282 (N_2282,In_799,In_61);
nor U2283 (N_2283,In_428,In_920);
nor U2284 (N_2284,In_275,In_341);
or U2285 (N_2285,In_339,In_852);
or U2286 (N_2286,In_409,In_423);
nand U2287 (N_2287,In_927,In_184);
nor U2288 (N_2288,In_371,In_462);
nor U2289 (N_2289,In_603,In_584);
or U2290 (N_2290,In_411,In_500);
nor U2291 (N_2291,In_28,In_870);
nand U2292 (N_2292,In_651,In_0);
or U2293 (N_2293,In_789,In_955);
and U2294 (N_2294,In_173,In_163);
nand U2295 (N_2295,In_22,In_328);
nor U2296 (N_2296,In_93,In_481);
nor U2297 (N_2297,In_502,In_349);
nand U2298 (N_2298,In_612,In_995);
nand U2299 (N_2299,In_356,In_886);
and U2300 (N_2300,In_894,In_622);
nand U2301 (N_2301,In_632,In_13);
nand U2302 (N_2302,In_816,In_311);
nand U2303 (N_2303,In_700,In_988);
or U2304 (N_2304,In_402,In_94);
nor U2305 (N_2305,In_777,In_539);
and U2306 (N_2306,In_410,In_867);
and U2307 (N_2307,In_870,In_482);
nand U2308 (N_2308,In_292,In_764);
nor U2309 (N_2309,In_775,In_956);
or U2310 (N_2310,In_961,In_209);
or U2311 (N_2311,In_776,In_857);
and U2312 (N_2312,In_593,In_453);
nor U2313 (N_2313,In_110,In_599);
or U2314 (N_2314,In_935,In_142);
and U2315 (N_2315,In_674,In_135);
and U2316 (N_2316,In_33,In_54);
and U2317 (N_2317,In_221,In_356);
or U2318 (N_2318,In_398,In_438);
or U2319 (N_2319,In_721,In_994);
nand U2320 (N_2320,In_742,In_995);
or U2321 (N_2321,In_295,In_666);
and U2322 (N_2322,In_500,In_688);
or U2323 (N_2323,In_849,In_13);
and U2324 (N_2324,In_544,In_229);
or U2325 (N_2325,In_842,In_518);
xnor U2326 (N_2326,In_364,In_311);
or U2327 (N_2327,In_97,In_316);
and U2328 (N_2328,In_670,In_512);
nand U2329 (N_2329,In_636,In_190);
nand U2330 (N_2330,In_673,In_487);
nand U2331 (N_2331,In_268,In_611);
nand U2332 (N_2332,In_327,In_464);
and U2333 (N_2333,In_518,In_614);
or U2334 (N_2334,In_140,In_990);
and U2335 (N_2335,In_825,In_363);
nor U2336 (N_2336,In_418,In_720);
nand U2337 (N_2337,In_452,In_666);
and U2338 (N_2338,In_628,In_753);
and U2339 (N_2339,In_217,In_586);
xor U2340 (N_2340,In_986,In_670);
and U2341 (N_2341,In_509,In_687);
and U2342 (N_2342,In_619,In_911);
nor U2343 (N_2343,In_58,In_586);
or U2344 (N_2344,In_114,In_100);
nand U2345 (N_2345,In_825,In_797);
and U2346 (N_2346,In_292,In_445);
nor U2347 (N_2347,In_159,In_66);
nor U2348 (N_2348,In_831,In_923);
nand U2349 (N_2349,In_612,In_335);
nor U2350 (N_2350,In_795,In_314);
nand U2351 (N_2351,In_805,In_892);
or U2352 (N_2352,In_666,In_886);
nor U2353 (N_2353,In_730,In_412);
nor U2354 (N_2354,In_286,In_703);
or U2355 (N_2355,In_784,In_50);
nor U2356 (N_2356,In_389,In_187);
nand U2357 (N_2357,In_397,In_198);
and U2358 (N_2358,In_191,In_939);
or U2359 (N_2359,In_860,In_799);
nor U2360 (N_2360,In_315,In_10);
nand U2361 (N_2361,In_348,In_857);
nand U2362 (N_2362,In_108,In_964);
and U2363 (N_2363,In_370,In_688);
nor U2364 (N_2364,In_291,In_691);
or U2365 (N_2365,In_236,In_115);
nand U2366 (N_2366,In_887,In_854);
or U2367 (N_2367,In_990,In_435);
or U2368 (N_2368,In_28,In_811);
or U2369 (N_2369,In_752,In_894);
or U2370 (N_2370,In_510,In_910);
or U2371 (N_2371,In_693,In_77);
and U2372 (N_2372,In_396,In_593);
and U2373 (N_2373,In_424,In_812);
and U2374 (N_2374,In_60,In_769);
nor U2375 (N_2375,In_926,In_992);
nand U2376 (N_2376,In_694,In_635);
nand U2377 (N_2377,In_994,In_191);
nand U2378 (N_2378,In_389,In_732);
or U2379 (N_2379,In_16,In_405);
and U2380 (N_2380,In_856,In_948);
or U2381 (N_2381,In_203,In_389);
nand U2382 (N_2382,In_611,In_125);
nor U2383 (N_2383,In_485,In_797);
nor U2384 (N_2384,In_536,In_347);
nor U2385 (N_2385,In_525,In_868);
nor U2386 (N_2386,In_27,In_153);
and U2387 (N_2387,In_237,In_763);
or U2388 (N_2388,In_982,In_519);
nand U2389 (N_2389,In_66,In_414);
nand U2390 (N_2390,In_266,In_306);
nor U2391 (N_2391,In_428,In_820);
or U2392 (N_2392,In_966,In_44);
nor U2393 (N_2393,In_15,In_973);
or U2394 (N_2394,In_716,In_934);
or U2395 (N_2395,In_236,In_692);
or U2396 (N_2396,In_756,In_278);
nor U2397 (N_2397,In_569,In_51);
nand U2398 (N_2398,In_698,In_835);
and U2399 (N_2399,In_953,In_717);
and U2400 (N_2400,In_606,In_41);
nor U2401 (N_2401,In_127,In_835);
and U2402 (N_2402,In_258,In_841);
nand U2403 (N_2403,In_723,In_45);
nand U2404 (N_2404,In_228,In_892);
nand U2405 (N_2405,In_241,In_428);
and U2406 (N_2406,In_36,In_229);
nand U2407 (N_2407,In_837,In_326);
nand U2408 (N_2408,In_288,In_465);
nand U2409 (N_2409,In_86,In_407);
and U2410 (N_2410,In_452,In_61);
nand U2411 (N_2411,In_686,In_645);
nor U2412 (N_2412,In_611,In_218);
or U2413 (N_2413,In_582,In_818);
and U2414 (N_2414,In_861,In_683);
nor U2415 (N_2415,In_211,In_997);
and U2416 (N_2416,In_503,In_120);
nor U2417 (N_2417,In_874,In_244);
nor U2418 (N_2418,In_68,In_177);
nor U2419 (N_2419,In_573,In_977);
or U2420 (N_2420,In_865,In_506);
xnor U2421 (N_2421,In_223,In_295);
or U2422 (N_2422,In_459,In_360);
nand U2423 (N_2423,In_350,In_111);
and U2424 (N_2424,In_745,In_650);
nand U2425 (N_2425,In_813,In_164);
and U2426 (N_2426,In_283,In_498);
and U2427 (N_2427,In_93,In_817);
and U2428 (N_2428,In_241,In_666);
or U2429 (N_2429,In_648,In_259);
nor U2430 (N_2430,In_193,In_691);
and U2431 (N_2431,In_348,In_43);
and U2432 (N_2432,In_310,In_853);
nor U2433 (N_2433,In_563,In_833);
and U2434 (N_2434,In_344,In_656);
and U2435 (N_2435,In_707,In_902);
xor U2436 (N_2436,In_507,In_252);
and U2437 (N_2437,In_789,In_394);
and U2438 (N_2438,In_145,In_798);
nor U2439 (N_2439,In_39,In_852);
nand U2440 (N_2440,In_542,In_39);
nor U2441 (N_2441,In_656,In_433);
or U2442 (N_2442,In_689,In_475);
or U2443 (N_2443,In_406,In_594);
nand U2444 (N_2444,In_481,In_991);
nand U2445 (N_2445,In_616,In_108);
and U2446 (N_2446,In_234,In_830);
nand U2447 (N_2447,In_652,In_475);
nand U2448 (N_2448,In_819,In_420);
nor U2449 (N_2449,In_658,In_986);
and U2450 (N_2450,In_536,In_240);
nand U2451 (N_2451,In_402,In_387);
or U2452 (N_2452,In_715,In_988);
and U2453 (N_2453,In_921,In_875);
nand U2454 (N_2454,In_235,In_913);
or U2455 (N_2455,In_594,In_152);
nand U2456 (N_2456,In_38,In_468);
nor U2457 (N_2457,In_120,In_597);
nor U2458 (N_2458,In_939,In_119);
and U2459 (N_2459,In_863,In_312);
and U2460 (N_2460,In_34,In_911);
or U2461 (N_2461,In_444,In_807);
and U2462 (N_2462,In_369,In_439);
nor U2463 (N_2463,In_226,In_744);
nor U2464 (N_2464,In_218,In_774);
or U2465 (N_2465,In_73,In_400);
nand U2466 (N_2466,In_879,In_110);
or U2467 (N_2467,In_502,In_487);
nand U2468 (N_2468,In_351,In_773);
nand U2469 (N_2469,In_246,In_366);
or U2470 (N_2470,In_222,In_285);
nand U2471 (N_2471,In_344,In_559);
nor U2472 (N_2472,In_110,In_236);
nor U2473 (N_2473,In_905,In_983);
or U2474 (N_2474,In_965,In_426);
nand U2475 (N_2475,In_783,In_518);
nand U2476 (N_2476,In_317,In_364);
or U2477 (N_2477,In_688,In_2);
nor U2478 (N_2478,In_701,In_249);
and U2479 (N_2479,In_88,In_857);
or U2480 (N_2480,In_842,In_426);
nor U2481 (N_2481,In_337,In_560);
nand U2482 (N_2482,In_416,In_252);
nand U2483 (N_2483,In_867,In_938);
or U2484 (N_2484,In_691,In_648);
or U2485 (N_2485,In_887,In_665);
or U2486 (N_2486,In_389,In_942);
or U2487 (N_2487,In_895,In_622);
or U2488 (N_2488,In_143,In_224);
nand U2489 (N_2489,In_467,In_918);
or U2490 (N_2490,In_652,In_904);
nand U2491 (N_2491,In_780,In_785);
and U2492 (N_2492,In_465,In_250);
nand U2493 (N_2493,In_394,In_154);
and U2494 (N_2494,In_816,In_606);
or U2495 (N_2495,In_561,In_431);
or U2496 (N_2496,In_443,In_425);
xnor U2497 (N_2497,In_974,In_849);
or U2498 (N_2498,In_704,In_594);
and U2499 (N_2499,In_75,In_351);
and U2500 (N_2500,In_251,In_314);
or U2501 (N_2501,In_762,In_860);
or U2502 (N_2502,In_520,In_45);
or U2503 (N_2503,In_482,In_508);
and U2504 (N_2504,In_708,In_912);
nor U2505 (N_2505,In_449,In_819);
and U2506 (N_2506,In_892,In_215);
or U2507 (N_2507,In_985,In_212);
nand U2508 (N_2508,In_412,In_844);
nor U2509 (N_2509,In_809,In_923);
nor U2510 (N_2510,In_827,In_324);
or U2511 (N_2511,In_712,In_608);
and U2512 (N_2512,In_549,In_488);
or U2513 (N_2513,In_109,In_380);
nand U2514 (N_2514,In_726,In_772);
nand U2515 (N_2515,In_549,In_884);
nand U2516 (N_2516,In_910,In_179);
and U2517 (N_2517,In_507,In_880);
nand U2518 (N_2518,In_229,In_239);
and U2519 (N_2519,In_981,In_130);
and U2520 (N_2520,In_864,In_354);
nor U2521 (N_2521,In_477,In_909);
nor U2522 (N_2522,In_198,In_853);
nor U2523 (N_2523,In_273,In_366);
nor U2524 (N_2524,In_375,In_216);
and U2525 (N_2525,In_386,In_314);
and U2526 (N_2526,In_289,In_618);
nand U2527 (N_2527,In_341,In_824);
or U2528 (N_2528,In_445,In_110);
or U2529 (N_2529,In_276,In_518);
nor U2530 (N_2530,In_594,In_380);
or U2531 (N_2531,In_926,In_997);
or U2532 (N_2532,In_107,In_871);
or U2533 (N_2533,In_10,In_497);
nor U2534 (N_2534,In_607,In_540);
and U2535 (N_2535,In_601,In_577);
and U2536 (N_2536,In_313,In_720);
nor U2537 (N_2537,In_985,In_949);
and U2538 (N_2538,In_630,In_117);
and U2539 (N_2539,In_110,In_720);
nand U2540 (N_2540,In_33,In_147);
or U2541 (N_2541,In_850,In_113);
nor U2542 (N_2542,In_19,In_440);
and U2543 (N_2543,In_466,In_235);
and U2544 (N_2544,In_551,In_701);
or U2545 (N_2545,In_606,In_405);
nor U2546 (N_2546,In_190,In_114);
or U2547 (N_2547,In_831,In_111);
nand U2548 (N_2548,In_209,In_230);
nor U2549 (N_2549,In_134,In_423);
nand U2550 (N_2550,In_223,In_555);
or U2551 (N_2551,In_833,In_492);
and U2552 (N_2552,In_593,In_741);
and U2553 (N_2553,In_894,In_65);
and U2554 (N_2554,In_449,In_954);
and U2555 (N_2555,In_72,In_11);
and U2556 (N_2556,In_65,In_557);
nand U2557 (N_2557,In_260,In_817);
or U2558 (N_2558,In_62,In_508);
or U2559 (N_2559,In_686,In_514);
nor U2560 (N_2560,In_111,In_836);
and U2561 (N_2561,In_822,In_58);
and U2562 (N_2562,In_123,In_810);
and U2563 (N_2563,In_765,In_192);
and U2564 (N_2564,In_674,In_286);
or U2565 (N_2565,In_836,In_694);
nor U2566 (N_2566,In_164,In_73);
and U2567 (N_2567,In_417,In_679);
or U2568 (N_2568,In_823,In_192);
or U2569 (N_2569,In_474,In_551);
and U2570 (N_2570,In_419,In_732);
and U2571 (N_2571,In_626,In_314);
or U2572 (N_2572,In_698,In_678);
or U2573 (N_2573,In_878,In_739);
nor U2574 (N_2574,In_746,In_247);
nor U2575 (N_2575,In_855,In_901);
and U2576 (N_2576,In_155,In_509);
and U2577 (N_2577,In_556,In_288);
and U2578 (N_2578,In_910,In_202);
nor U2579 (N_2579,In_739,In_64);
and U2580 (N_2580,In_187,In_732);
nand U2581 (N_2581,In_841,In_944);
nand U2582 (N_2582,In_551,In_74);
nand U2583 (N_2583,In_431,In_740);
nand U2584 (N_2584,In_825,In_103);
xnor U2585 (N_2585,In_323,In_482);
nor U2586 (N_2586,In_59,In_560);
nand U2587 (N_2587,In_930,In_422);
nand U2588 (N_2588,In_140,In_822);
nor U2589 (N_2589,In_704,In_980);
and U2590 (N_2590,In_731,In_975);
nor U2591 (N_2591,In_53,In_318);
xor U2592 (N_2592,In_412,In_900);
and U2593 (N_2593,In_719,In_313);
and U2594 (N_2594,In_927,In_320);
nand U2595 (N_2595,In_222,In_606);
and U2596 (N_2596,In_433,In_192);
nand U2597 (N_2597,In_590,In_305);
nor U2598 (N_2598,In_391,In_557);
and U2599 (N_2599,In_539,In_187);
nand U2600 (N_2600,In_631,In_4);
or U2601 (N_2601,In_686,In_288);
nor U2602 (N_2602,In_568,In_77);
nor U2603 (N_2603,In_786,In_840);
and U2604 (N_2604,In_574,In_313);
or U2605 (N_2605,In_716,In_890);
and U2606 (N_2606,In_140,In_332);
and U2607 (N_2607,In_652,In_359);
nand U2608 (N_2608,In_659,In_881);
or U2609 (N_2609,In_75,In_528);
nand U2610 (N_2610,In_720,In_945);
nand U2611 (N_2611,In_366,In_916);
and U2612 (N_2612,In_639,In_575);
or U2613 (N_2613,In_117,In_832);
nand U2614 (N_2614,In_479,In_548);
nand U2615 (N_2615,In_218,In_236);
and U2616 (N_2616,In_683,In_740);
or U2617 (N_2617,In_220,In_408);
nand U2618 (N_2618,In_589,In_22);
nor U2619 (N_2619,In_905,In_329);
nor U2620 (N_2620,In_85,In_826);
and U2621 (N_2621,In_445,In_669);
nor U2622 (N_2622,In_738,In_343);
or U2623 (N_2623,In_500,In_959);
or U2624 (N_2624,In_92,In_730);
and U2625 (N_2625,In_546,In_967);
or U2626 (N_2626,In_115,In_181);
or U2627 (N_2627,In_884,In_305);
or U2628 (N_2628,In_178,In_768);
xor U2629 (N_2629,In_892,In_48);
nand U2630 (N_2630,In_558,In_444);
nor U2631 (N_2631,In_743,In_731);
xnor U2632 (N_2632,In_297,In_462);
and U2633 (N_2633,In_149,In_615);
or U2634 (N_2634,In_160,In_83);
or U2635 (N_2635,In_696,In_99);
nand U2636 (N_2636,In_190,In_775);
xor U2637 (N_2637,In_782,In_823);
and U2638 (N_2638,In_828,In_747);
nor U2639 (N_2639,In_748,In_742);
and U2640 (N_2640,In_840,In_6);
nand U2641 (N_2641,In_358,In_953);
and U2642 (N_2642,In_114,In_345);
and U2643 (N_2643,In_268,In_15);
and U2644 (N_2644,In_347,In_805);
nand U2645 (N_2645,In_842,In_54);
or U2646 (N_2646,In_700,In_663);
or U2647 (N_2647,In_942,In_999);
nand U2648 (N_2648,In_620,In_58);
nor U2649 (N_2649,In_411,In_398);
and U2650 (N_2650,In_729,In_15);
and U2651 (N_2651,In_878,In_382);
nand U2652 (N_2652,In_576,In_483);
nor U2653 (N_2653,In_634,In_236);
or U2654 (N_2654,In_886,In_29);
nand U2655 (N_2655,In_107,In_615);
nand U2656 (N_2656,In_747,In_420);
nand U2657 (N_2657,In_953,In_713);
and U2658 (N_2658,In_405,In_926);
nor U2659 (N_2659,In_961,In_286);
or U2660 (N_2660,In_474,In_535);
and U2661 (N_2661,In_764,In_922);
xnor U2662 (N_2662,In_790,In_249);
nand U2663 (N_2663,In_433,In_258);
or U2664 (N_2664,In_578,In_110);
xor U2665 (N_2665,In_710,In_838);
and U2666 (N_2666,In_764,In_872);
nand U2667 (N_2667,In_302,In_288);
nand U2668 (N_2668,In_41,In_288);
nand U2669 (N_2669,In_23,In_562);
nand U2670 (N_2670,In_264,In_530);
or U2671 (N_2671,In_48,In_74);
nand U2672 (N_2672,In_780,In_706);
and U2673 (N_2673,In_727,In_385);
and U2674 (N_2674,In_885,In_250);
or U2675 (N_2675,In_297,In_265);
or U2676 (N_2676,In_54,In_64);
nand U2677 (N_2677,In_256,In_938);
or U2678 (N_2678,In_965,In_683);
or U2679 (N_2679,In_541,In_821);
and U2680 (N_2680,In_871,In_497);
nand U2681 (N_2681,In_165,In_278);
and U2682 (N_2682,In_642,In_515);
nand U2683 (N_2683,In_769,In_181);
and U2684 (N_2684,In_623,In_42);
and U2685 (N_2685,In_7,In_120);
and U2686 (N_2686,In_811,In_905);
nand U2687 (N_2687,In_800,In_276);
nor U2688 (N_2688,In_565,In_171);
and U2689 (N_2689,In_52,In_345);
nor U2690 (N_2690,In_199,In_794);
nand U2691 (N_2691,In_151,In_84);
nor U2692 (N_2692,In_309,In_853);
nand U2693 (N_2693,In_50,In_822);
nor U2694 (N_2694,In_325,In_20);
nand U2695 (N_2695,In_198,In_708);
nor U2696 (N_2696,In_682,In_324);
and U2697 (N_2697,In_234,In_677);
nand U2698 (N_2698,In_175,In_591);
or U2699 (N_2699,In_261,In_857);
nand U2700 (N_2700,In_357,In_652);
and U2701 (N_2701,In_669,In_3);
nor U2702 (N_2702,In_161,In_444);
nand U2703 (N_2703,In_738,In_409);
nand U2704 (N_2704,In_30,In_345);
nand U2705 (N_2705,In_571,In_497);
or U2706 (N_2706,In_923,In_696);
and U2707 (N_2707,In_80,In_714);
or U2708 (N_2708,In_426,In_827);
or U2709 (N_2709,In_361,In_802);
nor U2710 (N_2710,In_151,In_189);
nor U2711 (N_2711,In_614,In_875);
nand U2712 (N_2712,In_747,In_530);
or U2713 (N_2713,In_470,In_418);
and U2714 (N_2714,In_78,In_512);
and U2715 (N_2715,In_440,In_43);
nor U2716 (N_2716,In_836,In_67);
nand U2717 (N_2717,In_882,In_260);
nand U2718 (N_2718,In_71,In_162);
or U2719 (N_2719,In_773,In_759);
and U2720 (N_2720,In_803,In_973);
and U2721 (N_2721,In_393,In_329);
nand U2722 (N_2722,In_274,In_138);
and U2723 (N_2723,In_74,In_929);
nand U2724 (N_2724,In_67,In_822);
nand U2725 (N_2725,In_205,In_307);
nand U2726 (N_2726,In_655,In_203);
nand U2727 (N_2727,In_817,In_382);
and U2728 (N_2728,In_495,In_826);
and U2729 (N_2729,In_259,In_99);
nor U2730 (N_2730,In_992,In_868);
and U2731 (N_2731,In_94,In_715);
and U2732 (N_2732,In_211,In_857);
nor U2733 (N_2733,In_338,In_453);
and U2734 (N_2734,In_413,In_821);
nand U2735 (N_2735,In_372,In_832);
or U2736 (N_2736,In_167,In_696);
or U2737 (N_2737,In_205,In_866);
or U2738 (N_2738,In_580,In_127);
nor U2739 (N_2739,In_909,In_296);
nor U2740 (N_2740,In_930,In_586);
and U2741 (N_2741,In_137,In_385);
nand U2742 (N_2742,In_684,In_313);
nand U2743 (N_2743,In_689,In_207);
and U2744 (N_2744,In_614,In_391);
or U2745 (N_2745,In_674,In_14);
nor U2746 (N_2746,In_811,In_264);
nand U2747 (N_2747,In_793,In_779);
and U2748 (N_2748,In_620,In_103);
nand U2749 (N_2749,In_138,In_944);
and U2750 (N_2750,In_973,In_665);
nor U2751 (N_2751,In_828,In_123);
nor U2752 (N_2752,In_44,In_193);
or U2753 (N_2753,In_428,In_627);
nand U2754 (N_2754,In_557,In_369);
and U2755 (N_2755,In_102,In_920);
or U2756 (N_2756,In_555,In_803);
and U2757 (N_2757,In_141,In_250);
and U2758 (N_2758,In_277,In_254);
and U2759 (N_2759,In_253,In_267);
nor U2760 (N_2760,In_65,In_139);
or U2761 (N_2761,In_305,In_856);
xnor U2762 (N_2762,In_814,In_337);
or U2763 (N_2763,In_885,In_384);
nand U2764 (N_2764,In_638,In_505);
and U2765 (N_2765,In_74,In_160);
and U2766 (N_2766,In_639,In_257);
nand U2767 (N_2767,In_349,In_708);
and U2768 (N_2768,In_326,In_189);
or U2769 (N_2769,In_947,In_108);
and U2770 (N_2770,In_800,In_827);
or U2771 (N_2771,In_198,In_155);
and U2772 (N_2772,In_447,In_406);
nand U2773 (N_2773,In_782,In_664);
and U2774 (N_2774,In_567,In_97);
xnor U2775 (N_2775,In_828,In_515);
nor U2776 (N_2776,In_828,In_28);
or U2777 (N_2777,In_760,In_179);
or U2778 (N_2778,In_516,In_710);
or U2779 (N_2779,In_577,In_397);
nor U2780 (N_2780,In_633,In_125);
nor U2781 (N_2781,In_399,In_878);
or U2782 (N_2782,In_506,In_65);
and U2783 (N_2783,In_343,In_447);
nor U2784 (N_2784,In_782,In_6);
nor U2785 (N_2785,In_249,In_669);
nand U2786 (N_2786,In_171,In_138);
and U2787 (N_2787,In_623,In_306);
nor U2788 (N_2788,In_398,In_539);
nand U2789 (N_2789,In_931,In_660);
and U2790 (N_2790,In_82,In_264);
or U2791 (N_2791,In_234,In_782);
and U2792 (N_2792,In_312,In_552);
and U2793 (N_2793,In_936,In_178);
nor U2794 (N_2794,In_135,In_481);
and U2795 (N_2795,In_539,In_769);
or U2796 (N_2796,In_275,In_340);
and U2797 (N_2797,In_502,In_18);
nor U2798 (N_2798,In_700,In_340);
nand U2799 (N_2799,In_403,In_565);
or U2800 (N_2800,In_807,In_571);
nor U2801 (N_2801,In_270,In_18);
nor U2802 (N_2802,In_340,In_139);
nor U2803 (N_2803,In_763,In_736);
and U2804 (N_2804,In_993,In_916);
or U2805 (N_2805,In_837,In_290);
or U2806 (N_2806,In_527,In_180);
nor U2807 (N_2807,In_701,In_687);
nor U2808 (N_2808,In_738,In_301);
and U2809 (N_2809,In_287,In_218);
or U2810 (N_2810,In_136,In_731);
nand U2811 (N_2811,In_458,In_799);
nor U2812 (N_2812,In_488,In_5);
nand U2813 (N_2813,In_969,In_25);
and U2814 (N_2814,In_730,In_544);
or U2815 (N_2815,In_433,In_268);
or U2816 (N_2816,In_35,In_785);
nand U2817 (N_2817,In_413,In_706);
and U2818 (N_2818,In_596,In_647);
and U2819 (N_2819,In_775,In_959);
and U2820 (N_2820,In_142,In_513);
and U2821 (N_2821,In_927,In_587);
nand U2822 (N_2822,In_161,In_145);
or U2823 (N_2823,In_758,In_340);
or U2824 (N_2824,In_585,In_938);
nand U2825 (N_2825,In_521,In_618);
or U2826 (N_2826,In_861,In_659);
or U2827 (N_2827,In_74,In_988);
nor U2828 (N_2828,In_746,In_497);
nand U2829 (N_2829,In_760,In_490);
and U2830 (N_2830,In_907,In_766);
nand U2831 (N_2831,In_301,In_618);
nor U2832 (N_2832,In_771,In_53);
and U2833 (N_2833,In_296,In_923);
nand U2834 (N_2834,In_921,In_166);
nand U2835 (N_2835,In_841,In_646);
and U2836 (N_2836,In_372,In_327);
nor U2837 (N_2837,In_583,In_718);
or U2838 (N_2838,In_841,In_329);
nand U2839 (N_2839,In_211,In_112);
or U2840 (N_2840,In_23,In_451);
and U2841 (N_2841,In_159,In_229);
nand U2842 (N_2842,In_256,In_549);
or U2843 (N_2843,In_812,In_838);
or U2844 (N_2844,In_142,In_51);
nand U2845 (N_2845,In_923,In_183);
or U2846 (N_2846,In_974,In_491);
nor U2847 (N_2847,In_769,In_716);
nand U2848 (N_2848,In_292,In_856);
nand U2849 (N_2849,In_59,In_833);
nor U2850 (N_2850,In_925,In_451);
or U2851 (N_2851,In_283,In_461);
and U2852 (N_2852,In_199,In_623);
nand U2853 (N_2853,In_979,In_405);
nand U2854 (N_2854,In_243,In_996);
nor U2855 (N_2855,In_338,In_393);
or U2856 (N_2856,In_330,In_699);
nand U2857 (N_2857,In_356,In_586);
and U2858 (N_2858,In_996,In_345);
or U2859 (N_2859,In_888,In_320);
or U2860 (N_2860,In_681,In_391);
nor U2861 (N_2861,In_632,In_958);
or U2862 (N_2862,In_686,In_692);
nand U2863 (N_2863,In_118,In_363);
or U2864 (N_2864,In_682,In_225);
or U2865 (N_2865,In_369,In_288);
and U2866 (N_2866,In_747,In_38);
or U2867 (N_2867,In_609,In_76);
nand U2868 (N_2868,In_429,In_169);
nor U2869 (N_2869,In_892,In_481);
nand U2870 (N_2870,In_682,In_875);
and U2871 (N_2871,In_42,In_590);
and U2872 (N_2872,In_267,In_411);
or U2873 (N_2873,In_739,In_74);
and U2874 (N_2874,In_817,In_151);
and U2875 (N_2875,In_8,In_759);
and U2876 (N_2876,In_583,In_889);
nor U2877 (N_2877,In_259,In_143);
or U2878 (N_2878,In_731,In_89);
or U2879 (N_2879,In_532,In_685);
or U2880 (N_2880,In_279,In_617);
nand U2881 (N_2881,In_729,In_35);
nand U2882 (N_2882,In_534,In_802);
and U2883 (N_2883,In_268,In_750);
and U2884 (N_2884,In_900,In_596);
nor U2885 (N_2885,In_584,In_475);
xnor U2886 (N_2886,In_954,In_760);
nor U2887 (N_2887,In_452,In_315);
nor U2888 (N_2888,In_374,In_539);
and U2889 (N_2889,In_302,In_836);
and U2890 (N_2890,In_368,In_535);
nor U2891 (N_2891,In_270,In_333);
nand U2892 (N_2892,In_315,In_81);
nor U2893 (N_2893,In_624,In_128);
nand U2894 (N_2894,In_775,In_61);
nor U2895 (N_2895,In_53,In_524);
nor U2896 (N_2896,In_100,In_728);
nor U2897 (N_2897,In_884,In_152);
nand U2898 (N_2898,In_409,In_427);
and U2899 (N_2899,In_715,In_84);
and U2900 (N_2900,In_386,In_616);
nand U2901 (N_2901,In_154,In_339);
nand U2902 (N_2902,In_153,In_289);
or U2903 (N_2903,In_509,In_99);
or U2904 (N_2904,In_699,In_421);
nand U2905 (N_2905,In_390,In_706);
nand U2906 (N_2906,In_14,In_660);
and U2907 (N_2907,In_22,In_134);
nand U2908 (N_2908,In_334,In_576);
and U2909 (N_2909,In_458,In_67);
nand U2910 (N_2910,In_460,In_257);
or U2911 (N_2911,In_758,In_574);
nor U2912 (N_2912,In_413,In_537);
and U2913 (N_2913,In_275,In_963);
nor U2914 (N_2914,In_858,In_168);
nand U2915 (N_2915,In_143,In_848);
or U2916 (N_2916,In_605,In_923);
nand U2917 (N_2917,In_6,In_596);
nand U2918 (N_2918,In_149,In_899);
nor U2919 (N_2919,In_830,In_910);
nor U2920 (N_2920,In_343,In_758);
and U2921 (N_2921,In_752,In_8);
nor U2922 (N_2922,In_508,In_341);
nor U2923 (N_2923,In_577,In_77);
and U2924 (N_2924,In_180,In_628);
nor U2925 (N_2925,In_598,In_267);
and U2926 (N_2926,In_523,In_992);
and U2927 (N_2927,In_930,In_866);
nand U2928 (N_2928,In_144,In_303);
or U2929 (N_2929,In_564,In_681);
nand U2930 (N_2930,In_748,In_689);
nor U2931 (N_2931,In_939,In_398);
nand U2932 (N_2932,In_573,In_130);
and U2933 (N_2933,In_773,In_974);
or U2934 (N_2934,In_874,In_300);
nand U2935 (N_2935,In_239,In_970);
xnor U2936 (N_2936,In_459,In_2);
and U2937 (N_2937,In_684,In_659);
nor U2938 (N_2938,In_889,In_248);
nand U2939 (N_2939,In_355,In_959);
nor U2940 (N_2940,In_709,In_153);
nor U2941 (N_2941,In_675,In_462);
nand U2942 (N_2942,In_13,In_448);
and U2943 (N_2943,In_983,In_916);
or U2944 (N_2944,In_337,In_431);
nor U2945 (N_2945,In_197,In_302);
or U2946 (N_2946,In_373,In_72);
xor U2947 (N_2947,In_926,In_564);
nor U2948 (N_2948,In_813,In_659);
or U2949 (N_2949,In_866,In_224);
nand U2950 (N_2950,In_273,In_943);
nor U2951 (N_2951,In_469,In_917);
or U2952 (N_2952,In_809,In_247);
or U2953 (N_2953,In_113,In_875);
or U2954 (N_2954,In_264,In_198);
or U2955 (N_2955,In_488,In_962);
nor U2956 (N_2956,In_470,In_922);
nand U2957 (N_2957,In_676,In_571);
or U2958 (N_2958,In_201,In_515);
or U2959 (N_2959,In_679,In_828);
or U2960 (N_2960,In_890,In_522);
nor U2961 (N_2961,In_518,In_600);
nor U2962 (N_2962,In_313,In_694);
nor U2963 (N_2963,In_10,In_628);
nand U2964 (N_2964,In_500,In_803);
and U2965 (N_2965,In_184,In_876);
nand U2966 (N_2966,In_913,In_710);
and U2967 (N_2967,In_826,In_343);
and U2968 (N_2968,In_386,In_488);
or U2969 (N_2969,In_805,In_268);
nand U2970 (N_2970,In_339,In_16);
or U2971 (N_2971,In_343,In_511);
and U2972 (N_2972,In_182,In_954);
nor U2973 (N_2973,In_176,In_291);
nor U2974 (N_2974,In_237,In_342);
nor U2975 (N_2975,In_680,In_141);
nand U2976 (N_2976,In_144,In_992);
nand U2977 (N_2977,In_186,In_955);
and U2978 (N_2978,In_139,In_69);
and U2979 (N_2979,In_717,In_75);
and U2980 (N_2980,In_652,In_546);
nand U2981 (N_2981,In_170,In_327);
and U2982 (N_2982,In_846,In_330);
or U2983 (N_2983,In_433,In_530);
or U2984 (N_2984,In_102,In_978);
and U2985 (N_2985,In_480,In_951);
nor U2986 (N_2986,In_428,In_793);
nor U2987 (N_2987,In_115,In_696);
nor U2988 (N_2988,In_846,In_650);
nand U2989 (N_2989,In_539,In_323);
nor U2990 (N_2990,In_169,In_991);
and U2991 (N_2991,In_893,In_29);
nand U2992 (N_2992,In_758,In_296);
nand U2993 (N_2993,In_597,In_90);
nor U2994 (N_2994,In_701,In_227);
nor U2995 (N_2995,In_64,In_409);
nand U2996 (N_2996,In_910,In_530);
or U2997 (N_2997,In_981,In_947);
or U2998 (N_2998,In_61,In_451);
nor U2999 (N_2999,In_397,In_757);
and U3000 (N_3000,In_670,In_935);
nand U3001 (N_3001,In_86,In_964);
and U3002 (N_3002,In_26,In_213);
nor U3003 (N_3003,In_126,In_559);
or U3004 (N_3004,In_261,In_738);
nand U3005 (N_3005,In_970,In_238);
nor U3006 (N_3006,In_156,In_887);
nand U3007 (N_3007,In_890,In_117);
nand U3008 (N_3008,In_122,In_798);
nand U3009 (N_3009,In_796,In_795);
or U3010 (N_3010,In_509,In_514);
nand U3011 (N_3011,In_152,In_204);
nor U3012 (N_3012,In_381,In_336);
nor U3013 (N_3013,In_562,In_782);
nand U3014 (N_3014,In_257,In_726);
nor U3015 (N_3015,In_637,In_407);
nand U3016 (N_3016,In_255,In_409);
nand U3017 (N_3017,In_624,In_316);
or U3018 (N_3018,In_341,In_635);
nor U3019 (N_3019,In_580,In_731);
or U3020 (N_3020,In_734,In_617);
nand U3021 (N_3021,In_27,In_875);
and U3022 (N_3022,In_288,In_78);
or U3023 (N_3023,In_188,In_99);
and U3024 (N_3024,In_580,In_685);
or U3025 (N_3025,In_445,In_120);
nor U3026 (N_3026,In_242,In_317);
and U3027 (N_3027,In_15,In_411);
and U3028 (N_3028,In_261,In_516);
nor U3029 (N_3029,In_705,In_218);
nand U3030 (N_3030,In_526,In_426);
nand U3031 (N_3031,In_925,In_975);
and U3032 (N_3032,In_848,In_529);
and U3033 (N_3033,In_120,In_812);
or U3034 (N_3034,In_578,In_840);
or U3035 (N_3035,In_827,In_147);
nor U3036 (N_3036,In_782,In_817);
and U3037 (N_3037,In_277,In_996);
nor U3038 (N_3038,In_336,In_878);
nand U3039 (N_3039,In_321,In_833);
or U3040 (N_3040,In_615,In_987);
nor U3041 (N_3041,In_661,In_270);
or U3042 (N_3042,In_853,In_424);
nand U3043 (N_3043,In_90,In_764);
and U3044 (N_3044,In_78,In_639);
and U3045 (N_3045,In_220,In_617);
nand U3046 (N_3046,In_592,In_422);
nor U3047 (N_3047,In_783,In_186);
and U3048 (N_3048,In_579,In_262);
nand U3049 (N_3049,In_479,In_537);
nand U3050 (N_3050,In_700,In_889);
nor U3051 (N_3051,In_494,In_769);
or U3052 (N_3052,In_63,In_854);
or U3053 (N_3053,In_190,In_384);
nand U3054 (N_3054,In_697,In_671);
nand U3055 (N_3055,In_808,In_895);
or U3056 (N_3056,In_410,In_535);
and U3057 (N_3057,In_887,In_283);
nand U3058 (N_3058,In_672,In_832);
nor U3059 (N_3059,In_231,In_497);
nor U3060 (N_3060,In_557,In_735);
and U3061 (N_3061,In_207,In_656);
nor U3062 (N_3062,In_618,In_294);
or U3063 (N_3063,In_346,In_562);
nand U3064 (N_3064,In_143,In_127);
nand U3065 (N_3065,In_868,In_27);
and U3066 (N_3066,In_366,In_557);
and U3067 (N_3067,In_123,In_674);
nor U3068 (N_3068,In_27,In_671);
nand U3069 (N_3069,In_86,In_699);
nor U3070 (N_3070,In_947,In_337);
nor U3071 (N_3071,In_405,In_415);
nor U3072 (N_3072,In_961,In_839);
nor U3073 (N_3073,In_737,In_153);
or U3074 (N_3074,In_915,In_898);
nand U3075 (N_3075,In_670,In_983);
and U3076 (N_3076,In_832,In_794);
nor U3077 (N_3077,In_318,In_292);
nor U3078 (N_3078,In_917,In_101);
nor U3079 (N_3079,In_437,In_377);
or U3080 (N_3080,In_112,In_264);
nand U3081 (N_3081,In_340,In_818);
nor U3082 (N_3082,In_403,In_172);
nand U3083 (N_3083,In_411,In_720);
and U3084 (N_3084,In_939,In_425);
or U3085 (N_3085,In_279,In_601);
nor U3086 (N_3086,In_674,In_697);
nand U3087 (N_3087,In_662,In_787);
or U3088 (N_3088,In_255,In_821);
or U3089 (N_3089,In_911,In_858);
and U3090 (N_3090,In_564,In_805);
nand U3091 (N_3091,In_482,In_806);
nand U3092 (N_3092,In_800,In_182);
nor U3093 (N_3093,In_758,In_3);
and U3094 (N_3094,In_456,In_383);
or U3095 (N_3095,In_516,In_326);
or U3096 (N_3096,In_213,In_121);
and U3097 (N_3097,In_637,In_141);
nand U3098 (N_3098,In_661,In_712);
nand U3099 (N_3099,In_78,In_590);
and U3100 (N_3100,In_38,In_953);
and U3101 (N_3101,In_978,In_345);
nor U3102 (N_3102,In_769,In_721);
nand U3103 (N_3103,In_358,In_259);
and U3104 (N_3104,In_725,In_152);
or U3105 (N_3105,In_746,In_951);
nand U3106 (N_3106,In_194,In_179);
nand U3107 (N_3107,In_217,In_567);
nand U3108 (N_3108,In_869,In_525);
nor U3109 (N_3109,In_245,In_896);
and U3110 (N_3110,In_860,In_338);
nor U3111 (N_3111,In_32,In_898);
nand U3112 (N_3112,In_919,In_763);
nand U3113 (N_3113,In_844,In_830);
nand U3114 (N_3114,In_762,In_368);
or U3115 (N_3115,In_182,In_96);
nor U3116 (N_3116,In_41,In_293);
or U3117 (N_3117,In_359,In_192);
or U3118 (N_3118,In_520,In_510);
and U3119 (N_3119,In_17,In_761);
and U3120 (N_3120,In_654,In_751);
nor U3121 (N_3121,In_0,In_239);
or U3122 (N_3122,In_259,In_228);
or U3123 (N_3123,In_548,In_871);
nand U3124 (N_3124,In_179,In_49);
or U3125 (N_3125,In_615,In_913);
and U3126 (N_3126,In_194,In_814);
nor U3127 (N_3127,In_223,In_647);
nand U3128 (N_3128,In_836,In_841);
nand U3129 (N_3129,In_148,In_603);
and U3130 (N_3130,In_357,In_670);
nand U3131 (N_3131,In_376,In_214);
or U3132 (N_3132,In_189,In_627);
nand U3133 (N_3133,In_938,In_311);
nand U3134 (N_3134,In_78,In_145);
or U3135 (N_3135,In_103,In_907);
and U3136 (N_3136,In_215,In_532);
nand U3137 (N_3137,In_507,In_196);
nand U3138 (N_3138,In_543,In_259);
nand U3139 (N_3139,In_873,In_867);
nor U3140 (N_3140,In_25,In_670);
nand U3141 (N_3141,In_753,In_717);
and U3142 (N_3142,In_285,In_596);
and U3143 (N_3143,In_775,In_395);
and U3144 (N_3144,In_665,In_163);
and U3145 (N_3145,In_213,In_823);
nor U3146 (N_3146,In_906,In_63);
or U3147 (N_3147,In_20,In_316);
nor U3148 (N_3148,In_519,In_125);
or U3149 (N_3149,In_658,In_678);
nor U3150 (N_3150,In_681,In_7);
nor U3151 (N_3151,In_972,In_629);
nand U3152 (N_3152,In_783,In_538);
and U3153 (N_3153,In_277,In_832);
or U3154 (N_3154,In_699,In_559);
nor U3155 (N_3155,In_939,In_404);
nand U3156 (N_3156,In_715,In_49);
nand U3157 (N_3157,In_799,In_217);
nand U3158 (N_3158,In_197,In_734);
or U3159 (N_3159,In_554,In_565);
nand U3160 (N_3160,In_287,In_784);
or U3161 (N_3161,In_27,In_30);
nand U3162 (N_3162,In_248,In_392);
and U3163 (N_3163,In_436,In_980);
nor U3164 (N_3164,In_677,In_357);
or U3165 (N_3165,In_309,In_105);
nand U3166 (N_3166,In_143,In_79);
nor U3167 (N_3167,In_156,In_550);
nand U3168 (N_3168,In_383,In_535);
nand U3169 (N_3169,In_390,In_986);
xnor U3170 (N_3170,In_935,In_977);
or U3171 (N_3171,In_647,In_233);
nand U3172 (N_3172,In_304,In_431);
or U3173 (N_3173,In_707,In_970);
nor U3174 (N_3174,In_76,In_13);
or U3175 (N_3175,In_388,In_796);
or U3176 (N_3176,In_369,In_908);
or U3177 (N_3177,In_826,In_268);
nand U3178 (N_3178,In_724,In_471);
nand U3179 (N_3179,In_33,In_851);
nor U3180 (N_3180,In_76,In_18);
or U3181 (N_3181,In_120,In_700);
or U3182 (N_3182,In_9,In_638);
or U3183 (N_3183,In_724,In_180);
nand U3184 (N_3184,In_244,In_339);
nand U3185 (N_3185,In_875,In_554);
nor U3186 (N_3186,In_147,In_384);
or U3187 (N_3187,In_519,In_108);
and U3188 (N_3188,In_853,In_930);
or U3189 (N_3189,In_577,In_553);
and U3190 (N_3190,In_479,In_945);
or U3191 (N_3191,In_992,In_332);
or U3192 (N_3192,In_391,In_862);
nand U3193 (N_3193,In_248,In_852);
or U3194 (N_3194,In_187,In_259);
nor U3195 (N_3195,In_35,In_496);
nand U3196 (N_3196,In_51,In_864);
or U3197 (N_3197,In_784,In_526);
and U3198 (N_3198,In_383,In_492);
or U3199 (N_3199,In_721,In_164);
and U3200 (N_3200,In_14,In_312);
or U3201 (N_3201,In_148,In_713);
nor U3202 (N_3202,In_642,In_695);
and U3203 (N_3203,In_33,In_737);
nand U3204 (N_3204,In_628,In_144);
nand U3205 (N_3205,In_803,In_782);
nand U3206 (N_3206,In_760,In_551);
nor U3207 (N_3207,In_480,In_637);
xnor U3208 (N_3208,In_298,In_259);
or U3209 (N_3209,In_877,In_395);
nor U3210 (N_3210,In_47,In_18);
or U3211 (N_3211,In_702,In_946);
nand U3212 (N_3212,In_949,In_386);
nor U3213 (N_3213,In_79,In_387);
or U3214 (N_3214,In_761,In_527);
and U3215 (N_3215,In_765,In_145);
nor U3216 (N_3216,In_828,In_480);
nand U3217 (N_3217,In_197,In_401);
and U3218 (N_3218,In_920,In_829);
and U3219 (N_3219,In_304,In_948);
or U3220 (N_3220,In_612,In_536);
nand U3221 (N_3221,In_834,In_863);
and U3222 (N_3222,In_208,In_521);
or U3223 (N_3223,In_566,In_637);
and U3224 (N_3224,In_918,In_706);
or U3225 (N_3225,In_129,In_53);
and U3226 (N_3226,In_201,In_582);
and U3227 (N_3227,In_65,In_300);
nand U3228 (N_3228,In_322,In_628);
nor U3229 (N_3229,In_320,In_89);
nor U3230 (N_3230,In_990,In_699);
nor U3231 (N_3231,In_21,In_510);
nand U3232 (N_3232,In_145,In_417);
nand U3233 (N_3233,In_723,In_287);
nand U3234 (N_3234,In_428,In_519);
or U3235 (N_3235,In_339,In_978);
nand U3236 (N_3236,In_408,In_551);
nor U3237 (N_3237,In_400,In_114);
and U3238 (N_3238,In_431,In_420);
nor U3239 (N_3239,In_999,In_594);
nor U3240 (N_3240,In_476,In_359);
nand U3241 (N_3241,In_595,In_490);
nand U3242 (N_3242,In_146,In_112);
or U3243 (N_3243,In_97,In_398);
nor U3244 (N_3244,In_384,In_406);
nor U3245 (N_3245,In_114,In_561);
nor U3246 (N_3246,In_953,In_858);
and U3247 (N_3247,In_316,In_682);
nand U3248 (N_3248,In_862,In_546);
nand U3249 (N_3249,In_506,In_585);
or U3250 (N_3250,In_489,In_947);
or U3251 (N_3251,In_830,In_707);
and U3252 (N_3252,In_187,In_301);
nand U3253 (N_3253,In_69,In_868);
or U3254 (N_3254,In_931,In_564);
and U3255 (N_3255,In_218,In_680);
nand U3256 (N_3256,In_856,In_563);
and U3257 (N_3257,In_987,In_212);
nor U3258 (N_3258,In_711,In_347);
and U3259 (N_3259,In_416,In_318);
or U3260 (N_3260,In_743,In_155);
nor U3261 (N_3261,In_60,In_880);
nor U3262 (N_3262,In_204,In_347);
nand U3263 (N_3263,In_276,In_929);
or U3264 (N_3264,In_62,In_39);
nand U3265 (N_3265,In_945,In_961);
nand U3266 (N_3266,In_123,In_17);
and U3267 (N_3267,In_475,In_870);
and U3268 (N_3268,In_856,In_743);
and U3269 (N_3269,In_924,In_75);
or U3270 (N_3270,In_938,In_109);
and U3271 (N_3271,In_279,In_71);
or U3272 (N_3272,In_49,In_807);
or U3273 (N_3273,In_964,In_732);
nor U3274 (N_3274,In_899,In_181);
or U3275 (N_3275,In_731,In_475);
and U3276 (N_3276,In_531,In_54);
nand U3277 (N_3277,In_481,In_770);
or U3278 (N_3278,In_887,In_3);
nor U3279 (N_3279,In_555,In_462);
or U3280 (N_3280,In_148,In_944);
nor U3281 (N_3281,In_552,In_750);
or U3282 (N_3282,In_392,In_38);
nor U3283 (N_3283,In_218,In_747);
nor U3284 (N_3284,In_717,In_159);
nor U3285 (N_3285,In_733,In_303);
nand U3286 (N_3286,In_646,In_614);
nand U3287 (N_3287,In_401,In_178);
nor U3288 (N_3288,In_232,In_848);
and U3289 (N_3289,In_653,In_257);
and U3290 (N_3290,In_981,In_487);
nand U3291 (N_3291,In_328,In_6);
nand U3292 (N_3292,In_371,In_105);
or U3293 (N_3293,In_701,In_763);
nor U3294 (N_3294,In_575,In_736);
or U3295 (N_3295,In_257,In_301);
or U3296 (N_3296,In_114,In_704);
and U3297 (N_3297,In_982,In_45);
and U3298 (N_3298,In_939,In_77);
nor U3299 (N_3299,In_613,In_511);
nor U3300 (N_3300,In_57,In_991);
nand U3301 (N_3301,In_631,In_525);
nand U3302 (N_3302,In_136,In_561);
and U3303 (N_3303,In_212,In_785);
and U3304 (N_3304,In_568,In_52);
nor U3305 (N_3305,In_876,In_955);
or U3306 (N_3306,In_153,In_536);
nor U3307 (N_3307,In_158,In_186);
nor U3308 (N_3308,In_599,In_425);
nor U3309 (N_3309,In_210,In_165);
or U3310 (N_3310,In_921,In_602);
nor U3311 (N_3311,In_275,In_488);
nand U3312 (N_3312,In_437,In_469);
or U3313 (N_3313,In_421,In_404);
nor U3314 (N_3314,In_529,In_18);
or U3315 (N_3315,In_398,In_962);
xnor U3316 (N_3316,In_732,In_463);
nor U3317 (N_3317,In_227,In_275);
or U3318 (N_3318,In_170,In_981);
nor U3319 (N_3319,In_229,In_815);
nor U3320 (N_3320,In_560,In_12);
and U3321 (N_3321,In_951,In_276);
and U3322 (N_3322,In_649,In_483);
and U3323 (N_3323,In_52,In_411);
nor U3324 (N_3324,In_659,In_991);
and U3325 (N_3325,In_874,In_282);
or U3326 (N_3326,In_799,In_459);
and U3327 (N_3327,In_886,In_460);
or U3328 (N_3328,In_973,In_524);
or U3329 (N_3329,In_34,In_226);
nand U3330 (N_3330,In_65,In_428);
and U3331 (N_3331,In_672,In_627);
nor U3332 (N_3332,In_102,In_868);
or U3333 (N_3333,In_709,In_688);
and U3334 (N_3334,In_158,In_993);
nand U3335 (N_3335,In_82,In_49);
and U3336 (N_3336,In_510,In_182);
and U3337 (N_3337,In_996,In_981);
nor U3338 (N_3338,In_253,In_389);
and U3339 (N_3339,In_777,In_367);
nand U3340 (N_3340,In_468,In_832);
and U3341 (N_3341,In_996,In_515);
or U3342 (N_3342,In_814,In_748);
nand U3343 (N_3343,In_266,In_842);
and U3344 (N_3344,In_819,In_13);
or U3345 (N_3345,In_145,In_63);
and U3346 (N_3346,In_957,In_119);
nor U3347 (N_3347,In_891,In_616);
nand U3348 (N_3348,In_963,In_677);
nand U3349 (N_3349,In_359,In_132);
nand U3350 (N_3350,In_635,In_431);
nand U3351 (N_3351,In_250,In_491);
and U3352 (N_3352,In_750,In_811);
and U3353 (N_3353,In_280,In_440);
nor U3354 (N_3354,In_740,In_711);
or U3355 (N_3355,In_888,In_67);
nand U3356 (N_3356,In_207,In_831);
and U3357 (N_3357,In_606,In_885);
and U3358 (N_3358,In_96,In_784);
or U3359 (N_3359,In_209,In_122);
or U3360 (N_3360,In_331,In_407);
nor U3361 (N_3361,In_101,In_902);
nand U3362 (N_3362,In_81,In_638);
nand U3363 (N_3363,In_412,In_141);
and U3364 (N_3364,In_678,In_680);
nor U3365 (N_3365,In_218,In_173);
nand U3366 (N_3366,In_951,In_19);
nor U3367 (N_3367,In_447,In_955);
and U3368 (N_3368,In_359,In_622);
nand U3369 (N_3369,In_110,In_596);
nor U3370 (N_3370,In_702,In_894);
nand U3371 (N_3371,In_773,In_991);
and U3372 (N_3372,In_151,In_58);
nand U3373 (N_3373,In_351,In_922);
nor U3374 (N_3374,In_969,In_637);
and U3375 (N_3375,In_128,In_626);
or U3376 (N_3376,In_868,In_427);
and U3377 (N_3377,In_134,In_352);
nor U3378 (N_3378,In_704,In_984);
and U3379 (N_3379,In_506,In_281);
nand U3380 (N_3380,In_468,In_81);
and U3381 (N_3381,In_422,In_601);
or U3382 (N_3382,In_573,In_186);
nand U3383 (N_3383,In_3,In_420);
nor U3384 (N_3384,In_312,In_363);
nand U3385 (N_3385,In_400,In_403);
xor U3386 (N_3386,In_441,In_471);
nand U3387 (N_3387,In_655,In_856);
and U3388 (N_3388,In_934,In_395);
and U3389 (N_3389,In_916,In_318);
nor U3390 (N_3390,In_851,In_393);
or U3391 (N_3391,In_726,In_74);
or U3392 (N_3392,In_31,In_245);
nand U3393 (N_3393,In_279,In_147);
nor U3394 (N_3394,In_116,In_722);
nand U3395 (N_3395,In_656,In_190);
xor U3396 (N_3396,In_792,In_684);
nand U3397 (N_3397,In_913,In_423);
nor U3398 (N_3398,In_323,In_279);
nand U3399 (N_3399,In_192,In_247);
nor U3400 (N_3400,In_619,In_995);
and U3401 (N_3401,In_84,In_609);
and U3402 (N_3402,In_791,In_55);
and U3403 (N_3403,In_525,In_276);
nor U3404 (N_3404,In_755,In_540);
and U3405 (N_3405,In_669,In_901);
and U3406 (N_3406,In_934,In_269);
and U3407 (N_3407,In_765,In_962);
nand U3408 (N_3408,In_384,In_961);
nand U3409 (N_3409,In_115,In_523);
and U3410 (N_3410,In_401,In_379);
or U3411 (N_3411,In_467,In_682);
nand U3412 (N_3412,In_866,In_129);
xnor U3413 (N_3413,In_363,In_542);
or U3414 (N_3414,In_832,In_66);
or U3415 (N_3415,In_450,In_955);
or U3416 (N_3416,In_643,In_781);
nor U3417 (N_3417,In_416,In_738);
or U3418 (N_3418,In_482,In_295);
nand U3419 (N_3419,In_236,In_585);
and U3420 (N_3420,In_723,In_805);
nor U3421 (N_3421,In_851,In_21);
and U3422 (N_3422,In_230,In_234);
nor U3423 (N_3423,In_595,In_124);
nand U3424 (N_3424,In_415,In_963);
or U3425 (N_3425,In_198,In_953);
or U3426 (N_3426,In_723,In_931);
and U3427 (N_3427,In_607,In_541);
nand U3428 (N_3428,In_324,In_159);
or U3429 (N_3429,In_359,In_672);
nand U3430 (N_3430,In_654,In_260);
nor U3431 (N_3431,In_861,In_820);
or U3432 (N_3432,In_779,In_747);
and U3433 (N_3433,In_532,In_698);
and U3434 (N_3434,In_779,In_356);
nand U3435 (N_3435,In_744,In_156);
nand U3436 (N_3436,In_601,In_386);
or U3437 (N_3437,In_410,In_159);
nor U3438 (N_3438,In_652,In_202);
or U3439 (N_3439,In_199,In_717);
or U3440 (N_3440,In_376,In_778);
and U3441 (N_3441,In_383,In_316);
and U3442 (N_3442,In_859,In_473);
and U3443 (N_3443,In_388,In_612);
nand U3444 (N_3444,In_593,In_820);
and U3445 (N_3445,In_204,In_743);
or U3446 (N_3446,In_803,In_644);
nand U3447 (N_3447,In_745,In_882);
nand U3448 (N_3448,In_25,In_841);
or U3449 (N_3449,In_185,In_802);
nand U3450 (N_3450,In_15,In_17);
nor U3451 (N_3451,In_464,In_823);
nor U3452 (N_3452,In_422,In_112);
or U3453 (N_3453,In_583,In_860);
and U3454 (N_3454,In_682,In_490);
and U3455 (N_3455,In_971,In_393);
and U3456 (N_3456,In_501,In_259);
nor U3457 (N_3457,In_729,In_86);
and U3458 (N_3458,In_242,In_415);
nand U3459 (N_3459,In_273,In_352);
or U3460 (N_3460,In_241,In_409);
nand U3461 (N_3461,In_351,In_649);
nand U3462 (N_3462,In_225,In_736);
and U3463 (N_3463,In_156,In_981);
and U3464 (N_3464,In_959,In_508);
and U3465 (N_3465,In_863,In_334);
or U3466 (N_3466,In_776,In_685);
and U3467 (N_3467,In_100,In_476);
or U3468 (N_3468,In_487,In_666);
nor U3469 (N_3469,In_1,In_284);
and U3470 (N_3470,In_695,In_710);
or U3471 (N_3471,In_53,In_566);
nor U3472 (N_3472,In_610,In_704);
or U3473 (N_3473,In_155,In_361);
nand U3474 (N_3474,In_375,In_51);
or U3475 (N_3475,In_6,In_413);
nor U3476 (N_3476,In_219,In_138);
nand U3477 (N_3477,In_107,In_848);
nor U3478 (N_3478,In_191,In_382);
xnor U3479 (N_3479,In_357,In_591);
nand U3480 (N_3480,In_176,In_827);
and U3481 (N_3481,In_352,In_486);
nand U3482 (N_3482,In_42,In_556);
or U3483 (N_3483,In_628,In_444);
or U3484 (N_3484,In_0,In_414);
or U3485 (N_3485,In_266,In_506);
nor U3486 (N_3486,In_139,In_953);
nor U3487 (N_3487,In_770,In_465);
or U3488 (N_3488,In_999,In_737);
and U3489 (N_3489,In_958,In_228);
nor U3490 (N_3490,In_717,In_228);
nand U3491 (N_3491,In_885,In_959);
or U3492 (N_3492,In_51,In_97);
and U3493 (N_3493,In_1,In_171);
nor U3494 (N_3494,In_420,In_939);
nand U3495 (N_3495,In_444,In_269);
nor U3496 (N_3496,In_242,In_156);
or U3497 (N_3497,In_454,In_45);
nor U3498 (N_3498,In_993,In_427);
and U3499 (N_3499,In_797,In_251);
and U3500 (N_3500,In_425,In_389);
nor U3501 (N_3501,In_268,In_759);
and U3502 (N_3502,In_598,In_572);
or U3503 (N_3503,In_632,In_876);
nor U3504 (N_3504,In_869,In_624);
nand U3505 (N_3505,In_515,In_494);
nor U3506 (N_3506,In_4,In_472);
and U3507 (N_3507,In_116,In_657);
nand U3508 (N_3508,In_58,In_924);
nand U3509 (N_3509,In_883,In_884);
nand U3510 (N_3510,In_6,In_301);
nand U3511 (N_3511,In_48,In_735);
nand U3512 (N_3512,In_185,In_463);
or U3513 (N_3513,In_431,In_761);
or U3514 (N_3514,In_881,In_429);
nor U3515 (N_3515,In_488,In_487);
nor U3516 (N_3516,In_730,In_243);
or U3517 (N_3517,In_222,In_577);
nand U3518 (N_3518,In_436,In_310);
or U3519 (N_3519,In_595,In_526);
and U3520 (N_3520,In_473,In_836);
nor U3521 (N_3521,In_73,In_437);
or U3522 (N_3522,In_211,In_698);
or U3523 (N_3523,In_515,In_798);
nor U3524 (N_3524,In_541,In_711);
nor U3525 (N_3525,In_34,In_147);
nor U3526 (N_3526,In_568,In_367);
or U3527 (N_3527,In_47,In_124);
nor U3528 (N_3528,In_451,In_223);
nor U3529 (N_3529,In_262,In_222);
or U3530 (N_3530,In_564,In_789);
and U3531 (N_3531,In_285,In_636);
nand U3532 (N_3532,In_91,In_995);
or U3533 (N_3533,In_337,In_304);
and U3534 (N_3534,In_373,In_198);
nand U3535 (N_3535,In_153,In_679);
nor U3536 (N_3536,In_237,In_648);
nand U3537 (N_3537,In_688,In_752);
or U3538 (N_3538,In_905,In_280);
and U3539 (N_3539,In_383,In_873);
nand U3540 (N_3540,In_48,In_151);
and U3541 (N_3541,In_132,In_444);
and U3542 (N_3542,In_375,In_256);
nor U3543 (N_3543,In_868,In_83);
or U3544 (N_3544,In_782,In_357);
nand U3545 (N_3545,In_362,In_87);
and U3546 (N_3546,In_213,In_633);
and U3547 (N_3547,In_78,In_268);
nor U3548 (N_3548,In_281,In_37);
nor U3549 (N_3549,In_709,In_776);
nor U3550 (N_3550,In_112,In_312);
nand U3551 (N_3551,In_844,In_396);
and U3552 (N_3552,In_50,In_470);
nor U3553 (N_3553,In_332,In_184);
and U3554 (N_3554,In_546,In_475);
nor U3555 (N_3555,In_801,In_170);
and U3556 (N_3556,In_598,In_656);
nor U3557 (N_3557,In_235,In_334);
nor U3558 (N_3558,In_967,In_811);
nand U3559 (N_3559,In_397,In_792);
or U3560 (N_3560,In_277,In_248);
or U3561 (N_3561,In_407,In_761);
nand U3562 (N_3562,In_101,In_883);
and U3563 (N_3563,In_541,In_0);
nor U3564 (N_3564,In_287,In_224);
nor U3565 (N_3565,In_691,In_289);
nor U3566 (N_3566,In_900,In_180);
nand U3567 (N_3567,In_12,In_422);
and U3568 (N_3568,In_911,In_624);
nand U3569 (N_3569,In_406,In_938);
or U3570 (N_3570,In_70,In_34);
nand U3571 (N_3571,In_294,In_954);
or U3572 (N_3572,In_589,In_387);
nor U3573 (N_3573,In_969,In_874);
and U3574 (N_3574,In_957,In_636);
nand U3575 (N_3575,In_892,In_6);
nor U3576 (N_3576,In_388,In_978);
and U3577 (N_3577,In_10,In_16);
nor U3578 (N_3578,In_980,In_346);
or U3579 (N_3579,In_240,In_830);
or U3580 (N_3580,In_81,In_574);
and U3581 (N_3581,In_430,In_405);
nor U3582 (N_3582,In_529,In_488);
nand U3583 (N_3583,In_507,In_976);
nor U3584 (N_3584,In_593,In_412);
nor U3585 (N_3585,In_455,In_105);
nor U3586 (N_3586,In_985,In_243);
and U3587 (N_3587,In_200,In_810);
nor U3588 (N_3588,In_817,In_811);
and U3589 (N_3589,In_361,In_341);
nand U3590 (N_3590,In_277,In_143);
nand U3591 (N_3591,In_177,In_387);
or U3592 (N_3592,In_109,In_801);
and U3593 (N_3593,In_537,In_637);
nor U3594 (N_3594,In_134,In_519);
or U3595 (N_3595,In_234,In_410);
or U3596 (N_3596,In_587,In_219);
and U3597 (N_3597,In_565,In_59);
or U3598 (N_3598,In_160,In_585);
nand U3599 (N_3599,In_741,In_828);
nor U3600 (N_3600,In_690,In_364);
nand U3601 (N_3601,In_679,In_553);
nand U3602 (N_3602,In_150,In_329);
or U3603 (N_3603,In_344,In_462);
and U3604 (N_3604,In_616,In_681);
or U3605 (N_3605,In_809,In_420);
and U3606 (N_3606,In_210,In_826);
and U3607 (N_3607,In_954,In_884);
and U3608 (N_3608,In_564,In_405);
and U3609 (N_3609,In_742,In_501);
nor U3610 (N_3610,In_106,In_49);
nand U3611 (N_3611,In_792,In_85);
nor U3612 (N_3612,In_318,In_127);
and U3613 (N_3613,In_341,In_906);
nand U3614 (N_3614,In_77,In_428);
and U3615 (N_3615,In_788,In_440);
and U3616 (N_3616,In_270,In_23);
and U3617 (N_3617,In_681,In_552);
and U3618 (N_3618,In_272,In_693);
nor U3619 (N_3619,In_362,In_216);
and U3620 (N_3620,In_257,In_823);
nor U3621 (N_3621,In_1,In_257);
nand U3622 (N_3622,In_838,In_744);
and U3623 (N_3623,In_612,In_356);
nor U3624 (N_3624,In_410,In_331);
nand U3625 (N_3625,In_200,In_951);
or U3626 (N_3626,In_310,In_429);
nand U3627 (N_3627,In_808,In_334);
nand U3628 (N_3628,In_495,In_498);
nand U3629 (N_3629,In_824,In_852);
nand U3630 (N_3630,In_683,In_999);
or U3631 (N_3631,In_916,In_57);
nand U3632 (N_3632,In_586,In_577);
or U3633 (N_3633,In_14,In_47);
and U3634 (N_3634,In_75,In_875);
and U3635 (N_3635,In_816,In_296);
nand U3636 (N_3636,In_38,In_762);
or U3637 (N_3637,In_924,In_120);
or U3638 (N_3638,In_160,In_153);
nand U3639 (N_3639,In_979,In_777);
nand U3640 (N_3640,In_168,In_531);
or U3641 (N_3641,In_799,In_212);
nor U3642 (N_3642,In_91,In_265);
nor U3643 (N_3643,In_976,In_47);
or U3644 (N_3644,In_790,In_829);
nand U3645 (N_3645,In_998,In_325);
or U3646 (N_3646,In_806,In_52);
and U3647 (N_3647,In_470,In_680);
and U3648 (N_3648,In_508,In_720);
or U3649 (N_3649,In_239,In_760);
or U3650 (N_3650,In_695,In_746);
and U3651 (N_3651,In_263,In_340);
or U3652 (N_3652,In_97,In_245);
and U3653 (N_3653,In_435,In_843);
or U3654 (N_3654,In_39,In_938);
and U3655 (N_3655,In_129,In_967);
nand U3656 (N_3656,In_906,In_559);
nor U3657 (N_3657,In_886,In_250);
nor U3658 (N_3658,In_840,In_168);
or U3659 (N_3659,In_289,In_419);
or U3660 (N_3660,In_46,In_316);
or U3661 (N_3661,In_12,In_866);
and U3662 (N_3662,In_878,In_368);
or U3663 (N_3663,In_4,In_726);
xnor U3664 (N_3664,In_4,In_629);
and U3665 (N_3665,In_384,In_505);
nor U3666 (N_3666,In_313,In_744);
and U3667 (N_3667,In_105,In_368);
and U3668 (N_3668,In_281,In_542);
and U3669 (N_3669,In_449,In_700);
or U3670 (N_3670,In_75,In_782);
or U3671 (N_3671,In_328,In_530);
nand U3672 (N_3672,In_609,In_713);
nor U3673 (N_3673,In_740,In_24);
nand U3674 (N_3674,In_304,In_869);
nand U3675 (N_3675,In_586,In_923);
nor U3676 (N_3676,In_311,In_265);
nor U3677 (N_3677,In_123,In_420);
nor U3678 (N_3678,In_581,In_479);
nand U3679 (N_3679,In_995,In_285);
nand U3680 (N_3680,In_577,In_664);
and U3681 (N_3681,In_679,In_450);
or U3682 (N_3682,In_909,In_918);
nand U3683 (N_3683,In_941,In_529);
and U3684 (N_3684,In_803,In_395);
and U3685 (N_3685,In_406,In_402);
nor U3686 (N_3686,In_649,In_444);
and U3687 (N_3687,In_596,In_449);
nand U3688 (N_3688,In_287,In_80);
and U3689 (N_3689,In_127,In_434);
nand U3690 (N_3690,In_191,In_49);
nand U3691 (N_3691,In_893,In_377);
nor U3692 (N_3692,In_177,In_585);
nand U3693 (N_3693,In_698,In_119);
and U3694 (N_3694,In_581,In_534);
nand U3695 (N_3695,In_770,In_531);
and U3696 (N_3696,In_693,In_758);
and U3697 (N_3697,In_546,In_207);
or U3698 (N_3698,In_945,In_711);
xnor U3699 (N_3699,In_481,In_514);
or U3700 (N_3700,In_512,In_954);
or U3701 (N_3701,In_346,In_908);
nor U3702 (N_3702,In_375,In_413);
nor U3703 (N_3703,In_879,In_768);
or U3704 (N_3704,In_878,In_801);
or U3705 (N_3705,In_598,In_532);
nand U3706 (N_3706,In_268,In_153);
nor U3707 (N_3707,In_238,In_866);
and U3708 (N_3708,In_605,In_541);
nand U3709 (N_3709,In_209,In_547);
nor U3710 (N_3710,In_520,In_262);
or U3711 (N_3711,In_858,In_98);
nor U3712 (N_3712,In_952,In_580);
nand U3713 (N_3713,In_553,In_199);
nor U3714 (N_3714,In_728,In_609);
nand U3715 (N_3715,In_62,In_835);
nor U3716 (N_3716,In_750,In_321);
nor U3717 (N_3717,In_650,In_250);
nand U3718 (N_3718,In_790,In_192);
or U3719 (N_3719,In_280,In_361);
nor U3720 (N_3720,In_569,In_671);
and U3721 (N_3721,In_595,In_533);
nand U3722 (N_3722,In_649,In_770);
nand U3723 (N_3723,In_417,In_361);
and U3724 (N_3724,In_127,In_810);
nor U3725 (N_3725,In_43,In_258);
and U3726 (N_3726,In_57,In_903);
or U3727 (N_3727,In_508,In_975);
nand U3728 (N_3728,In_331,In_126);
nor U3729 (N_3729,In_821,In_462);
nand U3730 (N_3730,In_468,In_698);
nor U3731 (N_3731,In_52,In_399);
and U3732 (N_3732,In_993,In_431);
nor U3733 (N_3733,In_156,In_12);
nand U3734 (N_3734,In_328,In_278);
or U3735 (N_3735,In_645,In_43);
or U3736 (N_3736,In_272,In_915);
nand U3737 (N_3737,In_492,In_537);
nand U3738 (N_3738,In_943,In_189);
and U3739 (N_3739,In_760,In_229);
or U3740 (N_3740,In_900,In_483);
or U3741 (N_3741,In_726,In_348);
or U3742 (N_3742,In_945,In_936);
or U3743 (N_3743,In_672,In_619);
nor U3744 (N_3744,In_386,In_954);
or U3745 (N_3745,In_966,In_92);
or U3746 (N_3746,In_104,In_205);
nor U3747 (N_3747,In_477,In_707);
nand U3748 (N_3748,In_596,In_378);
nand U3749 (N_3749,In_686,In_911);
or U3750 (N_3750,In_493,In_545);
and U3751 (N_3751,In_517,In_97);
nand U3752 (N_3752,In_870,In_470);
or U3753 (N_3753,In_315,In_708);
or U3754 (N_3754,In_791,In_837);
and U3755 (N_3755,In_268,In_643);
nand U3756 (N_3756,In_349,In_479);
nand U3757 (N_3757,In_166,In_915);
and U3758 (N_3758,In_7,In_353);
and U3759 (N_3759,In_845,In_542);
nor U3760 (N_3760,In_767,In_329);
nand U3761 (N_3761,In_665,In_408);
nor U3762 (N_3762,In_391,In_70);
and U3763 (N_3763,In_111,In_410);
and U3764 (N_3764,In_82,In_848);
and U3765 (N_3765,In_477,In_585);
xor U3766 (N_3766,In_82,In_344);
nor U3767 (N_3767,In_663,In_306);
or U3768 (N_3768,In_75,In_706);
nand U3769 (N_3769,In_104,In_773);
and U3770 (N_3770,In_725,In_666);
nor U3771 (N_3771,In_37,In_109);
and U3772 (N_3772,In_978,In_412);
nor U3773 (N_3773,In_746,In_108);
and U3774 (N_3774,In_411,In_150);
nor U3775 (N_3775,In_123,In_574);
nand U3776 (N_3776,In_186,In_325);
nor U3777 (N_3777,In_607,In_413);
nand U3778 (N_3778,In_518,In_727);
nand U3779 (N_3779,In_73,In_224);
and U3780 (N_3780,In_245,In_504);
or U3781 (N_3781,In_973,In_286);
nor U3782 (N_3782,In_251,In_542);
and U3783 (N_3783,In_758,In_429);
and U3784 (N_3784,In_233,In_153);
nand U3785 (N_3785,In_553,In_314);
nand U3786 (N_3786,In_532,In_382);
nor U3787 (N_3787,In_659,In_81);
nor U3788 (N_3788,In_51,In_953);
nor U3789 (N_3789,In_266,In_757);
or U3790 (N_3790,In_649,In_153);
nand U3791 (N_3791,In_467,In_304);
nand U3792 (N_3792,In_790,In_180);
nand U3793 (N_3793,In_208,In_515);
nor U3794 (N_3794,In_811,In_742);
and U3795 (N_3795,In_233,In_722);
or U3796 (N_3796,In_199,In_311);
or U3797 (N_3797,In_428,In_653);
nand U3798 (N_3798,In_764,In_193);
nor U3799 (N_3799,In_105,In_389);
nand U3800 (N_3800,In_249,In_879);
nand U3801 (N_3801,In_100,In_828);
nor U3802 (N_3802,In_833,In_99);
or U3803 (N_3803,In_309,In_995);
and U3804 (N_3804,In_481,In_477);
nand U3805 (N_3805,In_727,In_686);
nand U3806 (N_3806,In_282,In_279);
and U3807 (N_3807,In_204,In_34);
and U3808 (N_3808,In_964,In_755);
or U3809 (N_3809,In_226,In_627);
or U3810 (N_3810,In_943,In_328);
and U3811 (N_3811,In_481,In_540);
and U3812 (N_3812,In_112,In_423);
nand U3813 (N_3813,In_205,In_344);
or U3814 (N_3814,In_490,In_163);
nor U3815 (N_3815,In_170,In_657);
or U3816 (N_3816,In_134,In_637);
and U3817 (N_3817,In_748,In_425);
nand U3818 (N_3818,In_423,In_243);
and U3819 (N_3819,In_261,In_106);
nor U3820 (N_3820,In_749,In_569);
nand U3821 (N_3821,In_997,In_425);
nor U3822 (N_3822,In_451,In_854);
and U3823 (N_3823,In_48,In_107);
nor U3824 (N_3824,In_311,In_720);
and U3825 (N_3825,In_577,In_591);
or U3826 (N_3826,In_614,In_306);
or U3827 (N_3827,In_914,In_104);
xor U3828 (N_3828,In_348,In_351);
and U3829 (N_3829,In_306,In_340);
and U3830 (N_3830,In_444,In_233);
nor U3831 (N_3831,In_252,In_912);
and U3832 (N_3832,In_239,In_383);
nand U3833 (N_3833,In_433,In_719);
and U3834 (N_3834,In_371,In_973);
nand U3835 (N_3835,In_463,In_539);
nor U3836 (N_3836,In_975,In_427);
nor U3837 (N_3837,In_121,In_459);
nand U3838 (N_3838,In_538,In_529);
and U3839 (N_3839,In_106,In_912);
or U3840 (N_3840,In_569,In_286);
nand U3841 (N_3841,In_419,In_731);
xnor U3842 (N_3842,In_621,In_958);
nor U3843 (N_3843,In_252,In_264);
nand U3844 (N_3844,In_873,In_605);
and U3845 (N_3845,In_99,In_713);
or U3846 (N_3846,In_677,In_554);
nand U3847 (N_3847,In_568,In_499);
nor U3848 (N_3848,In_38,In_360);
nor U3849 (N_3849,In_913,In_742);
nor U3850 (N_3850,In_578,In_318);
xnor U3851 (N_3851,In_72,In_13);
nor U3852 (N_3852,In_348,In_471);
nor U3853 (N_3853,In_991,In_565);
or U3854 (N_3854,In_703,In_131);
nor U3855 (N_3855,In_796,In_408);
and U3856 (N_3856,In_114,In_821);
nand U3857 (N_3857,In_810,In_608);
nor U3858 (N_3858,In_351,In_529);
or U3859 (N_3859,In_976,In_614);
xnor U3860 (N_3860,In_276,In_635);
and U3861 (N_3861,In_596,In_135);
nand U3862 (N_3862,In_69,In_373);
nor U3863 (N_3863,In_309,In_638);
or U3864 (N_3864,In_628,In_954);
or U3865 (N_3865,In_173,In_70);
nand U3866 (N_3866,In_516,In_341);
nand U3867 (N_3867,In_260,In_850);
nor U3868 (N_3868,In_160,In_402);
and U3869 (N_3869,In_432,In_678);
or U3870 (N_3870,In_922,In_97);
and U3871 (N_3871,In_884,In_52);
nor U3872 (N_3872,In_706,In_928);
and U3873 (N_3873,In_137,In_352);
or U3874 (N_3874,In_67,In_871);
or U3875 (N_3875,In_345,In_198);
nand U3876 (N_3876,In_989,In_201);
nor U3877 (N_3877,In_390,In_885);
or U3878 (N_3878,In_295,In_849);
nand U3879 (N_3879,In_980,In_86);
or U3880 (N_3880,In_31,In_894);
nor U3881 (N_3881,In_798,In_312);
nor U3882 (N_3882,In_296,In_751);
nand U3883 (N_3883,In_933,In_664);
nor U3884 (N_3884,In_109,In_418);
or U3885 (N_3885,In_27,In_443);
nand U3886 (N_3886,In_829,In_355);
nor U3887 (N_3887,In_473,In_116);
nand U3888 (N_3888,In_259,In_112);
nand U3889 (N_3889,In_77,In_656);
nand U3890 (N_3890,In_865,In_868);
or U3891 (N_3891,In_131,In_857);
or U3892 (N_3892,In_418,In_986);
nand U3893 (N_3893,In_722,In_750);
or U3894 (N_3894,In_298,In_911);
or U3895 (N_3895,In_611,In_103);
or U3896 (N_3896,In_101,In_269);
and U3897 (N_3897,In_891,In_248);
nand U3898 (N_3898,In_109,In_932);
and U3899 (N_3899,In_582,In_525);
and U3900 (N_3900,In_388,In_193);
nand U3901 (N_3901,In_631,In_240);
and U3902 (N_3902,In_123,In_499);
nor U3903 (N_3903,In_397,In_628);
or U3904 (N_3904,In_199,In_78);
nand U3905 (N_3905,In_391,In_271);
and U3906 (N_3906,In_118,In_89);
or U3907 (N_3907,In_803,In_651);
nand U3908 (N_3908,In_538,In_355);
and U3909 (N_3909,In_652,In_635);
and U3910 (N_3910,In_684,In_397);
and U3911 (N_3911,In_855,In_659);
nand U3912 (N_3912,In_399,In_220);
and U3913 (N_3913,In_598,In_497);
and U3914 (N_3914,In_527,In_785);
nor U3915 (N_3915,In_94,In_875);
and U3916 (N_3916,In_734,In_991);
nand U3917 (N_3917,In_35,In_243);
or U3918 (N_3918,In_297,In_920);
nand U3919 (N_3919,In_219,In_691);
and U3920 (N_3920,In_927,In_353);
nand U3921 (N_3921,In_382,In_898);
nor U3922 (N_3922,In_755,In_819);
nor U3923 (N_3923,In_384,In_533);
and U3924 (N_3924,In_323,In_194);
or U3925 (N_3925,In_915,In_94);
nor U3926 (N_3926,In_49,In_859);
nand U3927 (N_3927,In_641,In_976);
and U3928 (N_3928,In_706,In_144);
or U3929 (N_3929,In_434,In_12);
and U3930 (N_3930,In_456,In_982);
nand U3931 (N_3931,In_210,In_695);
and U3932 (N_3932,In_320,In_285);
and U3933 (N_3933,In_656,In_649);
and U3934 (N_3934,In_84,In_983);
nor U3935 (N_3935,In_532,In_411);
or U3936 (N_3936,In_431,In_608);
or U3937 (N_3937,In_933,In_209);
nor U3938 (N_3938,In_360,In_29);
nor U3939 (N_3939,In_757,In_698);
nor U3940 (N_3940,In_668,In_813);
or U3941 (N_3941,In_374,In_412);
xor U3942 (N_3942,In_247,In_774);
and U3943 (N_3943,In_789,In_489);
nand U3944 (N_3944,In_544,In_724);
or U3945 (N_3945,In_267,In_295);
and U3946 (N_3946,In_509,In_861);
or U3947 (N_3947,In_935,In_887);
nor U3948 (N_3948,In_564,In_701);
nand U3949 (N_3949,In_215,In_386);
or U3950 (N_3950,In_433,In_714);
nand U3951 (N_3951,In_258,In_120);
nor U3952 (N_3952,In_408,In_564);
and U3953 (N_3953,In_609,In_928);
or U3954 (N_3954,In_307,In_521);
or U3955 (N_3955,In_84,In_460);
nor U3956 (N_3956,In_402,In_561);
nand U3957 (N_3957,In_763,In_332);
nor U3958 (N_3958,In_595,In_588);
nor U3959 (N_3959,In_695,In_535);
nor U3960 (N_3960,In_142,In_763);
and U3961 (N_3961,In_812,In_941);
nor U3962 (N_3962,In_19,In_608);
nand U3963 (N_3963,In_37,In_633);
or U3964 (N_3964,In_950,In_921);
and U3965 (N_3965,In_69,In_993);
nand U3966 (N_3966,In_586,In_269);
nand U3967 (N_3967,In_209,In_498);
or U3968 (N_3968,In_231,In_867);
nor U3969 (N_3969,In_979,In_758);
nor U3970 (N_3970,In_893,In_330);
nor U3971 (N_3971,In_584,In_302);
nand U3972 (N_3972,In_520,In_992);
or U3973 (N_3973,In_647,In_386);
and U3974 (N_3974,In_263,In_415);
and U3975 (N_3975,In_373,In_336);
or U3976 (N_3976,In_373,In_412);
nand U3977 (N_3977,In_775,In_745);
nand U3978 (N_3978,In_681,In_818);
and U3979 (N_3979,In_183,In_68);
nor U3980 (N_3980,In_696,In_582);
xor U3981 (N_3981,In_423,In_543);
and U3982 (N_3982,In_829,In_704);
nand U3983 (N_3983,In_30,In_487);
nand U3984 (N_3984,In_192,In_639);
or U3985 (N_3985,In_56,In_789);
nor U3986 (N_3986,In_179,In_608);
nor U3987 (N_3987,In_345,In_825);
and U3988 (N_3988,In_602,In_611);
or U3989 (N_3989,In_73,In_94);
xnor U3990 (N_3990,In_789,In_765);
and U3991 (N_3991,In_823,In_87);
nand U3992 (N_3992,In_707,In_312);
nor U3993 (N_3993,In_73,In_640);
and U3994 (N_3994,In_34,In_938);
nand U3995 (N_3995,In_267,In_870);
nor U3996 (N_3996,In_440,In_586);
or U3997 (N_3997,In_870,In_15);
or U3998 (N_3998,In_680,In_151);
nand U3999 (N_3999,In_775,In_632);
or U4000 (N_4000,In_401,In_113);
and U4001 (N_4001,In_478,In_648);
or U4002 (N_4002,In_745,In_653);
nor U4003 (N_4003,In_855,In_168);
or U4004 (N_4004,In_886,In_981);
nor U4005 (N_4005,In_887,In_748);
nand U4006 (N_4006,In_910,In_344);
nand U4007 (N_4007,In_419,In_501);
nor U4008 (N_4008,In_725,In_891);
nor U4009 (N_4009,In_538,In_517);
and U4010 (N_4010,In_417,In_308);
xnor U4011 (N_4011,In_923,In_519);
nand U4012 (N_4012,In_271,In_452);
and U4013 (N_4013,In_989,In_830);
nand U4014 (N_4014,In_556,In_954);
nand U4015 (N_4015,In_310,In_542);
nand U4016 (N_4016,In_69,In_856);
nand U4017 (N_4017,In_175,In_38);
or U4018 (N_4018,In_841,In_996);
and U4019 (N_4019,In_122,In_316);
xor U4020 (N_4020,In_357,In_459);
or U4021 (N_4021,In_443,In_417);
nand U4022 (N_4022,In_383,In_306);
nand U4023 (N_4023,In_925,In_212);
or U4024 (N_4024,In_948,In_338);
nand U4025 (N_4025,In_168,In_472);
or U4026 (N_4026,In_956,In_318);
and U4027 (N_4027,In_874,In_442);
and U4028 (N_4028,In_447,In_149);
or U4029 (N_4029,In_225,In_649);
nor U4030 (N_4030,In_506,In_717);
nand U4031 (N_4031,In_746,In_67);
nand U4032 (N_4032,In_591,In_667);
or U4033 (N_4033,In_470,In_794);
nor U4034 (N_4034,In_791,In_326);
or U4035 (N_4035,In_291,In_984);
nor U4036 (N_4036,In_325,In_495);
nor U4037 (N_4037,In_101,In_514);
and U4038 (N_4038,In_847,In_557);
or U4039 (N_4039,In_43,In_171);
nor U4040 (N_4040,In_77,In_235);
and U4041 (N_4041,In_439,In_363);
nand U4042 (N_4042,In_745,In_864);
or U4043 (N_4043,In_763,In_729);
nor U4044 (N_4044,In_286,In_600);
and U4045 (N_4045,In_365,In_207);
and U4046 (N_4046,In_353,In_337);
or U4047 (N_4047,In_270,In_212);
nand U4048 (N_4048,In_889,In_319);
and U4049 (N_4049,In_808,In_281);
and U4050 (N_4050,In_890,In_707);
nor U4051 (N_4051,In_522,In_357);
and U4052 (N_4052,In_660,In_146);
or U4053 (N_4053,In_826,In_865);
or U4054 (N_4054,In_525,In_250);
nor U4055 (N_4055,In_256,In_3);
or U4056 (N_4056,In_988,In_992);
or U4057 (N_4057,In_333,In_564);
or U4058 (N_4058,In_953,In_371);
and U4059 (N_4059,In_764,In_289);
nand U4060 (N_4060,In_131,In_513);
or U4061 (N_4061,In_704,In_9);
nor U4062 (N_4062,In_460,In_122);
and U4063 (N_4063,In_194,In_698);
nand U4064 (N_4064,In_44,In_34);
nor U4065 (N_4065,In_410,In_465);
and U4066 (N_4066,In_792,In_499);
xnor U4067 (N_4067,In_399,In_71);
or U4068 (N_4068,In_853,In_355);
nor U4069 (N_4069,In_124,In_639);
nand U4070 (N_4070,In_340,In_288);
or U4071 (N_4071,In_762,In_471);
nand U4072 (N_4072,In_3,In_139);
nand U4073 (N_4073,In_42,In_140);
nand U4074 (N_4074,In_563,In_591);
or U4075 (N_4075,In_559,In_973);
or U4076 (N_4076,In_894,In_247);
and U4077 (N_4077,In_333,In_187);
nor U4078 (N_4078,In_24,In_685);
or U4079 (N_4079,In_41,In_680);
or U4080 (N_4080,In_930,In_476);
or U4081 (N_4081,In_373,In_160);
nor U4082 (N_4082,In_298,In_293);
and U4083 (N_4083,In_117,In_75);
nand U4084 (N_4084,In_419,In_618);
and U4085 (N_4085,In_238,In_555);
and U4086 (N_4086,In_351,In_831);
or U4087 (N_4087,In_241,In_321);
or U4088 (N_4088,In_347,In_767);
nand U4089 (N_4089,In_236,In_99);
xor U4090 (N_4090,In_207,In_269);
nor U4091 (N_4091,In_197,In_955);
and U4092 (N_4092,In_897,In_23);
nand U4093 (N_4093,In_351,In_161);
nor U4094 (N_4094,In_616,In_962);
nand U4095 (N_4095,In_649,In_624);
and U4096 (N_4096,In_451,In_934);
nand U4097 (N_4097,In_83,In_588);
and U4098 (N_4098,In_113,In_941);
or U4099 (N_4099,In_794,In_926);
nor U4100 (N_4100,In_875,In_429);
and U4101 (N_4101,In_982,In_773);
and U4102 (N_4102,In_351,In_890);
or U4103 (N_4103,In_408,In_224);
or U4104 (N_4104,In_924,In_476);
nor U4105 (N_4105,In_10,In_763);
or U4106 (N_4106,In_979,In_907);
nand U4107 (N_4107,In_687,In_625);
nand U4108 (N_4108,In_99,In_101);
or U4109 (N_4109,In_501,In_679);
and U4110 (N_4110,In_587,In_527);
nand U4111 (N_4111,In_226,In_665);
or U4112 (N_4112,In_621,In_664);
or U4113 (N_4113,In_470,In_458);
and U4114 (N_4114,In_99,In_200);
and U4115 (N_4115,In_129,In_142);
or U4116 (N_4116,In_90,In_250);
nor U4117 (N_4117,In_840,In_475);
and U4118 (N_4118,In_547,In_748);
nand U4119 (N_4119,In_963,In_657);
or U4120 (N_4120,In_120,In_149);
and U4121 (N_4121,In_989,In_760);
and U4122 (N_4122,In_217,In_279);
nor U4123 (N_4123,In_292,In_662);
nor U4124 (N_4124,In_941,In_312);
nand U4125 (N_4125,In_588,In_811);
and U4126 (N_4126,In_357,In_621);
and U4127 (N_4127,In_302,In_238);
nand U4128 (N_4128,In_428,In_57);
nand U4129 (N_4129,In_745,In_755);
nor U4130 (N_4130,In_340,In_861);
and U4131 (N_4131,In_530,In_369);
nor U4132 (N_4132,In_894,In_502);
and U4133 (N_4133,In_737,In_735);
or U4134 (N_4134,In_754,In_262);
or U4135 (N_4135,In_892,In_845);
and U4136 (N_4136,In_903,In_849);
nor U4137 (N_4137,In_534,In_538);
or U4138 (N_4138,In_966,In_350);
or U4139 (N_4139,In_923,In_338);
nand U4140 (N_4140,In_568,In_603);
or U4141 (N_4141,In_654,In_749);
nor U4142 (N_4142,In_935,In_162);
or U4143 (N_4143,In_531,In_557);
and U4144 (N_4144,In_919,In_40);
nor U4145 (N_4145,In_581,In_49);
nand U4146 (N_4146,In_437,In_885);
xor U4147 (N_4147,In_195,In_137);
nor U4148 (N_4148,In_460,In_502);
nand U4149 (N_4149,In_727,In_883);
xnor U4150 (N_4150,In_724,In_661);
or U4151 (N_4151,In_660,In_9);
and U4152 (N_4152,In_518,In_514);
xor U4153 (N_4153,In_563,In_285);
nand U4154 (N_4154,In_667,In_125);
or U4155 (N_4155,In_845,In_376);
and U4156 (N_4156,In_331,In_391);
nor U4157 (N_4157,In_405,In_316);
nand U4158 (N_4158,In_279,In_956);
nand U4159 (N_4159,In_905,In_498);
and U4160 (N_4160,In_681,In_105);
nor U4161 (N_4161,In_361,In_906);
nor U4162 (N_4162,In_379,In_577);
or U4163 (N_4163,In_532,In_285);
nor U4164 (N_4164,In_600,In_732);
and U4165 (N_4165,In_683,In_25);
and U4166 (N_4166,In_71,In_888);
nand U4167 (N_4167,In_226,In_909);
or U4168 (N_4168,In_584,In_828);
nor U4169 (N_4169,In_968,In_887);
nor U4170 (N_4170,In_213,In_162);
nand U4171 (N_4171,In_303,In_431);
or U4172 (N_4172,In_209,In_640);
nor U4173 (N_4173,In_414,In_140);
and U4174 (N_4174,In_122,In_937);
and U4175 (N_4175,In_473,In_654);
or U4176 (N_4176,In_790,In_809);
or U4177 (N_4177,In_205,In_496);
or U4178 (N_4178,In_866,In_789);
nand U4179 (N_4179,In_144,In_630);
and U4180 (N_4180,In_930,In_460);
nor U4181 (N_4181,In_169,In_118);
nor U4182 (N_4182,In_803,In_991);
nor U4183 (N_4183,In_574,In_183);
and U4184 (N_4184,In_881,In_479);
nand U4185 (N_4185,In_153,In_174);
nand U4186 (N_4186,In_61,In_190);
and U4187 (N_4187,In_617,In_685);
and U4188 (N_4188,In_826,In_93);
or U4189 (N_4189,In_893,In_721);
and U4190 (N_4190,In_156,In_235);
or U4191 (N_4191,In_672,In_408);
nor U4192 (N_4192,In_25,In_956);
nand U4193 (N_4193,In_291,In_681);
nor U4194 (N_4194,In_524,In_769);
or U4195 (N_4195,In_323,In_519);
nor U4196 (N_4196,In_424,In_54);
nand U4197 (N_4197,In_536,In_870);
nor U4198 (N_4198,In_619,In_231);
and U4199 (N_4199,In_975,In_624);
nand U4200 (N_4200,In_328,In_793);
nand U4201 (N_4201,In_555,In_447);
nor U4202 (N_4202,In_824,In_964);
and U4203 (N_4203,In_363,In_278);
nand U4204 (N_4204,In_374,In_23);
and U4205 (N_4205,In_311,In_271);
nand U4206 (N_4206,In_632,In_633);
nand U4207 (N_4207,In_564,In_795);
or U4208 (N_4208,In_521,In_920);
nand U4209 (N_4209,In_185,In_552);
nor U4210 (N_4210,In_395,In_176);
and U4211 (N_4211,In_11,In_703);
or U4212 (N_4212,In_898,In_374);
or U4213 (N_4213,In_638,In_52);
nand U4214 (N_4214,In_806,In_962);
or U4215 (N_4215,In_402,In_218);
and U4216 (N_4216,In_580,In_781);
nor U4217 (N_4217,In_593,In_876);
nor U4218 (N_4218,In_535,In_403);
nand U4219 (N_4219,In_616,In_497);
and U4220 (N_4220,In_727,In_440);
and U4221 (N_4221,In_405,In_960);
and U4222 (N_4222,In_769,In_606);
or U4223 (N_4223,In_241,In_895);
xnor U4224 (N_4224,In_175,In_46);
nor U4225 (N_4225,In_408,In_678);
or U4226 (N_4226,In_949,In_727);
and U4227 (N_4227,In_397,In_836);
nand U4228 (N_4228,In_587,In_4);
nand U4229 (N_4229,In_220,In_721);
and U4230 (N_4230,In_402,In_120);
nand U4231 (N_4231,In_291,In_621);
nor U4232 (N_4232,In_902,In_206);
nand U4233 (N_4233,In_372,In_82);
nand U4234 (N_4234,In_783,In_129);
or U4235 (N_4235,In_511,In_215);
nor U4236 (N_4236,In_671,In_483);
and U4237 (N_4237,In_223,In_154);
or U4238 (N_4238,In_604,In_34);
nor U4239 (N_4239,In_231,In_253);
nand U4240 (N_4240,In_999,In_883);
nand U4241 (N_4241,In_713,In_213);
nor U4242 (N_4242,In_12,In_889);
or U4243 (N_4243,In_381,In_417);
or U4244 (N_4244,In_603,In_39);
or U4245 (N_4245,In_490,In_963);
nand U4246 (N_4246,In_588,In_203);
and U4247 (N_4247,In_491,In_434);
nand U4248 (N_4248,In_148,In_753);
and U4249 (N_4249,In_482,In_368);
or U4250 (N_4250,In_872,In_403);
or U4251 (N_4251,In_485,In_519);
nor U4252 (N_4252,In_347,In_778);
nor U4253 (N_4253,In_368,In_624);
and U4254 (N_4254,In_706,In_299);
nor U4255 (N_4255,In_593,In_903);
nand U4256 (N_4256,In_89,In_154);
or U4257 (N_4257,In_415,In_899);
nand U4258 (N_4258,In_28,In_928);
or U4259 (N_4259,In_851,In_846);
and U4260 (N_4260,In_227,In_635);
nor U4261 (N_4261,In_803,In_509);
or U4262 (N_4262,In_742,In_438);
nand U4263 (N_4263,In_579,In_448);
nand U4264 (N_4264,In_429,In_590);
and U4265 (N_4265,In_109,In_419);
nor U4266 (N_4266,In_370,In_609);
or U4267 (N_4267,In_55,In_964);
or U4268 (N_4268,In_334,In_545);
nand U4269 (N_4269,In_42,In_877);
nor U4270 (N_4270,In_386,In_51);
and U4271 (N_4271,In_771,In_914);
and U4272 (N_4272,In_252,In_37);
nand U4273 (N_4273,In_262,In_922);
nor U4274 (N_4274,In_810,In_203);
or U4275 (N_4275,In_243,In_179);
and U4276 (N_4276,In_270,In_677);
nand U4277 (N_4277,In_580,In_147);
or U4278 (N_4278,In_361,In_291);
and U4279 (N_4279,In_645,In_400);
or U4280 (N_4280,In_755,In_215);
or U4281 (N_4281,In_347,In_602);
or U4282 (N_4282,In_568,In_924);
nor U4283 (N_4283,In_765,In_742);
nor U4284 (N_4284,In_930,In_139);
nor U4285 (N_4285,In_616,In_51);
and U4286 (N_4286,In_180,In_213);
nor U4287 (N_4287,In_411,In_890);
nand U4288 (N_4288,In_134,In_973);
nand U4289 (N_4289,In_585,In_816);
nand U4290 (N_4290,In_649,In_840);
nand U4291 (N_4291,In_931,In_145);
nor U4292 (N_4292,In_558,In_855);
nand U4293 (N_4293,In_250,In_486);
and U4294 (N_4294,In_220,In_864);
nor U4295 (N_4295,In_130,In_380);
and U4296 (N_4296,In_688,In_769);
xnor U4297 (N_4297,In_289,In_568);
nand U4298 (N_4298,In_299,In_870);
or U4299 (N_4299,In_455,In_569);
nor U4300 (N_4300,In_80,In_263);
and U4301 (N_4301,In_55,In_966);
or U4302 (N_4302,In_813,In_144);
and U4303 (N_4303,In_189,In_569);
and U4304 (N_4304,In_467,In_432);
nor U4305 (N_4305,In_783,In_499);
or U4306 (N_4306,In_651,In_656);
and U4307 (N_4307,In_955,In_324);
and U4308 (N_4308,In_37,In_465);
nand U4309 (N_4309,In_689,In_665);
or U4310 (N_4310,In_358,In_705);
nand U4311 (N_4311,In_316,In_342);
or U4312 (N_4312,In_916,In_787);
nand U4313 (N_4313,In_426,In_930);
nor U4314 (N_4314,In_193,In_798);
and U4315 (N_4315,In_97,In_697);
nor U4316 (N_4316,In_347,In_422);
xor U4317 (N_4317,In_248,In_453);
nand U4318 (N_4318,In_264,In_438);
nor U4319 (N_4319,In_811,In_604);
and U4320 (N_4320,In_829,In_527);
nor U4321 (N_4321,In_567,In_710);
and U4322 (N_4322,In_769,In_849);
nor U4323 (N_4323,In_900,In_750);
nor U4324 (N_4324,In_541,In_178);
nand U4325 (N_4325,In_286,In_238);
nand U4326 (N_4326,In_213,In_151);
or U4327 (N_4327,In_439,In_15);
and U4328 (N_4328,In_140,In_49);
or U4329 (N_4329,In_127,In_171);
or U4330 (N_4330,In_569,In_926);
and U4331 (N_4331,In_549,In_554);
and U4332 (N_4332,In_678,In_8);
and U4333 (N_4333,In_964,In_772);
and U4334 (N_4334,In_981,In_339);
nand U4335 (N_4335,In_634,In_546);
or U4336 (N_4336,In_925,In_359);
nand U4337 (N_4337,In_767,In_337);
nor U4338 (N_4338,In_731,In_886);
nand U4339 (N_4339,In_728,In_139);
nor U4340 (N_4340,In_100,In_537);
nor U4341 (N_4341,In_800,In_924);
nor U4342 (N_4342,In_795,In_551);
nor U4343 (N_4343,In_976,In_379);
nor U4344 (N_4344,In_620,In_759);
and U4345 (N_4345,In_984,In_230);
nand U4346 (N_4346,In_683,In_736);
nand U4347 (N_4347,In_145,In_782);
or U4348 (N_4348,In_61,In_683);
and U4349 (N_4349,In_87,In_24);
nor U4350 (N_4350,In_209,In_805);
and U4351 (N_4351,In_317,In_998);
nand U4352 (N_4352,In_651,In_198);
or U4353 (N_4353,In_991,In_72);
nor U4354 (N_4354,In_683,In_439);
nand U4355 (N_4355,In_266,In_979);
or U4356 (N_4356,In_397,In_168);
or U4357 (N_4357,In_632,In_669);
or U4358 (N_4358,In_97,In_851);
and U4359 (N_4359,In_517,In_474);
nand U4360 (N_4360,In_558,In_841);
and U4361 (N_4361,In_83,In_290);
nor U4362 (N_4362,In_950,In_350);
nand U4363 (N_4363,In_531,In_569);
and U4364 (N_4364,In_606,In_824);
and U4365 (N_4365,In_371,In_372);
and U4366 (N_4366,In_922,In_49);
nand U4367 (N_4367,In_755,In_925);
nand U4368 (N_4368,In_498,In_234);
nand U4369 (N_4369,In_16,In_940);
or U4370 (N_4370,In_437,In_583);
nor U4371 (N_4371,In_731,In_597);
nand U4372 (N_4372,In_702,In_98);
nor U4373 (N_4373,In_780,In_992);
and U4374 (N_4374,In_694,In_220);
nor U4375 (N_4375,In_709,In_789);
nand U4376 (N_4376,In_285,In_738);
or U4377 (N_4377,In_914,In_517);
nand U4378 (N_4378,In_21,In_976);
and U4379 (N_4379,In_840,In_43);
nand U4380 (N_4380,In_762,In_469);
and U4381 (N_4381,In_252,In_678);
and U4382 (N_4382,In_277,In_268);
nand U4383 (N_4383,In_375,In_155);
and U4384 (N_4384,In_867,In_839);
nand U4385 (N_4385,In_174,In_250);
or U4386 (N_4386,In_622,In_398);
nand U4387 (N_4387,In_934,In_902);
or U4388 (N_4388,In_442,In_39);
or U4389 (N_4389,In_785,In_572);
nand U4390 (N_4390,In_765,In_416);
and U4391 (N_4391,In_72,In_805);
nor U4392 (N_4392,In_56,In_572);
and U4393 (N_4393,In_368,In_222);
or U4394 (N_4394,In_583,In_666);
nand U4395 (N_4395,In_18,In_645);
or U4396 (N_4396,In_791,In_866);
nor U4397 (N_4397,In_276,In_688);
or U4398 (N_4398,In_514,In_761);
nor U4399 (N_4399,In_598,In_746);
or U4400 (N_4400,In_921,In_133);
nand U4401 (N_4401,In_745,In_790);
or U4402 (N_4402,In_373,In_143);
nor U4403 (N_4403,In_3,In_356);
nand U4404 (N_4404,In_602,In_457);
nand U4405 (N_4405,In_648,In_927);
nand U4406 (N_4406,In_114,In_265);
or U4407 (N_4407,In_828,In_39);
and U4408 (N_4408,In_726,In_943);
xor U4409 (N_4409,In_781,In_164);
nand U4410 (N_4410,In_33,In_895);
and U4411 (N_4411,In_605,In_254);
or U4412 (N_4412,In_327,In_686);
nand U4413 (N_4413,In_730,In_232);
or U4414 (N_4414,In_59,In_737);
nor U4415 (N_4415,In_91,In_154);
nand U4416 (N_4416,In_65,In_237);
nand U4417 (N_4417,In_273,In_969);
or U4418 (N_4418,In_204,In_460);
nand U4419 (N_4419,In_420,In_963);
nor U4420 (N_4420,In_643,In_952);
nand U4421 (N_4421,In_823,In_811);
nor U4422 (N_4422,In_368,In_823);
nand U4423 (N_4423,In_95,In_720);
nand U4424 (N_4424,In_75,In_64);
nor U4425 (N_4425,In_411,In_245);
and U4426 (N_4426,In_177,In_207);
xor U4427 (N_4427,In_427,In_1);
or U4428 (N_4428,In_505,In_47);
and U4429 (N_4429,In_134,In_635);
nand U4430 (N_4430,In_652,In_793);
nor U4431 (N_4431,In_913,In_332);
and U4432 (N_4432,In_792,In_179);
or U4433 (N_4433,In_309,In_938);
nand U4434 (N_4434,In_402,In_473);
or U4435 (N_4435,In_36,In_211);
or U4436 (N_4436,In_352,In_378);
or U4437 (N_4437,In_616,In_600);
and U4438 (N_4438,In_861,In_748);
nor U4439 (N_4439,In_551,In_361);
nand U4440 (N_4440,In_697,In_423);
nor U4441 (N_4441,In_823,In_661);
and U4442 (N_4442,In_976,In_965);
and U4443 (N_4443,In_963,In_128);
nor U4444 (N_4444,In_580,In_918);
and U4445 (N_4445,In_700,In_118);
and U4446 (N_4446,In_382,In_524);
nand U4447 (N_4447,In_367,In_403);
or U4448 (N_4448,In_628,In_122);
nand U4449 (N_4449,In_418,In_474);
or U4450 (N_4450,In_303,In_219);
nor U4451 (N_4451,In_342,In_122);
nand U4452 (N_4452,In_483,In_818);
nand U4453 (N_4453,In_348,In_314);
or U4454 (N_4454,In_114,In_601);
nand U4455 (N_4455,In_591,In_428);
or U4456 (N_4456,In_406,In_269);
and U4457 (N_4457,In_181,In_8);
nor U4458 (N_4458,In_639,In_96);
nor U4459 (N_4459,In_286,In_576);
nand U4460 (N_4460,In_505,In_596);
or U4461 (N_4461,In_860,In_731);
nor U4462 (N_4462,In_39,In_977);
nor U4463 (N_4463,In_739,In_628);
nand U4464 (N_4464,In_103,In_395);
and U4465 (N_4465,In_82,In_580);
nand U4466 (N_4466,In_180,In_994);
or U4467 (N_4467,In_384,In_71);
nor U4468 (N_4468,In_447,In_987);
and U4469 (N_4469,In_404,In_417);
and U4470 (N_4470,In_22,In_695);
nor U4471 (N_4471,In_553,In_735);
or U4472 (N_4472,In_839,In_485);
and U4473 (N_4473,In_134,In_843);
and U4474 (N_4474,In_801,In_53);
nand U4475 (N_4475,In_636,In_176);
and U4476 (N_4476,In_518,In_777);
or U4477 (N_4477,In_474,In_920);
nor U4478 (N_4478,In_997,In_765);
or U4479 (N_4479,In_533,In_958);
or U4480 (N_4480,In_278,In_316);
or U4481 (N_4481,In_5,In_388);
or U4482 (N_4482,In_758,In_920);
nor U4483 (N_4483,In_625,In_227);
and U4484 (N_4484,In_872,In_460);
nand U4485 (N_4485,In_950,In_609);
nand U4486 (N_4486,In_511,In_562);
nor U4487 (N_4487,In_61,In_804);
nor U4488 (N_4488,In_497,In_675);
and U4489 (N_4489,In_865,In_852);
nor U4490 (N_4490,In_976,In_28);
and U4491 (N_4491,In_258,In_103);
nor U4492 (N_4492,In_514,In_742);
or U4493 (N_4493,In_424,In_743);
and U4494 (N_4494,In_912,In_775);
nor U4495 (N_4495,In_750,In_873);
nand U4496 (N_4496,In_782,In_146);
nand U4497 (N_4497,In_496,In_208);
nor U4498 (N_4498,In_542,In_492);
and U4499 (N_4499,In_366,In_565);
nor U4500 (N_4500,In_720,In_560);
and U4501 (N_4501,In_376,In_185);
and U4502 (N_4502,In_451,In_24);
or U4503 (N_4503,In_992,In_920);
and U4504 (N_4504,In_612,In_16);
and U4505 (N_4505,In_14,In_997);
nor U4506 (N_4506,In_728,In_885);
nand U4507 (N_4507,In_96,In_825);
and U4508 (N_4508,In_969,In_590);
or U4509 (N_4509,In_910,In_743);
nor U4510 (N_4510,In_275,In_240);
or U4511 (N_4511,In_88,In_332);
nand U4512 (N_4512,In_828,In_699);
and U4513 (N_4513,In_707,In_878);
or U4514 (N_4514,In_188,In_950);
nand U4515 (N_4515,In_294,In_650);
or U4516 (N_4516,In_391,In_170);
nand U4517 (N_4517,In_613,In_266);
nor U4518 (N_4518,In_635,In_495);
nand U4519 (N_4519,In_270,In_30);
nor U4520 (N_4520,In_105,In_724);
nor U4521 (N_4521,In_674,In_81);
nand U4522 (N_4522,In_307,In_564);
or U4523 (N_4523,In_633,In_358);
and U4524 (N_4524,In_590,In_538);
nor U4525 (N_4525,In_543,In_427);
nor U4526 (N_4526,In_56,In_779);
nor U4527 (N_4527,In_899,In_122);
and U4528 (N_4528,In_798,In_318);
nor U4529 (N_4529,In_541,In_24);
and U4530 (N_4530,In_456,In_863);
nor U4531 (N_4531,In_3,In_408);
nor U4532 (N_4532,In_478,In_899);
and U4533 (N_4533,In_739,In_253);
nor U4534 (N_4534,In_96,In_966);
nor U4535 (N_4535,In_282,In_50);
or U4536 (N_4536,In_380,In_329);
nor U4537 (N_4537,In_198,In_427);
nor U4538 (N_4538,In_422,In_850);
nor U4539 (N_4539,In_650,In_743);
or U4540 (N_4540,In_245,In_982);
nand U4541 (N_4541,In_943,In_512);
or U4542 (N_4542,In_366,In_835);
nor U4543 (N_4543,In_578,In_906);
nand U4544 (N_4544,In_959,In_697);
or U4545 (N_4545,In_388,In_30);
or U4546 (N_4546,In_273,In_542);
and U4547 (N_4547,In_369,In_601);
nand U4548 (N_4548,In_650,In_733);
or U4549 (N_4549,In_734,In_891);
nand U4550 (N_4550,In_302,In_337);
nand U4551 (N_4551,In_325,In_73);
nand U4552 (N_4552,In_234,In_175);
nor U4553 (N_4553,In_707,In_320);
nand U4554 (N_4554,In_50,In_106);
or U4555 (N_4555,In_596,In_970);
or U4556 (N_4556,In_269,In_592);
and U4557 (N_4557,In_811,In_475);
nor U4558 (N_4558,In_140,In_152);
or U4559 (N_4559,In_875,In_604);
or U4560 (N_4560,In_516,In_10);
nand U4561 (N_4561,In_616,In_396);
and U4562 (N_4562,In_114,In_528);
nor U4563 (N_4563,In_120,In_718);
nor U4564 (N_4564,In_158,In_576);
nand U4565 (N_4565,In_229,In_886);
nor U4566 (N_4566,In_5,In_736);
nor U4567 (N_4567,In_581,In_579);
nand U4568 (N_4568,In_520,In_340);
or U4569 (N_4569,In_796,In_973);
and U4570 (N_4570,In_525,In_183);
or U4571 (N_4571,In_602,In_814);
nand U4572 (N_4572,In_739,In_434);
nand U4573 (N_4573,In_647,In_805);
nor U4574 (N_4574,In_778,In_964);
nor U4575 (N_4575,In_324,In_984);
nor U4576 (N_4576,In_475,In_703);
and U4577 (N_4577,In_141,In_653);
nor U4578 (N_4578,In_225,In_934);
nand U4579 (N_4579,In_341,In_330);
and U4580 (N_4580,In_920,In_624);
and U4581 (N_4581,In_912,In_967);
nor U4582 (N_4582,In_989,In_615);
and U4583 (N_4583,In_928,In_606);
and U4584 (N_4584,In_330,In_584);
and U4585 (N_4585,In_974,In_249);
or U4586 (N_4586,In_546,In_13);
and U4587 (N_4587,In_407,In_502);
nand U4588 (N_4588,In_380,In_637);
and U4589 (N_4589,In_353,In_327);
nor U4590 (N_4590,In_373,In_21);
and U4591 (N_4591,In_452,In_111);
nor U4592 (N_4592,In_183,In_756);
nor U4593 (N_4593,In_911,In_803);
nand U4594 (N_4594,In_645,In_574);
or U4595 (N_4595,In_921,In_354);
nand U4596 (N_4596,In_872,In_290);
and U4597 (N_4597,In_510,In_752);
nand U4598 (N_4598,In_346,In_497);
or U4599 (N_4599,In_856,In_825);
and U4600 (N_4600,In_654,In_993);
and U4601 (N_4601,In_710,In_972);
or U4602 (N_4602,In_761,In_248);
nand U4603 (N_4603,In_775,In_860);
nand U4604 (N_4604,In_233,In_872);
and U4605 (N_4605,In_559,In_994);
or U4606 (N_4606,In_504,In_536);
or U4607 (N_4607,In_871,In_406);
nand U4608 (N_4608,In_814,In_835);
or U4609 (N_4609,In_926,In_78);
and U4610 (N_4610,In_6,In_768);
nor U4611 (N_4611,In_968,In_560);
nor U4612 (N_4612,In_292,In_526);
or U4613 (N_4613,In_978,In_89);
or U4614 (N_4614,In_259,In_730);
nand U4615 (N_4615,In_967,In_874);
or U4616 (N_4616,In_664,In_803);
nand U4617 (N_4617,In_819,In_704);
nor U4618 (N_4618,In_56,In_299);
nor U4619 (N_4619,In_83,In_214);
nand U4620 (N_4620,In_154,In_377);
or U4621 (N_4621,In_670,In_927);
nand U4622 (N_4622,In_56,In_781);
nand U4623 (N_4623,In_415,In_907);
or U4624 (N_4624,In_40,In_778);
nand U4625 (N_4625,In_354,In_41);
and U4626 (N_4626,In_898,In_77);
or U4627 (N_4627,In_0,In_760);
and U4628 (N_4628,In_527,In_781);
nand U4629 (N_4629,In_805,In_492);
nor U4630 (N_4630,In_731,In_644);
and U4631 (N_4631,In_958,In_305);
nor U4632 (N_4632,In_721,In_256);
or U4633 (N_4633,In_884,In_421);
nand U4634 (N_4634,In_266,In_230);
nand U4635 (N_4635,In_53,In_44);
or U4636 (N_4636,In_293,In_530);
and U4637 (N_4637,In_569,In_420);
nand U4638 (N_4638,In_601,In_408);
nand U4639 (N_4639,In_694,In_986);
nand U4640 (N_4640,In_892,In_190);
nand U4641 (N_4641,In_19,In_86);
or U4642 (N_4642,In_228,In_911);
or U4643 (N_4643,In_823,In_786);
nand U4644 (N_4644,In_623,In_144);
nand U4645 (N_4645,In_339,In_819);
or U4646 (N_4646,In_367,In_965);
nor U4647 (N_4647,In_650,In_131);
or U4648 (N_4648,In_911,In_414);
and U4649 (N_4649,In_354,In_114);
and U4650 (N_4650,In_825,In_416);
and U4651 (N_4651,In_32,In_364);
nand U4652 (N_4652,In_958,In_860);
nand U4653 (N_4653,In_595,In_181);
or U4654 (N_4654,In_863,In_891);
and U4655 (N_4655,In_440,In_576);
nor U4656 (N_4656,In_828,In_244);
and U4657 (N_4657,In_108,In_300);
and U4658 (N_4658,In_838,In_290);
nand U4659 (N_4659,In_717,In_45);
and U4660 (N_4660,In_340,In_533);
nand U4661 (N_4661,In_13,In_471);
nand U4662 (N_4662,In_200,In_323);
or U4663 (N_4663,In_590,In_387);
or U4664 (N_4664,In_982,In_830);
nor U4665 (N_4665,In_638,In_868);
and U4666 (N_4666,In_954,In_673);
or U4667 (N_4667,In_875,In_83);
or U4668 (N_4668,In_241,In_301);
nand U4669 (N_4669,In_146,In_295);
nand U4670 (N_4670,In_339,In_351);
nor U4671 (N_4671,In_751,In_340);
nand U4672 (N_4672,In_502,In_879);
nand U4673 (N_4673,In_855,In_396);
nand U4674 (N_4674,In_116,In_907);
xor U4675 (N_4675,In_729,In_322);
nor U4676 (N_4676,In_899,In_292);
or U4677 (N_4677,In_135,In_139);
or U4678 (N_4678,In_918,In_845);
and U4679 (N_4679,In_693,In_160);
nand U4680 (N_4680,In_565,In_75);
and U4681 (N_4681,In_857,In_363);
nand U4682 (N_4682,In_378,In_618);
or U4683 (N_4683,In_760,In_65);
nand U4684 (N_4684,In_429,In_46);
and U4685 (N_4685,In_330,In_561);
or U4686 (N_4686,In_569,In_359);
and U4687 (N_4687,In_683,In_907);
nand U4688 (N_4688,In_608,In_391);
nand U4689 (N_4689,In_622,In_98);
nor U4690 (N_4690,In_717,In_523);
and U4691 (N_4691,In_638,In_432);
or U4692 (N_4692,In_205,In_0);
nand U4693 (N_4693,In_970,In_535);
and U4694 (N_4694,In_283,In_395);
nand U4695 (N_4695,In_23,In_525);
or U4696 (N_4696,In_201,In_200);
and U4697 (N_4697,In_922,In_574);
nor U4698 (N_4698,In_194,In_765);
and U4699 (N_4699,In_511,In_233);
and U4700 (N_4700,In_775,In_142);
nor U4701 (N_4701,In_350,In_236);
nor U4702 (N_4702,In_576,In_835);
nor U4703 (N_4703,In_280,In_633);
nand U4704 (N_4704,In_542,In_371);
nand U4705 (N_4705,In_958,In_947);
and U4706 (N_4706,In_704,In_910);
nor U4707 (N_4707,In_314,In_618);
or U4708 (N_4708,In_64,In_435);
and U4709 (N_4709,In_182,In_515);
or U4710 (N_4710,In_393,In_923);
nand U4711 (N_4711,In_633,In_341);
or U4712 (N_4712,In_574,In_136);
and U4713 (N_4713,In_51,In_237);
xnor U4714 (N_4714,In_68,In_544);
nor U4715 (N_4715,In_463,In_159);
nand U4716 (N_4716,In_598,In_212);
nor U4717 (N_4717,In_728,In_709);
or U4718 (N_4718,In_427,In_126);
nand U4719 (N_4719,In_811,In_966);
nor U4720 (N_4720,In_144,In_462);
or U4721 (N_4721,In_388,In_937);
and U4722 (N_4722,In_113,In_798);
nor U4723 (N_4723,In_10,In_17);
nor U4724 (N_4724,In_448,In_835);
and U4725 (N_4725,In_979,In_239);
xor U4726 (N_4726,In_63,In_237);
and U4727 (N_4727,In_558,In_397);
xnor U4728 (N_4728,In_413,In_384);
or U4729 (N_4729,In_219,In_533);
and U4730 (N_4730,In_911,In_856);
or U4731 (N_4731,In_114,In_535);
nor U4732 (N_4732,In_932,In_989);
and U4733 (N_4733,In_686,In_81);
or U4734 (N_4734,In_310,In_932);
or U4735 (N_4735,In_116,In_608);
and U4736 (N_4736,In_410,In_286);
or U4737 (N_4737,In_884,In_51);
or U4738 (N_4738,In_826,In_144);
and U4739 (N_4739,In_731,In_285);
or U4740 (N_4740,In_839,In_644);
nor U4741 (N_4741,In_263,In_326);
nor U4742 (N_4742,In_174,In_474);
nand U4743 (N_4743,In_322,In_558);
nor U4744 (N_4744,In_97,In_134);
nor U4745 (N_4745,In_980,In_34);
nand U4746 (N_4746,In_981,In_208);
nor U4747 (N_4747,In_121,In_445);
or U4748 (N_4748,In_417,In_49);
nand U4749 (N_4749,In_851,In_859);
and U4750 (N_4750,In_91,In_203);
or U4751 (N_4751,In_113,In_23);
or U4752 (N_4752,In_743,In_344);
nor U4753 (N_4753,In_627,In_388);
and U4754 (N_4754,In_427,In_137);
and U4755 (N_4755,In_886,In_22);
and U4756 (N_4756,In_175,In_415);
and U4757 (N_4757,In_997,In_217);
and U4758 (N_4758,In_480,In_866);
and U4759 (N_4759,In_991,In_407);
or U4760 (N_4760,In_926,In_813);
or U4761 (N_4761,In_549,In_34);
nand U4762 (N_4762,In_631,In_174);
nand U4763 (N_4763,In_518,In_743);
nor U4764 (N_4764,In_749,In_65);
nand U4765 (N_4765,In_561,In_255);
nor U4766 (N_4766,In_699,In_259);
nor U4767 (N_4767,In_483,In_795);
nor U4768 (N_4768,In_24,In_515);
nand U4769 (N_4769,In_722,In_871);
nor U4770 (N_4770,In_603,In_51);
nand U4771 (N_4771,In_117,In_42);
nor U4772 (N_4772,In_610,In_294);
nand U4773 (N_4773,In_105,In_757);
or U4774 (N_4774,In_395,In_370);
nor U4775 (N_4775,In_898,In_506);
or U4776 (N_4776,In_442,In_556);
and U4777 (N_4777,In_7,In_24);
nand U4778 (N_4778,In_895,In_711);
and U4779 (N_4779,In_178,In_585);
and U4780 (N_4780,In_410,In_548);
and U4781 (N_4781,In_810,In_673);
nor U4782 (N_4782,In_599,In_199);
nor U4783 (N_4783,In_477,In_982);
or U4784 (N_4784,In_202,In_258);
and U4785 (N_4785,In_124,In_259);
and U4786 (N_4786,In_888,In_987);
nand U4787 (N_4787,In_771,In_423);
and U4788 (N_4788,In_36,In_58);
or U4789 (N_4789,In_745,In_424);
nand U4790 (N_4790,In_966,In_237);
xor U4791 (N_4791,In_741,In_796);
or U4792 (N_4792,In_259,In_875);
and U4793 (N_4793,In_406,In_584);
or U4794 (N_4794,In_885,In_707);
or U4795 (N_4795,In_10,In_54);
and U4796 (N_4796,In_235,In_488);
nor U4797 (N_4797,In_559,In_124);
nand U4798 (N_4798,In_369,In_132);
nand U4799 (N_4799,In_795,In_322);
or U4800 (N_4800,In_373,In_774);
nand U4801 (N_4801,In_4,In_130);
and U4802 (N_4802,In_317,In_973);
and U4803 (N_4803,In_263,In_407);
nor U4804 (N_4804,In_106,In_455);
nor U4805 (N_4805,In_40,In_310);
and U4806 (N_4806,In_163,In_443);
and U4807 (N_4807,In_554,In_355);
nand U4808 (N_4808,In_285,In_175);
and U4809 (N_4809,In_422,In_531);
nor U4810 (N_4810,In_590,In_622);
nand U4811 (N_4811,In_130,In_19);
or U4812 (N_4812,In_812,In_214);
and U4813 (N_4813,In_42,In_458);
nand U4814 (N_4814,In_227,In_738);
nand U4815 (N_4815,In_88,In_893);
and U4816 (N_4816,In_512,In_869);
and U4817 (N_4817,In_857,In_432);
nor U4818 (N_4818,In_591,In_804);
and U4819 (N_4819,In_989,In_327);
and U4820 (N_4820,In_112,In_272);
nor U4821 (N_4821,In_768,In_697);
and U4822 (N_4822,In_801,In_626);
or U4823 (N_4823,In_389,In_186);
nor U4824 (N_4824,In_809,In_556);
and U4825 (N_4825,In_573,In_372);
and U4826 (N_4826,In_183,In_462);
and U4827 (N_4827,In_187,In_85);
or U4828 (N_4828,In_672,In_760);
nand U4829 (N_4829,In_75,In_678);
or U4830 (N_4830,In_891,In_315);
or U4831 (N_4831,In_36,In_610);
nor U4832 (N_4832,In_49,In_328);
nor U4833 (N_4833,In_390,In_956);
or U4834 (N_4834,In_182,In_857);
nor U4835 (N_4835,In_581,In_730);
nand U4836 (N_4836,In_878,In_968);
nor U4837 (N_4837,In_461,In_516);
and U4838 (N_4838,In_69,In_399);
and U4839 (N_4839,In_194,In_738);
nand U4840 (N_4840,In_418,In_328);
nand U4841 (N_4841,In_152,In_42);
nand U4842 (N_4842,In_53,In_36);
and U4843 (N_4843,In_750,In_575);
nand U4844 (N_4844,In_831,In_747);
nor U4845 (N_4845,In_670,In_998);
nand U4846 (N_4846,In_852,In_112);
nor U4847 (N_4847,In_791,In_24);
nand U4848 (N_4848,In_147,In_627);
and U4849 (N_4849,In_709,In_564);
nand U4850 (N_4850,In_799,In_923);
nand U4851 (N_4851,In_836,In_553);
and U4852 (N_4852,In_148,In_167);
and U4853 (N_4853,In_651,In_199);
or U4854 (N_4854,In_318,In_455);
nand U4855 (N_4855,In_711,In_752);
nand U4856 (N_4856,In_546,In_891);
nor U4857 (N_4857,In_10,In_725);
and U4858 (N_4858,In_498,In_303);
or U4859 (N_4859,In_409,In_183);
nand U4860 (N_4860,In_661,In_216);
nor U4861 (N_4861,In_49,In_379);
nand U4862 (N_4862,In_590,In_525);
or U4863 (N_4863,In_4,In_406);
and U4864 (N_4864,In_203,In_157);
nor U4865 (N_4865,In_957,In_639);
and U4866 (N_4866,In_739,In_479);
nand U4867 (N_4867,In_660,In_491);
and U4868 (N_4868,In_764,In_499);
nor U4869 (N_4869,In_612,In_735);
nor U4870 (N_4870,In_948,In_270);
nand U4871 (N_4871,In_929,In_314);
and U4872 (N_4872,In_122,In_927);
and U4873 (N_4873,In_8,In_679);
and U4874 (N_4874,In_858,In_419);
nor U4875 (N_4875,In_453,In_329);
or U4876 (N_4876,In_499,In_296);
or U4877 (N_4877,In_224,In_264);
xnor U4878 (N_4878,In_77,In_906);
and U4879 (N_4879,In_650,In_284);
and U4880 (N_4880,In_690,In_184);
nor U4881 (N_4881,In_176,In_915);
nor U4882 (N_4882,In_969,In_234);
xor U4883 (N_4883,In_284,In_263);
or U4884 (N_4884,In_459,In_130);
or U4885 (N_4885,In_968,In_427);
and U4886 (N_4886,In_418,In_66);
nor U4887 (N_4887,In_333,In_721);
and U4888 (N_4888,In_153,In_444);
nor U4889 (N_4889,In_933,In_170);
or U4890 (N_4890,In_498,In_555);
and U4891 (N_4891,In_943,In_641);
and U4892 (N_4892,In_92,In_804);
nor U4893 (N_4893,In_726,In_438);
nor U4894 (N_4894,In_109,In_638);
nand U4895 (N_4895,In_348,In_112);
or U4896 (N_4896,In_71,In_938);
nand U4897 (N_4897,In_992,In_265);
nor U4898 (N_4898,In_990,In_208);
xor U4899 (N_4899,In_204,In_836);
or U4900 (N_4900,In_17,In_763);
nand U4901 (N_4901,In_961,In_718);
nor U4902 (N_4902,In_321,In_544);
or U4903 (N_4903,In_297,In_506);
and U4904 (N_4904,In_520,In_841);
nor U4905 (N_4905,In_612,In_310);
nand U4906 (N_4906,In_665,In_444);
nor U4907 (N_4907,In_232,In_287);
nor U4908 (N_4908,In_960,In_186);
or U4909 (N_4909,In_179,In_828);
nor U4910 (N_4910,In_318,In_790);
and U4911 (N_4911,In_528,In_362);
nand U4912 (N_4912,In_340,In_229);
and U4913 (N_4913,In_162,In_962);
xor U4914 (N_4914,In_465,In_596);
or U4915 (N_4915,In_597,In_96);
nand U4916 (N_4916,In_400,In_746);
nor U4917 (N_4917,In_778,In_737);
nor U4918 (N_4918,In_250,In_343);
or U4919 (N_4919,In_213,In_549);
xnor U4920 (N_4920,In_2,In_508);
nor U4921 (N_4921,In_642,In_635);
and U4922 (N_4922,In_709,In_118);
and U4923 (N_4923,In_244,In_788);
nand U4924 (N_4924,In_108,In_392);
nand U4925 (N_4925,In_693,In_997);
nand U4926 (N_4926,In_996,In_822);
or U4927 (N_4927,In_16,In_683);
or U4928 (N_4928,In_52,In_814);
xor U4929 (N_4929,In_813,In_279);
nand U4930 (N_4930,In_155,In_920);
or U4931 (N_4931,In_871,In_280);
nor U4932 (N_4932,In_478,In_993);
or U4933 (N_4933,In_42,In_681);
or U4934 (N_4934,In_151,In_696);
nor U4935 (N_4935,In_39,In_24);
nand U4936 (N_4936,In_791,In_95);
nand U4937 (N_4937,In_971,In_525);
nand U4938 (N_4938,In_31,In_702);
nor U4939 (N_4939,In_533,In_606);
and U4940 (N_4940,In_394,In_689);
nor U4941 (N_4941,In_798,In_631);
and U4942 (N_4942,In_791,In_731);
nor U4943 (N_4943,In_535,In_52);
nor U4944 (N_4944,In_906,In_682);
nor U4945 (N_4945,In_604,In_832);
and U4946 (N_4946,In_88,In_912);
nor U4947 (N_4947,In_132,In_642);
nand U4948 (N_4948,In_999,In_376);
or U4949 (N_4949,In_624,In_155);
nand U4950 (N_4950,In_262,In_810);
and U4951 (N_4951,In_578,In_444);
nand U4952 (N_4952,In_581,In_177);
or U4953 (N_4953,In_751,In_896);
nand U4954 (N_4954,In_640,In_272);
and U4955 (N_4955,In_770,In_121);
or U4956 (N_4956,In_212,In_854);
nand U4957 (N_4957,In_575,In_448);
or U4958 (N_4958,In_724,In_854);
and U4959 (N_4959,In_266,In_70);
nor U4960 (N_4960,In_488,In_773);
nand U4961 (N_4961,In_93,In_292);
nand U4962 (N_4962,In_767,In_69);
and U4963 (N_4963,In_521,In_900);
nand U4964 (N_4964,In_20,In_797);
nor U4965 (N_4965,In_96,In_820);
nor U4966 (N_4966,In_43,In_740);
nor U4967 (N_4967,In_700,In_942);
and U4968 (N_4968,In_701,In_350);
nor U4969 (N_4969,In_289,In_666);
nand U4970 (N_4970,In_637,In_677);
nand U4971 (N_4971,In_967,In_795);
nand U4972 (N_4972,In_674,In_630);
nor U4973 (N_4973,In_214,In_311);
and U4974 (N_4974,In_656,In_28);
nand U4975 (N_4975,In_401,In_94);
nand U4976 (N_4976,In_841,In_459);
nor U4977 (N_4977,In_123,In_796);
nor U4978 (N_4978,In_100,In_217);
nand U4979 (N_4979,In_174,In_922);
nand U4980 (N_4980,In_91,In_83);
nor U4981 (N_4981,In_675,In_455);
nand U4982 (N_4982,In_676,In_289);
and U4983 (N_4983,In_581,In_592);
nand U4984 (N_4984,In_239,In_563);
and U4985 (N_4985,In_784,In_235);
or U4986 (N_4986,In_327,In_601);
nand U4987 (N_4987,In_596,In_470);
nor U4988 (N_4988,In_902,In_615);
and U4989 (N_4989,In_570,In_583);
or U4990 (N_4990,In_566,In_689);
and U4991 (N_4991,In_958,In_963);
nand U4992 (N_4992,In_142,In_32);
xnor U4993 (N_4993,In_53,In_105);
nand U4994 (N_4994,In_871,In_382);
or U4995 (N_4995,In_311,In_770);
nor U4996 (N_4996,In_714,In_745);
nand U4997 (N_4997,In_849,In_771);
or U4998 (N_4998,In_405,In_318);
nand U4999 (N_4999,In_413,In_502);
or U5000 (N_5000,N_3443,N_3974);
or U5001 (N_5001,N_175,N_2870);
and U5002 (N_5002,N_2993,N_4687);
nand U5003 (N_5003,N_3206,N_4275);
or U5004 (N_5004,N_2953,N_780);
nor U5005 (N_5005,N_1159,N_2478);
or U5006 (N_5006,N_3970,N_4419);
and U5007 (N_5007,N_3652,N_4625);
or U5008 (N_5008,N_1180,N_4676);
or U5009 (N_5009,N_2711,N_4128);
and U5010 (N_5010,N_3382,N_712);
nand U5011 (N_5011,N_1178,N_3101);
nand U5012 (N_5012,N_3327,N_3370);
or U5013 (N_5013,N_3483,N_1068);
nand U5014 (N_5014,N_3339,N_287);
or U5015 (N_5015,N_2011,N_4018);
and U5016 (N_5016,N_2551,N_2607);
or U5017 (N_5017,N_1481,N_4445);
nor U5018 (N_5018,N_3631,N_3819);
and U5019 (N_5019,N_3980,N_726);
and U5020 (N_5020,N_2901,N_172);
nand U5021 (N_5021,N_4241,N_995);
nor U5022 (N_5022,N_3184,N_1256);
nand U5023 (N_5023,N_2097,N_3310);
nor U5024 (N_5024,N_2727,N_3222);
nand U5025 (N_5025,N_3262,N_4670);
and U5026 (N_5026,N_4347,N_2562);
and U5027 (N_5027,N_4292,N_2776);
nand U5028 (N_5028,N_1577,N_2396);
nor U5029 (N_5029,N_4796,N_4645);
nand U5030 (N_5030,N_1172,N_3848);
or U5031 (N_5031,N_2112,N_4455);
or U5032 (N_5032,N_4972,N_3984);
nor U5033 (N_5033,N_499,N_2881);
or U5034 (N_5034,N_2026,N_4284);
and U5035 (N_5035,N_2905,N_2247);
nor U5036 (N_5036,N_1800,N_2018);
nand U5037 (N_5037,N_316,N_4016);
nor U5038 (N_5038,N_4374,N_326);
or U5039 (N_5039,N_1297,N_3938);
and U5040 (N_5040,N_993,N_3643);
or U5041 (N_5041,N_3764,N_3473);
and U5042 (N_5042,N_1824,N_3426);
nor U5043 (N_5043,N_1326,N_1215);
and U5044 (N_5044,N_796,N_1455);
or U5045 (N_5045,N_1850,N_2684);
or U5046 (N_5046,N_2992,N_3889);
and U5047 (N_5047,N_4431,N_2348);
nand U5048 (N_5048,N_4742,N_3890);
nor U5049 (N_5049,N_2811,N_1301);
nor U5050 (N_5050,N_4504,N_4767);
xnor U5051 (N_5051,N_945,N_14);
and U5052 (N_5052,N_3562,N_1035);
nor U5053 (N_5053,N_3728,N_2340);
and U5054 (N_5054,N_1640,N_3045);
nand U5055 (N_5055,N_1737,N_4956);
or U5056 (N_5056,N_2998,N_1945);
xnor U5057 (N_5057,N_134,N_2492);
nor U5058 (N_5058,N_4780,N_3242);
nor U5059 (N_5059,N_4962,N_504);
nand U5060 (N_5060,N_1152,N_2165);
and U5061 (N_5061,N_1928,N_3857);
and U5062 (N_5062,N_782,N_74);
and U5063 (N_5063,N_1994,N_3670);
nor U5064 (N_5064,N_3903,N_120);
and U5065 (N_5065,N_4808,N_2922);
and U5066 (N_5066,N_2481,N_4614);
or U5067 (N_5067,N_4847,N_1637);
or U5068 (N_5068,N_2500,N_256);
nor U5069 (N_5069,N_3604,N_2140);
and U5070 (N_5070,N_606,N_4566);
nand U5071 (N_5071,N_2185,N_2154);
nor U5072 (N_5072,N_1106,N_2055);
and U5073 (N_5073,N_3065,N_4531);
or U5074 (N_5074,N_3041,N_1132);
and U5075 (N_5075,N_2847,N_3172);
nand U5076 (N_5076,N_4832,N_705);
or U5077 (N_5077,N_937,N_103);
and U5078 (N_5078,N_3605,N_1200);
and U5079 (N_5079,N_4945,N_1656);
xnor U5080 (N_5080,N_981,N_4436);
nor U5081 (N_5081,N_4203,N_3733);
nand U5082 (N_5082,N_2818,N_3695);
nor U5083 (N_5083,N_3132,N_37);
and U5084 (N_5084,N_1440,N_4496);
or U5085 (N_5085,N_1175,N_3480);
nand U5086 (N_5086,N_27,N_797);
or U5087 (N_5087,N_4405,N_3094);
or U5088 (N_5088,N_2136,N_1558);
and U5089 (N_5089,N_1907,N_4830);
or U5090 (N_5090,N_2316,N_4151);
and U5091 (N_5091,N_655,N_450);
nor U5092 (N_5092,N_1587,N_624);
and U5093 (N_5093,N_1211,N_405);
or U5094 (N_5094,N_2582,N_1);
nand U5095 (N_5095,N_2276,N_1602);
nor U5096 (N_5096,N_4433,N_3878);
nor U5097 (N_5097,N_832,N_1551);
and U5098 (N_5098,N_2131,N_2495);
nand U5099 (N_5099,N_3859,N_2969);
and U5100 (N_5100,N_3161,N_1920);
nand U5101 (N_5101,N_813,N_1729);
and U5102 (N_5102,N_3260,N_3667);
or U5103 (N_5103,N_4365,N_577);
or U5104 (N_5104,N_1310,N_2884);
nand U5105 (N_5105,N_2332,N_1545);
and U5106 (N_5106,N_2634,N_1606);
nand U5107 (N_5107,N_1259,N_264);
nand U5108 (N_5108,N_2898,N_3359);
nor U5109 (N_5109,N_2821,N_4589);
and U5110 (N_5110,N_2549,N_2401);
or U5111 (N_5111,N_2725,N_3781);
and U5112 (N_5112,N_2854,N_2312);
nand U5113 (N_5113,N_4593,N_4535);
or U5114 (N_5114,N_878,N_866);
nand U5115 (N_5115,N_58,N_858);
or U5116 (N_5116,N_3498,N_2911);
or U5117 (N_5117,N_3245,N_2469);
nand U5118 (N_5118,N_127,N_955);
nor U5119 (N_5119,N_1071,N_641);
or U5120 (N_5120,N_776,N_2490);
or U5121 (N_5121,N_756,N_2822);
or U5122 (N_5122,N_4314,N_790);
nor U5123 (N_5123,N_3055,N_1880);
nand U5124 (N_5124,N_3309,N_2861);
nor U5125 (N_5125,N_2566,N_1862);
nor U5126 (N_5126,N_4121,N_1216);
nor U5127 (N_5127,N_144,N_2690);
or U5128 (N_5128,N_3300,N_2016);
or U5129 (N_5129,N_4865,N_2516);
or U5130 (N_5130,N_1527,N_4929);
nand U5131 (N_5131,N_3545,N_483);
and U5132 (N_5132,N_4852,N_918);
and U5133 (N_5133,N_2614,N_1348);
and U5134 (N_5134,N_1380,N_2604);
nand U5135 (N_5135,N_3778,N_130);
nor U5136 (N_5136,N_2240,N_1779);
or U5137 (N_5137,N_2271,N_4541);
nand U5138 (N_5138,N_1258,N_1407);
and U5139 (N_5139,N_1472,N_2730);
and U5140 (N_5140,N_3739,N_1794);
nor U5141 (N_5141,N_4935,N_458);
or U5142 (N_5142,N_3745,N_2683);
or U5143 (N_5143,N_3662,N_136);
and U5144 (N_5144,N_2095,N_2245);
nor U5145 (N_5145,N_3989,N_3962);
nor U5146 (N_5146,N_2761,N_4007);
nor U5147 (N_5147,N_1869,N_4675);
nand U5148 (N_5148,N_4877,N_2246);
nor U5149 (N_5149,N_4751,N_4249);
and U5150 (N_5150,N_4940,N_3690);
or U5151 (N_5151,N_1955,N_1155);
nor U5152 (N_5152,N_4738,N_1377);
nor U5153 (N_5153,N_3634,N_4825);
and U5154 (N_5154,N_779,N_366);
or U5155 (N_5155,N_1365,N_2534);
and U5156 (N_5156,N_318,N_3455);
and U5157 (N_5157,N_2351,N_3806);
nand U5158 (N_5158,N_893,N_387);
and U5159 (N_5159,N_4991,N_2065);
nand U5160 (N_5160,N_3237,N_551);
and U5161 (N_5161,N_1055,N_2897);
and U5162 (N_5162,N_1921,N_1898);
nor U5163 (N_5163,N_1217,N_3356);
and U5164 (N_5164,N_1744,N_244);
nor U5165 (N_5165,N_3106,N_3911);
nand U5166 (N_5166,N_4286,N_2060);
nor U5167 (N_5167,N_4824,N_2793);
nor U5168 (N_5168,N_3429,N_4019);
or U5169 (N_5169,N_4305,N_924);
or U5170 (N_5170,N_1619,N_2256);
nand U5171 (N_5171,N_1784,N_923);
nor U5172 (N_5172,N_1636,N_4210);
or U5173 (N_5173,N_2651,N_1160);
nand U5174 (N_5174,N_1494,N_3821);
nand U5175 (N_5175,N_1074,N_3074);
and U5176 (N_5176,N_2278,N_3870);
nor U5177 (N_5177,N_3615,N_2813);
and U5178 (N_5178,N_3507,N_422);
nand U5179 (N_5179,N_2523,N_4047);
nor U5180 (N_5180,N_2184,N_1147);
nor U5181 (N_5181,N_1873,N_3759);
nor U5182 (N_5182,N_3828,N_642);
or U5183 (N_5183,N_791,N_4);
and U5184 (N_5184,N_2198,N_2708);
or U5185 (N_5185,N_4871,N_4976);
nand U5186 (N_5186,N_676,N_2941);
and U5187 (N_5187,N_3367,N_365);
and U5188 (N_5188,N_2522,N_668);
nand U5189 (N_5189,N_3230,N_2287);
or U5190 (N_5190,N_4639,N_4350);
nor U5191 (N_5191,N_1020,N_1290);
nor U5192 (N_5192,N_856,N_3969);
or U5193 (N_5193,N_30,N_1442);
and U5194 (N_5194,N_4409,N_12);
nor U5195 (N_5195,N_4234,N_714);
nor U5196 (N_5196,N_3121,N_804);
or U5197 (N_5197,N_2099,N_834);
and U5198 (N_5198,N_3597,N_2638);
and U5199 (N_5199,N_105,N_1177);
and U5200 (N_5200,N_1505,N_2641);
nand U5201 (N_5201,N_608,N_3246);
or U5202 (N_5202,N_2857,N_2594);
nor U5203 (N_5203,N_913,N_713);
nand U5204 (N_5204,N_2622,N_2034);
nand U5205 (N_5205,N_4612,N_3375);
and U5206 (N_5206,N_1449,N_930);
nand U5207 (N_5207,N_3433,N_3624);
nand U5208 (N_5208,N_3381,N_4366);
nor U5209 (N_5209,N_4402,N_1241);
or U5210 (N_5210,N_2294,N_4957);
or U5211 (N_5211,N_4147,N_3808);
nor U5212 (N_5212,N_1519,N_4490);
and U5213 (N_5213,N_2749,N_4897);
nor U5214 (N_5214,N_1446,N_1702);
or U5215 (N_5215,N_2239,N_3664);
and U5216 (N_5216,N_3353,N_1716);
or U5217 (N_5217,N_1401,N_2559);
and U5218 (N_5218,N_3823,N_4242);
or U5219 (N_5219,N_4046,N_4560);
or U5220 (N_5220,N_336,N_2028);
nor U5221 (N_5221,N_4831,N_4107);
and U5222 (N_5222,N_3713,N_2723);
or U5223 (N_5223,N_3398,N_117);
nor U5224 (N_5224,N_4231,N_2451);
and U5225 (N_5225,N_3743,N_972);
nand U5226 (N_5226,N_4885,N_2342);
or U5227 (N_5227,N_1003,N_3525);
or U5228 (N_5228,N_696,N_59);
xnor U5229 (N_5229,N_3145,N_182);
nor U5230 (N_5230,N_1239,N_3863);
nand U5231 (N_5231,N_512,N_1304);
or U5232 (N_5232,N_4067,N_1633);
or U5233 (N_5233,N_3686,N_2605);
nand U5234 (N_5234,N_1052,N_688);
nand U5235 (N_5235,N_691,N_2296);
nand U5236 (N_5236,N_1000,N_2611);
nor U5237 (N_5237,N_3136,N_1009);
nor U5238 (N_5238,N_4734,N_3419);
or U5239 (N_5239,N_4174,N_4201);
or U5240 (N_5240,N_652,N_1571);
or U5241 (N_5241,N_4728,N_1815);
or U5242 (N_5242,N_1727,N_4931);
nor U5243 (N_5243,N_2606,N_3154);
nor U5244 (N_5244,N_132,N_2688);
nand U5245 (N_5245,N_811,N_3193);
nor U5246 (N_5246,N_11,N_1684);
and U5247 (N_5247,N_3082,N_709);
nor U5248 (N_5248,N_2865,N_4761);
or U5249 (N_5249,N_833,N_386);
and U5250 (N_5250,N_958,N_4993);
nor U5251 (N_5251,N_2731,N_1166);
or U5252 (N_5252,N_4156,N_2387);
nor U5253 (N_5253,N_4892,N_1146);
nand U5254 (N_5254,N_575,N_4696);
nor U5255 (N_5255,N_4828,N_307);
nor U5256 (N_5256,N_2000,N_2568);
nor U5257 (N_5257,N_3166,N_2480);
or U5258 (N_5258,N_4100,N_2781);
nand U5259 (N_5259,N_2120,N_300);
or U5260 (N_5260,N_76,N_3089);
or U5261 (N_5261,N_4873,N_741);
nor U5262 (N_5262,N_4724,N_1162);
nand U5263 (N_5263,N_4634,N_3302);
and U5264 (N_5264,N_1228,N_4886);
and U5265 (N_5265,N_396,N_4766);
or U5266 (N_5266,N_3285,N_1432);
nand U5267 (N_5267,N_4605,N_2828);
or U5268 (N_5268,N_1411,N_1375);
nor U5269 (N_5269,N_4212,N_4494);
nand U5270 (N_5270,N_3772,N_1654);
and U5271 (N_5271,N_513,N_1661);
or U5272 (N_5272,N_508,N_3152);
nor U5273 (N_5273,N_2970,N_4966);
nor U5274 (N_5274,N_2827,N_4503);
and U5275 (N_5275,N_4500,N_2447);
and U5276 (N_5276,N_926,N_3040);
or U5277 (N_5277,N_1057,N_2915);
or U5278 (N_5278,N_232,N_1080);
and U5279 (N_5279,N_2610,N_2974);
nor U5280 (N_5280,N_3732,N_4530);
nor U5281 (N_5281,N_531,N_1047);
and U5282 (N_5282,N_1552,N_911);
or U5283 (N_5283,N_3740,N_2216);
and U5284 (N_5284,N_1087,N_3592);
and U5285 (N_5285,N_1930,N_410);
or U5286 (N_5286,N_1666,N_2843);
nand U5287 (N_5287,N_1987,N_1368);
nand U5288 (N_5288,N_1832,N_479);
and U5289 (N_5289,N_2473,N_2357);
nor U5290 (N_5290,N_891,N_3031);
nand U5291 (N_5291,N_3872,N_4334);
or U5292 (N_5292,N_61,N_1980);
nor U5293 (N_5293,N_230,N_4992);
nand U5294 (N_5294,N_4204,N_594);
and U5295 (N_5295,N_4272,N_306);
or U5296 (N_5296,N_3815,N_63);
nand U5297 (N_5297,N_3307,N_2300);
or U5298 (N_5298,N_670,N_1110);
nand U5299 (N_5299,N_1439,N_4418);
and U5300 (N_5300,N_1932,N_2472);
nor U5301 (N_5301,N_3407,N_1381);
nand U5302 (N_5302,N_272,N_277);
nand U5303 (N_5303,N_1818,N_54);
nand U5304 (N_5304,N_408,N_4768);
nor U5305 (N_5305,N_2710,N_2038);
nand U5306 (N_5306,N_2601,N_2106);
or U5307 (N_5307,N_4632,N_3033);
or U5308 (N_5308,N_4616,N_4983);
nand U5309 (N_5309,N_578,N_2207);
nand U5310 (N_5310,N_3163,N_4125);
and U5311 (N_5311,N_4792,N_3746);
nor U5312 (N_5312,N_1475,N_3060);
nor U5313 (N_5313,N_1791,N_83);
nand U5314 (N_5314,N_1409,N_963);
nand U5315 (N_5315,N_4096,N_4458);
nand U5316 (N_5316,N_2518,N_3936);
or U5317 (N_5317,N_2051,N_3199);
and U5318 (N_5318,N_4754,N_3767);
or U5319 (N_5319,N_1938,N_1740);
or U5320 (N_5320,N_1101,N_3174);
nor U5321 (N_5321,N_2874,N_2996);
and U5322 (N_5322,N_4222,N_4164);
nand U5323 (N_5323,N_3202,N_1329);
nand U5324 (N_5324,N_1685,N_494);
nor U5325 (N_5325,N_3044,N_4452);
nand U5326 (N_5326,N_3408,N_403);
nor U5327 (N_5327,N_4731,N_460);
nor U5328 (N_5328,N_2595,N_4951);
or U5329 (N_5329,N_3501,N_3973);
or U5330 (N_5330,N_4679,N_3757);
nor U5331 (N_5331,N_2766,N_1575);
nand U5332 (N_5332,N_4420,N_2100);
or U5333 (N_5333,N_1512,N_4225);
or U5334 (N_5334,N_4622,N_1051);
or U5335 (N_5335,N_3576,N_3410);
and U5336 (N_5336,N_3275,N_4099);
and U5337 (N_5337,N_2780,N_2524);
nor U5338 (N_5338,N_3918,N_3569);
nand U5339 (N_5339,N_3709,N_3494);
and U5340 (N_5340,N_4088,N_3452);
and U5341 (N_5341,N_3528,N_149);
and U5342 (N_5342,N_4556,N_1487);
xnor U5343 (N_5343,N_2629,N_4785);
or U5344 (N_5344,N_4706,N_2121);
or U5345 (N_5345,N_3614,N_3721);
and U5346 (N_5346,N_4540,N_2415);
and U5347 (N_5347,N_4006,N_1856);
or U5348 (N_5348,N_2274,N_4481);
and U5349 (N_5349,N_3156,N_3627);
or U5350 (N_5350,N_4089,N_1530);
nor U5351 (N_5351,N_3761,N_3876);
nor U5352 (N_5352,N_3578,N_2747);
or U5353 (N_5353,N_3608,N_456);
and U5354 (N_5354,N_1708,N_2751);
nand U5355 (N_5355,N_4689,N_1991);
nand U5356 (N_5356,N_2815,N_397);
nand U5357 (N_5357,N_1075,N_2588);
nand U5358 (N_5358,N_2712,N_3028);
nor U5359 (N_5359,N_910,N_3510);
and U5360 (N_5360,N_3929,N_125);
and U5361 (N_5361,N_3406,N_1183);
nand U5362 (N_5362,N_2410,N_4258);
nand U5363 (N_5363,N_219,N_587);
and U5364 (N_5364,N_4516,N_2226);
and U5365 (N_5365,N_1845,N_382);
nor U5366 (N_5366,N_4788,N_1711);
or U5367 (N_5367,N_1676,N_3682);
nor U5368 (N_5368,N_3742,N_1677);
or U5369 (N_5369,N_2254,N_3514);
nor U5370 (N_5370,N_3247,N_3794);
and U5371 (N_5371,N_3189,N_4414);
nor U5372 (N_5372,N_3651,N_4860);
or U5373 (N_5373,N_2691,N_3434);
nand U5374 (N_5374,N_3641,N_660);
nor U5375 (N_5375,N_4971,N_2868);
or U5376 (N_5376,N_475,N_1027);
and U5377 (N_5377,N_4457,N_2521);
nor U5378 (N_5378,N_2372,N_2114);
and U5379 (N_5379,N_2042,N_2275);
nor U5380 (N_5380,N_60,N_2738);
or U5381 (N_5381,N_2315,N_781);
nor U5382 (N_5382,N_2540,N_3798);
nor U5383 (N_5383,N_2616,N_36);
nor U5384 (N_5384,N_2252,N_323);
nand U5385 (N_5385,N_3020,N_1039);
or U5386 (N_5386,N_895,N_1400);
or U5387 (N_5387,N_1879,N_4341);
nand U5388 (N_5388,N_4319,N_1557);
or U5389 (N_5389,N_845,N_279);
nor U5390 (N_5390,N_2115,N_2942);
nand U5391 (N_5391,N_2334,N_4776);
nor U5392 (N_5392,N_583,N_2201);
nand U5393 (N_5393,N_444,N_2409);
nand U5394 (N_5394,N_186,N_275);
or U5395 (N_5395,N_1371,N_2264);
nor U5396 (N_5396,N_2758,N_3666);
and U5397 (N_5397,N_1145,N_4671);
xor U5398 (N_5398,N_2900,N_1788);
nor U5399 (N_5399,N_4941,N_1761);
nor U5400 (N_5400,N_3617,N_3553);
nand U5401 (N_5401,N_3414,N_4545);
or U5402 (N_5402,N_1315,N_3684);
or U5403 (N_5403,N_138,N_4185);
nand U5404 (N_5404,N_4674,N_2541);
nor U5405 (N_5405,N_4802,N_141);
or U5406 (N_5406,N_4783,N_2117);
or U5407 (N_5407,N_4590,N_3413);
nor U5408 (N_5408,N_3344,N_3960);
nor U5409 (N_5409,N_4399,N_2452);
nand U5410 (N_5410,N_784,N_3008);
and U5411 (N_5411,N_975,N_3844);
nand U5412 (N_5412,N_1291,N_1628);
nand U5413 (N_5413,N_2966,N_1163);
nor U5414 (N_5414,N_4032,N_2726);
and U5415 (N_5415,N_4926,N_4188);
and U5416 (N_5416,N_2146,N_2531);
and U5417 (N_5417,N_1975,N_1648);
nor U5418 (N_5418,N_1870,N_2448);
nand U5419 (N_5419,N_179,N_4663);
and U5420 (N_5420,N_3793,N_2005);
nand U5421 (N_5421,N_2555,N_2772);
nor U5422 (N_5422,N_4838,N_909);
and U5423 (N_5423,N_4685,N_562);
nand U5424 (N_5424,N_1034,N_560);
or U5425 (N_5425,N_3602,N_3037);
and U5426 (N_5426,N_139,N_1427);
xor U5427 (N_5427,N_196,N_3807);
nor U5428 (N_5428,N_2831,N_1863);
nand U5429 (N_5429,N_4289,N_4138);
or U5430 (N_5430,N_476,N_2374);
nor U5431 (N_5431,N_346,N_4329);
nand U5432 (N_5432,N_3025,N_1060);
nand U5433 (N_5433,N_1583,N_4757);
and U5434 (N_5434,N_4143,N_1940);
nand U5435 (N_5435,N_4596,N_1668);
nand U5436 (N_5436,N_4369,N_1005);
or U5437 (N_5437,N_886,N_2875);
nor U5438 (N_5438,N_4421,N_916);
nor U5439 (N_5439,N_4661,N_4401);
nor U5440 (N_5440,N_4461,N_601);
nand U5441 (N_5441,N_4519,N_4577);
and U5442 (N_5442,N_2160,N_2093);
nand U5443 (N_5443,N_1169,N_4964);
or U5444 (N_5444,N_4740,N_880);
or U5445 (N_5445,N_2122,N_2754);
and U5446 (N_5446,N_592,N_1939);
nor U5447 (N_5447,N_372,N_1812);
nand U5448 (N_5448,N_2389,N_1548);
and U5449 (N_5449,N_4837,N_471);
nand U5450 (N_5450,N_4732,N_347);
and U5451 (N_5451,N_3536,N_505);
xor U5452 (N_5452,N_4554,N_708);
or U5453 (N_5453,N_2670,N_448);
nand U5454 (N_5454,N_481,N_1193);
or U5455 (N_5455,N_2685,N_2603);
nand U5456 (N_5456,N_3391,N_889);
nor U5457 (N_5457,N_4017,N_3591);
nor U5458 (N_5458,N_2260,N_2043);
nand U5459 (N_5459,N_638,N_4235);
nand U5460 (N_5460,N_1313,N_1396);
or U5461 (N_5461,N_500,N_459);
xnor U5462 (N_5462,N_2686,N_4563);
nand U5463 (N_5463,N_2623,N_1688);
and U5464 (N_5464,N_2295,N_4071);
nor U5465 (N_5465,N_4758,N_3477);
nand U5466 (N_5466,N_3446,N_4717);
nand U5467 (N_5467,N_1680,N_2999);
or U5468 (N_5468,N_812,N_4898);
nor U5469 (N_5469,N_2569,N_4909);
nor U5470 (N_5470,N_3268,N_3964);
and U5471 (N_5471,N_4442,N_2598);
nand U5472 (N_5472,N_4550,N_3751);
nor U5473 (N_5473,N_1953,N_4131);
nand U5474 (N_5474,N_1993,N_3365);
nor U5475 (N_5475,N_3683,N_3629);
and U5476 (N_5476,N_2666,N_2775);
nand U5477 (N_5477,N_4736,N_3000);
nor U5478 (N_5478,N_3255,N_4132);
nand U5479 (N_5479,N_566,N_687);
and U5480 (N_5480,N_4066,N_2362);
nand U5481 (N_5481,N_4763,N_29);
nand U5482 (N_5482,N_2398,N_4741);
nor U5483 (N_5483,N_229,N_976);
and U5484 (N_5484,N_1370,N_3702);
nand U5485 (N_5485,N_1140,N_1501);
nor U5486 (N_5486,N_3706,N_747);
nand U5487 (N_5487,N_4599,N_1434);
and U5488 (N_5488,N_4655,N_1626);
or U5489 (N_5489,N_2098,N_5);
nor U5490 (N_5490,N_2162,N_999);
nand U5491 (N_5491,N_3869,N_698);
and U5492 (N_5492,N_2113,N_4601);
nor U5493 (N_5493,N_4512,N_4382);
or U5494 (N_5494,N_2019,N_2001);
nor U5495 (N_5495,N_1268,N_3535);
and U5496 (N_5496,N_574,N_4975);
nor U5497 (N_5497,N_2774,N_1810);
and U5498 (N_5498,N_2816,N_2002);
or U5499 (N_5499,N_1032,N_735);
and U5500 (N_5500,N_4980,N_1883);
nand U5501 (N_5501,N_1531,N_2546);
nor U5502 (N_5502,N_489,N_1363);
nor U5503 (N_5503,N_2926,N_2411);
or U5504 (N_5504,N_4406,N_1949);
nor U5505 (N_5505,N_1762,N_1342);
or U5506 (N_5506,N_4184,N_1474);
nor U5507 (N_5507,N_827,N_4858);
or U5508 (N_5508,N_3780,N_4943);
or U5509 (N_5509,N_616,N_1164);
and U5510 (N_5510,N_3420,N_4580);
nor U5511 (N_5511,N_1963,N_1422);
nand U5512 (N_5512,N_514,N_1923);
nor U5513 (N_5513,N_1480,N_4509);
nor U5514 (N_5514,N_534,N_3467);
nand U5515 (N_5515,N_3990,N_4288);
and U5516 (N_5516,N_1157,N_4137);
and U5517 (N_5517,N_4228,N_3866);
or U5518 (N_5518,N_2350,N_1222);
nor U5519 (N_5519,N_1458,N_2885);
nor U5520 (N_5520,N_3099,N_135);
nand U5521 (N_5521,N_4364,N_265);
nand U5522 (N_5522,N_4283,N_3523);
nand U5523 (N_5523,N_1891,N_1141);
or U5524 (N_5524,N_2158,N_2647);
or U5525 (N_5525,N_226,N_4623);
nor U5526 (N_5526,N_2663,N_1192);
and U5527 (N_5527,N_4301,N_1059);
xor U5528 (N_5528,N_4705,N_710);
nand U5529 (N_5529,N_922,N_1105);
nand U5530 (N_5530,N_697,N_1260);
and U5531 (N_5531,N_3565,N_1604);
nand U5532 (N_5532,N_1042,N_4487);
or U5533 (N_5533,N_3810,N_3850);
or U5534 (N_5534,N_2429,N_2208);
and U5535 (N_5535,N_736,N_1817);
nor U5536 (N_5536,N_3383,N_4001);
nor U5537 (N_5537,N_4394,N_195);
and U5538 (N_5538,N_527,N_580);
nand U5539 (N_5539,N_2227,N_2058);
nand U5540 (N_5540,N_1002,N_1094);
nand U5541 (N_5541,N_3995,N_728);
and U5542 (N_5542,N_4627,N_2105);
or U5543 (N_5543,N_4846,N_2850);
and U5544 (N_5544,N_1097,N_795);
and U5545 (N_5545,N_1859,N_3933);
or U5546 (N_5546,N_1459,N_748);
and U5547 (N_5547,N_3376,N_760);
and U5548 (N_5548,N_537,N_1821);
or U5549 (N_5549,N_4899,N_4393);
nand U5550 (N_5550,N_3203,N_3920);
nand U5551 (N_5551,N_4404,N_2442);
or U5552 (N_5552,N_2759,N_4062);
and U5553 (N_5553,N_407,N_4063);
nand U5554 (N_5554,N_3063,N_2943);
and U5555 (N_5555,N_3871,N_2672);
nor U5556 (N_5556,N_2482,N_1232);
or U5557 (N_5557,N_2570,N_1154);
nor U5558 (N_5558,N_209,N_2778);
nor U5559 (N_5559,N_4323,N_3053);
nor U5560 (N_5560,N_3011,N_280);
or U5561 (N_5561,N_4355,N_635);
or U5562 (N_5562,N_178,N_3648);
nand U5563 (N_5563,N_902,N_818);
nand U5564 (N_5564,N_3186,N_4986);
and U5565 (N_5565,N_2318,N_3500);
and U5566 (N_5566,N_48,N_903);
nor U5567 (N_5567,N_2925,N_4397);
and U5568 (N_5568,N_722,N_4699);
or U5569 (N_5569,N_1369,N_3577);
and U5570 (N_5570,N_4604,N_53);
and U5571 (N_5571,N_4948,N_2373);
and U5572 (N_5572,N_3660,N_3762);
and U5573 (N_5573,N_3860,N_2762);
nor U5574 (N_5574,N_1317,N_4715);
nand U5575 (N_5575,N_3803,N_4324);
nor U5576 (N_5576,N_4022,N_1168);
nand U5577 (N_5577,N_4160,N_4984);
nand U5578 (N_5578,N_338,N_581);
and U5579 (N_5579,N_4070,N_140);
nor U5580 (N_5580,N_3428,N_2346);
nor U5581 (N_5581,N_1943,N_4815);
nor U5582 (N_5582,N_767,N_4023);
or U5583 (N_5583,N_3379,N_3265);
and U5584 (N_5584,N_2196,N_3979);
nand U5585 (N_5585,N_2225,N_3093);
or U5586 (N_5586,N_3491,N_4779);
and U5587 (N_5587,N_2840,N_3522);
or U5588 (N_5588,N_4223,N_1790);
nor U5589 (N_5589,N_1756,N_851);
nor U5590 (N_5590,N_4459,N_806);
nand U5591 (N_5591,N_118,N_1414);
and U5592 (N_5592,N_2963,N_2491);
or U5593 (N_5593,N_2560,N_3766);
or U5594 (N_5594,N_246,N_4408);
nand U5595 (N_5595,N_1743,N_4575);
nand U5596 (N_5596,N_2917,N_3546);
and U5597 (N_5597,N_3114,N_3179);
and U5598 (N_5598,N_4340,N_4801);
or U5599 (N_5599,N_3516,N_389);
and U5600 (N_5600,N_1293,N_4666);
or U5601 (N_5601,N_4011,N_4267);
or U5602 (N_5602,N_3061,N_2344);
and U5603 (N_5603,N_2356,N_3517);
or U5604 (N_5604,N_2037,N_2565);
or U5605 (N_5605,N_1410,N_3291);
or U5606 (N_5606,N_4692,N_4480);
nor U5607 (N_5607,N_1428,N_4643);
nor U5608 (N_5608,N_1186,N_314);
nor U5609 (N_5609,N_2866,N_2767);
or U5610 (N_5610,N_992,N_2972);
and U5611 (N_5611,N_1423,N_4139);
xor U5612 (N_5612,N_2199,N_2657);
nor U5613 (N_5613,N_455,N_820);
nand U5614 (N_5614,N_904,N_1782);
or U5615 (N_5615,N_73,N_1805);
nor U5616 (N_5616,N_2581,N_2845);
nand U5617 (N_5617,N_80,N_2982);
or U5618 (N_5618,N_3100,N_2771);
nand U5619 (N_5619,N_1906,N_2558);
nand U5620 (N_5620,N_1436,N_3372);
nand U5621 (N_5621,N_3883,N_3315);
nor U5622 (N_5622,N_4168,N_3665);
xnor U5623 (N_5623,N_2052,N_1622);
nor U5624 (N_5624,N_3418,N_369);
nor U5625 (N_5625,N_3688,N_1251);
and U5626 (N_5626,N_987,N_378);
nand U5627 (N_5627,N_3143,N_3158);
nand U5628 (N_5628,N_1892,N_3812);
and U5629 (N_5629,N_4921,N_1629);
nand U5630 (N_5630,N_4733,N_3185);
and U5631 (N_5631,N_4484,N_778);
nor U5632 (N_5632,N_3588,N_350);
or U5633 (N_5633,N_1764,N_3924);
or U5634 (N_5634,N_1798,N_1406);
and U5635 (N_5635,N_3397,N_720);
and U5636 (N_5636,N_4735,N_4638);
nor U5637 (N_5637,N_3583,N_2292);
or U5638 (N_5638,N_2326,N_2814);
nand U5639 (N_5639,N_4528,N_3852);
nor U5640 (N_5640,N_3105,N_1662);
nor U5641 (N_5641,N_596,N_840);
nand U5642 (N_5642,N_4179,N_825);
nand U5643 (N_5643,N_3693,N_4040);
nand U5644 (N_5644,N_968,N_3947);
nand U5645 (N_5645,N_2143,N_3953);
or U5646 (N_5646,N_4515,N_284);
or U5647 (N_5647,N_4498,N_2659);
nand U5648 (N_5648,N_2147,N_200);
and U5649 (N_5649,N_2538,N_1015);
nor U5650 (N_5650,N_2740,N_2231);
or U5651 (N_5651,N_1714,N_2674);
nand U5652 (N_5652,N_4471,N_1829);
nand U5653 (N_5653,N_2552,N_1483);
nand U5654 (N_5654,N_385,N_4015);
nand U5655 (N_5655,N_876,N_4300);
and U5656 (N_5656,N_519,N_707);
nand U5657 (N_5657,N_3405,N_2682);
and U5658 (N_5658,N_570,N_3563);
nor U5659 (N_5659,N_3320,N_1934);
nand U5660 (N_5660,N_1240,N_2249);
nor U5661 (N_5661,N_2343,N_4224);
or U5662 (N_5662,N_4262,N_3646);
nand U5663 (N_5663,N_3590,N_3625);
nor U5664 (N_5664,N_617,N_2177);
or U5665 (N_5665,N_3554,N_593);
nor U5666 (N_5666,N_45,N_2211);
nand U5667 (N_5667,N_1524,N_496);
or U5668 (N_5668,N_1300,N_4237);
or U5669 (N_5669,N_4844,N_4771);
nand U5670 (N_5670,N_3775,N_3396);
and U5671 (N_5671,N_3293,N_4908);
nand U5672 (N_5672,N_4360,N_3904);
and U5673 (N_5673,N_3120,N_563);
and U5674 (N_5674,N_4973,N_2062);
nand U5675 (N_5675,N_2689,N_2180);
nand U5676 (N_5676,N_1710,N_984);
or U5677 (N_5677,N_1792,N_2989);
and U5678 (N_5678,N_176,N_1759);
and U5679 (N_5679,N_1470,N_730);
and U5680 (N_5680,N_1012,N_19);
nand U5681 (N_5681,N_4571,N_831);
or U5682 (N_5682,N_3575,N_1497);
or U5683 (N_5683,N_3016,N_3873);
nor U5684 (N_5684,N_2844,N_672);
xor U5685 (N_5685,N_3714,N_1367);
or U5686 (N_5686,N_1273,N_2450);
xor U5687 (N_5687,N_2206,N_2745);
and U5688 (N_5688,N_337,N_4477);
and U5689 (N_5689,N_2561,N_967);
nor U5690 (N_5690,N_1111,N_158);
or U5691 (N_5691,N_4875,N_4118);
nand U5692 (N_5692,N_3972,N_2054);
and U5693 (N_5693,N_57,N_4920);
and U5694 (N_5694,N_3897,N_1617);
nand U5695 (N_5695,N_1874,N_2465);
nor U5696 (N_5696,N_4558,N_4887);
nand U5697 (N_5697,N_1539,N_3613);
and U5698 (N_5698,N_4486,N_4669);
nor U5699 (N_5699,N_2200,N_1245);
nor U5700 (N_5700,N_4805,N_3888);
nor U5701 (N_5701,N_3140,N_2585);
or U5702 (N_5702,N_3305,N_4370);
or U5703 (N_5703,N_2640,N_1220);
or U5704 (N_5704,N_4906,N_4136);
or U5705 (N_5705,N_2134,N_222);
or U5706 (N_5706,N_1072,N_2694);
nor U5707 (N_5707,N_2487,N_1965);
nand U5708 (N_5708,N_2156,N_253);
or U5709 (N_5709,N_2625,N_2798);
xnor U5710 (N_5710,N_355,N_1670);
nor U5711 (N_5711,N_2234,N_964);
or U5712 (N_5712,N_1757,N_2528);
nor U5713 (N_5713,N_1871,N_4398);
nor U5714 (N_5714,N_2337,N_683);
or U5715 (N_5715,N_3943,N_842);
nor U5716 (N_5716,N_3109,N_1901);
nand U5717 (N_5717,N_618,N_42);
or U5718 (N_5718,N_4764,N_4192);
nor U5719 (N_5719,N_1749,N_4009);
nand U5720 (N_5720,N_2457,N_4748);
or U5721 (N_5721,N_507,N_1738);
nor U5722 (N_5722,N_4633,N_4045);
nor U5723 (N_5723,N_807,N_2855);
nor U5724 (N_5724,N_2191,N_869);
and U5725 (N_5725,N_1144,N_4915);
and U5726 (N_5726,N_4183,N_3950);
and U5727 (N_5727,N_304,N_1195);
nor U5728 (N_5728,N_66,N_114);
nand U5729 (N_5729,N_361,N_1701);
or U5730 (N_5730,N_1773,N_2126);
or U5731 (N_5731,N_3551,N_1130);
nand U5732 (N_5732,N_3123,N_3997);
nand U5733 (N_5733,N_4848,N_2152);
and U5734 (N_5734,N_4356,N_695);
and U5735 (N_5735,N_4456,N_506);
or U5736 (N_5736,N_217,N_2434);
nor U5737 (N_5737,N_4000,N_3326);
nor U5738 (N_5738,N_2536,N_4995);
or U5739 (N_5739,N_4432,N_1373);
nand U5740 (N_5740,N_803,N_351);
or U5741 (N_5741,N_4255,N_4804);
or U5742 (N_5742,N_4325,N_3809);
and U5743 (N_5743,N_324,N_2338);
nor U5744 (N_5744,N_2413,N_2498);
nor U5745 (N_5745,N_2912,N_2354);
nor U5746 (N_5746,N_1615,N_4059);
nand U5747 (N_5747,N_1090,N_977);
nor U5748 (N_5748,N_328,N_4043);
and U5749 (N_5749,N_261,N_4119);
nand U5750 (N_5750,N_4389,N_379);
or U5751 (N_5751,N_934,N_1206);
and U5752 (N_5752,N_2222,N_4576);
and U5753 (N_5753,N_1452,N_3113);
and U5754 (N_5754,N_2994,N_2737);
and U5755 (N_5755,N_250,N_109);
and U5756 (N_5756,N_3760,N_3080);
nand U5757 (N_5757,N_520,N_1843);
xnor U5758 (N_5758,N_1777,N_3478);
and U5759 (N_5759,N_4158,N_529);
and U5760 (N_5760,N_3650,N_692);
and U5761 (N_5761,N_4977,N_663);
nor U5762 (N_5762,N_2391,N_3773);
or U5763 (N_5763,N_2515,N_1624);
nor U5764 (N_5764,N_585,N_104);
and U5765 (N_5765,N_2946,N_3463);
nand U5766 (N_5766,N_1150,N_234);
nand U5767 (N_5767,N_4229,N_4690);
nand U5768 (N_5768,N_4197,N_556);
and U5769 (N_5769,N_965,N_3159);
and U5770 (N_5770,N_775,N_941);
nor U5771 (N_5771,N_2809,N_3280);
and U5772 (N_5772,N_1108,N_1352);
or U5773 (N_5773,N_3734,N_3010);
and U5774 (N_5774,N_586,N_155);
nand U5775 (N_5775,N_3308,N_4507);
nand U5776 (N_5776,N_218,N_108);
nor U5777 (N_5777,N_947,N_828);
nor U5778 (N_5778,N_2236,N_2212);
nor U5779 (N_5779,N_3017,N_1210);
nand U5780 (N_5780,N_1208,N_2700);
and U5781 (N_5781,N_686,N_3930);
nor U5782 (N_5782,N_4020,N_1589);
nor U5783 (N_5783,N_1056,N_2909);
nand U5784 (N_5784,N_4981,N_919);
and U5785 (N_5785,N_4219,N_1642);
and U5786 (N_5786,N_3620,N_1627);
or U5787 (N_5787,N_3699,N_4075);
nand U5788 (N_5788,N_1058,N_165);
or U5789 (N_5789,N_3630,N_2084);
nand U5790 (N_5790,N_1104,N_393);
and U5791 (N_5791,N_3070,N_2376);
or U5792 (N_5792,N_3574,N_4523);
nor U5793 (N_5793,N_3529,N_2799);
nand U5794 (N_5794,N_3538,N_564);
or U5795 (N_5795,N_3839,N_848);
nor U5796 (N_5796,N_1511,N_2835);
nand U5797 (N_5797,N_1667,N_1468);
nor U5798 (N_5798,N_1588,N_400);
or U5799 (N_5799,N_2041,N_210);
nand U5800 (N_5800,N_2483,N_849);
or U5801 (N_5801,N_2349,N_4533);
nand U5802 (N_5802,N_1437,N_3824);
nor U5803 (N_5803,N_1610,N_932);
nor U5804 (N_5804,N_1223,N_3236);
and U5805 (N_5805,N_262,N_4230);
and U5806 (N_5806,N_743,N_644);
nand U5807 (N_5807,N_2864,N_4363);
or U5808 (N_5808,N_3566,N_1465);
nor U5809 (N_5809,N_95,N_152);
or U5810 (N_5810,N_4548,N_2443);
nand U5811 (N_5811,N_4620,N_4817);
nor U5812 (N_5812,N_2586,N_4726);
nand U5813 (N_5813,N_1231,N_3378);
nand U5814 (N_5814,N_4791,N_2834);
nor U5815 (N_5815,N_2235,N_896);
nand U5816 (N_5816,N_33,N_1786);
nor U5817 (N_5817,N_765,N_985);
nor U5818 (N_5818,N_296,N_1807);
nand U5819 (N_5819,N_675,N_1698);
and U5820 (N_5820,N_2488,N_308);
nor U5821 (N_5821,N_1353,N_2223);
or U5822 (N_5822,N_774,N_3847);
nand U5823 (N_5823,N_1844,N_4553);
and U5824 (N_5824,N_2921,N_4911);
nand U5825 (N_5825,N_900,N_1438);
or U5826 (N_5826,N_3243,N_3350);
or U5827 (N_5827,N_417,N_2453);
and U5828 (N_5828,N_2263,N_3654);
and U5829 (N_5829,N_4745,N_2291);
nand U5830 (N_5830,N_4178,N_1896);
nand U5831 (N_5831,N_4647,N_208);
nand U5832 (N_5832,N_2554,N_3907);
or U5833 (N_5833,N_8,N_997);
nand U5834 (N_5834,N_2892,N_3254);
and U5835 (N_5835,N_85,N_1019);
nand U5836 (N_5836,N_4819,N_2503);
nor U5837 (N_5837,N_4205,N_4569);
or U5838 (N_5838,N_2829,N_462);
or U5839 (N_5839,N_1121,N_1608);
nor U5840 (N_5840,N_751,N_4033);
nand U5841 (N_5841,N_1522,N_3362);
and U5842 (N_5842,N_415,N_3559);
and U5843 (N_5843,N_1593,N_1201);
nor U5844 (N_5844,N_4057,N_1490);
nand U5845 (N_5845,N_4664,N_2303);
and U5846 (N_5846,N_4681,N_3676);
and U5847 (N_5847,N_2430,N_2405);
and U5848 (N_5848,N_439,N_2388);
or U5849 (N_5849,N_463,N_2192);
nand U5850 (N_5850,N_1196,N_290);
nor U5851 (N_5851,N_1248,N_4232);
nand U5852 (N_5852,N_3050,N_4221);
and U5853 (N_5853,N_1246,N_3282);
or U5854 (N_5854,N_1357,N_1281);
nand U5855 (N_5855,N_406,N_4799);
nor U5856 (N_5856,N_6,N_3609);
or U5857 (N_5857,N_2907,N_3217);
or U5858 (N_5858,N_3330,N_4893);
nor U5859 (N_5859,N_1809,N_3877);
or U5860 (N_5860,N_1521,N_3225);
and U5861 (N_5861,N_3024,N_819);
nand U5862 (N_5862,N_3448,N_2456);
nand U5863 (N_5863,N_847,N_3226);
nor U5864 (N_5864,N_4083,N_3486);
nor U5865 (N_5865,N_3084,N_2049);
nand U5866 (N_5866,N_436,N_4826);
nor U5867 (N_5867,N_2703,N_390);
nor U5868 (N_5868,N_2382,N_2139);
nand U5869 (N_5869,N_4239,N_1116);
and U5870 (N_5870,N_432,N_1046);
or U5871 (N_5871,N_4211,N_1878);
nand U5872 (N_5872,N_1537,N_2671);
nor U5873 (N_5873,N_1509,N_1050);
or U5874 (N_5874,N_4924,N_794);
or U5875 (N_5875,N_4279,N_523);
or U5876 (N_5876,N_4439,N_1271);
and U5877 (N_5877,N_1804,N_4508);
and U5878 (N_5878,N_4322,N_443);
or U5879 (N_5879,N_3502,N_4214);
or U5880 (N_5880,N_3073,N_4371);
nand U5881 (N_5881,N_2927,N_3657);
nand U5882 (N_5882,N_952,N_3496);
or U5883 (N_5883,N_3299,N_888);
or U5884 (N_5884,N_4628,N_2692);
nand U5885 (N_5885,N_4561,N_1203);
nor U5886 (N_5886,N_3840,N_3377);
or U5887 (N_5887,N_4318,N_1614);
or U5888 (N_5888,N_787,N_733);
and U5889 (N_5889,N_3219,N_3244);
or U5890 (N_5890,N_3616,N_3795);
nor U5891 (N_5891,N_690,N_4998);
nand U5892 (N_5892,N_503,N_3306);
nor U5893 (N_5893,N_1793,N_2046);
or U5894 (N_5894,N_2741,N_3416);
nand U5895 (N_5895,N_2807,N_3898);
or U5896 (N_5896,N_3490,N_437);
or U5897 (N_5897,N_761,N_4444);
and U5898 (N_5898,N_1946,N_4381);
and U5899 (N_5899,N_1758,N_3891);
nand U5900 (N_5900,N_1204,N_3825);
nor U5901 (N_5901,N_1412,N_4207);
or U5902 (N_5902,N_3599,N_4198);
or U5903 (N_5903,N_173,N_3048);
nand U5904 (N_5904,N_928,N_2612);
nor U5905 (N_5905,N_451,N_3301);
or U5906 (N_5906,N_1568,N_3552);
or U5907 (N_5907,N_2363,N_4965);
nor U5908 (N_5908,N_4954,N_3354);
nor U5909 (N_5909,N_2257,N_3831);
or U5910 (N_5910,N_3432,N_700);
and U5911 (N_5911,N_1387,N_3727);
and U5912 (N_5912,N_3313,N_2186);
nand U5913 (N_5913,N_3926,N_1335);
nand U5914 (N_5914,N_2313,N_912);
and U5915 (N_5915,N_1725,N_2768);
nand U5916 (N_5916,N_3484,N_4642);
nand U5917 (N_5917,N_4693,N_3311);
nor U5918 (N_5918,N_3176,N_1433);
nor U5919 (N_5919,N_3270,N_2288);
nand U5920 (N_5920,N_2722,N_4181);
nor U5921 (N_5921,N_557,N_2981);
nor U5922 (N_5922,N_3191,N_4722);
nand U5923 (N_5923,N_1594,N_664);
nor U5924 (N_5924,N_2244,N_98);
and U5925 (N_5925,N_850,N_399);
and U5926 (N_5926,N_942,N_3137);
nand U5927 (N_5927,N_1238,N_97);
and U5928 (N_5928,N_561,N_3438);
or U5929 (N_5929,N_3965,N_498);
nand U5930 (N_5930,N_4227,N_4428);
nor U5931 (N_5931,N_1705,N_1999);
or U5932 (N_5932,N_3865,N_18);
nor U5933 (N_5933,N_1219,N_988);
nor U5934 (N_5934,N_4772,N_1279);
and U5935 (N_5935,N_1650,N_1482);
and U5936 (N_5936,N_4209,N_2251);
nand U5937 (N_5937,N_1499,N_2736);
or U5938 (N_5938,N_3036,N_1734);
or U5939 (N_5939,N_1362,N_4154);
and U5940 (N_5940,N_2395,N_3437);
or U5941 (N_5941,N_521,N_1767);
or U5942 (N_5942,N_729,N_2331);
or U5943 (N_5943,N_2102,N_1603);
and U5944 (N_5944,N_2204,N_2760);
and U5945 (N_5945,N_3568,N_424);
and U5946 (N_5946,N_2895,N_122);
nor U5947 (N_5947,N_283,N_3687);
nor U5948 (N_5948,N_2646,N_1523);
nand U5949 (N_5949,N_1886,N_2377);
and U5950 (N_5950,N_633,N_2130);
or U5951 (N_5951,N_255,N_1471);
nor U5952 (N_5952,N_3987,N_93);
nor U5953 (N_5953,N_1855,N_846);
or U5954 (N_5954,N_4737,N_2658);
nand U5955 (N_5955,N_258,N_452);
and U5956 (N_5956,N_4747,N_2979);
and U5957 (N_5957,N_1112,N_2510);
or U5958 (N_5958,N_4328,N_626);
nor U5959 (N_5959,N_1851,N_2393);
and U5960 (N_5960,N_1276,N_4248);
xnor U5961 (N_5961,N_2111,N_4123);
nand U5962 (N_5962,N_4859,N_1720);
nor U5963 (N_5963,N_613,N_658);
and U5964 (N_5964,N_62,N_4567);
nor U5965 (N_5965,N_1026,N_4862);
or U5966 (N_5966,N_1283,N_2101);
and U5967 (N_5967,N_4526,N_357);
nand U5968 (N_5968,N_1795,N_1579);
xnor U5969 (N_5969,N_2036,N_3661);
nor U5970 (N_5970,N_1171,N_2526);
nor U5971 (N_5971,N_2779,N_1540);
or U5972 (N_5972,N_3487,N_2833);
and U5973 (N_5973,N_3636,N_879);
nor U5974 (N_5974,N_2678,N_4814);
nand U5975 (N_5975,N_192,N_4277);
xor U5976 (N_5976,N_2944,N_510);
nand U5977 (N_5977,N_3967,N_2951);
and U5978 (N_5978,N_4144,N_3038);
nand U5979 (N_5979,N_96,N_2379);
nor U5980 (N_5980,N_1445,N_4048);
or U5981 (N_5981,N_3298,N_3548);
or U5982 (N_5982,N_4104,N_2717);
and U5983 (N_5983,N_1227,N_1613);
and U5984 (N_5984,N_1914,N_885);
and U5985 (N_5985,N_727,N_4881);
nor U5986 (N_5986,N_1919,N_983);
or U5987 (N_5987,N_685,N_1467);
nor U5988 (N_5988,N_4529,N_1644);
nor U5989 (N_5989,N_4261,N_4437);
or U5990 (N_5990,N_1866,N_4266);
or U5991 (N_5991,N_1925,N_605);
nor U5992 (N_5992,N_3263,N_4390);
nor U5993 (N_5993,N_4163,N_1405);
and U5994 (N_5994,N_3035,N_3141);
nor U5995 (N_5995,N_3064,N_1100);
nand U5996 (N_5996,N_1674,N_3983);
nor U5997 (N_5997,N_569,N_362);
nor U5998 (N_5998,N_1393,N_1573);
and U5999 (N_5999,N_4856,N_4760);
and U6000 (N_6000,N_1093,N_2321);
and U6001 (N_6001,N_2218,N_4343);
nor U6002 (N_6002,N_1823,N_2985);
nor U6003 (N_6003,N_2439,N_2455);
nor U6004 (N_6004,N_2851,N_1564);
nor U6005 (N_6005,N_901,N_64);
or U6006 (N_6006,N_470,N_3493);
or U6007 (N_6007,N_4574,N_855);
and U6008 (N_6008,N_682,N_1036);
nor U6009 (N_6009,N_1783,N_3091);
or U6010 (N_6010,N_3587,N_4090);
nor U6011 (N_6011,N_228,N_867);
nor U6012 (N_6012,N_2704,N_4309);
and U6013 (N_6013,N_1366,N_3400);
nor U6014 (N_6014,N_4053,N_2527);
nand U6015 (N_6015,N_2888,N_1355);
nand U6016 (N_6016,N_1631,N_515);
nand U6017 (N_6017,N_548,N_2360);
nand U6018 (N_6018,N_4247,N_4251);
nand U6019 (N_6019,N_546,N_4467);
or U6020 (N_6020,N_113,N_2151);
nor U6021 (N_6021,N_211,N_2720);
and U6022 (N_6022,N_2964,N_3043);
and U6023 (N_6023,N_2935,N_2617);
nand U6024 (N_6024,N_719,N_4110);
nand U6025 (N_6025,N_409,N_299);
nor U6026 (N_6026,N_4506,N_1378);
or U6027 (N_6027,N_3875,N_3014);
nand U6028 (N_6028,N_2592,N_4233);
nor U6029 (N_6029,N_203,N_4617);
and U6030 (N_6030,N_3469,N_1682);
nor U6031 (N_6031,N_4485,N_1978);
nor U6032 (N_6032,N_2417,N_4105);
and U6033 (N_6033,N_2980,N_433);
or U6034 (N_6034,N_1502,N_809);
nand U6035 (N_6035,N_3817,N_550);
or U6036 (N_6036,N_4037,N_46);
nand U6037 (N_6037,N_2869,N_1316);
or U6038 (N_6038,N_1119,N_4624);
and U6039 (N_6039,N_4520,N_3119);
nor U6040 (N_6040,N_3677,N_2027);
nand U6041 (N_6041,N_4282,N_4026);
and U6042 (N_6042,N_3153,N_2496);
nand U6043 (N_6043,N_3090,N_2166);
or U6044 (N_6044,N_2369,N_4493);
nand U6045 (N_6045,N_4492,N_2578);
or U6046 (N_6046,N_3021,N_2632);
nor U6047 (N_6047,N_1935,N_2652);
or U6048 (N_6048,N_77,N_2407);
nand U6049 (N_6049,N_2135,N_764);
and U6050 (N_6050,N_2397,N_1951);
nor U6051 (N_6051,N_654,N_2792);
nand U6052 (N_6052,N_2602,N_3736);
nor U6053 (N_6053,N_4996,N_1462);
xnor U6054 (N_6054,N_1826,N_3986);
and U6055 (N_6055,N_3409,N_547);
or U6056 (N_6056,N_738,N_3194);
nor U6057 (N_6057,N_2542,N_2);
or U6058 (N_6058,N_457,N_4335);
or U6059 (N_6059,N_3248,N_1528);
nand U6060 (N_6060,N_3134,N_3292);
nand U6061 (N_6061,N_4362,N_1950);
and U6062 (N_6062,N_4514,N_4342);
nor U6063 (N_6063,N_2422,N_2035);
or U6064 (N_6064,N_4077,N_4117);
nand U6065 (N_6065,N_3151,N_1813);
nand U6066 (N_6066,N_2902,N_4646);
nand U6067 (N_6067,N_2017,N_2716);
nor U6068 (N_6068,N_4400,N_3009);
nor U6069 (N_6069,N_1485,N_2209);
nor U6070 (N_6070,N_2461,N_3102);
nor U6071 (N_6071,N_1820,N_3589);
nand U6072 (N_6072,N_914,N_4672);
nor U6073 (N_6073,N_1911,N_419);
and U6074 (N_6074,N_711,N_4036);
nor U6075 (N_6075,N_3341,N_4890);
and U6076 (N_6076,N_2599,N_2173);
nand U6077 (N_6077,N_4385,N_2127);
nor U6078 (N_6078,N_973,N_2765);
and U6079 (N_6079,N_263,N_4712);
or U6080 (N_6080,N_3811,N_600);
nand U6081 (N_6081,N_1952,N_1612);
nand U6082 (N_6082,N_2933,N_2735);
nor U6083 (N_6083,N_640,N_890);
nor U6084 (N_6084,N_646,N_3471);
nor U6085 (N_6085,N_3934,N_4613);
nor U6086 (N_6086,N_4134,N_1971);
and U6087 (N_6087,N_2012,N_4175);
nor U6088 (N_6088,N_3204,N_1565);
and U6089 (N_6089,N_9,N_1017);
nand U6090 (N_6090,N_4425,N_4108);
or U6091 (N_6091,N_1498,N_3133);
nor U6092 (N_6092,N_3595,N_3251);
or U6093 (N_6093,N_2817,N_4937);
nand U6094 (N_6094,N_4903,N_94);
nor U6095 (N_6095,N_2050,N_4055);
or U6096 (N_6096,N_1118,N_3635);
nor U6097 (N_6097,N_4629,N_2476);
and U6098 (N_6098,N_2977,N_4478);
or U6099 (N_6099,N_1148,N_4358);
nand U6100 (N_6100,N_1974,N_1324);
or U6101 (N_6101,N_2841,N_50);
and U6102 (N_6102,N_3192,N_837);
nor U6103 (N_6103,N_4176,N_2609);
or U6104 (N_6104,N_2750,N_1634);
nor U6105 (N_6105,N_699,N_2630);
nor U6106 (N_6106,N_4263,N_2583);
or U6107 (N_6107,N_395,N_4656);
or U6108 (N_6108,N_892,N_2262);
or U6109 (N_6109,N_4586,N_749);
nand U6110 (N_6110,N_1696,N_2194);
nor U6111 (N_6111,N_3111,N_3129);
or U6112 (N_6112,N_3976,N_1143);
and U6113 (N_6113,N_4330,N_2368);
or U6114 (N_6114,N_4426,N_438);
nand U6115 (N_6115,N_2826,N_4085);
xor U6116 (N_6116,N_2299,N_1972);
and U6117 (N_6117,N_3142,N_2971);
and U6118 (N_6118,N_1867,N_3741);
or U6119 (N_6119,N_2109,N_2141);
and U6120 (N_6120,N_4967,N_2230);
nand U6121 (N_6121,N_1985,N_3700);
or U6122 (N_6122,N_4377,N_1833);
nand U6123 (N_6123,N_2424,N_368);
xnor U6124 (N_6124,N_2918,N_2728);
and U6125 (N_6125,N_2370,N_3674);
and U6126 (N_6126,N_2319,N_3394);
nor U6127 (N_6127,N_1836,N_2361);
and U6128 (N_6128,N_4466,N_2988);
nand U6129 (N_6129,N_4153,N_953);
and U6130 (N_6130,N_1827,N_3543);
and U6131 (N_6131,N_4332,N_4756);
nand U6132 (N_6132,N_2032,N_2145);
nor U6133 (N_6133,N_982,N_3239);
or U6134 (N_6134,N_1010,N_4746);
nor U6135 (N_6135,N_746,N_4191);
nor U6136 (N_6136,N_2040,N_1479);
nand U6137 (N_6137,N_623,N_3223);
nand U6138 (N_6138,N_870,N_2215);
and U6139 (N_6139,N_4004,N_2464);
nor U6140 (N_6140,N_231,N_247);
or U6141 (N_6141,N_3393,N_4346);
nand U6142 (N_6142,N_4928,N_1916);
and U6143 (N_6143,N_1213,N_2463);
nand U6144 (N_6144,N_4299,N_4052);
nor U6145 (N_6145,N_1165,N_2421);
nor U6146 (N_6146,N_2233,N_4082);
nand U6147 (N_6147,N_2732,N_1802);
or U6148 (N_6148,N_148,N_3540);
and U6149 (N_6149,N_4895,N_3294);
nor U6150 (N_6150,N_4578,N_1419);
and U6151 (N_6151,N_4811,N_881);
nand U6152 (N_6152,N_1763,N_3719);
or U6153 (N_6153,N_1389,N_2284);
and U6154 (N_6154,N_4677,N_4997);
nor U6155 (N_6155,N_3131,N_3822);
and U6156 (N_6156,N_4602,N_2330);
and U6157 (N_6157,N_2323,N_3003);
or U6158 (N_6158,N_969,N_4502);
nand U6159 (N_6159,N_3977,N_1842);
nand U6160 (N_6160,N_1429,N_2073);
nand U6161 (N_6161,N_2129,N_816);
and U6162 (N_6162,N_4568,N_525);
and U6163 (N_6163,N_4126,N_4003);
and U6164 (N_6164,N_1550,N_2579);
nand U6165 (N_6165,N_2695,N_3858);
nand U6166 (N_6166,N_3731,N_763);
nand U6167 (N_6167,N_3047,N_4583);
and U6168 (N_6168,N_3533,N_3066);
nand U6169 (N_6169,N_3384,N_342);
nand U6170 (N_6170,N_3692,N_1295);
nor U6171 (N_6171,N_1450,N_3335);
and U6172 (N_6172,N_1176,N_2250);
and U6173 (N_6173,N_164,N_4611);
and U6174 (N_6174,N_3790,N_4076);
or U6175 (N_6175,N_3442,N_2801);
nor U6176 (N_6176,N_3753,N_905);
nand U6177 (N_6177,N_4253,N_1464);
or U6178 (N_6178,N_1247,N_1835);
nor U6179 (N_6179,N_2248,N_1235);
xnor U6180 (N_6180,N_4658,N_2283);
and U6181 (N_6181,N_2837,N_3782);
or U6182 (N_6182,N_1325,N_3233);
nor U6183 (N_6183,N_1254,N_28);
or U6184 (N_6184,N_3925,N_1221);
nand U6185 (N_6185,N_4424,N_3966);
nor U6186 (N_6186,N_25,N_1979);
nand U6187 (N_6187,N_2636,N_3892);
nand U6188 (N_6188,N_3334,N_1305);
or U6189 (N_6189,N_4649,N_677);
nor U6190 (N_6190,N_4902,N_286);
and U6191 (N_6191,N_4727,N_959);
nor U6192 (N_6192,N_1444,N_3949);
xor U6193 (N_6193,N_2939,N_1649);
nand U6194 (N_6194,N_2390,N_4313);
and U6195 (N_6195,N_2673,N_4065);
or U6196 (N_6196,N_4546,N_3081);
or U6197 (N_6197,N_2782,N_4970);
or U6198 (N_6198,N_21,N_3593);
nor U6199 (N_6199,N_3582,N_961);
nor U6200 (N_6200,N_2635,N_1806);
nor U6201 (N_6201,N_4130,N_1605);
nor U6202 (N_6202,N_4074,N_2243);
nor U6203 (N_6203,N_1889,N_1541);
nor U6204 (N_6204,N_1515,N_394);
and U6205 (N_6205,N_4631,N_777);
or U6206 (N_6206,N_801,N_1070);
or U6207 (N_6207,N_1707,N_2539);
or U6208 (N_6208,N_2272,N_100);
or U6209 (N_6209,N_2934,N_3187);
and U6210 (N_6210,N_1430,N_980);
nand U6211 (N_6211,N_4375,N_3006);
nor U6212 (N_6212,N_3916,N_2076);
or U6213 (N_6213,N_4694,N_1173);
and U6214 (N_6214,N_3910,N_3290);
and U6215 (N_6215,N_3125,N_4918);
nor U6216 (N_6216,N_1503,N_4961);
or U6217 (N_6217,N_518,N_1785);
nor U6218 (N_6218,N_1997,N_2438);
and U6219 (N_6219,N_3283,N_3796);
nand U6220 (N_6220,N_829,N_358);
nor U6221 (N_6221,N_4148,N_4974);
nand U6222 (N_6222,N_908,N_1318);
nor U6223 (N_6223,N_979,N_863);
nor U6224 (N_6224,N_2408,N_4876);
nand U6225 (N_6225,N_4648,N_4304);
or U6226 (N_6226,N_645,N_2653);
nor U6227 (N_6227,N_986,N_1024);
nand U6228 (N_6228,N_2384,N_4344);
nand U6229 (N_6229,N_3205,N_3758);
nand U6230 (N_6230,N_2577,N_4598);
or U6231 (N_6231,N_4152,N_3098);
nor U6232 (N_6232,N_1418,N_1686);
nor U6233 (N_6233,N_572,N_1484);
xor U6234 (N_6234,N_2083,N_4985);
and U6235 (N_6235,N_3632,N_740);
and U6236 (N_6236,N_4660,N_1292);
and U6237 (N_6237,N_1995,N_1536);
nor U6238 (N_6238,N_752,N_4818);
and U6239 (N_6239,N_1167,N_1447);
nand U6240 (N_6240,N_3207,N_330);
or U6241 (N_6241,N_2214,N_1252);
nand U6242 (N_6242,N_487,N_1337);
and U6243 (N_6243,N_4990,N_2628);
nor U6244 (N_6244,N_1226,N_2832);
nor U6245 (N_6245,N_2182,N_31);
and U6246 (N_6246,N_388,N_236);
or U6247 (N_6247,N_2358,N_2400);
and U6248 (N_6248,N_1286,N_2976);
and U6249 (N_6249,N_3445,N_3642);
nand U6250 (N_6250,N_1234,N_3791);
nand U6251 (N_6251,N_1321,N_2931);
or U6252 (N_6252,N_2876,N_206);
or U6253 (N_6253,N_1772,N_4353);
or U6254 (N_6254,N_269,N_3770);
and U6255 (N_6255,N_1244,N_4925);
nand U6256 (N_6256,N_1947,N_1719);
and U6257 (N_6257,N_1905,N_2030);
nand U6258 (N_6258,N_4348,N_4462);
nor U6259 (N_6259,N_2183,N_4581);
nor U6260 (N_6260,N_4349,N_3395);
and U6261 (N_6261,N_352,N_3399);
nand U6262 (N_6262,N_1089,N_871);
or U6263 (N_6263,N_1658,N_4460);
nand U6264 (N_6264,N_1095,N_2947);
or U6265 (N_6265,N_3214,N_4905);
nand U6266 (N_6266,N_4652,N_2936);
or U6267 (N_6267,N_4901,N_4678);
and U6268 (N_6268,N_799,N_3628);
xnor U6269 (N_6269,N_3069,N_3466);
nand U6270 (N_6270,N_1635,N_4710);
nand U6271 (N_6271,N_2619,N_82);
and U6272 (N_6272,N_3701,N_3978);
nor U6273 (N_6273,N_2133,N_3638);
and U6274 (N_6274,N_4278,N_3333);
and U6275 (N_6275,N_2157,N_1372);
and U6276 (N_6276,N_4226,N_800);
and U6277 (N_6277,N_1302,N_1079);
and U6278 (N_6278,N_238,N_2836);
nor U6279 (N_6279,N_4416,N_3544);
nand U6280 (N_6280,N_4880,N_1086);
nand U6281 (N_6281,N_2756,N_3558);
or U6282 (N_6282,N_4547,N_4058);
nand U6283 (N_6283,N_3178,N_4636);
nand U6284 (N_6284,N_3697,N_431);
nand U6285 (N_6285,N_4942,N_673);
nand U6286 (N_6286,N_684,N_4041);
or U6287 (N_6287,N_225,N_3716);
nor U6288 (N_6288,N_2639,N_3985);
nand U6289 (N_6289,N_3843,N_3289);
and U6290 (N_6290,N_35,N_177);
nand U6291 (N_6291,N_423,N_3564);
nor U6292 (N_6292,N_1822,N_861);
and U6293 (N_6293,N_332,N_404);
nor U6294 (N_6294,N_2548,N_354);
or U6295 (N_6295,N_1516,N_3177);
nor U6296 (N_6296,N_17,N_339);
or U6297 (N_6297,N_4008,N_4167);
and U6298 (N_6298,N_1895,N_830);
and U6299 (N_6299,N_1021,N_3919);
nand U6300 (N_6300,N_143,N_4762);
nand U6301 (N_6301,N_167,N_3385);
and U6302 (N_6302,N_3457,N_343);
nand U6303 (N_6303,N_2167,N_65);
nor U6304 (N_6304,N_312,N_1182);
nand U6305 (N_6305,N_4798,N_1161);
nor U6306 (N_6306,N_1641,N_1630);
or U6307 (N_6307,N_3485,N_3276);
nand U6308 (N_6308,N_1796,N_3287);
and U6309 (N_6309,N_4522,N_906);
nor U6310 (N_6310,N_1620,N_1402);
nand U6311 (N_6311,N_4579,N_3046);
xor U6312 (N_6312,N_951,N_602);
nor U6313 (N_6313,N_2010,N_4719);
nor U6314 (N_6314,N_1425,N_473);
and U6315 (N_6315,N_2477,N_4667);
nor U6316 (N_6316,N_2431,N_3729);
nor U6317 (N_6317,N_4129,N_4410);
or U6318 (N_6318,N_4331,N_4206);
and U6319 (N_6319,N_4013,N_2593);
nor U6320 (N_6320,N_2882,N_1689);
and U6321 (N_6321,N_2164,N_3886);
nand U6322 (N_6322,N_1741,N_344);
nand U6323 (N_6323,N_3511,N_4376);
or U6324 (N_6324,N_1954,N_4443);
or U6325 (N_6325,N_4874,N_191);
and U6326 (N_6326,N_4327,N_2267);
or U6327 (N_6327,N_621,N_2219);
nor U6328 (N_6328,N_533,N_1016);
nand U6329 (N_6329,N_1023,N_2896);
nor U6330 (N_6330,N_3940,N_3019);
nand U6331 (N_6331,N_3110,N_3425);
and U6332 (N_6332,N_1336,N_474);
nor U6333 (N_6333,N_3744,N_224);
nand U6334 (N_6334,N_2752,N_4122);
or U6335 (N_6335,N_759,N_4651);
or U6336 (N_6336,N_3087,N_3982);
nor U6337 (N_6337,N_721,N_715);
and U6338 (N_6338,N_4551,N_2285);
and U6339 (N_6339,N_4312,N_4097);
and U6340 (N_6340,N_4752,N_3722);
and U6341 (N_6341,N_1142,N_2545);
and U6342 (N_6342,N_335,N_1706);
and U6343 (N_6343,N_2345,N_3644);
and U6344 (N_6344,N_946,N_39);
and U6345 (N_6345,N_1319,N_723);
or U6346 (N_6346,N_2916,N_2015);
nand U6347 (N_6347,N_4952,N_3303);
or U6348 (N_6348,N_4870,N_4944);
and U6349 (N_6349,N_3725,N_3837);
and U6350 (N_6350,N_1595,N_1903);
or U6351 (N_6351,N_3838,N_3901);
nor U6352 (N_6352,N_3042,N_1237);
or U6353 (N_6353,N_1123,N_2094);
nor U6354 (N_6354,N_2945,N_3267);
and U6355 (N_6355,N_1736,N_2645);
and U6356 (N_6356,N_3835,N_4027);
nor U6357 (N_6357,N_420,N_3057);
nand U6358 (N_6358,N_3612,N_920);
nand U6359 (N_6359,N_24,N_3296);
nor U6360 (N_6360,N_2433,N_2458);
nand U6361 (N_6361,N_2009,N_3998);
nand U6362 (N_6362,N_1973,N_3160);
xnor U6363 (N_6363,N_4697,N_1904);
nand U6364 (N_6364,N_4585,N_174);
nor U6365 (N_6365,N_309,N_1374);
nor U6366 (N_6366,N_823,N_2795);
nand U6367 (N_6367,N_1025,N_3756);
nor U6368 (N_6368,N_2092,N_1416);
or U6369 (N_6369,N_3787,N_4882);
nor U6370 (N_6370,N_814,N_4960);
and U6371 (N_6371,N_4260,N_1298);
or U6372 (N_6372,N_3447,N_940);
or U6373 (N_6373,N_1586,N_2937);
nand U6374 (N_6374,N_603,N_2047);
and U6375 (N_6375,N_2889,N_2702);
nand U6376 (N_6376,N_3723,N_4307);
and U6377 (N_6377,N_3519,N_4417);
and U6378 (N_6378,N_2474,N_2729);
or U6379 (N_6379,N_744,N_1673);
nand U6380 (N_6380,N_3439,N_87);
and U6381 (N_6381,N_4254,N_3598);
and U6382 (N_6382,N_1384,N_2824);
or U6383 (N_6383,N_2224,N_2858);
nand U6384 (N_6384,N_4827,N_2573);
and U6385 (N_6385,N_2906,N_1616);
nand U6386 (N_6386,N_3779,N_4038);
nand U6387 (N_6387,N_4695,N_3062);
or U6388 (N_6388,N_750,N_1597);
or U6389 (N_6389,N_2403,N_607);
nand U6390 (N_6390,N_4109,N_1224);
nand U6391 (N_6391,N_3606,N_1350);
nand U6392 (N_6392,N_4857,N_844);
nor U6393 (N_6393,N_1066,N_47);
or U6394 (N_6394,N_3273,N_3879);
or U6395 (N_6395,N_2852,N_1998);
nor U6396 (N_6396,N_3792,N_1261);
or U6397 (N_6397,N_1691,N_718);
nand U6398 (N_6398,N_2494,N_3711);
and U6399 (N_6399,N_4938,N_1255);
or U6400 (N_6400,N_3637,N_4713);
or U6401 (N_6401,N_3015,N_1776);
xor U6402 (N_6402,N_4615,N_2203);
nor U6403 (N_6403,N_1198,N_52);
nand U6404 (N_6404,N_3963,N_2504);
nand U6405 (N_6405,N_3622,N_2664);
and U6406 (N_6406,N_1081,N_1088);
nor U6407 (N_6407,N_2024,N_4028);
or U6408 (N_6408,N_2501,N_2910);
nand U6409 (N_6409,N_2983,N_2887);
and U6410 (N_6410,N_3424,N_1726);
nand U6411 (N_6411,N_2613,N_4782);
nand U6412 (N_6412,N_3703,N_1018);
nor U6413 (N_6413,N_2304,N_4927);
nor U6414 (N_6414,N_2950,N_434);
and U6415 (N_6415,N_4208,N_446);
and U6416 (N_6416,N_1598,N_3763);
nor U6417 (N_6417,N_4562,N_1109);
nand U6418 (N_6418,N_4111,N_3067);
or U6419 (N_6419,N_1188,N_2724);
nor U6420 (N_6420,N_1578,N_3475);
nand U6421 (N_6421,N_1054,N_2550);
nor U6422 (N_6422,N_1924,N_2519);
and U6423 (N_6423,N_4035,N_3412);
nand U6424 (N_6424,N_3512,N_3470);
or U6425 (N_6425,N_4216,N_3961);
and U6426 (N_6426,N_2879,N_4790);
nor U6427 (N_6427,N_1549,N_2061);
nor U6428 (N_6428,N_4680,N_2399);
nand U6429 (N_6429,N_4049,N_1263);
nor U6430 (N_6430,N_1133,N_1852);
nor U6431 (N_6431,N_1538,N_4354);
and U6432 (N_6432,N_2003,N_1961);
and U6433 (N_6433,N_4468,N_970);
or U6434 (N_6434,N_1746,N_3103);
and U6435 (N_6435,N_1797,N_212);
nor U6436 (N_6436,N_41,N_4161);
nor U6437 (N_6437,N_591,N_4359);
or U6438 (N_6438,N_3197,N_3076);
nor U6439 (N_6439,N_445,N_1601);
nor U6440 (N_6440,N_3909,N_3816);
and U6441 (N_6441,N_4213,N_4068);
and U6442 (N_6442,N_4361,N_824);
or U6443 (N_6443,N_2784,N_1968);
or U6444 (N_6444,N_4930,N_2502);
and U6445 (N_6445,N_374,N_2328);
xnor U6446 (N_6446,N_3023,N_2924);
and U6447 (N_6447,N_3171,N_4483);
nor U6448 (N_6448,N_2499,N_3144);
and U6449 (N_6449,N_598,N_3659);
nor U6450 (N_6450,N_2873,N_3324);
nor U6451 (N_6451,N_2863,N_4285);
nand U6452 (N_6452,N_2960,N_3836);
or U6453 (N_6453,N_327,N_1392);
nor U6454 (N_6454,N_480,N_2289);
nor U6455 (N_6455,N_3148,N_4171);
or U6456 (N_6456,N_3468,N_4030);
nor U6457 (N_6457,N_4820,N_1695);
nand U6458 (N_6458,N_935,N_2514);
nand U6459 (N_6459,N_4955,N_3402);
nor U6460 (N_6460,N_4591,N_2627);
nor U6461 (N_6461,N_1839,N_3083);
nand U6462 (N_6462,N_994,N_4907);
and U6463 (N_6463,N_4316,N_2608);
nor U6464 (N_6464,N_421,N_4800);
nand U6465 (N_6465,N_3894,N_243);
nor U6466 (N_6466,N_3968,N_2668);
and U6467 (N_6467,N_4034,N_3389);
and U6468 (N_6468,N_4499,N_2086);
or U6469 (N_6469,N_492,N_1500);
nand U6470 (N_6470,N_1694,N_3357);
nand U6471 (N_6471,N_2168,N_3472);
nand U6472 (N_6472,N_3231,N_2584);
nand U6473 (N_6473,N_4592,N_4116);
xor U6474 (N_6474,N_1881,N_4187);
nor U6475 (N_6475,N_485,N_3750);
or U6476 (N_6476,N_1388,N_665);
nor U6477 (N_6477,N_2965,N_662);
nor U6478 (N_6478,N_3338,N_3216);
nand U6479 (N_6479,N_2045,N_716);
nor U6480 (N_6480,N_1840,N_1831);
nor U6481 (N_6481,N_3227,N_1265);
or U6482 (N_6482,N_4265,N_1526);
nand U6483 (N_6483,N_3325,N_1376);
and U6484 (N_6484,N_1861,N_3948);
or U6485 (N_6485,N_3827,N_2791);
nor U6486 (N_6486,N_2091,N_2991);
and U6487 (N_6487,N_4872,N_1048);
or U6488 (N_6488,N_2650,N_1828);
or U6489 (N_6489,N_4744,N_3235);
or U6490 (N_6490,N_205,N_3318);
nand U6491 (N_6491,N_2423,N_356);
and U6492 (N_6492,N_4293,N_3051);
nor U6493 (N_6493,N_2270,N_106);
nor U6494 (N_6494,N_1207,N_4570);
and U6495 (N_6495,N_1158,N_1660);
or U6496 (N_6496,N_4268,N_3450);
nand U6497 (N_6497,N_3258,N_3680);
or U6498 (N_6498,N_4302,N_815);
nand U6499 (N_6499,N_2788,N_2556);
nand U6500 (N_6500,N_1507,N_2919);
or U6501 (N_6501,N_3801,N_2642);
or U6502 (N_6502,N_3504,N_3431);
nand U6503 (N_6503,N_4584,N_2590);
and U6504 (N_6504,N_4947,N_2085);
nand U6505 (N_6505,N_4157,N_3541);
and U6506 (N_6506,N_371,N_2530);
nand U6507 (N_6507,N_310,N_4098);
nor U6508 (N_6508,N_1659,N_1045);
and U6509 (N_6509,N_1011,N_786);
or U6510 (N_6510,N_315,N_428);
and U6511 (N_6511,N_2755,N_1534);
or U6512 (N_6512,N_2893,N_70);
or U6513 (N_6513,N_4177,N_3992);
nor U6514 (N_6514,N_3749,N_3531);
and U6515 (N_6515,N_2178,N_1918);
and U6516 (N_6516,N_3621,N_1728);
nand U6517 (N_6517,N_147,N_1766);
or U6518 (N_6518,N_3288,N_2878);
nor U6519 (N_6519,N_1514,N_1136);
nand U6520 (N_6520,N_1948,N_4112);
or U6521 (N_6521,N_3571,N_1780);
nor U6522 (N_6522,N_1356,N_2575);
and U6523 (N_6523,N_643,N_3956);
nor U6524 (N_6524,N_1931,N_1343);
and U6525 (N_6525,N_110,N_4626);
nand U6526 (N_6526,N_364,N_568);
nand U6527 (N_6527,N_1651,N_936);
nand U6528 (N_6528,N_706,N_111);
and U6529 (N_6529,N_3240,N_2667);
nand U6530 (N_6530,N_2392,N_874);
nand U6531 (N_6531,N_1679,N_3738);
nand U6532 (N_6532,N_3374,N_1181);
and U6533 (N_6533,N_4703,N_1775);
nand U6534 (N_6534,N_907,N_3527);
and U6535 (N_6535,N_3639,N_1781);
nor U6536 (N_6536,N_3958,N_3882);
nor U6537 (N_6537,N_3127,N_2535);
and U6538 (N_6538,N_2587,N_2589);
and U6539 (N_6539,N_3180,N_3130);
nor U6540 (N_6540,N_4609,N_1078);
or U6541 (N_6541,N_2090,N_4641);
nor U6542 (N_6542,N_1894,N_1771);
and U6543 (N_6543,N_3880,N_1209);
nand U6544 (N_6544,N_4449,N_3908);
nor U6545 (N_6545,N_3603,N_3201);
and U6546 (N_6546,N_2677,N_154);
or U6547 (N_6547,N_4005,N_555);
nor U6548 (N_6548,N_3002,N_412);
and U6549 (N_6549,N_1134,N_3971);
nor U6550 (N_6550,N_3663,N_2508);
nand U6551 (N_6551,N_1681,N_241);
or U6552 (N_6552,N_123,N_4988);
or U6553 (N_6553,N_491,N_4684);
or U6554 (N_6554,N_273,N_3830);
nor U6555 (N_6555,N_4463,N_862);
nor U6556 (N_6556,N_1730,N_2967);
nand U6557 (N_6557,N_681,N_2088);
and U6558 (N_6558,N_971,N_1264);
nand U6559 (N_6559,N_1600,N_4453);
or U6560 (N_6560,N_4557,N_2493);
nor U6561 (N_6561,N_3032,N_1653);
nor U6562 (N_6562,N_3215,N_3645);
or U6563 (N_6563,N_4718,N_3107);
nand U6564 (N_6564,N_2367,N_2574);
nor U6565 (N_6565,N_333,N_2880);
nor U6566 (N_6566,N_289,N_2547);
nand U6567 (N_6567,N_116,N_4464);
nor U6568 (N_6568,N_2311,N_3681);
nand U6569 (N_6569,N_943,N_376);
and U6570 (N_6570,N_524,N_2679);
or U6571 (N_6571,N_4465,N_2329);
nor U6572 (N_6572,N_1908,N_2195);
and U6573 (N_6573,N_1983,N_1632);
nand U6574 (N_6574,N_1692,N_4702);
and U6575 (N_6575,N_4473,N_3034);
and U6576 (N_6576,N_3369,N_1493);
and U6577 (N_6577,N_2159,N_1194);
nand U6578 (N_6578,N_532,N_4807);
or U6579 (N_6579,N_3917,N_544);
xor U6580 (N_6580,N_2341,N_1643);
and U6581 (N_6581,N_3135,N_4413);
nor U6582 (N_6582,N_2155,N_3182);
and U6583 (N_6583,N_2335,N_4919);
or U6584 (N_6584,N_3058,N_4145);
nor U6585 (N_6585,N_4565,N_2984);
nand U6586 (N_6586,N_4333,N_133);
nand U6587 (N_6587,N_1403,N_216);
nor U6588 (N_6588,N_4124,N_931);
nor U6589 (N_6589,N_1022,N_2347);
or U6590 (N_6590,N_1199,N_648);
or U6591 (N_6591,N_1646,N_2365);
and U6592 (N_6592,N_2383,N_4454);
nor U6593 (N_6593,N_770,N_659);
nand U6594 (N_6594,N_3249,N_2903);
and U6595 (N_6595,N_1609,N_2637);
nand U6596 (N_6596,N_20,N_576);
nand U6597 (N_6597,N_4162,N_3771);
or U6598 (N_6598,N_497,N_1218);
or U6599 (N_6599,N_2459,N_3422);
nor U6600 (N_6600,N_1853,N_2733);
nand U6601 (N_6601,N_2056,N_235);
and U6602 (N_6602,N_2014,N_2229);
nand U6603 (N_6603,N_2281,N_305);
or U6604 (N_6604,N_2952,N_477);
nor U6605 (N_6605,N_3115,N_4220);
and U6606 (N_6606,N_1117,N_2068);
nand U6607 (N_6607,N_2181,N_3804);
nand U6608 (N_6608,N_3183,N_2891);
nand U6609 (N_6609,N_2718,N_615);
nand U6610 (N_6610,N_4923,N_3039);
or U6611 (N_6611,N_84,N_2808);
or U6612 (N_6612,N_488,N_1294);
or U6613 (N_6613,N_921,N_425);
or U6614 (N_6614,N_1513,N_3257);
nand U6615 (N_6615,N_2366,N_894);
and U6616 (N_6616,N_771,N_1457);
and U6617 (N_6617,N_1395,N_4542);
or U6618 (N_6618,N_3675,N_2886);
nor U6619 (N_6619,N_611,N_3211);
nor U6620 (N_6620,N_4559,N_1488);
or U6621 (N_6621,N_3453,N_1189);
nand U6622 (N_6622,N_3281,N_3440);
nand U6623 (N_6623,N_1417,N_2420);
or U6624 (N_6624,N_4795,N_3928);
nor U6625 (N_6625,N_1460,N_1137);
nor U6626 (N_6626,N_1657,N_3557);
xor U6627 (N_6627,N_4054,N_2987);
nand U6628 (N_6628,N_3623,N_2962);
nand U6629 (N_6629,N_3253,N_1747);
nor U6630 (N_6630,N_4595,N_4326);
nor U6631 (N_6631,N_2371,N_1040);
nor U6632 (N_6632,N_1028,N_1477);
or U6633 (N_6633,N_3188,N_3092);
nor U6634 (N_6634,N_3579,N_4256);
nand U6635 (N_6635,N_954,N_2309);
or U6636 (N_6636,N_124,N_1693);
or U6637 (N_6637,N_2454,N_278);
nor U6638 (N_6638,N_1149,N_1574);
nand U6639 (N_6639,N_1584,N_3079);
nand U6640 (N_6640,N_3351,N_2220);
and U6641 (N_6641,N_4555,N_429);
nand U6642 (N_6642,N_2713,N_414);
xnor U6643 (N_6643,N_2820,N_3195);
nor U6644 (N_6644,N_1745,N_3482);
or U6645 (N_6645,N_4888,N_1876);
nand U6646 (N_6646,N_2175,N_4380);
nand U6647 (N_6647,N_3332,N_2419);
and U6648 (N_6648,N_2044,N_4849);
nand U6649 (N_6649,N_1655,N_2137);
xnor U6650 (N_6650,N_1915,N_1340);
nand U6651 (N_6651,N_4833,N_3927);
nand U6652 (N_6652,N_4939,N_128);
or U6653 (N_6653,N_2890,N_2082);
and U6654 (N_6654,N_2161,N_1486);
and U6655 (N_6655,N_3001,N_56);
and U6656 (N_6656,N_1672,N_298);
nor U6657 (N_6657,N_1077,N_4823);
or U6658 (N_6658,N_1858,N_2261);
nor U6659 (N_6659,N_2096,N_2072);
nand U6660 (N_6660,N_4215,N_4441);
nand U6661 (N_6661,N_1243,N_2110);
and U6662 (N_6662,N_2255,N_4269);
or U6663 (N_6663,N_2957,N_4470);
nor U6664 (N_6664,N_288,N_2810);
nor U6665 (N_6665,N_1718,N_4513);
nor U6666 (N_6666,N_2475,N_2687);
or U6667 (N_6667,N_590,N_753);
nor U6668 (N_6668,N_2543,N_991);
nand U6669 (N_6669,N_4474,N_67);
or U6670 (N_6670,N_1399,N_3685);
or U6671 (N_6671,N_2352,N_1580);
nor U6672 (N_6672,N_3435,N_927);
and U6673 (N_6673,N_249,N_2468);
or U6674 (N_6674,N_1277,N_1229);
or U6675 (N_6675,N_2860,N_2039);
nand U6676 (N_6676,N_4103,N_2849);
nor U6677 (N_6677,N_724,N_3611);
nor U6678 (N_6678,N_1765,N_2355);
and U6679 (N_6679,N_392,N_704);
nor U6680 (N_6680,N_899,N_1752);
and U6681 (N_6681,N_620,N_3252);
and U6682 (N_6682,N_4730,N_4524);
nand U6683 (N_6683,N_260,N_2802);
nand U6684 (N_6684,N_3096,N_517);
nor U6685 (N_6685,N_3704,N_313);
nor U6686 (N_6686,N_1671,N_4423);
or U6687 (N_6687,N_2512,N_4539);
nand U6688 (N_6688,N_2059,N_3071);
nor U6689 (N_6689,N_4843,N_1280);
nor U6690 (N_6690,N_2197,N_2307);
nor U6691 (N_6691,N_2529,N_2325);
nor U6692 (N_6692,N_1091,N_1320);
nand U6693 (N_6693,N_2618,N_2763);
nor U6694 (N_6694,N_2648,N_4987);
and U6695 (N_6695,N_2205,N_2266);
nand U6696 (N_6696,N_2785,N_1992);
and U6697 (N_6697,N_2406,N_188);
and U6698 (N_6698,N_3570,N_2701);
or U6699 (N_6699,N_944,N_75);
or U6700 (N_6700,N_957,N_198);
nor U6701 (N_6701,N_3618,N_3056);
and U6702 (N_6702,N_3415,N_2949);
or U6703 (N_6703,N_1900,N_4190);
or U6704 (N_6704,N_3476,N_2557);
or U6705 (N_6705,N_187,N_1197);
or U6706 (N_6706,N_4707,N_2580);
or U6707 (N_6707,N_237,N_4564);
and U6708 (N_6708,N_4829,N_1569);
nand U6709 (N_6709,N_4959,N_4999);
or U6710 (N_6710,N_2238,N_1413);
and U6711 (N_6711,N_3117,N_4056);
and U6712 (N_6712,N_4337,N_3118);
or U6713 (N_6713,N_4182,N_3549);
nand U6714 (N_6714,N_3656,N_2171);
nand U6715 (N_6715,N_2128,N_4430);
or U6716 (N_6716,N_2412,N_4682);
nor U6717 (N_6717,N_4534,N_628);
nand U6718 (N_6718,N_2237,N_2830);
nor U6719 (N_6719,N_2928,N_1466);
and U6720 (N_6720,N_996,N_2631);
and U6721 (N_6721,N_1678,N_4501);
or U6722 (N_6722,N_1299,N_4630);
xor U6723 (N_6723,N_3181,N_4193);
nor U6724 (N_6724,N_3347,N_4159);
nand U6725 (N_6725,N_3826,N_359);
or U6726 (N_6726,N_3856,N_1029);
nor U6727 (N_6727,N_1581,N_1769);
nand U6728 (N_6728,N_3833,N_1884);
nor U6729 (N_6729,N_4582,N_1073);
nand U6730 (N_6730,N_3586,N_4412);
nor U6731 (N_6731,N_1570,N_4238);
and U6732 (N_6732,N_4982,N_4989);
nor U6733 (N_6733,N_2437,N_1755);
xnor U6734 (N_6734,N_2908,N_271);
or U6735 (N_6735,N_1083,N_1687);
nor U6736 (N_6736,N_1556,N_2080);
or U6737 (N_6737,N_4294,N_1591);
nand U6738 (N_6738,N_2914,N_3392);
nand U6739 (N_6739,N_3754,N_1272);
nor U6740 (N_6740,N_754,N_4434);
xnor U6741 (N_6741,N_1454,N_2948);
and U6742 (N_6742,N_4775,N_2179);
and U6743 (N_6743,N_331,N_1085);
nand U6744 (N_6744,N_2353,N_2020);
or U6745 (N_6745,N_1723,N_4701);
and U6746 (N_6746,N_3818,N_413);
nor U6747 (N_6747,N_769,N_1332);
or U6748 (N_6748,N_4904,N_3673);
nand U6749 (N_6749,N_2812,N_3095);
nor U6750 (N_6750,N_1559,N_112);
or U6751 (N_6751,N_2862,N_3059);
or U6752 (N_6752,N_2633,N_367);
or U6753 (N_6753,N_1451,N_1787);
or U6754 (N_6754,N_4900,N_1967);
or U6755 (N_6755,N_3797,N_71);
nand U6756 (N_6756,N_3534,N_119);
xnor U6757 (N_6757,N_1043,N_1156);
or U6758 (N_6758,N_3698,N_3139);
or U6759 (N_6759,N_2460,N_3049);
and U6760 (N_6760,N_2380,N_4688);
or U6761 (N_6761,N_166,N_157);
nor U6762 (N_6762,N_631,N_3765);
and U6763 (N_6763,N_1582,N_454);
nand U6764 (N_6764,N_3165,N_3013);
nor U6765 (N_6765,N_1561,N_3717);
or U6766 (N_6766,N_126,N_2572);
and U6767 (N_6767,N_55,N_3212);
or U6768 (N_6768,N_4698,N_3884);
nand U6769 (N_6769,N_2789,N_1103);
nand U6770 (N_6770,N_884,N_4386);
nand U6771 (N_6771,N_466,N_2805);
nor U6772 (N_6772,N_4720,N_44);
and U6773 (N_6773,N_4822,N_3241);
and U6774 (N_6774,N_1098,N_3672);
or U6775 (N_6775,N_4411,N_599);
nand U6776 (N_6776,N_873,N_1638);
nor U6777 (N_6777,N_4291,N_1735);
nor U6778 (N_6778,N_571,N_2932);
or U6779 (N_6779,N_501,N_2955);
nor U6780 (N_6780,N_4841,N_1274);
or U6781 (N_6781,N_3449,N_3007);
or U6782 (N_6782,N_1067,N_1379);
or U6783 (N_6783,N_2620,N_2404);
and U6784 (N_6784,N_4039,N_3314);
xnor U6785 (N_6785,N_1518,N_785);
or U6786 (N_6786,N_3855,N_1958);
nand U6787 (N_6787,N_925,N_1282);
and U6788 (N_6788,N_4072,N_3464);
nor U6789 (N_6789,N_4497,N_441);
nor U6790 (N_6790,N_4835,N_4450);
nor U6791 (N_6791,N_4781,N_3404);
and U6792 (N_6792,N_1327,N_3368);
nor U6793 (N_6793,N_1846,N_3694);
and U6794 (N_6794,N_2444,N_1359);
and U6795 (N_6795,N_453,N_2306);
or U6796 (N_6796,N_1970,N_3077);
xnor U6797 (N_6797,N_2232,N_1107);
nor U6798 (N_6798,N_989,N_2069);
and U6799 (N_6799,N_4368,N_962);
nor U6800 (N_6800,N_251,N_1739);
nand U6801 (N_6801,N_15,N_3885);
nor U6802 (N_6802,N_3229,N_4543);
or U6803 (N_6803,N_2571,N_2385);
nor U6804 (N_6804,N_1857,N_1977);
nand U6805 (N_6805,N_4750,N_1964);
nor U6806 (N_6806,N_4387,N_1102);
nand U6807 (N_6807,N_2273,N_72);
or U6808 (N_6808,N_1754,N_1699);
nand U6809 (N_6809,N_4240,N_4297);
nand U6810 (N_6810,N_4427,N_3752);
and U6811 (N_6811,N_4711,N_4517);
nand U6812 (N_6812,N_2057,N_838);
nand U6813 (N_6813,N_270,N_1543);
nor U6814 (N_6814,N_3678,N_2656);
or U6815 (N_6815,N_3259,N_1391);
nor U6816 (N_6816,N_242,N_373);
or U6817 (N_6817,N_2975,N_3596);
nor U6818 (N_6818,N_3068,N_3864);
or U6819 (N_6819,N_1253,N_4842);
and U6820 (N_6820,N_2228,N_2721);
or U6821 (N_6821,N_1124,N_3893);
nand U6822 (N_6822,N_522,N_411);
nand U6823 (N_6823,N_3423,N_4864);
and U6824 (N_6824,N_2470,N_3994);
and U6825 (N_6825,N_1212,N_1532);
and U6826 (N_6826,N_1721,N_3626);
nor U6827 (N_6827,N_353,N_4079);
nor U6828 (N_6828,N_656,N_159);
nand U6829 (N_6829,N_3881,N_2564);
nor U6830 (N_6830,N_349,N_215);
nor U6831 (N_6831,N_2877,N_650);
nor U6832 (N_6832,N_3345,N_2938);
nor U6833 (N_6833,N_4778,N_2418);
or U6834 (N_6834,N_1669,N_2803);
or U6835 (N_6835,N_1860,N_4700);
or U6836 (N_6836,N_4024,N_1732);
nor U6837 (N_6837,N_4729,N_2621);
or U6838 (N_6838,N_1344,N_4894);
nor U6839 (N_6839,N_185,N_2172);
and U6840 (N_6840,N_883,N_214);
nand U6841 (N_6841,N_1962,N_4014);
nor U6842 (N_6842,N_636,N_2696);
nor U6843 (N_6843,N_1888,N_502);
nand U6844 (N_6844,N_762,N_402);
and U6845 (N_6845,N_766,N_4933);
and U6846 (N_6846,N_2597,N_1383);
nor U6847 (N_6847,N_1875,N_86);
and U6848 (N_6848,N_1269,N_4588);
or U6849 (N_6849,N_4064,N_1311);
or U6850 (N_6850,N_1960,N_2116);
and U6851 (N_6851,N_1652,N_1546);
and U6852 (N_6852,N_2089,N_170);
and U6853 (N_6853,N_1205,N_2441);
nor U6854 (N_6854,N_3832,N_4367);
and U6855 (N_6855,N_3086,N_703);
or U6856 (N_6856,N_4403,N_3647);
or U6857 (N_6857,N_3506,N_92);
nor U6858 (N_6858,N_2119,N_661);
nand U6859 (N_6859,N_3403,N_4753);
or U6860 (N_6860,N_543,N_939);
nor U6861 (N_6861,N_317,N_34);
nor U6862 (N_6862,N_865,N_836);
or U6863 (N_6863,N_788,N_4797);
nor U6864 (N_6864,N_3513,N_653);
nand U6865 (N_6865,N_614,N_1751);
nand U6866 (N_6866,N_3346,N_4755);
or U6867 (N_6867,N_4429,N_4889);
nor U6868 (N_6868,N_558,N_3846);
nand U6869 (N_6869,N_4115,N_1420);
and U6870 (N_6870,N_281,N_4891);
or U6871 (N_6871,N_4668,N_449);
nor U6872 (N_6872,N_2804,N_321);
nand U6873 (N_6873,N_435,N_3784);
nand U6874 (N_6874,N_363,N_2954);
nand U6875 (N_6875,N_4769,N_1267);
or U6876 (N_6876,N_4510,N_4913);
or U6877 (N_6877,N_3027,N_4149);
or U6878 (N_6878,N_2402,N_4194);
or U6879 (N_6879,N_2615,N_89);
nand U6880 (N_6880,N_619,N_302);
xor U6881 (N_6881,N_2681,N_1742);
or U6882 (N_6882,N_802,N_4958);
and U6883 (N_6883,N_4384,N_345);
nor U6884 (N_6884,N_789,N_2719);
or U6885 (N_6885,N_4317,N_2007);
or U6886 (N_6886,N_3004,N_3157);
nand U6887 (N_6887,N_3286,N_1242);
nand U6888 (N_6888,N_4867,N_1065);
nor U6889 (N_6889,N_4787,N_2435);
or U6890 (N_6890,N_4855,N_4435);
nor U6891 (N_6891,N_1041,N_3360);
or U6892 (N_6892,N_1700,N_4840);
nand U6893 (N_6893,N_3799,N_3430);
and U6894 (N_6894,N_301,N_1496);
or U6895 (N_6895,N_2923,N_4708);
and U6896 (N_6896,N_4186,N_183);
and U6897 (N_6897,N_3167,N_4308);
xor U6898 (N_6898,N_3649,N_78);
nor U6899 (N_6899,N_220,N_3169);
or U6900 (N_6900,N_4521,N_2378);
and U6901 (N_6901,N_2066,N_1517);
and U6902 (N_6902,N_40,N_4495);
and U6903 (N_6903,N_1944,N_1233);
nand U6904 (N_6904,N_142,N_4786);
nand U6905 (N_6905,N_3820,N_567);
nor U6906 (N_6906,N_4714,N_461);
or U6907 (N_6907,N_1690,N_401);
nand U6908 (N_6908,N_4310,N_3515);
nor U6909 (N_6909,N_1214,N_2006);
nor U6910 (N_6910,N_1902,N_717);
or U6911 (N_6911,N_3556,N_929);
or U6912 (N_6912,N_3380,N_1837);
nor U6913 (N_6913,N_276,N_4610);
nand U6914 (N_6914,N_1841,N_3567);
or U6915 (N_6915,N_1722,N_90);
nand U6916 (N_6916,N_1435,N_1847);
nor U6917 (N_6917,N_1683,N_4968);
nor U6918 (N_6918,N_609,N_2675);
and U6919 (N_6919,N_4806,N_233);
or U6920 (N_6920,N_1115,N_2317);
nand U6921 (N_6921,N_3427,N_3954);
and U6922 (N_6922,N_632,N_3691);
nand U6923 (N_6923,N_3168,N_2517);
and U6924 (N_6924,N_4422,N_3921);
xor U6925 (N_6925,N_1555,N_4407);
xnor U6926 (N_6926,N_2142,N_4080);
nor U6927 (N_6927,N_4774,N_4489);
nor U6928 (N_6928,N_2213,N_974);
and U6929 (N_6929,N_4884,N_1492);
nor U6930 (N_6930,N_4969,N_4217);
nand U6931 (N_6931,N_2894,N_915);
and U6932 (N_6932,N_3146,N_2839);
nor U6933 (N_6933,N_2537,N_3124);
or U6934 (N_6934,N_737,N_1030);
and U6935 (N_6935,N_3323,N_639);
nor U6936 (N_6936,N_2769,N_3104);
nor U6937 (N_6937,N_146,N_1596);
nor U6938 (N_6938,N_2699,N_1476);
or U6939 (N_6939,N_4488,N_4793);
or U6940 (N_6940,N_1489,N_4600);
nor U6941 (N_6941,N_1364,N_3874);
nand U6942 (N_6942,N_582,N_4922);
nor U6943 (N_6943,N_1984,N_584);
nand U6944 (N_6944,N_322,N_2655);
and U6945 (N_6945,N_1287,N_3669);
nand U6946 (N_6946,N_3800,N_2787);
nor U6947 (N_6947,N_2823,N_4084);
nor U6948 (N_6948,N_783,N_1333);
or U6949 (N_6949,N_2064,N_822);
nand U6950 (N_6950,N_4280,N_26);
or U6951 (N_6951,N_3671,N_3600);
nand U6952 (N_6952,N_3988,N_3220);
nand U6953 (N_6953,N_3777,N_2301);
nand U6954 (N_6954,N_731,N_3905);
or U6955 (N_6955,N_4654,N_3861);
nand U6956 (N_6956,N_4650,N_3304);
nor U6957 (N_6957,N_10,N_2705);
or U6958 (N_6958,N_163,N_1225);
nor U6959 (N_6959,N_4723,N_3951);
nand U6960 (N_6960,N_540,N_1448);
or U6961 (N_6961,N_4142,N_805);
or U6962 (N_6962,N_3550,N_4315);
nor U6963 (N_6963,N_3317,N_2995);
nor U6964 (N_6964,N_3581,N_3679);
nand U6965 (N_6965,N_651,N_3278);
and U6966 (N_6966,N_2509,N_1848);
nand U6967 (N_6967,N_1153,N_3530);
nand U6968 (N_6968,N_3887,N_4587);
nor U6969 (N_6969,N_2484,N_3232);
nand U6970 (N_6970,N_3441,N_1184);
and U6971 (N_6971,N_375,N_3696);
or U6972 (N_6972,N_4320,N_2021);
nor U6973 (N_6973,N_2553,N_3261);
nor U6974 (N_6974,N_2265,N_2364);
and U6975 (N_6975,N_3867,N_391);
or U6976 (N_6976,N_1328,N_2990);
or U6977 (N_6977,N_4094,N_4140);
nand U6978 (N_6978,N_3316,N_3218);
or U6979 (N_6979,N_857,N_1390);
and U6980 (N_6980,N_2777,N_535);
or U6981 (N_6981,N_101,N_3342);
or U6982 (N_6982,N_573,N_4029);
nor U6983 (N_6983,N_184,N_3497);
nor U6984 (N_6984,N_4549,N_4784);
nor U6985 (N_6985,N_4395,N_91);
and U6986 (N_6986,N_4946,N_1789);
nand U6987 (N_6987,N_3272,N_1351);
or U6988 (N_6988,N_2280,N_3560);
nand U6989 (N_6989,N_2567,N_2485);
and U6990 (N_6990,N_2104,N_511);
nor U6991 (N_6991,N_1639,N_2697);
and U6992 (N_6992,N_4061,N_758);
nor U6993 (N_6993,N_3724,N_2913);
or U6994 (N_6994,N_917,N_137);
nor U6995 (N_6995,N_88,N_956);
nor U6996 (N_6996,N_4511,N_2174);
or U6997 (N_6997,N_1262,N_23);
and U6998 (N_6998,N_853,N_3312);
and U6999 (N_6999,N_3735,N_4794);
and U7000 (N_7000,N_1289,N_3122);
nand U7001 (N_7001,N_1709,N_1122);
nor U7002 (N_7002,N_1322,N_1007);
nor U7003 (N_7003,N_1174,N_2744);
nand U7004 (N_7004,N_4199,N_49);
nand U7005 (N_7005,N_3720,N_2268);
or U7006 (N_7006,N_2698,N_4173);
nor U7007 (N_7007,N_4172,N_4743);
or U7008 (N_7008,N_1338,N_2031);
or U7009 (N_7009,N_3328,N_3594);
nand U7010 (N_7010,N_1819,N_4716);
nor U7011 (N_7011,N_4202,N_1076);
nor U7012 (N_7012,N_4095,N_1285);
nand U7013 (N_7013,N_2715,N_245);
and U7014 (N_7014,N_3914,N_3584);
or U7015 (N_7015,N_1760,N_3768);
nor U7016 (N_7016,N_3851,N_4653);
or U7017 (N_7017,N_1129,N_4683);
or U7018 (N_7018,N_380,N_1917);
nand U7019 (N_7019,N_4127,N_1990);
xnor U7020 (N_7020,N_329,N_3479);
or U7021 (N_7021,N_3942,N_1064);
and U7022 (N_7022,N_4392,N_1887);
nand U7023 (N_7023,N_2660,N_2764);
or U7024 (N_7024,N_1625,N_1431);
and U7025 (N_7025,N_257,N_430);
or U7026 (N_7026,N_3532,N_4120);
nand U7027 (N_7027,N_3922,N_898);
nand U7028 (N_7028,N_2693,N_3005);
nand U7029 (N_7029,N_160,N_1415);
nand U7030 (N_7030,N_4518,N_3895);
nand U7031 (N_7031,N_3018,N_793);
nor U7032 (N_7032,N_1306,N_340);
and U7033 (N_7033,N_745,N_1834);
nor U7034 (N_7034,N_189,N_4704);
and U7035 (N_7035,N_3054,N_2124);
and U7036 (N_7036,N_3337,N_207);
nor U7037 (N_7037,N_1929,N_4290);
or U7038 (N_7038,N_2467,N_2269);
nor U7039 (N_7039,N_1801,N_2103);
nor U7040 (N_7040,N_4243,N_1061);
nand U7041 (N_7041,N_2416,N_3783);
nand U7042 (N_7042,N_1044,N_938);
and U7043 (N_7043,N_1717,N_3813);
or U7044 (N_7044,N_295,N_2308);
nor U7045 (N_7045,N_0,N_3658);
or U7046 (N_7046,N_674,N_267);
and U7047 (N_7047,N_3488,N_528);
or U7048 (N_7048,N_3112,N_2221);
nor U7049 (N_7049,N_2190,N_4866);
and U7050 (N_7050,N_102,N_1982);
nor U7051 (N_7051,N_115,N_1611);
and U7052 (N_7052,N_1854,N_348);
nor U7053 (N_7053,N_334,N_472);
or U7054 (N_7054,N_3149,N_4777);
nand U7055 (N_7055,N_647,N_2187);
nand U7056 (N_7056,N_254,N_4770);
nor U7057 (N_7057,N_2770,N_4196);
nor U7058 (N_7058,N_612,N_3481);
and U7059 (N_7059,N_597,N_3981);
or U7060 (N_7060,N_319,N_1814);
and U7061 (N_7061,N_3474,N_2462);
nand U7062 (N_7062,N_1404,N_197);
or U7063 (N_7063,N_370,N_2258);
or U7064 (N_7064,N_150,N_3708);
and U7065 (N_7065,N_1341,N_4505);
nor U7066 (N_7066,N_162,N_2242);
and U7067 (N_7067,N_1284,N_3072);
nor U7068 (N_7068,N_1525,N_2339);
nand U7069 (N_7069,N_4619,N_2025);
and U7070 (N_7070,N_1394,N_3284);
nor U7071 (N_7071,N_2930,N_4081);
nand U7072 (N_7072,N_3250,N_3126);
nor U7073 (N_7073,N_3329,N_4446);
nor U7074 (N_7074,N_1120,N_1981);
and U7075 (N_7075,N_2794,N_680);
or U7076 (N_7076,N_4438,N_3454);
nor U7077 (N_7077,N_3386,N_2170);
nand U7078 (N_7078,N_1567,N_3601);
nor U7079 (N_7079,N_725,N_4270);
nand U7080 (N_7080,N_4195,N_2624);
nand U7081 (N_7081,N_3955,N_1697);
nand U7082 (N_7082,N_2445,N_4607);
nand U7083 (N_7083,N_3561,N_1909);
nor U7084 (N_7084,N_3200,N_3238);
and U7085 (N_7085,N_742,N_3902);
and U7086 (N_7086,N_1799,N_1607);
and U7087 (N_7087,N_2314,N_3458);
or U7088 (N_7088,N_2662,N_1504);
nand U7089 (N_7089,N_1382,N_2132);
and U7090 (N_7090,N_1868,N_4739);
nand U7091 (N_7091,N_3937,N_4281);
or U7092 (N_7092,N_3444,N_3991);
nor U7093 (N_7093,N_2070,N_3);
xnor U7094 (N_7094,N_3834,N_1544);
nand U7095 (N_7095,N_579,N_4869);
nand U7096 (N_7096,N_3173,N_4879);
nand U7097 (N_7097,N_1976,N_4536);
or U7098 (N_7098,N_3208,N_1572);
nand U7099 (N_7099,N_3712,N_2333);
and U7100 (N_7100,N_447,N_4532);
or U7101 (N_7101,N_4608,N_4635);
nand U7102 (N_7102,N_1585,N_3769);
or U7103 (N_7103,N_3776,N_464);
nand U7104 (N_7104,N_4073,N_4618);
nor U7105 (N_7105,N_4868,N_1397);
or U7106 (N_7106,N_3209,N_1927);
or U7107 (N_7107,N_2746,N_4060);
or U7108 (N_7108,N_2883,N_1989);
nand U7109 (N_7109,N_1331,N_2425);
nand U7110 (N_7110,N_2071,N_3266);
or U7111 (N_7111,N_4821,N_4659);
nor U7112 (N_7112,N_7,N_841);
or U7113 (N_7113,N_1986,N_107);
and U7114 (N_7114,N_2176,N_32);
and U7115 (N_7115,N_671,N_1001);
and U7116 (N_7116,N_542,N_4851);
and U7117 (N_7117,N_4812,N_877);
and U7118 (N_7118,N_3518,N_1774);
nand U7119 (N_7119,N_3228,N_897);
nor U7120 (N_7120,N_2676,N_4597);
nand U7121 (N_7121,N_1441,N_1135);
nor U7122 (N_7122,N_1936,N_1443);
and U7123 (N_7123,N_1956,N_1250);
or U7124 (N_7124,N_2739,N_398);
nor U7125 (N_7125,N_4953,N_1957);
or U7126 (N_7126,N_3845,N_2489);
and U7127 (N_7127,N_1185,N_3331);
or U7128 (N_7128,N_4252,N_860);
or U7129 (N_7129,N_3164,N_835);
nor U7130 (N_7130,N_4594,N_3633);
nand U7131 (N_7131,N_2576,N_1191);
nand U7132 (N_7132,N_4573,N_3841);
nor U7133 (N_7133,N_3495,N_4691);
and U7134 (N_7134,N_2471,N_553);
nand U7135 (N_7135,N_442,N_4388);
and U7136 (N_7136,N_1724,N_4912);
nand U7137 (N_7137,N_4321,N_1542);
xnor U7138 (N_7138,N_4709,N_469);
nor U7139 (N_7139,N_3401,N_3465);
nand U7140 (N_7140,N_1926,N_495);
nand U7141 (N_7141,N_637,N_4276);
nor U7142 (N_7142,N_2997,N_1988);
nor U7143 (N_7143,N_4244,N_2324);
or U7144 (N_7144,N_4773,N_221);
xnor U7145 (N_7145,N_2029,N_4311);
and U7146 (N_7146,N_248,N_3150);
nor U7147 (N_7147,N_1803,N_3542);
nor U7148 (N_7148,N_4934,N_4101);
and U7149 (N_7149,N_1308,N_1768);
or U7150 (N_7150,N_3336,N_202);
or U7151 (N_7151,N_701,N_1408);
or U7152 (N_7152,N_2210,N_320);
and U7153 (N_7153,N_3213,N_4306);
nor U7154 (N_7154,N_3147,N_1560);
nor U7155 (N_7155,N_2150,N_3975);
nand U7156 (N_7156,N_3489,N_4845);
or U7157 (N_7157,N_1139,N_3295);
and U7158 (N_7158,N_4686,N_4725);
nor U7159 (N_7159,N_1554,N_3352);
or U7160 (N_7160,N_3436,N_1547);
and U7161 (N_7161,N_2643,N_4861);
nor U7162 (N_7162,N_990,N_1910);
or U7163 (N_7163,N_4092,N_69);
and U7164 (N_7164,N_554,N_1830);
or U7165 (N_7165,N_3210,N_193);
nand U7166 (N_7166,N_1922,N_2773);
or U7167 (N_7167,N_3640,N_2505);
or U7168 (N_7168,N_1049,N_43);
nand U7169 (N_7169,N_1314,N_1421);
and U7170 (N_7170,N_1996,N_3999);
nand U7171 (N_7171,N_792,N_1131);
and U7172 (N_7172,N_933,N_4839);
nor U7173 (N_7173,N_2286,N_38);
or U7174 (N_7174,N_679,N_1893);
nand U7175 (N_7175,N_1125,N_1748);
or U7176 (N_7176,N_2426,N_2743);
xor U7177 (N_7177,N_4087,N_622);
nand U7178 (N_7178,N_190,N_3789);
nor U7179 (N_7179,N_1170,N_2796);
nor U7180 (N_7180,N_1288,N_3805);
nor U7181 (N_7181,N_4765,N_79);
nor U7182 (N_7182,N_2436,N_2511);
nand U7183 (N_7183,N_1278,N_4603);
and U7184 (N_7184,N_3503,N_4527);
or U7185 (N_7185,N_325,N_839);
nand U7186 (N_7186,N_4078,N_427);
and U7187 (N_7187,N_3340,N_3196);
nor U7188 (N_7188,N_630,N_2440);
nand U7189 (N_7189,N_3175,N_3945);
nor U7190 (N_7190,N_2067,N_3361);
nand U7191 (N_7191,N_2497,N_3829);
nor U7192 (N_7192,N_2479,N_4637);
and U7193 (N_7193,N_2940,N_2899);
nand U7194 (N_7194,N_4910,N_4476);
or U7195 (N_7195,N_2709,N_171);
nand U7196 (N_7196,N_2108,N_1249);
and U7197 (N_7197,N_541,N_1811);
or U7198 (N_7198,N_3417,N_2956);
or U7199 (N_7199,N_2507,N_1899);
or U7200 (N_7200,N_99,N_2081);
nand U7201 (N_7201,N_2596,N_4994);
or U7202 (N_7202,N_4883,N_4789);
nor U7203 (N_7203,N_1138,N_2241);
or U7204 (N_7204,N_1937,N_2665);
and U7205 (N_7205,N_2188,N_3451);
and U7206 (N_7206,N_3913,N_2259);
or U7207 (N_7207,N_3364,N_2600);
nor U7208 (N_7208,N_1562,N_843);
nor U7209 (N_7209,N_1275,N_274);
and U7210 (N_7210,N_121,N_3138);
nor U7211 (N_7211,N_2842,N_4950);
nand U7212 (N_7212,N_3539,N_798);
and U7213 (N_7213,N_2087,N_1013);
or U7214 (N_7214,N_2414,N_3931);
nor U7215 (N_7215,N_808,N_3755);
nand U7216 (N_7216,N_1004,N_3322);
and U7217 (N_7217,N_887,N_4245);
or U7218 (N_7218,N_4914,N_3842);
nor U7219 (N_7219,N_3524,N_3462);
nand U7220 (N_7220,N_213,N_2217);
nor U7221 (N_7221,N_2806,N_3718);
or U7222 (N_7222,N_4091,N_1675);
nand U7223 (N_7223,N_3387,N_2123);
or U7224 (N_7224,N_2513,N_2381);
nor U7225 (N_7225,N_2986,N_666);
or U7226 (N_7226,N_3689,N_3748);
and U7227 (N_7227,N_4863,N_625);
and U7228 (N_7228,N_1190,N_4850);
and U7229 (N_7229,N_4025,N_1770);
nand U7230 (N_7230,N_3088,N_3747);
or U7231 (N_7231,N_4257,N_2734);
nand U7232 (N_7232,N_1959,N_1386);
nor U7233 (N_7233,N_341,N_1334);
and U7234 (N_7234,N_4809,N_526);
or U7235 (N_7235,N_1913,N_1099);
nand U7236 (N_7236,N_4165,N_3555);
nor U7237 (N_7237,N_360,N_3814);
or U7238 (N_7238,N_1520,N_2591);
nand U7239 (N_7239,N_3085,N_3710);
and U7240 (N_7240,N_4816,N_3520);
nor U7241 (N_7241,N_4979,N_2298);
or U7242 (N_7242,N_978,N_1345);
and U7243 (N_7243,N_2748,N_3012);
or U7244 (N_7244,N_1713,N_3959);
nor U7245 (N_7245,N_381,N_3957);
or U7246 (N_7246,N_1202,N_383);
nand U7247 (N_7247,N_4472,N_68);
or U7248 (N_7248,N_2800,N_4086);
and U7249 (N_7249,N_153,N_536);
and U7250 (N_7250,N_303,N_4836);
nand U7251 (N_7251,N_1566,N_2867);
nand U7252 (N_7252,N_493,N_852);
or U7253 (N_7253,N_4538,N_678);
nor U7254 (N_7254,N_2958,N_2394);
or U7255 (N_7255,N_4218,N_2193);
nor U7256 (N_7256,N_2706,N_1885);
nor U7257 (N_7257,N_2118,N_3198);
nand U7258 (N_7258,N_22,N_2359);
nor U7259 (N_7259,N_627,N_4114);
and U7260 (N_7260,N_773,N_2432);
nor U7261 (N_7261,N_2033,N_1664);
and U7262 (N_7262,N_240,N_268);
or U7263 (N_7263,N_2302,N_1599);
nand U7264 (N_7264,N_2742,N_4657);
nand U7265 (N_7265,N_418,N_734);
and U7266 (N_7266,N_2525,N_549);
and U7267 (N_7267,N_4640,N_3319);
or U7268 (N_7268,N_2322,N_3264);
nor U7269 (N_7269,N_4896,N_2253);
or U7270 (N_7270,N_1053,N_2819);
nor U7271 (N_7271,N_156,N_2202);
or U7272 (N_7272,N_1230,N_2644);
or U7273 (N_7273,N_3170,N_1533);
or U7274 (N_7274,N_1354,N_3116);
or U7275 (N_7275,N_3996,N_2282);
or U7276 (N_7276,N_3521,N_1187);
or U7277 (N_7277,N_1838,N_3358);
or U7278 (N_7278,N_4469,N_285);
or U7279 (N_7279,N_2074,N_1096);
nand U7280 (N_7280,N_1006,N_3774);
nand U7281 (N_7281,N_702,N_3363);
and U7282 (N_7282,N_1592,N_2661);
nor U7283 (N_7283,N_1330,N_950);
nand U7284 (N_7284,N_604,N_3932);
nor U7285 (N_7285,N_1535,N_1750);
or U7286 (N_7286,N_181,N_1126);
and U7287 (N_7287,N_3271,N_3607);
or U7288 (N_7288,N_13,N_4274);
nor U7289 (N_7289,N_1339,N_2310);
xor U7290 (N_7290,N_4357,N_3162);
and U7291 (N_7291,N_3786,N_3108);
and U7292 (N_7292,N_1062,N_2297);
nand U7293 (N_7293,N_3941,N_882);
and U7294 (N_7294,N_2786,N_1361);
and U7295 (N_7295,N_3221,N_4936);
or U7296 (N_7296,N_2023,N_1358);
nand U7297 (N_7297,N_1621,N_2872);
nand U7298 (N_7298,N_4180,N_3029);
or U7299 (N_7299,N_872,N_516);
or U7300 (N_7300,N_4606,N_1808);
nor U7301 (N_7301,N_4621,N_1179);
nand U7302 (N_7302,N_634,N_538);
and U7303 (N_7303,N_266,N_1424);
or U7304 (N_7304,N_4673,N_1508);
or U7305 (N_7305,N_4189,N_960);
nor U7306 (N_7306,N_3653,N_2680);
or U7307 (N_7307,N_2428,N_3388);
nor U7308 (N_7308,N_4012,N_1296);
nor U7309 (N_7309,N_1151,N_1865);
nand U7310 (N_7310,N_4440,N_4853);
nor U7311 (N_7311,N_2848,N_3421);
nand U7312 (N_7312,N_4298,N_2856);
nor U7313 (N_7313,N_1576,N_3862);
and U7314 (N_7314,N_739,N_199);
nand U7315 (N_7315,N_3868,N_2654);
nor U7316 (N_7316,N_4351,N_151);
and U7317 (N_7317,N_1715,N_440);
and U7318 (N_7318,N_4200,N_2077);
or U7319 (N_7319,N_4813,N_3355);
and U7320 (N_7320,N_490,N_4396);
and U7321 (N_7321,N_4303,N_4552);
nor U7322 (N_7322,N_3580,N_2846);
or U7323 (N_7323,N_1665,N_1966);
or U7324 (N_7324,N_3912,N_180);
nand U7325 (N_7325,N_4916,N_2707);
and U7326 (N_7326,N_1082,N_530);
nand U7327 (N_7327,N_3030,N_966);
or U7328 (N_7328,N_2293,N_1753);
nand U7329 (N_7329,N_2153,N_2853);
or U7330 (N_7330,N_2753,N_2626);
nor U7331 (N_7331,N_3371,N_4917);
nor U7332 (N_7332,N_1360,N_1270);
nand U7333 (N_7333,N_948,N_3573);
or U7334 (N_7334,N_4339,N_3610);
or U7335 (N_7335,N_486,N_1647);
xor U7336 (N_7336,N_1506,N_4451);
nand U7337 (N_7337,N_3900,N_3097);
nor U7338 (N_7338,N_1128,N_3993);
nand U7339 (N_7339,N_3026,N_51);
and U7340 (N_7340,N_1347,N_416);
nand U7341 (N_7341,N_1663,N_2008);
or U7342 (N_7342,N_1733,N_2022);
or U7343 (N_7343,N_3456,N_2048);
nand U7344 (N_7344,N_949,N_667);
nand U7345 (N_7345,N_2125,N_1912);
nor U7346 (N_7346,N_694,N_3715);
and U7347 (N_7347,N_2978,N_204);
and U7348 (N_7348,N_1309,N_2797);
or U7349 (N_7349,N_3726,N_3075);
and U7350 (N_7350,N_1712,N_1323);
and U7351 (N_7351,N_2520,N_3849);
nor U7352 (N_7352,N_4749,N_4544);
or U7353 (N_7353,N_4854,N_2075);
and U7354 (N_7354,N_1008,N_4345);
nor U7355 (N_7355,N_1127,N_4259);
nor U7356 (N_7356,N_4042,N_3899);
nor U7357 (N_7357,N_1553,N_4834);
or U7358 (N_7358,N_3526,N_3155);
nand U7359 (N_7359,N_131,N_4295);
or U7360 (N_7360,N_2929,N_482);
or U7361 (N_7361,N_1897,N_2290);
nor U7362 (N_7362,N_2920,N_1645);
or U7363 (N_7363,N_2757,N_2959);
nand U7364 (N_7364,N_1872,N_3668);
or U7365 (N_7365,N_293,N_3923);
and U7366 (N_7366,N_1969,N_4721);
nor U7367 (N_7367,N_3279,N_4246);
nor U7368 (N_7368,N_2533,N_2149);
nor U7369 (N_7369,N_294,N_4133);
and U7370 (N_7370,N_3343,N_3939);
nor U7371 (N_7371,N_3915,N_4093);
nor U7372 (N_7372,N_559,N_201);
nand U7373 (N_7373,N_4021,N_129);
or U7374 (N_7374,N_3508,N_3348);
nand U7375 (N_7375,N_2305,N_4113);
and U7376 (N_7376,N_826,N_1703);
and U7377 (N_7377,N_2327,N_1491);
nand U7378 (N_7378,N_3944,N_4051);
xnor U7379 (N_7379,N_3022,N_1426);
or U7380 (N_7380,N_649,N_1877);
nand U7381 (N_7381,N_2859,N_484);
nand U7382 (N_7382,N_4572,N_1266);
xnor U7383 (N_7383,N_854,N_3547);
nand U7384 (N_7384,N_3509,N_3190);
or U7385 (N_7385,N_817,N_4662);
nand U7386 (N_7386,N_1529,N_4759);
and U7387 (N_7387,N_4287,N_545);
nor U7388 (N_7388,N_565,N_810);
nand U7389 (N_7389,N_3373,N_4963);
nand U7390 (N_7390,N_1469,N_227);
or U7391 (N_7391,N_4264,N_4150);
and U7392 (N_7392,N_757,N_223);
and U7393 (N_7393,N_732,N_4336);
and U7394 (N_7394,N_2063,N_1033);
nor U7395 (N_7395,N_552,N_2169);
nor U7396 (N_7396,N_2871,N_3461);
nand U7397 (N_7397,N_4102,N_2466);
or U7398 (N_7398,N_4146,N_1563);
and U7399 (N_7399,N_864,N_3321);
or U7400 (N_7400,N_4479,N_1618);
or U7401 (N_7401,N_4803,N_465);
nor U7402 (N_7402,N_768,N_1623);
nor U7403 (N_7403,N_4949,N_3705);
or U7404 (N_7404,N_689,N_2189);
or U7405 (N_7405,N_2825,N_2649);
nor U7406 (N_7406,N_145,N_1063);
or U7407 (N_7407,N_2904,N_426);
nand U7408 (N_7408,N_657,N_4141);
or U7409 (N_7409,N_2973,N_3802);
or U7410 (N_7410,N_81,N_4170);
nand U7411 (N_7411,N_3707,N_2427);
nor U7412 (N_7412,N_772,N_1113);
nand U7413 (N_7413,N_3078,N_2790);
nor U7414 (N_7414,N_384,N_4378);
nor U7415 (N_7415,N_4169,N_3537);
or U7416 (N_7416,N_1014,N_2163);
and U7417 (N_7417,N_16,N_3655);
and U7418 (N_7418,N_4166,N_3585);
or U7419 (N_7419,N_3935,N_377);
or U7420 (N_7420,N_2669,N_2449);
and U7421 (N_7421,N_3256,N_2544);
or U7422 (N_7422,N_3366,N_4352);
or U7423 (N_7423,N_1495,N_2279);
or U7424 (N_7424,N_2783,N_2968);
nand U7425 (N_7425,N_4296,N_1882);
nand U7426 (N_7426,N_4810,N_4383);
nand U7427 (N_7427,N_468,N_1864);
or U7428 (N_7428,N_2013,N_1473);
or U7429 (N_7429,N_875,N_1778);
nor U7430 (N_7430,N_610,N_3572);
or U7431 (N_7431,N_4391,N_821);
and U7432 (N_7432,N_2486,N_3411);
and U7433 (N_7433,N_4044,N_3460);
nand U7434 (N_7434,N_4338,N_1510);
nor U7435 (N_7435,N_1461,N_2838);
or U7436 (N_7436,N_1312,N_509);
nand U7437 (N_7437,N_589,N_4379);
or U7438 (N_7438,N_3390,N_3224);
and U7439 (N_7439,N_4537,N_239);
or U7440 (N_7440,N_168,N_4250);
nand U7441 (N_7441,N_4010,N_4447);
nor U7442 (N_7442,N_2078,N_4050);
and U7443 (N_7443,N_2107,N_4271);
or U7444 (N_7444,N_291,N_467);
nor U7445 (N_7445,N_3297,N_3052);
or U7446 (N_7446,N_3619,N_755);
or U7447 (N_7447,N_1398,N_1307);
and U7448 (N_7448,N_1092,N_3277);
nand U7449 (N_7449,N_292,N_4491);
nand U7450 (N_7450,N_1816,N_1037);
and U7451 (N_7451,N_4135,N_3269);
nor U7452 (N_7452,N_2138,N_2079);
nand U7453 (N_7453,N_3499,N_3492);
and U7454 (N_7454,N_3730,N_282);
nand U7455 (N_7455,N_669,N_478);
nor U7456 (N_7456,N_3128,N_4373);
or U7457 (N_7457,N_2714,N_1890);
and U7458 (N_7458,N_252,N_1084);
nor U7459 (N_7459,N_1038,N_2320);
nor U7460 (N_7460,N_629,N_868);
and U7461 (N_7461,N_1933,N_1385);
and U7462 (N_7462,N_1590,N_3788);
nor U7463 (N_7463,N_4878,N_2506);
or U7464 (N_7464,N_4031,N_2148);
nor U7465 (N_7465,N_1731,N_2961);
or U7466 (N_7466,N_595,N_3505);
and U7467 (N_7467,N_1346,N_1825);
and U7468 (N_7468,N_1114,N_2053);
and U7469 (N_7469,N_3906,N_998);
and U7470 (N_7470,N_3349,N_3853);
or U7471 (N_7471,N_2375,N_259);
nand U7472 (N_7472,N_1349,N_4448);
and U7473 (N_7473,N_3274,N_4415);
nand U7474 (N_7474,N_1453,N_4932);
and U7475 (N_7475,N_3234,N_1463);
nor U7476 (N_7476,N_1456,N_4106);
nand U7477 (N_7477,N_4372,N_539);
and U7478 (N_7478,N_588,N_2277);
or U7479 (N_7479,N_3854,N_4525);
or U7480 (N_7480,N_4644,N_4069);
or U7481 (N_7481,N_297,N_2532);
nand U7482 (N_7482,N_693,N_1849);
or U7483 (N_7483,N_4273,N_2336);
nand U7484 (N_7484,N_1941,N_1257);
and U7485 (N_7485,N_4475,N_2004);
nor U7486 (N_7486,N_311,N_2386);
and U7487 (N_7487,N_2446,N_4002);
and U7488 (N_7488,N_1031,N_3896);
nand U7489 (N_7489,N_4236,N_3459);
nand U7490 (N_7490,N_2144,N_1236);
and U7491 (N_7491,N_3946,N_4665);
nand U7492 (N_7492,N_1704,N_1069);
or U7493 (N_7493,N_1942,N_1303);
or U7494 (N_7494,N_2563,N_3785);
nand U7495 (N_7495,N_4155,N_3737);
and U7496 (N_7496,N_161,N_194);
or U7497 (N_7497,N_169,N_1478);
or U7498 (N_7498,N_4978,N_859);
nand U7499 (N_7499,N_4482,N_3952);
and U7500 (N_7500,N_3733,N_867);
or U7501 (N_7501,N_1054,N_1537);
nand U7502 (N_7502,N_719,N_4401);
or U7503 (N_7503,N_98,N_1876);
or U7504 (N_7504,N_4022,N_1883);
xnor U7505 (N_7505,N_246,N_3960);
nor U7506 (N_7506,N_4684,N_3134);
and U7507 (N_7507,N_1656,N_4245);
nand U7508 (N_7508,N_2472,N_2935);
nor U7509 (N_7509,N_202,N_4285);
or U7510 (N_7510,N_3844,N_4371);
nor U7511 (N_7511,N_3052,N_4135);
nand U7512 (N_7512,N_668,N_1283);
and U7513 (N_7513,N_3197,N_3265);
nor U7514 (N_7514,N_556,N_4899);
and U7515 (N_7515,N_4287,N_3796);
and U7516 (N_7516,N_1901,N_1300);
nand U7517 (N_7517,N_4807,N_3987);
or U7518 (N_7518,N_1970,N_853);
nor U7519 (N_7519,N_2010,N_4433);
or U7520 (N_7520,N_4348,N_611);
and U7521 (N_7521,N_2840,N_1251);
nand U7522 (N_7522,N_4997,N_1782);
or U7523 (N_7523,N_1935,N_4476);
and U7524 (N_7524,N_2780,N_1443);
or U7525 (N_7525,N_1800,N_1171);
and U7526 (N_7526,N_990,N_4611);
nand U7527 (N_7527,N_942,N_2721);
nand U7528 (N_7528,N_4599,N_3231);
nor U7529 (N_7529,N_803,N_1453);
nand U7530 (N_7530,N_2161,N_4071);
and U7531 (N_7531,N_1809,N_1125);
and U7532 (N_7532,N_1152,N_3698);
nor U7533 (N_7533,N_4161,N_4115);
and U7534 (N_7534,N_1740,N_840);
nor U7535 (N_7535,N_867,N_1835);
nand U7536 (N_7536,N_1649,N_4469);
or U7537 (N_7537,N_309,N_1759);
or U7538 (N_7538,N_718,N_2248);
and U7539 (N_7539,N_1272,N_1303);
xnor U7540 (N_7540,N_2199,N_2400);
nand U7541 (N_7541,N_3691,N_2247);
and U7542 (N_7542,N_3729,N_4855);
nor U7543 (N_7543,N_1272,N_369);
or U7544 (N_7544,N_2872,N_4458);
or U7545 (N_7545,N_4238,N_1203);
nand U7546 (N_7546,N_2677,N_2143);
and U7547 (N_7547,N_2110,N_3241);
nor U7548 (N_7548,N_1543,N_4402);
and U7549 (N_7549,N_1448,N_1798);
nand U7550 (N_7550,N_1766,N_4086);
nand U7551 (N_7551,N_2312,N_4176);
or U7552 (N_7552,N_825,N_3123);
xnor U7553 (N_7553,N_4163,N_692);
nand U7554 (N_7554,N_3295,N_3711);
and U7555 (N_7555,N_2286,N_4580);
and U7556 (N_7556,N_1923,N_2517);
nor U7557 (N_7557,N_4651,N_4632);
nor U7558 (N_7558,N_4959,N_2296);
nor U7559 (N_7559,N_1861,N_2624);
and U7560 (N_7560,N_2951,N_2608);
and U7561 (N_7561,N_4610,N_2361);
or U7562 (N_7562,N_2851,N_1642);
nor U7563 (N_7563,N_1579,N_823);
and U7564 (N_7564,N_2200,N_4204);
and U7565 (N_7565,N_1401,N_4891);
nor U7566 (N_7566,N_4297,N_4967);
nand U7567 (N_7567,N_2688,N_2228);
or U7568 (N_7568,N_1302,N_4864);
or U7569 (N_7569,N_691,N_462);
nand U7570 (N_7570,N_2522,N_1672);
and U7571 (N_7571,N_3782,N_2838);
or U7572 (N_7572,N_3372,N_3102);
nand U7573 (N_7573,N_147,N_4553);
or U7574 (N_7574,N_4871,N_1153);
or U7575 (N_7575,N_285,N_4020);
nor U7576 (N_7576,N_1514,N_1199);
and U7577 (N_7577,N_880,N_3860);
or U7578 (N_7578,N_3439,N_4558);
and U7579 (N_7579,N_2491,N_3306);
nor U7580 (N_7580,N_3191,N_3592);
and U7581 (N_7581,N_1096,N_4290);
nand U7582 (N_7582,N_3546,N_2159);
or U7583 (N_7583,N_1926,N_4412);
nand U7584 (N_7584,N_864,N_2273);
nand U7585 (N_7585,N_3861,N_3272);
nand U7586 (N_7586,N_3056,N_4727);
or U7587 (N_7587,N_2676,N_1335);
or U7588 (N_7588,N_4038,N_3005);
nor U7589 (N_7589,N_1124,N_3909);
and U7590 (N_7590,N_4408,N_3152);
or U7591 (N_7591,N_3373,N_3994);
nor U7592 (N_7592,N_2862,N_757);
or U7593 (N_7593,N_1127,N_783);
or U7594 (N_7594,N_4001,N_1988);
and U7595 (N_7595,N_251,N_1649);
nor U7596 (N_7596,N_3246,N_3938);
and U7597 (N_7597,N_2575,N_4142);
and U7598 (N_7598,N_2094,N_2463);
and U7599 (N_7599,N_4879,N_3474);
or U7600 (N_7600,N_1580,N_2398);
nand U7601 (N_7601,N_1854,N_1166);
nand U7602 (N_7602,N_3041,N_4301);
nand U7603 (N_7603,N_3753,N_2694);
or U7604 (N_7604,N_140,N_1569);
and U7605 (N_7605,N_3582,N_1458);
nor U7606 (N_7606,N_1646,N_458);
nor U7607 (N_7607,N_351,N_2873);
and U7608 (N_7608,N_950,N_957);
and U7609 (N_7609,N_2227,N_3363);
or U7610 (N_7610,N_4536,N_1493);
and U7611 (N_7611,N_3803,N_553);
and U7612 (N_7612,N_1793,N_2315);
nand U7613 (N_7613,N_1937,N_2326);
nor U7614 (N_7614,N_4301,N_1668);
and U7615 (N_7615,N_2266,N_4271);
nor U7616 (N_7616,N_88,N_4376);
nor U7617 (N_7617,N_3673,N_3070);
or U7618 (N_7618,N_1640,N_3399);
nor U7619 (N_7619,N_3468,N_474);
nor U7620 (N_7620,N_331,N_510);
nand U7621 (N_7621,N_1465,N_1723);
or U7622 (N_7622,N_1835,N_4232);
nor U7623 (N_7623,N_3214,N_3494);
and U7624 (N_7624,N_448,N_3565);
or U7625 (N_7625,N_3571,N_3891);
nand U7626 (N_7626,N_213,N_1119);
nand U7627 (N_7627,N_2234,N_2411);
nor U7628 (N_7628,N_332,N_1470);
and U7629 (N_7629,N_3065,N_2992);
or U7630 (N_7630,N_4800,N_2299);
and U7631 (N_7631,N_1336,N_4988);
nand U7632 (N_7632,N_4475,N_4225);
nor U7633 (N_7633,N_2096,N_3521);
and U7634 (N_7634,N_6,N_4789);
or U7635 (N_7635,N_1914,N_4516);
nor U7636 (N_7636,N_3431,N_3700);
nand U7637 (N_7637,N_3163,N_1071);
or U7638 (N_7638,N_826,N_3140);
and U7639 (N_7639,N_1384,N_1402);
and U7640 (N_7640,N_1248,N_3508);
or U7641 (N_7641,N_3389,N_1636);
nand U7642 (N_7642,N_3308,N_519);
nor U7643 (N_7643,N_3626,N_4954);
or U7644 (N_7644,N_3851,N_894);
and U7645 (N_7645,N_2666,N_1095);
or U7646 (N_7646,N_4498,N_2102);
and U7647 (N_7647,N_4335,N_1591);
or U7648 (N_7648,N_2833,N_1693);
nor U7649 (N_7649,N_255,N_4869);
or U7650 (N_7650,N_3804,N_2954);
nand U7651 (N_7651,N_1002,N_4811);
nand U7652 (N_7652,N_1230,N_670);
and U7653 (N_7653,N_1368,N_2420);
or U7654 (N_7654,N_2007,N_1043);
nor U7655 (N_7655,N_3193,N_1716);
nand U7656 (N_7656,N_2289,N_2409);
and U7657 (N_7657,N_4296,N_817);
or U7658 (N_7658,N_1683,N_1926);
nand U7659 (N_7659,N_1012,N_4762);
nor U7660 (N_7660,N_2227,N_1538);
and U7661 (N_7661,N_1920,N_2776);
or U7662 (N_7662,N_4104,N_4242);
and U7663 (N_7663,N_316,N_3405);
or U7664 (N_7664,N_2125,N_44);
nor U7665 (N_7665,N_2898,N_963);
nand U7666 (N_7666,N_2615,N_2123);
or U7667 (N_7667,N_2895,N_3570);
or U7668 (N_7668,N_4303,N_582);
nor U7669 (N_7669,N_701,N_4645);
or U7670 (N_7670,N_1407,N_1849);
nor U7671 (N_7671,N_4335,N_756);
and U7672 (N_7672,N_3429,N_1273);
and U7673 (N_7673,N_1928,N_3372);
or U7674 (N_7674,N_3032,N_2355);
and U7675 (N_7675,N_3091,N_512);
and U7676 (N_7676,N_490,N_51);
or U7677 (N_7677,N_197,N_1518);
or U7678 (N_7678,N_1521,N_3059);
and U7679 (N_7679,N_1173,N_1073);
nor U7680 (N_7680,N_2560,N_2259);
nor U7681 (N_7681,N_767,N_3834);
nor U7682 (N_7682,N_2996,N_3241);
or U7683 (N_7683,N_1862,N_2199);
nand U7684 (N_7684,N_4496,N_2954);
nand U7685 (N_7685,N_3135,N_4120);
or U7686 (N_7686,N_1955,N_447);
and U7687 (N_7687,N_3101,N_4186);
and U7688 (N_7688,N_2681,N_1330);
nand U7689 (N_7689,N_2968,N_3203);
or U7690 (N_7690,N_2599,N_279);
or U7691 (N_7691,N_4454,N_2689);
or U7692 (N_7692,N_335,N_2223);
nand U7693 (N_7693,N_3324,N_2112);
or U7694 (N_7694,N_1546,N_3760);
nand U7695 (N_7695,N_1740,N_1314);
nor U7696 (N_7696,N_3564,N_4321);
and U7697 (N_7697,N_2172,N_2019);
or U7698 (N_7698,N_4904,N_957);
and U7699 (N_7699,N_3321,N_3369);
or U7700 (N_7700,N_3994,N_3560);
and U7701 (N_7701,N_4024,N_3303);
nand U7702 (N_7702,N_4604,N_974);
or U7703 (N_7703,N_471,N_4033);
nor U7704 (N_7704,N_1256,N_2952);
nor U7705 (N_7705,N_313,N_4466);
nor U7706 (N_7706,N_3052,N_1003);
and U7707 (N_7707,N_3718,N_839);
and U7708 (N_7708,N_3447,N_1468);
nand U7709 (N_7709,N_1884,N_2540);
nor U7710 (N_7710,N_4240,N_992);
nor U7711 (N_7711,N_1548,N_4765);
and U7712 (N_7712,N_4171,N_3604);
nor U7713 (N_7713,N_3451,N_2140);
nor U7714 (N_7714,N_4795,N_3051);
and U7715 (N_7715,N_4108,N_1915);
and U7716 (N_7716,N_396,N_1657);
nand U7717 (N_7717,N_791,N_1500);
or U7718 (N_7718,N_4500,N_3337);
or U7719 (N_7719,N_2856,N_775);
nor U7720 (N_7720,N_2055,N_4387);
xnor U7721 (N_7721,N_710,N_4645);
or U7722 (N_7722,N_1527,N_786);
and U7723 (N_7723,N_3294,N_4474);
nor U7724 (N_7724,N_563,N_2429);
nor U7725 (N_7725,N_1817,N_1693);
nand U7726 (N_7726,N_1486,N_683);
nor U7727 (N_7727,N_4734,N_2529);
nand U7728 (N_7728,N_2863,N_3598);
or U7729 (N_7729,N_160,N_4837);
nor U7730 (N_7730,N_3710,N_2016);
nor U7731 (N_7731,N_1617,N_3205);
nand U7732 (N_7732,N_3691,N_2422);
and U7733 (N_7733,N_4287,N_3504);
and U7734 (N_7734,N_3886,N_3728);
and U7735 (N_7735,N_2332,N_43);
nor U7736 (N_7736,N_1074,N_37);
nand U7737 (N_7737,N_4684,N_1741);
and U7738 (N_7738,N_2685,N_3720);
or U7739 (N_7739,N_3326,N_3992);
nor U7740 (N_7740,N_2080,N_2883);
nor U7741 (N_7741,N_26,N_411);
nand U7742 (N_7742,N_399,N_1163);
nor U7743 (N_7743,N_3721,N_287);
or U7744 (N_7744,N_1429,N_1306);
or U7745 (N_7745,N_3709,N_4389);
or U7746 (N_7746,N_3355,N_3056);
and U7747 (N_7747,N_3383,N_1921);
and U7748 (N_7748,N_3699,N_1358);
and U7749 (N_7749,N_1155,N_4897);
nand U7750 (N_7750,N_1685,N_3023);
or U7751 (N_7751,N_3949,N_3487);
or U7752 (N_7752,N_890,N_4072);
and U7753 (N_7753,N_4637,N_2345);
nor U7754 (N_7754,N_1876,N_2312);
nor U7755 (N_7755,N_439,N_2195);
and U7756 (N_7756,N_4700,N_2156);
nor U7757 (N_7757,N_3893,N_925);
and U7758 (N_7758,N_324,N_2633);
nand U7759 (N_7759,N_1257,N_2764);
and U7760 (N_7760,N_2928,N_447);
or U7761 (N_7761,N_1712,N_656);
nor U7762 (N_7762,N_1947,N_730);
nor U7763 (N_7763,N_1241,N_3594);
nand U7764 (N_7764,N_1143,N_298);
and U7765 (N_7765,N_218,N_2131);
and U7766 (N_7766,N_189,N_4718);
nor U7767 (N_7767,N_1571,N_2684);
or U7768 (N_7768,N_603,N_4698);
or U7769 (N_7769,N_4205,N_1475);
nand U7770 (N_7770,N_1511,N_2082);
or U7771 (N_7771,N_605,N_4560);
xor U7772 (N_7772,N_2033,N_2733);
and U7773 (N_7773,N_3250,N_3124);
nor U7774 (N_7774,N_2649,N_2259);
nand U7775 (N_7775,N_2063,N_4955);
nor U7776 (N_7776,N_3074,N_4647);
nand U7777 (N_7777,N_4986,N_3334);
nor U7778 (N_7778,N_2923,N_2065);
or U7779 (N_7779,N_1647,N_208);
xor U7780 (N_7780,N_989,N_1342);
nand U7781 (N_7781,N_3965,N_69);
nor U7782 (N_7782,N_1661,N_4645);
nor U7783 (N_7783,N_878,N_4890);
xor U7784 (N_7784,N_972,N_20);
nor U7785 (N_7785,N_2921,N_1532);
nor U7786 (N_7786,N_3090,N_347);
nand U7787 (N_7787,N_1001,N_385);
or U7788 (N_7788,N_395,N_3122);
nor U7789 (N_7789,N_3239,N_1996);
or U7790 (N_7790,N_730,N_3175);
nand U7791 (N_7791,N_2768,N_1564);
and U7792 (N_7792,N_3746,N_2581);
nand U7793 (N_7793,N_1541,N_4515);
xnor U7794 (N_7794,N_387,N_559);
and U7795 (N_7795,N_3203,N_348);
and U7796 (N_7796,N_4381,N_3228);
nand U7797 (N_7797,N_1704,N_3776);
or U7798 (N_7798,N_3308,N_228);
nor U7799 (N_7799,N_2481,N_1021);
or U7800 (N_7800,N_2867,N_3667);
and U7801 (N_7801,N_1454,N_3104);
and U7802 (N_7802,N_2095,N_3404);
nand U7803 (N_7803,N_3765,N_4942);
or U7804 (N_7804,N_4672,N_3570);
nand U7805 (N_7805,N_10,N_676);
or U7806 (N_7806,N_4507,N_1718);
nand U7807 (N_7807,N_698,N_4160);
nand U7808 (N_7808,N_2823,N_1167);
nand U7809 (N_7809,N_1331,N_1662);
and U7810 (N_7810,N_531,N_94);
nand U7811 (N_7811,N_265,N_3833);
nand U7812 (N_7812,N_518,N_4008);
nor U7813 (N_7813,N_2926,N_358);
or U7814 (N_7814,N_548,N_1833);
and U7815 (N_7815,N_4197,N_2995);
nor U7816 (N_7816,N_2584,N_4051);
nor U7817 (N_7817,N_3103,N_3931);
and U7818 (N_7818,N_2005,N_967);
nor U7819 (N_7819,N_3428,N_3644);
nor U7820 (N_7820,N_1365,N_951);
and U7821 (N_7821,N_3683,N_4124);
and U7822 (N_7822,N_2664,N_4734);
nor U7823 (N_7823,N_2740,N_3745);
nand U7824 (N_7824,N_483,N_785);
or U7825 (N_7825,N_73,N_1245);
nand U7826 (N_7826,N_3004,N_2710);
or U7827 (N_7827,N_4286,N_3716);
nor U7828 (N_7828,N_4063,N_2662);
nor U7829 (N_7829,N_4728,N_3205);
and U7830 (N_7830,N_2554,N_1435);
and U7831 (N_7831,N_1190,N_4879);
nor U7832 (N_7832,N_4548,N_2777);
nor U7833 (N_7833,N_3547,N_1780);
nand U7834 (N_7834,N_3548,N_676);
nor U7835 (N_7835,N_2734,N_4994);
xor U7836 (N_7836,N_741,N_4941);
and U7837 (N_7837,N_4560,N_1797);
and U7838 (N_7838,N_1175,N_4215);
nand U7839 (N_7839,N_728,N_2791);
and U7840 (N_7840,N_3429,N_3774);
nor U7841 (N_7841,N_4832,N_1213);
or U7842 (N_7842,N_4541,N_2551);
and U7843 (N_7843,N_288,N_508);
and U7844 (N_7844,N_1853,N_2805);
and U7845 (N_7845,N_1465,N_3014);
nor U7846 (N_7846,N_2487,N_2772);
nand U7847 (N_7847,N_2522,N_4864);
and U7848 (N_7848,N_2600,N_1474);
and U7849 (N_7849,N_28,N_1238);
nand U7850 (N_7850,N_1460,N_364);
nor U7851 (N_7851,N_57,N_2691);
or U7852 (N_7852,N_257,N_4252);
and U7853 (N_7853,N_3755,N_3632);
nand U7854 (N_7854,N_1502,N_3757);
and U7855 (N_7855,N_2350,N_1756);
nor U7856 (N_7856,N_2799,N_2681);
nor U7857 (N_7857,N_2597,N_4192);
nor U7858 (N_7858,N_1351,N_4865);
nand U7859 (N_7859,N_2118,N_4689);
and U7860 (N_7860,N_1652,N_2423);
nor U7861 (N_7861,N_4888,N_1332);
nand U7862 (N_7862,N_2130,N_3343);
and U7863 (N_7863,N_3575,N_4879);
or U7864 (N_7864,N_2502,N_405);
nor U7865 (N_7865,N_611,N_976);
nor U7866 (N_7866,N_4739,N_1438);
nand U7867 (N_7867,N_1344,N_524);
nand U7868 (N_7868,N_805,N_2899);
nor U7869 (N_7869,N_1236,N_2986);
nor U7870 (N_7870,N_1236,N_2083);
or U7871 (N_7871,N_4545,N_2369);
and U7872 (N_7872,N_1438,N_4226);
nand U7873 (N_7873,N_2665,N_4446);
nand U7874 (N_7874,N_1682,N_883);
nand U7875 (N_7875,N_1610,N_4992);
nand U7876 (N_7876,N_3737,N_4125);
or U7877 (N_7877,N_4492,N_806);
or U7878 (N_7878,N_964,N_50);
nand U7879 (N_7879,N_432,N_3881);
nand U7880 (N_7880,N_1609,N_3154);
or U7881 (N_7881,N_4507,N_4401);
or U7882 (N_7882,N_558,N_4853);
nand U7883 (N_7883,N_3020,N_4458);
and U7884 (N_7884,N_2136,N_464);
nand U7885 (N_7885,N_3731,N_4192);
or U7886 (N_7886,N_1081,N_3233);
or U7887 (N_7887,N_4173,N_1579);
and U7888 (N_7888,N_166,N_4579);
and U7889 (N_7889,N_2169,N_4289);
or U7890 (N_7890,N_4750,N_4599);
or U7891 (N_7891,N_1016,N_4762);
xnor U7892 (N_7892,N_3196,N_4266);
or U7893 (N_7893,N_4342,N_1231);
or U7894 (N_7894,N_3976,N_645);
or U7895 (N_7895,N_1571,N_2329);
or U7896 (N_7896,N_1763,N_4462);
nand U7897 (N_7897,N_56,N_3099);
or U7898 (N_7898,N_997,N_3140);
or U7899 (N_7899,N_1105,N_4938);
nor U7900 (N_7900,N_3195,N_1477);
nor U7901 (N_7901,N_2832,N_1464);
nor U7902 (N_7902,N_4965,N_1919);
nand U7903 (N_7903,N_3432,N_3693);
nor U7904 (N_7904,N_2992,N_1591);
and U7905 (N_7905,N_4274,N_1207);
nand U7906 (N_7906,N_1736,N_1005);
nor U7907 (N_7907,N_20,N_2679);
nand U7908 (N_7908,N_3953,N_1243);
and U7909 (N_7909,N_2437,N_2999);
nand U7910 (N_7910,N_4,N_2990);
and U7911 (N_7911,N_377,N_1826);
nand U7912 (N_7912,N_1968,N_843);
nand U7913 (N_7913,N_1397,N_3102);
and U7914 (N_7914,N_3126,N_805);
or U7915 (N_7915,N_3914,N_2245);
and U7916 (N_7916,N_2514,N_2481);
and U7917 (N_7917,N_534,N_1137);
nor U7918 (N_7918,N_3457,N_1934);
nand U7919 (N_7919,N_1877,N_4666);
nor U7920 (N_7920,N_805,N_626);
nand U7921 (N_7921,N_894,N_1580);
and U7922 (N_7922,N_2270,N_1907);
nand U7923 (N_7923,N_399,N_4387);
nand U7924 (N_7924,N_3518,N_4854);
nor U7925 (N_7925,N_2092,N_3431);
nand U7926 (N_7926,N_1245,N_4735);
nand U7927 (N_7927,N_4281,N_4248);
and U7928 (N_7928,N_2048,N_3851);
and U7929 (N_7929,N_4228,N_309);
or U7930 (N_7930,N_897,N_3329);
and U7931 (N_7931,N_3900,N_3122);
nor U7932 (N_7932,N_4150,N_3110);
and U7933 (N_7933,N_1948,N_1479);
nand U7934 (N_7934,N_3706,N_4176);
xnor U7935 (N_7935,N_3853,N_2253);
nor U7936 (N_7936,N_775,N_2891);
nand U7937 (N_7937,N_2299,N_2222);
nor U7938 (N_7938,N_3836,N_3493);
and U7939 (N_7939,N_4250,N_3007);
nor U7940 (N_7940,N_980,N_3828);
and U7941 (N_7941,N_2447,N_2638);
nor U7942 (N_7942,N_1853,N_3967);
and U7943 (N_7943,N_3543,N_247);
or U7944 (N_7944,N_3840,N_4264);
and U7945 (N_7945,N_463,N_3745);
nor U7946 (N_7946,N_3425,N_3887);
nand U7947 (N_7947,N_728,N_399);
nand U7948 (N_7948,N_1051,N_68);
nand U7949 (N_7949,N_3753,N_4933);
and U7950 (N_7950,N_1164,N_4687);
or U7951 (N_7951,N_3870,N_3349);
nand U7952 (N_7952,N_1448,N_1694);
nor U7953 (N_7953,N_4161,N_554);
nand U7954 (N_7954,N_1681,N_930);
nor U7955 (N_7955,N_918,N_3212);
and U7956 (N_7956,N_1884,N_227);
nor U7957 (N_7957,N_3404,N_979);
nand U7958 (N_7958,N_4658,N_3103);
nor U7959 (N_7959,N_434,N_2733);
nor U7960 (N_7960,N_1386,N_3312);
nor U7961 (N_7961,N_145,N_4908);
and U7962 (N_7962,N_1616,N_2863);
or U7963 (N_7963,N_4227,N_555);
nor U7964 (N_7964,N_3866,N_852);
and U7965 (N_7965,N_3526,N_292);
or U7966 (N_7966,N_1101,N_2169);
nor U7967 (N_7967,N_676,N_2898);
or U7968 (N_7968,N_3643,N_4837);
and U7969 (N_7969,N_272,N_4261);
and U7970 (N_7970,N_461,N_4429);
and U7971 (N_7971,N_562,N_395);
and U7972 (N_7972,N_3874,N_1059);
or U7973 (N_7973,N_23,N_823);
nor U7974 (N_7974,N_1207,N_1863);
nor U7975 (N_7975,N_2983,N_3827);
nand U7976 (N_7976,N_3937,N_3178);
and U7977 (N_7977,N_731,N_3622);
nand U7978 (N_7978,N_3916,N_4804);
nand U7979 (N_7979,N_4200,N_2699);
nor U7980 (N_7980,N_741,N_3887);
nor U7981 (N_7981,N_4110,N_4367);
or U7982 (N_7982,N_3502,N_1504);
and U7983 (N_7983,N_428,N_214);
nor U7984 (N_7984,N_4336,N_1482);
or U7985 (N_7985,N_2589,N_1977);
and U7986 (N_7986,N_4077,N_1334);
and U7987 (N_7987,N_1492,N_2060);
and U7988 (N_7988,N_3068,N_1319);
nor U7989 (N_7989,N_3279,N_4369);
and U7990 (N_7990,N_660,N_3812);
nor U7991 (N_7991,N_3165,N_4424);
nand U7992 (N_7992,N_4753,N_1571);
nor U7993 (N_7993,N_1043,N_853);
and U7994 (N_7994,N_4816,N_3543);
nor U7995 (N_7995,N_3339,N_4088);
nor U7996 (N_7996,N_1213,N_345);
or U7997 (N_7997,N_1600,N_1638);
nand U7998 (N_7998,N_3705,N_3956);
and U7999 (N_7999,N_2052,N_4218);
nand U8000 (N_8000,N_834,N_2113);
nand U8001 (N_8001,N_2126,N_4122);
and U8002 (N_8002,N_3865,N_4956);
and U8003 (N_8003,N_4664,N_228);
and U8004 (N_8004,N_1622,N_4082);
nand U8005 (N_8005,N_4844,N_68);
xor U8006 (N_8006,N_4108,N_66);
nand U8007 (N_8007,N_3488,N_758);
or U8008 (N_8008,N_3254,N_514);
nand U8009 (N_8009,N_1256,N_4478);
and U8010 (N_8010,N_3745,N_1996);
and U8011 (N_8011,N_3751,N_2687);
nand U8012 (N_8012,N_850,N_4134);
nor U8013 (N_8013,N_1477,N_968);
and U8014 (N_8014,N_4703,N_1012);
and U8015 (N_8015,N_4552,N_4309);
or U8016 (N_8016,N_3071,N_4452);
nand U8017 (N_8017,N_473,N_4497);
nand U8018 (N_8018,N_3402,N_2391);
nor U8019 (N_8019,N_324,N_1286);
nand U8020 (N_8020,N_4680,N_113);
nand U8021 (N_8021,N_1772,N_4260);
and U8022 (N_8022,N_388,N_3958);
nor U8023 (N_8023,N_4006,N_4186);
and U8024 (N_8024,N_4444,N_2027);
and U8025 (N_8025,N_4687,N_2652);
and U8026 (N_8026,N_70,N_663);
and U8027 (N_8027,N_4384,N_4393);
and U8028 (N_8028,N_1989,N_4810);
or U8029 (N_8029,N_3146,N_1014);
or U8030 (N_8030,N_3919,N_3647);
and U8031 (N_8031,N_1657,N_2635);
nand U8032 (N_8032,N_4172,N_2346);
nand U8033 (N_8033,N_2682,N_1427);
or U8034 (N_8034,N_936,N_804);
or U8035 (N_8035,N_2946,N_2951);
nand U8036 (N_8036,N_4954,N_2766);
and U8037 (N_8037,N_225,N_893);
nor U8038 (N_8038,N_4754,N_2731);
or U8039 (N_8039,N_121,N_607);
nor U8040 (N_8040,N_4878,N_3315);
nand U8041 (N_8041,N_3206,N_1853);
or U8042 (N_8042,N_4486,N_1640);
or U8043 (N_8043,N_4731,N_2607);
nor U8044 (N_8044,N_2380,N_2039);
and U8045 (N_8045,N_1941,N_927);
and U8046 (N_8046,N_4290,N_1039);
and U8047 (N_8047,N_4793,N_4553);
or U8048 (N_8048,N_1637,N_1757);
and U8049 (N_8049,N_683,N_1773);
or U8050 (N_8050,N_206,N_4766);
nand U8051 (N_8051,N_38,N_4749);
nor U8052 (N_8052,N_3805,N_3395);
nand U8053 (N_8053,N_4448,N_3759);
and U8054 (N_8054,N_300,N_4205);
and U8055 (N_8055,N_2744,N_4745);
or U8056 (N_8056,N_1657,N_3105);
nand U8057 (N_8057,N_2867,N_4394);
or U8058 (N_8058,N_3060,N_1589);
nand U8059 (N_8059,N_290,N_1);
and U8060 (N_8060,N_1842,N_4);
or U8061 (N_8061,N_4352,N_4368);
nor U8062 (N_8062,N_4330,N_1440);
and U8063 (N_8063,N_2946,N_4432);
and U8064 (N_8064,N_3678,N_4698);
and U8065 (N_8065,N_4532,N_4465);
and U8066 (N_8066,N_3256,N_143);
and U8067 (N_8067,N_4984,N_1578);
nor U8068 (N_8068,N_1904,N_901);
and U8069 (N_8069,N_3454,N_707);
nand U8070 (N_8070,N_692,N_2564);
and U8071 (N_8071,N_2496,N_3162);
nor U8072 (N_8072,N_1819,N_2972);
and U8073 (N_8073,N_2633,N_818);
nand U8074 (N_8074,N_3293,N_1213);
nand U8075 (N_8075,N_3687,N_448);
and U8076 (N_8076,N_4417,N_1621);
and U8077 (N_8077,N_542,N_963);
nor U8078 (N_8078,N_2052,N_4041);
nor U8079 (N_8079,N_194,N_43);
nor U8080 (N_8080,N_4965,N_4184);
and U8081 (N_8081,N_3477,N_3219);
nor U8082 (N_8082,N_2999,N_1176);
or U8083 (N_8083,N_515,N_702);
nor U8084 (N_8084,N_4311,N_4998);
and U8085 (N_8085,N_127,N_4534);
nand U8086 (N_8086,N_449,N_2419);
nand U8087 (N_8087,N_3639,N_4993);
nand U8088 (N_8088,N_1734,N_1797);
nand U8089 (N_8089,N_3327,N_2450);
nor U8090 (N_8090,N_4842,N_4541);
nor U8091 (N_8091,N_1267,N_2205);
or U8092 (N_8092,N_3238,N_2057);
or U8093 (N_8093,N_4128,N_598);
and U8094 (N_8094,N_2976,N_4889);
nor U8095 (N_8095,N_4196,N_4135);
or U8096 (N_8096,N_4316,N_4444);
nand U8097 (N_8097,N_4876,N_2592);
or U8098 (N_8098,N_4408,N_1048);
or U8099 (N_8099,N_1814,N_3807);
and U8100 (N_8100,N_4225,N_3355);
nand U8101 (N_8101,N_4213,N_1273);
nor U8102 (N_8102,N_4344,N_4941);
nand U8103 (N_8103,N_3371,N_1306);
nand U8104 (N_8104,N_2286,N_1589);
nand U8105 (N_8105,N_2210,N_1965);
nand U8106 (N_8106,N_1821,N_1962);
or U8107 (N_8107,N_2501,N_4705);
or U8108 (N_8108,N_1142,N_4613);
and U8109 (N_8109,N_1827,N_2350);
nand U8110 (N_8110,N_3430,N_1428);
nand U8111 (N_8111,N_4188,N_3218);
nor U8112 (N_8112,N_3250,N_2525);
nor U8113 (N_8113,N_2973,N_2344);
nand U8114 (N_8114,N_734,N_511);
nand U8115 (N_8115,N_2540,N_3345);
nand U8116 (N_8116,N_2687,N_1493);
nor U8117 (N_8117,N_3226,N_2942);
nand U8118 (N_8118,N_3077,N_2645);
nor U8119 (N_8119,N_4874,N_264);
or U8120 (N_8120,N_82,N_310);
nand U8121 (N_8121,N_2604,N_2997);
nand U8122 (N_8122,N_4153,N_2066);
and U8123 (N_8123,N_2768,N_3037);
nor U8124 (N_8124,N_1576,N_4823);
nor U8125 (N_8125,N_4514,N_1615);
xor U8126 (N_8126,N_4657,N_1324);
nand U8127 (N_8127,N_1022,N_2154);
or U8128 (N_8128,N_2422,N_4001);
nand U8129 (N_8129,N_1710,N_3249);
or U8130 (N_8130,N_3747,N_1173);
nor U8131 (N_8131,N_2572,N_911);
and U8132 (N_8132,N_3966,N_3526);
nor U8133 (N_8133,N_4177,N_4823);
and U8134 (N_8134,N_3311,N_3966);
nand U8135 (N_8135,N_2570,N_713);
nand U8136 (N_8136,N_1062,N_3796);
and U8137 (N_8137,N_2256,N_3705);
or U8138 (N_8138,N_2348,N_4955);
and U8139 (N_8139,N_1319,N_4350);
nand U8140 (N_8140,N_1989,N_1909);
nor U8141 (N_8141,N_4162,N_3392);
or U8142 (N_8142,N_3348,N_1931);
nor U8143 (N_8143,N_1874,N_288);
nor U8144 (N_8144,N_2534,N_2524);
or U8145 (N_8145,N_741,N_1235);
nand U8146 (N_8146,N_1917,N_1542);
and U8147 (N_8147,N_1386,N_2604);
nor U8148 (N_8148,N_1044,N_4264);
or U8149 (N_8149,N_2624,N_721);
nand U8150 (N_8150,N_1219,N_1641);
and U8151 (N_8151,N_2042,N_4292);
nor U8152 (N_8152,N_3602,N_1722);
or U8153 (N_8153,N_4219,N_1888);
and U8154 (N_8154,N_454,N_2915);
and U8155 (N_8155,N_240,N_2539);
nand U8156 (N_8156,N_1389,N_1213);
or U8157 (N_8157,N_145,N_2300);
nand U8158 (N_8158,N_3478,N_2315);
nand U8159 (N_8159,N_2403,N_4625);
or U8160 (N_8160,N_2422,N_2077);
and U8161 (N_8161,N_2422,N_4343);
xnor U8162 (N_8162,N_3518,N_1799);
and U8163 (N_8163,N_3585,N_1118);
nor U8164 (N_8164,N_3503,N_4683);
and U8165 (N_8165,N_559,N_3652);
nor U8166 (N_8166,N_3796,N_4339);
nand U8167 (N_8167,N_2766,N_3753);
or U8168 (N_8168,N_4117,N_2051);
nand U8169 (N_8169,N_2882,N_4223);
and U8170 (N_8170,N_1384,N_3792);
and U8171 (N_8171,N_2130,N_4880);
and U8172 (N_8172,N_2589,N_3145);
nand U8173 (N_8173,N_177,N_358);
and U8174 (N_8174,N_4674,N_2076);
nand U8175 (N_8175,N_1985,N_4857);
or U8176 (N_8176,N_1363,N_3919);
nand U8177 (N_8177,N_1956,N_4612);
or U8178 (N_8178,N_1423,N_4865);
or U8179 (N_8179,N_4352,N_189);
and U8180 (N_8180,N_4253,N_1964);
nor U8181 (N_8181,N_4938,N_36);
or U8182 (N_8182,N_2408,N_616);
nor U8183 (N_8183,N_3649,N_3398);
and U8184 (N_8184,N_3937,N_2310);
nor U8185 (N_8185,N_2001,N_2939);
nor U8186 (N_8186,N_787,N_3263);
or U8187 (N_8187,N_1260,N_580);
and U8188 (N_8188,N_2139,N_2254);
nor U8189 (N_8189,N_3975,N_1349);
nor U8190 (N_8190,N_189,N_217);
and U8191 (N_8191,N_3325,N_2357);
and U8192 (N_8192,N_4254,N_14);
and U8193 (N_8193,N_4216,N_4700);
nor U8194 (N_8194,N_2865,N_1161);
nand U8195 (N_8195,N_696,N_226);
nand U8196 (N_8196,N_3971,N_4365);
and U8197 (N_8197,N_26,N_591);
nand U8198 (N_8198,N_867,N_4065);
nand U8199 (N_8199,N_1752,N_1316);
or U8200 (N_8200,N_87,N_1231);
and U8201 (N_8201,N_3867,N_3180);
and U8202 (N_8202,N_892,N_4651);
nor U8203 (N_8203,N_355,N_1366);
nand U8204 (N_8204,N_4878,N_3894);
nand U8205 (N_8205,N_1118,N_2349);
nand U8206 (N_8206,N_3502,N_2458);
or U8207 (N_8207,N_3467,N_2198);
or U8208 (N_8208,N_24,N_2124);
or U8209 (N_8209,N_4313,N_2143);
or U8210 (N_8210,N_1141,N_295);
and U8211 (N_8211,N_1016,N_3825);
nor U8212 (N_8212,N_3336,N_1534);
nand U8213 (N_8213,N_3508,N_2552);
nor U8214 (N_8214,N_4630,N_231);
and U8215 (N_8215,N_330,N_3147);
nand U8216 (N_8216,N_4633,N_929);
or U8217 (N_8217,N_2340,N_3236);
nor U8218 (N_8218,N_4120,N_3963);
and U8219 (N_8219,N_3169,N_3492);
and U8220 (N_8220,N_1343,N_3291);
nand U8221 (N_8221,N_3542,N_2464);
or U8222 (N_8222,N_3860,N_4951);
nor U8223 (N_8223,N_4567,N_2938);
and U8224 (N_8224,N_3676,N_2149);
and U8225 (N_8225,N_467,N_1);
nand U8226 (N_8226,N_3601,N_94);
and U8227 (N_8227,N_3755,N_920);
or U8228 (N_8228,N_2651,N_3538);
and U8229 (N_8229,N_3017,N_3827);
nor U8230 (N_8230,N_1403,N_1450);
or U8231 (N_8231,N_125,N_3806);
nor U8232 (N_8232,N_1857,N_1693);
nor U8233 (N_8233,N_3357,N_3004);
nor U8234 (N_8234,N_4158,N_682);
nand U8235 (N_8235,N_2863,N_4580);
or U8236 (N_8236,N_1512,N_2080);
or U8237 (N_8237,N_2888,N_319);
and U8238 (N_8238,N_4638,N_2017);
or U8239 (N_8239,N_2314,N_4174);
or U8240 (N_8240,N_1378,N_933);
nor U8241 (N_8241,N_3272,N_606);
or U8242 (N_8242,N_3353,N_1712);
nor U8243 (N_8243,N_4513,N_371);
nand U8244 (N_8244,N_1690,N_4687);
or U8245 (N_8245,N_3913,N_2509);
or U8246 (N_8246,N_940,N_4470);
or U8247 (N_8247,N_301,N_2599);
and U8248 (N_8248,N_3440,N_1429);
nand U8249 (N_8249,N_3829,N_3499);
nor U8250 (N_8250,N_4148,N_2042);
nand U8251 (N_8251,N_4671,N_3051);
and U8252 (N_8252,N_532,N_3369);
or U8253 (N_8253,N_2502,N_930);
nand U8254 (N_8254,N_611,N_3025);
nor U8255 (N_8255,N_3841,N_2230);
and U8256 (N_8256,N_1766,N_4850);
nor U8257 (N_8257,N_3315,N_2033);
or U8258 (N_8258,N_1905,N_1774);
nor U8259 (N_8259,N_1689,N_2030);
and U8260 (N_8260,N_2155,N_4017);
or U8261 (N_8261,N_2891,N_4914);
nand U8262 (N_8262,N_598,N_99);
or U8263 (N_8263,N_1470,N_1099);
nor U8264 (N_8264,N_581,N_2957);
nand U8265 (N_8265,N_973,N_1317);
nand U8266 (N_8266,N_542,N_2664);
nor U8267 (N_8267,N_2296,N_2904);
nand U8268 (N_8268,N_1336,N_1994);
nand U8269 (N_8269,N_4341,N_489);
and U8270 (N_8270,N_550,N_3903);
nand U8271 (N_8271,N_2910,N_206);
or U8272 (N_8272,N_4270,N_3265);
and U8273 (N_8273,N_1022,N_1094);
nand U8274 (N_8274,N_1495,N_4245);
or U8275 (N_8275,N_1029,N_2507);
nand U8276 (N_8276,N_1333,N_2445);
nand U8277 (N_8277,N_2810,N_242);
nand U8278 (N_8278,N_3432,N_3911);
or U8279 (N_8279,N_840,N_33);
nor U8280 (N_8280,N_2714,N_789);
and U8281 (N_8281,N_4111,N_3719);
and U8282 (N_8282,N_4012,N_1686);
and U8283 (N_8283,N_4026,N_2227);
nand U8284 (N_8284,N_4498,N_178);
or U8285 (N_8285,N_2284,N_3365);
or U8286 (N_8286,N_4360,N_3388);
and U8287 (N_8287,N_259,N_3637);
xnor U8288 (N_8288,N_2137,N_3756);
nor U8289 (N_8289,N_3490,N_968);
or U8290 (N_8290,N_4238,N_1919);
and U8291 (N_8291,N_2981,N_2488);
nor U8292 (N_8292,N_1850,N_3107);
nor U8293 (N_8293,N_3957,N_3695);
nand U8294 (N_8294,N_445,N_2052);
nor U8295 (N_8295,N_2038,N_2797);
or U8296 (N_8296,N_3374,N_4451);
or U8297 (N_8297,N_1882,N_4338);
and U8298 (N_8298,N_3817,N_1598);
or U8299 (N_8299,N_2362,N_2399);
nand U8300 (N_8300,N_1322,N_463);
and U8301 (N_8301,N_4825,N_4205);
or U8302 (N_8302,N_3966,N_2604);
nand U8303 (N_8303,N_452,N_3508);
or U8304 (N_8304,N_1162,N_3462);
or U8305 (N_8305,N_486,N_3953);
nand U8306 (N_8306,N_2442,N_36);
and U8307 (N_8307,N_4020,N_3205);
or U8308 (N_8308,N_529,N_253);
nand U8309 (N_8309,N_597,N_2297);
nand U8310 (N_8310,N_3099,N_3017);
nand U8311 (N_8311,N_123,N_3179);
and U8312 (N_8312,N_4648,N_1676);
or U8313 (N_8313,N_1240,N_530);
nand U8314 (N_8314,N_1452,N_4452);
nor U8315 (N_8315,N_947,N_4845);
and U8316 (N_8316,N_4890,N_158);
or U8317 (N_8317,N_4403,N_1005);
and U8318 (N_8318,N_41,N_2701);
nand U8319 (N_8319,N_1030,N_787);
or U8320 (N_8320,N_4335,N_3993);
nor U8321 (N_8321,N_1936,N_2382);
nor U8322 (N_8322,N_1857,N_4719);
nor U8323 (N_8323,N_3935,N_1459);
and U8324 (N_8324,N_807,N_2053);
nor U8325 (N_8325,N_3632,N_2702);
or U8326 (N_8326,N_846,N_2385);
or U8327 (N_8327,N_648,N_3838);
and U8328 (N_8328,N_4488,N_3385);
nand U8329 (N_8329,N_2653,N_4559);
nand U8330 (N_8330,N_2943,N_1150);
nor U8331 (N_8331,N_3364,N_989);
nor U8332 (N_8332,N_2557,N_861);
and U8333 (N_8333,N_2143,N_3683);
nor U8334 (N_8334,N_3655,N_1297);
nand U8335 (N_8335,N_3470,N_1165);
or U8336 (N_8336,N_2028,N_207);
and U8337 (N_8337,N_564,N_4323);
nor U8338 (N_8338,N_1324,N_579);
nor U8339 (N_8339,N_203,N_263);
nor U8340 (N_8340,N_582,N_4001);
nand U8341 (N_8341,N_2030,N_4238);
nor U8342 (N_8342,N_4866,N_3831);
nor U8343 (N_8343,N_4735,N_1861);
or U8344 (N_8344,N_2314,N_2390);
and U8345 (N_8345,N_1608,N_4150);
nand U8346 (N_8346,N_2177,N_399);
and U8347 (N_8347,N_1813,N_2452);
nand U8348 (N_8348,N_1698,N_3069);
and U8349 (N_8349,N_2699,N_4014);
nand U8350 (N_8350,N_3030,N_633);
nand U8351 (N_8351,N_1859,N_2606);
or U8352 (N_8352,N_598,N_509);
or U8353 (N_8353,N_1070,N_1225);
nor U8354 (N_8354,N_3928,N_1829);
or U8355 (N_8355,N_2390,N_1652);
or U8356 (N_8356,N_1815,N_698);
nand U8357 (N_8357,N_2321,N_3739);
nand U8358 (N_8358,N_4912,N_4735);
nand U8359 (N_8359,N_4367,N_2113);
nand U8360 (N_8360,N_1856,N_3507);
nand U8361 (N_8361,N_1482,N_1377);
nand U8362 (N_8362,N_1964,N_1416);
nor U8363 (N_8363,N_205,N_2583);
nor U8364 (N_8364,N_3974,N_3783);
nand U8365 (N_8365,N_1105,N_3874);
nor U8366 (N_8366,N_2344,N_4952);
nor U8367 (N_8367,N_1255,N_4967);
and U8368 (N_8368,N_3793,N_1335);
nor U8369 (N_8369,N_1414,N_4609);
nand U8370 (N_8370,N_2512,N_4315);
nand U8371 (N_8371,N_678,N_1237);
nor U8372 (N_8372,N_2188,N_3469);
nor U8373 (N_8373,N_3967,N_1517);
and U8374 (N_8374,N_1927,N_2905);
nor U8375 (N_8375,N_4154,N_605);
or U8376 (N_8376,N_1542,N_2792);
and U8377 (N_8377,N_1244,N_4394);
nor U8378 (N_8378,N_1842,N_2052);
or U8379 (N_8379,N_289,N_3036);
or U8380 (N_8380,N_3444,N_2341);
nor U8381 (N_8381,N_3824,N_3731);
or U8382 (N_8382,N_1407,N_1434);
nor U8383 (N_8383,N_3859,N_4534);
or U8384 (N_8384,N_993,N_1595);
and U8385 (N_8385,N_1539,N_4724);
nor U8386 (N_8386,N_1997,N_1552);
or U8387 (N_8387,N_3975,N_1597);
nor U8388 (N_8388,N_4563,N_4196);
nand U8389 (N_8389,N_4675,N_3601);
nand U8390 (N_8390,N_4187,N_2969);
nor U8391 (N_8391,N_229,N_2983);
or U8392 (N_8392,N_3693,N_1264);
nand U8393 (N_8393,N_1407,N_4567);
and U8394 (N_8394,N_2984,N_1618);
and U8395 (N_8395,N_1654,N_1755);
and U8396 (N_8396,N_2320,N_776);
nand U8397 (N_8397,N_3435,N_3292);
or U8398 (N_8398,N_2744,N_1710);
and U8399 (N_8399,N_393,N_4573);
or U8400 (N_8400,N_2724,N_1466);
or U8401 (N_8401,N_2417,N_4455);
or U8402 (N_8402,N_728,N_3987);
nand U8403 (N_8403,N_1141,N_3081);
and U8404 (N_8404,N_1666,N_3751);
and U8405 (N_8405,N_474,N_4557);
nand U8406 (N_8406,N_2587,N_1181);
nand U8407 (N_8407,N_338,N_3671);
or U8408 (N_8408,N_629,N_4727);
and U8409 (N_8409,N_888,N_3889);
nand U8410 (N_8410,N_3977,N_1500);
nor U8411 (N_8411,N_2053,N_320);
nor U8412 (N_8412,N_1289,N_1508);
nor U8413 (N_8413,N_2303,N_784);
nand U8414 (N_8414,N_4116,N_3955);
and U8415 (N_8415,N_1048,N_637);
nand U8416 (N_8416,N_1770,N_3260);
or U8417 (N_8417,N_3973,N_1814);
and U8418 (N_8418,N_729,N_1470);
xor U8419 (N_8419,N_1481,N_712);
nor U8420 (N_8420,N_2811,N_1391);
or U8421 (N_8421,N_4403,N_283);
and U8422 (N_8422,N_2115,N_1970);
nand U8423 (N_8423,N_3705,N_2228);
or U8424 (N_8424,N_1922,N_4673);
or U8425 (N_8425,N_4598,N_2336);
or U8426 (N_8426,N_3628,N_3387);
nor U8427 (N_8427,N_154,N_1016);
nand U8428 (N_8428,N_2565,N_4182);
nor U8429 (N_8429,N_4385,N_2471);
or U8430 (N_8430,N_4163,N_664);
or U8431 (N_8431,N_3354,N_262);
and U8432 (N_8432,N_3642,N_3618);
nand U8433 (N_8433,N_1869,N_219);
and U8434 (N_8434,N_3433,N_3494);
and U8435 (N_8435,N_1535,N_3647);
nor U8436 (N_8436,N_910,N_3736);
nand U8437 (N_8437,N_3324,N_870);
or U8438 (N_8438,N_2419,N_1420);
nand U8439 (N_8439,N_1552,N_385);
and U8440 (N_8440,N_1732,N_84);
nor U8441 (N_8441,N_3131,N_3741);
nor U8442 (N_8442,N_3781,N_564);
nor U8443 (N_8443,N_3140,N_1480);
or U8444 (N_8444,N_2964,N_2768);
or U8445 (N_8445,N_1397,N_4584);
and U8446 (N_8446,N_2154,N_2459);
nand U8447 (N_8447,N_4917,N_2680);
nor U8448 (N_8448,N_2961,N_589);
and U8449 (N_8449,N_2777,N_2158);
nor U8450 (N_8450,N_2681,N_2335);
and U8451 (N_8451,N_1725,N_3570);
and U8452 (N_8452,N_3211,N_1280);
or U8453 (N_8453,N_2813,N_4619);
or U8454 (N_8454,N_3848,N_1160);
and U8455 (N_8455,N_1663,N_2109);
xor U8456 (N_8456,N_4994,N_1486);
and U8457 (N_8457,N_2286,N_2755);
and U8458 (N_8458,N_2417,N_4130);
nor U8459 (N_8459,N_3158,N_2504);
nand U8460 (N_8460,N_2434,N_1902);
and U8461 (N_8461,N_3488,N_917);
nor U8462 (N_8462,N_3011,N_1903);
or U8463 (N_8463,N_1732,N_3269);
and U8464 (N_8464,N_3306,N_4709);
and U8465 (N_8465,N_4812,N_84);
and U8466 (N_8466,N_715,N_2630);
and U8467 (N_8467,N_4405,N_225);
or U8468 (N_8468,N_2832,N_619);
or U8469 (N_8469,N_2841,N_768);
and U8470 (N_8470,N_4113,N_3299);
nor U8471 (N_8471,N_4984,N_1418);
and U8472 (N_8472,N_2551,N_742);
nand U8473 (N_8473,N_2637,N_3469);
nor U8474 (N_8474,N_2674,N_4512);
and U8475 (N_8475,N_1172,N_164);
nor U8476 (N_8476,N_3899,N_781);
nor U8477 (N_8477,N_581,N_2254);
nand U8478 (N_8478,N_3372,N_4554);
and U8479 (N_8479,N_3217,N_4223);
and U8480 (N_8480,N_2108,N_2827);
or U8481 (N_8481,N_611,N_4624);
or U8482 (N_8482,N_524,N_4710);
nand U8483 (N_8483,N_1448,N_2835);
and U8484 (N_8484,N_1189,N_423);
or U8485 (N_8485,N_4860,N_1078);
nand U8486 (N_8486,N_2386,N_4298);
or U8487 (N_8487,N_4112,N_249);
or U8488 (N_8488,N_1212,N_4077);
nand U8489 (N_8489,N_717,N_1069);
and U8490 (N_8490,N_3587,N_1452);
or U8491 (N_8491,N_4490,N_4819);
nor U8492 (N_8492,N_2249,N_4531);
or U8493 (N_8493,N_4626,N_4542);
nor U8494 (N_8494,N_3560,N_2470);
or U8495 (N_8495,N_1842,N_3841);
nor U8496 (N_8496,N_726,N_3607);
or U8497 (N_8497,N_734,N_1771);
nand U8498 (N_8498,N_2573,N_1801);
nand U8499 (N_8499,N_34,N_2602);
nor U8500 (N_8500,N_1044,N_3281);
or U8501 (N_8501,N_3640,N_109);
nand U8502 (N_8502,N_2124,N_115);
and U8503 (N_8503,N_3664,N_3329);
or U8504 (N_8504,N_704,N_3034);
nor U8505 (N_8505,N_2882,N_4677);
and U8506 (N_8506,N_1429,N_3446);
and U8507 (N_8507,N_2494,N_1899);
nor U8508 (N_8508,N_271,N_3404);
or U8509 (N_8509,N_2079,N_1085);
nand U8510 (N_8510,N_399,N_4229);
or U8511 (N_8511,N_194,N_119);
and U8512 (N_8512,N_1853,N_1671);
nor U8513 (N_8513,N_3366,N_3345);
nand U8514 (N_8514,N_3313,N_488);
and U8515 (N_8515,N_1261,N_1374);
nor U8516 (N_8516,N_1826,N_593);
or U8517 (N_8517,N_2386,N_839);
nor U8518 (N_8518,N_2362,N_1127);
or U8519 (N_8519,N_2945,N_92);
and U8520 (N_8520,N_4851,N_4700);
nor U8521 (N_8521,N_3533,N_1257);
nand U8522 (N_8522,N_1069,N_884);
or U8523 (N_8523,N_2468,N_1021);
or U8524 (N_8524,N_3458,N_1436);
and U8525 (N_8525,N_4839,N_4607);
or U8526 (N_8526,N_3218,N_1516);
and U8527 (N_8527,N_1112,N_3849);
or U8528 (N_8528,N_4795,N_1443);
nand U8529 (N_8529,N_1335,N_4423);
or U8530 (N_8530,N_16,N_1560);
nand U8531 (N_8531,N_3895,N_1337);
or U8532 (N_8532,N_445,N_3984);
nor U8533 (N_8533,N_1373,N_1004);
nor U8534 (N_8534,N_161,N_3750);
or U8535 (N_8535,N_4733,N_3719);
and U8536 (N_8536,N_1446,N_3729);
xnor U8537 (N_8537,N_3465,N_2935);
nor U8538 (N_8538,N_3583,N_968);
nand U8539 (N_8539,N_1441,N_3485);
and U8540 (N_8540,N_2412,N_1075);
nand U8541 (N_8541,N_391,N_2734);
nor U8542 (N_8542,N_1820,N_1822);
and U8543 (N_8543,N_918,N_2888);
nand U8544 (N_8544,N_4633,N_4923);
or U8545 (N_8545,N_2392,N_3942);
and U8546 (N_8546,N_1148,N_1567);
nand U8547 (N_8547,N_4612,N_4736);
nor U8548 (N_8548,N_1477,N_4672);
nand U8549 (N_8549,N_3055,N_2614);
or U8550 (N_8550,N_3388,N_4964);
and U8551 (N_8551,N_668,N_137);
and U8552 (N_8552,N_2955,N_3676);
nand U8553 (N_8553,N_4833,N_3778);
nor U8554 (N_8554,N_2270,N_4827);
and U8555 (N_8555,N_882,N_975);
nand U8556 (N_8556,N_2394,N_4099);
and U8557 (N_8557,N_1342,N_3590);
or U8558 (N_8558,N_1764,N_455);
nand U8559 (N_8559,N_4352,N_4302);
nand U8560 (N_8560,N_205,N_697);
or U8561 (N_8561,N_4653,N_356);
nand U8562 (N_8562,N_2773,N_3636);
or U8563 (N_8563,N_3330,N_2889);
and U8564 (N_8564,N_1540,N_1611);
and U8565 (N_8565,N_1924,N_1564);
nor U8566 (N_8566,N_4984,N_4372);
and U8567 (N_8567,N_880,N_2617);
or U8568 (N_8568,N_4007,N_3793);
or U8569 (N_8569,N_4994,N_3880);
and U8570 (N_8570,N_1198,N_2556);
or U8571 (N_8571,N_2314,N_3137);
nand U8572 (N_8572,N_4880,N_725);
or U8573 (N_8573,N_677,N_4319);
and U8574 (N_8574,N_1296,N_984);
and U8575 (N_8575,N_4904,N_2080);
and U8576 (N_8576,N_3328,N_2575);
and U8577 (N_8577,N_1626,N_1928);
and U8578 (N_8578,N_4596,N_4946);
or U8579 (N_8579,N_3211,N_843);
and U8580 (N_8580,N_4780,N_4785);
nand U8581 (N_8581,N_3726,N_2177);
and U8582 (N_8582,N_1840,N_431);
nand U8583 (N_8583,N_3458,N_4058);
nor U8584 (N_8584,N_358,N_991);
nor U8585 (N_8585,N_4624,N_4448);
nand U8586 (N_8586,N_156,N_3820);
nor U8587 (N_8587,N_2513,N_2354);
nor U8588 (N_8588,N_3701,N_1054);
and U8589 (N_8589,N_3082,N_41);
nand U8590 (N_8590,N_588,N_3553);
or U8591 (N_8591,N_2291,N_1773);
or U8592 (N_8592,N_2713,N_1531);
or U8593 (N_8593,N_2984,N_4299);
nand U8594 (N_8594,N_434,N_568);
or U8595 (N_8595,N_620,N_4722);
nor U8596 (N_8596,N_1136,N_354);
nor U8597 (N_8597,N_4454,N_2369);
and U8598 (N_8598,N_2636,N_2123);
nand U8599 (N_8599,N_1377,N_337);
and U8600 (N_8600,N_4751,N_3422);
nand U8601 (N_8601,N_1320,N_2350);
nand U8602 (N_8602,N_1955,N_611);
nor U8603 (N_8603,N_2579,N_1318);
and U8604 (N_8604,N_3179,N_632);
xor U8605 (N_8605,N_3313,N_2713);
or U8606 (N_8606,N_1848,N_2504);
and U8607 (N_8607,N_1030,N_4031);
or U8608 (N_8608,N_2980,N_2816);
nor U8609 (N_8609,N_4581,N_4355);
nand U8610 (N_8610,N_1141,N_2842);
xnor U8611 (N_8611,N_1199,N_2562);
nand U8612 (N_8612,N_1062,N_1758);
and U8613 (N_8613,N_4856,N_1150);
nand U8614 (N_8614,N_4252,N_985);
nor U8615 (N_8615,N_2423,N_34);
nor U8616 (N_8616,N_2422,N_1389);
and U8617 (N_8617,N_4478,N_2612);
and U8618 (N_8618,N_562,N_2935);
or U8619 (N_8619,N_224,N_983);
nor U8620 (N_8620,N_845,N_3395);
and U8621 (N_8621,N_4926,N_328);
nor U8622 (N_8622,N_2513,N_927);
nor U8623 (N_8623,N_1277,N_2394);
xnor U8624 (N_8624,N_584,N_2373);
or U8625 (N_8625,N_4534,N_116);
nor U8626 (N_8626,N_4201,N_65);
and U8627 (N_8627,N_4707,N_1699);
or U8628 (N_8628,N_4683,N_1874);
and U8629 (N_8629,N_2230,N_1656);
or U8630 (N_8630,N_2981,N_1457);
and U8631 (N_8631,N_803,N_7);
nor U8632 (N_8632,N_2600,N_1503);
and U8633 (N_8633,N_3944,N_1700);
nand U8634 (N_8634,N_4570,N_1488);
nand U8635 (N_8635,N_605,N_4292);
and U8636 (N_8636,N_332,N_896);
or U8637 (N_8637,N_880,N_854);
nor U8638 (N_8638,N_1415,N_2865);
nand U8639 (N_8639,N_338,N_2931);
and U8640 (N_8640,N_304,N_4509);
nor U8641 (N_8641,N_3654,N_1732);
and U8642 (N_8642,N_342,N_4496);
or U8643 (N_8643,N_3652,N_3672);
nor U8644 (N_8644,N_3769,N_4936);
nand U8645 (N_8645,N_2355,N_946);
nor U8646 (N_8646,N_4289,N_581);
or U8647 (N_8647,N_2253,N_1904);
nor U8648 (N_8648,N_4611,N_378);
and U8649 (N_8649,N_3911,N_196);
nand U8650 (N_8650,N_1038,N_3166);
nand U8651 (N_8651,N_1376,N_935);
or U8652 (N_8652,N_2471,N_4845);
or U8653 (N_8653,N_4570,N_2910);
nand U8654 (N_8654,N_3663,N_3151);
and U8655 (N_8655,N_367,N_1734);
and U8656 (N_8656,N_1336,N_3367);
nor U8657 (N_8657,N_2915,N_3948);
xor U8658 (N_8658,N_2329,N_3543);
or U8659 (N_8659,N_1315,N_1526);
nor U8660 (N_8660,N_3732,N_3000);
nor U8661 (N_8661,N_939,N_2042);
and U8662 (N_8662,N_222,N_464);
or U8663 (N_8663,N_3228,N_2187);
nand U8664 (N_8664,N_3352,N_682);
and U8665 (N_8665,N_2851,N_721);
nor U8666 (N_8666,N_4658,N_3285);
or U8667 (N_8667,N_3152,N_4886);
and U8668 (N_8668,N_4634,N_4530);
or U8669 (N_8669,N_78,N_2783);
and U8670 (N_8670,N_232,N_2624);
nand U8671 (N_8671,N_1246,N_2767);
and U8672 (N_8672,N_1843,N_4640);
or U8673 (N_8673,N_4683,N_1314);
nor U8674 (N_8674,N_2338,N_4771);
nor U8675 (N_8675,N_2518,N_1650);
nand U8676 (N_8676,N_3149,N_206);
nand U8677 (N_8677,N_1069,N_2924);
nand U8678 (N_8678,N_4273,N_440);
and U8679 (N_8679,N_4612,N_898);
nand U8680 (N_8680,N_4166,N_1333);
and U8681 (N_8681,N_4813,N_651);
xor U8682 (N_8682,N_2053,N_2104);
nand U8683 (N_8683,N_2889,N_2693);
nor U8684 (N_8684,N_51,N_1494);
nand U8685 (N_8685,N_3249,N_1733);
or U8686 (N_8686,N_520,N_19);
or U8687 (N_8687,N_1325,N_81);
nor U8688 (N_8688,N_4761,N_2258);
nor U8689 (N_8689,N_4967,N_4496);
nand U8690 (N_8690,N_2053,N_742);
nand U8691 (N_8691,N_3061,N_586);
nor U8692 (N_8692,N_137,N_3359);
nor U8693 (N_8693,N_928,N_1536);
and U8694 (N_8694,N_674,N_4406);
nor U8695 (N_8695,N_3267,N_906);
nor U8696 (N_8696,N_3992,N_2800);
or U8697 (N_8697,N_1562,N_3354);
and U8698 (N_8698,N_782,N_4091);
nand U8699 (N_8699,N_3324,N_4512);
and U8700 (N_8700,N_3566,N_893);
nor U8701 (N_8701,N_4085,N_4135);
nor U8702 (N_8702,N_3156,N_4885);
and U8703 (N_8703,N_503,N_1333);
or U8704 (N_8704,N_2825,N_1483);
nor U8705 (N_8705,N_4985,N_3043);
and U8706 (N_8706,N_3575,N_3450);
nand U8707 (N_8707,N_4662,N_2829);
and U8708 (N_8708,N_3060,N_683);
and U8709 (N_8709,N_4052,N_4631);
and U8710 (N_8710,N_1530,N_1386);
or U8711 (N_8711,N_2864,N_3423);
nor U8712 (N_8712,N_3209,N_3182);
and U8713 (N_8713,N_689,N_1103);
or U8714 (N_8714,N_753,N_318);
and U8715 (N_8715,N_949,N_1352);
or U8716 (N_8716,N_2354,N_4533);
nor U8717 (N_8717,N_3957,N_609);
or U8718 (N_8718,N_1789,N_2619);
or U8719 (N_8719,N_2069,N_3928);
nand U8720 (N_8720,N_172,N_3900);
nand U8721 (N_8721,N_3636,N_284);
nor U8722 (N_8722,N_1445,N_2657);
or U8723 (N_8723,N_1114,N_792);
nand U8724 (N_8724,N_4636,N_1561);
and U8725 (N_8725,N_1953,N_4504);
nor U8726 (N_8726,N_2853,N_263);
and U8727 (N_8727,N_1778,N_4546);
or U8728 (N_8728,N_2438,N_1454);
nand U8729 (N_8729,N_1776,N_3582);
and U8730 (N_8730,N_2593,N_3119);
or U8731 (N_8731,N_153,N_4320);
nor U8732 (N_8732,N_3184,N_3588);
nor U8733 (N_8733,N_2703,N_671);
or U8734 (N_8734,N_4019,N_3063);
nor U8735 (N_8735,N_892,N_686);
or U8736 (N_8736,N_2308,N_2771);
nand U8737 (N_8737,N_1790,N_3673);
nand U8738 (N_8738,N_1800,N_3982);
nand U8739 (N_8739,N_3632,N_1001);
nand U8740 (N_8740,N_3185,N_2006);
and U8741 (N_8741,N_3017,N_586);
nor U8742 (N_8742,N_3444,N_3433);
xnor U8743 (N_8743,N_3694,N_609);
and U8744 (N_8744,N_532,N_4408);
or U8745 (N_8745,N_4097,N_2388);
nand U8746 (N_8746,N_4752,N_1040);
nor U8747 (N_8747,N_1958,N_96);
nor U8748 (N_8748,N_2126,N_4983);
and U8749 (N_8749,N_4240,N_2836);
nor U8750 (N_8750,N_2892,N_779);
and U8751 (N_8751,N_3788,N_3339);
and U8752 (N_8752,N_1274,N_467);
and U8753 (N_8753,N_755,N_3537);
nand U8754 (N_8754,N_4526,N_833);
and U8755 (N_8755,N_3691,N_3171);
nand U8756 (N_8756,N_3924,N_1525);
nand U8757 (N_8757,N_3299,N_1323);
or U8758 (N_8758,N_1495,N_3813);
nand U8759 (N_8759,N_1374,N_741);
or U8760 (N_8760,N_2790,N_3435);
and U8761 (N_8761,N_9,N_1358);
nor U8762 (N_8762,N_3336,N_2936);
and U8763 (N_8763,N_2374,N_4626);
and U8764 (N_8764,N_1962,N_2242);
xnor U8765 (N_8765,N_3145,N_4649);
nand U8766 (N_8766,N_4376,N_1099);
and U8767 (N_8767,N_1073,N_3027);
nand U8768 (N_8768,N_4895,N_1287);
and U8769 (N_8769,N_2419,N_3493);
or U8770 (N_8770,N_4034,N_4904);
nand U8771 (N_8771,N_4304,N_2671);
and U8772 (N_8772,N_4396,N_710);
nor U8773 (N_8773,N_541,N_4522);
or U8774 (N_8774,N_4807,N_4956);
or U8775 (N_8775,N_2647,N_3995);
nor U8776 (N_8776,N_1401,N_3978);
nand U8777 (N_8777,N_4965,N_752);
nor U8778 (N_8778,N_1766,N_799);
and U8779 (N_8779,N_3111,N_281);
nand U8780 (N_8780,N_2353,N_299);
or U8781 (N_8781,N_771,N_4272);
nor U8782 (N_8782,N_19,N_4885);
nor U8783 (N_8783,N_188,N_3658);
nand U8784 (N_8784,N_2527,N_4168);
nor U8785 (N_8785,N_1629,N_3946);
or U8786 (N_8786,N_1591,N_2591);
and U8787 (N_8787,N_3536,N_4668);
and U8788 (N_8788,N_2905,N_4795);
or U8789 (N_8789,N_785,N_337);
nor U8790 (N_8790,N_1560,N_2911);
and U8791 (N_8791,N_111,N_4334);
and U8792 (N_8792,N_2648,N_256);
or U8793 (N_8793,N_604,N_2623);
nand U8794 (N_8794,N_2693,N_57);
and U8795 (N_8795,N_1868,N_4780);
nor U8796 (N_8796,N_1812,N_3301);
and U8797 (N_8797,N_504,N_4886);
or U8798 (N_8798,N_2425,N_1004);
and U8799 (N_8799,N_424,N_3772);
nor U8800 (N_8800,N_3338,N_4492);
nand U8801 (N_8801,N_2368,N_1455);
and U8802 (N_8802,N_932,N_4501);
nand U8803 (N_8803,N_2141,N_177);
and U8804 (N_8804,N_1881,N_2107);
nor U8805 (N_8805,N_1680,N_4767);
nor U8806 (N_8806,N_4850,N_778);
nor U8807 (N_8807,N_221,N_2218);
or U8808 (N_8808,N_0,N_2460);
nand U8809 (N_8809,N_4563,N_2349);
or U8810 (N_8810,N_4937,N_2133);
and U8811 (N_8811,N_2355,N_943);
nand U8812 (N_8812,N_4046,N_1078);
or U8813 (N_8813,N_37,N_3037);
nor U8814 (N_8814,N_4185,N_3362);
xor U8815 (N_8815,N_1496,N_1604);
nand U8816 (N_8816,N_3473,N_733);
and U8817 (N_8817,N_2691,N_2790);
or U8818 (N_8818,N_3920,N_1553);
and U8819 (N_8819,N_2217,N_4330);
or U8820 (N_8820,N_589,N_1831);
and U8821 (N_8821,N_1335,N_746);
nand U8822 (N_8822,N_2166,N_1822);
and U8823 (N_8823,N_3939,N_3817);
or U8824 (N_8824,N_310,N_1547);
or U8825 (N_8825,N_3775,N_1782);
nand U8826 (N_8826,N_2986,N_3497);
and U8827 (N_8827,N_4621,N_3742);
or U8828 (N_8828,N_3537,N_1053);
nand U8829 (N_8829,N_1735,N_467);
nand U8830 (N_8830,N_1115,N_4005);
nand U8831 (N_8831,N_2990,N_2226);
and U8832 (N_8832,N_2753,N_3192);
or U8833 (N_8833,N_4619,N_4779);
and U8834 (N_8834,N_3152,N_1825);
nor U8835 (N_8835,N_1167,N_3390);
nand U8836 (N_8836,N_4961,N_3976);
nor U8837 (N_8837,N_2956,N_4716);
and U8838 (N_8838,N_4786,N_1241);
nor U8839 (N_8839,N_709,N_1855);
nor U8840 (N_8840,N_2612,N_4329);
and U8841 (N_8841,N_1919,N_2494);
nor U8842 (N_8842,N_1192,N_1591);
and U8843 (N_8843,N_4254,N_4822);
or U8844 (N_8844,N_3961,N_803);
and U8845 (N_8845,N_1424,N_1616);
nor U8846 (N_8846,N_2856,N_2404);
nand U8847 (N_8847,N_1143,N_879);
nand U8848 (N_8848,N_3866,N_4144);
nor U8849 (N_8849,N_2952,N_3400);
or U8850 (N_8850,N_3004,N_3554);
and U8851 (N_8851,N_1627,N_463);
nor U8852 (N_8852,N_1190,N_3237);
nand U8853 (N_8853,N_3031,N_3824);
xor U8854 (N_8854,N_4222,N_962);
nor U8855 (N_8855,N_2380,N_1673);
or U8856 (N_8856,N_3947,N_1523);
nand U8857 (N_8857,N_3220,N_4859);
and U8858 (N_8858,N_2402,N_3416);
nand U8859 (N_8859,N_88,N_3120);
nor U8860 (N_8860,N_3669,N_3376);
and U8861 (N_8861,N_4943,N_2396);
or U8862 (N_8862,N_2481,N_1517);
nand U8863 (N_8863,N_4602,N_4590);
nor U8864 (N_8864,N_4432,N_4119);
or U8865 (N_8865,N_282,N_3932);
nor U8866 (N_8866,N_611,N_3098);
nand U8867 (N_8867,N_4849,N_266);
or U8868 (N_8868,N_3232,N_687);
nor U8869 (N_8869,N_4423,N_2843);
nor U8870 (N_8870,N_4965,N_3164);
and U8871 (N_8871,N_3495,N_3208);
nor U8872 (N_8872,N_3600,N_1992);
and U8873 (N_8873,N_1180,N_2294);
or U8874 (N_8874,N_3850,N_2423);
or U8875 (N_8875,N_2474,N_1239);
nor U8876 (N_8876,N_4076,N_1976);
or U8877 (N_8877,N_143,N_1904);
and U8878 (N_8878,N_2889,N_581);
nor U8879 (N_8879,N_636,N_463);
nor U8880 (N_8880,N_2160,N_4569);
or U8881 (N_8881,N_4866,N_950);
nand U8882 (N_8882,N_1946,N_2125);
nand U8883 (N_8883,N_2618,N_327);
nor U8884 (N_8884,N_2167,N_2842);
or U8885 (N_8885,N_995,N_2890);
or U8886 (N_8886,N_3239,N_310);
or U8887 (N_8887,N_2865,N_2049);
nor U8888 (N_8888,N_360,N_607);
nor U8889 (N_8889,N_2783,N_4788);
and U8890 (N_8890,N_4229,N_4396);
nor U8891 (N_8891,N_4331,N_4896);
nor U8892 (N_8892,N_1066,N_3355);
nor U8893 (N_8893,N_3337,N_1289);
or U8894 (N_8894,N_4019,N_3393);
nand U8895 (N_8895,N_1007,N_7);
nor U8896 (N_8896,N_4625,N_3437);
or U8897 (N_8897,N_2852,N_2993);
or U8898 (N_8898,N_710,N_1513);
nand U8899 (N_8899,N_3645,N_4276);
and U8900 (N_8900,N_3367,N_4684);
nand U8901 (N_8901,N_1502,N_4061);
and U8902 (N_8902,N_2390,N_4871);
and U8903 (N_8903,N_3348,N_2262);
nor U8904 (N_8904,N_3941,N_363);
xnor U8905 (N_8905,N_4751,N_187);
nand U8906 (N_8906,N_3255,N_3555);
and U8907 (N_8907,N_2278,N_1850);
nor U8908 (N_8908,N_2603,N_2628);
xnor U8909 (N_8909,N_2158,N_3238);
and U8910 (N_8910,N_3499,N_568);
nand U8911 (N_8911,N_2880,N_3316);
and U8912 (N_8912,N_2601,N_3237);
nand U8913 (N_8913,N_567,N_3410);
nand U8914 (N_8914,N_1778,N_1513);
nor U8915 (N_8915,N_4730,N_99);
nor U8916 (N_8916,N_151,N_1411);
and U8917 (N_8917,N_1825,N_2269);
and U8918 (N_8918,N_4995,N_2730);
or U8919 (N_8919,N_498,N_4898);
nor U8920 (N_8920,N_4597,N_805);
nand U8921 (N_8921,N_4622,N_2727);
or U8922 (N_8922,N_4942,N_3487);
nand U8923 (N_8923,N_1402,N_2653);
nand U8924 (N_8924,N_3585,N_3873);
and U8925 (N_8925,N_3514,N_3816);
nor U8926 (N_8926,N_1675,N_3182);
nand U8927 (N_8927,N_3427,N_278);
nand U8928 (N_8928,N_1263,N_1942);
nand U8929 (N_8929,N_4918,N_1366);
and U8930 (N_8930,N_2691,N_990);
nor U8931 (N_8931,N_3936,N_1865);
nand U8932 (N_8932,N_4688,N_2695);
xor U8933 (N_8933,N_3746,N_276);
nor U8934 (N_8934,N_4855,N_3567);
or U8935 (N_8935,N_2898,N_939);
and U8936 (N_8936,N_2076,N_324);
or U8937 (N_8937,N_4572,N_4251);
nor U8938 (N_8938,N_1832,N_36);
nand U8939 (N_8939,N_632,N_4080);
and U8940 (N_8940,N_2102,N_2697);
nor U8941 (N_8941,N_3688,N_703);
and U8942 (N_8942,N_3515,N_1674);
nand U8943 (N_8943,N_4886,N_145);
nor U8944 (N_8944,N_1547,N_1461);
and U8945 (N_8945,N_1404,N_3485);
nand U8946 (N_8946,N_1224,N_4644);
nand U8947 (N_8947,N_1395,N_2740);
nor U8948 (N_8948,N_2924,N_4972);
nand U8949 (N_8949,N_2245,N_1854);
or U8950 (N_8950,N_4896,N_3583);
and U8951 (N_8951,N_1368,N_837);
or U8952 (N_8952,N_1924,N_3756);
and U8953 (N_8953,N_4338,N_730);
xnor U8954 (N_8954,N_1268,N_1438);
or U8955 (N_8955,N_2476,N_3429);
nand U8956 (N_8956,N_3052,N_3187);
nor U8957 (N_8957,N_237,N_3092);
or U8958 (N_8958,N_1837,N_2574);
nor U8959 (N_8959,N_240,N_404);
nor U8960 (N_8960,N_667,N_4472);
nand U8961 (N_8961,N_3275,N_4544);
nand U8962 (N_8962,N_4712,N_2106);
or U8963 (N_8963,N_3713,N_4885);
nand U8964 (N_8964,N_396,N_4212);
nand U8965 (N_8965,N_4004,N_4370);
nor U8966 (N_8966,N_2569,N_993);
or U8967 (N_8967,N_789,N_2631);
or U8968 (N_8968,N_3905,N_2902);
nand U8969 (N_8969,N_1367,N_82);
nand U8970 (N_8970,N_4798,N_207);
nand U8971 (N_8971,N_2548,N_1557);
nand U8972 (N_8972,N_4624,N_1369);
nor U8973 (N_8973,N_3381,N_3596);
and U8974 (N_8974,N_1826,N_249);
and U8975 (N_8975,N_4833,N_4549);
and U8976 (N_8976,N_708,N_2742);
nor U8977 (N_8977,N_2494,N_1866);
or U8978 (N_8978,N_3294,N_2917);
and U8979 (N_8979,N_3236,N_1692);
or U8980 (N_8980,N_3582,N_3773);
or U8981 (N_8981,N_4656,N_3641);
nand U8982 (N_8982,N_1109,N_2489);
nand U8983 (N_8983,N_3864,N_733);
or U8984 (N_8984,N_2668,N_2947);
nor U8985 (N_8985,N_2632,N_1583);
nor U8986 (N_8986,N_921,N_1913);
or U8987 (N_8987,N_4169,N_1419);
nor U8988 (N_8988,N_379,N_775);
or U8989 (N_8989,N_2598,N_4537);
nor U8990 (N_8990,N_3689,N_3306);
nand U8991 (N_8991,N_1659,N_2400);
nand U8992 (N_8992,N_4530,N_4456);
nor U8993 (N_8993,N_4764,N_3963);
and U8994 (N_8994,N_1064,N_3005);
and U8995 (N_8995,N_519,N_2514);
nand U8996 (N_8996,N_2978,N_3112);
or U8997 (N_8997,N_2746,N_792);
and U8998 (N_8998,N_1289,N_3623);
nor U8999 (N_8999,N_2702,N_4774);
nor U9000 (N_9000,N_1461,N_1232);
or U9001 (N_9001,N_691,N_4109);
or U9002 (N_9002,N_1,N_2538);
nand U9003 (N_9003,N_1919,N_4256);
or U9004 (N_9004,N_420,N_3201);
or U9005 (N_9005,N_491,N_2750);
and U9006 (N_9006,N_1552,N_794);
or U9007 (N_9007,N_3819,N_1595);
and U9008 (N_9008,N_3733,N_2407);
or U9009 (N_9009,N_4508,N_4331);
nor U9010 (N_9010,N_3245,N_4147);
nor U9011 (N_9011,N_954,N_1767);
nand U9012 (N_9012,N_2438,N_3013);
or U9013 (N_9013,N_1498,N_2723);
or U9014 (N_9014,N_77,N_4139);
nor U9015 (N_9015,N_3625,N_4139);
nor U9016 (N_9016,N_75,N_2857);
nand U9017 (N_9017,N_4476,N_1892);
and U9018 (N_9018,N_2625,N_4604);
or U9019 (N_9019,N_1375,N_1436);
nor U9020 (N_9020,N_2938,N_4056);
nor U9021 (N_9021,N_3367,N_4394);
or U9022 (N_9022,N_2392,N_1814);
or U9023 (N_9023,N_602,N_3300);
nand U9024 (N_9024,N_4048,N_2275);
and U9025 (N_9025,N_2230,N_905);
nor U9026 (N_9026,N_384,N_1434);
nor U9027 (N_9027,N_323,N_1583);
nor U9028 (N_9028,N_1820,N_3611);
nor U9029 (N_9029,N_3106,N_58);
and U9030 (N_9030,N_918,N_1802);
and U9031 (N_9031,N_1305,N_539);
and U9032 (N_9032,N_1996,N_688);
or U9033 (N_9033,N_1255,N_2136);
or U9034 (N_9034,N_2230,N_4773);
or U9035 (N_9035,N_4870,N_1143);
or U9036 (N_9036,N_3509,N_4872);
or U9037 (N_9037,N_3682,N_4320);
or U9038 (N_9038,N_1381,N_4075);
nand U9039 (N_9039,N_3515,N_3641);
or U9040 (N_9040,N_1081,N_3371);
nand U9041 (N_9041,N_4087,N_4394);
nand U9042 (N_9042,N_1593,N_1764);
and U9043 (N_9043,N_801,N_2794);
nor U9044 (N_9044,N_20,N_3837);
and U9045 (N_9045,N_2716,N_2609);
and U9046 (N_9046,N_4798,N_3204);
or U9047 (N_9047,N_4569,N_2816);
and U9048 (N_9048,N_3779,N_347);
or U9049 (N_9049,N_2691,N_3160);
xor U9050 (N_9050,N_4844,N_2758);
nand U9051 (N_9051,N_868,N_1857);
and U9052 (N_9052,N_1422,N_1557);
nor U9053 (N_9053,N_2357,N_1434);
and U9054 (N_9054,N_453,N_2851);
and U9055 (N_9055,N_2066,N_4261);
nor U9056 (N_9056,N_4136,N_3317);
and U9057 (N_9057,N_1647,N_3323);
or U9058 (N_9058,N_232,N_4219);
nand U9059 (N_9059,N_806,N_2672);
nor U9060 (N_9060,N_1687,N_2833);
and U9061 (N_9061,N_1939,N_3862);
or U9062 (N_9062,N_1763,N_3919);
or U9063 (N_9063,N_4562,N_70);
nor U9064 (N_9064,N_1530,N_2602);
and U9065 (N_9065,N_936,N_1128);
and U9066 (N_9066,N_2714,N_4568);
nand U9067 (N_9067,N_1158,N_768);
nand U9068 (N_9068,N_2550,N_3145);
or U9069 (N_9069,N_1175,N_2700);
nor U9070 (N_9070,N_1511,N_2956);
nor U9071 (N_9071,N_3010,N_2636);
nor U9072 (N_9072,N_91,N_4888);
and U9073 (N_9073,N_153,N_961);
nor U9074 (N_9074,N_3224,N_1273);
or U9075 (N_9075,N_4802,N_2675);
or U9076 (N_9076,N_1426,N_2609);
and U9077 (N_9077,N_1476,N_1758);
nand U9078 (N_9078,N_4239,N_4924);
and U9079 (N_9079,N_2430,N_2116);
nand U9080 (N_9080,N_115,N_2915);
and U9081 (N_9081,N_4960,N_1681);
nor U9082 (N_9082,N_4840,N_2457);
or U9083 (N_9083,N_1809,N_3482);
and U9084 (N_9084,N_3753,N_4302);
and U9085 (N_9085,N_4725,N_4310);
and U9086 (N_9086,N_1950,N_1144);
and U9087 (N_9087,N_4403,N_3259);
and U9088 (N_9088,N_286,N_4992);
nor U9089 (N_9089,N_2489,N_1386);
nand U9090 (N_9090,N_236,N_87);
nand U9091 (N_9091,N_122,N_3469);
nor U9092 (N_9092,N_1098,N_2652);
and U9093 (N_9093,N_2872,N_3791);
nor U9094 (N_9094,N_841,N_2127);
nand U9095 (N_9095,N_2022,N_4876);
and U9096 (N_9096,N_3305,N_2341);
nor U9097 (N_9097,N_4901,N_2582);
or U9098 (N_9098,N_2057,N_1453);
nand U9099 (N_9099,N_1105,N_911);
and U9100 (N_9100,N_1888,N_3713);
or U9101 (N_9101,N_4975,N_3088);
and U9102 (N_9102,N_1801,N_1515);
nand U9103 (N_9103,N_4983,N_2875);
or U9104 (N_9104,N_2847,N_968);
or U9105 (N_9105,N_4617,N_4875);
or U9106 (N_9106,N_2353,N_4485);
or U9107 (N_9107,N_769,N_1957);
nor U9108 (N_9108,N_4519,N_2237);
nand U9109 (N_9109,N_3032,N_1229);
or U9110 (N_9110,N_3640,N_3388);
nor U9111 (N_9111,N_1139,N_4927);
and U9112 (N_9112,N_516,N_3087);
or U9113 (N_9113,N_3708,N_363);
nor U9114 (N_9114,N_4534,N_3148);
nor U9115 (N_9115,N_2842,N_1033);
nand U9116 (N_9116,N_3823,N_4143);
nand U9117 (N_9117,N_4408,N_4295);
or U9118 (N_9118,N_789,N_4694);
nor U9119 (N_9119,N_4434,N_4797);
nor U9120 (N_9120,N_377,N_3874);
and U9121 (N_9121,N_2052,N_1747);
nand U9122 (N_9122,N_4941,N_2050);
nor U9123 (N_9123,N_3436,N_4293);
nand U9124 (N_9124,N_3480,N_2728);
and U9125 (N_9125,N_4121,N_3760);
nor U9126 (N_9126,N_2957,N_2927);
or U9127 (N_9127,N_1609,N_4579);
nand U9128 (N_9128,N_820,N_2611);
nand U9129 (N_9129,N_1710,N_2315);
nand U9130 (N_9130,N_3587,N_1678);
or U9131 (N_9131,N_317,N_4845);
or U9132 (N_9132,N_1142,N_4243);
and U9133 (N_9133,N_4768,N_3774);
and U9134 (N_9134,N_2252,N_2895);
nor U9135 (N_9135,N_2325,N_1087);
and U9136 (N_9136,N_4765,N_4135);
and U9137 (N_9137,N_1461,N_90);
and U9138 (N_9138,N_1034,N_4189);
or U9139 (N_9139,N_4964,N_3488);
nor U9140 (N_9140,N_4983,N_465);
xor U9141 (N_9141,N_4906,N_4348);
nor U9142 (N_9142,N_1283,N_993);
nand U9143 (N_9143,N_442,N_2672);
nand U9144 (N_9144,N_572,N_2074);
and U9145 (N_9145,N_1132,N_2071);
nand U9146 (N_9146,N_1520,N_4791);
nor U9147 (N_9147,N_2219,N_3712);
or U9148 (N_9148,N_893,N_4016);
nor U9149 (N_9149,N_4941,N_3000);
nand U9150 (N_9150,N_991,N_1531);
or U9151 (N_9151,N_2489,N_3287);
and U9152 (N_9152,N_3889,N_230);
and U9153 (N_9153,N_3702,N_1200);
or U9154 (N_9154,N_2962,N_1366);
nand U9155 (N_9155,N_463,N_159);
and U9156 (N_9156,N_1555,N_1720);
nand U9157 (N_9157,N_2829,N_2480);
or U9158 (N_9158,N_3854,N_951);
nor U9159 (N_9159,N_3756,N_3902);
nand U9160 (N_9160,N_2605,N_1663);
nor U9161 (N_9161,N_3003,N_2160);
and U9162 (N_9162,N_3721,N_3498);
nor U9163 (N_9163,N_497,N_4344);
or U9164 (N_9164,N_3935,N_2584);
nand U9165 (N_9165,N_2145,N_2277);
and U9166 (N_9166,N_2537,N_2422);
or U9167 (N_9167,N_4677,N_2864);
or U9168 (N_9168,N_4669,N_3769);
or U9169 (N_9169,N_621,N_4794);
nor U9170 (N_9170,N_1986,N_3781);
nand U9171 (N_9171,N_3610,N_3472);
or U9172 (N_9172,N_4714,N_1009);
and U9173 (N_9173,N_4116,N_636);
or U9174 (N_9174,N_2162,N_4256);
or U9175 (N_9175,N_4118,N_826);
and U9176 (N_9176,N_2396,N_2405);
nor U9177 (N_9177,N_4898,N_4879);
and U9178 (N_9178,N_3389,N_1775);
nand U9179 (N_9179,N_625,N_3629);
nor U9180 (N_9180,N_1373,N_3835);
nand U9181 (N_9181,N_75,N_1974);
nand U9182 (N_9182,N_4195,N_2165);
nand U9183 (N_9183,N_3932,N_4514);
nand U9184 (N_9184,N_4016,N_1463);
and U9185 (N_9185,N_83,N_4148);
nand U9186 (N_9186,N_1696,N_300);
nor U9187 (N_9187,N_2134,N_4910);
or U9188 (N_9188,N_3659,N_3613);
nor U9189 (N_9189,N_322,N_606);
and U9190 (N_9190,N_678,N_1697);
nor U9191 (N_9191,N_1457,N_3511);
or U9192 (N_9192,N_810,N_3379);
nor U9193 (N_9193,N_3263,N_620);
or U9194 (N_9194,N_2513,N_1071);
nand U9195 (N_9195,N_912,N_3899);
nor U9196 (N_9196,N_3169,N_4286);
and U9197 (N_9197,N_4843,N_4767);
nor U9198 (N_9198,N_1293,N_4220);
and U9199 (N_9199,N_555,N_3965);
nor U9200 (N_9200,N_1814,N_4539);
and U9201 (N_9201,N_1824,N_81);
nor U9202 (N_9202,N_2061,N_2245);
or U9203 (N_9203,N_2020,N_4749);
and U9204 (N_9204,N_1567,N_2177);
and U9205 (N_9205,N_2666,N_3999);
and U9206 (N_9206,N_4392,N_2134);
nand U9207 (N_9207,N_20,N_4734);
nand U9208 (N_9208,N_497,N_658);
and U9209 (N_9209,N_3090,N_167);
or U9210 (N_9210,N_3263,N_4379);
nor U9211 (N_9211,N_1762,N_3373);
or U9212 (N_9212,N_328,N_1106);
nand U9213 (N_9213,N_2508,N_1525);
or U9214 (N_9214,N_3754,N_1523);
nand U9215 (N_9215,N_408,N_1878);
or U9216 (N_9216,N_4155,N_1896);
nand U9217 (N_9217,N_499,N_4933);
nor U9218 (N_9218,N_2272,N_4656);
or U9219 (N_9219,N_4550,N_1132);
and U9220 (N_9220,N_4375,N_1710);
and U9221 (N_9221,N_4494,N_1826);
nand U9222 (N_9222,N_467,N_3814);
nand U9223 (N_9223,N_4394,N_2930);
nand U9224 (N_9224,N_1938,N_2408);
or U9225 (N_9225,N_1880,N_2054);
nor U9226 (N_9226,N_3103,N_353);
nand U9227 (N_9227,N_675,N_1641);
or U9228 (N_9228,N_3449,N_295);
nor U9229 (N_9229,N_4797,N_4922);
or U9230 (N_9230,N_3361,N_2736);
or U9231 (N_9231,N_651,N_1975);
or U9232 (N_9232,N_2441,N_1395);
nand U9233 (N_9233,N_1462,N_4917);
nand U9234 (N_9234,N_1323,N_4481);
nor U9235 (N_9235,N_1415,N_717);
or U9236 (N_9236,N_3577,N_226);
or U9237 (N_9237,N_4587,N_1308);
or U9238 (N_9238,N_1157,N_3920);
and U9239 (N_9239,N_2584,N_3778);
nand U9240 (N_9240,N_2043,N_158);
nand U9241 (N_9241,N_1787,N_3183);
and U9242 (N_9242,N_3890,N_3262);
or U9243 (N_9243,N_3592,N_2890);
nand U9244 (N_9244,N_209,N_4640);
nand U9245 (N_9245,N_1674,N_3479);
nand U9246 (N_9246,N_3400,N_4885);
and U9247 (N_9247,N_116,N_4667);
or U9248 (N_9248,N_3899,N_4849);
or U9249 (N_9249,N_1382,N_739);
or U9250 (N_9250,N_1610,N_707);
or U9251 (N_9251,N_4343,N_994);
or U9252 (N_9252,N_1875,N_2700);
or U9253 (N_9253,N_583,N_839);
nand U9254 (N_9254,N_1261,N_1994);
and U9255 (N_9255,N_3841,N_4720);
and U9256 (N_9256,N_3576,N_1583);
and U9257 (N_9257,N_3064,N_2890);
or U9258 (N_9258,N_2630,N_274);
nor U9259 (N_9259,N_1218,N_224);
nor U9260 (N_9260,N_4028,N_913);
nor U9261 (N_9261,N_823,N_2392);
nand U9262 (N_9262,N_1946,N_3041);
nor U9263 (N_9263,N_3240,N_4618);
and U9264 (N_9264,N_3147,N_2670);
nand U9265 (N_9265,N_2036,N_978);
nand U9266 (N_9266,N_4435,N_1241);
and U9267 (N_9267,N_365,N_669);
or U9268 (N_9268,N_4694,N_2742);
nor U9269 (N_9269,N_3258,N_4187);
and U9270 (N_9270,N_3957,N_4799);
nand U9271 (N_9271,N_3932,N_2472);
and U9272 (N_9272,N_2187,N_4882);
and U9273 (N_9273,N_430,N_3679);
or U9274 (N_9274,N_4457,N_1502);
and U9275 (N_9275,N_3574,N_714);
xor U9276 (N_9276,N_1919,N_4352);
or U9277 (N_9277,N_319,N_2182);
and U9278 (N_9278,N_3912,N_218);
nor U9279 (N_9279,N_244,N_3875);
nor U9280 (N_9280,N_2018,N_3552);
and U9281 (N_9281,N_2709,N_1267);
nand U9282 (N_9282,N_4611,N_2964);
and U9283 (N_9283,N_1564,N_674);
or U9284 (N_9284,N_1956,N_4290);
nor U9285 (N_9285,N_3621,N_472);
nand U9286 (N_9286,N_4136,N_2632);
or U9287 (N_9287,N_1617,N_4415);
nor U9288 (N_9288,N_2479,N_95);
nand U9289 (N_9289,N_1759,N_4833);
or U9290 (N_9290,N_784,N_3023);
nand U9291 (N_9291,N_4126,N_3540);
nand U9292 (N_9292,N_1095,N_3244);
and U9293 (N_9293,N_3229,N_1172);
nor U9294 (N_9294,N_724,N_1259);
or U9295 (N_9295,N_1603,N_1823);
nor U9296 (N_9296,N_4442,N_2686);
nor U9297 (N_9297,N_515,N_2907);
or U9298 (N_9298,N_786,N_2925);
nand U9299 (N_9299,N_2896,N_2384);
or U9300 (N_9300,N_4640,N_3995);
nor U9301 (N_9301,N_3462,N_4759);
nand U9302 (N_9302,N_3858,N_3477);
nor U9303 (N_9303,N_2994,N_1367);
and U9304 (N_9304,N_3498,N_1798);
nor U9305 (N_9305,N_2007,N_1927);
nand U9306 (N_9306,N_3099,N_1863);
nand U9307 (N_9307,N_1336,N_2756);
nand U9308 (N_9308,N_3917,N_3044);
nand U9309 (N_9309,N_3684,N_2738);
or U9310 (N_9310,N_2946,N_1256);
nor U9311 (N_9311,N_1346,N_1539);
and U9312 (N_9312,N_1100,N_3432);
or U9313 (N_9313,N_2895,N_3801);
nand U9314 (N_9314,N_2281,N_3411);
and U9315 (N_9315,N_4854,N_1973);
nand U9316 (N_9316,N_4009,N_4563);
nand U9317 (N_9317,N_4034,N_4613);
and U9318 (N_9318,N_2291,N_3787);
and U9319 (N_9319,N_347,N_3069);
or U9320 (N_9320,N_510,N_1991);
or U9321 (N_9321,N_3087,N_72);
and U9322 (N_9322,N_4531,N_1045);
nand U9323 (N_9323,N_74,N_4959);
or U9324 (N_9324,N_2233,N_1059);
nor U9325 (N_9325,N_4087,N_1067);
and U9326 (N_9326,N_2524,N_130);
and U9327 (N_9327,N_3252,N_723);
nor U9328 (N_9328,N_821,N_4921);
xor U9329 (N_9329,N_3665,N_1209);
nor U9330 (N_9330,N_4268,N_3925);
nor U9331 (N_9331,N_288,N_381);
and U9332 (N_9332,N_3675,N_988);
nand U9333 (N_9333,N_492,N_2659);
nor U9334 (N_9334,N_2288,N_4867);
and U9335 (N_9335,N_4777,N_2967);
nor U9336 (N_9336,N_1783,N_763);
nor U9337 (N_9337,N_78,N_2554);
nor U9338 (N_9338,N_2382,N_4489);
or U9339 (N_9339,N_1864,N_1695);
nor U9340 (N_9340,N_1121,N_1825);
nor U9341 (N_9341,N_622,N_4726);
or U9342 (N_9342,N_638,N_1094);
nand U9343 (N_9343,N_3232,N_4899);
nor U9344 (N_9344,N_2196,N_82);
or U9345 (N_9345,N_2878,N_2177);
nor U9346 (N_9346,N_3904,N_2428);
nand U9347 (N_9347,N_317,N_1290);
nor U9348 (N_9348,N_2909,N_2934);
or U9349 (N_9349,N_787,N_2791);
nand U9350 (N_9350,N_4069,N_3674);
or U9351 (N_9351,N_4412,N_4210);
and U9352 (N_9352,N_1625,N_3123);
nand U9353 (N_9353,N_3793,N_4554);
nand U9354 (N_9354,N_3279,N_877);
nand U9355 (N_9355,N_3686,N_4710);
nor U9356 (N_9356,N_2763,N_3752);
nand U9357 (N_9357,N_4862,N_4119);
xnor U9358 (N_9358,N_3174,N_1065);
nand U9359 (N_9359,N_3371,N_4289);
and U9360 (N_9360,N_1977,N_3388);
nand U9361 (N_9361,N_3004,N_2178);
nand U9362 (N_9362,N_1344,N_1117);
nor U9363 (N_9363,N_1316,N_4293);
nand U9364 (N_9364,N_710,N_695);
nor U9365 (N_9365,N_4958,N_1514);
nor U9366 (N_9366,N_2464,N_1495);
nor U9367 (N_9367,N_3635,N_1809);
or U9368 (N_9368,N_1040,N_249);
or U9369 (N_9369,N_3554,N_569);
and U9370 (N_9370,N_3503,N_1731);
or U9371 (N_9371,N_3651,N_1230);
and U9372 (N_9372,N_1404,N_4510);
or U9373 (N_9373,N_1849,N_269);
and U9374 (N_9374,N_903,N_1012);
and U9375 (N_9375,N_4444,N_2934);
nand U9376 (N_9376,N_3308,N_2101);
or U9377 (N_9377,N_1509,N_4643);
nand U9378 (N_9378,N_1887,N_352);
and U9379 (N_9379,N_172,N_1338);
nand U9380 (N_9380,N_654,N_3941);
or U9381 (N_9381,N_2125,N_923);
or U9382 (N_9382,N_1058,N_637);
and U9383 (N_9383,N_2129,N_284);
nand U9384 (N_9384,N_638,N_3025);
or U9385 (N_9385,N_1052,N_1606);
nand U9386 (N_9386,N_2823,N_4549);
and U9387 (N_9387,N_4908,N_1740);
and U9388 (N_9388,N_2681,N_3116);
or U9389 (N_9389,N_1943,N_571);
nor U9390 (N_9390,N_2702,N_2638);
nand U9391 (N_9391,N_1979,N_951);
nor U9392 (N_9392,N_2856,N_4557);
nor U9393 (N_9393,N_4573,N_2402);
or U9394 (N_9394,N_660,N_2900);
nand U9395 (N_9395,N_3242,N_587);
or U9396 (N_9396,N_1084,N_1257);
and U9397 (N_9397,N_806,N_1496);
or U9398 (N_9398,N_662,N_4564);
or U9399 (N_9399,N_4964,N_3253);
nor U9400 (N_9400,N_4099,N_3103);
nand U9401 (N_9401,N_1102,N_1861);
or U9402 (N_9402,N_1543,N_2230);
nor U9403 (N_9403,N_97,N_3259);
or U9404 (N_9404,N_87,N_4478);
or U9405 (N_9405,N_4003,N_1320);
nor U9406 (N_9406,N_73,N_3629);
and U9407 (N_9407,N_4068,N_273);
nand U9408 (N_9408,N_2892,N_3215);
nand U9409 (N_9409,N_3797,N_4737);
or U9410 (N_9410,N_2187,N_3036);
nor U9411 (N_9411,N_594,N_3721);
nand U9412 (N_9412,N_1828,N_1899);
nand U9413 (N_9413,N_3250,N_4090);
and U9414 (N_9414,N_359,N_3135);
nor U9415 (N_9415,N_1538,N_1763);
and U9416 (N_9416,N_1198,N_2786);
xor U9417 (N_9417,N_4843,N_1660);
nand U9418 (N_9418,N_2740,N_1524);
and U9419 (N_9419,N_2883,N_2213);
nor U9420 (N_9420,N_1689,N_4132);
nor U9421 (N_9421,N_3142,N_4152);
nor U9422 (N_9422,N_2085,N_1477);
nor U9423 (N_9423,N_4388,N_2271);
nor U9424 (N_9424,N_1599,N_3902);
or U9425 (N_9425,N_528,N_4168);
or U9426 (N_9426,N_2417,N_4074);
nor U9427 (N_9427,N_661,N_1624);
nor U9428 (N_9428,N_2506,N_1735);
nor U9429 (N_9429,N_177,N_113);
nor U9430 (N_9430,N_3549,N_567);
nor U9431 (N_9431,N_1903,N_4902);
nor U9432 (N_9432,N_1268,N_1315);
and U9433 (N_9433,N_3781,N_2735);
or U9434 (N_9434,N_4116,N_1380);
and U9435 (N_9435,N_4140,N_4453);
and U9436 (N_9436,N_2042,N_4830);
nand U9437 (N_9437,N_2083,N_4883);
nand U9438 (N_9438,N_3867,N_4448);
or U9439 (N_9439,N_2554,N_1744);
nand U9440 (N_9440,N_1594,N_4643);
and U9441 (N_9441,N_2427,N_4498);
nor U9442 (N_9442,N_3843,N_791);
and U9443 (N_9443,N_4254,N_1965);
or U9444 (N_9444,N_2492,N_1829);
nor U9445 (N_9445,N_4134,N_4192);
and U9446 (N_9446,N_2601,N_4098);
or U9447 (N_9447,N_733,N_1106);
and U9448 (N_9448,N_4864,N_3090);
nor U9449 (N_9449,N_4668,N_1831);
nor U9450 (N_9450,N_4405,N_380);
or U9451 (N_9451,N_2359,N_4122);
and U9452 (N_9452,N_3727,N_463);
nor U9453 (N_9453,N_1805,N_138);
nand U9454 (N_9454,N_2262,N_2632);
nand U9455 (N_9455,N_4863,N_1524);
and U9456 (N_9456,N_2053,N_2563);
or U9457 (N_9457,N_3601,N_1693);
and U9458 (N_9458,N_4871,N_1725);
nor U9459 (N_9459,N_3709,N_2255);
or U9460 (N_9460,N_4374,N_4651);
or U9461 (N_9461,N_2786,N_4303);
or U9462 (N_9462,N_226,N_1607);
nor U9463 (N_9463,N_747,N_3471);
or U9464 (N_9464,N_551,N_1631);
nor U9465 (N_9465,N_2023,N_3972);
or U9466 (N_9466,N_4958,N_2083);
nor U9467 (N_9467,N_512,N_1163);
or U9468 (N_9468,N_4708,N_4125);
nand U9469 (N_9469,N_381,N_1500);
and U9470 (N_9470,N_1661,N_4225);
nor U9471 (N_9471,N_576,N_2752);
or U9472 (N_9472,N_3305,N_233);
and U9473 (N_9473,N_2562,N_2397);
nor U9474 (N_9474,N_438,N_2231);
and U9475 (N_9475,N_2070,N_2862);
nand U9476 (N_9476,N_1476,N_387);
and U9477 (N_9477,N_1497,N_1873);
and U9478 (N_9478,N_2295,N_1969);
nor U9479 (N_9479,N_3751,N_84);
nor U9480 (N_9480,N_1596,N_3563);
nor U9481 (N_9481,N_4033,N_569);
or U9482 (N_9482,N_3701,N_1653);
and U9483 (N_9483,N_1663,N_1269);
nand U9484 (N_9484,N_2658,N_3363);
and U9485 (N_9485,N_4252,N_2036);
nand U9486 (N_9486,N_3757,N_3277);
nand U9487 (N_9487,N_393,N_2554);
nand U9488 (N_9488,N_4377,N_1494);
and U9489 (N_9489,N_3722,N_2602);
or U9490 (N_9490,N_4591,N_3078);
nand U9491 (N_9491,N_2997,N_4842);
nor U9492 (N_9492,N_330,N_3464);
and U9493 (N_9493,N_2444,N_3395);
or U9494 (N_9494,N_2237,N_1635);
and U9495 (N_9495,N_4914,N_1339);
nand U9496 (N_9496,N_3921,N_953);
and U9497 (N_9497,N_2074,N_3850);
or U9498 (N_9498,N_1206,N_1717);
nor U9499 (N_9499,N_872,N_123);
nor U9500 (N_9500,N_1752,N_719);
and U9501 (N_9501,N_2580,N_2280);
nor U9502 (N_9502,N_2972,N_2169);
or U9503 (N_9503,N_1754,N_892);
or U9504 (N_9504,N_1540,N_3850);
or U9505 (N_9505,N_4541,N_3070);
nor U9506 (N_9506,N_4735,N_2276);
nor U9507 (N_9507,N_2885,N_4323);
and U9508 (N_9508,N_1223,N_941);
and U9509 (N_9509,N_4088,N_2263);
and U9510 (N_9510,N_4854,N_1472);
or U9511 (N_9511,N_4754,N_4265);
xnor U9512 (N_9512,N_1753,N_3011);
or U9513 (N_9513,N_812,N_3482);
nand U9514 (N_9514,N_2980,N_4899);
or U9515 (N_9515,N_3504,N_48);
or U9516 (N_9516,N_2203,N_2848);
nand U9517 (N_9517,N_4248,N_1129);
nand U9518 (N_9518,N_2438,N_1457);
nand U9519 (N_9519,N_1225,N_4395);
nor U9520 (N_9520,N_809,N_2496);
nand U9521 (N_9521,N_1867,N_1965);
or U9522 (N_9522,N_3554,N_2830);
or U9523 (N_9523,N_691,N_248);
or U9524 (N_9524,N_1870,N_631);
and U9525 (N_9525,N_3578,N_1845);
nor U9526 (N_9526,N_3706,N_356);
or U9527 (N_9527,N_137,N_3516);
nand U9528 (N_9528,N_3398,N_2523);
and U9529 (N_9529,N_428,N_794);
and U9530 (N_9530,N_39,N_2658);
nor U9531 (N_9531,N_555,N_3715);
nand U9532 (N_9532,N_798,N_1230);
and U9533 (N_9533,N_4260,N_2437);
or U9534 (N_9534,N_4169,N_2555);
or U9535 (N_9535,N_1162,N_1064);
or U9536 (N_9536,N_112,N_232);
and U9537 (N_9537,N_1708,N_1908);
and U9538 (N_9538,N_1029,N_3828);
and U9539 (N_9539,N_2684,N_2640);
and U9540 (N_9540,N_530,N_1051);
nor U9541 (N_9541,N_3806,N_226);
nor U9542 (N_9542,N_2815,N_79);
nor U9543 (N_9543,N_935,N_1482);
and U9544 (N_9544,N_2030,N_793);
and U9545 (N_9545,N_3892,N_2925);
or U9546 (N_9546,N_4710,N_6);
nor U9547 (N_9547,N_1553,N_466);
or U9548 (N_9548,N_3136,N_2292);
nor U9549 (N_9549,N_3127,N_1807);
nor U9550 (N_9550,N_4954,N_4765);
and U9551 (N_9551,N_2463,N_1477);
nor U9552 (N_9552,N_2512,N_3224);
nand U9553 (N_9553,N_391,N_4604);
and U9554 (N_9554,N_4095,N_917);
nand U9555 (N_9555,N_1103,N_4211);
xor U9556 (N_9556,N_1668,N_3966);
or U9557 (N_9557,N_125,N_4863);
nor U9558 (N_9558,N_3678,N_1021);
nor U9559 (N_9559,N_1099,N_2543);
or U9560 (N_9560,N_2825,N_313);
xnor U9561 (N_9561,N_3533,N_283);
nand U9562 (N_9562,N_995,N_4498);
and U9563 (N_9563,N_1958,N_2414);
or U9564 (N_9564,N_3332,N_4636);
nor U9565 (N_9565,N_3598,N_575);
or U9566 (N_9566,N_2246,N_3298);
and U9567 (N_9567,N_1754,N_2024);
nor U9568 (N_9568,N_1295,N_3057);
nand U9569 (N_9569,N_4964,N_335);
or U9570 (N_9570,N_4774,N_4914);
or U9571 (N_9571,N_2188,N_4327);
and U9572 (N_9572,N_3495,N_54);
and U9573 (N_9573,N_2345,N_4130);
or U9574 (N_9574,N_3042,N_2431);
nor U9575 (N_9575,N_1213,N_1266);
nor U9576 (N_9576,N_3400,N_579);
and U9577 (N_9577,N_4662,N_4393);
nor U9578 (N_9578,N_1893,N_4698);
or U9579 (N_9579,N_1722,N_1023);
and U9580 (N_9580,N_176,N_286);
and U9581 (N_9581,N_2002,N_2092);
and U9582 (N_9582,N_4419,N_2305);
nor U9583 (N_9583,N_4007,N_3084);
nand U9584 (N_9584,N_1075,N_1078);
nand U9585 (N_9585,N_62,N_4538);
nor U9586 (N_9586,N_1793,N_2339);
and U9587 (N_9587,N_3213,N_3400);
and U9588 (N_9588,N_2423,N_1358);
or U9589 (N_9589,N_4160,N_2264);
nand U9590 (N_9590,N_4009,N_1305);
and U9591 (N_9591,N_3586,N_4593);
nand U9592 (N_9592,N_1376,N_406);
and U9593 (N_9593,N_4685,N_851);
nand U9594 (N_9594,N_2482,N_2884);
or U9595 (N_9595,N_495,N_4229);
nand U9596 (N_9596,N_3114,N_4099);
nor U9597 (N_9597,N_949,N_1684);
and U9598 (N_9598,N_3479,N_986);
nand U9599 (N_9599,N_289,N_2368);
nand U9600 (N_9600,N_2656,N_3803);
or U9601 (N_9601,N_1206,N_1301);
and U9602 (N_9602,N_116,N_1307);
and U9603 (N_9603,N_1841,N_2023);
nand U9604 (N_9604,N_3700,N_2451);
and U9605 (N_9605,N_4444,N_3793);
or U9606 (N_9606,N_3790,N_3583);
nand U9607 (N_9607,N_4853,N_4239);
or U9608 (N_9608,N_264,N_3877);
and U9609 (N_9609,N_121,N_742);
nor U9610 (N_9610,N_74,N_2017);
nor U9611 (N_9611,N_1492,N_1530);
and U9612 (N_9612,N_4627,N_4827);
nand U9613 (N_9613,N_3683,N_343);
nor U9614 (N_9614,N_4259,N_569);
nor U9615 (N_9615,N_1864,N_3731);
nor U9616 (N_9616,N_2036,N_1255);
or U9617 (N_9617,N_457,N_1942);
and U9618 (N_9618,N_1419,N_3829);
nand U9619 (N_9619,N_1413,N_1498);
and U9620 (N_9620,N_4148,N_1473);
or U9621 (N_9621,N_2165,N_642);
nand U9622 (N_9622,N_3125,N_2769);
and U9623 (N_9623,N_2964,N_4485);
nor U9624 (N_9624,N_77,N_2777);
nand U9625 (N_9625,N_3317,N_1997);
nand U9626 (N_9626,N_977,N_1151);
and U9627 (N_9627,N_4538,N_369);
xor U9628 (N_9628,N_2687,N_4728);
nor U9629 (N_9629,N_1093,N_1448);
nor U9630 (N_9630,N_371,N_4547);
or U9631 (N_9631,N_2959,N_4359);
and U9632 (N_9632,N_720,N_1568);
and U9633 (N_9633,N_4776,N_514);
nand U9634 (N_9634,N_451,N_2052);
or U9635 (N_9635,N_2798,N_576);
and U9636 (N_9636,N_3296,N_60);
nand U9637 (N_9637,N_173,N_3998);
nor U9638 (N_9638,N_3675,N_3538);
and U9639 (N_9639,N_2945,N_91);
or U9640 (N_9640,N_2053,N_181);
or U9641 (N_9641,N_4309,N_1545);
or U9642 (N_9642,N_256,N_3123);
nand U9643 (N_9643,N_4701,N_1953);
nor U9644 (N_9644,N_2234,N_998);
and U9645 (N_9645,N_4921,N_919);
nor U9646 (N_9646,N_2398,N_3064);
and U9647 (N_9647,N_2222,N_4985);
and U9648 (N_9648,N_1893,N_2272);
nor U9649 (N_9649,N_134,N_4963);
nand U9650 (N_9650,N_3919,N_1890);
nor U9651 (N_9651,N_3939,N_2056);
nand U9652 (N_9652,N_1128,N_2182);
or U9653 (N_9653,N_255,N_4134);
nand U9654 (N_9654,N_2371,N_2979);
xnor U9655 (N_9655,N_2498,N_2038);
nor U9656 (N_9656,N_2915,N_2978);
and U9657 (N_9657,N_2906,N_4674);
or U9658 (N_9658,N_2070,N_3767);
nand U9659 (N_9659,N_2689,N_3705);
nor U9660 (N_9660,N_4878,N_1950);
and U9661 (N_9661,N_3018,N_4760);
nor U9662 (N_9662,N_2661,N_4635);
nor U9663 (N_9663,N_1354,N_3909);
and U9664 (N_9664,N_1004,N_2468);
nor U9665 (N_9665,N_2767,N_541);
nand U9666 (N_9666,N_3326,N_1538);
nand U9667 (N_9667,N_22,N_238);
nor U9668 (N_9668,N_4489,N_828);
or U9669 (N_9669,N_4430,N_3294);
or U9670 (N_9670,N_1763,N_4523);
nand U9671 (N_9671,N_2294,N_3608);
nand U9672 (N_9672,N_3455,N_3581);
or U9673 (N_9673,N_708,N_3206);
nor U9674 (N_9674,N_3828,N_2219);
nand U9675 (N_9675,N_371,N_845);
and U9676 (N_9676,N_1549,N_3816);
nor U9677 (N_9677,N_525,N_2775);
and U9678 (N_9678,N_521,N_4322);
nor U9679 (N_9679,N_1863,N_4231);
or U9680 (N_9680,N_4517,N_741);
xor U9681 (N_9681,N_1644,N_4681);
and U9682 (N_9682,N_1324,N_417);
and U9683 (N_9683,N_1829,N_3667);
and U9684 (N_9684,N_1200,N_42);
and U9685 (N_9685,N_4880,N_3869);
and U9686 (N_9686,N_4166,N_3807);
nand U9687 (N_9687,N_2623,N_4981);
nor U9688 (N_9688,N_2453,N_2823);
or U9689 (N_9689,N_3621,N_2374);
nor U9690 (N_9690,N_4111,N_4062);
and U9691 (N_9691,N_3759,N_1834);
and U9692 (N_9692,N_384,N_3686);
or U9693 (N_9693,N_1376,N_3778);
or U9694 (N_9694,N_1543,N_3153);
or U9695 (N_9695,N_482,N_197);
nand U9696 (N_9696,N_3275,N_4836);
and U9697 (N_9697,N_1692,N_76);
nand U9698 (N_9698,N_2713,N_4778);
and U9699 (N_9699,N_3787,N_1605);
or U9700 (N_9700,N_1276,N_4705);
and U9701 (N_9701,N_513,N_4445);
nand U9702 (N_9702,N_666,N_1890);
nand U9703 (N_9703,N_201,N_132);
and U9704 (N_9704,N_3112,N_4895);
nand U9705 (N_9705,N_3015,N_3457);
and U9706 (N_9706,N_4378,N_20);
or U9707 (N_9707,N_1097,N_1231);
nor U9708 (N_9708,N_1003,N_2643);
and U9709 (N_9709,N_3513,N_1848);
nor U9710 (N_9710,N_3789,N_4385);
nor U9711 (N_9711,N_24,N_1612);
or U9712 (N_9712,N_1380,N_2085);
nor U9713 (N_9713,N_3768,N_3844);
nand U9714 (N_9714,N_1929,N_1846);
nand U9715 (N_9715,N_4423,N_3645);
nand U9716 (N_9716,N_2681,N_3950);
nand U9717 (N_9717,N_819,N_4209);
or U9718 (N_9718,N_1743,N_1855);
or U9719 (N_9719,N_257,N_3290);
nor U9720 (N_9720,N_4953,N_2437);
nand U9721 (N_9721,N_3051,N_3480);
nand U9722 (N_9722,N_1611,N_3946);
nand U9723 (N_9723,N_2321,N_3075);
nand U9724 (N_9724,N_3823,N_2080);
and U9725 (N_9725,N_2537,N_100);
nand U9726 (N_9726,N_41,N_4680);
or U9727 (N_9727,N_2168,N_3918);
or U9728 (N_9728,N_1430,N_4887);
nor U9729 (N_9729,N_571,N_3478);
or U9730 (N_9730,N_810,N_3768);
nor U9731 (N_9731,N_3590,N_2931);
nand U9732 (N_9732,N_3153,N_4051);
nor U9733 (N_9733,N_3159,N_904);
or U9734 (N_9734,N_14,N_1305);
or U9735 (N_9735,N_4319,N_4724);
nor U9736 (N_9736,N_150,N_4356);
nand U9737 (N_9737,N_1215,N_785);
and U9738 (N_9738,N_1009,N_2598);
nand U9739 (N_9739,N_4035,N_985);
nand U9740 (N_9740,N_4308,N_231);
and U9741 (N_9741,N_825,N_4754);
nand U9742 (N_9742,N_531,N_1689);
and U9743 (N_9743,N_252,N_1730);
nand U9744 (N_9744,N_888,N_3853);
nor U9745 (N_9745,N_4964,N_1902);
nor U9746 (N_9746,N_3580,N_2163);
and U9747 (N_9747,N_1428,N_3412);
nor U9748 (N_9748,N_230,N_1717);
nor U9749 (N_9749,N_3733,N_2759);
nor U9750 (N_9750,N_4358,N_3377);
nor U9751 (N_9751,N_758,N_2535);
nor U9752 (N_9752,N_902,N_2625);
or U9753 (N_9753,N_1893,N_1542);
or U9754 (N_9754,N_2038,N_4114);
or U9755 (N_9755,N_1843,N_2280);
and U9756 (N_9756,N_21,N_281);
nor U9757 (N_9757,N_3782,N_344);
or U9758 (N_9758,N_3017,N_401);
or U9759 (N_9759,N_4456,N_4526);
or U9760 (N_9760,N_4149,N_346);
nand U9761 (N_9761,N_3219,N_51);
nor U9762 (N_9762,N_904,N_3507);
and U9763 (N_9763,N_50,N_4287);
or U9764 (N_9764,N_4049,N_1884);
and U9765 (N_9765,N_1815,N_3244);
and U9766 (N_9766,N_590,N_2653);
nor U9767 (N_9767,N_785,N_4642);
xor U9768 (N_9768,N_215,N_802);
or U9769 (N_9769,N_1123,N_1931);
or U9770 (N_9770,N_3580,N_3690);
nor U9771 (N_9771,N_2740,N_1978);
or U9772 (N_9772,N_3319,N_798);
nor U9773 (N_9773,N_626,N_2256);
or U9774 (N_9774,N_4020,N_4186);
nor U9775 (N_9775,N_3667,N_1146);
nand U9776 (N_9776,N_4784,N_4470);
nand U9777 (N_9777,N_2369,N_3968);
nand U9778 (N_9778,N_4508,N_4156);
nand U9779 (N_9779,N_291,N_2445);
or U9780 (N_9780,N_3827,N_1562);
nand U9781 (N_9781,N_2514,N_2925);
and U9782 (N_9782,N_2685,N_3884);
and U9783 (N_9783,N_2834,N_980);
nand U9784 (N_9784,N_3062,N_4966);
or U9785 (N_9785,N_989,N_557);
or U9786 (N_9786,N_3625,N_3492);
nor U9787 (N_9787,N_3823,N_263);
nor U9788 (N_9788,N_3434,N_2034);
nand U9789 (N_9789,N_3203,N_4395);
nor U9790 (N_9790,N_3457,N_579);
nand U9791 (N_9791,N_880,N_694);
and U9792 (N_9792,N_1285,N_2477);
and U9793 (N_9793,N_2790,N_4524);
and U9794 (N_9794,N_1573,N_4395);
and U9795 (N_9795,N_4951,N_493);
nand U9796 (N_9796,N_1850,N_2805);
or U9797 (N_9797,N_767,N_3503);
and U9798 (N_9798,N_49,N_1747);
or U9799 (N_9799,N_1268,N_794);
nand U9800 (N_9800,N_2009,N_3305);
nand U9801 (N_9801,N_803,N_3058);
nor U9802 (N_9802,N_4757,N_295);
or U9803 (N_9803,N_697,N_4011);
and U9804 (N_9804,N_992,N_1699);
nor U9805 (N_9805,N_1613,N_2027);
nor U9806 (N_9806,N_4943,N_3769);
or U9807 (N_9807,N_3471,N_1224);
and U9808 (N_9808,N_1785,N_1600);
nor U9809 (N_9809,N_2064,N_3361);
and U9810 (N_9810,N_626,N_2394);
and U9811 (N_9811,N_3082,N_725);
nor U9812 (N_9812,N_195,N_1685);
and U9813 (N_9813,N_2765,N_3663);
and U9814 (N_9814,N_433,N_3347);
nor U9815 (N_9815,N_2556,N_3542);
nor U9816 (N_9816,N_4789,N_549);
xor U9817 (N_9817,N_3499,N_1308);
nor U9818 (N_9818,N_4219,N_2632);
nand U9819 (N_9819,N_847,N_470);
nand U9820 (N_9820,N_606,N_33);
or U9821 (N_9821,N_2897,N_4784);
and U9822 (N_9822,N_711,N_4862);
or U9823 (N_9823,N_2230,N_1740);
nand U9824 (N_9824,N_2292,N_243);
and U9825 (N_9825,N_543,N_2357);
nor U9826 (N_9826,N_4150,N_2566);
or U9827 (N_9827,N_397,N_2276);
nand U9828 (N_9828,N_1602,N_1563);
and U9829 (N_9829,N_3323,N_2487);
nor U9830 (N_9830,N_4968,N_4907);
and U9831 (N_9831,N_4144,N_4946);
nand U9832 (N_9832,N_70,N_3308);
nand U9833 (N_9833,N_3204,N_4858);
xor U9834 (N_9834,N_2691,N_2322);
or U9835 (N_9835,N_301,N_2530);
nor U9836 (N_9836,N_845,N_1689);
and U9837 (N_9837,N_3712,N_2830);
or U9838 (N_9838,N_2966,N_825);
and U9839 (N_9839,N_4412,N_4719);
nand U9840 (N_9840,N_4378,N_1923);
and U9841 (N_9841,N_3271,N_4577);
or U9842 (N_9842,N_2816,N_4884);
or U9843 (N_9843,N_1941,N_3943);
xnor U9844 (N_9844,N_2943,N_3476);
xnor U9845 (N_9845,N_1192,N_1932);
or U9846 (N_9846,N_3794,N_853);
nor U9847 (N_9847,N_1261,N_3284);
or U9848 (N_9848,N_4736,N_480);
or U9849 (N_9849,N_1180,N_966);
or U9850 (N_9850,N_697,N_4372);
and U9851 (N_9851,N_1464,N_4818);
or U9852 (N_9852,N_4000,N_3531);
or U9853 (N_9853,N_1392,N_124);
or U9854 (N_9854,N_4259,N_3405);
and U9855 (N_9855,N_931,N_1570);
and U9856 (N_9856,N_2991,N_2760);
or U9857 (N_9857,N_1234,N_4423);
nand U9858 (N_9858,N_2157,N_2471);
nor U9859 (N_9859,N_3308,N_4630);
or U9860 (N_9860,N_2537,N_4322);
and U9861 (N_9861,N_577,N_623);
nand U9862 (N_9862,N_4636,N_2595);
nand U9863 (N_9863,N_4245,N_4736);
xnor U9864 (N_9864,N_4116,N_1573);
nor U9865 (N_9865,N_1484,N_1129);
or U9866 (N_9866,N_4307,N_1857);
or U9867 (N_9867,N_2648,N_2863);
nor U9868 (N_9868,N_1090,N_4565);
nand U9869 (N_9869,N_4766,N_1200);
nand U9870 (N_9870,N_4213,N_200);
nand U9871 (N_9871,N_3505,N_4892);
nand U9872 (N_9872,N_1573,N_135);
nor U9873 (N_9873,N_3016,N_4665);
nand U9874 (N_9874,N_1153,N_1595);
or U9875 (N_9875,N_2492,N_560);
nand U9876 (N_9876,N_2166,N_4881);
nor U9877 (N_9877,N_4812,N_4591);
nand U9878 (N_9878,N_3508,N_3196);
nand U9879 (N_9879,N_4129,N_3548);
nand U9880 (N_9880,N_3686,N_2784);
or U9881 (N_9881,N_158,N_4385);
nor U9882 (N_9882,N_982,N_2930);
or U9883 (N_9883,N_4086,N_2586);
or U9884 (N_9884,N_2325,N_23);
nor U9885 (N_9885,N_3375,N_3446);
and U9886 (N_9886,N_935,N_3091);
or U9887 (N_9887,N_4659,N_1584);
and U9888 (N_9888,N_4446,N_3527);
and U9889 (N_9889,N_748,N_2498);
and U9890 (N_9890,N_211,N_4092);
xor U9891 (N_9891,N_2595,N_3207);
or U9892 (N_9892,N_648,N_1519);
or U9893 (N_9893,N_3743,N_300);
and U9894 (N_9894,N_100,N_4108);
nor U9895 (N_9895,N_271,N_1891);
and U9896 (N_9896,N_1785,N_262);
or U9897 (N_9897,N_3764,N_4110);
nor U9898 (N_9898,N_2224,N_1482);
and U9899 (N_9899,N_2173,N_3479);
or U9900 (N_9900,N_4226,N_4726);
or U9901 (N_9901,N_3397,N_425);
or U9902 (N_9902,N_1061,N_3721);
nand U9903 (N_9903,N_3599,N_158);
nor U9904 (N_9904,N_2463,N_1870);
or U9905 (N_9905,N_4726,N_582);
nor U9906 (N_9906,N_1277,N_227);
or U9907 (N_9907,N_4950,N_3842);
or U9908 (N_9908,N_450,N_975);
nand U9909 (N_9909,N_753,N_4213);
or U9910 (N_9910,N_1004,N_2590);
or U9911 (N_9911,N_1002,N_4320);
or U9912 (N_9912,N_1641,N_2302);
nor U9913 (N_9913,N_1501,N_2482);
nor U9914 (N_9914,N_2674,N_1226);
and U9915 (N_9915,N_3573,N_4776);
nand U9916 (N_9916,N_1060,N_2726);
nand U9917 (N_9917,N_2385,N_2225);
nor U9918 (N_9918,N_3911,N_74);
xor U9919 (N_9919,N_4020,N_1626);
and U9920 (N_9920,N_2868,N_1241);
and U9921 (N_9921,N_4191,N_864);
nor U9922 (N_9922,N_3705,N_2104);
nand U9923 (N_9923,N_2374,N_4448);
nand U9924 (N_9924,N_2735,N_2695);
xor U9925 (N_9925,N_3997,N_1650);
nor U9926 (N_9926,N_1168,N_1095);
or U9927 (N_9927,N_4073,N_3952);
or U9928 (N_9928,N_4454,N_1807);
nor U9929 (N_9929,N_3669,N_4651);
nand U9930 (N_9930,N_4566,N_1607);
or U9931 (N_9931,N_3625,N_1664);
nor U9932 (N_9932,N_4807,N_4628);
and U9933 (N_9933,N_3137,N_3803);
nor U9934 (N_9934,N_1630,N_4333);
nand U9935 (N_9935,N_3889,N_1172);
or U9936 (N_9936,N_979,N_1070);
nand U9937 (N_9937,N_803,N_1648);
nor U9938 (N_9938,N_1961,N_2894);
or U9939 (N_9939,N_2205,N_3788);
or U9940 (N_9940,N_1573,N_2325);
xnor U9941 (N_9941,N_2525,N_1771);
nor U9942 (N_9942,N_3428,N_4181);
nand U9943 (N_9943,N_698,N_4796);
or U9944 (N_9944,N_257,N_2763);
and U9945 (N_9945,N_1807,N_3537);
and U9946 (N_9946,N_3918,N_716);
and U9947 (N_9947,N_540,N_853);
and U9948 (N_9948,N_1230,N_4994);
xor U9949 (N_9949,N_260,N_1432);
nor U9950 (N_9950,N_716,N_2586);
nand U9951 (N_9951,N_4500,N_2828);
nand U9952 (N_9952,N_2648,N_3174);
and U9953 (N_9953,N_4042,N_1166);
or U9954 (N_9954,N_1708,N_2406);
nor U9955 (N_9955,N_1827,N_4468);
or U9956 (N_9956,N_4905,N_4709);
nand U9957 (N_9957,N_2133,N_689);
and U9958 (N_9958,N_1910,N_2059);
and U9959 (N_9959,N_638,N_1063);
nand U9960 (N_9960,N_2550,N_3539);
nor U9961 (N_9961,N_3538,N_3912);
and U9962 (N_9962,N_3517,N_212);
nor U9963 (N_9963,N_3368,N_299);
nand U9964 (N_9964,N_2034,N_4625);
and U9965 (N_9965,N_2945,N_2456);
nor U9966 (N_9966,N_4192,N_1015);
and U9967 (N_9967,N_2854,N_2280);
or U9968 (N_9968,N_4953,N_126);
or U9969 (N_9969,N_334,N_3915);
nand U9970 (N_9970,N_2394,N_4421);
and U9971 (N_9971,N_750,N_3956);
or U9972 (N_9972,N_2917,N_4897);
nand U9973 (N_9973,N_1331,N_1207);
nand U9974 (N_9974,N_3010,N_946);
nor U9975 (N_9975,N_3232,N_730);
or U9976 (N_9976,N_1498,N_1011);
or U9977 (N_9977,N_375,N_2974);
nand U9978 (N_9978,N_494,N_832);
or U9979 (N_9979,N_4916,N_1958);
or U9980 (N_9980,N_3234,N_1727);
nand U9981 (N_9981,N_181,N_4895);
nor U9982 (N_9982,N_502,N_1952);
or U9983 (N_9983,N_3714,N_1845);
nand U9984 (N_9984,N_2823,N_4151);
or U9985 (N_9985,N_3551,N_1329);
or U9986 (N_9986,N_4732,N_3584);
or U9987 (N_9987,N_1482,N_1570);
or U9988 (N_9988,N_940,N_2285);
nand U9989 (N_9989,N_1660,N_3320);
nand U9990 (N_9990,N_3288,N_1894);
nor U9991 (N_9991,N_3962,N_1696);
and U9992 (N_9992,N_2161,N_1474);
nor U9993 (N_9993,N_4020,N_1795);
or U9994 (N_9994,N_2800,N_4110);
or U9995 (N_9995,N_3454,N_963);
nor U9996 (N_9996,N_413,N_1420);
or U9997 (N_9997,N_4090,N_2709);
and U9998 (N_9998,N_4258,N_1502);
xnor U9999 (N_9999,N_2578,N_3587);
and UO_0 (O_0,N_7309,N_9845);
or UO_1 (O_1,N_6183,N_9142);
nand UO_2 (O_2,N_5558,N_7695);
nor UO_3 (O_3,N_7175,N_9097);
or UO_4 (O_4,N_9315,N_9925);
nor UO_5 (O_5,N_7582,N_5698);
or UO_6 (O_6,N_7438,N_5522);
or UO_7 (O_7,N_8842,N_5668);
nor UO_8 (O_8,N_5954,N_6749);
nand UO_9 (O_9,N_5692,N_7296);
nand UO_10 (O_10,N_9150,N_6496);
nor UO_11 (O_11,N_9206,N_7214);
and UO_12 (O_12,N_5133,N_8803);
nor UO_13 (O_13,N_9641,N_8782);
or UO_14 (O_14,N_9589,N_5766);
or UO_15 (O_15,N_5422,N_7389);
nand UO_16 (O_16,N_7152,N_8183);
and UO_17 (O_17,N_7629,N_5852);
and UO_18 (O_18,N_9327,N_7996);
or UO_19 (O_19,N_5441,N_7725);
or UO_20 (O_20,N_7418,N_7074);
or UO_21 (O_21,N_6083,N_7312);
and UO_22 (O_22,N_6740,N_7326);
or UO_23 (O_23,N_6484,N_5138);
nand UO_24 (O_24,N_5278,N_6337);
nor UO_25 (O_25,N_5065,N_6011);
and UO_26 (O_26,N_9603,N_7843);
nor UO_27 (O_27,N_9779,N_6179);
and UO_28 (O_28,N_5232,N_6344);
nand UO_29 (O_29,N_7627,N_6043);
or UO_30 (O_30,N_5959,N_5417);
and UO_31 (O_31,N_7887,N_8736);
nand UO_32 (O_32,N_8438,N_6644);
nor UO_33 (O_33,N_7058,N_9463);
nor UO_34 (O_34,N_5564,N_8668);
or UO_35 (O_35,N_9165,N_8332);
nand UO_36 (O_36,N_8885,N_5219);
nand UO_37 (O_37,N_7940,N_7886);
and UO_38 (O_38,N_6068,N_7789);
or UO_39 (O_39,N_5205,N_7170);
or UO_40 (O_40,N_9352,N_6826);
nand UO_41 (O_41,N_5448,N_5914);
nor UO_42 (O_42,N_7426,N_7733);
nand UO_43 (O_43,N_5689,N_8952);
xor UO_44 (O_44,N_6023,N_5270);
or UO_45 (O_45,N_5351,N_8994);
nor UO_46 (O_46,N_6797,N_9990);
nand UO_47 (O_47,N_9303,N_8236);
nor UO_48 (O_48,N_6794,N_7933);
nor UO_49 (O_49,N_7363,N_7604);
and UO_50 (O_50,N_6709,N_8533);
nand UO_51 (O_51,N_9083,N_7117);
nand UO_52 (O_52,N_6902,N_8433);
xor UO_53 (O_53,N_9469,N_8238);
or UO_54 (O_54,N_6099,N_7970);
nor UO_55 (O_55,N_6110,N_7249);
nor UO_56 (O_56,N_9955,N_5454);
nor UO_57 (O_57,N_6837,N_5934);
or UO_58 (O_58,N_5268,N_6795);
and UO_59 (O_59,N_7470,N_6674);
nand UO_60 (O_60,N_7535,N_8463);
nand UO_61 (O_61,N_7145,N_9601);
or UO_62 (O_62,N_5674,N_7279);
and UO_63 (O_63,N_6578,N_5030);
and UO_64 (O_64,N_7476,N_9489);
and UO_65 (O_65,N_9975,N_5924);
nand UO_66 (O_66,N_9154,N_8748);
or UO_67 (O_67,N_6014,N_6132);
and UO_68 (O_68,N_5590,N_9542);
nand UO_69 (O_69,N_9284,N_7376);
and UO_70 (O_70,N_6671,N_8865);
nand UO_71 (O_71,N_5817,N_5895);
nor UO_72 (O_72,N_5007,N_8930);
or UO_73 (O_73,N_9400,N_8279);
nor UO_74 (O_74,N_5166,N_9246);
nand UO_75 (O_75,N_7202,N_6333);
or UO_76 (O_76,N_9385,N_5555);
and UO_77 (O_77,N_7223,N_8143);
nor UO_78 (O_78,N_6645,N_6200);
nand UO_79 (O_79,N_8794,N_6154);
or UO_80 (O_80,N_8811,N_6699);
nor UO_81 (O_81,N_9379,N_9768);
or UO_82 (O_82,N_5778,N_6045);
or UO_83 (O_83,N_8773,N_8336);
nor UO_84 (O_84,N_7751,N_9293);
and UO_85 (O_85,N_7248,N_6426);
nand UO_86 (O_86,N_6760,N_6691);
nor UO_87 (O_87,N_6577,N_6679);
nand UO_88 (O_88,N_9449,N_6391);
or UO_89 (O_89,N_9612,N_7514);
nor UO_90 (O_90,N_5032,N_6159);
or UO_91 (O_91,N_8593,N_7678);
nor UO_92 (O_92,N_7115,N_7784);
and UO_93 (O_93,N_7599,N_6713);
nand UO_94 (O_94,N_7664,N_5231);
nand UO_95 (O_95,N_9608,N_7100);
or UO_96 (O_96,N_7052,N_9319);
nor UO_97 (O_97,N_9045,N_5458);
nand UO_98 (O_98,N_8379,N_8979);
nand UO_99 (O_99,N_8455,N_9010);
nor UO_100 (O_100,N_9640,N_6726);
nor UO_101 (O_101,N_8339,N_7464);
and UO_102 (O_102,N_7301,N_8522);
and UO_103 (O_103,N_6448,N_5662);
nand UO_104 (O_104,N_8389,N_8701);
nand UO_105 (O_105,N_8771,N_6685);
and UO_106 (O_106,N_9733,N_6285);
or UO_107 (O_107,N_5480,N_8967);
nor UO_108 (O_108,N_8318,N_7203);
and UO_109 (O_109,N_6584,N_8902);
and UO_110 (O_110,N_8933,N_7785);
and UO_111 (O_111,N_9860,N_9967);
or UO_112 (O_112,N_9238,N_8059);
or UO_113 (O_113,N_5896,N_7496);
and UO_114 (O_114,N_6234,N_9981);
nor UO_115 (O_115,N_6602,N_8664);
or UO_116 (O_116,N_5712,N_6474);
nor UO_117 (O_117,N_8950,N_7455);
or UO_118 (O_118,N_8937,N_8819);
or UO_119 (O_119,N_5728,N_9953);
or UO_120 (O_120,N_9487,N_9310);
or UO_121 (O_121,N_9633,N_5220);
nand UO_122 (O_122,N_8047,N_8833);
nand UO_123 (O_123,N_8008,N_7701);
nor UO_124 (O_124,N_5946,N_9921);
nor UO_125 (O_125,N_6847,N_5251);
nand UO_126 (O_126,N_8739,N_6239);
nand UO_127 (O_127,N_6279,N_6431);
nor UO_128 (O_128,N_6737,N_6956);
nor UO_129 (O_129,N_9059,N_9948);
or UO_130 (O_130,N_8978,N_8619);
nor UO_131 (O_131,N_8537,N_8239);
nor UO_132 (O_132,N_8767,N_5247);
or UO_133 (O_133,N_8982,N_9203);
or UO_134 (O_134,N_6774,N_5572);
and UO_135 (O_135,N_9875,N_5354);
or UO_136 (O_136,N_8275,N_9823);
or UO_137 (O_137,N_7798,N_6326);
and UO_138 (O_138,N_6890,N_8689);
nand UO_139 (O_139,N_8620,N_8523);
and UO_140 (O_140,N_5675,N_5071);
nor UO_141 (O_141,N_9596,N_6753);
nand UO_142 (O_142,N_7821,N_8812);
nor UO_143 (O_143,N_6813,N_9757);
or UO_144 (O_144,N_6966,N_9357);
or UO_145 (O_145,N_6944,N_8650);
nand UO_146 (O_146,N_5253,N_5989);
nor UO_147 (O_147,N_7349,N_8906);
nand UO_148 (O_148,N_6204,N_9676);
xnor UO_149 (O_149,N_6127,N_6784);
nand UO_150 (O_150,N_5210,N_6149);
nand UO_151 (O_151,N_9871,N_8569);
and UO_152 (O_152,N_6403,N_9978);
xnor UO_153 (O_153,N_5055,N_7261);
nand UO_154 (O_154,N_6913,N_7596);
nor UO_155 (O_155,N_9190,N_6935);
and UO_156 (O_156,N_8372,N_9917);
nand UO_157 (O_157,N_9015,N_8805);
nor UO_158 (O_158,N_8185,N_6485);
and UO_159 (O_159,N_8447,N_8639);
nor UO_160 (O_160,N_5443,N_7792);
and UO_161 (O_161,N_5399,N_5579);
and UO_162 (O_162,N_7558,N_9996);
nor UO_163 (O_163,N_6963,N_8205);
and UO_164 (O_164,N_6152,N_6687);
nor UO_165 (O_165,N_8016,N_8211);
nand UO_166 (O_166,N_6829,N_6102);
nor UO_167 (O_167,N_7468,N_6503);
and UO_168 (O_168,N_6938,N_9699);
or UO_169 (O_169,N_9139,N_9202);
and UO_170 (O_170,N_7027,N_5949);
nor UO_171 (O_171,N_6056,N_7055);
nand UO_172 (O_172,N_6475,N_5792);
nor UO_173 (O_173,N_9679,N_8674);
nor UO_174 (O_174,N_9896,N_9667);
or UO_175 (O_175,N_5812,N_5343);
nor UO_176 (O_176,N_6762,N_8139);
or UO_177 (O_177,N_5486,N_6281);
and UO_178 (O_178,N_9496,N_8848);
and UO_179 (O_179,N_5338,N_6734);
nand UO_180 (O_180,N_7890,N_7098);
nand UO_181 (O_181,N_7350,N_8095);
and UO_182 (O_182,N_5808,N_5902);
nor UO_183 (O_183,N_7589,N_8167);
nor UO_184 (O_184,N_6723,N_5068);
nand UO_185 (O_185,N_5434,N_6061);
and UO_186 (O_186,N_5403,N_9692);
or UO_187 (O_187,N_7667,N_8255);
nor UO_188 (O_188,N_5722,N_7646);
or UO_189 (O_189,N_5608,N_8041);
nor UO_190 (O_190,N_7765,N_5716);
and UO_191 (O_191,N_8749,N_8464);
nand UO_192 (O_192,N_6288,N_7592);
and UO_193 (O_193,N_7416,N_9773);
or UO_194 (O_194,N_8964,N_5525);
and UO_195 (O_195,N_8955,N_5687);
and UO_196 (O_196,N_7869,N_9974);
nor UO_197 (O_197,N_7022,N_7262);
nor UO_198 (O_198,N_8995,N_5661);
nor UO_199 (O_199,N_7670,N_8690);
and UO_200 (O_200,N_8957,N_9250);
and UO_201 (O_201,N_5666,N_7269);
nor UO_202 (O_202,N_5705,N_9588);
or UO_203 (O_203,N_7083,N_7194);
or UO_204 (O_204,N_6271,N_5189);
or UO_205 (O_205,N_8925,N_7953);
nand UO_206 (O_206,N_9636,N_5016);
nor UO_207 (O_207,N_8165,N_8350);
and UO_208 (O_208,N_7804,N_6157);
nand UO_209 (O_209,N_5039,N_5015);
nor UO_210 (O_210,N_6747,N_9895);
nor UO_211 (O_211,N_7057,N_7607);
and UO_212 (O_212,N_5286,N_9611);
and UO_213 (O_213,N_8900,N_7985);
or UO_214 (O_214,N_5412,N_6901);
or UO_215 (O_215,N_7803,N_5112);
nor UO_216 (O_216,N_7734,N_7884);
nor UO_217 (O_217,N_7503,N_7918);
or UO_218 (O_218,N_7114,N_5288);
or UO_219 (O_219,N_6903,N_5145);
nor UO_220 (O_220,N_7227,N_8570);
and UO_221 (O_221,N_9812,N_5521);
or UO_222 (O_222,N_5164,N_9763);
and UO_223 (O_223,N_9623,N_7963);
and UO_224 (O_224,N_5489,N_6064);
nand UO_225 (O_225,N_8262,N_9941);
nand UO_226 (O_226,N_9394,N_9582);
nand UO_227 (O_227,N_9701,N_6143);
nor UO_228 (O_228,N_5549,N_8691);
or UO_229 (O_229,N_5394,N_9970);
nand UO_230 (O_230,N_7896,N_6112);
nand UO_231 (O_231,N_8948,N_7037);
nand UO_232 (O_232,N_6545,N_5141);
nand UO_233 (O_233,N_5764,N_9678);
and UO_234 (O_234,N_6251,N_5361);
nand UO_235 (O_235,N_8324,N_6319);
nand UO_236 (O_236,N_6155,N_9005);
nor UO_237 (O_237,N_5762,N_6994);
nor UO_238 (O_238,N_6821,N_8150);
or UO_239 (O_239,N_5474,N_9865);
or UO_240 (O_240,N_7439,N_7984);
nor UO_241 (O_241,N_9041,N_8234);
nor UO_242 (O_242,N_7957,N_9034);
nand UO_243 (O_243,N_9700,N_7532);
nor UO_244 (O_244,N_9006,N_7533);
nand UO_245 (O_245,N_5965,N_7338);
nand UO_246 (O_246,N_8477,N_8171);
and UO_247 (O_247,N_6409,N_6752);
and UO_248 (O_248,N_9770,N_8097);
and UO_249 (O_249,N_7714,N_8932);
nor UO_250 (O_250,N_6062,N_7505);
or UO_251 (O_251,N_7322,N_8385);
and UO_252 (O_252,N_8855,N_5804);
and UO_253 (O_253,N_6688,N_9138);
xnor UO_254 (O_254,N_9342,N_7436);
nor UO_255 (O_255,N_5156,N_5851);
and UO_256 (O_256,N_5658,N_8910);
nand UO_257 (O_257,N_5309,N_5952);
nor UO_258 (O_258,N_5727,N_6856);
or UO_259 (O_259,N_8270,N_5799);
and UO_260 (O_260,N_7539,N_5693);
or UO_261 (O_261,N_7165,N_9543);
nand UO_262 (O_262,N_5150,N_7679);
nor UO_263 (O_263,N_6429,N_7873);
and UO_264 (O_264,N_7289,N_6611);
and UO_265 (O_265,N_5957,N_6582);
and UO_266 (O_266,N_8525,N_9291);
or UO_267 (O_267,N_5240,N_7240);
nor UO_268 (O_268,N_9862,N_8904);
nand UO_269 (O_269,N_6437,N_5123);
nor UO_270 (O_270,N_6990,N_6601);
and UO_271 (O_271,N_5456,N_9513);
nor UO_272 (O_272,N_8248,N_7857);
nor UO_273 (O_273,N_7507,N_8138);
nor UO_274 (O_274,N_7731,N_7020);
or UO_275 (O_275,N_6523,N_7467);
nor UO_276 (O_276,N_5969,N_9366);
nor UO_277 (O_277,N_7851,N_7563);
nand UO_278 (O_278,N_9090,N_6539);
or UO_279 (O_279,N_6399,N_5697);
or UO_280 (O_280,N_5181,N_8109);
nor UO_281 (O_281,N_8965,N_8624);
nand UO_282 (O_282,N_8382,N_9423);
nand UO_283 (O_283,N_7244,N_5002);
or UO_284 (O_284,N_7945,N_6759);
nand UO_285 (O_285,N_6369,N_5225);
or UO_286 (O_286,N_8297,N_5463);
nand UO_287 (O_287,N_9816,N_8401);
or UO_288 (O_288,N_9961,N_5892);
nand UO_289 (O_289,N_7614,N_8181);
nand UO_290 (O_290,N_8936,N_5711);
and UO_291 (O_291,N_8424,N_9220);
or UO_292 (O_292,N_7591,N_5641);
nand UO_293 (O_293,N_8366,N_6883);
and UO_294 (O_294,N_7264,N_8212);
nor UO_295 (O_295,N_9704,N_6838);
nor UO_296 (O_296,N_7384,N_6035);
nand UO_297 (O_297,N_6930,N_9703);
and UO_298 (O_298,N_9952,N_6291);
nor UO_299 (O_299,N_5328,N_5102);
nand UO_300 (O_300,N_6280,N_5890);
and UO_301 (O_301,N_7064,N_8408);
nand UO_302 (O_302,N_6019,N_5879);
or UO_303 (O_303,N_5206,N_8201);
or UO_304 (O_304,N_7474,N_5339);
nand UO_305 (O_305,N_8617,N_6318);
or UO_306 (O_306,N_7245,N_7780);
nor UO_307 (O_307,N_8963,N_7878);
and UO_308 (O_308,N_7043,N_7555);
or UO_309 (O_309,N_9539,N_8316);
and UO_310 (O_310,N_5273,N_7764);
and UO_311 (O_311,N_8162,N_9118);
and UO_312 (O_312,N_7587,N_5857);
nor UO_313 (O_313,N_6446,N_5910);
or UO_314 (O_314,N_8053,N_5152);
nand UO_315 (O_315,N_8449,N_8622);
nor UO_316 (O_316,N_9986,N_6568);
or UO_317 (O_317,N_5483,N_7317);
xnor UO_318 (O_318,N_7618,N_6401);
nand UO_319 (O_319,N_9485,N_8945);
nand UO_320 (O_320,N_9082,N_9268);
or UO_321 (O_321,N_9499,N_8699);
nor UO_322 (O_322,N_7366,N_8997);
or UO_323 (O_323,N_5903,N_6609);
nor UO_324 (O_324,N_5807,N_8352);
and UO_325 (O_325,N_6690,N_5545);
or UO_326 (O_326,N_8943,N_9916);
or UO_327 (O_327,N_6007,N_9200);
or UO_328 (O_328,N_7480,N_8026);
nor UO_329 (O_329,N_8608,N_8498);
or UO_330 (O_330,N_6000,N_5921);
or UO_331 (O_331,N_5287,N_8891);
xnor UO_332 (O_332,N_6900,N_5344);
nor UO_333 (O_333,N_7808,N_8500);
and UO_334 (O_334,N_7707,N_8200);
or UO_335 (O_335,N_9419,N_8241);
nor UO_336 (O_336,N_6819,N_6668);
nand UO_337 (O_337,N_7965,N_9124);
nand UO_338 (O_338,N_8027,N_8705);
and UO_339 (O_339,N_9519,N_9782);
and UO_340 (O_340,N_5743,N_5080);
nor UO_341 (O_341,N_7966,N_9558);
nand UO_342 (O_342,N_5535,N_6241);
nand UO_343 (O_343,N_6015,N_8312);
xor UO_344 (O_344,N_7872,N_9905);
or UO_345 (O_345,N_6163,N_5096);
nand UO_346 (O_346,N_5647,N_6355);
nor UO_347 (O_347,N_8418,N_9120);
and UO_348 (O_348,N_7982,N_5517);
and UO_349 (O_349,N_8081,N_8453);
and UO_350 (O_350,N_9890,N_8293);
nor UO_351 (O_351,N_9758,N_6248);
or UO_352 (O_352,N_6140,N_9966);
or UO_353 (O_353,N_8244,N_8566);
or UO_354 (O_354,N_5236,N_5638);
and UO_355 (O_355,N_8815,N_7133);
and UO_356 (O_356,N_9654,N_6621);
and UO_357 (O_357,N_6698,N_5085);
nand UO_358 (O_358,N_8349,N_8415);
or UO_359 (O_359,N_7750,N_6458);
nand UO_360 (O_360,N_7981,N_8804);
nand UO_361 (O_361,N_7809,N_5214);
or UO_362 (O_362,N_6918,N_5173);
nand UO_363 (O_363,N_5614,N_8197);
or UO_364 (O_364,N_9557,N_8613);
nor UO_365 (O_365,N_9559,N_8562);
or UO_366 (O_366,N_5054,N_7566);
xnor UO_367 (O_367,N_7934,N_9964);
and UO_368 (O_368,N_6673,N_5859);
and UO_369 (O_369,N_9874,N_7706);
or UO_370 (O_370,N_5410,N_6208);
or UO_371 (O_371,N_6864,N_7415);
nand UO_372 (O_372,N_9395,N_7682);
or UO_373 (O_373,N_7360,N_5373);
nor UO_374 (O_374,N_6150,N_6686);
and UO_375 (O_375,N_8246,N_7989);
and UO_376 (O_376,N_9289,N_6806);
and UO_377 (O_377,N_5868,N_9755);
and UO_378 (O_378,N_9164,N_8683);
or UO_379 (O_379,N_8412,N_7613);
nand UO_380 (O_380,N_8494,N_5269);
and UO_381 (O_381,N_9659,N_7396);
or UO_382 (O_382,N_9383,N_5739);
nand UO_383 (O_383,N_5767,N_7700);
and UO_384 (O_384,N_8961,N_7755);
and UO_385 (O_385,N_9831,N_7754);
and UO_386 (O_386,N_7685,N_6495);
and UO_387 (O_387,N_6246,N_5073);
nand UO_388 (O_388,N_5050,N_9889);
nor UO_389 (O_389,N_8511,N_9438);
nor UO_390 (O_390,N_5745,N_8716);
or UO_391 (O_391,N_5255,N_5585);
nand UO_392 (O_392,N_9348,N_7010);
or UO_393 (O_393,N_6696,N_7325);
nand UO_394 (O_394,N_9044,N_8695);
and UO_395 (O_395,N_7458,N_5595);
or UO_396 (O_396,N_8506,N_9957);
nor UO_397 (O_397,N_6413,N_8715);
nor UO_398 (O_398,N_8659,N_8417);
or UO_399 (O_399,N_8540,N_8721);
and UO_400 (O_400,N_8756,N_7550);
nand UO_401 (O_401,N_6257,N_8103);
and UO_402 (O_402,N_5140,N_5818);
and UO_403 (O_403,N_5644,N_5221);
and UO_404 (O_404,N_6270,N_5217);
nor UO_405 (O_405,N_9219,N_9067);
nor UO_406 (O_406,N_9280,N_5654);
and UO_407 (O_407,N_6788,N_5188);
or UO_408 (O_408,N_7377,N_8021);
or UO_409 (O_409,N_5627,N_7369);
and UO_410 (O_410,N_5127,N_7747);
or UO_411 (O_411,N_6512,N_8439);
nand UO_412 (O_412,N_9017,N_9573);
nor UO_413 (O_413,N_9590,N_5971);
nand UO_414 (O_414,N_9218,N_9781);
and UO_415 (O_415,N_9838,N_5772);
nor UO_416 (O_416,N_8012,N_7071);
nand UO_417 (O_417,N_8051,N_9924);
or UO_418 (O_418,N_8552,N_6261);
nand UO_419 (O_419,N_5299,N_9520);
nand UO_420 (O_420,N_9373,N_5770);
or UO_421 (O_421,N_8557,N_8931);
nor UO_422 (O_422,N_9922,N_9294);
nor UO_423 (O_423,N_8751,N_9424);
or UO_424 (O_424,N_5368,N_8868);
nor UO_425 (O_425,N_8939,N_8131);
and UO_426 (O_426,N_7140,N_7839);
nand UO_427 (O_427,N_5865,N_8240);
and UO_428 (O_428,N_9851,N_6173);
or UO_429 (O_429,N_9767,N_9468);
nand UO_430 (O_430,N_6438,N_7688);
nor UO_431 (O_431,N_9465,N_5784);
nor UO_432 (O_432,N_8375,N_8208);
or UO_433 (O_433,N_9617,N_5191);
nand UO_434 (O_434,N_7182,N_5186);
nand UO_435 (O_435,N_8284,N_8680);
or UO_436 (O_436,N_9455,N_8213);
nand UO_437 (O_437,N_9618,N_6879);
nor UO_438 (O_438,N_8086,N_5567);
and UO_439 (O_439,N_7815,N_8652);
nor UO_440 (O_440,N_8899,N_7522);
nor UO_441 (O_441,N_7216,N_7572);
and UO_442 (O_442,N_6616,N_8547);
nor UO_443 (O_443,N_8431,N_9840);
or UO_444 (O_444,N_9182,N_5519);
and UO_445 (O_445,N_9512,N_8295);
or UO_446 (O_446,N_7229,N_7072);
or UO_447 (O_447,N_6427,N_9856);
and UO_448 (O_448,N_7274,N_7164);
nand UO_449 (O_449,N_5538,N_7846);
xnor UO_450 (O_450,N_9314,N_5795);
nand UO_451 (O_451,N_7411,N_5475);
nand UO_452 (O_452,N_8517,N_5659);
and UO_453 (O_453,N_6334,N_5295);
nand UO_454 (O_454,N_5996,N_9025);
nor UO_455 (O_455,N_5021,N_5045);
nor UO_456 (O_456,N_9929,N_5616);
nor UO_457 (O_457,N_7882,N_5708);
nor UO_458 (O_458,N_9761,N_5732);
nand UO_459 (O_459,N_5497,N_8437);
nand UO_460 (O_460,N_8376,N_7266);
and UO_461 (O_461,N_7299,N_9391);
nand UO_462 (O_462,N_9933,N_9076);
and UO_463 (O_463,N_9121,N_9191);
nor UO_464 (O_464,N_6224,N_9783);
and UO_465 (O_465,N_5856,N_9686);
nor UO_466 (O_466,N_8632,N_7868);
nand UO_467 (O_467,N_5117,N_7016);
nor UO_468 (O_468,N_7546,N_8578);
or UO_469 (O_469,N_5599,N_9134);
or UO_470 (O_470,N_8538,N_6050);
or UO_471 (O_471,N_7028,N_8959);
nand UO_472 (O_472,N_6195,N_9613);
nand UO_473 (O_473,N_7597,N_5835);
and UO_474 (O_474,N_5259,N_7447);
nor UO_475 (O_475,N_5803,N_5227);
nand UO_476 (O_476,N_8610,N_7178);
and UO_477 (O_477,N_8858,N_6799);
nor UO_478 (O_478,N_7569,N_8018);
nand UO_479 (O_479,N_6400,N_8543);
nand UO_480 (O_480,N_8919,N_6388);
or UO_481 (O_481,N_5837,N_8402);
nand UO_482 (O_482,N_9508,N_6217);
or UO_483 (O_483,N_6121,N_5063);
and UO_484 (O_484,N_8230,N_7257);
nand UO_485 (O_485,N_8450,N_5059);
nand UO_486 (O_486,N_6999,N_7761);
and UO_487 (O_487,N_7631,N_7654);
nand UO_488 (O_488,N_6805,N_8137);
and UO_489 (O_489,N_6849,N_5153);
or UO_490 (O_490,N_6634,N_5128);
nor UO_491 (O_491,N_7307,N_9409);
and UO_492 (O_492,N_9995,N_6655);
nor UO_493 (O_493,N_9443,N_5298);
and UO_494 (O_494,N_9046,N_8170);
and UO_495 (O_495,N_6404,N_9149);
or UO_496 (O_496,N_8445,N_5898);
nor UO_497 (O_497,N_6459,N_9673);
and UO_498 (O_498,N_7703,N_8663);
nand UO_499 (O_499,N_7446,N_5175);
or UO_500 (O_500,N_7814,N_9392);
nand UO_501 (O_501,N_5577,N_8345);
nand UO_502 (O_502,N_5825,N_9115);
and UO_503 (O_503,N_7916,N_7838);
nor UO_504 (O_504,N_8269,N_7235);
or UO_505 (O_505,N_5999,N_9942);
nor UO_506 (O_506,N_9926,N_6518);
or UO_507 (O_507,N_5980,N_8132);
nand UO_508 (O_508,N_9376,N_8675);
or UO_509 (O_509,N_5547,N_6160);
nand UO_510 (O_510,N_9891,N_8795);
nor UO_511 (O_511,N_7720,N_7427);
nand UO_512 (O_512,N_5176,N_7290);
nor UO_513 (O_513,N_9035,N_6211);
nand UO_514 (O_514,N_6510,N_8274);
or UO_515 (O_515,N_8268,N_8198);
or UO_516 (O_516,N_7961,N_6840);
nand UO_517 (O_517,N_5755,N_7078);
or UO_518 (O_518,N_7802,N_8231);
and UO_519 (O_519,N_7051,N_8281);
and UO_520 (O_520,N_9965,N_7404);
nand UO_521 (O_521,N_6046,N_7158);
nand UO_522 (O_522,N_9070,N_5704);
and UO_523 (O_523,N_5347,N_5904);
nor UO_524 (O_524,N_8962,N_8727);
nand UO_525 (O_525,N_9266,N_8017);
or UO_526 (O_526,N_7180,N_8656);
or UO_527 (O_527,N_8100,N_8115);
nor UO_528 (O_528,N_8688,N_7344);
and UO_529 (O_529,N_7930,N_7786);
nor UO_530 (O_530,N_7845,N_5509);
or UO_531 (O_531,N_8296,N_9039);
nand UO_532 (O_532,N_6284,N_9864);
and UO_533 (O_533,N_8993,N_9664);
nand UO_534 (O_534,N_5963,N_5466);
nor UO_535 (O_535,N_7241,N_8813);
or UO_536 (O_536,N_5469,N_9014);
nand UO_537 (O_537,N_8763,N_8406);
and UO_538 (O_538,N_6460,N_9466);
nand UO_539 (O_539,N_6632,N_5402);
nand UO_540 (O_540,N_7161,N_5115);
nor UO_541 (O_541,N_8823,N_7060);
or UO_542 (O_542,N_7520,N_6220);
nand UO_543 (O_543,N_5108,N_9047);
nor UO_544 (O_544,N_7017,N_5439);
nand UO_545 (O_545,N_6165,N_6743);
or UO_546 (O_546,N_8479,N_8696);
and UO_547 (O_547,N_9359,N_6259);
and UO_548 (O_548,N_5089,N_6415);
and UO_549 (O_549,N_9746,N_8738);
or UO_550 (O_550,N_9074,N_8847);
or UO_551 (O_551,N_8435,N_8119);
nor UO_552 (O_552,N_9677,N_9811);
or UO_553 (O_553,N_6192,N_8713);
and UO_554 (O_554,N_8820,N_9578);
nand UO_555 (O_555,N_8574,N_5507);
nand UO_556 (O_556,N_6920,N_6330);
and UO_557 (O_557,N_5400,N_9936);
nor UO_558 (O_558,N_5651,N_5012);
or UO_559 (O_559,N_5782,N_6769);
and UO_560 (O_560,N_6715,N_8067);
nand UO_561 (O_561,N_7691,N_7900);
nand UO_562 (O_562,N_9696,N_8911);
or UO_563 (O_563,N_7199,N_9585);
nand UO_564 (O_564,N_9658,N_8698);
or UO_565 (O_565,N_7041,N_9137);
and UO_566 (O_566,N_8707,N_6595);
and UO_567 (O_567,N_6801,N_8254);
and UO_568 (O_568,N_5215,N_5933);
nor UO_569 (O_569,N_5578,N_6542);
and UO_570 (O_570,N_8340,N_8377);
or UO_571 (O_571,N_7823,N_6885);
and UO_572 (O_572,N_7888,N_9053);
and UO_573 (O_573,N_7205,N_9902);
and UO_574 (O_574,N_6931,N_7144);
and UO_575 (O_575,N_6010,N_9222);
and UO_576 (O_576,N_6719,N_7221);
nor UO_577 (O_577,N_9939,N_6469);
nand UO_578 (O_578,N_7907,N_7645);
and UO_579 (O_579,N_5453,N_7944);
and UO_580 (O_580,N_9054,N_6543);
nand UO_581 (O_581,N_6708,N_7757);
or UO_582 (O_582,N_6447,N_5562);
and UO_583 (O_583,N_7334,N_8010);
nor UO_584 (O_584,N_6044,N_7774);
and UO_585 (O_585,N_5861,N_5022);
and UO_586 (O_586,N_8810,N_7659);
and UO_587 (O_587,N_9774,N_6250);
nor UO_588 (O_588,N_8907,N_8797);
and UO_589 (O_589,N_5544,N_6054);
nor UO_590 (O_590,N_9287,N_9461);
nor UO_591 (O_591,N_9426,N_8070);
or UO_592 (O_592,N_6978,N_7323);
and UO_593 (O_593,N_8974,N_5660);
and UO_594 (O_594,N_8459,N_5719);
nand UO_595 (O_595,N_6471,N_7457);
nand UO_596 (O_596,N_8307,N_6638);
nor UO_597 (O_597,N_8971,N_5994);
and UO_598 (O_598,N_6746,N_7867);
nand UO_599 (O_599,N_9073,N_5875);
or UO_600 (O_600,N_7603,N_6449);
and UO_601 (O_601,N_9243,N_5640);
or UO_602 (O_602,N_5067,N_5318);
nand UO_603 (O_603,N_5682,N_7038);
and UO_604 (O_604,N_6934,N_6287);
or UO_605 (O_605,N_6586,N_8667);
nor UO_606 (O_606,N_8423,N_7378);
xnor UO_607 (O_607,N_7897,N_6094);
nand UO_608 (O_608,N_7414,N_9788);
and UO_609 (O_609,N_7138,N_8083);
nand UO_610 (O_610,N_6228,N_7531);
and UO_611 (O_611,N_7915,N_5560);
and UO_612 (O_612,N_8153,N_8968);
and UO_613 (O_613,N_8840,N_9393);
and UO_614 (O_614,N_7473,N_9769);
and UO_615 (O_615,N_7450,N_6335);
or UO_616 (O_616,N_5498,N_6858);
and UO_617 (O_617,N_7488,N_9019);
nor UO_618 (O_618,N_5091,N_5293);
nand UO_619 (O_619,N_9217,N_8863);
or UO_620 (O_620,N_9476,N_9486);
nand UO_621 (O_621,N_7988,N_7722);
and UO_622 (O_622,N_8087,N_6957);
nor UO_623 (O_623,N_6328,N_7837);
and UO_624 (O_624,N_7186,N_7920);
nor UO_625 (O_625,N_9358,N_6873);
or UO_626 (O_626,N_8286,N_5097);
and UO_627 (O_627,N_6905,N_6812);
nand UO_628 (O_628,N_9307,N_8140);
or UO_629 (O_629,N_5828,N_6051);
nand UO_630 (O_630,N_9886,N_6343);
and UO_631 (O_631,N_6996,N_5436);
or UO_632 (O_632,N_8876,N_6393);
or UO_633 (O_633,N_7025,N_5192);
and UO_634 (O_634,N_9281,N_6350);
nand UO_635 (O_635,N_6764,N_8549);
and UO_636 (O_636,N_6598,N_7954);
or UO_637 (O_637,N_8934,N_7238);
nor UO_638 (O_638,N_5876,N_7434);
or UO_639 (O_639,N_5718,N_5995);
nand UO_640 (O_640,N_5964,N_5033);
and UO_641 (O_641,N_8020,N_9368);
nor UO_642 (O_642,N_9112,N_9598);
nand UO_643 (O_643,N_8023,N_6700);
nand UO_644 (O_644,N_9146,N_6465);
and UO_645 (O_645,N_7537,N_5609);
nand UO_646 (O_646,N_8542,N_6114);
and UO_647 (O_647,N_6915,N_7652);
nor UO_648 (O_648,N_8353,N_6134);
nor UO_649 (O_649,N_5199,N_6077);
and UO_650 (O_650,N_9707,N_8660);
and UO_651 (O_651,N_6186,N_5118);
and UO_652 (O_652,N_5315,N_8251);
nor UO_653 (O_653,N_5322,N_6610);
nor UO_654 (O_654,N_6950,N_8529);
nor UO_655 (O_655,N_6472,N_6336);
and UO_656 (O_656,N_8730,N_9710);
and UO_657 (O_657,N_7065,N_9272);
or UO_658 (O_658,N_5596,N_9065);
nor UO_659 (O_659,N_7895,N_5779);
nand UO_660 (O_660,N_6048,N_7743);
nand UO_661 (O_661,N_8942,N_5556);
and UO_662 (O_662,N_9403,N_8554);
nand UO_663 (O_663,N_7459,N_6131);
nor UO_664 (O_664,N_6570,N_5332);
nand UO_665 (O_665,N_7270,N_7622);
nor UO_666 (O_666,N_6363,N_8036);
or UO_667 (O_667,N_7387,N_9467);
or UO_668 (O_668,N_9495,N_6809);
nor UO_669 (O_669,N_8768,N_6153);
nor UO_670 (O_670,N_5729,N_7960);
and UO_671 (O_671,N_7737,N_6254);
nor UO_672 (O_672,N_7424,N_9412);
nand UO_673 (O_673,N_5975,N_6745);
nand UO_674 (O_674,N_7139,N_6814);
nand UO_675 (O_675,N_5356,N_5187);
nand UO_676 (O_676,N_5473,N_7593);
nand UO_677 (O_677,N_6193,N_9003);
nor UO_678 (O_678,N_6206,N_6509);
or UO_679 (O_679,N_9249,N_5487);
and UO_680 (O_680,N_9308,N_6807);
or UO_681 (O_681,N_5296,N_6825);
nor UO_682 (O_682,N_9607,N_7362);
nand UO_683 (O_683,N_5974,N_5927);
and UO_684 (O_684,N_6293,N_6435);
or UO_685 (O_685,N_6126,N_9609);
nand UO_686 (O_686,N_8766,N_7509);
nor UO_687 (O_687,N_5204,N_9702);
nor UO_688 (O_688,N_5447,N_6002);
nor UO_689 (O_689,N_9340,N_5314);
nor UO_690 (O_690,N_7011,N_7819);
and UO_691 (O_691,N_8309,N_7493);
nor UO_692 (O_692,N_9602,N_5249);
or UO_693 (O_693,N_6122,N_6818);
nor UO_694 (O_694,N_8099,N_9894);
xnor UO_695 (O_695,N_5131,N_5084);
or UO_696 (O_696,N_5284,N_6617);
and UO_697 (O_697,N_7380,N_7210);
and UO_698 (O_698,N_8466,N_7687);
and UO_699 (O_699,N_7177,N_6776);
nor UO_700 (O_700,N_8643,N_7498);
nand UO_701 (O_701,N_9853,N_9197);
and UO_702 (O_702,N_7588,N_5028);
nand UO_703 (O_703,N_5636,N_5137);
nand UO_704 (O_704,N_7914,N_5126);
and UO_705 (O_705,N_9144,N_9906);
nand UO_706 (O_706,N_7409,N_8348);
and UO_707 (O_707,N_5703,N_5731);
nand UO_708 (O_708,N_8069,N_6939);
nor UO_709 (O_709,N_9532,N_9080);
or UO_710 (O_710,N_6124,N_7385);
and UO_711 (O_711,N_8034,N_6269);
and UO_712 (O_712,N_8129,N_7841);
and UO_713 (O_713,N_7651,N_6922);
or UO_714 (O_714,N_5363,N_7319);
or UO_715 (O_715,N_9346,N_8623);
and UO_716 (O_716,N_8544,N_8242);
or UO_717 (O_717,N_9444,N_5816);
nand UO_718 (O_718,N_9668,N_5094);
or UO_719 (O_719,N_6286,N_9796);
nor UO_720 (O_720,N_8889,N_9835);
and UO_721 (O_721,N_8913,N_9572);
or UO_722 (O_722,N_9274,N_7142);
and UO_723 (O_723,N_6536,N_5680);
nand UO_724 (O_724,N_7425,N_6262);
nor UO_725 (O_725,N_8184,N_7119);
nand UO_726 (O_726,N_7413,N_9982);
or UO_727 (O_727,N_7339,N_8050);
nor UO_728 (O_728,N_6566,N_6483);
nor UO_729 (O_729,N_5694,N_8460);
and UO_730 (O_730,N_7054,N_6078);
nor UO_731 (O_731,N_8969,N_6354);
nand UO_732 (O_732,N_5529,N_6376);
or UO_733 (O_733,N_9415,N_7306);
nand UO_734 (O_734,N_8743,N_5981);
or UO_735 (O_735,N_7719,N_8555);
nand UO_736 (O_736,N_5391,N_8215);
nor UO_737 (O_737,N_7925,N_6130);
and UO_738 (O_738,N_5093,N_6249);
nand UO_739 (O_739,N_5673,N_8058);
nor UO_740 (O_740,N_9550,N_6025);
and UO_741 (O_741,N_6717,N_6962);
or UO_742 (O_742,N_8612,N_8661);
and UO_743 (O_743,N_5077,N_6741);
or UO_744 (O_744,N_6727,N_6406);
nor UO_745 (O_745,N_6973,N_9363);
nor UO_746 (O_746,N_7273,N_9656);
or UO_747 (O_747,N_5573,N_8386);
nand UO_748 (O_748,N_9949,N_8563);
and UO_749 (O_749,N_9718,N_6505);
or UO_750 (O_750,N_7936,N_9960);
or UO_751 (O_751,N_6887,N_5031);
nor UO_752 (O_752,N_6706,N_8457);
and UO_753 (O_753,N_5446,N_6170);
and UO_754 (O_754,N_7643,N_7889);
nand UO_755 (O_755,N_8976,N_9051);
or UO_756 (O_756,N_8720,N_5276);
and UO_757 (O_757,N_7541,N_7939);
nor UO_758 (O_758,N_8553,N_6697);
or UO_759 (O_759,N_8285,N_9265);
xnor UO_760 (O_760,N_9436,N_6695);
or UO_761 (O_761,N_6384,N_8223);
and UO_762 (O_762,N_8966,N_8280);
or UO_763 (O_763,N_6704,N_8019);
nor UO_764 (O_764,N_9038,N_8793);
nor UO_765 (O_765,N_7718,N_8779);
and UO_766 (O_766,N_9007,N_6171);
nor UO_767 (O_767,N_6971,N_9096);
or UO_768 (O_768,N_9093,N_6804);
or UO_769 (O_769,N_7176,N_9538);
and UO_770 (O_770,N_9167,N_7574);
or UO_771 (O_771,N_9242,N_6628);
and UO_772 (O_772,N_6817,N_6428);
nor UO_773 (O_773,N_8774,N_6237);
nor UO_774 (O_774,N_8785,N_6940);
and UO_775 (O_775,N_6936,N_9911);
nand UO_776 (O_776,N_8387,N_6041);
nand UO_777 (O_777,N_6863,N_6266);
or UO_778 (O_778,N_8647,N_7716);
and UO_779 (O_779,N_9971,N_8029);
nor UO_780 (O_780,N_9504,N_9793);
nor UO_781 (O_781,N_8163,N_8894);
and UO_782 (O_782,N_6862,N_8780);
and UO_783 (O_783,N_9026,N_9836);
nand UO_784 (O_784,N_5348,N_6898);
nand UO_785 (O_785,N_8259,N_6842);
or UO_786 (O_786,N_6226,N_5375);
and UO_787 (O_787,N_7642,N_8078);
nand UO_788 (O_788,N_5581,N_5366);
or UO_789 (O_789,N_7070,N_7777);
nand UO_790 (O_790,N_8534,N_9077);
or UO_791 (O_791,N_6878,N_9951);
and UO_792 (O_792,N_9312,N_6120);
nand UO_793 (O_793,N_5615,N_9555);
and UO_794 (O_794,N_8719,N_6853);
nand UO_795 (O_795,N_6325,N_7428);
or UO_796 (O_796,N_5208,N_7258);
and UO_797 (O_797,N_5194,N_7090);
and UO_798 (O_798,N_6057,N_7335);
nor UO_799 (O_799,N_8179,N_5738);
nor UO_800 (O_800,N_8323,N_9361);
or UO_801 (O_801,N_9160,N_8605);
and UO_802 (O_802,N_5679,N_8442);
nor UO_803 (O_803,N_8388,N_7073);
and UO_804 (O_804,N_5069,N_8325);
nand UO_805 (O_805,N_6635,N_9434);
and UO_806 (O_806,N_5576,N_7542);
or UO_807 (O_807,N_8972,N_7817);
nor UO_808 (O_808,N_7668,N_6091);
nand UO_809 (O_809,N_6424,N_8783);
nor UO_810 (O_810,N_8261,N_8399);
and UO_811 (O_811,N_5721,N_6511);
nand UO_812 (O_812,N_7373,N_9899);
and UO_813 (O_813,N_8545,N_5183);
nand UO_814 (O_814,N_9569,N_9128);
and UO_815 (O_815,N_5484,N_9878);
or UO_816 (O_816,N_6310,N_6982);
nor UO_817 (O_817,N_7137,N_5834);
and UO_818 (O_818,N_5292,N_7732);
and UO_819 (O_819,N_8784,N_9113);
nand UO_820 (O_820,N_9013,N_6347);
nor UO_821 (O_821,N_8927,N_7513);
nor UO_822 (O_822,N_5991,N_5926);
and UO_823 (O_823,N_6216,N_9544);
nor UO_824 (O_824,N_6932,N_6166);
nor UO_825 (O_825,N_6755,N_6049);
nand UO_826 (O_826,N_7268,N_6763);
nand UO_827 (O_827,N_9141,N_7247);
nor UO_828 (O_828,N_9233,N_7508);
and UO_829 (O_829,N_7222,N_8194);
and UO_830 (O_830,N_8735,N_8603);
and UO_831 (O_831,N_5053,N_5306);
and UO_832 (O_832,N_6808,N_9126);
nor UO_833 (O_833,N_6653,N_6299);
nor UO_834 (O_834,N_6277,N_9048);
or UO_835 (O_835,N_8174,N_6989);
or UO_836 (O_836,N_8597,N_9753);
or UO_837 (O_837,N_6658,N_8616);
or UO_838 (O_838,N_9216,N_9241);
and UO_839 (O_839,N_5008,N_7026);
nand UO_840 (O_840,N_7421,N_7316);
nand UO_841 (O_841,N_8322,N_6434);
and UO_842 (O_842,N_8890,N_5515);
nor UO_843 (O_843,N_7260,N_5303);
nand UO_844 (O_844,N_8596,N_8214);
or UO_845 (O_845,N_8807,N_5548);
nand UO_846 (O_846,N_7233,N_5737);
or UO_847 (O_847,N_7640,N_7958);
or UO_848 (O_848,N_9213,N_7174);
and UO_849 (O_849,N_5340,N_7305);
and UO_850 (O_850,N_6870,N_6162);
and UO_851 (O_851,N_9565,N_8836);
nor UO_852 (O_852,N_8074,N_9004);
nor UO_853 (O_853,N_9068,N_9801);
and UO_854 (O_854,N_7665,N_5998);
nor UO_855 (O_855,N_5124,N_9105);
nand UO_856 (O_856,N_7433,N_7616);
or UO_857 (O_857,N_7567,N_5211);
or UO_858 (O_858,N_8277,N_9169);
nor UO_859 (O_859,N_6524,N_7927);
nor UO_860 (O_860,N_8499,N_8302);
or UO_861 (O_861,N_6298,N_5510);
nand UO_862 (O_862,N_8722,N_8877);
or UO_863 (O_863,N_8762,N_5855);
and UO_864 (O_864,N_7909,N_9850);
nor UO_865 (O_865,N_8428,N_7677);
and UO_866 (O_866,N_6722,N_7692);
nand UO_867 (O_867,N_5777,N_6569);
or UO_868 (O_868,N_9567,N_5823);
nand UO_869 (O_869,N_8657,N_7198);
or UO_870 (O_870,N_7968,N_6079);
or UO_871 (O_871,N_7336,N_9843);
or UO_872 (O_872,N_7254,N_5425);
nand UO_873 (O_873,N_9229,N_5461);
nand UO_874 (O_874,N_9586,N_7093);
or UO_875 (O_875,N_8590,N_6500);
nor UO_876 (O_876,N_7002,N_9804);
nor UO_877 (O_877,N_6089,N_8191);
or UO_878 (O_878,N_5805,N_8627);
nor UO_879 (O_879,N_7584,N_9992);
nor UO_880 (O_880,N_5814,N_9107);
and UO_881 (O_881,N_9713,N_8600);
nor UO_882 (O_882,N_7091,N_6798);
nor UO_883 (O_883,N_5200,N_7412);
or UO_884 (O_884,N_8592,N_7465);
nor UO_885 (O_885,N_5539,N_7661);
and UO_886 (O_886,N_9305,N_7500);
or UO_887 (O_887,N_8520,N_5178);
nor UO_888 (O_888,N_9697,N_5985);
or UO_889 (O_889,N_5815,N_9300);
or UO_890 (O_890,N_6662,N_8677);
and UO_891 (O_891,N_9020,N_9847);
nand UO_892 (O_892,N_6608,N_8337);
nand UO_893 (O_893,N_5844,N_7168);
nand UO_894 (O_894,N_8458,N_7173);
and UO_895 (O_895,N_6977,N_9062);
or UO_896 (O_896,N_9791,N_8940);
and UO_897 (O_897,N_8973,N_8828);
nand UO_898 (O_898,N_9251,N_7181);
nor UO_899 (O_899,N_7810,N_7902);
and UO_900 (O_900,N_7556,N_9869);
nand UO_901 (O_901,N_8491,N_9151);
and UO_902 (O_902,N_5180,N_9604);
nor UO_903 (O_903,N_7056,N_9347);
nand UO_904 (O_904,N_9817,N_7374);
nor UO_905 (O_905,N_9102,N_6327);
or UO_906 (O_906,N_6710,N_8055);
or UO_907 (O_907,N_7580,N_9109);
or UO_908 (O_908,N_8844,N_7949);
and UO_909 (O_909,N_7689,N_5747);
or UO_910 (O_910,N_8519,N_6624);
nor UO_911 (O_911,N_9691,N_8568);
and UO_912 (O_912,N_8022,N_8539);
and UO_913 (O_913,N_6919,N_5559);
or UO_914 (O_914,N_9842,N_7368);
nor UO_915 (O_915,N_8374,N_6564);
nand UO_916 (O_916,N_7187,N_8392);
or UO_917 (O_917,N_9515,N_7294);
nand UO_918 (O_918,N_8501,N_6282);
and UO_919 (O_919,N_8960,N_7752);
nand UO_920 (O_920,N_5334,N_6470);
and UO_921 (O_921,N_6442,N_7189);
nand UO_922 (O_922,N_8032,N_5646);
and UO_923 (O_923,N_9135,N_5566);
nor UO_924 (O_924,N_6063,N_9828);
nand UO_925 (O_925,N_5610,N_7669);
or UO_926 (O_926,N_5442,N_8649);
nand UO_927 (O_927,N_9326,N_7069);
nor UO_928 (O_928,N_8178,N_8249);
nand UO_929 (O_929,N_6383,N_5759);
and UO_930 (O_930,N_6053,N_7885);
nor UO_931 (O_931,N_6824,N_6304);
or UO_932 (O_932,N_5900,N_7109);
or UO_933 (O_933,N_6623,N_8892);
nor UO_934 (O_934,N_6387,N_7284);
or UO_935 (O_935,N_9762,N_8648);
nor UO_936 (O_936,N_8104,N_6482);
nor UO_937 (O_937,N_7400,N_9125);
or UO_938 (O_938,N_8257,N_5657);
nand UO_939 (O_939,N_5430,N_7353);
nor UO_940 (O_940,N_5907,N_6906);
or UO_941 (O_941,N_9397,N_8625);
nor UO_942 (O_942,N_5499,N_8703);
nand UO_943 (O_943,N_5628,N_9442);
or UO_944 (O_944,N_5631,N_6909);
nor UO_945 (O_945,N_6087,N_7225);
nand UO_946 (O_946,N_8887,N_6692);
and UO_947 (O_947,N_7234,N_6309);
nor UO_948 (O_948,N_9694,N_8761);
and UO_949 (O_949,N_7285,N_6412);
nand UO_950 (O_950,N_6756,N_9927);
or UO_951 (O_951,N_9260,N_7463);
nand UO_952 (O_952,N_8124,N_9945);
nand UO_953 (O_953,N_9143,N_5571);
or UO_954 (O_954,N_5829,N_5025);
and UO_955 (O_955,N_5301,N_9410);
nor UO_956 (O_956,N_6480,N_7259);
or UO_957 (O_957,N_9711,N_5941);
nor UO_958 (O_958,N_6499,N_6620);
and UO_959 (O_959,N_6223,N_6141);
and UO_960 (O_960,N_6232,N_9173);
nor UO_961 (O_961,N_5017,N_6839);
nand UO_962 (O_962,N_7617,N_7200);
or UO_963 (O_963,N_6783,N_5049);
or UO_964 (O_964,N_6560,N_9079);
and UO_965 (O_965,N_5238,N_8169);
nand UO_966 (O_966,N_5972,N_8260);
and UO_967 (O_967,N_5976,N_8923);
nor UO_968 (O_968,N_5906,N_8577);
nor UO_969 (O_969,N_7372,N_6615);
and UO_970 (O_970,N_6661,N_5516);
nand UO_971 (O_971,N_9171,N_6161);
nor UO_972 (O_972,N_5316,N_5966);
or UO_973 (O_973,N_8777,N_7302);
or UO_974 (O_974,N_8983,N_6657);
and UO_975 (O_975,N_9175,N_5100);
nor UO_976 (O_976,N_6952,N_9683);
and UO_977 (O_977,N_5182,N_5471);
and UO_978 (O_978,N_9375,N_6528);
nor UO_979 (O_979,N_5881,N_9040);
nor UO_980 (O_980,N_6835,N_5882);
nor UO_981 (O_981,N_5960,N_7715);
nand UO_982 (O_982,N_6561,N_5569);
or UO_983 (O_983,N_9988,N_6521);
nor UO_984 (O_984,N_8045,N_7807);
nand UO_985 (O_985,N_6313,N_7850);
nor UO_986 (O_986,N_8835,N_6275);
and UO_987 (O_987,N_8796,N_6238);
nand UO_988 (O_988,N_5656,N_8127);
and UO_989 (O_989,N_6714,N_7636);
and UO_990 (O_990,N_9369,N_5754);
and UO_991 (O_991,N_6572,N_7104);
nand UO_992 (O_992,N_5677,N_9646);
nand UO_993 (O_993,N_9522,N_8484);
nor UO_994 (O_994,N_6874,N_7085);
nand UO_995 (O_995,N_8422,N_5736);
and UO_996 (O_996,N_7297,N_7125);
nor UO_997 (O_997,N_5230,N_8859);
or UO_998 (O_998,N_9159,N_8975);
and UO_999 (O_999,N_5457,N_5688);
or UO_1000 (O_1000,N_9275,N_7686);
nor UO_1001 (O_1001,N_6559,N_9259);
nor UO_1002 (O_1002,N_8420,N_8986);
nand UO_1003 (O_1003,N_8313,N_6072);
nand UO_1004 (O_1004,N_6382,N_9012);
or UO_1005 (O_1005,N_5154,N_6683);
or UO_1006 (O_1006,N_7858,N_9194);
and UO_1007 (O_1007,N_8253,N_5321);
nor UO_1008 (O_1008,N_7863,N_5920);
and UO_1009 (O_1009,N_8755,N_6498);
and UO_1010 (O_1010,N_5665,N_7106);
and UO_1011 (O_1011,N_8130,N_5237);
or UO_1012 (O_1012,N_8634,N_9561);
and UO_1013 (O_1013,N_7403,N_5177);
nor UO_1014 (O_1014,N_9599,N_7813);
or UO_1015 (O_1015,N_6802,N_5676);
and UO_1016 (O_1016,N_6882,N_9994);
nand UO_1017 (O_1017,N_9060,N_8362);
nor UO_1018 (O_1018,N_8452,N_7608);
nor UO_1019 (O_1019,N_8938,N_5203);
and UO_1020 (O_1020,N_8485,N_7481);
or UO_1021 (O_1021,N_8149,N_5901);
or UO_1022 (O_1022,N_7560,N_8001);
nor UO_1023 (O_1023,N_6843,N_5114);
nand UO_1024 (O_1024,N_9204,N_9301);
nand UO_1025 (O_1025,N_9130,N_5163);
nand UO_1026 (O_1026,N_9634,N_9931);
nand UO_1027 (O_1027,N_6767,N_9011);
xor UO_1028 (O_1028,N_5526,N_5720);
and UO_1029 (O_1029,N_7736,N_6476);
and UO_1030 (O_1030,N_5243,N_8291);
nand UO_1031 (O_1031,N_6985,N_5377);
or UO_1032 (O_1032,N_5162,N_8471);
and UO_1033 (O_1033,N_9876,N_9750);
or UO_1034 (O_1034,N_9638,N_9433);
nor UO_1035 (O_1035,N_5407,N_6027);
nor UO_1036 (O_1036,N_6828,N_6891);
and UO_1037 (O_1037,N_7634,N_8356);
and UO_1038 (O_1038,N_7554,N_5602);
and UO_1039 (O_1039,N_5723,N_9343);
nor UO_1040 (O_1040,N_6599,N_9560);
nor UO_1041 (O_1041,N_6332,N_7964);
nand UO_1042 (O_1042,N_6329,N_7834);
nand UO_1043 (O_1043,N_8225,N_7741);
nand UO_1044 (O_1044,N_9271,N_8953);
nor UO_1045 (O_1045,N_8156,N_5423);
or UO_1046 (O_1046,N_9893,N_5490);
and UO_1047 (O_1047,N_5151,N_8723);
nand UO_1048 (O_1048,N_7926,N_6975);
nand UO_1049 (O_1049,N_5197,N_9627);
nand UO_1050 (O_1050,N_8841,N_9518);
or UO_1051 (O_1051,N_9108,N_6182);
or UO_1052 (O_1052,N_5034,N_7975);
and UO_1053 (O_1053,N_5839,N_6703);
or UO_1054 (O_1054,N_5532,N_8071);
and UO_1055 (O_1055,N_8250,N_6375);
nor UO_1056 (O_1056,N_6876,N_6253);
and UO_1057 (O_1057,N_7523,N_9632);
or UO_1058 (O_1058,N_7393,N_8470);
nand UO_1059 (O_1059,N_6941,N_7352);
or UO_1060 (O_1060,N_6855,N_7799);
nor UO_1061 (O_1061,N_6198,N_9475);
and UO_1062 (O_1062,N_7893,N_5537);
or UO_1063 (O_1063,N_6292,N_8929);
and UO_1064 (O_1064,N_9778,N_5843);
and UO_1065 (O_1065,N_5905,N_9337);
nor UO_1066 (O_1066,N_5184,N_6410);
nor UO_1067 (O_1067,N_8326,N_9098);
or UO_1068 (O_1068,N_5300,N_6605);
nor UO_1069 (O_1069,N_9803,N_5493);
nor UO_1070 (O_1070,N_6927,N_5263);
or UO_1071 (O_1071,N_6006,N_7623);
nand UO_1072 (O_1072,N_5035,N_8496);
nand UO_1073 (O_1073,N_5864,N_7159);
or UO_1074 (O_1074,N_8681,N_8072);
xor UO_1075 (O_1075,N_7763,N_9180);
or UO_1076 (O_1076,N_7871,N_7001);
and UO_1077 (O_1077,N_5841,N_9248);
and UO_1078 (O_1078,N_7392,N_7962);
and UO_1079 (O_1079,N_5038,N_7097);
and UO_1080 (O_1080,N_9396,N_8048);
nand UO_1081 (O_1081,N_6832,N_8073);
nor UO_1082 (O_1082,N_7482,N_8671);
or UO_1083 (O_1083,N_6423,N_6295);
or UO_1084 (O_1084,N_6402,N_6771);
nor UO_1085 (O_1085,N_6827,N_9309);
or UO_1086 (O_1086,N_9661,N_9728);
or UO_1087 (O_1087,N_9775,N_6467);
and UO_1088 (O_1088,N_9325,N_5401);
nor UO_1089 (O_1089,N_7304,N_6177);
or UO_1090 (O_1090,N_7635,N_8486);
nand UO_1091 (O_1091,N_7475,N_6185);
nor UO_1092 (O_1092,N_9662,N_6433);
and UO_1093 (O_1093,N_5451,N_6139);
nand UO_1094 (O_1094,N_8535,N_6959);
or UO_1095 (O_1095,N_8693,N_9324);
nor UO_1096 (O_1096,N_6744,N_5740);
nor UO_1097 (O_1097,N_6579,N_5863);
nor UO_1098 (O_1098,N_7320,N_7862);
and UO_1099 (O_1099,N_8830,N_8717);
or UO_1100 (O_1100,N_8068,N_6751);
nor UO_1101 (O_1101,N_6255,N_6654);
and UO_1102 (O_1102,N_9690,N_9072);
or UO_1103 (O_1103,N_5958,N_6263);
and UO_1104 (O_1104,N_6414,N_9030);
or UO_1105 (O_1105,N_8333,N_7135);
nand UO_1106 (O_1106,N_8065,N_9441);
and UO_1107 (O_1107,N_5383,N_5500);
and UO_1108 (O_1108,N_5169,N_8040);
nand UO_1109 (O_1109,N_9365,N_7195);
nor UO_1110 (O_1110,N_6884,N_8474);
nor UO_1111 (O_1111,N_7021,N_9672);
nand UO_1112 (O_1112,N_5226,N_8176);
nand UO_1113 (O_1113,N_6169,N_8654);
or UO_1114 (O_1114,N_6664,N_5813);
and UO_1115 (O_1115,N_9269,N_7499);
nand UO_1116 (O_1116,N_7663,N_7534);
xnor UO_1117 (O_1117,N_6067,N_8788);
nor UO_1118 (O_1118,N_7218,N_6397);
nor UO_1119 (O_1119,N_8258,N_7030);
or UO_1120 (O_1120,N_8928,N_8896);
or UO_1121 (O_1121,N_6841,N_9479);
and UO_1122 (O_1122,N_6353,N_5540);
nand UO_1123 (O_1123,N_9754,N_8837);
or UO_1124 (O_1124,N_9533,N_8808);
nand UO_1125 (O_1125,N_5013,N_5826);
and UO_1126 (O_1126,N_8586,N_6831);
nor UO_1127 (O_1127,N_9470,N_5623);
and UO_1128 (O_1128,N_5130,N_7937);
or UO_1129 (O_1129,N_5380,N_8113);
nand UO_1130 (O_1130,N_5565,N_9078);
and UO_1131 (O_1131,N_6172,N_6718);
nand UO_1132 (O_1132,N_5432,N_6158);
nor UO_1133 (O_1133,N_8878,N_9516);
or UO_1134 (O_1134,N_9670,N_6948);
and UO_1135 (O_1135,N_9553,N_8136);
or UO_1136 (O_1136,N_5786,N_6071);
nor UO_1137 (O_1137,N_9193,N_9328);
nand UO_1138 (O_1138,N_8154,N_7379);
nor UO_1139 (O_1139,N_6720,N_7711);
nand UO_1140 (O_1140,N_5756,N_5413);
xnor UO_1141 (O_1141,N_5076,N_5239);
nor UO_1142 (O_1142,N_7553,N_9503);
nand UO_1143 (O_1143,N_5752,N_6525);
nand UO_1144 (O_1144,N_8327,N_8924);
nand UO_1145 (O_1145,N_6738,N_8706);
or UO_1146 (O_1146,N_7228,N_7704);
nor UO_1147 (O_1147,N_8092,N_7120);
and UO_1148 (O_1148,N_5603,N_5866);
nand UO_1149 (O_1149,N_9132,N_9158);
nor UO_1150 (O_1150,N_8528,N_8321);
nand UO_1151 (O_1151,N_8227,N_8226);
and UO_1152 (O_1152,N_5279,N_6316);
nor UO_1153 (O_1153,N_8120,N_7277);
nand UO_1154 (O_1154,N_7787,N_5869);
or UO_1155 (O_1155,N_6677,N_7976);
nor UO_1156 (O_1156,N_8101,N_9094);
or UO_1157 (O_1157,N_7059,N_9036);
or UO_1158 (O_1158,N_8390,N_9846);
nor UO_1159 (O_1159,N_9527,N_5838);
and UO_1160 (O_1160,N_5046,N_8503);
or UO_1161 (O_1161,N_9873,N_6964);
nand UO_1162 (O_1162,N_6534,N_7053);
nand UO_1163 (O_1163,N_6836,N_8502);
nor UO_1164 (O_1164,N_5018,N_6380);
nor UO_1165 (O_1165,N_7987,N_7521);
and UO_1166 (O_1166,N_9081,N_6364);
nor UO_1167 (O_1167,N_5557,N_6487);
nand UO_1168 (O_1168,N_7921,N_8678);
nor UO_1169 (O_1169,N_9480,N_9212);
and UO_1170 (O_1170,N_8117,N_9744);
or UO_1171 (O_1171,N_5342,N_6272);
and UO_1172 (O_1172,N_6943,N_6240);
nand UO_1173 (O_1173,N_6381,N_8888);
nand UO_1174 (O_1174,N_5337,N_6492);
nand UO_1175 (O_1175,N_5364,N_5272);
or UO_1176 (O_1176,N_7612,N_8595);
or UO_1177 (O_1177,N_8883,N_9439);
and UO_1178 (O_1178,N_5090,N_9920);
or UO_1179 (O_1179,N_9535,N_8448);
nand UO_1180 (O_1180,N_8278,N_9153);
nor UO_1181 (O_1181,N_5761,N_9306);
nor UO_1182 (O_1182,N_5918,N_9698);
or UO_1183 (O_1183,N_9619,N_6540);
nor UO_1184 (O_1184,N_6419,N_6980);
xnor UO_1185 (O_1185,N_6175,N_7952);
nand UO_1186 (O_1186,N_7950,N_8728);
or UO_1187 (O_1187,N_6306,N_6880);
or UO_1188 (O_1188,N_8609,N_7805);
or UO_1189 (O_1189,N_6219,N_5250);
nand UO_1190 (O_1190,N_7324,N_5618);
nand UO_1191 (O_1191,N_6047,N_9844);
and UO_1192 (O_1192,N_5757,N_7063);
nor UO_1193 (O_1193,N_9071,N_5612);
nor UO_1194 (O_1194,N_8359,N_8852);
nand UO_1195 (O_1195,N_7812,N_9841);
nand UO_1196 (O_1196,N_6965,N_6868);
nand UO_1197 (O_1197,N_5681,N_5170);
or UO_1198 (O_1198,N_6535,N_5324);
and UO_1199 (O_1199,N_9181,N_6486);
or UO_1200 (O_1200,N_9888,N_9509);
nand UO_1201 (O_1201,N_8054,N_5320);
nor UO_1202 (O_1202,N_9883,N_6390);
nor UO_1203 (O_1203,N_6080,N_9417);
nand UO_1204 (O_1204,N_6450,N_5887);
nor UO_1205 (O_1205,N_6086,N_5043);
and UO_1206 (O_1206,N_9825,N_8031);
nor UO_1207 (O_1207,N_8247,N_6118);
or UO_1208 (O_1208,N_5248,N_8473);
nor UO_1209 (O_1209,N_8588,N_5552);
or UO_1210 (O_1210,N_9705,N_9901);
and UO_1211 (O_1211,N_5582,N_7672);
nand UO_1212 (O_1212,N_9932,N_6454);
or UO_1213 (O_1213,N_5734,N_9207);
and UO_1214 (O_1214,N_6297,N_6942);
nand UO_1215 (O_1215,N_8395,N_8801);
or UO_1216 (O_1216,N_5925,N_5554);
or UO_1217 (O_1217,N_7746,N_6107);
or UO_1218 (O_1218,N_8398,N_8080);
nand UO_1219 (O_1219,N_5508,N_6725);
and UO_1220 (O_1220,N_9174,N_8187);
nand UO_1221 (O_1221,N_8772,N_7793);
xor UO_1222 (O_1222,N_6946,N_6367);
and UO_1223 (O_1223,N_8984,N_7171);
nand UO_1224 (O_1224,N_8741,N_7417);
nor UO_1225 (O_1225,N_5455,N_8116);
nor UO_1226 (O_1226,N_5106,N_7877);
nor UO_1227 (O_1227,N_8252,N_6229);
and UO_1228 (O_1228,N_5266,N_7391);
or UO_1229 (O_1229,N_7111,N_9549);
and UO_1230 (O_1230,N_7794,N_9937);
nor UO_1231 (O_1231,N_5267,N_8264);
nand UO_1232 (O_1232,N_8237,N_7684);
or UO_1233 (O_1233,N_5004,N_9784);
and UO_1234 (O_1234,N_9708,N_5074);
nand UO_1235 (O_1235,N_5671,N_6852);
nand UO_1236 (O_1236,N_7931,N_5798);
nor UO_1237 (O_1237,N_7674,N_8015);
and UO_1238 (O_1238,N_6225,N_9655);
and UO_1239 (O_1239,N_7441,N_5686);
or UO_1240 (O_1240,N_8220,N_6468);
and UO_1241 (O_1241,N_7536,N_9998);
or UO_1242 (O_1242,N_5993,N_5052);
and UO_1243 (O_1243,N_7358,N_7023);
or UO_1244 (O_1244,N_6607,N_5860);
nor UO_1245 (O_1245,N_6897,N_9240);
nor UO_1246 (O_1246,N_8641,N_6547);
and UO_1247 (O_1247,N_9264,N_5670);
and UO_1248 (O_1248,N_5159,N_7990);
nand UO_1249 (O_1249,N_9168,N_7491);
nor UO_1250 (O_1250,N_6574,N_5171);
nand UO_1251 (O_1251,N_7429,N_6859);
nand UO_1252 (O_1252,N_6614,N_9063);
nand UO_1253 (O_1253,N_8918,N_6820);
or UO_1254 (O_1254,N_9111,N_5956);
nor UO_1255 (O_1255,N_7770,N_7477);
nand UO_1256 (O_1256,N_7594,N_6247);
or UO_1257 (O_1257,N_5622,N_5801);
nor UO_1258 (O_1258,N_8469,N_8289);
nor UO_1259 (O_1259,N_7318,N_9915);
or UO_1260 (O_1260,N_6368,N_5939);
nor UO_1261 (O_1261,N_8505,N_8867);
and UO_1262 (O_1262,N_6742,N_6473);
nor UO_1263 (O_1263,N_8786,N_6178);
or UO_1264 (O_1264,N_6789,N_5639);
and UO_1265 (O_1265,N_9820,N_6912);
or UO_1266 (O_1266,N_7694,N_8495);
or UO_1267 (O_1267,N_9622,N_7730);
nand UO_1268 (O_1268,N_9739,N_7955);
and UO_1269 (O_1269,N_8427,N_8196);
nand UO_1270 (O_1270,N_9792,N_7232);
nor UO_1271 (O_1271,N_9946,N_8282);
nor UO_1272 (O_1272,N_9374,N_9231);
xor UO_1273 (O_1273,N_6585,N_7974);
or UO_1274 (O_1274,N_5940,N_6218);
nand UO_1275 (O_1275,N_9239,N_8951);
or UO_1276 (O_1276,N_7905,N_6109);
nor UO_1277 (O_1277,N_7611,N_7551);
or UO_1278 (O_1278,N_8462,N_6005);
and UO_1279 (O_1279,N_7275,N_5105);
and UO_1280 (O_1280,N_5409,N_7408);
nor UO_1281 (O_1281,N_7924,N_9866);
nand UO_1282 (O_1282,N_7544,N_7031);
xor UO_1283 (O_1283,N_6904,N_7132);
nor UO_1284 (O_1284,N_8151,N_6639);
or UO_1285 (O_1285,N_6630,N_5629);
nand UO_1286 (O_1286,N_5438,N_5228);
and UO_1287 (O_1287,N_8219,N_8585);
or UO_1288 (O_1288,N_6070,N_8790);
and UO_1289 (O_1289,N_5044,N_7625);
nor UO_1290 (O_1290,N_6519,N_6439);
nor UO_1291 (O_1291,N_7790,N_8224);
and UO_1292 (O_1292,N_8381,N_8343);
nand UO_1293 (O_1293,N_5889,N_9766);
nor UO_1294 (O_1294,N_9923,N_6554);
or UO_1295 (O_1295,N_9360,N_7797);
and UO_1296 (O_1296,N_8665,N_7148);
and UO_1297 (O_1297,N_7995,N_5769);
or UO_1298 (O_1298,N_8365,N_8028);
nand UO_1299 (O_1299,N_9511,N_9738);
and UO_1300 (O_1300,N_7951,N_8591);
and UO_1301 (O_1301,N_5135,N_9977);
and UO_1302 (O_1302,N_7847,N_7451);
or UO_1303 (O_1303,N_5781,N_9564);
nand UO_1304 (O_1304,N_9176,N_6589);
or UO_1305 (O_1305,N_7255,N_9635);
nor UO_1306 (O_1306,N_5335,N_8884);
nand UO_1307 (O_1307,N_8371,N_7443);
and UO_1308 (O_1308,N_7283,N_9649);
nor UO_1309 (O_1309,N_9029,N_8879);
nor UO_1310 (O_1310,N_5357,N_9056);
nand UO_1311 (O_1311,N_8606,N_6090);
or UO_1312 (O_1312,N_8292,N_6958);
or UO_1313 (O_1313,N_9650,N_5908);
nand UO_1314 (O_1314,N_6105,N_5110);
nor UO_1315 (O_1315,N_6676,N_9406);
nor UO_1316 (O_1316,N_9223,N_5282);
or UO_1317 (O_1317,N_8300,N_9628);
nor UO_1318 (O_1318,N_6315,N_5809);
nand UO_1319 (O_1319,N_9706,N_7094);
and UO_1320 (O_1320,N_9962,N_8456);
nand UO_1321 (O_1321,N_9205,N_8410);
nand UO_1322 (O_1322,N_8988,N_6895);
or UO_1323 (O_1323,N_6892,N_7971);
and UO_1324 (O_1324,N_9918,N_8524);
and UO_1325 (O_1325,N_9285,N_5075);
or UO_1326 (O_1326,N_7776,N_8311);
nor UO_1327 (O_1327,N_9726,N_7998);
and UO_1328 (O_1328,N_5504,N_6576);
or UO_1329 (O_1329,N_6420,N_7696);
nor UO_1330 (O_1330,N_8331,N_9478);
nor UO_1331 (O_1331,N_9198,N_9351);
and UO_1332 (O_1332,N_6810,N_9161);
nor UO_1333 (O_1333,N_9335,N_6084);
nand UO_1334 (O_1334,N_7942,N_6846);
nand UO_1335 (O_1335,N_7673,N_7681);
nand UO_1336 (O_1336,N_7075,N_7959);
nor UO_1337 (O_1337,N_5858,N_6098);
nor UO_1338 (O_1338,N_6648,N_5735);
and UO_1339 (O_1339,N_8614,N_8303);
nor UO_1340 (O_1340,N_6386,N_6998);
nand UO_1341 (O_1341,N_6694,N_5997);
and UO_1342 (O_1342,N_9934,N_7049);
and UO_1343 (O_1343,N_5271,N_5709);
or UO_1344 (O_1344,N_7538,N_5874);
or UO_1345 (O_1345,N_5794,N_8221);
nor UO_1346 (O_1346,N_5824,N_5027);
nor UO_1347 (O_1347,N_7365,N_8635);
nor UO_1348 (O_1348,N_8922,N_8306);
nand UO_1349 (O_1349,N_8824,N_5872);
and UO_1350 (O_1350,N_7230,N_5379);
and UO_1351 (O_1351,N_5749,N_6612);
nor UO_1352 (O_1352,N_5244,N_5415);
and UO_1353 (O_1353,N_9621,N_5209);
nand UO_1354 (O_1354,N_8210,N_9681);
and UO_1355 (O_1355,N_9714,N_6001);
or UO_1356 (O_1356,N_6732,N_6575);
nor UO_1357 (O_1357,N_6636,N_6712);
or UO_1358 (O_1358,N_9329,N_5632);
or UO_1359 (O_1359,N_6059,N_5437);
and UO_1360 (O_1360,N_7146,N_8869);
nor UO_1361 (O_1361,N_5973,N_6021);
and UO_1362 (O_1362,N_6033,N_7050);
nor UO_1363 (O_1363,N_8866,N_5932);
or UO_1364 (O_1364,N_6451,N_7598);
xor UO_1365 (O_1365,N_9234,N_9574);
nand UO_1366 (O_1366,N_8114,N_9189);
or UO_1367 (O_1367,N_6032,N_6790);
or UO_1368 (O_1368,N_7656,N_7407);
nand UO_1369 (O_1369,N_5936,N_9665);
nand UO_1370 (O_1370,N_6866,N_9556);
and UO_1371 (O_1371,N_8467,N_5598);
nand UO_1372 (O_1372,N_7830,N_5358);
and UO_1373 (O_1373,N_5986,N_5116);
and UO_1374 (O_1374,N_6385,N_7009);
nand UO_1375 (O_1375,N_5481,N_8003);
and UO_1376 (O_1376,N_8228,N_7086);
and UO_1377 (O_1377,N_8558,N_8864);
and UO_1378 (O_1378,N_9095,N_7250);
nor UO_1379 (O_1379,N_9790,N_9023);
nor UO_1380 (O_1380,N_9106,N_6522);
nor UO_1381 (O_1381,N_9689,N_5842);
or UO_1382 (O_1382,N_8159,N_7345);
and UO_1383 (O_1383,N_7024,N_8682);
nor UO_1384 (O_1384,N_5800,N_6181);
nand UO_1385 (O_1385,N_7295,N_5543);
and UO_1386 (O_1386,N_6022,N_9380);
nand UO_1387 (O_1387,N_7831,N_5751);
nand UO_1388 (O_1388,N_7127,N_6348);
and UO_1389 (O_1389,N_9919,N_7394);
or UO_1390 (O_1390,N_5003,N_5583);
nand UO_1391 (O_1391,N_5947,N_5758);
nand UO_1392 (O_1392,N_8177,N_8006);
nand UO_1393 (O_1393,N_8670,N_6210);
nand UO_1394 (O_1394,N_8397,N_8754);
and UO_1395 (O_1395,N_8175,N_6066);
nor UO_1396 (O_1396,N_9378,N_7956);
or UO_1397 (O_1397,N_8207,N_6013);
or UO_1398 (O_1398,N_8344,N_6558);
nand UO_1399 (O_1399,N_8843,N_6871);
nand UO_1400 (O_1400,N_7048,N_8854);
nand UO_1401 (O_1401,N_6689,N_9829);
and UO_1402 (O_1402,N_9752,N_6640);
or UO_1403 (O_1403,N_5699,N_5542);
or UO_1404 (O_1404,N_9321,N_6256);
and UO_1405 (O_1405,N_6707,N_7479);
nand UO_1406 (O_1406,N_7671,N_5992);
nand UO_1407 (O_1407,N_5382,N_5104);
nand UO_1408 (O_1408,N_7252,N_6678);
nand UO_1409 (O_1409,N_5312,N_7620);
nand UO_1410 (O_1410,N_7778,N_5536);
nor UO_1411 (O_1411,N_6613,N_6730);
nand UO_1412 (O_1412,N_7842,N_5329);
nor UO_1413 (O_1413,N_7134,N_9583);
or UO_1414 (O_1414,N_9484,N_6037);
nand UO_1415 (O_1415,N_9472,N_7928);
or UO_1416 (O_1416,N_8405,N_6538);
and UO_1417 (O_1417,N_9477,N_6191);
nor UO_1418 (O_1418,N_7015,N_9277);
and UO_1419 (O_1419,N_9450,N_8049);
nor UO_1420 (O_1420,N_6125,N_8789);
nand UO_1421 (O_1421,N_8118,N_6514);
nor UO_1422 (O_1422,N_7226,N_7321);
and UO_1423 (O_1423,N_7406,N_8513);
nand UO_1424 (O_1424,N_7912,N_8687);
nand UO_1425 (O_1425,N_9089,N_6541);
and UO_1426 (O_1426,N_5899,N_6432);
or UO_1427 (O_1427,N_5854,N_9145);
or UO_1428 (O_1428,N_5424,N_5378);
nor UO_1429 (O_1429,N_8845,N_9416);
nor UO_1430 (O_1430,N_5185,N_5011);
and UO_1431 (O_1431,N_9279,N_9909);
nand UO_1432 (O_1432,N_5763,N_9684);
nand UO_1433 (O_1433,N_9270,N_9104);
nor UO_1434 (O_1434,N_8141,N_7130);
and UO_1435 (O_1435,N_6779,N_6981);
nor UO_1436 (O_1436,N_6580,N_5290);
or UO_1437 (O_1437,N_7355,N_8834);
or UO_1438 (O_1438,N_7442,N_6017);
or UO_1439 (O_1439,N_7088,N_9092);
nand UO_1440 (O_1440,N_5283,N_7630);
and UO_1441 (O_1441,N_7271,N_9488);
nand UO_1442 (O_1442,N_8514,N_7118);
or UO_1443 (O_1443,N_6925,N_8903);
or UO_1444 (O_1444,N_6951,N_6455);
and UO_1445 (O_1445,N_6629,N_9614);
or UO_1446 (O_1446,N_6289,N_8806);
and UO_1447 (O_1447,N_8391,N_9252);
or UO_1448 (O_1448,N_8853,N_5867);
nand UO_1449 (O_1449,N_7906,N_5155);
nand UO_1450 (O_1450,N_7136,N_5398);
nor UO_1451 (O_1451,N_9099,N_6205);
nor UO_1452 (O_1452,N_9867,N_5047);
and UO_1453 (O_1453,N_5435,N_8582);
and UO_1454 (O_1454,N_8527,N_8358);
nand UO_1455 (O_1455,N_9297,N_8342);
nor UO_1456 (O_1456,N_6872,N_5951);
nor UO_1457 (O_1457,N_5216,N_6308);
and UO_1458 (O_1458,N_7832,N_7729);
nand UO_1459 (O_1459,N_7601,N_8035);
or UO_1460 (O_1460,N_8363,N_7032);
nor UO_1461 (O_1461,N_6362,N_7511);
nor UO_1462 (O_1462,N_5411,N_6544);
nand UO_1463 (O_1463,N_6278,N_5099);
nand UO_1464 (O_1464,N_5849,N_7007);
or UO_1465 (O_1465,N_9133,N_7973);
or UO_1466 (O_1466,N_7573,N_8245);
nor UO_1467 (O_1467,N_6038,N_9043);
or UO_1468 (O_1468,N_5776,N_8084);
and UO_1469 (O_1469,N_7478,N_7641);
and UO_1470 (O_1470,N_8583,N_7006);
or UO_1471 (O_1471,N_5222,N_6096);
nand UO_1472 (O_1472,N_5962,N_6914);
nor UO_1473 (O_1473,N_6167,N_5523);
or UO_1474 (O_1474,N_6009,N_9123);
or UO_1475 (O_1475,N_8787,N_9446);
nor UO_1476 (O_1476,N_9258,N_9798);
and UO_1477 (O_1477,N_7899,N_9460);
or UO_1478 (O_1478,N_9908,N_7497);
and UO_1479 (O_1479,N_5280,N_9453);
or UO_1480 (O_1480,N_6373,N_5381);
and UO_1481 (O_1481,N_9904,N_7769);
nor UO_1482 (O_1482,N_8798,N_5546);
nand UO_1483 (O_1483,N_6494,N_8946);
or UO_1484 (O_1484,N_8916,N_6073);
nand UO_1485 (O_1485,N_5948,N_7448);
nand UO_1486 (O_1486,N_9666,N_5485);
nor UO_1487 (O_1487,N_9581,N_9210);
and UO_1488 (O_1488,N_7501,N_8105);
and UO_1489 (O_1489,N_7903,N_7579);
nand UO_1490 (O_1490,N_6830,N_5871);
nand UO_1491 (O_1491,N_5733,N_6775);
nand UO_1492 (O_1492,N_6324,N_8731);
xor UO_1493 (O_1493,N_9912,N_8256);
or UO_1494 (O_1494,N_6552,N_9600);
nor UO_1495 (O_1495,N_6896,N_6422);
nand UO_1496 (O_1496,N_8383,N_9521);
or UO_1497 (O_1497,N_6101,N_6212);
or UO_1498 (O_1498,N_5285,N_5405);
nor UO_1499 (O_1499,N_6865,N_5790);
endmodule