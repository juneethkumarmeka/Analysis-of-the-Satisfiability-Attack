module basic_1500_15000_2000_5_levels_1xor_1(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999;
nand U0 (N_0,In_1053,In_1319);
and U1 (N_1,In_1123,In_1455);
and U2 (N_2,In_848,In_958);
nor U3 (N_3,In_1449,In_1022);
nand U4 (N_4,In_1441,In_1120);
nand U5 (N_5,In_130,In_1219);
nor U6 (N_6,In_80,In_676);
or U7 (N_7,In_1097,In_452);
nand U8 (N_8,In_77,In_1253);
or U9 (N_9,In_497,In_1045);
nor U10 (N_10,In_1243,In_793);
nor U11 (N_11,In_1408,In_1018);
or U12 (N_12,In_44,In_121);
nor U13 (N_13,In_562,In_720);
nand U14 (N_14,In_237,In_1397);
nor U15 (N_15,In_1148,In_1398);
nand U16 (N_16,In_964,In_1459);
nor U17 (N_17,In_253,In_525);
and U18 (N_18,In_565,In_1347);
xnor U19 (N_19,In_470,In_1165);
nor U20 (N_20,In_1341,In_630);
and U21 (N_21,In_1412,In_1021);
or U22 (N_22,In_750,In_193);
nand U23 (N_23,In_297,In_409);
nor U24 (N_24,In_1477,In_1247);
and U25 (N_25,In_1246,In_1060);
and U26 (N_26,In_1199,In_415);
or U27 (N_27,In_126,In_191);
or U28 (N_28,In_1065,In_941);
nand U29 (N_29,In_263,In_312);
or U30 (N_30,In_1089,In_187);
or U31 (N_31,In_891,In_867);
xor U32 (N_32,In_151,In_1350);
or U33 (N_33,In_384,In_56);
or U34 (N_34,In_1265,In_524);
nor U35 (N_35,In_257,In_117);
nor U36 (N_36,In_267,In_337);
nand U37 (N_37,In_1187,In_291);
or U38 (N_38,In_1016,In_1365);
nor U39 (N_39,In_316,In_731);
or U40 (N_40,In_1302,In_993);
and U41 (N_41,In_490,In_785);
and U42 (N_42,In_535,In_655);
nand U43 (N_43,In_498,In_1234);
or U44 (N_44,In_325,In_275);
nor U45 (N_45,In_102,In_840);
nand U46 (N_46,In_310,In_741);
or U47 (N_47,In_1289,In_134);
and U48 (N_48,In_603,In_38);
or U49 (N_49,In_1076,In_26);
and U50 (N_50,In_1332,In_1066);
nand U51 (N_51,In_1027,In_335);
or U52 (N_52,In_1079,In_1049);
or U53 (N_53,In_206,In_854);
nor U54 (N_54,In_919,In_296);
nand U55 (N_55,In_268,In_1117);
and U56 (N_56,In_1404,In_1254);
and U57 (N_57,In_737,In_1370);
nor U58 (N_58,In_46,In_1450);
nor U59 (N_59,In_601,In_1196);
and U60 (N_60,In_13,In_1036);
and U61 (N_61,In_120,In_1447);
or U62 (N_62,In_683,In_903);
nor U63 (N_63,In_314,In_342);
nor U64 (N_64,In_155,In_1373);
nand U65 (N_65,In_186,In_775);
or U66 (N_66,In_1485,In_22);
nand U67 (N_67,In_114,In_899);
or U68 (N_68,In_236,In_1479);
or U69 (N_69,In_1340,In_1052);
nor U70 (N_70,In_1285,In_625);
nor U71 (N_71,In_1106,In_256);
nand U72 (N_72,In_177,In_241);
and U73 (N_73,In_823,In_1180);
nand U74 (N_74,In_1236,In_507);
nand U75 (N_75,In_907,In_397);
nor U76 (N_76,In_1181,In_512);
nor U77 (N_77,In_154,In_961);
xor U78 (N_78,In_135,In_1394);
and U79 (N_79,In_1420,In_1354);
and U80 (N_80,In_1034,In_1393);
nor U81 (N_81,In_1282,In_1040);
or U82 (N_82,In_363,In_650);
and U83 (N_83,In_804,In_1058);
or U84 (N_84,In_707,In_1290);
and U85 (N_85,In_617,In_230);
nor U86 (N_86,In_349,In_1328);
nand U87 (N_87,In_560,In_53);
nand U88 (N_88,In_833,In_500);
and U89 (N_89,In_588,In_534);
nor U90 (N_90,In_1382,In_1320);
and U91 (N_91,In_566,In_887);
nor U92 (N_92,In_718,In_1258);
nor U93 (N_93,In_865,In_1316);
and U94 (N_94,In_381,In_19);
or U95 (N_95,In_940,In_1272);
or U96 (N_96,In_1407,In_111);
nor U97 (N_97,In_776,In_311);
nand U98 (N_98,In_1466,In_1442);
and U99 (N_99,In_320,In_675);
nand U100 (N_100,In_1378,In_1233);
and U101 (N_101,In_1464,In_298);
or U102 (N_102,In_678,In_165);
or U103 (N_103,In_686,In_465);
nand U104 (N_104,In_491,In_1077);
and U105 (N_105,In_1200,In_1020);
nand U106 (N_106,In_845,In_736);
or U107 (N_107,In_1298,In_289);
nor U108 (N_108,In_602,In_351);
and U109 (N_109,In_223,In_1114);
nor U110 (N_110,In_450,In_1405);
nor U111 (N_111,In_133,In_423);
and U112 (N_112,In_233,In_668);
nor U113 (N_113,In_1151,In_1264);
and U114 (N_114,In_406,In_1000);
nand U115 (N_115,In_996,In_1164);
or U116 (N_116,In_1483,In_172);
nand U117 (N_117,In_1379,In_835);
nand U118 (N_118,In_1067,In_375);
nor U119 (N_119,In_986,In_1498);
or U120 (N_120,In_1299,In_471);
and U121 (N_121,In_369,In_439);
and U122 (N_122,In_510,In_136);
and U123 (N_123,In_1063,In_331);
nor U124 (N_124,In_364,In_382);
nor U125 (N_125,In_182,In_1166);
nand U126 (N_126,In_112,In_677);
nor U127 (N_127,In_921,In_59);
or U128 (N_128,In_266,In_95);
nor U129 (N_129,In_511,In_561);
nand U130 (N_130,In_672,In_1396);
nand U131 (N_131,In_569,In_1057);
nand U132 (N_132,In_383,In_1140);
or U133 (N_133,In_248,In_299);
and U134 (N_134,In_11,In_635);
nor U135 (N_135,In_544,In_1098);
and U136 (N_136,In_1,In_5);
nand U137 (N_137,In_445,In_1071);
nand U138 (N_138,In_1336,In_73);
and U139 (N_139,In_710,In_679);
nor U140 (N_140,In_24,In_777);
nand U141 (N_141,In_1143,In_122);
or U142 (N_142,In_817,In_189);
nand U143 (N_143,In_1222,In_1383);
or U144 (N_144,In_596,In_540);
and U145 (N_145,In_25,In_956);
or U146 (N_146,In_1361,In_340);
nand U147 (N_147,In_1059,In_481);
or U148 (N_148,In_1260,In_417);
and U149 (N_149,In_1266,In_1352);
nor U150 (N_150,In_766,In_391);
and U151 (N_151,In_579,In_82);
xnor U152 (N_152,In_324,In_702);
nor U153 (N_153,In_425,In_781);
nand U154 (N_154,In_242,In_1314);
nand U155 (N_155,In_1287,In_100);
xnor U156 (N_156,In_938,In_945);
nor U157 (N_157,In_12,In_502);
or U158 (N_158,In_692,In_664);
nor U159 (N_159,In_606,In_492);
and U160 (N_160,In_265,In_438);
and U161 (N_161,In_219,In_179);
nand U162 (N_162,In_691,In_515);
or U163 (N_163,In_770,In_15);
or U164 (N_164,In_1101,In_1342);
nor U165 (N_165,In_499,In_453);
or U166 (N_166,In_942,In_106);
and U167 (N_167,In_1154,In_1168);
and U168 (N_168,In_1488,In_254);
or U169 (N_169,In_764,In_605);
and U170 (N_170,In_1139,In_478);
nor U171 (N_171,In_173,In_8);
nor U172 (N_172,In_123,In_505);
and U173 (N_173,In_380,In_1118);
and U174 (N_174,In_1232,In_568);
and U175 (N_175,In_595,In_1113);
nor U176 (N_176,In_1482,In_140);
xnor U177 (N_177,In_751,In_1146);
nand U178 (N_178,In_1309,In_831);
and U179 (N_179,In_763,In_1192);
nor U180 (N_180,In_727,In_604);
nor U181 (N_181,In_794,In_926);
or U182 (N_182,In_1388,In_1267);
or U183 (N_183,In_559,In_98);
and U184 (N_184,In_728,In_713);
and U185 (N_185,In_378,In_1155);
nand U186 (N_186,In_101,In_460);
or U187 (N_187,In_846,In_1206);
nor U188 (N_188,In_284,In_698);
or U189 (N_189,In_488,In_1262);
nor U190 (N_190,In_489,In_530);
or U191 (N_191,In_730,In_959);
nor U192 (N_192,In_700,In_1014);
and U193 (N_193,In_957,In_113);
nor U194 (N_194,In_935,In_440);
and U195 (N_195,In_1300,In_552);
nand U196 (N_196,In_771,In_851);
or U197 (N_197,In_449,In_1417);
nand U198 (N_198,In_924,In_575);
and U199 (N_199,In_1297,In_1241);
or U200 (N_200,In_322,In_1346);
nor U201 (N_201,In_564,In_828);
and U202 (N_202,In_124,In_580);
or U203 (N_203,In_1434,In_1137);
nand U204 (N_204,In_212,In_1339);
nor U205 (N_205,In_1499,In_1338);
nand U206 (N_206,In_243,In_14);
nor U207 (N_207,In_871,In_558);
or U208 (N_208,In_1132,In_317);
or U209 (N_209,In_1303,In_1245);
and U210 (N_210,In_1252,In_612);
and U211 (N_211,In_570,In_647);
nand U212 (N_212,In_795,In_772);
xnor U213 (N_213,In_295,In_859);
nor U214 (N_214,In_939,In_832);
nand U215 (N_215,In_301,In_600);
nor U216 (N_216,In_1448,In_207);
or U217 (N_217,In_1472,In_79);
and U218 (N_218,In_66,In_721);
nand U219 (N_219,In_1223,In_1431);
nor U220 (N_220,In_799,In_900);
nand U221 (N_221,In_767,In_873);
nor U222 (N_222,In_894,In_103);
and U223 (N_223,In_387,In_1446);
or U224 (N_224,In_508,In_1463);
or U225 (N_225,In_598,In_318);
nand U226 (N_226,In_856,In_1322);
and U227 (N_227,In_1047,In_674);
or U228 (N_228,In_834,In_156);
or U229 (N_229,In_1145,In_567);
nand U230 (N_230,In_537,In_980);
and U231 (N_231,In_1011,In_27);
and U232 (N_232,In_1153,In_461);
or U233 (N_233,In_1451,In_620);
nand U234 (N_234,In_1366,In_180);
nor U235 (N_235,In_673,In_1315);
nand U236 (N_236,In_222,In_214);
nand U237 (N_237,In_695,In_656);
and U238 (N_238,In_1104,In_1188);
and U239 (N_239,In_780,In_487);
nand U240 (N_240,In_687,In_472);
nand U241 (N_241,In_1471,In_1134);
or U242 (N_242,In_755,In_1013);
nand U243 (N_243,In_71,In_348);
and U244 (N_244,In_1390,In_1185);
or U245 (N_245,In_1017,In_354);
and U246 (N_246,In_352,In_838);
nor U247 (N_247,In_994,In_1128);
nand U248 (N_248,In_626,In_1116);
and U249 (N_249,In_1093,In_110);
or U250 (N_250,In_23,In_43);
nor U251 (N_251,In_1368,In_979);
and U252 (N_252,In_1364,In_395);
and U253 (N_253,In_158,In_809);
or U254 (N_254,In_792,In_609);
nand U255 (N_255,In_1456,In_1226);
and U256 (N_256,In_1130,In_424);
nor U257 (N_257,In_593,In_195);
nor U258 (N_258,In_1046,In_1306);
and U259 (N_259,In_473,In_629);
or U260 (N_260,In_506,In_1371);
nor U261 (N_261,In_693,In_1411);
nand U262 (N_262,In_1278,In_141);
nand U263 (N_263,In_1227,In_1028);
or U264 (N_264,In_1475,In_1268);
and U265 (N_265,In_334,In_85);
nand U266 (N_266,In_495,In_662);
or U267 (N_267,In_878,In_270);
nor U268 (N_268,In_1119,In_345);
and U269 (N_269,In_261,In_174);
and U270 (N_270,In_1248,In_282);
or U271 (N_271,In_213,In_1044);
nand U272 (N_272,In_479,In_716);
nand U273 (N_273,In_533,In_60);
and U274 (N_274,In_818,In_408);
and U275 (N_275,In_105,In_426);
or U276 (N_276,In_1269,In_1062);
or U277 (N_277,In_1457,In_1279);
and U278 (N_278,In_294,In_773);
and U279 (N_279,In_84,In_1088);
or U280 (N_280,In_1492,In_1129);
nor U281 (N_281,In_1194,In_1392);
or U282 (N_282,In_51,In_714);
nand U283 (N_283,In_654,In_285);
and U284 (N_284,In_368,In_538);
or U285 (N_285,In_1176,In_614);
and U286 (N_286,In_874,In_1184);
and U287 (N_287,In_661,In_861);
or U288 (N_288,In_463,In_176);
nor U289 (N_289,In_246,In_16);
or U290 (N_290,In_1374,In_928);
xnor U291 (N_291,In_974,In_347);
and U292 (N_292,In_45,In_1249);
or U293 (N_293,In_1144,In_912);
and U294 (N_294,In_476,In_1256);
and U295 (N_295,In_1286,In_247);
nor U296 (N_296,In_1231,In_125);
and U297 (N_297,In_1377,In_1075);
or U298 (N_298,In_1197,In_1074);
nand U299 (N_299,In_684,In_91);
nor U300 (N_300,In_1109,In_509);
nand U301 (N_301,In_144,In_875);
nor U302 (N_302,In_868,In_201);
nand U303 (N_303,In_1344,In_1102);
and U304 (N_304,In_1478,In_658);
nor U305 (N_305,In_469,In_1461);
nand U306 (N_306,In_1318,In_797);
or U307 (N_307,In_493,In_1462);
and U308 (N_308,In_1147,In_1195);
nand U309 (N_309,In_843,In_951);
or U310 (N_310,In_379,In_215);
or U311 (N_311,In_644,In_597);
or U312 (N_312,In_402,In_1133);
nor U313 (N_313,In_1413,In_549);
nor U314 (N_314,In_362,In_1415);
nand U315 (N_315,In_1201,In_902);
and U316 (N_316,In_960,In_1325);
nand U317 (N_317,In_769,In_1496);
or U318 (N_318,In_467,In_358);
and U319 (N_319,In_1112,In_1096);
nand U320 (N_320,In_396,In_1418);
or U321 (N_321,In_639,In_343);
and U322 (N_322,In_883,In_1351);
nor U323 (N_323,In_985,In_705);
and U324 (N_324,In_264,In_286);
nor U325 (N_325,In_1032,In_738);
nor U326 (N_326,In_1242,In_610);
nor U327 (N_327,In_401,In_962);
or U328 (N_328,In_968,In_376);
nand U329 (N_329,In_997,In_782);
or U330 (N_330,In_455,In_701);
or U331 (N_331,In_1141,In_587);
nand U332 (N_332,In_860,In_1427);
nor U333 (N_333,In_870,In_55);
nand U334 (N_334,In_866,In_966);
nor U335 (N_335,In_1082,In_1080);
or U336 (N_336,In_836,In_518);
and U337 (N_337,In_313,In_734);
or U338 (N_338,In_231,In_1476);
nand U339 (N_339,In_594,In_64);
and U340 (N_340,In_1438,In_385);
nand U341 (N_341,In_1326,In_815);
or U342 (N_342,In_1384,In_39);
or U343 (N_343,In_21,In_1291);
or U344 (N_344,In_258,In_1225);
nand U345 (N_345,In_578,In_1095);
and U346 (N_346,In_234,In_1470);
nand U347 (N_347,In_404,In_72);
nand U348 (N_348,In_885,In_1183);
or U349 (N_349,In_740,In_1257);
nand U350 (N_350,In_539,In_227);
nor U351 (N_351,In_753,In_709);
and U352 (N_352,In_589,In_858);
and U353 (N_353,In_1419,In_480);
nor U354 (N_354,In_555,In_447);
nor U355 (N_355,In_1048,In_955);
nor U356 (N_356,In_1310,In_657);
or U357 (N_357,In_1235,In_735);
or U358 (N_358,In_855,In_880);
nand U359 (N_359,In_1171,In_826);
nor U360 (N_360,In_431,In_1167);
nand U361 (N_361,In_1142,In_290);
and U362 (N_362,In_882,In_1426);
and U363 (N_363,In_1004,In_1386);
nor U364 (N_364,In_1400,In_143);
nor U365 (N_365,In_1280,In_315);
nor U366 (N_366,In_359,In_1073);
nor U367 (N_367,In_269,In_287);
or U368 (N_368,In_58,In_666);
or U369 (N_369,In_896,In_681);
and U370 (N_370,In_171,In_631);
nand U371 (N_371,In_969,In_228);
and U372 (N_372,In_1432,In_576);
and U373 (N_373,In_30,In_905);
nor U374 (N_374,In_392,In_571);
nand U375 (N_375,In_305,In_821);
and U376 (N_376,In_1409,In_618);
nand U377 (N_377,In_1440,In_699);
nor U378 (N_378,In_1439,In_1281);
nor U379 (N_379,In_330,In_982);
and U380 (N_380,In_200,In_138);
or U381 (N_381,In_585,In_1375);
nor U382 (N_382,In_532,In_1162);
or U383 (N_383,In_167,In_1480);
or U384 (N_384,In_1465,In_1061);
xor U385 (N_385,In_279,In_262);
nand U386 (N_386,In_1138,In_18);
and U387 (N_387,In_1295,In_806);
nand U388 (N_388,In_554,In_1433);
nand U389 (N_389,In_947,In_965);
and U390 (N_390,In_1007,In_590);
and U391 (N_391,In_1209,In_1015);
or U392 (N_392,In_178,In_1072);
nand U393 (N_393,In_468,In_844);
nand U394 (N_394,In_872,In_1178);
and U395 (N_395,In_1395,In_967);
and U396 (N_396,In_1251,In_1237);
or U397 (N_397,In_99,In_104);
nor U398 (N_398,In_436,In_162);
nand U399 (N_399,In_685,In_733);
or U400 (N_400,In_1399,In_1213);
and U401 (N_401,In_743,In_688);
xnor U402 (N_402,In_943,In_723);
nor U403 (N_403,In_157,In_474);
and U404 (N_404,In_628,In_7);
nand U405 (N_405,In_542,In_749);
nand U406 (N_406,In_801,In_332);
and U407 (N_407,In_759,In_170);
nand U408 (N_408,In_852,In_1430);
and U409 (N_409,In_527,In_147);
nand U410 (N_410,In_652,In_280);
nand U411 (N_411,In_633,In_403);
or U412 (N_412,In_169,In_520);
nand U413 (N_413,In_811,In_198);
nor U414 (N_414,In_1026,In_669);
and U415 (N_415,In_459,In_249);
and U416 (N_416,In_194,In_646);
or U417 (N_417,In_37,In_922);
and U418 (N_418,In_483,In_1308);
nor U419 (N_419,In_235,In_67);
nor U420 (N_420,In_485,In_1064);
nand U421 (N_421,In_1008,In_1050);
and U422 (N_422,In_107,In_1042);
xor U423 (N_423,In_784,In_820);
or U424 (N_424,In_20,In_1038);
or U425 (N_425,In_128,In_1068);
or U426 (N_426,In_1169,In_341);
nand U427 (N_427,In_886,In_1103);
nor U428 (N_428,In_192,In_703);
and U429 (N_429,In_33,In_225);
or U430 (N_430,In_153,In_999);
xor U431 (N_431,In_1131,In_184);
nand U432 (N_432,In_87,In_909);
and U433 (N_433,In_197,In_950);
nand U434 (N_434,In_1292,In_803);
nand U435 (N_435,In_1255,In_726);
nand U436 (N_436,In_9,In_1311);
and U437 (N_437,In_627,In_1321);
nor U438 (N_438,In_747,In_1039);
nand U439 (N_439,In_205,In_758);
nor U440 (N_440,In_1406,In_88);
nand U441 (N_441,In_1170,In_484);
or U442 (N_442,In_188,In_790);
nor U443 (N_443,In_1150,In_446);
nand U444 (N_444,In_1220,In_971);
or U445 (N_445,In_798,In_339);
nor U446 (N_446,In_411,In_190);
and U447 (N_447,In_1244,In_869);
nor U448 (N_448,In_812,In_150);
nand U449 (N_449,In_1469,In_1274);
nor U450 (N_450,In_889,In_76);
nand U451 (N_451,In_127,In_1273);
and U452 (N_452,In_94,In_410);
nand U453 (N_453,In_218,In_970);
and U454 (N_454,In_934,In_637);
and U455 (N_455,In_591,In_304);
nand U456 (N_456,In_1362,In_464);
nand U457 (N_457,In_1041,In_1259);
nand U458 (N_458,In_309,In_857);
nand U459 (N_459,In_1452,In_917);
nor U460 (N_460,In_910,In_1084);
or U461 (N_461,In_152,In_659);
and U462 (N_462,In_1006,In_1107);
nor U463 (N_463,In_245,In_665);
nand U464 (N_464,In_884,In_90);
or U465 (N_465,In_338,In_429);
or U466 (N_466,In_390,In_422);
and U467 (N_467,In_1163,In_1161);
nand U468 (N_468,In_642,In_582);
nor U469 (N_469,In_1468,In_41);
nand U470 (N_470,In_789,In_199);
nand U471 (N_471,In_1005,In_414);
nand U472 (N_472,In_1182,In_1435);
nor U473 (N_473,In_220,In_1228);
and U474 (N_474,In_161,In_17);
nand U475 (N_475,In_42,In_1177);
or U476 (N_476,In_521,In_901);
nand U477 (N_477,In_768,In_1402);
nor U478 (N_478,In_2,In_448);
and U479 (N_479,In_466,In_432);
nor U480 (N_480,In_877,In_779);
xor U481 (N_481,In_1312,In_407);
or U482 (N_482,In_645,In_1085);
or U483 (N_483,In_1090,In_78);
and U484 (N_484,In_1410,In_1422);
or U485 (N_485,In_1356,In_388);
nand U486 (N_486,In_636,In_451);
nand U487 (N_487,In_54,In_1250);
nand U488 (N_488,In_1296,In_259);
nor U489 (N_489,In_302,In_355);
nand U490 (N_490,In_948,In_791);
nor U491 (N_491,In_708,In_1385);
or U492 (N_492,In_1174,In_813);
nor U493 (N_493,In_1494,In_118);
and U494 (N_494,In_952,In_514);
and U495 (N_495,In_1051,In_300);
nand U496 (N_496,In_306,In_386);
nand U497 (N_497,In_1111,In_739);
and U498 (N_498,In_166,In_973);
nand U499 (N_499,In_1056,In_1493);
nand U500 (N_500,In_944,In_208);
nor U501 (N_501,In_1349,In_573);
nor U502 (N_502,In_1126,In_1473);
or U503 (N_503,In_1158,In_1214);
or U504 (N_504,In_689,In_86);
and U505 (N_505,In_913,In_357);
nand U506 (N_506,In_932,In_221);
nor U507 (N_507,In_1424,In_168);
and U508 (N_508,In_904,In_550);
nand U509 (N_509,In_667,In_1453);
nor U510 (N_510,In_1108,In_1348);
and U511 (N_511,In_802,In_931);
nand U512 (N_512,In_816,In_1009);
or U513 (N_513,In_1087,In_1094);
and U514 (N_514,In_496,In_1210);
nor U515 (N_515,In_839,In_372);
nand U516 (N_516,In_1202,In_1486);
nand U517 (N_517,In_563,In_526);
and U518 (N_518,In_651,In_240);
or U519 (N_519,In_760,In_216);
nand U520 (N_520,In_336,In_1327);
or U521 (N_521,In_1389,In_273);
nand U522 (N_522,In_599,In_1156);
nand U523 (N_523,In_1125,In_10);
nand U524 (N_524,In_1191,In_454);
xor U525 (N_525,In_303,In_1324);
or U526 (N_526,In_1305,In_978);
or U527 (N_527,In_762,In_96);
and U528 (N_528,In_954,In_584);
or U529 (N_529,In_1460,In_517);
nor U530 (N_530,In_987,In_946);
or U531 (N_531,In_293,In_1497);
nor U532 (N_532,In_853,In_1127);
nand U533 (N_533,In_3,In_308);
and U534 (N_534,In_1122,In_641);
nor U535 (N_535,In_371,In_1270);
and U536 (N_536,In_1293,In_433);
nor U537 (N_537,In_732,In_437);
nand U538 (N_538,In_1301,In_319);
and U539 (N_539,In_1335,In_1261);
nor U540 (N_540,In_906,In_748);
or U541 (N_541,In_995,In_1224);
nor U542 (N_542,In_70,In_1345);
or U543 (N_543,In_373,In_1491);
xor U544 (N_544,In_1193,In_837);
nand U545 (N_545,In_796,In_890);
nor U546 (N_546,In_81,In_185);
nor U547 (N_547,In_634,In_1414);
nand U548 (N_548,In_34,In_613);
and U549 (N_549,In_788,In_1437);
nor U550 (N_550,In_260,In_494);
and U551 (N_551,In_1221,In_892);
or U552 (N_552,In_711,In_653);
or U553 (N_553,In_35,In_47);
and U554 (N_554,In_288,In_1179);
nand U555 (N_555,In_1115,In_31);
nand U556 (N_556,In_250,In_546);
or U557 (N_557,In_327,In_210);
or U558 (N_558,In_1358,In_572);
nor U559 (N_559,In_984,In_1190);
or U560 (N_560,In_536,In_211);
or U561 (N_561,In_501,In_1330);
and U562 (N_562,In_405,In_89);
nor U563 (N_563,In_807,In_671);
nand U564 (N_564,In_774,In_643);
nor U565 (N_565,In_529,In_462);
and U566 (N_566,In_988,In_949);
and U567 (N_567,In_420,In_927);
nor U568 (N_568,In_29,In_83);
nand U569 (N_569,In_616,In_975);
nand U570 (N_570,In_523,In_930);
and U571 (N_571,In_516,In_648);
nor U572 (N_572,In_757,In_367);
or U573 (N_573,In_841,In_93);
nor U574 (N_574,In_1333,In_160);
nor U575 (N_575,In_366,In_911);
or U576 (N_576,In_825,In_933);
or U577 (N_577,In_649,In_1238);
nor U578 (N_578,In_1230,In_1489);
and U579 (N_579,In_40,In_1484);
nand U580 (N_580,In_1100,In_992);
nand U581 (N_581,In_283,In_1331);
nand U582 (N_582,In_1217,In_6);
or U583 (N_583,In_74,In_547);
or U584 (N_584,In_204,In_808);
and U585 (N_585,In_864,In_830);
nand U586 (N_586,In_418,In_1323);
nor U587 (N_587,In_255,In_1070);
nand U588 (N_588,In_914,In_232);
nand U589 (N_589,In_48,In_1329);
or U590 (N_590,In_660,In_346);
nand U591 (N_591,In_1211,In_805);
or U592 (N_592,In_1172,In_435);
and U593 (N_593,In_430,In_531);
nor U594 (N_594,In_953,In_1454);
and U595 (N_595,In_1421,In_1033);
nor U596 (N_596,In_413,In_1229);
nor U597 (N_597,In_1294,In_1029);
nand U598 (N_598,In_202,In_360);
nand U599 (N_599,In_196,In_923);
and U600 (N_600,In_756,In_1086);
nand U601 (N_601,In_1376,In_1423);
nor U602 (N_602,In_990,In_482);
and U603 (N_603,In_963,In_1010);
nand U604 (N_604,In_742,In_75);
or U605 (N_605,In_139,In_1110);
nor U606 (N_606,In_356,In_203);
or U607 (N_607,In_1444,In_109);
xor U608 (N_608,In_209,In_183);
or U609 (N_609,In_1436,In_765);
nand U610 (N_610,In_1490,In_754);
nor U611 (N_611,In_146,In_1288);
or U612 (N_612,In_389,In_52);
nor U613 (N_613,In_1239,In_1391);
nand U614 (N_614,In_581,In_722);
nand U615 (N_615,In_1069,In_553);
nand U616 (N_616,In_778,In_876);
and U617 (N_617,In_361,In_374);
nand U618 (N_618,In_274,In_682);
and U619 (N_619,In_814,In_1481);
or U620 (N_620,In_329,In_1189);
nand U621 (N_621,In_442,In_1078);
nor U622 (N_622,In_244,In_670);
nand U623 (N_623,In_1055,In_632);
nor U624 (N_624,In_1360,In_1208);
nand U625 (N_625,In_624,In_925);
and U626 (N_626,In_217,In_68);
or U627 (N_627,In_292,In_719);
nor U628 (N_628,In_281,In_1428);
nor U629 (N_629,In_323,In_393);
or U630 (N_630,In_849,In_1002);
nand U631 (N_631,In_1207,In_1307);
nor U632 (N_632,In_444,In_937);
nor U633 (N_633,In_800,In_1212);
nor U634 (N_634,In_456,In_1467);
nand U635 (N_635,In_1043,In_1263);
nor U636 (N_636,In_862,In_706);
and U637 (N_637,In_1275,In_50);
or U638 (N_638,In_619,In_1175);
or U639 (N_639,In_746,In_989);
nand U640 (N_640,In_1024,In_1277);
nor U641 (N_641,In_513,In_725);
or U642 (N_642,In_1276,In_1487);
or U643 (N_643,In_1019,In_920);
or U644 (N_644,In_847,In_1136);
or U645 (N_645,In_129,In_557);
nand U646 (N_646,In_119,In_421);
or U647 (N_647,In_1359,In_1380);
or U648 (N_648,In_1157,In_522);
or U649 (N_649,In_1204,In_271);
and U650 (N_650,In_419,In_551);
and U651 (N_651,In_694,In_224);
and U652 (N_652,In_724,In_434);
xnor U653 (N_653,In_1023,In_1198);
or U654 (N_654,In_583,In_377);
nor U655 (N_655,In_1001,In_1240);
nor U656 (N_656,In_850,In_1083);
nor U657 (N_657,In_879,In_398);
nor U658 (N_658,In_272,In_49);
and U659 (N_659,In_1355,In_164);
nand U660 (N_660,In_412,In_908);
nand U661 (N_661,In_1081,In_1025);
or U662 (N_662,In_819,In_229);
or U663 (N_663,In_163,In_929);
and U664 (N_664,In_991,In_1216);
nand U665 (N_665,In_1030,In_881);
nand U666 (N_666,In_916,In_36);
and U667 (N_667,In_745,In_696);
nor U668 (N_668,In_640,In_475);
and U669 (N_669,In_556,In_61);
and U670 (N_670,In_108,In_1031);
nor U671 (N_671,In_1353,In_344);
or U672 (N_672,In_824,In_148);
and U673 (N_673,In_400,In_690);
nor U674 (N_674,In_1357,In_1381);
and U675 (N_675,In_895,In_32);
and U676 (N_676,In_1124,In_615);
nor U677 (N_677,In_822,In_1218);
nand U678 (N_678,In_1205,In_829);
nor U679 (N_679,In_1012,In_1416);
nor U680 (N_680,In_898,In_399);
nor U681 (N_681,In_680,In_428);
nand U682 (N_682,In_1363,In_998);
nor U683 (N_683,In_1313,In_545);
or U684 (N_684,In_503,In_441);
nand U685 (N_685,In_1159,In_717);
nand U686 (N_686,In_842,In_586);
or U687 (N_687,In_697,In_1173);
and U688 (N_688,In_251,In_729);
and U689 (N_689,In_277,In_226);
or U690 (N_690,In_761,In_621);
or U691 (N_691,In_977,In_1445);
nor U692 (N_692,In_1387,In_541);
or U693 (N_693,In_1149,In_115);
nor U694 (N_694,In_592,In_863);
nor U695 (N_695,In_827,In_365);
nand U696 (N_696,In_574,In_321);
and U697 (N_697,In_116,In_981);
nor U698 (N_698,In_145,In_458);
or U699 (N_699,In_1003,In_350);
and U700 (N_700,In_638,In_65);
and U701 (N_701,In_1317,In_238);
and U702 (N_702,In_328,In_1337);
nor U703 (N_703,In_69,In_239);
nor U704 (N_704,In_752,In_1403);
nand U705 (N_705,In_252,In_548);
nand U706 (N_706,In_608,In_0);
nand U707 (N_707,In_97,In_1186);
or U708 (N_708,In_1334,In_744);
nor U709 (N_709,In_1474,In_1099);
and U710 (N_710,In_1160,In_132);
nand U711 (N_711,In_1283,In_137);
nor U712 (N_712,In_1215,In_175);
nor U713 (N_713,In_888,In_326);
nor U714 (N_714,In_1091,In_783);
nand U715 (N_715,In_57,In_394);
nand U716 (N_716,In_142,In_1203);
nand U717 (N_717,In_131,In_1495);
and U718 (N_718,In_1121,In_893);
nand U719 (N_719,In_4,In_443);
and U720 (N_720,In_577,In_159);
and U721 (N_721,In_28,In_1304);
nand U722 (N_722,In_477,In_1105);
and U723 (N_723,In_1284,In_607);
nand U724 (N_724,In_1035,In_972);
nand U725 (N_725,In_897,In_810);
and U726 (N_726,In_92,In_457);
nor U727 (N_727,In_1343,In_307);
or U728 (N_728,In_915,In_663);
or U729 (N_729,In_519,In_622);
and U730 (N_730,In_353,In_976);
nand U731 (N_731,In_1037,In_278);
nor U732 (N_732,In_611,In_528);
nor U733 (N_733,In_786,In_543);
nand U734 (N_734,In_712,In_416);
nand U735 (N_735,In_333,In_936);
or U736 (N_736,In_787,In_1458);
nor U737 (N_737,In_1443,In_983);
or U738 (N_738,In_276,In_1401);
or U739 (N_739,In_1271,In_504);
nand U740 (N_740,In_427,In_181);
nand U741 (N_741,In_1152,In_1429);
and U742 (N_742,In_1425,In_1092);
nand U743 (N_743,In_1135,In_486);
nand U744 (N_744,In_62,In_1054);
and U745 (N_745,In_704,In_918);
and U746 (N_746,In_1367,In_63);
and U747 (N_747,In_623,In_715);
nor U748 (N_748,In_1372,In_149);
nand U749 (N_749,In_1369,In_370);
nor U750 (N_750,In_678,In_181);
and U751 (N_751,In_608,In_396);
nor U752 (N_752,In_730,In_1384);
nor U753 (N_753,In_1220,In_348);
nand U754 (N_754,In_288,In_1470);
and U755 (N_755,In_1036,In_363);
nor U756 (N_756,In_232,In_459);
nand U757 (N_757,In_700,In_1355);
nor U758 (N_758,In_711,In_79);
nand U759 (N_759,In_1119,In_1497);
xor U760 (N_760,In_1227,In_1468);
nand U761 (N_761,In_1251,In_1214);
nor U762 (N_762,In_1315,In_730);
nand U763 (N_763,In_16,In_341);
and U764 (N_764,In_287,In_364);
and U765 (N_765,In_465,In_371);
nor U766 (N_766,In_1330,In_365);
and U767 (N_767,In_1110,In_1364);
or U768 (N_768,In_1197,In_250);
and U769 (N_769,In_825,In_1398);
or U770 (N_770,In_345,In_402);
nor U771 (N_771,In_1456,In_279);
and U772 (N_772,In_564,In_439);
or U773 (N_773,In_350,In_6);
nor U774 (N_774,In_254,In_268);
xnor U775 (N_775,In_407,In_1005);
xnor U776 (N_776,In_1439,In_1385);
nand U777 (N_777,In_401,In_630);
nor U778 (N_778,In_811,In_778);
and U779 (N_779,In_951,In_708);
or U780 (N_780,In_435,In_436);
nor U781 (N_781,In_1025,In_489);
and U782 (N_782,In_479,In_343);
nor U783 (N_783,In_800,In_257);
nand U784 (N_784,In_448,In_1193);
nand U785 (N_785,In_804,In_698);
or U786 (N_786,In_100,In_301);
and U787 (N_787,In_1324,In_1242);
or U788 (N_788,In_815,In_561);
or U789 (N_789,In_93,In_494);
or U790 (N_790,In_1191,In_1448);
or U791 (N_791,In_1001,In_757);
and U792 (N_792,In_1133,In_357);
nand U793 (N_793,In_1295,In_623);
or U794 (N_794,In_1222,In_890);
or U795 (N_795,In_774,In_239);
nand U796 (N_796,In_1102,In_490);
and U797 (N_797,In_693,In_347);
or U798 (N_798,In_1377,In_42);
nor U799 (N_799,In_1322,In_653);
nand U800 (N_800,In_38,In_732);
nand U801 (N_801,In_1109,In_203);
nand U802 (N_802,In_36,In_669);
nor U803 (N_803,In_1177,In_155);
or U804 (N_804,In_795,In_1369);
nand U805 (N_805,In_986,In_759);
or U806 (N_806,In_19,In_1423);
nor U807 (N_807,In_1195,In_1253);
or U808 (N_808,In_273,In_1402);
and U809 (N_809,In_1047,In_710);
or U810 (N_810,In_84,In_190);
nor U811 (N_811,In_440,In_41);
nor U812 (N_812,In_363,In_659);
nor U813 (N_813,In_1161,In_317);
or U814 (N_814,In_1253,In_1268);
nand U815 (N_815,In_1424,In_485);
and U816 (N_816,In_1239,In_1207);
and U817 (N_817,In_723,In_270);
and U818 (N_818,In_1053,In_1249);
nand U819 (N_819,In_1290,In_1407);
nor U820 (N_820,In_1016,In_672);
and U821 (N_821,In_76,In_596);
and U822 (N_822,In_533,In_139);
or U823 (N_823,In_620,In_1289);
nand U824 (N_824,In_781,In_480);
nor U825 (N_825,In_701,In_619);
or U826 (N_826,In_715,In_1466);
and U827 (N_827,In_998,In_748);
and U828 (N_828,In_696,In_713);
and U829 (N_829,In_50,In_805);
nand U830 (N_830,In_449,In_106);
nand U831 (N_831,In_837,In_64);
or U832 (N_832,In_1322,In_1016);
nor U833 (N_833,In_809,In_94);
or U834 (N_834,In_993,In_759);
nand U835 (N_835,In_267,In_236);
xor U836 (N_836,In_380,In_1051);
nor U837 (N_837,In_1239,In_136);
nor U838 (N_838,In_1484,In_752);
nand U839 (N_839,In_260,In_34);
nor U840 (N_840,In_1365,In_642);
nand U841 (N_841,In_652,In_308);
nand U842 (N_842,In_238,In_1443);
and U843 (N_843,In_619,In_147);
nand U844 (N_844,In_1438,In_216);
and U845 (N_845,In_391,In_705);
and U846 (N_846,In_403,In_684);
nand U847 (N_847,In_673,In_441);
and U848 (N_848,In_1293,In_1020);
nor U849 (N_849,In_533,In_1464);
nor U850 (N_850,In_935,In_1039);
and U851 (N_851,In_937,In_806);
or U852 (N_852,In_376,In_70);
nand U853 (N_853,In_123,In_21);
and U854 (N_854,In_263,In_595);
nand U855 (N_855,In_406,In_1134);
or U856 (N_856,In_1164,In_901);
nand U857 (N_857,In_258,In_1281);
nor U858 (N_858,In_38,In_1110);
and U859 (N_859,In_242,In_1024);
and U860 (N_860,In_656,In_930);
and U861 (N_861,In_89,In_872);
or U862 (N_862,In_999,In_1103);
nor U863 (N_863,In_1073,In_406);
or U864 (N_864,In_1375,In_1180);
nand U865 (N_865,In_964,In_882);
nor U866 (N_866,In_959,In_985);
nor U867 (N_867,In_10,In_1314);
nand U868 (N_868,In_929,In_325);
nand U869 (N_869,In_618,In_901);
or U870 (N_870,In_855,In_214);
nand U871 (N_871,In_828,In_1344);
or U872 (N_872,In_1169,In_1451);
nand U873 (N_873,In_1270,In_1100);
nand U874 (N_874,In_882,In_493);
and U875 (N_875,In_379,In_791);
nand U876 (N_876,In_723,In_1170);
nor U877 (N_877,In_190,In_1481);
nand U878 (N_878,In_1180,In_358);
nor U879 (N_879,In_5,In_921);
nand U880 (N_880,In_805,In_1207);
nand U881 (N_881,In_1436,In_494);
and U882 (N_882,In_417,In_1060);
and U883 (N_883,In_1219,In_687);
nand U884 (N_884,In_1310,In_1308);
nand U885 (N_885,In_760,In_1208);
nor U886 (N_886,In_233,In_741);
and U887 (N_887,In_514,In_1070);
or U888 (N_888,In_630,In_356);
or U889 (N_889,In_65,In_1469);
and U890 (N_890,In_686,In_1259);
xnor U891 (N_891,In_1226,In_381);
or U892 (N_892,In_249,In_145);
or U893 (N_893,In_994,In_1245);
and U894 (N_894,In_226,In_231);
or U895 (N_895,In_412,In_240);
nor U896 (N_896,In_1223,In_1225);
nand U897 (N_897,In_127,In_118);
nand U898 (N_898,In_1313,In_127);
or U899 (N_899,In_647,In_887);
or U900 (N_900,In_1076,In_378);
nand U901 (N_901,In_506,In_118);
and U902 (N_902,In_1120,In_1093);
and U903 (N_903,In_771,In_1081);
and U904 (N_904,In_331,In_1030);
and U905 (N_905,In_1083,In_1003);
nor U906 (N_906,In_834,In_20);
or U907 (N_907,In_800,In_223);
and U908 (N_908,In_858,In_1132);
nor U909 (N_909,In_299,In_556);
or U910 (N_910,In_456,In_829);
or U911 (N_911,In_951,In_845);
or U912 (N_912,In_252,In_906);
nand U913 (N_913,In_709,In_476);
or U914 (N_914,In_1400,In_391);
nor U915 (N_915,In_1328,In_91);
and U916 (N_916,In_780,In_539);
or U917 (N_917,In_491,In_324);
nor U918 (N_918,In_6,In_943);
or U919 (N_919,In_631,In_1148);
xor U920 (N_920,In_1194,In_397);
nor U921 (N_921,In_720,In_629);
and U922 (N_922,In_687,In_289);
nor U923 (N_923,In_113,In_1459);
nor U924 (N_924,In_688,In_1238);
or U925 (N_925,In_1047,In_461);
nor U926 (N_926,In_1312,In_621);
nor U927 (N_927,In_1086,In_84);
nor U928 (N_928,In_959,In_1078);
or U929 (N_929,In_1342,In_1327);
nand U930 (N_930,In_200,In_685);
or U931 (N_931,In_627,In_1475);
and U932 (N_932,In_965,In_1369);
nor U933 (N_933,In_1339,In_620);
or U934 (N_934,In_240,In_396);
nor U935 (N_935,In_910,In_1240);
or U936 (N_936,In_770,In_805);
and U937 (N_937,In_164,In_38);
and U938 (N_938,In_367,In_410);
nand U939 (N_939,In_793,In_129);
and U940 (N_940,In_1193,In_763);
or U941 (N_941,In_531,In_125);
or U942 (N_942,In_1320,In_1313);
and U943 (N_943,In_278,In_1029);
or U944 (N_944,In_613,In_673);
and U945 (N_945,In_478,In_195);
or U946 (N_946,In_275,In_16);
or U947 (N_947,In_137,In_142);
nor U948 (N_948,In_932,In_645);
and U949 (N_949,In_1150,In_985);
nor U950 (N_950,In_279,In_1330);
and U951 (N_951,In_1368,In_821);
nand U952 (N_952,In_812,In_1397);
nor U953 (N_953,In_1012,In_690);
nand U954 (N_954,In_75,In_954);
or U955 (N_955,In_717,In_1109);
nor U956 (N_956,In_1403,In_308);
or U957 (N_957,In_1140,In_367);
nor U958 (N_958,In_262,In_889);
nand U959 (N_959,In_829,In_277);
nor U960 (N_960,In_1404,In_383);
or U961 (N_961,In_501,In_1003);
nor U962 (N_962,In_229,In_154);
and U963 (N_963,In_241,In_1461);
or U964 (N_964,In_754,In_276);
or U965 (N_965,In_361,In_335);
nor U966 (N_966,In_1493,In_473);
nand U967 (N_967,In_300,In_662);
or U968 (N_968,In_640,In_693);
nor U969 (N_969,In_1186,In_566);
nand U970 (N_970,In_1095,In_1042);
and U971 (N_971,In_1325,In_215);
and U972 (N_972,In_81,In_862);
nand U973 (N_973,In_1298,In_1122);
and U974 (N_974,In_354,In_750);
nand U975 (N_975,In_975,In_1052);
and U976 (N_976,In_1241,In_348);
nor U977 (N_977,In_437,In_27);
xnor U978 (N_978,In_521,In_404);
or U979 (N_979,In_930,In_1358);
nor U980 (N_980,In_1499,In_977);
or U981 (N_981,In_20,In_305);
nor U982 (N_982,In_697,In_336);
nand U983 (N_983,In_172,In_1339);
or U984 (N_984,In_471,In_626);
and U985 (N_985,In_889,In_803);
or U986 (N_986,In_766,In_1273);
nand U987 (N_987,In_1140,In_804);
nor U988 (N_988,In_647,In_523);
or U989 (N_989,In_540,In_718);
nand U990 (N_990,In_474,In_410);
nor U991 (N_991,In_1411,In_1417);
and U992 (N_992,In_858,In_577);
nand U993 (N_993,In_600,In_449);
nand U994 (N_994,In_265,In_787);
nor U995 (N_995,In_1055,In_1334);
nand U996 (N_996,In_476,In_255);
nand U997 (N_997,In_1062,In_528);
nor U998 (N_998,In_576,In_223);
and U999 (N_999,In_1438,In_663);
and U1000 (N_1000,In_432,In_521);
nand U1001 (N_1001,In_1107,In_63);
or U1002 (N_1002,In_1479,In_279);
and U1003 (N_1003,In_971,In_1437);
or U1004 (N_1004,In_499,In_459);
or U1005 (N_1005,In_1419,In_260);
and U1006 (N_1006,In_459,In_660);
or U1007 (N_1007,In_337,In_477);
nand U1008 (N_1008,In_900,In_448);
or U1009 (N_1009,In_353,In_43);
or U1010 (N_1010,In_268,In_140);
or U1011 (N_1011,In_49,In_1140);
nor U1012 (N_1012,In_1316,In_1187);
nand U1013 (N_1013,In_1073,In_736);
or U1014 (N_1014,In_1229,In_263);
or U1015 (N_1015,In_1225,In_1120);
and U1016 (N_1016,In_870,In_605);
and U1017 (N_1017,In_1420,In_797);
or U1018 (N_1018,In_1342,In_1417);
nand U1019 (N_1019,In_854,In_176);
nand U1020 (N_1020,In_1119,In_71);
or U1021 (N_1021,In_1049,In_1020);
nor U1022 (N_1022,In_1318,In_500);
or U1023 (N_1023,In_741,In_1374);
xnor U1024 (N_1024,In_998,In_424);
and U1025 (N_1025,In_362,In_82);
and U1026 (N_1026,In_1114,In_963);
and U1027 (N_1027,In_1170,In_1237);
nor U1028 (N_1028,In_775,In_1356);
nor U1029 (N_1029,In_651,In_251);
or U1030 (N_1030,In_869,In_1439);
nand U1031 (N_1031,In_733,In_579);
or U1032 (N_1032,In_1499,In_21);
and U1033 (N_1033,In_1447,In_654);
or U1034 (N_1034,In_1068,In_380);
nand U1035 (N_1035,In_1480,In_441);
or U1036 (N_1036,In_1360,In_1022);
and U1037 (N_1037,In_304,In_887);
and U1038 (N_1038,In_1052,In_78);
or U1039 (N_1039,In_960,In_597);
nor U1040 (N_1040,In_230,In_75);
nor U1041 (N_1041,In_616,In_377);
nand U1042 (N_1042,In_1104,In_569);
and U1043 (N_1043,In_958,In_786);
and U1044 (N_1044,In_1327,In_471);
nand U1045 (N_1045,In_30,In_841);
or U1046 (N_1046,In_117,In_1407);
nor U1047 (N_1047,In_1467,In_453);
nand U1048 (N_1048,In_900,In_1113);
or U1049 (N_1049,In_959,In_1378);
or U1050 (N_1050,In_702,In_526);
and U1051 (N_1051,In_759,In_1351);
nor U1052 (N_1052,In_916,In_139);
nor U1053 (N_1053,In_1426,In_1126);
nand U1054 (N_1054,In_1031,In_441);
and U1055 (N_1055,In_783,In_1460);
nor U1056 (N_1056,In_264,In_1157);
or U1057 (N_1057,In_1304,In_234);
nand U1058 (N_1058,In_24,In_1161);
nor U1059 (N_1059,In_681,In_446);
nand U1060 (N_1060,In_616,In_447);
or U1061 (N_1061,In_411,In_740);
nand U1062 (N_1062,In_421,In_94);
nand U1063 (N_1063,In_547,In_1200);
nor U1064 (N_1064,In_589,In_953);
nor U1065 (N_1065,In_417,In_1435);
or U1066 (N_1066,In_1482,In_827);
nand U1067 (N_1067,In_141,In_1412);
nor U1068 (N_1068,In_1149,In_214);
and U1069 (N_1069,In_1002,In_349);
nand U1070 (N_1070,In_47,In_510);
or U1071 (N_1071,In_1213,In_242);
nand U1072 (N_1072,In_771,In_1276);
nand U1073 (N_1073,In_832,In_777);
nor U1074 (N_1074,In_1123,In_502);
xnor U1075 (N_1075,In_1123,In_443);
and U1076 (N_1076,In_48,In_1421);
nor U1077 (N_1077,In_1195,In_788);
or U1078 (N_1078,In_542,In_1349);
nor U1079 (N_1079,In_639,In_689);
nor U1080 (N_1080,In_688,In_255);
nor U1081 (N_1081,In_1011,In_764);
nor U1082 (N_1082,In_552,In_557);
or U1083 (N_1083,In_87,In_1432);
xor U1084 (N_1084,In_117,In_888);
nor U1085 (N_1085,In_1437,In_279);
nand U1086 (N_1086,In_710,In_838);
and U1087 (N_1087,In_1473,In_848);
nand U1088 (N_1088,In_172,In_910);
and U1089 (N_1089,In_336,In_988);
and U1090 (N_1090,In_422,In_23);
nand U1091 (N_1091,In_1061,In_1247);
nor U1092 (N_1092,In_1142,In_622);
nand U1093 (N_1093,In_1328,In_723);
nor U1094 (N_1094,In_1182,In_213);
nand U1095 (N_1095,In_869,In_111);
nand U1096 (N_1096,In_408,In_1065);
nand U1097 (N_1097,In_459,In_901);
and U1098 (N_1098,In_382,In_745);
nor U1099 (N_1099,In_856,In_810);
nand U1100 (N_1100,In_798,In_829);
nand U1101 (N_1101,In_189,In_118);
or U1102 (N_1102,In_55,In_195);
nand U1103 (N_1103,In_355,In_625);
and U1104 (N_1104,In_907,In_396);
and U1105 (N_1105,In_819,In_300);
nor U1106 (N_1106,In_78,In_782);
or U1107 (N_1107,In_966,In_971);
or U1108 (N_1108,In_184,In_481);
and U1109 (N_1109,In_992,In_735);
xor U1110 (N_1110,In_10,In_1296);
nor U1111 (N_1111,In_1258,In_451);
nand U1112 (N_1112,In_3,In_473);
and U1113 (N_1113,In_52,In_1001);
nand U1114 (N_1114,In_1067,In_1495);
nand U1115 (N_1115,In_1233,In_1446);
nand U1116 (N_1116,In_311,In_782);
or U1117 (N_1117,In_162,In_773);
nand U1118 (N_1118,In_1001,In_227);
or U1119 (N_1119,In_605,In_1105);
nand U1120 (N_1120,In_739,In_761);
nand U1121 (N_1121,In_974,In_1259);
or U1122 (N_1122,In_1067,In_132);
and U1123 (N_1123,In_906,In_884);
nor U1124 (N_1124,In_669,In_1165);
nor U1125 (N_1125,In_594,In_525);
and U1126 (N_1126,In_250,In_598);
and U1127 (N_1127,In_1150,In_967);
and U1128 (N_1128,In_1485,In_1444);
or U1129 (N_1129,In_219,In_1396);
nor U1130 (N_1130,In_610,In_733);
and U1131 (N_1131,In_1421,In_1427);
and U1132 (N_1132,In_300,In_793);
nand U1133 (N_1133,In_783,In_672);
or U1134 (N_1134,In_528,In_152);
nor U1135 (N_1135,In_1288,In_500);
and U1136 (N_1136,In_251,In_1065);
nand U1137 (N_1137,In_324,In_888);
nand U1138 (N_1138,In_1087,In_1430);
and U1139 (N_1139,In_1441,In_851);
or U1140 (N_1140,In_58,In_1038);
nor U1141 (N_1141,In_1475,In_1026);
or U1142 (N_1142,In_1328,In_879);
nor U1143 (N_1143,In_984,In_545);
and U1144 (N_1144,In_1416,In_1427);
nand U1145 (N_1145,In_337,In_379);
or U1146 (N_1146,In_193,In_1345);
nand U1147 (N_1147,In_475,In_1060);
or U1148 (N_1148,In_687,In_1233);
nand U1149 (N_1149,In_305,In_483);
xor U1150 (N_1150,In_881,In_1155);
nand U1151 (N_1151,In_495,In_1426);
nand U1152 (N_1152,In_1079,In_58);
nand U1153 (N_1153,In_749,In_583);
and U1154 (N_1154,In_394,In_314);
nand U1155 (N_1155,In_899,In_559);
nor U1156 (N_1156,In_321,In_752);
or U1157 (N_1157,In_221,In_133);
or U1158 (N_1158,In_594,In_1359);
or U1159 (N_1159,In_845,In_639);
nand U1160 (N_1160,In_442,In_409);
and U1161 (N_1161,In_1460,In_425);
or U1162 (N_1162,In_514,In_62);
or U1163 (N_1163,In_1311,In_276);
or U1164 (N_1164,In_1215,In_82);
and U1165 (N_1165,In_372,In_1308);
nand U1166 (N_1166,In_647,In_941);
nor U1167 (N_1167,In_875,In_514);
nand U1168 (N_1168,In_450,In_1136);
nand U1169 (N_1169,In_1061,In_1324);
and U1170 (N_1170,In_683,In_372);
or U1171 (N_1171,In_1339,In_94);
nor U1172 (N_1172,In_1434,In_268);
nor U1173 (N_1173,In_411,In_928);
nand U1174 (N_1174,In_68,In_190);
and U1175 (N_1175,In_239,In_547);
and U1176 (N_1176,In_541,In_58);
nor U1177 (N_1177,In_294,In_45);
or U1178 (N_1178,In_1303,In_548);
and U1179 (N_1179,In_103,In_1224);
xnor U1180 (N_1180,In_32,In_155);
nor U1181 (N_1181,In_994,In_25);
nor U1182 (N_1182,In_186,In_535);
and U1183 (N_1183,In_676,In_721);
and U1184 (N_1184,In_1085,In_1404);
or U1185 (N_1185,In_1061,In_1454);
or U1186 (N_1186,In_845,In_998);
and U1187 (N_1187,In_1067,In_1302);
nand U1188 (N_1188,In_635,In_605);
and U1189 (N_1189,In_1299,In_594);
and U1190 (N_1190,In_449,In_302);
and U1191 (N_1191,In_1138,In_1188);
or U1192 (N_1192,In_892,In_422);
or U1193 (N_1193,In_1178,In_736);
or U1194 (N_1194,In_1078,In_1184);
or U1195 (N_1195,In_308,In_62);
and U1196 (N_1196,In_45,In_20);
or U1197 (N_1197,In_15,In_1095);
or U1198 (N_1198,In_687,In_979);
or U1199 (N_1199,In_642,In_1453);
nor U1200 (N_1200,In_516,In_1285);
nand U1201 (N_1201,In_886,In_912);
nand U1202 (N_1202,In_773,In_1093);
nor U1203 (N_1203,In_569,In_1339);
and U1204 (N_1204,In_210,In_127);
nand U1205 (N_1205,In_472,In_1058);
nand U1206 (N_1206,In_809,In_1474);
nand U1207 (N_1207,In_369,In_1199);
nor U1208 (N_1208,In_1170,In_377);
nor U1209 (N_1209,In_425,In_382);
nor U1210 (N_1210,In_182,In_1381);
or U1211 (N_1211,In_1037,In_841);
nand U1212 (N_1212,In_19,In_653);
and U1213 (N_1213,In_1131,In_577);
xor U1214 (N_1214,In_637,In_241);
nand U1215 (N_1215,In_613,In_238);
and U1216 (N_1216,In_786,In_639);
and U1217 (N_1217,In_42,In_742);
and U1218 (N_1218,In_795,In_281);
and U1219 (N_1219,In_400,In_1280);
and U1220 (N_1220,In_807,In_1210);
or U1221 (N_1221,In_1346,In_435);
nor U1222 (N_1222,In_766,In_435);
nand U1223 (N_1223,In_42,In_134);
or U1224 (N_1224,In_533,In_1364);
nor U1225 (N_1225,In_370,In_164);
or U1226 (N_1226,In_340,In_1106);
or U1227 (N_1227,In_1117,In_1024);
nor U1228 (N_1228,In_366,In_1208);
or U1229 (N_1229,In_1247,In_647);
xnor U1230 (N_1230,In_1237,In_1494);
nand U1231 (N_1231,In_973,In_616);
or U1232 (N_1232,In_193,In_423);
nor U1233 (N_1233,In_1293,In_1277);
nor U1234 (N_1234,In_589,In_841);
or U1235 (N_1235,In_1385,In_530);
nor U1236 (N_1236,In_366,In_1063);
nor U1237 (N_1237,In_1292,In_1407);
nand U1238 (N_1238,In_854,In_441);
nor U1239 (N_1239,In_804,In_1392);
or U1240 (N_1240,In_1198,In_581);
and U1241 (N_1241,In_1485,In_114);
and U1242 (N_1242,In_584,In_959);
nand U1243 (N_1243,In_1148,In_158);
or U1244 (N_1244,In_65,In_260);
nand U1245 (N_1245,In_192,In_647);
or U1246 (N_1246,In_1169,In_1214);
or U1247 (N_1247,In_579,In_549);
or U1248 (N_1248,In_1152,In_39);
xor U1249 (N_1249,In_552,In_203);
nor U1250 (N_1250,In_288,In_1432);
or U1251 (N_1251,In_170,In_380);
and U1252 (N_1252,In_1234,In_1089);
and U1253 (N_1253,In_1004,In_46);
or U1254 (N_1254,In_1020,In_936);
nor U1255 (N_1255,In_1016,In_1020);
and U1256 (N_1256,In_762,In_1090);
nand U1257 (N_1257,In_1042,In_170);
and U1258 (N_1258,In_548,In_609);
nor U1259 (N_1259,In_926,In_181);
or U1260 (N_1260,In_974,In_1247);
and U1261 (N_1261,In_1040,In_1411);
nor U1262 (N_1262,In_368,In_942);
nand U1263 (N_1263,In_1063,In_330);
and U1264 (N_1264,In_1141,In_1328);
nand U1265 (N_1265,In_436,In_1470);
nor U1266 (N_1266,In_1160,In_505);
or U1267 (N_1267,In_166,In_1193);
nor U1268 (N_1268,In_1035,In_294);
or U1269 (N_1269,In_631,In_295);
and U1270 (N_1270,In_310,In_706);
or U1271 (N_1271,In_165,In_110);
nand U1272 (N_1272,In_613,In_1264);
or U1273 (N_1273,In_1422,In_1179);
or U1274 (N_1274,In_1282,In_144);
nand U1275 (N_1275,In_1216,In_1114);
nor U1276 (N_1276,In_132,In_261);
nand U1277 (N_1277,In_344,In_734);
nor U1278 (N_1278,In_777,In_1140);
nand U1279 (N_1279,In_1466,In_270);
nand U1280 (N_1280,In_179,In_710);
nor U1281 (N_1281,In_1298,In_820);
nor U1282 (N_1282,In_587,In_1403);
nand U1283 (N_1283,In_1324,In_307);
or U1284 (N_1284,In_1059,In_171);
nor U1285 (N_1285,In_1252,In_227);
nand U1286 (N_1286,In_1292,In_693);
xor U1287 (N_1287,In_174,In_683);
and U1288 (N_1288,In_431,In_1029);
nor U1289 (N_1289,In_777,In_702);
nand U1290 (N_1290,In_621,In_69);
nor U1291 (N_1291,In_415,In_1063);
nand U1292 (N_1292,In_125,In_45);
or U1293 (N_1293,In_925,In_1399);
nor U1294 (N_1294,In_1463,In_886);
nand U1295 (N_1295,In_753,In_426);
or U1296 (N_1296,In_436,In_749);
and U1297 (N_1297,In_145,In_1224);
nand U1298 (N_1298,In_1260,In_1154);
or U1299 (N_1299,In_870,In_241);
or U1300 (N_1300,In_976,In_259);
nor U1301 (N_1301,In_859,In_1272);
or U1302 (N_1302,In_1240,In_23);
nor U1303 (N_1303,In_1281,In_780);
and U1304 (N_1304,In_515,In_549);
and U1305 (N_1305,In_478,In_286);
nor U1306 (N_1306,In_83,In_1364);
or U1307 (N_1307,In_1086,In_987);
and U1308 (N_1308,In_751,In_1124);
nand U1309 (N_1309,In_207,In_703);
or U1310 (N_1310,In_1220,In_1410);
nor U1311 (N_1311,In_1181,In_1090);
nand U1312 (N_1312,In_1145,In_1134);
nand U1313 (N_1313,In_341,In_69);
nor U1314 (N_1314,In_1468,In_750);
nor U1315 (N_1315,In_869,In_819);
nand U1316 (N_1316,In_1492,In_1401);
or U1317 (N_1317,In_157,In_1416);
nand U1318 (N_1318,In_400,In_1445);
and U1319 (N_1319,In_960,In_1491);
nand U1320 (N_1320,In_125,In_1327);
nand U1321 (N_1321,In_976,In_1432);
and U1322 (N_1322,In_469,In_764);
nand U1323 (N_1323,In_3,In_795);
and U1324 (N_1324,In_954,In_873);
nor U1325 (N_1325,In_12,In_1159);
nand U1326 (N_1326,In_1079,In_989);
nor U1327 (N_1327,In_589,In_1201);
nor U1328 (N_1328,In_1083,In_404);
nand U1329 (N_1329,In_980,In_604);
nor U1330 (N_1330,In_1075,In_807);
nor U1331 (N_1331,In_909,In_65);
or U1332 (N_1332,In_237,In_844);
and U1333 (N_1333,In_389,In_495);
or U1334 (N_1334,In_812,In_713);
nor U1335 (N_1335,In_923,In_255);
nor U1336 (N_1336,In_840,In_503);
nor U1337 (N_1337,In_427,In_242);
nor U1338 (N_1338,In_1445,In_1204);
nand U1339 (N_1339,In_737,In_630);
nor U1340 (N_1340,In_1351,In_118);
and U1341 (N_1341,In_1468,In_513);
nand U1342 (N_1342,In_514,In_825);
and U1343 (N_1343,In_1074,In_110);
nor U1344 (N_1344,In_1134,In_1303);
nand U1345 (N_1345,In_772,In_1260);
nor U1346 (N_1346,In_1146,In_787);
xor U1347 (N_1347,In_1403,In_1267);
nor U1348 (N_1348,In_1394,In_497);
nand U1349 (N_1349,In_461,In_1477);
or U1350 (N_1350,In_662,In_85);
or U1351 (N_1351,In_1128,In_1132);
or U1352 (N_1352,In_42,In_1252);
and U1353 (N_1353,In_1110,In_1055);
and U1354 (N_1354,In_1390,In_24);
or U1355 (N_1355,In_784,In_1065);
nand U1356 (N_1356,In_723,In_1011);
nand U1357 (N_1357,In_996,In_1391);
nand U1358 (N_1358,In_891,In_994);
and U1359 (N_1359,In_271,In_982);
nor U1360 (N_1360,In_389,In_1224);
nand U1361 (N_1361,In_1405,In_927);
nand U1362 (N_1362,In_66,In_633);
or U1363 (N_1363,In_587,In_146);
or U1364 (N_1364,In_1413,In_953);
and U1365 (N_1365,In_3,In_1165);
and U1366 (N_1366,In_1365,In_974);
nor U1367 (N_1367,In_1354,In_880);
xor U1368 (N_1368,In_1120,In_60);
or U1369 (N_1369,In_555,In_946);
and U1370 (N_1370,In_578,In_259);
and U1371 (N_1371,In_1078,In_517);
nor U1372 (N_1372,In_1198,In_1454);
nor U1373 (N_1373,In_219,In_476);
nand U1374 (N_1374,In_1075,In_512);
nor U1375 (N_1375,In_1462,In_668);
nor U1376 (N_1376,In_741,In_607);
nand U1377 (N_1377,In_496,In_507);
nand U1378 (N_1378,In_340,In_850);
or U1379 (N_1379,In_590,In_1317);
nand U1380 (N_1380,In_474,In_428);
nor U1381 (N_1381,In_1443,In_164);
nand U1382 (N_1382,In_66,In_927);
or U1383 (N_1383,In_335,In_525);
nand U1384 (N_1384,In_784,In_1130);
nor U1385 (N_1385,In_629,In_60);
nand U1386 (N_1386,In_968,In_353);
nand U1387 (N_1387,In_1138,In_587);
or U1388 (N_1388,In_1322,In_1105);
nand U1389 (N_1389,In_629,In_218);
or U1390 (N_1390,In_1401,In_356);
nand U1391 (N_1391,In_519,In_1189);
and U1392 (N_1392,In_359,In_766);
or U1393 (N_1393,In_1432,In_1193);
nor U1394 (N_1394,In_1198,In_658);
nor U1395 (N_1395,In_1411,In_890);
or U1396 (N_1396,In_1128,In_1465);
or U1397 (N_1397,In_864,In_925);
nor U1398 (N_1398,In_341,In_526);
nor U1399 (N_1399,In_1160,In_1041);
or U1400 (N_1400,In_130,In_548);
or U1401 (N_1401,In_82,In_137);
and U1402 (N_1402,In_1187,In_831);
nand U1403 (N_1403,In_417,In_1225);
nor U1404 (N_1404,In_1235,In_1174);
xnor U1405 (N_1405,In_186,In_1343);
xnor U1406 (N_1406,In_90,In_1205);
nand U1407 (N_1407,In_726,In_635);
nand U1408 (N_1408,In_520,In_1478);
or U1409 (N_1409,In_526,In_552);
and U1410 (N_1410,In_504,In_441);
and U1411 (N_1411,In_393,In_1291);
nand U1412 (N_1412,In_772,In_970);
or U1413 (N_1413,In_830,In_761);
nor U1414 (N_1414,In_133,In_1166);
and U1415 (N_1415,In_124,In_425);
or U1416 (N_1416,In_212,In_730);
nor U1417 (N_1417,In_1065,In_65);
or U1418 (N_1418,In_426,In_225);
nand U1419 (N_1419,In_934,In_1159);
nor U1420 (N_1420,In_1167,In_460);
or U1421 (N_1421,In_472,In_1306);
and U1422 (N_1422,In_1001,In_1142);
nor U1423 (N_1423,In_1330,In_108);
nand U1424 (N_1424,In_177,In_839);
nand U1425 (N_1425,In_172,In_1214);
and U1426 (N_1426,In_131,In_744);
nand U1427 (N_1427,In_1028,In_1126);
nand U1428 (N_1428,In_992,In_885);
nor U1429 (N_1429,In_883,In_645);
or U1430 (N_1430,In_782,In_490);
nor U1431 (N_1431,In_1263,In_824);
and U1432 (N_1432,In_266,In_34);
or U1433 (N_1433,In_834,In_782);
nor U1434 (N_1434,In_351,In_593);
xor U1435 (N_1435,In_1389,In_793);
or U1436 (N_1436,In_866,In_1136);
nor U1437 (N_1437,In_677,In_1233);
nor U1438 (N_1438,In_947,In_1208);
nand U1439 (N_1439,In_1252,In_279);
or U1440 (N_1440,In_175,In_1117);
and U1441 (N_1441,In_176,In_1363);
or U1442 (N_1442,In_540,In_1147);
nor U1443 (N_1443,In_579,In_1066);
xnor U1444 (N_1444,In_1493,In_973);
nor U1445 (N_1445,In_390,In_1107);
nor U1446 (N_1446,In_806,In_795);
nor U1447 (N_1447,In_1492,In_427);
or U1448 (N_1448,In_156,In_228);
and U1449 (N_1449,In_1084,In_169);
nor U1450 (N_1450,In_642,In_996);
nor U1451 (N_1451,In_343,In_285);
or U1452 (N_1452,In_367,In_158);
nor U1453 (N_1453,In_708,In_1378);
and U1454 (N_1454,In_358,In_829);
nand U1455 (N_1455,In_323,In_95);
or U1456 (N_1456,In_557,In_1444);
nor U1457 (N_1457,In_221,In_24);
and U1458 (N_1458,In_1380,In_1372);
nor U1459 (N_1459,In_951,In_1267);
or U1460 (N_1460,In_1089,In_744);
nor U1461 (N_1461,In_489,In_174);
nand U1462 (N_1462,In_1007,In_1335);
and U1463 (N_1463,In_1443,In_513);
or U1464 (N_1464,In_604,In_395);
nand U1465 (N_1465,In_1218,In_60);
and U1466 (N_1466,In_1424,In_543);
or U1467 (N_1467,In_1401,In_980);
and U1468 (N_1468,In_56,In_1026);
nand U1469 (N_1469,In_657,In_511);
or U1470 (N_1470,In_329,In_449);
or U1471 (N_1471,In_1209,In_355);
nand U1472 (N_1472,In_1084,In_264);
and U1473 (N_1473,In_141,In_315);
nor U1474 (N_1474,In_1045,In_335);
xnor U1475 (N_1475,In_1240,In_1440);
nand U1476 (N_1476,In_1319,In_1029);
or U1477 (N_1477,In_21,In_1048);
nor U1478 (N_1478,In_1313,In_631);
or U1479 (N_1479,In_56,In_908);
or U1480 (N_1480,In_1494,In_144);
or U1481 (N_1481,In_114,In_427);
or U1482 (N_1482,In_1103,In_1469);
nor U1483 (N_1483,In_1023,In_1205);
or U1484 (N_1484,In_1430,In_657);
nand U1485 (N_1485,In_1016,In_1242);
nor U1486 (N_1486,In_1486,In_1214);
or U1487 (N_1487,In_193,In_1492);
and U1488 (N_1488,In_1466,In_1143);
or U1489 (N_1489,In_1096,In_788);
xnor U1490 (N_1490,In_1034,In_350);
xnor U1491 (N_1491,In_683,In_1108);
or U1492 (N_1492,In_1240,In_1041);
or U1493 (N_1493,In_999,In_1378);
nand U1494 (N_1494,In_1019,In_956);
and U1495 (N_1495,In_1176,In_1348);
and U1496 (N_1496,In_1429,In_1446);
or U1497 (N_1497,In_862,In_1413);
nor U1498 (N_1498,In_51,In_977);
and U1499 (N_1499,In_361,In_738);
and U1500 (N_1500,In_704,In_468);
or U1501 (N_1501,In_1061,In_238);
and U1502 (N_1502,In_348,In_742);
or U1503 (N_1503,In_40,In_453);
or U1504 (N_1504,In_148,In_546);
xnor U1505 (N_1505,In_542,In_1240);
or U1506 (N_1506,In_1236,In_43);
and U1507 (N_1507,In_824,In_649);
or U1508 (N_1508,In_807,In_996);
nand U1509 (N_1509,In_1192,In_675);
or U1510 (N_1510,In_531,In_707);
nor U1511 (N_1511,In_229,In_1403);
and U1512 (N_1512,In_1111,In_562);
nor U1513 (N_1513,In_252,In_1);
nand U1514 (N_1514,In_534,In_685);
nand U1515 (N_1515,In_985,In_800);
nand U1516 (N_1516,In_1127,In_119);
nand U1517 (N_1517,In_165,In_251);
or U1518 (N_1518,In_798,In_719);
nand U1519 (N_1519,In_499,In_813);
nor U1520 (N_1520,In_1367,In_837);
nand U1521 (N_1521,In_474,In_515);
or U1522 (N_1522,In_709,In_1279);
and U1523 (N_1523,In_1122,In_601);
nand U1524 (N_1524,In_1381,In_1147);
or U1525 (N_1525,In_628,In_1380);
nand U1526 (N_1526,In_802,In_868);
nand U1527 (N_1527,In_632,In_689);
nor U1528 (N_1528,In_1122,In_439);
nor U1529 (N_1529,In_900,In_771);
or U1530 (N_1530,In_1167,In_714);
nand U1531 (N_1531,In_697,In_1284);
and U1532 (N_1532,In_640,In_1013);
and U1533 (N_1533,In_394,In_1477);
nand U1534 (N_1534,In_1325,In_1264);
and U1535 (N_1535,In_24,In_1382);
or U1536 (N_1536,In_638,In_1445);
xor U1537 (N_1537,In_1458,In_542);
or U1538 (N_1538,In_341,In_1271);
or U1539 (N_1539,In_631,In_61);
nand U1540 (N_1540,In_142,In_67);
nor U1541 (N_1541,In_727,In_1086);
or U1542 (N_1542,In_1348,In_51);
nor U1543 (N_1543,In_1358,In_224);
nor U1544 (N_1544,In_1368,In_1317);
nand U1545 (N_1545,In_171,In_1225);
nand U1546 (N_1546,In_1369,In_658);
nor U1547 (N_1547,In_520,In_180);
nor U1548 (N_1548,In_480,In_297);
nand U1549 (N_1549,In_5,In_401);
nand U1550 (N_1550,In_197,In_960);
and U1551 (N_1551,In_861,In_89);
nor U1552 (N_1552,In_1126,In_965);
and U1553 (N_1553,In_123,In_1228);
nor U1554 (N_1554,In_79,In_1425);
and U1555 (N_1555,In_227,In_321);
nor U1556 (N_1556,In_329,In_38);
or U1557 (N_1557,In_563,In_41);
nor U1558 (N_1558,In_917,In_886);
or U1559 (N_1559,In_102,In_439);
nand U1560 (N_1560,In_187,In_1485);
or U1561 (N_1561,In_68,In_121);
and U1562 (N_1562,In_1335,In_172);
nor U1563 (N_1563,In_331,In_774);
or U1564 (N_1564,In_1468,In_396);
nor U1565 (N_1565,In_796,In_786);
nor U1566 (N_1566,In_1113,In_901);
nor U1567 (N_1567,In_238,In_471);
and U1568 (N_1568,In_225,In_496);
nor U1569 (N_1569,In_796,In_319);
or U1570 (N_1570,In_698,In_1148);
or U1571 (N_1571,In_1470,In_1264);
and U1572 (N_1572,In_265,In_1108);
nand U1573 (N_1573,In_667,In_1337);
nor U1574 (N_1574,In_580,In_1313);
nor U1575 (N_1575,In_1363,In_1043);
and U1576 (N_1576,In_1006,In_968);
or U1577 (N_1577,In_846,In_780);
or U1578 (N_1578,In_1101,In_581);
nor U1579 (N_1579,In_219,In_21);
and U1580 (N_1580,In_1321,In_1487);
or U1581 (N_1581,In_43,In_887);
nand U1582 (N_1582,In_706,In_467);
or U1583 (N_1583,In_1020,In_116);
nand U1584 (N_1584,In_168,In_59);
nand U1585 (N_1585,In_698,In_75);
or U1586 (N_1586,In_300,In_77);
nor U1587 (N_1587,In_655,In_480);
nand U1588 (N_1588,In_300,In_653);
and U1589 (N_1589,In_135,In_996);
or U1590 (N_1590,In_327,In_1104);
nand U1591 (N_1591,In_823,In_261);
and U1592 (N_1592,In_717,In_1186);
or U1593 (N_1593,In_133,In_1007);
and U1594 (N_1594,In_729,In_1480);
and U1595 (N_1595,In_181,In_492);
xnor U1596 (N_1596,In_311,In_420);
and U1597 (N_1597,In_203,In_441);
nor U1598 (N_1598,In_494,In_990);
nor U1599 (N_1599,In_1370,In_1384);
or U1600 (N_1600,In_615,In_493);
nand U1601 (N_1601,In_877,In_375);
nand U1602 (N_1602,In_527,In_1484);
nor U1603 (N_1603,In_1412,In_134);
or U1604 (N_1604,In_761,In_95);
or U1605 (N_1605,In_1432,In_869);
nor U1606 (N_1606,In_1299,In_1133);
nand U1607 (N_1607,In_823,In_1213);
nand U1608 (N_1608,In_877,In_1355);
nor U1609 (N_1609,In_425,In_533);
nor U1610 (N_1610,In_199,In_1080);
nand U1611 (N_1611,In_295,In_810);
or U1612 (N_1612,In_666,In_891);
nor U1613 (N_1613,In_1305,In_271);
or U1614 (N_1614,In_239,In_127);
nor U1615 (N_1615,In_595,In_972);
nand U1616 (N_1616,In_1385,In_486);
and U1617 (N_1617,In_230,In_1449);
nor U1618 (N_1618,In_848,In_28);
nand U1619 (N_1619,In_102,In_680);
nor U1620 (N_1620,In_422,In_180);
xnor U1621 (N_1621,In_1100,In_1420);
nand U1622 (N_1622,In_1426,In_540);
and U1623 (N_1623,In_690,In_316);
and U1624 (N_1624,In_81,In_250);
and U1625 (N_1625,In_1230,In_624);
or U1626 (N_1626,In_801,In_739);
nand U1627 (N_1627,In_631,In_91);
nor U1628 (N_1628,In_1214,In_1355);
and U1629 (N_1629,In_407,In_1304);
nand U1630 (N_1630,In_1478,In_903);
and U1631 (N_1631,In_30,In_1482);
and U1632 (N_1632,In_60,In_1051);
or U1633 (N_1633,In_205,In_138);
or U1634 (N_1634,In_290,In_468);
or U1635 (N_1635,In_685,In_175);
nor U1636 (N_1636,In_1006,In_209);
and U1637 (N_1637,In_1125,In_1102);
and U1638 (N_1638,In_709,In_1490);
or U1639 (N_1639,In_1307,In_840);
nand U1640 (N_1640,In_423,In_1439);
and U1641 (N_1641,In_598,In_1326);
or U1642 (N_1642,In_287,In_89);
and U1643 (N_1643,In_1174,In_684);
or U1644 (N_1644,In_63,In_1209);
and U1645 (N_1645,In_876,In_1093);
and U1646 (N_1646,In_1147,In_32);
nor U1647 (N_1647,In_730,In_32);
nor U1648 (N_1648,In_886,In_376);
nand U1649 (N_1649,In_957,In_236);
or U1650 (N_1650,In_1203,In_1284);
nand U1651 (N_1651,In_400,In_410);
nor U1652 (N_1652,In_44,In_678);
nand U1653 (N_1653,In_628,In_1171);
nor U1654 (N_1654,In_753,In_1);
nand U1655 (N_1655,In_268,In_106);
nor U1656 (N_1656,In_365,In_174);
or U1657 (N_1657,In_525,In_156);
or U1658 (N_1658,In_381,In_536);
or U1659 (N_1659,In_971,In_1075);
or U1660 (N_1660,In_95,In_1089);
nor U1661 (N_1661,In_568,In_503);
or U1662 (N_1662,In_1333,In_577);
nor U1663 (N_1663,In_123,In_93);
nor U1664 (N_1664,In_1311,In_762);
nand U1665 (N_1665,In_582,In_1391);
or U1666 (N_1666,In_994,In_314);
nand U1667 (N_1667,In_1406,In_220);
and U1668 (N_1668,In_1455,In_36);
nor U1669 (N_1669,In_913,In_68);
nor U1670 (N_1670,In_765,In_1315);
or U1671 (N_1671,In_677,In_1119);
and U1672 (N_1672,In_90,In_126);
and U1673 (N_1673,In_85,In_3);
nand U1674 (N_1674,In_1482,In_787);
nor U1675 (N_1675,In_1298,In_323);
nand U1676 (N_1676,In_501,In_802);
nor U1677 (N_1677,In_815,In_1034);
or U1678 (N_1678,In_745,In_62);
nor U1679 (N_1679,In_1205,In_218);
and U1680 (N_1680,In_695,In_686);
or U1681 (N_1681,In_127,In_922);
and U1682 (N_1682,In_650,In_1317);
and U1683 (N_1683,In_1148,In_18);
nand U1684 (N_1684,In_399,In_268);
nand U1685 (N_1685,In_1352,In_878);
nor U1686 (N_1686,In_957,In_421);
or U1687 (N_1687,In_184,In_186);
or U1688 (N_1688,In_956,In_591);
nor U1689 (N_1689,In_1366,In_1035);
nor U1690 (N_1690,In_1422,In_337);
nand U1691 (N_1691,In_50,In_712);
nand U1692 (N_1692,In_638,In_803);
and U1693 (N_1693,In_905,In_470);
nor U1694 (N_1694,In_1031,In_1209);
nor U1695 (N_1695,In_1161,In_1301);
and U1696 (N_1696,In_747,In_888);
and U1697 (N_1697,In_323,In_797);
nor U1698 (N_1698,In_1389,In_140);
nor U1699 (N_1699,In_931,In_984);
or U1700 (N_1700,In_1406,In_366);
and U1701 (N_1701,In_895,In_1318);
nand U1702 (N_1702,In_1378,In_1027);
and U1703 (N_1703,In_653,In_737);
and U1704 (N_1704,In_255,In_676);
and U1705 (N_1705,In_1149,In_1166);
or U1706 (N_1706,In_908,In_1020);
and U1707 (N_1707,In_652,In_363);
nand U1708 (N_1708,In_1131,In_1007);
nand U1709 (N_1709,In_1413,In_1224);
and U1710 (N_1710,In_682,In_247);
nand U1711 (N_1711,In_310,In_704);
nand U1712 (N_1712,In_293,In_1158);
nor U1713 (N_1713,In_542,In_580);
nand U1714 (N_1714,In_57,In_1018);
or U1715 (N_1715,In_466,In_1450);
nand U1716 (N_1716,In_1318,In_1146);
nand U1717 (N_1717,In_1432,In_898);
and U1718 (N_1718,In_725,In_1068);
nor U1719 (N_1719,In_1214,In_522);
nand U1720 (N_1720,In_19,In_676);
or U1721 (N_1721,In_257,In_413);
and U1722 (N_1722,In_176,In_1277);
or U1723 (N_1723,In_1497,In_1340);
nor U1724 (N_1724,In_347,In_225);
or U1725 (N_1725,In_1324,In_508);
nand U1726 (N_1726,In_831,In_1370);
or U1727 (N_1727,In_1103,In_1280);
nor U1728 (N_1728,In_1108,In_648);
or U1729 (N_1729,In_1426,In_829);
nand U1730 (N_1730,In_1495,In_977);
or U1731 (N_1731,In_660,In_1007);
or U1732 (N_1732,In_1340,In_1138);
and U1733 (N_1733,In_339,In_865);
nor U1734 (N_1734,In_320,In_598);
nor U1735 (N_1735,In_981,In_509);
or U1736 (N_1736,In_47,In_766);
and U1737 (N_1737,In_893,In_364);
or U1738 (N_1738,In_1088,In_910);
and U1739 (N_1739,In_441,In_1414);
or U1740 (N_1740,In_1490,In_1029);
nor U1741 (N_1741,In_565,In_1404);
nand U1742 (N_1742,In_1348,In_490);
nor U1743 (N_1743,In_719,In_82);
and U1744 (N_1744,In_1219,In_870);
nor U1745 (N_1745,In_431,In_239);
and U1746 (N_1746,In_1347,In_1154);
and U1747 (N_1747,In_860,In_475);
nor U1748 (N_1748,In_306,In_1137);
or U1749 (N_1749,In_326,In_845);
nand U1750 (N_1750,In_829,In_709);
nor U1751 (N_1751,In_163,In_478);
nand U1752 (N_1752,In_299,In_1270);
and U1753 (N_1753,In_1028,In_399);
or U1754 (N_1754,In_1486,In_1100);
and U1755 (N_1755,In_1248,In_1186);
nor U1756 (N_1756,In_37,In_1135);
or U1757 (N_1757,In_1363,In_575);
nor U1758 (N_1758,In_1468,In_294);
nand U1759 (N_1759,In_259,In_1396);
or U1760 (N_1760,In_211,In_274);
and U1761 (N_1761,In_180,In_752);
and U1762 (N_1762,In_583,In_1136);
or U1763 (N_1763,In_1305,In_880);
or U1764 (N_1764,In_1159,In_1172);
and U1765 (N_1765,In_33,In_515);
nor U1766 (N_1766,In_1175,In_610);
or U1767 (N_1767,In_217,In_1340);
and U1768 (N_1768,In_421,In_1088);
or U1769 (N_1769,In_824,In_557);
nor U1770 (N_1770,In_905,In_330);
or U1771 (N_1771,In_587,In_1280);
or U1772 (N_1772,In_810,In_334);
and U1773 (N_1773,In_1478,In_36);
nor U1774 (N_1774,In_1279,In_255);
nand U1775 (N_1775,In_347,In_45);
and U1776 (N_1776,In_919,In_992);
and U1777 (N_1777,In_1315,In_114);
nor U1778 (N_1778,In_967,In_641);
nand U1779 (N_1779,In_432,In_1277);
or U1780 (N_1780,In_638,In_493);
and U1781 (N_1781,In_475,In_284);
or U1782 (N_1782,In_606,In_207);
nor U1783 (N_1783,In_403,In_74);
or U1784 (N_1784,In_1419,In_756);
or U1785 (N_1785,In_887,In_162);
and U1786 (N_1786,In_1056,In_1265);
nand U1787 (N_1787,In_1123,In_329);
and U1788 (N_1788,In_864,In_1335);
nand U1789 (N_1789,In_1292,In_100);
and U1790 (N_1790,In_1060,In_406);
and U1791 (N_1791,In_450,In_929);
nand U1792 (N_1792,In_321,In_185);
or U1793 (N_1793,In_854,In_1495);
nor U1794 (N_1794,In_240,In_1431);
and U1795 (N_1795,In_1140,In_805);
and U1796 (N_1796,In_1244,In_195);
nand U1797 (N_1797,In_1083,In_227);
nand U1798 (N_1798,In_428,In_1440);
and U1799 (N_1799,In_830,In_493);
nand U1800 (N_1800,In_358,In_1016);
and U1801 (N_1801,In_888,In_1297);
or U1802 (N_1802,In_336,In_344);
and U1803 (N_1803,In_561,In_737);
and U1804 (N_1804,In_736,In_609);
nand U1805 (N_1805,In_776,In_957);
and U1806 (N_1806,In_992,In_331);
nor U1807 (N_1807,In_151,In_938);
and U1808 (N_1808,In_99,In_820);
and U1809 (N_1809,In_1007,In_156);
or U1810 (N_1810,In_1161,In_295);
nor U1811 (N_1811,In_1131,In_1423);
or U1812 (N_1812,In_360,In_825);
nor U1813 (N_1813,In_1368,In_587);
nand U1814 (N_1814,In_648,In_1078);
or U1815 (N_1815,In_723,In_239);
or U1816 (N_1816,In_1240,In_319);
nor U1817 (N_1817,In_423,In_1013);
nor U1818 (N_1818,In_1419,In_785);
nor U1819 (N_1819,In_94,In_131);
or U1820 (N_1820,In_621,In_1190);
or U1821 (N_1821,In_735,In_145);
nor U1822 (N_1822,In_891,In_560);
nor U1823 (N_1823,In_310,In_96);
nand U1824 (N_1824,In_1309,In_861);
or U1825 (N_1825,In_1295,In_202);
xnor U1826 (N_1826,In_231,In_437);
nor U1827 (N_1827,In_1319,In_486);
and U1828 (N_1828,In_106,In_189);
or U1829 (N_1829,In_1473,In_1192);
nand U1830 (N_1830,In_679,In_1457);
or U1831 (N_1831,In_586,In_902);
or U1832 (N_1832,In_932,In_508);
and U1833 (N_1833,In_1405,In_1249);
or U1834 (N_1834,In_674,In_149);
nor U1835 (N_1835,In_926,In_1014);
and U1836 (N_1836,In_949,In_381);
nor U1837 (N_1837,In_1459,In_147);
or U1838 (N_1838,In_794,In_115);
and U1839 (N_1839,In_1324,In_157);
nor U1840 (N_1840,In_1059,In_266);
or U1841 (N_1841,In_218,In_1191);
or U1842 (N_1842,In_683,In_379);
nor U1843 (N_1843,In_1019,In_653);
or U1844 (N_1844,In_632,In_621);
or U1845 (N_1845,In_247,In_1310);
or U1846 (N_1846,In_692,In_613);
nand U1847 (N_1847,In_215,In_1094);
nand U1848 (N_1848,In_91,In_1178);
and U1849 (N_1849,In_679,In_433);
nand U1850 (N_1850,In_130,In_1325);
or U1851 (N_1851,In_238,In_197);
and U1852 (N_1852,In_433,In_1335);
or U1853 (N_1853,In_251,In_205);
nor U1854 (N_1854,In_1019,In_346);
and U1855 (N_1855,In_645,In_293);
nand U1856 (N_1856,In_703,In_1022);
and U1857 (N_1857,In_806,In_264);
or U1858 (N_1858,In_1096,In_1328);
nor U1859 (N_1859,In_373,In_1190);
and U1860 (N_1860,In_1417,In_1083);
and U1861 (N_1861,In_1437,In_940);
and U1862 (N_1862,In_242,In_1381);
or U1863 (N_1863,In_732,In_1141);
nand U1864 (N_1864,In_123,In_1412);
nor U1865 (N_1865,In_1489,In_1102);
and U1866 (N_1866,In_1151,In_168);
and U1867 (N_1867,In_656,In_1269);
nor U1868 (N_1868,In_564,In_217);
or U1869 (N_1869,In_133,In_703);
nand U1870 (N_1870,In_971,In_846);
or U1871 (N_1871,In_461,In_631);
and U1872 (N_1872,In_1170,In_263);
nor U1873 (N_1873,In_1434,In_174);
or U1874 (N_1874,In_777,In_892);
or U1875 (N_1875,In_992,In_1384);
or U1876 (N_1876,In_365,In_79);
nor U1877 (N_1877,In_737,In_674);
nor U1878 (N_1878,In_384,In_323);
nand U1879 (N_1879,In_725,In_218);
nor U1880 (N_1880,In_340,In_22);
xor U1881 (N_1881,In_647,In_303);
nor U1882 (N_1882,In_2,In_1052);
nand U1883 (N_1883,In_91,In_319);
or U1884 (N_1884,In_134,In_838);
nor U1885 (N_1885,In_45,In_761);
or U1886 (N_1886,In_879,In_917);
and U1887 (N_1887,In_298,In_159);
and U1888 (N_1888,In_976,In_463);
or U1889 (N_1889,In_680,In_920);
or U1890 (N_1890,In_844,In_978);
or U1891 (N_1891,In_541,In_1235);
nand U1892 (N_1892,In_472,In_1424);
nor U1893 (N_1893,In_595,In_233);
nor U1894 (N_1894,In_258,In_918);
nor U1895 (N_1895,In_585,In_538);
xnor U1896 (N_1896,In_1444,In_189);
nand U1897 (N_1897,In_1098,In_615);
nor U1898 (N_1898,In_1140,In_890);
xor U1899 (N_1899,In_1380,In_1141);
nand U1900 (N_1900,In_770,In_60);
or U1901 (N_1901,In_1354,In_1133);
nand U1902 (N_1902,In_740,In_621);
or U1903 (N_1903,In_788,In_735);
nand U1904 (N_1904,In_1338,In_1393);
and U1905 (N_1905,In_1398,In_660);
nor U1906 (N_1906,In_1107,In_252);
and U1907 (N_1907,In_798,In_872);
and U1908 (N_1908,In_658,In_491);
and U1909 (N_1909,In_1347,In_1493);
nor U1910 (N_1910,In_1058,In_1409);
and U1911 (N_1911,In_1083,In_1468);
and U1912 (N_1912,In_1422,In_1065);
or U1913 (N_1913,In_1147,In_511);
nor U1914 (N_1914,In_1354,In_64);
nor U1915 (N_1915,In_1340,In_1376);
and U1916 (N_1916,In_339,In_367);
and U1917 (N_1917,In_1064,In_1489);
and U1918 (N_1918,In_1215,In_1234);
nand U1919 (N_1919,In_415,In_1198);
and U1920 (N_1920,In_1301,In_986);
and U1921 (N_1921,In_466,In_1054);
nand U1922 (N_1922,In_173,In_567);
or U1923 (N_1923,In_67,In_488);
nand U1924 (N_1924,In_1348,In_112);
nor U1925 (N_1925,In_1359,In_212);
nand U1926 (N_1926,In_51,In_13);
or U1927 (N_1927,In_1316,In_945);
and U1928 (N_1928,In_236,In_1494);
nand U1929 (N_1929,In_875,In_852);
nand U1930 (N_1930,In_828,In_71);
nand U1931 (N_1931,In_1123,In_334);
or U1932 (N_1932,In_1399,In_1019);
nor U1933 (N_1933,In_188,In_889);
and U1934 (N_1934,In_190,In_431);
nand U1935 (N_1935,In_1067,In_1428);
and U1936 (N_1936,In_410,In_251);
or U1937 (N_1937,In_85,In_607);
nor U1938 (N_1938,In_1027,In_644);
or U1939 (N_1939,In_1018,In_1142);
and U1940 (N_1940,In_816,In_759);
nand U1941 (N_1941,In_865,In_1014);
nand U1942 (N_1942,In_726,In_1476);
nor U1943 (N_1943,In_479,In_584);
nand U1944 (N_1944,In_805,In_691);
and U1945 (N_1945,In_878,In_198);
or U1946 (N_1946,In_1416,In_590);
nor U1947 (N_1947,In_891,In_1135);
nand U1948 (N_1948,In_541,In_422);
nand U1949 (N_1949,In_1183,In_632);
and U1950 (N_1950,In_501,In_651);
nand U1951 (N_1951,In_229,In_82);
and U1952 (N_1952,In_500,In_445);
or U1953 (N_1953,In_886,In_623);
nor U1954 (N_1954,In_1434,In_454);
and U1955 (N_1955,In_1492,In_548);
nor U1956 (N_1956,In_53,In_541);
nand U1957 (N_1957,In_1268,In_1321);
and U1958 (N_1958,In_898,In_71);
or U1959 (N_1959,In_646,In_955);
and U1960 (N_1960,In_725,In_532);
or U1961 (N_1961,In_302,In_964);
nor U1962 (N_1962,In_50,In_1444);
and U1963 (N_1963,In_96,In_837);
nor U1964 (N_1964,In_681,In_377);
nor U1965 (N_1965,In_1089,In_466);
or U1966 (N_1966,In_1021,In_543);
and U1967 (N_1967,In_233,In_1223);
nand U1968 (N_1968,In_82,In_1172);
or U1969 (N_1969,In_396,In_312);
or U1970 (N_1970,In_1324,In_151);
or U1971 (N_1971,In_112,In_1235);
and U1972 (N_1972,In_1079,In_304);
and U1973 (N_1973,In_1382,In_1081);
nor U1974 (N_1974,In_1086,In_1434);
nand U1975 (N_1975,In_654,In_733);
and U1976 (N_1976,In_224,In_1294);
or U1977 (N_1977,In_828,In_538);
and U1978 (N_1978,In_985,In_1310);
nor U1979 (N_1979,In_612,In_90);
nand U1980 (N_1980,In_1231,In_600);
nand U1981 (N_1981,In_874,In_779);
nand U1982 (N_1982,In_881,In_579);
nor U1983 (N_1983,In_1226,In_783);
nor U1984 (N_1984,In_1481,In_788);
nand U1985 (N_1985,In_282,In_178);
or U1986 (N_1986,In_474,In_414);
or U1987 (N_1987,In_735,In_796);
nand U1988 (N_1988,In_291,In_494);
and U1989 (N_1989,In_284,In_397);
and U1990 (N_1990,In_1408,In_207);
and U1991 (N_1991,In_167,In_251);
nor U1992 (N_1992,In_522,In_1086);
nand U1993 (N_1993,In_1272,In_652);
nand U1994 (N_1994,In_1387,In_775);
nor U1995 (N_1995,In_1187,In_487);
and U1996 (N_1996,In_455,In_636);
nor U1997 (N_1997,In_1298,In_1192);
nand U1998 (N_1998,In_1134,In_1022);
nand U1999 (N_1999,In_784,In_1410);
or U2000 (N_2000,In_130,In_606);
nor U2001 (N_2001,In_33,In_1455);
nand U2002 (N_2002,In_1361,In_1186);
and U2003 (N_2003,In_1427,In_1455);
nand U2004 (N_2004,In_178,In_1282);
nor U2005 (N_2005,In_1170,In_1383);
and U2006 (N_2006,In_878,In_158);
nor U2007 (N_2007,In_794,In_684);
or U2008 (N_2008,In_110,In_441);
nor U2009 (N_2009,In_776,In_601);
nand U2010 (N_2010,In_1457,In_1327);
or U2011 (N_2011,In_1257,In_1270);
and U2012 (N_2012,In_1070,In_906);
and U2013 (N_2013,In_908,In_331);
or U2014 (N_2014,In_272,In_588);
nor U2015 (N_2015,In_208,In_716);
nand U2016 (N_2016,In_140,In_1254);
nor U2017 (N_2017,In_1413,In_1439);
nand U2018 (N_2018,In_402,In_475);
and U2019 (N_2019,In_314,In_1436);
and U2020 (N_2020,In_661,In_1016);
nor U2021 (N_2021,In_216,In_1458);
nor U2022 (N_2022,In_365,In_400);
nor U2023 (N_2023,In_653,In_680);
and U2024 (N_2024,In_18,In_492);
and U2025 (N_2025,In_185,In_1327);
or U2026 (N_2026,In_1309,In_1286);
nor U2027 (N_2027,In_776,In_169);
xor U2028 (N_2028,In_1379,In_720);
nor U2029 (N_2029,In_433,In_571);
nor U2030 (N_2030,In_1383,In_1458);
nand U2031 (N_2031,In_1021,In_232);
nor U2032 (N_2032,In_993,In_619);
or U2033 (N_2033,In_1188,In_1196);
nor U2034 (N_2034,In_736,In_468);
or U2035 (N_2035,In_2,In_1321);
nor U2036 (N_2036,In_31,In_997);
nor U2037 (N_2037,In_443,In_974);
and U2038 (N_2038,In_811,In_210);
and U2039 (N_2039,In_1434,In_845);
and U2040 (N_2040,In_775,In_153);
and U2041 (N_2041,In_1106,In_923);
and U2042 (N_2042,In_741,In_1042);
nand U2043 (N_2043,In_1296,In_1235);
nand U2044 (N_2044,In_1473,In_1296);
and U2045 (N_2045,In_938,In_388);
nor U2046 (N_2046,In_60,In_1457);
and U2047 (N_2047,In_1492,In_451);
nand U2048 (N_2048,In_1039,In_408);
or U2049 (N_2049,In_753,In_821);
and U2050 (N_2050,In_727,In_1449);
and U2051 (N_2051,In_988,In_404);
nor U2052 (N_2052,In_1272,In_198);
and U2053 (N_2053,In_122,In_288);
nand U2054 (N_2054,In_1408,In_1218);
or U2055 (N_2055,In_916,In_145);
or U2056 (N_2056,In_874,In_504);
or U2057 (N_2057,In_1473,In_1414);
nor U2058 (N_2058,In_1027,In_187);
nand U2059 (N_2059,In_991,In_983);
or U2060 (N_2060,In_347,In_747);
or U2061 (N_2061,In_443,In_1385);
nor U2062 (N_2062,In_974,In_775);
nand U2063 (N_2063,In_1340,In_551);
nor U2064 (N_2064,In_1019,In_614);
or U2065 (N_2065,In_353,In_736);
nor U2066 (N_2066,In_873,In_876);
nor U2067 (N_2067,In_1265,In_289);
nand U2068 (N_2068,In_432,In_526);
nor U2069 (N_2069,In_227,In_1204);
nor U2070 (N_2070,In_839,In_669);
and U2071 (N_2071,In_1470,In_643);
or U2072 (N_2072,In_84,In_682);
nand U2073 (N_2073,In_107,In_456);
or U2074 (N_2074,In_1072,In_110);
and U2075 (N_2075,In_1335,In_324);
and U2076 (N_2076,In_121,In_444);
nand U2077 (N_2077,In_566,In_411);
and U2078 (N_2078,In_829,In_1478);
or U2079 (N_2079,In_1295,In_1420);
and U2080 (N_2080,In_672,In_1130);
and U2081 (N_2081,In_407,In_1180);
nand U2082 (N_2082,In_1369,In_160);
xnor U2083 (N_2083,In_918,In_875);
and U2084 (N_2084,In_123,In_993);
and U2085 (N_2085,In_17,In_476);
and U2086 (N_2086,In_1095,In_888);
nand U2087 (N_2087,In_1209,In_552);
nand U2088 (N_2088,In_1276,In_1422);
nand U2089 (N_2089,In_298,In_227);
and U2090 (N_2090,In_1345,In_182);
or U2091 (N_2091,In_972,In_691);
nand U2092 (N_2092,In_337,In_898);
or U2093 (N_2093,In_230,In_1436);
nor U2094 (N_2094,In_213,In_233);
and U2095 (N_2095,In_432,In_242);
and U2096 (N_2096,In_668,In_306);
nand U2097 (N_2097,In_1183,In_1256);
nor U2098 (N_2098,In_200,In_1469);
and U2099 (N_2099,In_821,In_1044);
nand U2100 (N_2100,In_1171,In_1247);
or U2101 (N_2101,In_814,In_382);
and U2102 (N_2102,In_1488,In_1173);
nand U2103 (N_2103,In_55,In_874);
or U2104 (N_2104,In_1323,In_920);
and U2105 (N_2105,In_771,In_1092);
nand U2106 (N_2106,In_387,In_507);
nand U2107 (N_2107,In_602,In_1320);
nand U2108 (N_2108,In_65,In_563);
or U2109 (N_2109,In_732,In_156);
and U2110 (N_2110,In_124,In_158);
nor U2111 (N_2111,In_217,In_588);
nand U2112 (N_2112,In_135,In_1330);
or U2113 (N_2113,In_377,In_373);
or U2114 (N_2114,In_1392,In_299);
nor U2115 (N_2115,In_407,In_1459);
nand U2116 (N_2116,In_349,In_391);
or U2117 (N_2117,In_546,In_1295);
and U2118 (N_2118,In_1118,In_925);
nor U2119 (N_2119,In_280,In_198);
nand U2120 (N_2120,In_776,In_673);
and U2121 (N_2121,In_1268,In_135);
nand U2122 (N_2122,In_1140,In_866);
and U2123 (N_2123,In_1497,In_1352);
nor U2124 (N_2124,In_212,In_809);
nor U2125 (N_2125,In_687,In_1411);
and U2126 (N_2126,In_620,In_1146);
nand U2127 (N_2127,In_1400,In_1406);
nand U2128 (N_2128,In_346,In_1337);
nor U2129 (N_2129,In_119,In_941);
nor U2130 (N_2130,In_325,In_1185);
nor U2131 (N_2131,In_244,In_1273);
nand U2132 (N_2132,In_721,In_716);
nor U2133 (N_2133,In_907,In_1083);
or U2134 (N_2134,In_29,In_393);
nor U2135 (N_2135,In_599,In_634);
or U2136 (N_2136,In_749,In_461);
and U2137 (N_2137,In_213,In_1039);
or U2138 (N_2138,In_677,In_1351);
nand U2139 (N_2139,In_734,In_1455);
nor U2140 (N_2140,In_1494,In_1338);
or U2141 (N_2141,In_848,In_1165);
or U2142 (N_2142,In_1463,In_122);
nand U2143 (N_2143,In_1366,In_138);
nand U2144 (N_2144,In_520,In_375);
or U2145 (N_2145,In_1328,In_561);
or U2146 (N_2146,In_1057,In_548);
and U2147 (N_2147,In_1126,In_165);
nand U2148 (N_2148,In_1363,In_821);
nand U2149 (N_2149,In_1419,In_751);
nor U2150 (N_2150,In_1133,In_1380);
xnor U2151 (N_2151,In_87,In_334);
and U2152 (N_2152,In_656,In_1094);
or U2153 (N_2153,In_1212,In_1301);
or U2154 (N_2154,In_610,In_337);
or U2155 (N_2155,In_1282,In_1177);
or U2156 (N_2156,In_1198,In_187);
and U2157 (N_2157,In_945,In_1247);
and U2158 (N_2158,In_194,In_392);
nor U2159 (N_2159,In_1052,In_902);
nand U2160 (N_2160,In_493,In_273);
or U2161 (N_2161,In_1042,In_1138);
or U2162 (N_2162,In_821,In_400);
or U2163 (N_2163,In_192,In_687);
and U2164 (N_2164,In_1149,In_982);
and U2165 (N_2165,In_984,In_430);
or U2166 (N_2166,In_1006,In_1007);
and U2167 (N_2167,In_1117,In_867);
or U2168 (N_2168,In_384,In_272);
and U2169 (N_2169,In_12,In_501);
nand U2170 (N_2170,In_1166,In_158);
or U2171 (N_2171,In_983,In_172);
nand U2172 (N_2172,In_1245,In_910);
and U2173 (N_2173,In_956,In_589);
nor U2174 (N_2174,In_145,In_312);
and U2175 (N_2175,In_648,In_731);
nor U2176 (N_2176,In_1198,In_768);
nor U2177 (N_2177,In_1035,In_1072);
or U2178 (N_2178,In_137,In_1047);
or U2179 (N_2179,In_1120,In_484);
and U2180 (N_2180,In_162,In_1352);
nand U2181 (N_2181,In_795,In_78);
nand U2182 (N_2182,In_63,In_829);
nand U2183 (N_2183,In_429,In_539);
nand U2184 (N_2184,In_1325,In_197);
or U2185 (N_2185,In_636,In_1054);
and U2186 (N_2186,In_713,In_257);
nor U2187 (N_2187,In_977,In_237);
and U2188 (N_2188,In_832,In_1118);
nor U2189 (N_2189,In_637,In_521);
or U2190 (N_2190,In_650,In_393);
and U2191 (N_2191,In_349,In_871);
and U2192 (N_2192,In_142,In_662);
xor U2193 (N_2193,In_719,In_527);
or U2194 (N_2194,In_1462,In_10);
nor U2195 (N_2195,In_529,In_1294);
and U2196 (N_2196,In_864,In_901);
or U2197 (N_2197,In_1317,In_595);
or U2198 (N_2198,In_1327,In_389);
nor U2199 (N_2199,In_1428,In_540);
nand U2200 (N_2200,In_1423,In_1294);
or U2201 (N_2201,In_441,In_346);
nand U2202 (N_2202,In_781,In_1);
nand U2203 (N_2203,In_759,In_935);
and U2204 (N_2204,In_21,In_739);
nand U2205 (N_2205,In_947,In_527);
nand U2206 (N_2206,In_1006,In_799);
or U2207 (N_2207,In_1213,In_606);
nand U2208 (N_2208,In_407,In_1278);
and U2209 (N_2209,In_802,In_1270);
nand U2210 (N_2210,In_856,In_1226);
nand U2211 (N_2211,In_814,In_789);
and U2212 (N_2212,In_161,In_99);
nand U2213 (N_2213,In_164,In_613);
nand U2214 (N_2214,In_471,In_904);
or U2215 (N_2215,In_1255,In_874);
nand U2216 (N_2216,In_249,In_820);
nand U2217 (N_2217,In_92,In_74);
or U2218 (N_2218,In_1153,In_760);
nand U2219 (N_2219,In_869,In_148);
and U2220 (N_2220,In_916,In_408);
nor U2221 (N_2221,In_473,In_1499);
nand U2222 (N_2222,In_1419,In_748);
nor U2223 (N_2223,In_936,In_1014);
or U2224 (N_2224,In_1306,In_615);
nand U2225 (N_2225,In_732,In_1204);
nand U2226 (N_2226,In_1039,In_1369);
or U2227 (N_2227,In_1032,In_443);
and U2228 (N_2228,In_1104,In_586);
nor U2229 (N_2229,In_1291,In_1072);
nor U2230 (N_2230,In_672,In_1306);
or U2231 (N_2231,In_987,In_1181);
xnor U2232 (N_2232,In_1172,In_505);
and U2233 (N_2233,In_473,In_1201);
nand U2234 (N_2234,In_813,In_1257);
xor U2235 (N_2235,In_327,In_53);
and U2236 (N_2236,In_1174,In_428);
nor U2237 (N_2237,In_650,In_460);
and U2238 (N_2238,In_1218,In_510);
or U2239 (N_2239,In_186,In_803);
and U2240 (N_2240,In_209,In_579);
nand U2241 (N_2241,In_208,In_14);
nand U2242 (N_2242,In_110,In_856);
or U2243 (N_2243,In_406,In_1486);
or U2244 (N_2244,In_391,In_651);
nand U2245 (N_2245,In_63,In_718);
or U2246 (N_2246,In_1039,In_1361);
or U2247 (N_2247,In_263,In_1011);
nor U2248 (N_2248,In_1435,In_907);
nor U2249 (N_2249,In_1369,In_328);
nand U2250 (N_2250,In_208,In_933);
xor U2251 (N_2251,In_481,In_271);
nor U2252 (N_2252,In_921,In_1429);
and U2253 (N_2253,In_617,In_1284);
nand U2254 (N_2254,In_27,In_285);
or U2255 (N_2255,In_717,In_1009);
and U2256 (N_2256,In_1323,In_1387);
and U2257 (N_2257,In_227,In_185);
and U2258 (N_2258,In_139,In_647);
nand U2259 (N_2259,In_1483,In_1137);
nor U2260 (N_2260,In_909,In_1040);
and U2261 (N_2261,In_1284,In_79);
and U2262 (N_2262,In_1116,In_252);
and U2263 (N_2263,In_564,In_1055);
and U2264 (N_2264,In_10,In_770);
nor U2265 (N_2265,In_254,In_528);
nor U2266 (N_2266,In_213,In_495);
nand U2267 (N_2267,In_1059,In_1278);
nor U2268 (N_2268,In_1006,In_1427);
nor U2269 (N_2269,In_1051,In_730);
or U2270 (N_2270,In_27,In_104);
nand U2271 (N_2271,In_586,In_128);
nor U2272 (N_2272,In_140,In_1303);
nor U2273 (N_2273,In_1459,In_767);
nor U2274 (N_2274,In_1416,In_1200);
nand U2275 (N_2275,In_742,In_172);
or U2276 (N_2276,In_751,In_1214);
nand U2277 (N_2277,In_648,In_182);
and U2278 (N_2278,In_414,In_565);
nor U2279 (N_2279,In_1330,In_372);
nor U2280 (N_2280,In_1021,In_803);
nand U2281 (N_2281,In_333,In_962);
and U2282 (N_2282,In_1096,In_585);
or U2283 (N_2283,In_1151,In_478);
or U2284 (N_2284,In_1272,In_81);
nand U2285 (N_2285,In_1033,In_1293);
and U2286 (N_2286,In_50,In_209);
nor U2287 (N_2287,In_710,In_782);
nand U2288 (N_2288,In_127,In_621);
nand U2289 (N_2289,In_553,In_1446);
or U2290 (N_2290,In_952,In_523);
nand U2291 (N_2291,In_1490,In_501);
nor U2292 (N_2292,In_955,In_1122);
or U2293 (N_2293,In_910,In_1328);
xnor U2294 (N_2294,In_1358,In_494);
nor U2295 (N_2295,In_1198,In_490);
nor U2296 (N_2296,In_1489,In_398);
and U2297 (N_2297,In_1318,In_1124);
or U2298 (N_2298,In_759,In_401);
and U2299 (N_2299,In_430,In_126);
nor U2300 (N_2300,In_748,In_860);
nand U2301 (N_2301,In_1080,In_1112);
and U2302 (N_2302,In_965,In_669);
nor U2303 (N_2303,In_495,In_461);
or U2304 (N_2304,In_825,In_265);
nand U2305 (N_2305,In_1113,In_1017);
nand U2306 (N_2306,In_710,In_1027);
and U2307 (N_2307,In_899,In_420);
nor U2308 (N_2308,In_735,In_1171);
or U2309 (N_2309,In_722,In_1210);
nor U2310 (N_2310,In_879,In_1415);
nor U2311 (N_2311,In_1261,In_200);
or U2312 (N_2312,In_451,In_653);
nand U2313 (N_2313,In_378,In_1190);
or U2314 (N_2314,In_813,In_1296);
xnor U2315 (N_2315,In_932,In_399);
nand U2316 (N_2316,In_992,In_697);
or U2317 (N_2317,In_1264,In_1162);
or U2318 (N_2318,In_1363,In_997);
or U2319 (N_2319,In_539,In_1184);
and U2320 (N_2320,In_661,In_329);
and U2321 (N_2321,In_510,In_1498);
and U2322 (N_2322,In_384,In_1404);
and U2323 (N_2323,In_80,In_1110);
and U2324 (N_2324,In_918,In_822);
nand U2325 (N_2325,In_1101,In_1439);
nand U2326 (N_2326,In_619,In_17);
nor U2327 (N_2327,In_770,In_110);
nand U2328 (N_2328,In_120,In_744);
nor U2329 (N_2329,In_245,In_483);
or U2330 (N_2330,In_897,In_623);
nand U2331 (N_2331,In_573,In_1422);
nor U2332 (N_2332,In_461,In_289);
and U2333 (N_2333,In_1363,In_990);
nor U2334 (N_2334,In_335,In_41);
or U2335 (N_2335,In_372,In_1438);
nor U2336 (N_2336,In_345,In_56);
nand U2337 (N_2337,In_902,In_175);
nor U2338 (N_2338,In_1289,In_292);
nor U2339 (N_2339,In_29,In_57);
or U2340 (N_2340,In_266,In_105);
nor U2341 (N_2341,In_1287,In_868);
xor U2342 (N_2342,In_1193,In_340);
or U2343 (N_2343,In_848,In_784);
nor U2344 (N_2344,In_1154,In_1231);
or U2345 (N_2345,In_1273,In_667);
or U2346 (N_2346,In_13,In_1066);
or U2347 (N_2347,In_920,In_1216);
nor U2348 (N_2348,In_692,In_258);
or U2349 (N_2349,In_137,In_1480);
or U2350 (N_2350,In_909,In_837);
nor U2351 (N_2351,In_1274,In_440);
or U2352 (N_2352,In_366,In_834);
or U2353 (N_2353,In_999,In_567);
nor U2354 (N_2354,In_953,In_130);
nor U2355 (N_2355,In_485,In_81);
or U2356 (N_2356,In_1240,In_1254);
or U2357 (N_2357,In_100,In_818);
or U2358 (N_2358,In_1147,In_887);
or U2359 (N_2359,In_666,In_561);
nand U2360 (N_2360,In_284,In_710);
or U2361 (N_2361,In_416,In_669);
and U2362 (N_2362,In_1493,In_747);
xnor U2363 (N_2363,In_791,In_516);
nor U2364 (N_2364,In_1409,In_627);
or U2365 (N_2365,In_1300,In_743);
or U2366 (N_2366,In_1331,In_284);
nand U2367 (N_2367,In_1158,In_301);
or U2368 (N_2368,In_299,In_645);
and U2369 (N_2369,In_1450,In_697);
nand U2370 (N_2370,In_1281,In_1056);
nand U2371 (N_2371,In_896,In_582);
or U2372 (N_2372,In_706,In_577);
nand U2373 (N_2373,In_52,In_224);
and U2374 (N_2374,In_228,In_913);
nor U2375 (N_2375,In_149,In_770);
nand U2376 (N_2376,In_1484,In_1108);
nand U2377 (N_2377,In_59,In_108);
and U2378 (N_2378,In_1317,In_898);
and U2379 (N_2379,In_78,In_281);
or U2380 (N_2380,In_1301,In_1050);
nand U2381 (N_2381,In_549,In_1121);
or U2382 (N_2382,In_668,In_863);
and U2383 (N_2383,In_165,In_944);
and U2384 (N_2384,In_327,In_1168);
nor U2385 (N_2385,In_410,In_113);
nand U2386 (N_2386,In_832,In_603);
nand U2387 (N_2387,In_106,In_628);
nor U2388 (N_2388,In_819,In_799);
and U2389 (N_2389,In_923,In_378);
and U2390 (N_2390,In_823,In_1028);
or U2391 (N_2391,In_534,In_883);
and U2392 (N_2392,In_173,In_770);
nand U2393 (N_2393,In_361,In_291);
and U2394 (N_2394,In_97,In_1403);
or U2395 (N_2395,In_462,In_164);
and U2396 (N_2396,In_1010,In_1436);
nand U2397 (N_2397,In_1432,In_211);
nand U2398 (N_2398,In_1103,In_333);
and U2399 (N_2399,In_743,In_1313);
nor U2400 (N_2400,In_905,In_678);
nand U2401 (N_2401,In_364,In_395);
and U2402 (N_2402,In_1291,In_1086);
and U2403 (N_2403,In_86,In_663);
nand U2404 (N_2404,In_86,In_1075);
or U2405 (N_2405,In_816,In_998);
nand U2406 (N_2406,In_1183,In_1040);
nand U2407 (N_2407,In_70,In_1016);
nor U2408 (N_2408,In_212,In_903);
nor U2409 (N_2409,In_668,In_96);
and U2410 (N_2410,In_706,In_1017);
nor U2411 (N_2411,In_283,In_608);
nor U2412 (N_2412,In_986,In_360);
and U2413 (N_2413,In_40,In_1478);
nor U2414 (N_2414,In_1164,In_1079);
nor U2415 (N_2415,In_834,In_1448);
and U2416 (N_2416,In_709,In_1172);
and U2417 (N_2417,In_720,In_1350);
and U2418 (N_2418,In_1158,In_471);
nand U2419 (N_2419,In_293,In_1476);
or U2420 (N_2420,In_93,In_1327);
nand U2421 (N_2421,In_1383,In_142);
nand U2422 (N_2422,In_330,In_99);
and U2423 (N_2423,In_74,In_481);
nand U2424 (N_2424,In_118,In_1415);
and U2425 (N_2425,In_48,In_906);
nand U2426 (N_2426,In_1186,In_1105);
xor U2427 (N_2427,In_352,In_125);
or U2428 (N_2428,In_150,In_241);
nor U2429 (N_2429,In_1397,In_1265);
nor U2430 (N_2430,In_889,In_1149);
nand U2431 (N_2431,In_409,In_702);
nor U2432 (N_2432,In_1389,In_6);
or U2433 (N_2433,In_1199,In_994);
nand U2434 (N_2434,In_1346,In_539);
nor U2435 (N_2435,In_1188,In_1265);
nand U2436 (N_2436,In_130,In_1424);
nor U2437 (N_2437,In_58,In_1002);
nor U2438 (N_2438,In_560,In_141);
and U2439 (N_2439,In_817,In_17);
nor U2440 (N_2440,In_1209,In_1043);
or U2441 (N_2441,In_420,In_529);
and U2442 (N_2442,In_1465,In_200);
nand U2443 (N_2443,In_841,In_870);
nand U2444 (N_2444,In_662,In_43);
nor U2445 (N_2445,In_151,In_564);
or U2446 (N_2446,In_631,In_358);
or U2447 (N_2447,In_968,In_898);
and U2448 (N_2448,In_806,In_920);
nor U2449 (N_2449,In_95,In_572);
and U2450 (N_2450,In_1091,In_155);
nand U2451 (N_2451,In_952,In_766);
nor U2452 (N_2452,In_752,In_1234);
or U2453 (N_2453,In_386,In_706);
and U2454 (N_2454,In_1008,In_279);
nand U2455 (N_2455,In_637,In_42);
and U2456 (N_2456,In_1370,In_893);
and U2457 (N_2457,In_1068,In_945);
and U2458 (N_2458,In_528,In_1060);
and U2459 (N_2459,In_875,In_372);
nand U2460 (N_2460,In_1095,In_638);
nor U2461 (N_2461,In_608,In_1264);
and U2462 (N_2462,In_544,In_152);
nand U2463 (N_2463,In_1125,In_145);
and U2464 (N_2464,In_230,In_1265);
nand U2465 (N_2465,In_366,In_390);
or U2466 (N_2466,In_1198,In_940);
or U2467 (N_2467,In_412,In_808);
and U2468 (N_2468,In_1050,In_543);
and U2469 (N_2469,In_1075,In_910);
nand U2470 (N_2470,In_886,In_196);
or U2471 (N_2471,In_1379,In_584);
and U2472 (N_2472,In_709,In_458);
and U2473 (N_2473,In_1322,In_1225);
and U2474 (N_2474,In_548,In_576);
or U2475 (N_2475,In_158,In_572);
and U2476 (N_2476,In_1137,In_331);
nor U2477 (N_2477,In_1214,In_246);
or U2478 (N_2478,In_716,In_94);
nand U2479 (N_2479,In_701,In_667);
or U2480 (N_2480,In_92,In_1101);
and U2481 (N_2481,In_249,In_113);
and U2482 (N_2482,In_639,In_227);
nor U2483 (N_2483,In_204,In_962);
xor U2484 (N_2484,In_18,In_1206);
or U2485 (N_2485,In_573,In_1356);
nor U2486 (N_2486,In_233,In_1267);
and U2487 (N_2487,In_323,In_231);
nand U2488 (N_2488,In_645,In_323);
or U2489 (N_2489,In_1435,In_628);
or U2490 (N_2490,In_867,In_445);
nor U2491 (N_2491,In_996,In_23);
or U2492 (N_2492,In_278,In_105);
nand U2493 (N_2493,In_1483,In_1097);
nand U2494 (N_2494,In_700,In_1125);
or U2495 (N_2495,In_1424,In_959);
nand U2496 (N_2496,In_1337,In_1204);
and U2497 (N_2497,In_974,In_1284);
nor U2498 (N_2498,In_151,In_1284);
nand U2499 (N_2499,In_351,In_595);
or U2500 (N_2500,In_1294,In_1203);
nand U2501 (N_2501,In_53,In_614);
nand U2502 (N_2502,In_182,In_339);
and U2503 (N_2503,In_1202,In_934);
nand U2504 (N_2504,In_1217,In_830);
nand U2505 (N_2505,In_88,In_1083);
nor U2506 (N_2506,In_514,In_613);
and U2507 (N_2507,In_1143,In_1274);
or U2508 (N_2508,In_1141,In_645);
or U2509 (N_2509,In_261,In_430);
nor U2510 (N_2510,In_1122,In_1219);
or U2511 (N_2511,In_912,In_746);
and U2512 (N_2512,In_1423,In_810);
and U2513 (N_2513,In_1268,In_1327);
nand U2514 (N_2514,In_857,In_994);
nor U2515 (N_2515,In_1346,In_686);
nor U2516 (N_2516,In_650,In_842);
nand U2517 (N_2517,In_938,In_1019);
or U2518 (N_2518,In_120,In_841);
nand U2519 (N_2519,In_324,In_1163);
nor U2520 (N_2520,In_1259,In_1181);
nor U2521 (N_2521,In_643,In_756);
and U2522 (N_2522,In_911,In_443);
nor U2523 (N_2523,In_1143,In_1209);
nor U2524 (N_2524,In_383,In_7);
and U2525 (N_2525,In_593,In_955);
or U2526 (N_2526,In_947,In_530);
nand U2527 (N_2527,In_738,In_1430);
nand U2528 (N_2528,In_904,In_1283);
or U2529 (N_2529,In_58,In_1220);
and U2530 (N_2530,In_101,In_946);
nor U2531 (N_2531,In_177,In_694);
nand U2532 (N_2532,In_428,In_1138);
and U2533 (N_2533,In_305,In_623);
nand U2534 (N_2534,In_631,In_904);
and U2535 (N_2535,In_995,In_1247);
or U2536 (N_2536,In_55,In_1403);
nand U2537 (N_2537,In_463,In_1303);
nor U2538 (N_2538,In_868,In_332);
and U2539 (N_2539,In_19,In_545);
nor U2540 (N_2540,In_1305,In_244);
or U2541 (N_2541,In_988,In_426);
nand U2542 (N_2542,In_281,In_371);
or U2543 (N_2543,In_320,In_425);
or U2544 (N_2544,In_1218,In_741);
and U2545 (N_2545,In_900,In_1201);
nor U2546 (N_2546,In_808,In_803);
nor U2547 (N_2547,In_1479,In_1002);
and U2548 (N_2548,In_680,In_659);
nand U2549 (N_2549,In_1360,In_1289);
and U2550 (N_2550,In_105,In_451);
xnor U2551 (N_2551,In_100,In_117);
nand U2552 (N_2552,In_270,In_1121);
and U2553 (N_2553,In_227,In_981);
or U2554 (N_2554,In_3,In_889);
or U2555 (N_2555,In_45,In_669);
or U2556 (N_2556,In_582,In_562);
nand U2557 (N_2557,In_571,In_711);
nand U2558 (N_2558,In_960,In_763);
xnor U2559 (N_2559,In_1103,In_1002);
nand U2560 (N_2560,In_684,In_48);
or U2561 (N_2561,In_1175,In_13);
and U2562 (N_2562,In_1432,In_1451);
or U2563 (N_2563,In_641,In_1235);
nor U2564 (N_2564,In_1498,In_496);
and U2565 (N_2565,In_829,In_1258);
and U2566 (N_2566,In_1401,In_219);
nand U2567 (N_2567,In_49,In_1077);
nor U2568 (N_2568,In_539,In_590);
nand U2569 (N_2569,In_88,In_220);
nor U2570 (N_2570,In_443,In_324);
nand U2571 (N_2571,In_926,In_463);
nor U2572 (N_2572,In_560,In_325);
or U2573 (N_2573,In_462,In_315);
nand U2574 (N_2574,In_816,In_1441);
and U2575 (N_2575,In_1468,In_1107);
or U2576 (N_2576,In_115,In_2);
nor U2577 (N_2577,In_594,In_506);
or U2578 (N_2578,In_635,In_247);
nor U2579 (N_2579,In_327,In_94);
nand U2580 (N_2580,In_532,In_420);
and U2581 (N_2581,In_27,In_1211);
nand U2582 (N_2582,In_657,In_1082);
nand U2583 (N_2583,In_1280,In_45);
nand U2584 (N_2584,In_313,In_662);
or U2585 (N_2585,In_1147,In_1415);
or U2586 (N_2586,In_1291,In_1195);
and U2587 (N_2587,In_1047,In_1433);
or U2588 (N_2588,In_197,In_516);
and U2589 (N_2589,In_468,In_533);
nand U2590 (N_2590,In_755,In_1363);
and U2591 (N_2591,In_663,In_246);
xor U2592 (N_2592,In_1000,In_970);
and U2593 (N_2593,In_647,In_1003);
and U2594 (N_2594,In_892,In_723);
nand U2595 (N_2595,In_1199,In_891);
nand U2596 (N_2596,In_828,In_323);
and U2597 (N_2597,In_926,In_370);
and U2598 (N_2598,In_1436,In_39);
nand U2599 (N_2599,In_552,In_1446);
nand U2600 (N_2600,In_1317,In_832);
nor U2601 (N_2601,In_40,In_665);
and U2602 (N_2602,In_1274,In_558);
nor U2603 (N_2603,In_60,In_52);
nand U2604 (N_2604,In_496,In_876);
nor U2605 (N_2605,In_181,In_1423);
and U2606 (N_2606,In_887,In_1472);
and U2607 (N_2607,In_826,In_988);
and U2608 (N_2608,In_693,In_1451);
or U2609 (N_2609,In_545,In_1309);
nor U2610 (N_2610,In_1345,In_500);
and U2611 (N_2611,In_424,In_197);
and U2612 (N_2612,In_1489,In_216);
nand U2613 (N_2613,In_655,In_1389);
or U2614 (N_2614,In_1344,In_432);
and U2615 (N_2615,In_106,In_477);
and U2616 (N_2616,In_698,In_1357);
and U2617 (N_2617,In_96,In_127);
nor U2618 (N_2618,In_1182,In_836);
or U2619 (N_2619,In_1433,In_5);
nor U2620 (N_2620,In_1128,In_151);
nand U2621 (N_2621,In_236,In_1208);
or U2622 (N_2622,In_440,In_1405);
nand U2623 (N_2623,In_941,In_345);
nor U2624 (N_2624,In_312,In_126);
and U2625 (N_2625,In_1208,In_579);
or U2626 (N_2626,In_1069,In_1165);
nand U2627 (N_2627,In_602,In_989);
nor U2628 (N_2628,In_1470,In_1434);
or U2629 (N_2629,In_1466,In_357);
nor U2630 (N_2630,In_490,In_1143);
nand U2631 (N_2631,In_397,In_1155);
and U2632 (N_2632,In_15,In_212);
nor U2633 (N_2633,In_1173,In_904);
nand U2634 (N_2634,In_1162,In_819);
and U2635 (N_2635,In_785,In_41);
nor U2636 (N_2636,In_743,In_1052);
or U2637 (N_2637,In_514,In_713);
nor U2638 (N_2638,In_315,In_1185);
nand U2639 (N_2639,In_368,In_574);
or U2640 (N_2640,In_191,In_980);
nand U2641 (N_2641,In_1222,In_839);
nand U2642 (N_2642,In_1246,In_821);
nor U2643 (N_2643,In_1244,In_727);
or U2644 (N_2644,In_752,In_99);
nand U2645 (N_2645,In_388,In_573);
or U2646 (N_2646,In_1050,In_375);
or U2647 (N_2647,In_66,In_1001);
nor U2648 (N_2648,In_330,In_407);
and U2649 (N_2649,In_1138,In_75);
or U2650 (N_2650,In_710,In_1403);
and U2651 (N_2651,In_706,In_11);
or U2652 (N_2652,In_1274,In_760);
nand U2653 (N_2653,In_142,In_47);
nor U2654 (N_2654,In_675,In_936);
nor U2655 (N_2655,In_799,In_254);
xnor U2656 (N_2656,In_1123,In_1346);
or U2657 (N_2657,In_226,In_51);
or U2658 (N_2658,In_1351,In_54);
and U2659 (N_2659,In_371,In_1207);
or U2660 (N_2660,In_617,In_638);
nor U2661 (N_2661,In_926,In_1005);
and U2662 (N_2662,In_423,In_1365);
and U2663 (N_2663,In_959,In_1047);
or U2664 (N_2664,In_359,In_1252);
xnor U2665 (N_2665,In_949,In_687);
or U2666 (N_2666,In_417,In_459);
nor U2667 (N_2667,In_450,In_1251);
and U2668 (N_2668,In_1051,In_589);
nand U2669 (N_2669,In_1101,In_1299);
and U2670 (N_2670,In_436,In_432);
nand U2671 (N_2671,In_1494,In_252);
nor U2672 (N_2672,In_895,In_644);
nor U2673 (N_2673,In_533,In_702);
nand U2674 (N_2674,In_1055,In_1160);
or U2675 (N_2675,In_1260,In_568);
or U2676 (N_2676,In_1242,In_1453);
and U2677 (N_2677,In_1076,In_1241);
or U2678 (N_2678,In_755,In_442);
nor U2679 (N_2679,In_766,In_1134);
or U2680 (N_2680,In_333,In_255);
or U2681 (N_2681,In_115,In_313);
and U2682 (N_2682,In_1201,In_949);
nand U2683 (N_2683,In_529,In_59);
nand U2684 (N_2684,In_1108,In_652);
nor U2685 (N_2685,In_1381,In_571);
nor U2686 (N_2686,In_842,In_876);
nand U2687 (N_2687,In_666,In_437);
nand U2688 (N_2688,In_401,In_876);
nor U2689 (N_2689,In_389,In_1059);
or U2690 (N_2690,In_965,In_312);
nor U2691 (N_2691,In_373,In_880);
nand U2692 (N_2692,In_1025,In_1073);
nand U2693 (N_2693,In_900,In_1285);
and U2694 (N_2694,In_425,In_775);
and U2695 (N_2695,In_1027,In_1325);
nand U2696 (N_2696,In_517,In_412);
nor U2697 (N_2697,In_418,In_703);
nand U2698 (N_2698,In_91,In_870);
or U2699 (N_2699,In_674,In_180);
nor U2700 (N_2700,In_1106,In_1001);
and U2701 (N_2701,In_301,In_229);
or U2702 (N_2702,In_245,In_65);
or U2703 (N_2703,In_1356,In_458);
nand U2704 (N_2704,In_930,In_938);
nor U2705 (N_2705,In_1468,In_1178);
and U2706 (N_2706,In_43,In_1494);
and U2707 (N_2707,In_1235,In_738);
nand U2708 (N_2708,In_56,In_1366);
nor U2709 (N_2709,In_1114,In_1035);
xnor U2710 (N_2710,In_666,In_879);
or U2711 (N_2711,In_214,In_1002);
or U2712 (N_2712,In_816,In_490);
and U2713 (N_2713,In_292,In_891);
or U2714 (N_2714,In_584,In_1374);
or U2715 (N_2715,In_444,In_825);
or U2716 (N_2716,In_467,In_595);
nor U2717 (N_2717,In_188,In_210);
nor U2718 (N_2718,In_306,In_940);
nor U2719 (N_2719,In_741,In_297);
nor U2720 (N_2720,In_646,In_223);
nand U2721 (N_2721,In_60,In_1140);
and U2722 (N_2722,In_993,In_1276);
nand U2723 (N_2723,In_3,In_440);
and U2724 (N_2724,In_1282,In_853);
and U2725 (N_2725,In_449,In_687);
nand U2726 (N_2726,In_777,In_819);
and U2727 (N_2727,In_1259,In_750);
and U2728 (N_2728,In_504,In_1413);
nor U2729 (N_2729,In_60,In_551);
nand U2730 (N_2730,In_1315,In_515);
and U2731 (N_2731,In_688,In_105);
nand U2732 (N_2732,In_723,In_372);
or U2733 (N_2733,In_179,In_1461);
and U2734 (N_2734,In_1094,In_1297);
or U2735 (N_2735,In_854,In_58);
and U2736 (N_2736,In_45,In_633);
and U2737 (N_2737,In_332,In_1019);
and U2738 (N_2738,In_287,In_80);
and U2739 (N_2739,In_556,In_1003);
or U2740 (N_2740,In_679,In_354);
and U2741 (N_2741,In_1459,In_1443);
or U2742 (N_2742,In_96,In_410);
or U2743 (N_2743,In_448,In_740);
nand U2744 (N_2744,In_30,In_830);
nor U2745 (N_2745,In_1363,In_1326);
nor U2746 (N_2746,In_1308,In_168);
or U2747 (N_2747,In_1444,In_575);
xor U2748 (N_2748,In_825,In_1231);
nand U2749 (N_2749,In_879,In_532);
or U2750 (N_2750,In_607,In_406);
and U2751 (N_2751,In_1204,In_623);
or U2752 (N_2752,In_29,In_651);
nand U2753 (N_2753,In_1262,In_5);
and U2754 (N_2754,In_1304,In_780);
nor U2755 (N_2755,In_550,In_707);
nor U2756 (N_2756,In_894,In_845);
or U2757 (N_2757,In_1289,In_1499);
nand U2758 (N_2758,In_727,In_793);
nand U2759 (N_2759,In_543,In_628);
and U2760 (N_2760,In_845,In_661);
or U2761 (N_2761,In_1024,In_1093);
or U2762 (N_2762,In_527,In_1481);
and U2763 (N_2763,In_428,In_1092);
and U2764 (N_2764,In_11,In_1070);
nor U2765 (N_2765,In_215,In_611);
or U2766 (N_2766,In_1343,In_1413);
and U2767 (N_2767,In_797,In_107);
nand U2768 (N_2768,In_852,In_543);
or U2769 (N_2769,In_457,In_1210);
or U2770 (N_2770,In_252,In_665);
nand U2771 (N_2771,In_1471,In_890);
and U2772 (N_2772,In_76,In_33);
nor U2773 (N_2773,In_1150,In_284);
or U2774 (N_2774,In_389,In_27);
nand U2775 (N_2775,In_194,In_1461);
nor U2776 (N_2776,In_828,In_481);
nor U2777 (N_2777,In_170,In_1480);
nand U2778 (N_2778,In_17,In_1097);
or U2779 (N_2779,In_1040,In_1126);
nor U2780 (N_2780,In_551,In_230);
nand U2781 (N_2781,In_781,In_42);
or U2782 (N_2782,In_852,In_436);
or U2783 (N_2783,In_812,In_1240);
nand U2784 (N_2784,In_137,In_1289);
nand U2785 (N_2785,In_123,In_433);
nand U2786 (N_2786,In_1332,In_1222);
nand U2787 (N_2787,In_1230,In_680);
nand U2788 (N_2788,In_578,In_1237);
nand U2789 (N_2789,In_808,In_290);
or U2790 (N_2790,In_324,In_629);
or U2791 (N_2791,In_456,In_72);
nor U2792 (N_2792,In_1081,In_13);
xor U2793 (N_2793,In_184,In_1324);
and U2794 (N_2794,In_1133,In_201);
and U2795 (N_2795,In_109,In_985);
or U2796 (N_2796,In_963,In_614);
or U2797 (N_2797,In_1460,In_1153);
nand U2798 (N_2798,In_230,In_1315);
and U2799 (N_2799,In_571,In_367);
and U2800 (N_2800,In_509,In_308);
or U2801 (N_2801,In_475,In_119);
and U2802 (N_2802,In_359,In_28);
nand U2803 (N_2803,In_561,In_418);
nand U2804 (N_2804,In_1343,In_861);
or U2805 (N_2805,In_592,In_1127);
nand U2806 (N_2806,In_1219,In_373);
nor U2807 (N_2807,In_653,In_937);
nand U2808 (N_2808,In_1276,In_1334);
nor U2809 (N_2809,In_1144,In_1464);
nor U2810 (N_2810,In_249,In_328);
and U2811 (N_2811,In_403,In_1147);
nor U2812 (N_2812,In_987,In_1305);
and U2813 (N_2813,In_1439,In_362);
or U2814 (N_2814,In_501,In_1177);
nor U2815 (N_2815,In_223,In_130);
nor U2816 (N_2816,In_37,In_169);
and U2817 (N_2817,In_218,In_391);
nand U2818 (N_2818,In_791,In_147);
and U2819 (N_2819,In_878,In_999);
and U2820 (N_2820,In_916,In_1121);
nand U2821 (N_2821,In_1276,In_883);
and U2822 (N_2822,In_564,In_170);
or U2823 (N_2823,In_1451,In_181);
nor U2824 (N_2824,In_1268,In_1273);
or U2825 (N_2825,In_264,In_7);
nor U2826 (N_2826,In_215,In_1437);
nand U2827 (N_2827,In_526,In_813);
nor U2828 (N_2828,In_1329,In_432);
or U2829 (N_2829,In_838,In_1426);
nor U2830 (N_2830,In_567,In_1141);
and U2831 (N_2831,In_547,In_300);
nor U2832 (N_2832,In_695,In_318);
nand U2833 (N_2833,In_444,In_811);
nor U2834 (N_2834,In_490,In_819);
nand U2835 (N_2835,In_973,In_650);
nor U2836 (N_2836,In_1008,In_1190);
nand U2837 (N_2837,In_719,In_367);
nor U2838 (N_2838,In_445,In_1180);
and U2839 (N_2839,In_698,In_754);
and U2840 (N_2840,In_133,In_1324);
nand U2841 (N_2841,In_897,In_836);
nor U2842 (N_2842,In_648,In_1086);
and U2843 (N_2843,In_682,In_211);
nand U2844 (N_2844,In_466,In_1263);
and U2845 (N_2845,In_60,In_1019);
or U2846 (N_2846,In_846,In_1394);
or U2847 (N_2847,In_1167,In_954);
and U2848 (N_2848,In_1243,In_449);
nor U2849 (N_2849,In_108,In_623);
nor U2850 (N_2850,In_196,In_357);
nand U2851 (N_2851,In_1432,In_10);
or U2852 (N_2852,In_695,In_404);
nand U2853 (N_2853,In_360,In_924);
nor U2854 (N_2854,In_20,In_723);
and U2855 (N_2855,In_554,In_551);
nand U2856 (N_2856,In_80,In_583);
nand U2857 (N_2857,In_806,In_1181);
nand U2858 (N_2858,In_1398,In_545);
and U2859 (N_2859,In_1081,In_367);
and U2860 (N_2860,In_966,In_659);
nor U2861 (N_2861,In_29,In_1108);
and U2862 (N_2862,In_1268,In_652);
nand U2863 (N_2863,In_519,In_989);
nor U2864 (N_2864,In_191,In_908);
and U2865 (N_2865,In_1043,In_791);
and U2866 (N_2866,In_763,In_594);
and U2867 (N_2867,In_147,In_1284);
or U2868 (N_2868,In_693,In_759);
nand U2869 (N_2869,In_1329,In_1415);
or U2870 (N_2870,In_100,In_365);
or U2871 (N_2871,In_154,In_1293);
or U2872 (N_2872,In_307,In_111);
and U2873 (N_2873,In_1007,In_55);
or U2874 (N_2874,In_138,In_328);
and U2875 (N_2875,In_1126,In_983);
and U2876 (N_2876,In_1265,In_995);
xor U2877 (N_2877,In_972,In_678);
nand U2878 (N_2878,In_859,In_919);
nor U2879 (N_2879,In_1042,In_1380);
nor U2880 (N_2880,In_23,In_1054);
nor U2881 (N_2881,In_431,In_4);
or U2882 (N_2882,In_1482,In_1400);
and U2883 (N_2883,In_590,In_1108);
or U2884 (N_2884,In_1189,In_1299);
nor U2885 (N_2885,In_265,In_425);
nand U2886 (N_2886,In_1287,In_1467);
or U2887 (N_2887,In_957,In_280);
or U2888 (N_2888,In_217,In_119);
nand U2889 (N_2889,In_1479,In_634);
or U2890 (N_2890,In_787,In_977);
nand U2891 (N_2891,In_59,In_526);
or U2892 (N_2892,In_322,In_639);
nand U2893 (N_2893,In_1381,In_554);
or U2894 (N_2894,In_89,In_613);
or U2895 (N_2895,In_978,In_793);
xor U2896 (N_2896,In_1246,In_1293);
nand U2897 (N_2897,In_1087,In_970);
nand U2898 (N_2898,In_1440,In_962);
nand U2899 (N_2899,In_1033,In_1292);
nand U2900 (N_2900,In_228,In_1499);
or U2901 (N_2901,In_242,In_1323);
nand U2902 (N_2902,In_1228,In_313);
and U2903 (N_2903,In_475,In_1122);
nand U2904 (N_2904,In_514,In_1135);
nor U2905 (N_2905,In_891,In_1448);
nand U2906 (N_2906,In_764,In_963);
nand U2907 (N_2907,In_349,In_938);
and U2908 (N_2908,In_259,In_447);
nand U2909 (N_2909,In_1457,In_683);
nand U2910 (N_2910,In_414,In_377);
and U2911 (N_2911,In_665,In_1414);
nand U2912 (N_2912,In_786,In_768);
nor U2913 (N_2913,In_876,In_685);
or U2914 (N_2914,In_417,In_1461);
and U2915 (N_2915,In_582,In_563);
and U2916 (N_2916,In_926,In_1075);
and U2917 (N_2917,In_937,In_77);
and U2918 (N_2918,In_1034,In_1051);
nor U2919 (N_2919,In_114,In_1401);
and U2920 (N_2920,In_847,In_503);
nand U2921 (N_2921,In_987,In_1091);
and U2922 (N_2922,In_709,In_1220);
or U2923 (N_2923,In_1070,In_1030);
nor U2924 (N_2924,In_774,In_442);
or U2925 (N_2925,In_947,In_1220);
nand U2926 (N_2926,In_879,In_1232);
nand U2927 (N_2927,In_286,In_291);
and U2928 (N_2928,In_353,In_232);
or U2929 (N_2929,In_920,In_685);
or U2930 (N_2930,In_918,In_1304);
and U2931 (N_2931,In_156,In_1070);
nand U2932 (N_2932,In_877,In_1004);
or U2933 (N_2933,In_345,In_201);
and U2934 (N_2934,In_48,In_230);
or U2935 (N_2935,In_582,In_54);
or U2936 (N_2936,In_479,In_1051);
nor U2937 (N_2937,In_284,In_201);
or U2938 (N_2938,In_1283,In_993);
nor U2939 (N_2939,In_209,In_899);
xor U2940 (N_2940,In_684,In_844);
nand U2941 (N_2941,In_44,In_991);
and U2942 (N_2942,In_1322,In_19);
or U2943 (N_2943,In_1235,In_1009);
or U2944 (N_2944,In_184,In_1329);
nor U2945 (N_2945,In_1364,In_970);
nor U2946 (N_2946,In_1280,In_384);
or U2947 (N_2947,In_1101,In_452);
and U2948 (N_2948,In_830,In_159);
nand U2949 (N_2949,In_512,In_86);
or U2950 (N_2950,In_1243,In_140);
nand U2951 (N_2951,In_554,In_1280);
nand U2952 (N_2952,In_1130,In_14);
or U2953 (N_2953,In_1137,In_667);
or U2954 (N_2954,In_1116,In_851);
nand U2955 (N_2955,In_720,In_618);
nor U2956 (N_2956,In_46,In_559);
nor U2957 (N_2957,In_1182,In_1129);
nand U2958 (N_2958,In_490,In_995);
and U2959 (N_2959,In_950,In_1275);
and U2960 (N_2960,In_1127,In_964);
nor U2961 (N_2961,In_865,In_1374);
or U2962 (N_2962,In_804,In_80);
nor U2963 (N_2963,In_171,In_801);
nand U2964 (N_2964,In_96,In_1476);
nand U2965 (N_2965,In_1421,In_1355);
nand U2966 (N_2966,In_618,In_411);
nor U2967 (N_2967,In_1417,In_587);
and U2968 (N_2968,In_844,In_1209);
nand U2969 (N_2969,In_711,In_350);
and U2970 (N_2970,In_186,In_1421);
nor U2971 (N_2971,In_590,In_462);
and U2972 (N_2972,In_35,In_1079);
nand U2973 (N_2973,In_1033,In_952);
nor U2974 (N_2974,In_370,In_1019);
nor U2975 (N_2975,In_876,In_1126);
xor U2976 (N_2976,In_334,In_1350);
or U2977 (N_2977,In_682,In_672);
nor U2978 (N_2978,In_370,In_805);
and U2979 (N_2979,In_197,In_38);
and U2980 (N_2980,In_775,In_509);
or U2981 (N_2981,In_552,In_1387);
nor U2982 (N_2982,In_456,In_279);
and U2983 (N_2983,In_652,In_26);
or U2984 (N_2984,In_243,In_830);
nand U2985 (N_2985,In_1115,In_957);
nand U2986 (N_2986,In_1052,In_319);
or U2987 (N_2987,In_17,In_1072);
nor U2988 (N_2988,In_954,In_959);
nor U2989 (N_2989,In_143,In_268);
nand U2990 (N_2990,In_1361,In_1435);
and U2991 (N_2991,In_849,In_565);
nor U2992 (N_2992,In_961,In_998);
nand U2993 (N_2993,In_521,In_1193);
nand U2994 (N_2994,In_283,In_815);
and U2995 (N_2995,In_487,In_515);
nand U2996 (N_2996,In_1273,In_85);
or U2997 (N_2997,In_32,In_800);
and U2998 (N_2998,In_761,In_119);
nor U2999 (N_2999,In_666,In_1001);
or U3000 (N_3000,N_2899,N_2215);
nor U3001 (N_3001,N_1252,N_2465);
or U3002 (N_3002,N_2532,N_729);
and U3003 (N_3003,N_2754,N_1613);
nand U3004 (N_3004,N_1786,N_2699);
nand U3005 (N_3005,N_1530,N_2413);
or U3006 (N_3006,N_2974,N_9);
or U3007 (N_3007,N_2915,N_267);
xnor U3008 (N_3008,N_689,N_2193);
and U3009 (N_3009,N_2133,N_2401);
and U3010 (N_3010,N_2481,N_286);
nand U3011 (N_3011,N_2955,N_278);
or U3012 (N_3012,N_2728,N_858);
nand U3013 (N_3013,N_1555,N_698);
nor U3014 (N_3014,N_216,N_585);
or U3015 (N_3015,N_1924,N_438);
nor U3016 (N_3016,N_46,N_1358);
nand U3017 (N_3017,N_2039,N_1643);
nand U3018 (N_3018,N_1738,N_2781);
or U3019 (N_3019,N_2716,N_1879);
or U3020 (N_3020,N_1291,N_1344);
nor U3021 (N_3021,N_2403,N_621);
and U3022 (N_3022,N_569,N_2870);
or U3023 (N_3023,N_2521,N_1662);
or U3024 (N_3024,N_1255,N_1963);
or U3025 (N_3025,N_2795,N_2420);
or U3026 (N_3026,N_2200,N_1365);
nor U3027 (N_3027,N_1719,N_413);
nor U3028 (N_3028,N_847,N_882);
and U3029 (N_3029,N_1465,N_2898);
nand U3030 (N_3030,N_2230,N_269);
or U3031 (N_3031,N_2054,N_2216);
nand U3032 (N_3032,N_1265,N_2660);
nor U3033 (N_3033,N_1834,N_1002);
nand U3034 (N_3034,N_576,N_2609);
nor U3035 (N_3035,N_952,N_522);
nand U3036 (N_3036,N_2782,N_684);
nor U3037 (N_3037,N_2610,N_141);
or U3038 (N_3038,N_110,N_1121);
and U3039 (N_3039,N_505,N_2464);
nor U3040 (N_3040,N_1969,N_1029);
or U3041 (N_3041,N_776,N_1847);
nand U3042 (N_3042,N_59,N_2849);
or U3043 (N_3043,N_637,N_843);
and U3044 (N_3044,N_1778,N_2510);
nand U3045 (N_3045,N_1309,N_601);
and U3046 (N_3046,N_2491,N_214);
or U3047 (N_3047,N_398,N_51);
nand U3048 (N_3048,N_149,N_818);
and U3049 (N_3049,N_1559,N_1088);
nor U3050 (N_3050,N_2613,N_701);
and U3051 (N_3051,N_2984,N_2894);
or U3052 (N_3052,N_2385,N_1871);
or U3053 (N_3053,N_1954,N_2158);
and U3054 (N_3054,N_1878,N_2636);
nand U3055 (N_3055,N_2831,N_961);
nor U3056 (N_3056,N_2561,N_932);
or U3057 (N_3057,N_2218,N_2767);
and U3058 (N_3058,N_223,N_431);
or U3059 (N_3059,N_1189,N_2095);
or U3060 (N_3060,N_1330,N_2698);
nand U3061 (N_3061,N_193,N_2633);
nor U3062 (N_3062,N_1751,N_1135);
nand U3063 (N_3063,N_1113,N_960);
nor U3064 (N_3064,N_1663,N_1855);
nor U3065 (N_3065,N_1341,N_649);
xor U3066 (N_3066,N_1773,N_1950);
and U3067 (N_3067,N_1464,N_2222);
or U3068 (N_3068,N_2724,N_1056);
nor U3069 (N_3069,N_1168,N_1369);
or U3070 (N_3070,N_2626,N_2856);
or U3071 (N_3071,N_1357,N_1524);
nor U3072 (N_3072,N_645,N_2625);
nor U3073 (N_3073,N_382,N_2003);
nand U3074 (N_3074,N_2807,N_1030);
or U3075 (N_3075,N_1631,N_2505);
and U3076 (N_3076,N_325,N_2525);
nor U3077 (N_3077,N_2713,N_2307);
nor U3078 (N_3078,N_1755,N_936);
and U3079 (N_3079,N_548,N_995);
nand U3080 (N_3080,N_1196,N_298);
xor U3081 (N_3081,N_646,N_233);
and U3082 (N_3082,N_1597,N_1074);
or U3083 (N_3083,N_923,N_2140);
nor U3084 (N_3084,N_2747,N_2760);
and U3085 (N_3085,N_2169,N_2570);
or U3086 (N_3086,N_1355,N_1517);
or U3087 (N_3087,N_2273,N_468);
nor U3088 (N_3088,N_2298,N_941);
nand U3089 (N_3089,N_2501,N_559);
nand U3090 (N_3090,N_2280,N_2493);
nand U3091 (N_3091,N_1940,N_83);
and U3092 (N_3092,N_675,N_2500);
nor U3093 (N_3093,N_1491,N_368);
or U3094 (N_3094,N_1458,N_2542);
or U3095 (N_3095,N_2381,N_2722);
and U3096 (N_3096,N_887,N_308);
nor U3097 (N_3097,N_1959,N_1096);
and U3098 (N_3098,N_2995,N_2682);
or U3099 (N_3099,N_1649,N_2239);
or U3100 (N_3100,N_2847,N_1833);
nand U3101 (N_3101,N_2209,N_2400);
nand U3102 (N_3102,N_1201,N_2396);
nand U3103 (N_3103,N_1152,N_1138);
and U3104 (N_3104,N_929,N_2467);
nor U3105 (N_3105,N_629,N_801);
and U3106 (N_3106,N_1095,N_29);
or U3107 (N_3107,N_2873,N_1531);
or U3108 (N_3108,N_1478,N_1482);
nor U3109 (N_3109,N_1282,N_964);
nand U3110 (N_3110,N_360,N_2537);
nor U3111 (N_3111,N_1498,N_955);
or U3112 (N_3112,N_1655,N_432);
or U3113 (N_3113,N_547,N_2008);
nor U3114 (N_3114,N_1393,N_1703);
nor U3115 (N_3115,N_1173,N_2877);
or U3116 (N_3116,N_1714,N_156);
nand U3117 (N_3117,N_1034,N_473);
nand U3118 (N_3118,N_2811,N_1329);
and U3119 (N_3119,N_121,N_2349);
nor U3120 (N_3120,N_213,N_1274);
nand U3121 (N_3121,N_685,N_2253);
nor U3122 (N_3122,N_909,N_1716);
or U3123 (N_3123,N_1547,N_997);
and U3124 (N_3124,N_1296,N_951);
nor U3125 (N_3125,N_1301,N_2740);
and U3126 (N_3126,N_2549,N_1383);
nor U3127 (N_3127,N_1035,N_1960);
nand U3128 (N_3128,N_310,N_1251);
nor U3129 (N_3129,N_669,N_1585);
nand U3130 (N_3130,N_421,N_1466);
xnor U3131 (N_3131,N_1090,N_1133);
nor U3132 (N_3132,N_2842,N_915);
nor U3133 (N_3133,N_2937,N_2502);
and U3134 (N_3134,N_151,N_552);
nor U3135 (N_3135,N_2473,N_2659);
nor U3136 (N_3136,N_2271,N_2146);
and U3137 (N_3137,N_1368,N_2572);
or U3138 (N_3138,N_2233,N_2875);
nand U3139 (N_3139,N_2829,N_2766);
or U3140 (N_3140,N_2380,N_654);
nand U3141 (N_3141,N_2520,N_116);
nor U3142 (N_3142,N_289,N_190);
nor U3143 (N_3143,N_1302,N_900);
nand U3144 (N_3144,N_178,N_519);
nor U3145 (N_3145,N_856,N_195);
nand U3146 (N_3146,N_1541,N_926);
and U3147 (N_3147,N_219,N_677);
and U3148 (N_3148,N_1939,N_39);
nor U3149 (N_3149,N_2110,N_1205);
or U3150 (N_3150,N_2757,N_718);
nor U3151 (N_3151,N_876,N_2661);
nand U3152 (N_3152,N_2151,N_534);
nand U3153 (N_3153,N_2445,N_703);
xor U3154 (N_3154,N_469,N_1584);
nand U3155 (N_3155,N_1809,N_363);
or U3156 (N_3156,N_2,N_1499);
and U3157 (N_3157,N_1180,N_1408);
and U3158 (N_3158,N_2573,N_2076);
and U3159 (N_3159,N_697,N_1787);
nand U3160 (N_3160,N_2452,N_914);
nor U3161 (N_3161,N_1340,N_2485);
nand U3162 (N_3162,N_1492,N_1212);
or U3163 (N_3163,N_1112,N_2608);
nor U3164 (N_3164,N_1525,N_1403);
and U3165 (N_3165,N_1214,N_817);
and U3166 (N_3166,N_1399,N_1474);
nor U3167 (N_3167,N_1012,N_2615);
xnor U3168 (N_3168,N_2908,N_1798);
or U3169 (N_3169,N_667,N_772);
and U3170 (N_3170,N_1394,N_2334);
nor U3171 (N_3171,N_2021,N_1725);
and U3172 (N_3172,N_1389,N_614);
nor U3173 (N_3173,N_865,N_2592);
or U3174 (N_3174,N_1688,N_472);
nand U3175 (N_3175,N_1713,N_1268);
or U3176 (N_3176,N_2322,N_1682);
nor U3177 (N_3177,N_600,N_523);
xor U3178 (N_3178,N_165,N_55);
nor U3179 (N_3179,N_1974,N_1011);
and U3180 (N_3180,N_2045,N_303);
nor U3181 (N_3181,N_1164,N_92);
and U3182 (N_3182,N_68,N_1608);
and U3183 (N_3183,N_2614,N_1501);
nand U3184 (N_3184,N_602,N_1380);
nand U3185 (N_3185,N_890,N_2840);
nor U3186 (N_3186,N_1285,N_1417);
nor U3187 (N_3187,N_2835,N_2587);
nor U3188 (N_3188,N_2419,N_934);
and U3189 (N_3189,N_924,N_1920);
nand U3190 (N_3190,N_1768,N_925);
nand U3191 (N_3191,N_2191,N_895);
xor U3192 (N_3192,N_334,N_2341);
or U3193 (N_3193,N_482,N_2064);
or U3194 (N_3194,N_112,N_2606);
and U3195 (N_3195,N_1105,N_246);
nand U3196 (N_3196,N_768,N_2927);
or U3197 (N_3197,N_562,N_1653);
nand U3198 (N_3198,N_1862,N_2964);
or U3199 (N_3199,N_2836,N_1668);
and U3200 (N_3200,N_2611,N_2001);
or U3201 (N_3201,N_625,N_385);
or U3202 (N_3202,N_2292,N_810);
nand U3203 (N_3203,N_2707,N_2077);
or U3204 (N_3204,N_2965,N_2925);
or U3205 (N_3205,N_1992,N_1971);
nor U3206 (N_3206,N_226,N_1);
nand U3207 (N_3207,N_465,N_518);
and U3208 (N_3208,N_340,N_2142);
nor U3209 (N_3209,N_1518,N_1216);
nor U3210 (N_3210,N_588,N_2818);
or U3211 (N_3211,N_1005,N_2793);
nor U3212 (N_3212,N_2529,N_2255);
or U3213 (N_3213,N_1596,N_477);
nand U3214 (N_3214,N_714,N_168);
or U3215 (N_3215,N_2284,N_1063);
and U3216 (N_3216,N_2408,N_24);
xnor U3217 (N_3217,N_330,N_2675);
nand U3218 (N_3218,N_2571,N_2565);
and U3219 (N_3219,N_2617,N_447);
or U3220 (N_3220,N_2778,N_2123);
and U3221 (N_3221,N_1147,N_1219);
or U3222 (N_3222,N_832,N_1400);
and U3223 (N_3223,N_2941,N_1004);
nor U3224 (N_3224,N_1705,N_1313);
or U3225 (N_3225,N_1804,N_470);
or U3226 (N_3226,N_446,N_1933);
and U3227 (N_3227,N_492,N_1545);
and U3228 (N_3228,N_1733,N_1260);
and U3229 (N_3229,N_2906,N_2524);
nor U3230 (N_3230,N_1982,N_2460);
or U3231 (N_3231,N_795,N_917);
or U3232 (N_3232,N_2796,N_542);
nand U3233 (N_3233,N_1117,N_2632);
and U3234 (N_3234,N_2725,N_2701);
nor U3235 (N_3235,N_2597,N_2415);
nand U3236 (N_3236,N_130,N_533);
and U3237 (N_3237,N_619,N_555);
nand U3238 (N_3238,N_1103,N_782);
and U3239 (N_3239,N_1304,N_2933);
nor U3240 (N_3240,N_1576,N_1642);
nor U3241 (N_3241,N_2801,N_2189);
or U3242 (N_3242,N_1163,N_74);
nand U3243 (N_3243,N_2848,N_5);
or U3244 (N_3244,N_1925,N_963);
nor U3245 (N_3245,N_560,N_1727);
xnor U3246 (N_3246,N_1476,N_2240);
nand U3247 (N_3247,N_1704,N_2243);
or U3248 (N_3248,N_297,N_1896);
nand U3249 (N_3249,N_1336,N_1058);
xor U3250 (N_3250,N_574,N_814);
or U3251 (N_3251,N_665,N_1259);
nand U3252 (N_3252,N_991,N_475);
and U3253 (N_3253,N_1209,N_2961);
and U3254 (N_3254,N_1810,N_510);
and U3255 (N_3255,N_578,N_2872);
or U3256 (N_3256,N_2433,N_1072);
or U3257 (N_3257,N_1505,N_1983);
or U3258 (N_3258,N_692,N_607);
or U3259 (N_3259,N_2451,N_1297);
or U3260 (N_3260,N_2844,N_2731);
nand U3261 (N_3261,N_1527,N_2179);
nor U3262 (N_3262,N_2892,N_304);
and U3263 (N_3263,N_2543,N_1210);
and U3264 (N_3264,N_973,N_2553);
nor U3265 (N_3265,N_2210,N_1900);
and U3266 (N_3266,N_1588,N_2616);
xor U3267 (N_3267,N_2981,N_2670);
or U3268 (N_3268,N_892,N_2950);
nor U3269 (N_3269,N_1014,N_509);
and U3270 (N_3270,N_2862,N_906);
nor U3271 (N_3271,N_1069,N_1469);
or U3272 (N_3272,N_1027,N_2893);
nand U3273 (N_3273,N_2851,N_1680);
or U3274 (N_3274,N_16,N_2674);
nor U3275 (N_3275,N_2839,N_2258);
and U3276 (N_3276,N_2953,N_573);
nand U3277 (N_3277,N_1125,N_2669);
and U3278 (N_3278,N_383,N_1702);
and U3279 (N_3279,N_824,N_1911);
nand U3280 (N_3280,N_653,N_439);
and U3281 (N_3281,N_1529,N_2172);
nor U3282 (N_3282,N_1729,N_526);
and U3283 (N_3283,N_1182,N_2037);
nand U3284 (N_3284,N_2895,N_1762);
and U3285 (N_3285,N_828,N_612);
nor U3286 (N_3286,N_52,N_931);
nand U3287 (N_3287,N_2283,N_719);
or U3288 (N_3288,N_1534,N_616);
nand U3289 (N_3289,N_448,N_2512);
or U3290 (N_3290,N_1731,N_1685);
or U3291 (N_3291,N_631,N_496);
and U3292 (N_3292,N_830,N_2093);
nor U3293 (N_3293,N_579,N_638);
nand U3294 (N_3294,N_157,N_1289);
or U3295 (N_3295,N_798,N_1003);
and U3296 (N_3296,N_2990,N_2861);
nor U3297 (N_3297,N_1784,N_584);
nand U3298 (N_3298,N_927,N_2300);
nand U3299 (N_3299,N_132,N_1066);
or U3300 (N_3300,N_90,N_476);
and U3301 (N_3301,N_293,N_2013);
and U3302 (N_3302,N_591,N_1829);
nor U3303 (N_3303,N_1913,N_2921);
nand U3304 (N_3304,N_2639,N_1689);
nor U3305 (N_3305,N_1908,N_1536);
or U3306 (N_3306,N_537,N_2788);
nor U3307 (N_3307,N_2579,N_328);
and U3308 (N_3308,N_517,N_2676);
or U3309 (N_3309,N_1258,N_752);
nand U3310 (N_3310,N_2916,N_2315);
and U3311 (N_3311,N_49,N_133);
or U3312 (N_3312,N_1444,N_152);
nor U3313 (N_3313,N_2827,N_1735);
and U3314 (N_3314,N_1232,N_2643);
nand U3315 (N_3315,N_1697,N_1162);
nand U3316 (N_3316,N_1732,N_1238);
nand U3317 (N_3317,N_12,N_1347);
or U3318 (N_3318,N_1835,N_1799);
nor U3319 (N_3319,N_1230,N_1471);
nand U3320 (N_3320,N_984,N_145);
nor U3321 (N_3321,N_2320,N_811);
or U3322 (N_3322,N_2332,N_2254);
nand U3323 (N_3323,N_497,N_82);
or U3324 (N_3324,N_2448,N_1495);
nor U3325 (N_3325,N_1522,N_2453);
and U3326 (N_3326,N_153,N_2120);
or U3327 (N_3327,N_2407,N_1327);
nor U3328 (N_3328,N_1686,N_1695);
and U3329 (N_3329,N_2414,N_2227);
or U3330 (N_3330,N_1607,N_1549);
nor U3331 (N_3331,N_679,N_2028);
or U3332 (N_3332,N_2141,N_2548);
and U3333 (N_3333,N_1017,N_1594);
nor U3334 (N_3334,N_321,N_1627);
nand U3335 (N_3335,N_1049,N_1437);
and U3336 (N_3336,N_2441,N_415);
nor U3337 (N_3337,N_2780,N_388);
nand U3338 (N_3338,N_2582,N_243);
or U3339 (N_3339,N_1455,N_1262);
nand U3340 (N_3340,N_414,N_580);
nand U3341 (N_3341,N_624,N_1317);
nand U3342 (N_3342,N_660,N_2519);
or U3343 (N_3343,N_484,N_2858);
nor U3344 (N_3344,N_1544,N_524);
or U3345 (N_3345,N_1637,N_2486);
nand U3346 (N_3346,N_2683,N_1057);
and U3347 (N_3347,N_2034,N_2869);
or U3348 (N_3348,N_2577,N_486);
nand U3349 (N_3349,N_2359,N_381);
nand U3350 (N_3350,N_1061,N_1235);
or U3351 (N_3351,N_1757,N_613);
nor U3352 (N_3352,N_324,N_1178);
and U3353 (N_3353,N_140,N_77);
nand U3354 (N_3354,N_983,N_2952);
or U3355 (N_3355,N_1574,N_866);
nand U3356 (N_3356,N_459,N_418);
or U3357 (N_3357,N_2347,N_1957);
and U3358 (N_3358,N_2291,N_201);
and U3359 (N_3359,N_1428,N_1429);
and U3360 (N_3360,N_1550,N_910);
or U3361 (N_3361,N_261,N_2302);
nand U3362 (N_3362,N_2361,N_829);
or U3363 (N_3363,N_14,N_480);
and U3364 (N_3364,N_1987,N_2574);
or U3365 (N_3365,N_2823,N_1746);
nand U3366 (N_3366,N_1789,N_2352);
and U3367 (N_3367,N_1537,N_1333);
nand U3368 (N_3368,N_2337,N_2066);
or U3369 (N_3369,N_1569,N_1965);
nand U3370 (N_3370,N_2035,N_1816);
or U3371 (N_3371,N_2459,N_192);
nor U3372 (N_3372,N_1831,N_430);
and U3373 (N_3373,N_336,N_831);
and U3374 (N_3374,N_1456,N_2867);
and U3375 (N_3375,N_2695,N_912);
and U3376 (N_3376,N_626,N_1723);
or U3377 (N_3377,N_1823,N_295);
nand U3378 (N_3378,N_458,N_790);
and U3379 (N_3379,N_1488,N_1586);
and U3380 (N_3380,N_1460,N_1032);
or U3381 (N_3381,N_245,N_1221);
or U3382 (N_3382,N_1277,N_194);
nand U3383 (N_3383,N_2272,N_1877);
nand U3384 (N_3384,N_331,N_207);
or U3385 (N_3385,N_595,N_2876);
xor U3386 (N_3386,N_1053,N_2363);
or U3387 (N_3387,N_179,N_656);
and U3388 (N_3388,N_173,N_2723);
nand U3389 (N_3389,N_713,N_809);
nor U3390 (N_3390,N_1606,N_1308);
and U3391 (N_3391,N_1423,N_1207);
or U3392 (N_3392,N_28,N_690);
or U3393 (N_3393,N_1361,N_1667);
and U3394 (N_3394,N_350,N_1146);
and U3395 (N_3395,N_1967,N_1846);
and U3396 (N_3396,N_2299,N_1183);
nor U3397 (N_3397,N_2619,N_867);
nor U3398 (N_3398,N_707,N_1320);
nor U3399 (N_3399,N_2388,N_1116);
nor U3400 (N_3400,N_2604,N_1899);
and U3401 (N_3401,N_764,N_372);
and U3402 (N_3402,N_2094,N_1579);
and U3403 (N_3403,N_1276,N_2022);
or U3404 (N_3404,N_2988,N_322);
nor U3405 (N_3405,N_1354,N_124);
and U3406 (N_3406,N_546,N_1392);
nand U3407 (N_3407,N_115,N_1487);
nand U3408 (N_3408,N_2662,N_2742);
or U3409 (N_3409,N_23,N_2461);
nand U3410 (N_3410,N_873,N_1452);
nor U3411 (N_3411,N_1951,N_1721);
nor U3412 (N_3412,N_2833,N_2999);
nor U3413 (N_3413,N_1191,N_2103);
nand U3414 (N_3414,N_908,N_2009);
nor U3415 (N_3415,N_1629,N_109);
nand U3416 (N_3416,N_2353,N_1203);
or U3417 (N_3417,N_1507,N_1263);
nor U3418 (N_3418,N_1872,N_700);
and U3419 (N_3419,N_2161,N_1381);
nor U3420 (N_3420,N_2346,N_375);
nand U3421 (N_3421,N_2319,N_2497);
or U3422 (N_3422,N_1577,N_771);
and U3423 (N_3423,N_177,N_2350);
nor U3424 (N_3424,N_2329,N_203);
and U3425 (N_3425,N_2148,N_365);
and U3426 (N_3426,N_1071,N_928);
and U3427 (N_3427,N_2328,N_1440);
and U3428 (N_3428,N_1331,N_2260);
or U3429 (N_3429,N_225,N_2458);
or U3430 (N_3430,N_2081,N_174);
and U3431 (N_3431,N_797,N_1084);
nand U3432 (N_3432,N_4,N_864);
or U3433 (N_3433,N_235,N_403);
or U3434 (N_3434,N_2068,N_253);
and U3435 (N_3435,N_191,N_2427);
or U3436 (N_3436,N_1657,N_1165);
nand U3437 (N_3437,N_1827,N_292);
or U3438 (N_3438,N_1039,N_2507);
nand U3439 (N_3439,N_1472,N_66);
nand U3440 (N_3440,N_2362,N_392);
or U3441 (N_3441,N_2678,N_1848);
and U3442 (N_3442,N_1445,N_2217);
nor U3443 (N_3443,N_1759,N_1480);
or U3444 (N_3444,N_2905,N_1919);
nand U3445 (N_3445,N_1169,N_2228);
xor U3446 (N_3446,N_785,N_38);
nor U3447 (N_3447,N_2880,N_2390);
and U3448 (N_3448,N_1083,N_1947);
and U3449 (N_3449,N_1700,N_2330);
nor U3450 (N_3450,N_2603,N_1562);
nor U3451 (N_3451,N_581,N_182);
or U3452 (N_3452,N_1188,N_2826);
nand U3453 (N_3453,N_933,N_1136);
nand U3454 (N_3454,N_774,N_56);
nor U3455 (N_3455,N_256,N_2884);
nor U3456 (N_3456,N_640,N_2627);
nor U3457 (N_3457,N_2303,N_332);
and U3458 (N_3458,N_1928,N_1192);
or U3459 (N_3459,N_131,N_2371);
xnor U3460 (N_3460,N_957,N_661);
and U3461 (N_3461,N_979,N_69);
nand U3462 (N_3462,N_1640,N_96);
or U3463 (N_3463,N_311,N_842);
and U3464 (N_3464,N_301,N_2069);
or U3465 (N_3465,N_443,N_1325);
and U3466 (N_3466,N_312,N_2555);
or U3467 (N_3467,N_632,N_879);
nand U3468 (N_3468,N_67,N_85);
nand U3469 (N_3469,N_1931,N_590);
or U3470 (N_3470,N_2599,N_888);
nand U3471 (N_3471,N_1374,N_2855);
nand U3472 (N_3472,N_978,N_2259);
or U3473 (N_3473,N_2559,N_2986);
nand U3474 (N_3474,N_760,N_2137);
nor U3475 (N_3475,N_2846,N_1194);
nand U3476 (N_3476,N_239,N_853);
nand U3477 (N_3477,N_1793,N_1684);
nor U3478 (N_3478,N_1825,N_820);
nand U3479 (N_3479,N_2944,N_618);
nand U3480 (N_3480,N_1548,N_2078);
nand U3481 (N_3481,N_299,N_2373);
or U3482 (N_3482,N_2691,N_136);
and U3483 (N_3483,N_1275,N_1064);
nor U3484 (N_3484,N_2607,N_2992);
and U3485 (N_3485,N_323,N_2528);
nand U3486 (N_3486,N_1849,N_2192);
and U3487 (N_3487,N_2541,N_259);
nand U3488 (N_3488,N_990,N_544);
and U3489 (N_3489,N_2399,N_1587);
and U3490 (N_3490,N_346,N_949);
or U3491 (N_3491,N_1792,N_268);
nand U3492 (N_3492,N_2809,N_2374);
or U3493 (N_3493,N_1861,N_1788);
nand U3494 (N_3494,N_706,N_2263);
nand U3495 (N_3495,N_2206,N_2083);
nor U3496 (N_3496,N_582,N_784);
or U3497 (N_3497,N_2256,N_623);
nor U3498 (N_3498,N_2552,N_103);
and U3499 (N_3499,N_503,N_366);
and U3500 (N_3500,N_733,N_1625);
nor U3501 (N_3501,N_977,N_647);
or U3502 (N_3502,N_2679,N_1353);
nand U3503 (N_3503,N_1010,N_2494);
and U3504 (N_3504,N_274,N_833);
and U3505 (N_3505,N_462,N_1591);
or U3506 (N_3506,N_652,N_1915);
nand U3507 (N_3507,N_2018,N_1253);
and U3508 (N_3508,N_1973,N_1382);
nor U3509 (N_3509,N_2339,N_343);
nand U3510 (N_3510,N_1876,N_2602);
nor U3511 (N_3511,N_464,N_1828);
nand U3512 (N_3512,N_1051,N_2287);
or U3513 (N_3513,N_281,N_2717);
nand U3514 (N_3514,N_449,N_954);
or U3515 (N_3515,N_181,N_1434);
or U3516 (N_3516,N_1853,N_1019);
nand U3517 (N_3517,N_64,N_2113);
nor U3518 (N_3518,N_2170,N_1015);
nand U3519 (N_3519,N_702,N_2816);
nor U3520 (N_3520,N_994,N_1432);
or U3521 (N_3521,N_736,N_2276);
and U3522 (N_3522,N_2049,N_15);
or U3523 (N_3523,N_1181,N_2308);
nand U3524 (N_3524,N_2153,N_767);
nor U3525 (N_3525,N_1826,N_694);
and U3526 (N_3526,N_1479,N_2000);
or U3527 (N_3527,N_37,N_1946);
or U3528 (N_3528,N_884,N_127);
or U3529 (N_3529,N_1195,N_2741);
or U3530 (N_3530,N_2180,N_395);
nor U3531 (N_3531,N_881,N_1580);
nor U3532 (N_3532,N_2097,N_854);
nor U3533 (N_3533,N_1171,N_778);
or U3534 (N_3534,N_1237,N_2903);
nor U3535 (N_3535,N_2174,N_1601);
and U3536 (N_3536,N_1989,N_948);
and U3537 (N_3537,N_514,N_2687);
nand U3538 (N_3538,N_184,N_2434);
or U3539 (N_3539,N_1504,N_520);
nand U3540 (N_3540,N_2554,N_525);
nand U3541 (N_3541,N_2031,N_516);
or U3542 (N_3542,N_2483,N_370);
or U3543 (N_3543,N_568,N_1286);
nor U3544 (N_3544,N_2024,N_1822);
or U3545 (N_3545,N_1366,N_1885);
or U3546 (N_3546,N_780,N_2462);
and U3547 (N_3547,N_2994,N_2539);
nor U3548 (N_3548,N_1127,N_2223);
nand U3549 (N_3549,N_1615,N_359);
nor U3550 (N_3550,N_1351,N_586);
or U3551 (N_3551,N_980,N_1139);
nand U3552 (N_3552,N_1288,N_1620);
or U3553 (N_3553,N_2857,N_376);
and U3554 (N_3554,N_1018,N_2504);
nand U3555 (N_3555,N_6,N_2580);
or U3556 (N_3556,N_2423,N_2730);
and U3557 (N_3557,N_1687,N_2313);
nand U3558 (N_3558,N_1332,N_401);
nand U3559 (N_3559,N_1986,N_1770);
nor U3560 (N_3560,N_2694,N_2978);
or U3561 (N_3561,N_35,N_2377);
or U3562 (N_3562,N_845,N_455);
and U3563 (N_3563,N_1502,N_803);
nand U3564 (N_3564,N_1690,N_187);
xor U3565 (N_3565,N_2666,N_1709);
nor U3566 (N_3566,N_1054,N_2985);
nor U3567 (N_3567,N_185,N_11);
or U3568 (N_3568,N_2389,N_369);
nor U3569 (N_3569,N_2649,N_2321);
nor U3570 (N_3570,N_558,N_1820);
nor U3571 (N_3571,N_251,N_1228);
nand U3572 (N_3572,N_1953,N_1777);
nand U3573 (N_3573,N_1602,N_1184);
and U3574 (N_3574,N_604,N_1451);
and U3575 (N_3575,N_1172,N_862);
and U3576 (N_3576,N_1503,N_1363);
and U3577 (N_3577,N_339,N_1859);
and U3578 (N_3578,N_1886,N_2394);
nand U3579 (N_3579,N_1411,N_1486);
and U3580 (N_3580,N_2111,N_2325);
nand U3581 (N_3581,N_2144,N_2438);
nor U3582 (N_3582,N_2136,N_2027);
nor U3583 (N_3583,N_2108,N_88);
and U3584 (N_3584,N_450,N_2265);
and U3585 (N_3585,N_686,N_2783);
or U3586 (N_3586,N_1747,N_1819);
and U3587 (N_3587,N_2853,N_2221);
nand U3588 (N_3588,N_1186,N_2972);
and U3589 (N_3589,N_1665,N_2982);
xor U3590 (N_3590,N_839,N_2063);
nand U3591 (N_3591,N_1568,N_2358);
or U3592 (N_3592,N_389,N_2550);
or U3593 (N_3593,N_2168,N_1159);
nand U3594 (N_3594,N_95,N_2475);
nor U3595 (N_3595,N_2772,N_2923);
nand U3596 (N_3596,N_710,N_2951);
or U3597 (N_3597,N_1654,N_1050);
and U3598 (N_3598,N_1851,N_2454);
or U3599 (N_3599,N_2157,N_258);
or U3600 (N_3600,N_1857,N_1044);
nor U3601 (N_3601,N_746,N_2787);
and U3602 (N_3602,N_1991,N_1753);
nor U3603 (N_3603,N_2693,N_1160);
nor U3604 (N_3604,N_2245,N_2503);
and U3605 (N_3605,N_1632,N_1385);
nor U3606 (N_3606,N_2644,N_1672);
xnor U3607 (N_3607,N_1006,N_488);
nand U3608 (N_3608,N_1157,N_1889);
and U3609 (N_3609,N_2564,N_2262);
nand U3610 (N_3610,N_13,N_1553);
nor U3611 (N_3611,N_2530,N_358);
nor U3612 (N_3612,N_423,N_1538);
and U3613 (N_3613,N_2029,N_2264);
or U3614 (N_3614,N_2152,N_1890);
nand U3615 (N_3615,N_408,N_566);
or U3616 (N_3616,N_2712,N_512);
nor U3617 (N_3617,N_2004,N_2959);
nor U3618 (N_3618,N_2948,N_699);
nand U3619 (N_3619,N_1048,N_1204);
nand U3620 (N_3620,N_1717,N_1906);
and U3621 (N_3621,N_2885,N_1154);
nand U3622 (N_3622,N_155,N_2250);
or U3623 (N_3623,N_483,N_129);
nand U3624 (N_3624,N_2940,N_2680);
or U3625 (N_3625,N_1844,N_1808);
or U3626 (N_3626,N_32,N_2416);
and U3627 (N_3627,N_1185,N_2297);
or U3628 (N_3628,N_1158,N_2444);
nor U3629 (N_3629,N_822,N_1715);
nor U3630 (N_3630,N_1242,N_2968);
nor U3631 (N_3631,N_2977,N_390);
and U3632 (N_3632,N_1223,N_844);
nand U3633 (N_3633,N_2417,N_1055);
and U3634 (N_3634,N_1681,N_2718);
or U3635 (N_3635,N_756,N_1148);
or U3636 (N_3636,N_2336,N_169);
nand U3637 (N_3637,N_2719,N_904);
nor U3638 (N_3638,N_2088,N_2623);
or U3639 (N_3639,N_2122,N_2584);
nand U3640 (N_3640,N_605,N_1079);
nor U3641 (N_3641,N_2771,N_2038);
and U3642 (N_3642,N_1978,N_2668);
or U3643 (N_3643,N_2652,N_2932);
nor U3644 (N_3644,N_2756,N_2883);
or U3645 (N_3645,N_1500,N_2721);
nor U3646 (N_3646,N_143,N_2211);
nor U3647 (N_3647,N_1948,N_996);
or U3648 (N_3648,N_2020,N_766);
or U3649 (N_3649,N_2509,N_1818);
nor U3650 (N_3650,N_2980,N_2134);
nor U3651 (N_3651,N_1617,N_1321);
nor U3652 (N_3652,N_709,N_2897);
nor U3653 (N_3653,N_327,N_362);
nand U3654 (N_3654,N_2411,N_1093);
xor U3655 (N_3655,N_104,N_1187);
or U3656 (N_3656,N_1076,N_2803);
nor U3657 (N_3657,N_846,N_1750);
nand U3658 (N_3658,N_353,N_775);
and U3659 (N_3659,N_456,N_2917);
nor U3660 (N_3660,N_1952,N_1416);
or U3661 (N_3661,N_1901,N_1401);
and U3662 (N_3662,N_2479,N_1342);
and U3663 (N_3663,N_1560,N_2375);
nor U3664 (N_3664,N_2477,N_2640);
nand U3665 (N_3665,N_2738,N_236);
or U3666 (N_3666,N_1880,N_139);
nand U3667 (N_3667,N_2711,N_1623);
nand U3668 (N_3668,N_1244,N_1628);
nor U3669 (N_3669,N_893,N_314);
nand U3670 (N_3670,N_2446,N_474);
nor U3671 (N_3671,N_2929,N_1047);
and U3672 (N_3672,N_664,N_1763);
nand U3673 (N_3673,N_615,N_671);
nor U3674 (N_3674,N_2594,N_804);
nand U3675 (N_3675,N_1007,N_2071);
nand U3676 (N_3676,N_1509,N_241);
nand U3677 (N_3677,N_2014,N_1927);
nand U3678 (N_3678,N_2409,N_1803);
or U3679 (N_3679,N_2966,N_589);
nor U3680 (N_3680,N_454,N_1661);
nor U3681 (N_3681,N_2969,N_874);
nand U3682 (N_3682,N_1413,N_436);
and U3683 (N_3683,N_2079,N_2702);
or U3684 (N_3684,N_796,N_87);
or U3685 (N_3685,N_608,N_1790);
nor U3686 (N_3686,N_662,N_2422);
and U3687 (N_3687,N_2852,N_2736);
and U3688 (N_3688,N_1882,N_2251);
nor U3689 (N_3689,N_683,N_969);
or U3690 (N_3690,N_171,N_161);
and U3691 (N_3691,N_765,N_2798);
and U3692 (N_3692,N_2815,N_1106);
or U3693 (N_3693,N_1736,N_164);
nor U3694 (N_3694,N_2405,N_1272);
or U3695 (N_3695,N_2171,N_391);
nand U3696 (N_3696,N_2257,N_1592);
or U3697 (N_3697,N_341,N_1863);
nand U3698 (N_3698,N_2293,N_2187);
nand U3699 (N_3699,N_271,N_463);
or U3700 (N_3700,N_229,N_2007);
nand U3701 (N_3701,N_2650,N_1150);
nand U3702 (N_3702,N_10,N_2850);
and U3703 (N_3703,N_148,N_1122);
and U3704 (N_3704,N_1371,N_794);
nand U3705 (N_3705,N_2517,N_2457);
or U3706 (N_3706,N_1130,N_583);
nand U3707 (N_3707,N_531,N_1120);
or U3708 (N_3708,N_515,N_557);
and U3709 (N_3709,N_1250,N_1352);
or U3710 (N_3710,N_922,N_1712);
or U3711 (N_3711,N_606,N_1641);
and U3712 (N_3712,N_276,N_1459);
and U3713 (N_3713,N_435,N_1198);
xnor U3714 (N_3714,N_2436,N_918);
nor U3715 (N_3715,N_1001,N_479);
nand U3716 (N_3716,N_1026,N_396);
nand U3717 (N_3717,N_73,N_255);
nand U3718 (N_3718,N_761,N_564);
or U3719 (N_3719,N_1761,N_99);
and U3720 (N_3720,N_2547,N_2551);
or U3721 (N_3721,N_1766,N_1980);
nand U3722 (N_3722,N_2882,N_861);
and U3723 (N_3723,N_108,N_1619);
or U3724 (N_3724,N_642,N_2214);
nand U3725 (N_3725,N_2774,N_1025);
nand U3726 (N_3726,N_2891,N_1273);
nor U3727 (N_3727,N_1552,N_2514);
nor U3728 (N_3728,N_142,N_1418);
and U3729 (N_3729,N_1845,N_693);
and U3730 (N_3730,N_2620,N_1801);
or U3731 (N_3731,N_2372,N_1583);
nand U3732 (N_3732,N_1115,N_807);
or U3733 (N_3733,N_128,N_2490);
nor U3734 (N_3734,N_1081,N_2729);
and U3735 (N_3735,N_2804,N_357);
nor U3736 (N_3736,N_1231,N_114);
nor U3737 (N_3737,N_1837,N_1350);
nand U3738 (N_3738,N_2762,N_2348);
nor U3739 (N_3739,N_33,N_1461);
nor U3740 (N_3740,N_2946,N_1867);
and U3741 (N_3741,N_2005,N_2048);
and U3742 (N_3742,N_1838,N_2181);
nand U3743 (N_3743,N_1639,N_1449);
nor U3744 (N_3744,N_2967,N_2828);
nand U3745 (N_3745,N_2425,N_1683);
nor U3746 (N_3746,N_1243,N_593);
or U3747 (N_3747,N_97,N_2499);
nor U3748 (N_3748,N_1817,N_1995);
and U3749 (N_3749,N_2369,N_812);
and U3750 (N_3750,N_735,N_950);
nand U3751 (N_3751,N_1912,N_208);
nand U3752 (N_3752,N_309,N_1956);
nand U3753 (N_3753,N_1193,N_290);
or U3754 (N_3754,N_138,N_2357);
nor U3755 (N_3755,N_1021,N_2053);
and U3756 (N_3756,N_1441,N_1065);
or U3757 (N_3757,N_749,N_1170);
or U3758 (N_3758,N_1144,N_1294);
nand U3759 (N_3759,N_1305,N_2073);
or U3760 (N_3760,N_919,N_1131);
nor U3761 (N_3761,N_1557,N_970);
xnor U3762 (N_3762,N_1856,N_1454);
or U3763 (N_3763,N_1324,N_1779);
and U3764 (N_3764,N_2904,N_1475);
and U3765 (N_3765,N_2928,N_848);
and U3766 (N_3766,N_1390,N_1582);
and U3767 (N_3767,N_1462,N_441);
nand U3768 (N_3768,N_672,N_2125);
nand U3769 (N_3769,N_1865,N_726);
and U3770 (N_3770,N_2591,N_2051);
nor U3771 (N_3771,N_1671,N_953);
or U3772 (N_3772,N_1367,N_2086);
or U3773 (N_3773,N_2016,N_1624);
xnor U3774 (N_3774,N_1666,N_1299);
nor U3775 (N_3775,N_2041,N_2645);
and U3776 (N_3776,N_275,N_1558);
and U3777 (N_3777,N_1780,N_787);
or U3778 (N_3778,N_166,N_2791);
nand U3779 (N_3779,N_1614,N_1318);
or U3780 (N_3780,N_611,N_708);
and U3781 (N_3781,N_1903,N_222);
and U3782 (N_3782,N_875,N_294);
or U3783 (N_3783,N_2578,N_405);
nand U3784 (N_3784,N_2275,N_532);
nor U3785 (N_3785,N_1346,N_942);
nand U3786 (N_3786,N_2802,N_2468);
nand U3787 (N_3787,N_2601,N_1156);
nor U3788 (N_3788,N_1694,N_2700);
and U3789 (N_3789,N_1123,N_2241);
and U3790 (N_3790,N_891,N_789);
or U3791 (N_3791,N_2149,N_1881);
and U3792 (N_3792,N_1377,N_2688);
and U3793 (N_3793,N_2323,N_2991);
nor U3794 (N_3794,N_1395,N_1270);
and U3795 (N_3795,N_1921,N_424);
nor U3796 (N_3796,N_305,N_1009);
xor U3797 (N_3797,N_1636,N_499);
or U3798 (N_3798,N_1370,N_1384);
and U3799 (N_3799,N_404,N_2919);
and U3800 (N_3800,N_1758,N_2720);
or U3801 (N_3801,N_1740,N_221);
and U3802 (N_3802,N_2685,N_2019);
and U3803 (N_3803,N_1630,N_1744);
or U3804 (N_3804,N_2677,N_2044);
nor U3805 (N_3805,N_3,N_1234);
or U3806 (N_3806,N_2182,N_1679);
or U3807 (N_3807,N_1279,N_2768);
and U3808 (N_3808,N_2266,N_227);
xor U3809 (N_3809,N_1566,N_628);
and U3810 (N_3810,N_377,N_691);
or U3811 (N_3811,N_1651,N_1436);
nor U3812 (N_3812,N_427,N_326);
nand U3813 (N_3813,N_2267,N_1442);
and U3814 (N_3814,N_1045,N_1692);
nand U3815 (N_3815,N_407,N_1020);
nand U3816 (N_3816,N_453,N_1082);
nor U3817 (N_3817,N_999,N_2637);
nor U3818 (N_3818,N_1916,N_896);
nand U3819 (N_3819,N_1975,N_1328);
nand U3820 (N_3820,N_2817,N_808);
nor U3821 (N_3821,N_119,N_2518);
or U3822 (N_3822,N_2026,N_2672);
or U3823 (N_3823,N_1477,N_1433);
nor U3824 (N_3824,N_935,N_1022);
or U3825 (N_3825,N_2006,N_1080);
nor U3826 (N_3826,N_556,N_1388);
and U3827 (N_3827,N_2050,N_337);
or U3828 (N_3828,N_2585,N_1841);
and U3829 (N_3829,N_1658,N_1942);
and U3830 (N_3830,N_2526,N_1240);
or U3831 (N_3831,N_2040,N_412);
and U3832 (N_3832,N_2091,N_349);
or U3833 (N_3833,N_2197,N_1573);
or U3834 (N_3834,N_2080,N_306);
or U3835 (N_3835,N_1409,N_530);
and U3836 (N_3836,N_1791,N_687);
or U3837 (N_3837,N_2489,N_2655);
nor U3838 (N_3838,N_2709,N_2901);
nor U3839 (N_3839,N_2395,N_1407);
and U3840 (N_3840,N_821,N_880);
nor U3841 (N_3841,N_102,N_2631);
and U3842 (N_3842,N_1211,N_498);
and U3843 (N_3843,N_2622,N_826);
nor U3844 (N_3844,N_2646,N_2753);
nand U3845 (N_3845,N_2450,N_2665);
or U3846 (N_3846,N_800,N_1227);
nand U3847 (N_3847,N_1955,N_2987);
nor U3848 (N_3848,N_280,N_1129);
nor U3849 (N_3849,N_1463,N_163);
nor U3850 (N_3850,N_2703,N_2199);
and U3851 (N_3851,N_899,N_1128);
and U3852 (N_3852,N_1800,N_98);
nor U3853 (N_3853,N_2178,N_1241);
nand U3854 (N_3854,N_296,N_238);
nand U3855 (N_3855,N_723,N_902);
and U3856 (N_3856,N_799,N_2469);
or U3857 (N_3857,N_1806,N_2387);
or U3858 (N_3858,N_1533,N_859);
or U3859 (N_3859,N_791,N_2648);
or U3860 (N_3860,N_2428,N_1149);
nand U3861 (N_3861,N_125,N_371);
or U3862 (N_3862,N_2737,N_2112);
nand U3863 (N_3863,N_985,N_2203);
nor U3864 (N_3864,N_1783,N_2129);
nor U3865 (N_3865,N_1875,N_1378);
nor U3866 (N_3866,N_1563,N_19);
and U3867 (N_3867,N_2983,N_1646);
and U3868 (N_3868,N_2590,N_1316);
and U3869 (N_3869,N_2205,N_2588);
or U3870 (N_3870,N_2365,N_94);
nand U3871 (N_3871,N_2229,N_592);
and U3872 (N_3872,N_1737,N_2480);
or U3873 (N_3873,N_44,N_2705);
and U3874 (N_3874,N_1564,N_1008);
nand U3875 (N_3875,N_1612,N_2224);
and U3876 (N_3876,N_2492,N_2750);
nor U3877 (N_3877,N_356,N_1958);
and U3878 (N_3878,N_740,N_2268);
nand U3879 (N_3879,N_242,N_1497);
nand U3880 (N_3880,N_2343,N_1870);
nor U3881 (N_3881,N_2651,N_745);
and U3882 (N_3882,N_540,N_1600);
and U3883 (N_3883,N_1994,N_1981);
and U3884 (N_3884,N_2225,N_1599);
nand U3885 (N_3885,N_2121,N_2931);
and U3886 (N_3886,N_1239,N_461);
or U3887 (N_3887,N_2058,N_1042);
nand U3888 (N_3888,N_380,N_1795);
nand U3889 (N_3889,N_2331,N_1589);
nor U3890 (N_3890,N_2734,N_870);
or U3891 (N_3891,N_1581,N_1110);
and U3892 (N_3892,N_162,N_2085);
or U3893 (N_3893,N_2011,N_494);
xor U3894 (N_3894,N_738,N_2773);
nand U3895 (N_3895,N_2195,N_712);
or U3896 (N_3896,N_176,N_2102);
nor U3897 (N_3897,N_1373,N_1016);
or U3898 (N_3898,N_1909,N_2887);
nor U3899 (N_3899,N_1493,N_1830);
nand U3900 (N_3900,N_30,N_1676);
and U3901 (N_3901,N_2128,N_2527);
or U3902 (N_3902,N_150,N_2586);
nand U3903 (N_3903,N_428,N_2017);
nor U3904 (N_3904,N_1398,N_1167);
and U3905 (N_3905,N_731,N_1656);
or U3906 (N_3906,N_2455,N_2900);
nor U3907 (N_3907,N_444,N_2344);
or U3908 (N_3908,N_2997,N_663);
and U3909 (N_3909,N_1922,N_609);
or U3910 (N_3910,N_118,N_2746);
and U3911 (N_3911,N_2513,N_2800);
and U3912 (N_3912,N_42,N_2484);
and U3913 (N_3913,N_2131,N_1107);
and U3914 (N_3914,N_806,N_2805);
nand U3915 (N_3915,N_351,N_1375);
xor U3916 (N_3916,N_1339,N_1372);
and U3917 (N_3917,N_2775,N_2998);
and U3918 (N_3918,N_1561,N_335);
nor U3919 (N_3919,N_2278,N_333);
nor U3920 (N_3920,N_2794,N_2912);
and U3921 (N_3921,N_2871,N_2410);
nor U3922 (N_3922,N_670,N_1420);
or U3923 (N_3923,N_1938,N_2107);
and U3924 (N_3924,N_89,N_989);
nand U3925 (N_3925,N_897,N_2913);
or U3926 (N_3926,N_240,N_620);
nand U3927 (N_3927,N_2442,N_2059);
nand U3928 (N_3928,N_1073,N_2970);
or U3929 (N_3929,N_2378,N_1565);
and U3930 (N_3930,N_1767,N_1745);
nor U3931 (N_3931,N_577,N_2190);
nand U3932 (N_3932,N_958,N_1895);
nand U3933 (N_3933,N_1621,N_535);
nand U3934 (N_3934,N_777,N_400);
nor U3935 (N_3935,N_1932,N_1510);
xnor U3936 (N_3936,N_722,N_639);
or U3937 (N_3937,N_2384,N_41);
and U3938 (N_3938,N_871,N_1944);
or U3939 (N_3939,N_1515,N_1858);
and U3940 (N_3940,N_1781,N_2863);
nor U3941 (N_3941,N_2237,N_536);
nor U3942 (N_3942,N_1067,N_1315);
or U3943 (N_3943,N_282,N_2947);
or U3944 (N_3944,N_1284,N_2082);
xor U3945 (N_3945,N_2162,N_1894);
nand U3946 (N_3946,N_1868,N_2247);
and U3947 (N_3947,N_93,N_2671);
nor U3948 (N_3948,N_2084,N_2163);
nand U3949 (N_3949,N_1701,N_2010);
nor U3950 (N_3950,N_786,N_2176);
and U3951 (N_3951,N_160,N_2426);
or U3952 (N_3952,N_1166,N_575);
nor U3953 (N_3953,N_1448,N_1467);
nor U3954 (N_3954,N_2270,N_972);
nand U3955 (N_3955,N_1360,N_2938);
nor U3956 (N_3956,N_111,N_1349);
and U3957 (N_3957,N_1334,N_1650);
or U3958 (N_3958,N_2089,N_1199);
nor U3959 (N_3959,N_1739,N_113);
nor U3960 (N_3960,N_863,N_1485);
nor U3961 (N_3961,N_1893,N_1722);
or U3962 (N_3962,N_1945,N_1874);
and U3963 (N_3963,N_1698,N_597);
and U3964 (N_3964,N_857,N_204);
or U3965 (N_3965,N_855,N_1720);
and U3966 (N_3966,N_101,N_1450);
and U3967 (N_3967,N_2820,N_2326);
nor U3968 (N_3968,N_1961,N_1511);
or U3969 (N_3969,N_943,N_1752);
nand U3970 (N_3970,N_7,N_1376);
or U3971 (N_3971,N_1843,N_2656);
and U3972 (N_3972,N_1962,N_705);
nor U3973 (N_3973,N_402,N_2294);
nor U3974 (N_3974,N_2364,N_2447);
or U3975 (N_3975,N_1929,N_1618);
or U3976 (N_3976,N_1824,N_1410);
and U3977 (N_3977,N_2595,N_2508);
nand U3978 (N_3978,N_2317,N_452);
or U3979 (N_3979,N_263,N_1949);
and U3980 (N_3980,N_2515,N_1660);
or U3981 (N_3981,N_283,N_2301);
or U3982 (N_3982,N_2376,N_1114);
nand U3983 (N_3983,N_1897,N_1622);
nor U3984 (N_3984,N_1923,N_437);
nor U3985 (N_3985,N_2511,N_1314);
nor U3986 (N_3986,N_117,N_2540);
and U3987 (N_3987,N_2681,N_2789);
and U3988 (N_3988,N_501,N_2824);
nor U3989 (N_3989,N_1604,N_2733);
or U3990 (N_3990,N_1769,N_940);
nand U3991 (N_3991,N_1267,N_2269);
and U3992 (N_3992,N_1043,N_120);
nand U3993 (N_3993,N_1220,N_1869);
nand U3994 (N_3994,N_2101,N_27);
nand U3995 (N_3995,N_2575,N_2098);
nor U3996 (N_3996,N_877,N_2739);
and U3997 (N_3997,N_1280,N_1292);
and U3998 (N_3998,N_2830,N_348);
and U3999 (N_3999,N_2690,N_2440);
nand U4000 (N_4000,N_86,N_1040);
and U4001 (N_4001,N_783,N_2055);
and U4002 (N_4002,N_1696,N_2312);
nor U4003 (N_4003,N_2478,N_344);
nor U4004 (N_4004,N_183,N_755);
nor U4005 (N_4005,N_2686,N_2763);
or U4006 (N_4006,N_762,N_1206);
nand U4007 (N_4007,N_1542,N_287);
nand U4008 (N_4008,N_2911,N_1850);
and U4009 (N_4009,N_2126,N_1322);
nand U4010 (N_4010,N_976,N_1814);
or U4011 (N_4011,N_724,N_2704);
and U4012 (N_4012,N_2962,N_2360);
or U4013 (N_4013,N_1710,N_2100);
or U4014 (N_4014,N_627,N_230);
and U4015 (N_4015,N_2404,N_1293);
nand U4016 (N_4016,N_1902,N_211);
nand U4017 (N_4017,N_1771,N_758);
nor U4018 (N_4018,N_2567,N_122);
nand U4019 (N_4019,N_232,N_1405);
nand U4020 (N_4020,N_1326,N_2918);
and U4021 (N_4021,N_617,N_2368);
nor U4022 (N_4022,N_1970,N_959);
or U4023 (N_4023,N_2306,N_319);
and U4024 (N_4024,N_1261,N_1059);
and U4025 (N_4025,N_338,N_1764);
nor U4026 (N_4026,N_644,N_384);
nor U4027 (N_4027,N_2600,N_1248);
nor U4028 (N_4028,N_285,N_393);
and U4029 (N_4029,N_2506,N_2208);
and U4030 (N_4030,N_1078,N_1670);
nor U4031 (N_4031,N_2160,N_2285);
nor U4032 (N_4032,N_1590,N_2556);
or U4033 (N_4033,N_2236,N_1892);
or U4034 (N_4034,N_2155,N_2808);
or U4035 (N_4035,N_1998,N_1438);
or U4036 (N_4036,N_2759,N_2318);
and U4037 (N_4037,N_2533,N_2186);
nand U4038 (N_4038,N_146,N_1785);
xor U4039 (N_4039,N_504,N_2392);
nand U4040 (N_4040,N_175,N_1678);
nor U4041 (N_4041,N_1815,N_750);
nand U4042 (N_4042,N_2118,N_2370);
or U4043 (N_4043,N_1972,N_2822);
and U4044 (N_4044,N_2797,N_1718);
or U4045 (N_4045,N_2834,N_920);
nor U4046 (N_4046,N_1427,N_872);
nor U4047 (N_4047,N_416,N_2866);
nor U4048 (N_4048,N_2099,N_2166);
nand U4049 (N_4049,N_2673,N_1811);
nor U4050 (N_4050,N_2758,N_40);
and U4051 (N_4051,N_674,N_986);
nand U4052 (N_4052,N_2201,N_2279);
nand U4053 (N_4053,N_248,N_1312);
and U4054 (N_4054,N_2463,N_1177);
and U4055 (N_4055,N_1264,N_2327);
nor U4056 (N_4056,N_2406,N_1111);
or U4057 (N_4057,N_1634,N_47);
nor U4058 (N_4058,N_387,N_543);
nor U4059 (N_4059,N_1226,N_2838);
or U4060 (N_4060,N_1406,N_1097);
nor U4061 (N_4061,N_2926,N_2437);
nand U4062 (N_4062,N_364,N_2886);
and U4063 (N_4063,N_1421,N_2889);
or U4064 (N_4064,N_2012,N_1141);
nand U4065 (N_4065,N_2634,N_539);
nand U4066 (N_4066,N_1842,N_1610);
or U4067 (N_4067,N_1941,N_313);
nand U4068 (N_4068,N_1457,N_825);
nor U4069 (N_4069,N_206,N_657);
or U4070 (N_4070,N_91,N_747);
nor U4071 (N_4071,N_189,N_352);
nor U4072 (N_4072,N_1675,N_651);
nand U4073 (N_4073,N_2231,N_2910);
nand U4074 (N_4074,N_2316,N_254);
nor U4075 (N_4075,N_2234,N_2735);
and U4076 (N_4076,N_678,N_284);
nand U4077 (N_4077,N_1046,N_1528);
nor U4078 (N_4078,N_634,N_883);
nand U4079 (N_4079,N_1996,N_2132);
nor U4080 (N_4080,N_426,N_956);
and U4081 (N_4081,N_205,N_2583);
or U4082 (N_4082,N_2976,N_1888);
nor U4083 (N_4083,N_1760,N_1990);
or U4084 (N_4084,N_913,N_1023);
nor U4085 (N_4085,N_2443,N_2814);
xnor U4086 (N_4086,N_658,N_320);
or U4087 (N_4087,N_1068,N_1512);
nor U4088 (N_4088,N_753,N_2391);
nor U4089 (N_4089,N_273,N_397);
and U4090 (N_4090,N_840,N_2032);
or U4091 (N_4091,N_2274,N_2945);
nand U4092 (N_4092,N_2252,N_457);
and U4093 (N_4093,N_2664,N_1693);
and U4094 (N_4094,N_2367,N_471);
nand U4095 (N_4095,N_2745,N_2708);
and U4096 (N_4096,N_1283,N_2657);
or U4097 (N_4097,N_1821,N_1174);
and U4098 (N_4098,N_379,N_2498);
or U4099 (N_4099,N_975,N_751);
or U4100 (N_4100,N_666,N_105);
or U4101 (N_4101,N_968,N_272);
nand U4102 (N_4102,N_1520,N_2296);
nand U4103 (N_4103,N_759,N_65);
or U4104 (N_4104,N_1904,N_2647);
nand U4105 (N_4105,N_2092,N_367);
nand U4106 (N_4106,N_1222,N_1104);
nor U4107 (N_4107,N_2868,N_374);
xor U4108 (N_4108,N_2177,N_481);
nand U4109 (N_4109,N_841,N_2654);
or U4110 (N_4110,N_291,N_2167);
or U4111 (N_4111,N_1749,N_1236);
and U4112 (N_4112,N_123,N_1997);
or U4113 (N_4113,N_43,N_2127);
xor U4114 (N_4114,N_2070,N_2618);
nand U4115 (N_4115,N_1652,N_1387);
and U4116 (N_4116,N_2246,N_1988);
nor U4117 (N_4117,N_31,N_849);
nor U4118 (N_4118,N_2598,N_48);
nor U4119 (N_4119,N_2770,N_1807);
nand U4120 (N_4120,N_2430,N_636);
nor U4121 (N_4121,N_1099,N_1540);
nand U4122 (N_4122,N_838,N_937);
nand U4123 (N_4123,N_2924,N_2743);
or U4124 (N_4124,N_860,N_2067);
or U4125 (N_4125,N_2624,N_1935);
nand U4126 (N_4126,N_2311,N_134);
nand U4127 (N_4127,N_342,N_2355);
nor U4128 (N_4128,N_2939,N_2335);
or U4129 (N_4129,N_2562,N_2692);
and U4130 (N_4130,N_730,N_598);
or U4131 (N_4131,N_2825,N_433);
nand U4132 (N_4132,N_823,N_354);
nand U4133 (N_4133,N_355,N_988);
nand U4134 (N_4134,N_2560,N_61);
or U4135 (N_4135,N_2989,N_1179);
nor U4136 (N_4136,N_2290,N_1930);
nand U4137 (N_4137,N_885,N_2117);
nand U4138 (N_4138,N_2402,N_2638);
nand U4139 (N_4139,N_2036,N_2776);
and U4140 (N_4140,N_1140,N_553);
and U4141 (N_4141,N_2435,N_2482);
or U4142 (N_4142,N_1866,N_1839);
nor U4143 (N_4143,N_981,N_485);
or U4144 (N_4144,N_1249,N_930);
nor U4145 (N_4145,N_2145,N_2249);
nor U4146 (N_4146,N_1664,N_84);
or U4147 (N_4147,N_1483,N_987);
or U4148 (N_4148,N_1124,N_2878);
nand U4149 (N_4149,N_17,N_2202);
nor U4150 (N_4150,N_1215,N_231);
nor U4151 (N_4151,N_734,N_1190);
nand U4152 (N_4152,N_563,N_1898);
nand U4153 (N_4153,N_1295,N_1013);
nand U4154 (N_4154,N_1730,N_1496);
nand U4155 (N_4155,N_2874,N_491);
nor U4156 (N_4156,N_1570,N_2213);
or U4157 (N_4157,N_1245,N_2431);
nor U4158 (N_4158,N_315,N_528);
or U4159 (N_4159,N_22,N_754);
and U4160 (N_4160,N_1119,N_2879);
or U4161 (N_4161,N_137,N_1999);
nor U4162 (N_4162,N_218,N_2558);
or U4163 (N_4163,N_2147,N_2466);
nand U4164 (N_4164,N_257,N_2288);
and U4165 (N_4165,N_2057,N_992);
nor U4166 (N_4166,N_2033,N_549);
or U4167 (N_4167,N_2226,N_411);
nor U4168 (N_4168,N_1348,N_2748);
nor U4169 (N_4169,N_1151,N_779);
or U4170 (N_4170,N_594,N_815);
or U4171 (N_4171,N_2295,N_551);
nand U4172 (N_4172,N_2545,N_1521);
nor U4173 (N_4173,N_1706,N_680);
or U4174 (N_4174,N_2354,N_8);
or U4175 (N_4175,N_1873,N_1142);
or U4176 (N_4176,N_2907,N_1708);
and U4177 (N_4177,N_1000,N_1985);
nor U4178 (N_4178,N_1797,N_237);
and U4179 (N_4179,N_982,N_695);
and U4180 (N_4180,N_1310,N_1523);
nor U4181 (N_4181,N_62,N_1979);
and U4182 (N_4182,N_993,N_1578);
and U4183 (N_4183,N_200,N_1813);
nand U4184 (N_4184,N_1691,N_490);
and U4185 (N_4185,N_1748,N_1473);
and U4186 (N_4186,N_1287,N_1391);
or U4187 (N_4187,N_1062,N_493);
nand U4188 (N_4188,N_721,N_2065);
nand U4189 (N_4189,N_2832,N_425);
and U4190 (N_4190,N_1041,N_1290);
nand U4191 (N_4191,N_643,N_1155);
and U4192 (N_4192,N_2114,N_1426);
or U4193 (N_4193,N_1132,N_2752);
nand U4194 (N_4194,N_1519,N_2531);
nor U4195 (N_4195,N_2568,N_2470);
or U4196 (N_4196,N_1266,N_2393);
nand U4197 (N_4197,N_265,N_2119);
or U4198 (N_4198,N_1345,N_2449);
nor U4199 (N_4199,N_2338,N_244);
and U4200 (N_4200,N_944,N_1673);
nor U4201 (N_4201,N_1514,N_1137);
and U4202 (N_4202,N_1728,N_2630);
nor U4203 (N_4203,N_1805,N_2198);
nor U4204 (N_4204,N_596,N_696);
or U4205 (N_4205,N_302,N_2476);
or U4206 (N_4206,N_279,N_2104);
and U4207 (N_4207,N_2090,N_2960);
and U4208 (N_4208,N_2628,N_1508);
nand U4209 (N_4209,N_1424,N_2220);
and U4210 (N_4210,N_1598,N_2714);
nand U4211 (N_4211,N_2282,N_1575);
or U4212 (N_4212,N_1734,N_1964);
or U4213 (N_4213,N_72,N_2139);
xnor U4214 (N_4214,N_1153,N_2865);
nor U4215 (N_4215,N_1765,N_316);
and U4216 (N_4216,N_1633,N_508);
or U4217 (N_4217,N_2658,N_965);
and U4218 (N_4218,N_1422,N_781);
nor U4219 (N_4219,N_1419,N_2156);
nor U4220 (N_4220,N_1571,N_159);
nand U4221 (N_4221,N_1217,N_2663);
and U4222 (N_4222,N_2496,N_1086);
and U4223 (N_4223,N_1447,N_81);
or U4224 (N_4224,N_1224,N_2755);
and U4225 (N_4225,N_1968,N_507);
and U4226 (N_4226,N_2340,N_1775);
nand U4227 (N_4227,N_1092,N_318);
nand U4228 (N_4228,N_788,N_2185);
or U4229 (N_4229,N_440,N_2812);
nand U4230 (N_4230,N_1513,N_180);
nor U4231 (N_4231,N_2061,N_54);
nand U4232 (N_4232,N_2942,N_2860);
and U4233 (N_4233,N_386,N_2629);
nor U4234 (N_4234,N_1037,N_487);
or U4235 (N_4235,N_1435,N_2342);
nor U4236 (N_4236,N_1707,N_2383);
nor U4237 (N_4237,N_1966,N_2596);
nor U4238 (N_4238,N_1699,N_2074);
nand U4239 (N_4239,N_1028,N_264);
and U4240 (N_4240,N_998,N_2196);
nand U4241 (N_4241,N_1864,N_1918);
or U4242 (N_4242,N_2576,N_1645);
nor U4243 (N_4243,N_2954,N_378);
and U4244 (N_4244,N_2996,N_610);
nor U4245 (N_4245,N_1782,N_1840);
and U4246 (N_4246,N_212,N_2845);
and U4247 (N_4247,N_460,N_20);
nor U4248 (N_4248,N_1984,N_2957);
and U4249 (N_4249,N_260,N_2052);
or U4250 (N_4250,N_1638,N_158);
nor U4251 (N_4251,N_135,N_603);
nand U4252 (N_4252,N_1490,N_1335);
nand U4253 (N_4253,N_1269,N_2621);
and U4254 (N_4254,N_2238,N_2786);
nor U4255 (N_4255,N_2232,N_2366);
or U4256 (N_4256,N_1077,N_2248);
nor U4257 (N_4257,N_813,N_717);
or U4258 (N_4258,N_1145,N_1397);
or U4259 (N_4259,N_2432,N_1593);
nand U4260 (N_4260,N_217,N_2581);
and U4261 (N_4261,N_737,N_2314);
nand U4262 (N_4262,N_2456,N_2935);
nand U4263 (N_4263,N_394,N_633);
nand U4264 (N_4264,N_2043,N_1774);
nand U4265 (N_4265,N_1506,N_249);
or U4266 (N_4266,N_1572,N_1812);
and U4267 (N_4267,N_816,N_373);
or U4268 (N_4268,N_538,N_147);
and U4269 (N_4269,N_1470,N_1303);
nand U4270 (N_4270,N_1936,N_1364);
and U4271 (N_4271,N_345,N_947);
nand U4272 (N_4272,N_2936,N_2397);
nor U4273 (N_4273,N_172,N_650);
nor U4274 (N_4274,N_1431,N_1854);
nand U4275 (N_4275,N_71,N_725);
nor U4276 (N_4276,N_2785,N_2749);
or U4277 (N_4277,N_2920,N_1257);
nand U4278 (N_4278,N_1993,N_1143);
or U4279 (N_4279,N_1091,N_911);
nand U4280 (N_4280,N_1356,N_1647);
nor U4281 (N_4281,N_1098,N_2765);
nor U4282 (N_4282,N_2106,N_2281);
nor U4283 (N_4283,N_1108,N_773);
nor U4284 (N_4284,N_2424,N_1278);
or U4285 (N_4285,N_2075,N_2854);
nor U4286 (N_4286,N_2653,N_716);
nand U4287 (N_4287,N_0,N_228);
nor U4288 (N_4288,N_347,N_2569);
nor U4289 (N_4289,N_966,N_1208);
and U4290 (N_4290,N_1323,N_630);
and U4291 (N_4291,N_1176,N_2641);
and U4292 (N_4292,N_417,N_1311);
nand U4293 (N_4293,N_2975,N_2439);
and U4294 (N_4294,N_197,N_2934);
and U4295 (N_4295,N_1386,N_2184);
nor U4296 (N_4296,N_668,N_80);
and U4297 (N_4297,N_1934,N_1648);
nor U4298 (N_4298,N_2896,N_599);
and U4299 (N_4299,N_50,N_2706);
and U4300 (N_4300,N_2207,N_2212);
or U4301 (N_4301,N_451,N_1489);
xor U4302 (N_4302,N_2345,N_1891);
or U4303 (N_4303,N_1741,N_1319);
and U4304 (N_4304,N_743,N_1200);
or U4305 (N_4305,N_571,N_2109);
and U4306 (N_4306,N_741,N_1796);
nor U4307 (N_4307,N_1754,N_78);
nand U4308 (N_4308,N_894,N_2523);
nor U4309 (N_4309,N_659,N_2042);
nor U4310 (N_4310,N_2235,N_2837);
and U4311 (N_4311,N_1070,N_903);
or U4312 (N_4312,N_2351,N_1494);
nand U4313 (N_4313,N_2930,N_126);
nor U4314 (N_4314,N_434,N_1551);
nand U4315 (N_4315,N_727,N_2566);
and U4316 (N_4316,N_2286,N_198);
or U4317 (N_4317,N_79,N_1024);
or U4318 (N_4318,N_2841,N_2030);
nand U4319 (N_4319,N_2546,N_2261);
and U4320 (N_4320,N_2667,N_1794);
nor U4321 (N_4321,N_2183,N_1516);
xor U4322 (N_4322,N_1926,N_2799);
nand U4323 (N_4323,N_1674,N_262);
nand U4324 (N_4324,N_886,N_1446);
nand U4325 (N_4325,N_489,N_409);
and U4326 (N_4326,N_1175,N_742);
nor U4327 (N_4327,N_2979,N_1060);
nor U4328 (N_4328,N_2956,N_2150);
nand U4329 (N_4329,N_2888,N_1802);
nand U4330 (N_4330,N_676,N_1213);
and U4331 (N_4331,N_224,N_420);
nor U4332 (N_4332,N_1526,N_1836);
or U4333 (N_4333,N_1484,N_422);
nor U4334 (N_4334,N_971,N_25);
nor U4335 (N_4335,N_2777,N_2710);
or U4336 (N_4336,N_711,N_704);
nor U4337 (N_4337,N_209,N_1832);
and U4338 (N_4338,N_1271,N_511);
nand U4339 (N_4339,N_2474,N_554);
or U4340 (N_4340,N_2612,N_317);
nor U4341 (N_4341,N_1161,N_2922);
nand U4342 (N_4342,N_2993,N_1556);
or U4343 (N_4343,N_868,N_1543);
and U4344 (N_4344,N_2563,N_2333);
nand U4345 (N_4345,N_792,N_527);
nor U4346 (N_4346,N_1359,N_2696);
nand U4347 (N_4347,N_1860,N_1616);
nor U4348 (N_4348,N_2859,N_1425);
or U4349 (N_4349,N_1202,N_329);
or U4350 (N_4350,N_1306,N_106);
nor U4351 (N_4351,N_57,N_901);
nand U4352 (N_4352,N_2593,N_805);
nand U4353 (N_4353,N_748,N_467);
nand U4354 (N_4354,N_2421,N_1743);
and U4355 (N_4355,N_2495,N_186);
or U4356 (N_4356,N_1635,N_2471);
nand U4357 (N_4357,N_2379,N_2130);
nand U4358 (N_4358,N_2732,N_2813);
nand U4359 (N_4359,N_2277,N_2806);
and U4360 (N_4360,N_2219,N_1605);
nor U4361 (N_4361,N_419,N_2289);
and U4362 (N_4362,N_1075,N_2356);
nand U4363 (N_4363,N_1134,N_144);
nor U4364 (N_4364,N_1031,N_827);
nand U4365 (N_4365,N_2173,N_521);
nor U4366 (N_4366,N_541,N_478);
or U4367 (N_4367,N_2309,N_2792);
or U4368 (N_4368,N_1225,N_2382);
nand U4369 (N_4369,N_2060,N_21);
and U4370 (N_4370,N_2087,N_100);
and U4371 (N_4371,N_1412,N_570);
nor U4372 (N_4372,N_2779,N_2790);
nor U4373 (N_4373,N_852,N_2310);
or U4374 (N_4374,N_1724,N_270);
and U4375 (N_4375,N_2116,N_561);
and U4376 (N_4376,N_1229,N_2557);
nor U4377 (N_4377,N_2143,N_2244);
nand U4378 (N_4378,N_921,N_2023);
nand U4379 (N_4379,N_1914,N_641);
nor U4380 (N_4380,N_1338,N_550);
or U4381 (N_4381,N_1343,N_2429);
and U4382 (N_4382,N_170,N_45);
nor U4383 (N_4383,N_728,N_2135);
or U4384 (N_4384,N_2744,N_732);
nor U4385 (N_4385,N_2864,N_850);
and U4386 (N_4386,N_429,N_2175);
or U4387 (N_4387,N_1532,N_2516);
and U4388 (N_4388,N_2412,N_939);
and U4389 (N_4389,N_1118,N_869);
nand U4390 (N_4390,N_1109,N_1917);
and U4391 (N_4391,N_889,N_1254);
or U4392 (N_4392,N_622,N_2764);
nor U4393 (N_4393,N_506,N_1102);
or U4394 (N_4394,N_587,N_1247);
nor U4395 (N_4395,N_2056,N_837);
and U4396 (N_4396,N_2159,N_1300);
and U4397 (N_4397,N_1539,N_673);
or U4398 (N_4398,N_907,N_2821);
and U4399 (N_4399,N_2943,N_1726);
nand U4400 (N_4400,N_2536,N_2544);
nor U4401 (N_4401,N_361,N_2684);
or U4402 (N_4402,N_1481,N_2843);
nor U4403 (N_4403,N_1197,N_744);
nand U4404 (N_4404,N_2304,N_1085);
or U4405 (N_4405,N_1609,N_1659);
or U4406 (N_4406,N_1535,N_681);
nor U4407 (N_4407,N_938,N_1415);
nor U4408 (N_4408,N_2715,N_974);
nor U4409 (N_4409,N_36,N_188);
or U4410 (N_4410,N_1626,N_252);
nor U4411 (N_4411,N_1453,N_2046);
nor U4412 (N_4412,N_466,N_63);
or U4413 (N_4413,N_2689,N_1036);
nand U4414 (N_4414,N_770,N_1976);
nor U4415 (N_4415,N_70,N_2487);
and U4416 (N_4416,N_1414,N_1883);
nor U4417 (N_4417,N_2819,N_2810);
and U4418 (N_4418,N_58,N_1100);
and U4419 (N_4419,N_2165,N_2522);
nand U4420 (N_4420,N_769,N_1907);
nand U4421 (N_4421,N_1468,N_1362);
nand U4422 (N_4422,N_76,N_2909);
or U4423 (N_4423,N_2115,N_2096);
and U4424 (N_4424,N_739,N_1677);
nand U4425 (N_4425,N_2164,N_1402);
and U4426 (N_4426,N_1554,N_250);
or U4427 (N_4427,N_757,N_1404);
nand U4428 (N_4428,N_898,N_2902);
and U4429 (N_4429,N_2105,N_1246);
nor U4430 (N_4430,N_720,N_1089);
nor U4431 (N_4431,N_2418,N_445);
nand U4432 (N_4432,N_819,N_210);
and U4433 (N_4433,N_26,N_1443);
nor U4434 (N_4434,N_220,N_1256);
nand U4435 (N_4435,N_793,N_2697);
and U4436 (N_4436,N_1595,N_1396);
nand U4437 (N_4437,N_1772,N_75);
and U4438 (N_4438,N_60,N_715);
nand U4439 (N_4439,N_2188,N_2025);
nand U4440 (N_4440,N_2761,N_107);
and U4441 (N_4441,N_635,N_1852);
or U4442 (N_4442,N_196,N_154);
nor U4443 (N_4443,N_2727,N_2194);
xor U4444 (N_4444,N_34,N_851);
nand U4445 (N_4445,N_2751,N_1937);
and U4446 (N_4446,N_2535,N_1439);
and U4447 (N_4447,N_2324,N_905);
and U4448 (N_4448,N_406,N_2890);
and U4449 (N_4449,N_2971,N_529);
and U4450 (N_4450,N_167,N_215);
and U4451 (N_4451,N_2124,N_1711);
nor U4452 (N_4452,N_1218,N_2589);
nor U4453 (N_4453,N_288,N_2642);
nand U4454 (N_4454,N_916,N_2949);
nor U4455 (N_4455,N_1307,N_545);
nor U4456 (N_4456,N_410,N_962);
or U4457 (N_4457,N_655,N_1101);
nor U4458 (N_4458,N_1887,N_2398);
nand U4459 (N_4459,N_266,N_2305);
nor U4460 (N_4460,N_1052,N_688);
and U4461 (N_4461,N_1603,N_2635);
and U4462 (N_4462,N_567,N_1644);
or U4463 (N_4463,N_2242,N_682);
nand U4464 (N_4464,N_565,N_967);
or U4465 (N_4465,N_2015,N_2062);
nand U4466 (N_4466,N_202,N_307);
nor U4467 (N_4467,N_1884,N_1281);
and U4468 (N_4468,N_277,N_2386);
and U4469 (N_4469,N_1611,N_1742);
nor U4470 (N_4470,N_2072,N_399);
nor U4471 (N_4471,N_1977,N_199);
and U4472 (N_4472,N_2154,N_300);
nand U4473 (N_4473,N_2726,N_1087);
and U4474 (N_4474,N_1126,N_234);
or U4475 (N_4475,N_2769,N_1033);
and U4476 (N_4476,N_2002,N_945);
nor U4477 (N_4477,N_495,N_2204);
or U4478 (N_4478,N_18,N_1233);
and U4479 (N_4479,N_2605,N_2958);
nor U4480 (N_4480,N_1943,N_247);
nand U4481 (N_4481,N_2534,N_1756);
or U4482 (N_4482,N_500,N_502);
nor U4483 (N_4483,N_1905,N_1430);
or U4484 (N_4484,N_53,N_1669);
nor U4485 (N_4485,N_1776,N_2963);
nor U4486 (N_4486,N_1094,N_1298);
or U4487 (N_4487,N_1337,N_2047);
and U4488 (N_4488,N_835,N_878);
and U4489 (N_4489,N_572,N_802);
nor U4490 (N_4490,N_513,N_1546);
and U4491 (N_4491,N_2784,N_836);
nand U4492 (N_4492,N_2973,N_2914);
nor U4493 (N_4493,N_2538,N_442);
or U4494 (N_4494,N_1567,N_2138);
or U4495 (N_4495,N_1038,N_2488);
nor U4496 (N_4496,N_1379,N_2472);
or U4497 (N_4497,N_834,N_763);
and U4498 (N_4498,N_946,N_1910);
or U4499 (N_4499,N_648,N_2881);
nand U4500 (N_4500,N_2006,N_370);
and U4501 (N_4501,N_191,N_308);
and U4502 (N_4502,N_1268,N_2554);
or U4503 (N_4503,N_492,N_933);
nand U4504 (N_4504,N_497,N_962);
and U4505 (N_4505,N_1399,N_1559);
nand U4506 (N_4506,N_2046,N_192);
or U4507 (N_4507,N_2718,N_2164);
nand U4508 (N_4508,N_1822,N_1448);
and U4509 (N_4509,N_77,N_1354);
and U4510 (N_4510,N_736,N_1226);
and U4511 (N_4511,N_1392,N_1813);
or U4512 (N_4512,N_2418,N_2558);
and U4513 (N_4513,N_375,N_373);
and U4514 (N_4514,N_1554,N_639);
or U4515 (N_4515,N_1538,N_2319);
nand U4516 (N_4516,N_1415,N_102);
or U4517 (N_4517,N_2978,N_2308);
nand U4518 (N_4518,N_1767,N_196);
nor U4519 (N_4519,N_2937,N_1392);
nand U4520 (N_4520,N_294,N_428);
or U4521 (N_4521,N_2236,N_1103);
or U4522 (N_4522,N_1307,N_2452);
or U4523 (N_4523,N_2860,N_174);
nor U4524 (N_4524,N_1980,N_2126);
or U4525 (N_4525,N_2809,N_210);
or U4526 (N_4526,N_798,N_830);
xnor U4527 (N_4527,N_2773,N_1487);
nor U4528 (N_4528,N_2768,N_1774);
or U4529 (N_4529,N_1080,N_172);
nand U4530 (N_4530,N_894,N_1767);
nor U4531 (N_4531,N_1890,N_1578);
or U4532 (N_4532,N_1969,N_1470);
and U4533 (N_4533,N_2493,N_1892);
or U4534 (N_4534,N_2877,N_547);
and U4535 (N_4535,N_520,N_1929);
or U4536 (N_4536,N_1981,N_1724);
nor U4537 (N_4537,N_1783,N_2096);
or U4538 (N_4538,N_2722,N_2354);
and U4539 (N_4539,N_1855,N_375);
and U4540 (N_4540,N_249,N_272);
nor U4541 (N_4541,N_433,N_655);
and U4542 (N_4542,N_2274,N_2486);
and U4543 (N_4543,N_1168,N_1201);
nor U4544 (N_4544,N_2272,N_2842);
and U4545 (N_4545,N_860,N_84);
or U4546 (N_4546,N_2990,N_1600);
and U4547 (N_4547,N_658,N_2952);
nor U4548 (N_4548,N_1554,N_775);
nor U4549 (N_4549,N_2425,N_2359);
or U4550 (N_4550,N_641,N_2835);
or U4551 (N_4551,N_1711,N_2555);
nand U4552 (N_4552,N_996,N_1526);
nand U4553 (N_4553,N_158,N_2312);
and U4554 (N_4554,N_575,N_160);
nor U4555 (N_4555,N_884,N_2304);
and U4556 (N_4556,N_2114,N_11);
nor U4557 (N_4557,N_808,N_2726);
and U4558 (N_4558,N_2795,N_2881);
or U4559 (N_4559,N_956,N_2314);
nor U4560 (N_4560,N_1042,N_862);
or U4561 (N_4561,N_2106,N_528);
nand U4562 (N_4562,N_512,N_350);
nand U4563 (N_4563,N_1699,N_415);
nand U4564 (N_4564,N_765,N_2159);
nand U4565 (N_4565,N_1100,N_1017);
or U4566 (N_4566,N_525,N_2565);
nand U4567 (N_4567,N_1683,N_1964);
and U4568 (N_4568,N_2964,N_2873);
or U4569 (N_4569,N_2612,N_214);
and U4570 (N_4570,N_2751,N_682);
or U4571 (N_4571,N_380,N_2482);
nor U4572 (N_4572,N_819,N_2646);
and U4573 (N_4573,N_2142,N_1025);
nand U4574 (N_4574,N_579,N_2539);
nand U4575 (N_4575,N_891,N_2652);
nor U4576 (N_4576,N_2847,N_2221);
nor U4577 (N_4577,N_33,N_2216);
xor U4578 (N_4578,N_2355,N_206);
nand U4579 (N_4579,N_1585,N_2536);
nand U4580 (N_4580,N_949,N_1866);
nand U4581 (N_4581,N_1586,N_1216);
nor U4582 (N_4582,N_2594,N_850);
nand U4583 (N_4583,N_1392,N_69);
nand U4584 (N_4584,N_977,N_679);
and U4585 (N_4585,N_2837,N_1537);
nor U4586 (N_4586,N_2034,N_210);
or U4587 (N_4587,N_818,N_1750);
nand U4588 (N_4588,N_394,N_2139);
nand U4589 (N_4589,N_2488,N_1522);
and U4590 (N_4590,N_642,N_1175);
nor U4591 (N_4591,N_2176,N_948);
nor U4592 (N_4592,N_1089,N_708);
nand U4593 (N_4593,N_473,N_691);
nor U4594 (N_4594,N_1741,N_1756);
nand U4595 (N_4595,N_724,N_458);
nand U4596 (N_4596,N_2970,N_1640);
and U4597 (N_4597,N_1436,N_2389);
and U4598 (N_4598,N_1048,N_1309);
or U4599 (N_4599,N_2758,N_1015);
nand U4600 (N_4600,N_719,N_118);
nand U4601 (N_4601,N_606,N_1593);
or U4602 (N_4602,N_2001,N_554);
or U4603 (N_4603,N_2514,N_2745);
and U4604 (N_4604,N_445,N_1159);
or U4605 (N_4605,N_2931,N_2744);
and U4606 (N_4606,N_2536,N_1986);
and U4607 (N_4607,N_989,N_54);
nor U4608 (N_4608,N_474,N_1462);
or U4609 (N_4609,N_2526,N_589);
or U4610 (N_4610,N_2253,N_1084);
nor U4611 (N_4611,N_168,N_97);
nand U4612 (N_4612,N_496,N_2373);
and U4613 (N_4613,N_1102,N_627);
nand U4614 (N_4614,N_298,N_651);
and U4615 (N_4615,N_1351,N_907);
and U4616 (N_4616,N_48,N_2084);
and U4617 (N_4617,N_2358,N_1026);
nand U4618 (N_4618,N_2893,N_347);
or U4619 (N_4619,N_1560,N_2276);
or U4620 (N_4620,N_2900,N_2795);
and U4621 (N_4621,N_177,N_1584);
or U4622 (N_4622,N_1909,N_996);
or U4623 (N_4623,N_2431,N_2051);
or U4624 (N_4624,N_2024,N_886);
nor U4625 (N_4625,N_293,N_1856);
and U4626 (N_4626,N_1177,N_1569);
nor U4627 (N_4627,N_256,N_530);
nor U4628 (N_4628,N_716,N_2670);
or U4629 (N_4629,N_509,N_1365);
or U4630 (N_4630,N_455,N_407);
nand U4631 (N_4631,N_1023,N_2575);
nor U4632 (N_4632,N_2164,N_2734);
nor U4633 (N_4633,N_80,N_2387);
nor U4634 (N_4634,N_2618,N_2066);
and U4635 (N_4635,N_1442,N_2421);
nor U4636 (N_4636,N_1392,N_2330);
nand U4637 (N_4637,N_322,N_1324);
xnor U4638 (N_4638,N_1306,N_2946);
and U4639 (N_4639,N_1204,N_725);
and U4640 (N_4640,N_8,N_2346);
nand U4641 (N_4641,N_2471,N_1431);
nor U4642 (N_4642,N_730,N_1187);
nor U4643 (N_4643,N_200,N_2201);
nand U4644 (N_4644,N_2186,N_2699);
nand U4645 (N_4645,N_1554,N_2845);
or U4646 (N_4646,N_55,N_1102);
nand U4647 (N_4647,N_56,N_1918);
nand U4648 (N_4648,N_287,N_2323);
and U4649 (N_4649,N_16,N_1610);
nand U4650 (N_4650,N_492,N_116);
and U4651 (N_4651,N_2090,N_2820);
or U4652 (N_4652,N_1790,N_2155);
and U4653 (N_4653,N_615,N_1955);
nor U4654 (N_4654,N_240,N_1062);
or U4655 (N_4655,N_1904,N_2488);
or U4656 (N_4656,N_2669,N_2584);
nand U4657 (N_4657,N_2667,N_1383);
and U4658 (N_4658,N_2010,N_888);
or U4659 (N_4659,N_537,N_100);
or U4660 (N_4660,N_387,N_2457);
nand U4661 (N_4661,N_495,N_2830);
nor U4662 (N_4662,N_1740,N_1591);
or U4663 (N_4663,N_1274,N_1735);
and U4664 (N_4664,N_2597,N_997);
or U4665 (N_4665,N_165,N_2214);
and U4666 (N_4666,N_849,N_790);
or U4667 (N_4667,N_1163,N_78);
and U4668 (N_4668,N_2921,N_1563);
and U4669 (N_4669,N_653,N_1768);
and U4670 (N_4670,N_2871,N_1028);
and U4671 (N_4671,N_420,N_2288);
nor U4672 (N_4672,N_285,N_1248);
nor U4673 (N_4673,N_1935,N_620);
or U4674 (N_4674,N_2465,N_2079);
nand U4675 (N_4675,N_2231,N_612);
nand U4676 (N_4676,N_1912,N_429);
and U4677 (N_4677,N_1462,N_436);
and U4678 (N_4678,N_2218,N_1181);
and U4679 (N_4679,N_2324,N_1000);
nor U4680 (N_4680,N_1524,N_2384);
or U4681 (N_4681,N_2806,N_2785);
nand U4682 (N_4682,N_2359,N_1328);
or U4683 (N_4683,N_1572,N_2556);
or U4684 (N_4684,N_2317,N_677);
and U4685 (N_4685,N_647,N_1960);
and U4686 (N_4686,N_539,N_1272);
and U4687 (N_4687,N_1973,N_726);
nor U4688 (N_4688,N_1037,N_2120);
or U4689 (N_4689,N_2439,N_1981);
nand U4690 (N_4690,N_38,N_2240);
nor U4691 (N_4691,N_493,N_2833);
and U4692 (N_4692,N_2902,N_2668);
nor U4693 (N_4693,N_2290,N_2226);
or U4694 (N_4694,N_2168,N_1657);
xnor U4695 (N_4695,N_2231,N_1873);
or U4696 (N_4696,N_1496,N_1373);
or U4697 (N_4697,N_1182,N_400);
and U4698 (N_4698,N_1621,N_2966);
and U4699 (N_4699,N_2610,N_714);
and U4700 (N_4700,N_1456,N_2317);
nor U4701 (N_4701,N_545,N_2001);
nor U4702 (N_4702,N_1925,N_1262);
and U4703 (N_4703,N_2784,N_1936);
and U4704 (N_4704,N_2831,N_226);
nand U4705 (N_4705,N_403,N_256);
nor U4706 (N_4706,N_922,N_1091);
nor U4707 (N_4707,N_1549,N_2619);
and U4708 (N_4708,N_2191,N_2050);
nand U4709 (N_4709,N_1004,N_2217);
or U4710 (N_4710,N_1076,N_770);
and U4711 (N_4711,N_2468,N_2537);
nand U4712 (N_4712,N_935,N_717);
or U4713 (N_4713,N_1854,N_2517);
nor U4714 (N_4714,N_2101,N_1081);
nand U4715 (N_4715,N_2632,N_2693);
nor U4716 (N_4716,N_1443,N_2637);
or U4717 (N_4717,N_1573,N_2823);
nor U4718 (N_4718,N_1743,N_2632);
nor U4719 (N_4719,N_2065,N_307);
nor U4720 (N_4720,N_2385,N_1818);
and U4721 (N_4721,N_2383,N_255);
and U4722 (N_4722,N_1489,N_649);
or U4723 (N_4723,N_2517,N_792);
and U4724 (N_4724,N_10,N_2553);
or U4725 (N_4725,N_2250,N_127);
nor U4726 (N_4726,N_2825,N_1361);
nor U4727 (N_4727,N_63,N_1279);
nand U4728 (N_4728,N_472,N_2884);
nor U4729 (N_4729,N_2889,N_2620);
nor U4730 (N_4730,N_986,N_2168);
nor U4731 (N_4731,N_833,N_2305);
nand U4732 (N_4732,N_1394,N_1983);
or U4733 (N_4733,N_554,N_2476);
and U4734 (N_4734,N_1915,N_2517);
and U4735 (N_4735,N_230,N_755);
nor U4736 (N_4736,N_984,N_2156);
or U4737 (N_4737,N_1591,N_2294);
nand U4738 (N_4738,N_772,N_528);
nor U4739 (N_4739,N_368,N_2850);
or U4740 (N_4740,N_81,N_2668);
nand U4741 (N_4741,N_1723,N_552);
or U4742 (N_4742,N_2131,N_1975);
nand U4743 (N_4743,N_2398,N_1312);
nor U4744 (N_4744,N_2425,N_2773);
and U4745 (N_4745,N_318,N_1871);
and U4746 (N_4746,N_1856,N_1653);
or U4747 (N_4747,N_1122,N_554);
nor U4748 (N_4748,N_1021,N_1616);
nor U4749 (N_4749,N_311,N_2486);
or U4750 (N_4750,N_2425,N_701);
and U4751 (N_4751,N_215,N_1683);
nand U4752 (N_4752,N_2051,N_2410);
nand U4753 (N_4753,N_685,N_71);
nand U4754 (N_4754,N_2915,N_474);
nor U4755 (N_4755,N_2201,N_129);
or U4756 (N_4756,N_231,N_1105);
nor U4757 (N_4757,N_1591,N_471);
nor U4758 (N_4758,N_530,N_752);
nor U4759 (N_4759,N_203,N_2163);
nand U4760 (N_4760,N_1254,N_2805);
nor U4761 (N_4761,N_2107,N_1437);
nand U4762 (N_4762,N_2399,N_1874);
nor U4763 (N_4763,N_1823,N_2943);
nand U4764 (N_4764,N_490,N_640);
nand U4765 (N_4765,N_1642,N_761);
and U4766 (N_4766,N_884,N_236);
nand U4767 (N_4767,N_2751,N_1771);
and U4768 (N_4768,N_877,N_1728);
or U4769 (N_4769,N_784,N_666);
nand U4770 (N_4770,N_2212,N_243);
or U4771 (N_4771,N_1842,N_87);
nor U4772 (N_4772,N_2313,N_2965);
and U4773 (N_4773,N_392,N_1268);
or U4774 (N_4774,N_2431,N_2055);
nor U4775 (N_4775,N_371,N_50);
and U4776 (N_4776,N_677,N_1671);
and U4777 (N_4777,N_637,N_1325);
and U4778 (N_4778,N_845,N_1204);
or U4779 (N_4779,N_1096,N_4);
or U4780 (N_4780,N_571,N_453);
or U4781 (N_4781,N_1053,N_2436);
nand U4782 (N_4782,N_2436,N_2035);
nor U4783 (N_4783,N_2714,N_2019);
or U4784 (N_4784,N_1691,N_1839);
and U4785 (N_4785,N_2158,N_718);
nor U4786 (N_4786,N_2682,N_941);
nor U4787 (N_4787,N_997,N_1941);
nand U4788 (N_4788,N_875,N_298);
and U4789 (N_4789,N_436,N_190);
and U4790 (N_4790,N_836,N_1574);
nand U4791 (N_4791,N_2207,N_311);
nand U4792 (N_4792,N_230,N_354);
and U4793 (N_4793,N_2162,N_2112);
nor U4794 (N_4794,N_2219,N_2078);
nand U4795 (N_4795,N_254,N_1216);
nand U4796 (N_4796,N_1843,N_1595);
and U4797 (N_4797,N_2578,N_1367);
and U4798 (N_4798,N_397,N_890);
nor U4799 (N_4799,N_1228,N_810);
nor U4800 (N_4800,N_771,N_198);
or U4801 (N_4801,N_1703,N_1005);
nand U4802 (N_4802,N_2969,N_639);
nor U4803 (N_4803,N_1839,N_2346);
nand U4804 (N_4804,N_612,N_2908);
nor U4805 (N_4805,N_791,N_777);
or U4806 (N_4806,N_1241,N_2522);
nand U4807 (N_4807,N_1950,N_565);
and U4808 (N_4808,N_1882,N_1955);
nand U4809 (N_4809,N_488,N_2550);
nor U4810 (N_4810,N_1183,N_9);
xnor U4811 (N_4811,N_821,N_2849);
or U4812 (N_4812,N_626,N_2211);
nor U4813 (N_4813,N_2379,N_1533);
nor U4814 (N_4814,N_2231,N_2926);
or U4815 (N_4815,N_1192,N_2250);
nor U4816 (N_4816,N_2297,N_1514);
nand U4817 (N_4817,N_2689,N_2969);
nand U4818 (N_4818,N_33,N_127);
or U4819 (N_4819,N_307,N_1099);
and U4820 (N_4820,N_1130,N_152);
nor U4821 (N_4821,N_2129,N_308);
nor U4822 (N_4822,N_1965,N_2856);
or U4823 (N_4823,N_1121,N_691);
nand U4824 (N_4824,N_538,N_2309);
nand U4825 (N_4825,N_747,N_612);
xnor U4826 (N_4826,N_2342,N_1783);
or U4827 (N_4827,N_1110,N_1609);
or U4828 (N_4828,N_1359,N_1965);
nand U4829 (N_4829,N_724,N_1262);
nor U4830 (N_4830,N_2284,N_340);
nand U4831 (N_4831,N_410,N_2408);
and U4832 (N_4832,N_330,N_388);
nand U4833 (N_4833,N_1031,N_1121);
or U4834 (N_4834,N_2599,N_329);
or U4835 (N_4835,N_1695,N_2830);
and U4836 (N_4836,N_2553,N_2916);
or U4837 (N_4837,N_562,N_2669);
or U4838 (N_4838,N_665,N_1112);
nor U4839 (N_4839,N_978,N_968);
xnor U4840 (N_4840,N_1719,N_1117);
nand U4841 (N_4841,N_147,N_1571);
and U4842 (N_4842,N_2973,N_1030);
and U4843 (N_4843,N_1714,N_2684);
xor U4844 (N_4844,N_1098,N_1415);
or U4845 (N_4845,N_1104,N_1915);
nor U4846 (N_4846,N_2097,N_2654);
or U4847 (N_4847,N_25,N_1879);
nand U4848 (N_4848,N_1085,N_453);
and U4849 (N_4849,N_203,N_1012);
nor U4850 (N_4850,N_363,N_498);
or U4851 (N_4851,N_244,N_439);
and U4852 (N_4852,N_2088,N_783);
nor U4853 (N_4853,N_2672,N_651);
and U4854 (N_4854,N_2637,N_2651);
nor U4855 (N_4855,N_157,N_1022);
or U4856 (N_4856,N_78,N_2321);
or U4857 (N_4857,N_2275,N_723);
or U4858 (N_4858,N_2929,N_977);
nor U4859 (N_4859,N_2844,N_2556);
nor U4860 (N_4860,N_686,N_2104);
and U4861 (N_4861,N_714,N_1216);
and U4862 (N_4862,N_1091,N_2236);
and U4863 (N_4863,N_2148,N_1824);
and U4864 (N_4864,N_1216,N_246);
nor U4865 (N_4865,N_1863,N_2238);
and U4866 (N_4866,N_15,N_1967);
nor U4867 (N_4867,N_1326,N_608);
or U4868 (N_4868,N_2738,N_587);
or U4869 (N_4869,N_1594,N_1989);
or U4870 (N_4870,N_1119,N_1695);
nand U4871 (N_4871,N_362,N_2753);
xnor U4872 (N_4872,N_728,N_605);
and U4873 (N_4873,N_2815,N_884);
nand U4874 (N_4874,N_2968,N_571);
or U4875 (N_4875,N_961,N_1260);
nor U4876 (N_4876,N_1537,N_31);
nand U4877 (N_4877,N_2550,N_2818);
or U4878 (N_4878,N_2734,N_2785);
and U4879 (N_4879,N_1169,N_2915);
nor U4880 (N_4880,N_800,N_2935);
nor U4881 (N_4881,N_842,N_597);
nand U4882 (N_4882,N_1751,N_608);
nand U4883 (N_4883,N_789,N_247);
nor U4884 (N_4884,N_1014,N_2962);
nor U4885 (N_4885,N_1163,N_766);
nand U4886 (N_4886,N_1527,N_1850);
or U4887 (N_4887,N_2799,N_1539);
nor U4888 (N_4888,N_542,N_2192);
nand U4889 (N_4889,N_1868,N_1324);
nand U4890 (N_4890,N_290,N_343);
and U4891 (N_4891,N_514,N_1116);
or U4892 (N_4892,N_367,N_806);
nor U4893 (N_4893,N_2678,N_771);
nand U4894 (N_4894,N_1149,N_2192);
or U4895 (N_4895,N_2979,N_111);
or U4896 (N_4896,N_2792,N_2587);
nand U4897 (N_4897,N_162,N_1053);
nand U4898 (N_4898,N_2579,N_787);
nand U4899 (N_4899,N_189,N_1779);
nand U4900 (N_4900,N_1980,N_654);
nor U4901 (N_4901,N_2523,N_1671);
or U4902 (N_4902,N_1790,N_2674);
or U4903 (N_4903,N_2875,N_1790);
nor U4904 (N_4904,N_887,N_1622);
nand U4905 (N_4905,N_2773,N_888);
or U4906 (N_4906,N_1358,N_49);
nand U4907 (N_4907,N_1759,N_1188);
and U4908 (N_4908,N_1222,N_1774);
nand U4909 (N_4909,N_1957,N_743);
nand U4910 (N_4910,N_1876,N_2006);
and U4911 (N_4911,N_1548,N_2693);
nand U4912 (N_4912,N_1984,N_602);
and U4913 (N_4913,N_1678,N_514);
nor U4914 (N_4914,N_195,N_2014);
and U4915 (N_4915,N_2255,N_1148);
nand U4916 (N_4916,N_2574,N_920);
nor U4917 (N_4917,N_964,N_2787);
and U4918 (N_4918,N_895,N_894);
and U4919 (N_4919,N_468,N_778);
nand U4920 (N_4920,N_2766,N_1400);
nor U4921 (N_4921,N_2807,N_999);
nand U4922 (N_4922,N_759,N_28);
nand U4923 (N_4923,N_530,N_677);
nor U4924 (N_4924,N_1936,N_863);
nor U4925 (N_4925,N_1531,N_2361);
nand U4926 (N_4926,N_2679,N_1122);
nand U4927 (N_4927,N_2354,N_1750);
nor U4928 (N_4928,N_2333,N_1039);
nand U4929 (N_4929,N_2852,N_2168);
nor U4930 (N_4930,N_2981,N_1795);
nand U4931 (N_4931,N_1608,N_1387);
xor U4932 (N_4932,N_1752,N_337);
or U4933 (N_4933,N_1036,N_57);
nor U4934 (N_4934,N_2941,N_730);
or U4935 (N_4935,N_1634,N_1660);
or U4936 (N_4936,N_2389,N_1312);
nand U4937 (N_4937,N_864,N_2346);
or U4938 (N_4938,N_1128,N_2222);
nand U4939 (N_4939,N_2081,N_2573);
nor U4940 (N_4940,N_1023,N_2437);
and U4941 (N_4941,N_1214,N_1716);
and U4942 (N_4942,N_2109,N_2383);
nor U4943 (N_4943,N_2341,N_2003);
nand U4944 (N_4944,N_1375,N_385);
nand U4945 (N_4945,N_1287,N_802);
nand U4946 (N_4946,N_1282,N_2977);
or U4947 (N_4947,N_1977,N_2665);
and U4948 (N_4948,N_2783,N_1149);
and U4949 (N_4949,N_203,N_2229);
and U4950 (N_4950,N_173,N_9);
and U4951 (N_4951,N_1652,N_691);
nand U4952 (N_4952,N_851,N_1064);
nor U4953 (N_4953,N_378,N_662);
or U4954 (N_4954,N_1596,N_33);
or U4955 (N_4955,N_1829,N_635);
nand U4956 (N_4956,N_2809,N_1083);
nor U4957 (N_4957,N_2655,N_1596);
and U4958 (N_4958,N_2584,N_2869);
nand U4959 (N_4959,N_2050,N_1273);
nand U4960 (N_4960,N_1036,N_2188);
nor U4961 (N_4961,N_2814,N_2829);
nor U4962 (N_4962,N_1722,N_2525);
or U4963 (N_4963,N_736,N_2919);
nand U4964 (N_4964,N_2169,N_1740);
nor U4965 (N_4965,N_2888,N_1092);
nor U4966 (N_4966,N_24,N_1599);
or U4967 (N_4967,N_2944,N_1868);
nand U4968 (N_4968,N_1561,N_257);
xor U4969 (N_4969,N_644,N_1365);
or U4970 (N_4970,N_2378,N_1755);
nand U4971 (N_4971,N_2806,N_2228);
or U4972 (N_4972,N_2867,N_668);
nor U4973 (N_4973,N_404,N_2503);
nand U4974 (N_4974,N_2665,N_1947);
and U4975 (N_4975,N_1952,N_2562);
and U4976 (N_4976,N_1598,N_2809);
and U4977 (N_4977,N_2599,N_2523);
or U4978 (N_4978,N_1760,N_2963);
nand U4979 (N_4979,N_2975,N_2114);
or U4980 (N_4980,N_1733,N_283);
or U4981 (N_4981,N_1724,N_714);
nand U4982 (N_4982,N_480,N_2842);
nand U4983 (N_4983,N_481,N_1175);
nor U4984 (N_4984,N_1103,N_2587);
and U4985 (N_4985,N_477,N_211);
or U4986 (N_4986,N_2051,N_2642);
and U4987 (N_4987,N_1850,N_2102);
or U4988 (N_4988,N_1726,N_540);
nand U4989 (N_4989,N_2349,N_1430);
nor U4990 (N_4990,N_1234,N_1353);
nand U4991 (N_4991,N_2524,N_38);
nand U4992 (N_4992,N_1075,N_2646);
and U4993 (N_4993,N_705,N_431);
or U4994 (N_4994,N_1913,N_1524);
nor U4995 (N_4995,N_2896,N_1218);
and U4996 (N_4996,N_64,N_1268);
nand U4997 (N_4997,N_345,N_1272);
or U4998 (N_4998,N_2122,N_2793);
nor U4999 (N_4999,N_2753,N_1635);
and U5000 (N_5000,N_1039,N_2568);
nor U5001 (N_5001,N_355,N_812);
nand U5002 (N_5002,N_2422,N_1300);
or U5003 (N_5003,N_1330,N_2454);
or U5004 (N_5004,N_1306,N_716);
nand U5005 (N_5005,N_2044,N_2516);
nand U5006 (N_5006,N_2087,N_2564);
and U5007 (N_5007,N_2076,N_2127);
nor U5008 (N_5008,N_1783,N_632);
or U5009 (N_5009,N_257,N_1938);
or U5010 (N_5010,N_643,N_239);
nor U5011 (N_5011,N_725,N_1481);
nor U5012 (N_5012,N_2453,N_534);
and U5013 (N_5013,N_2062,N_1964);
nor U5014 (N_5014,N_2421,N_2730);
nor U5015 (N_5015,N_2748,N_1889);
nand U5016 (N_5016,N_2377,N_2042);
and U5017 (N_5017,N_1588,N_1817);
or U5018 (N_5018,N_73,N_2251);
or U5019 (N_5019,N_70,N_2313);
xnor U5020 (N_5020,N_1463,N_1449);
or U5021 (N_5021,N_270,N_1770);
nor U5022 (N_5022,N_510,N_1122);
and U5023 (N_5023,N_2755,N_1207);
nand U5024 (N_5024,N_330,N_371);
xor U5025 (N_5025,N_2479,N_2681);
and U5026 (N_5026,N_2927,N_880);
nand U5027 (N_5027,N_1848,N_2657);
or U5028 (N_5028,N_2319,N_1546);
nand U5029 (N_5029,N_1956,N_208);
nor U5030 (N_5030,N_2333,N_1183);
or U5031 (N_5031,N_2259,N_2129);
or U5032 (N_5032,N_375,N_2091);
or U5033 (N_5033,N_753,N_1215);
xor U5034 (N_5034,N_989,N_126);
and U5035 (N_5035,N_2874,N_1006);
and U5036 (N_5036,N_2897,N_1183);
nand U5037 (N_5037,N_46,N_306);
nand U5038 (N_5038,N_1452,N_1508);
nor U5039 (N_5039,N_2422,N_1079);
and U5040 (N_5040,N_1547,N_1466);
nor U5041 (N_5041,N_2437,N_2930);
and U5042 (N_5042,N_360,N_1814);
and U5043 (N_5043,N_726,N_2086);
and U5044 (N_5044,N_221,N_2656);
nand U5045 (N_5045,N_733,N_345);
nand U5046 (N_5046,N_897,N_2384);
nor U5047 (N_5047,N_1057,N_2491);
and U5048 (N_5048,N_956,N_1874);
nor U5049 (N_5049,N_1588,N_230);
or U5050 (N_5050,N_2518,N_2975);
and U5051 (N_5051,N_911,N_1826);
nor U5052 (N_5052,N_2129,N_2637);
nor U5053 (N_5053,N_1968,N_1306);
nor U5054 (N_5054,N_654,N_1956);
nor U5055 (N_5055,N_1270,N_2960);
or U5056 (N_5056,N_2500,N_1042);
nand U5057 (N_5057,N_238,N_645);
and U5058 (N_5058,N_2782,N_1125);
nor U5059 (N_5059,N_2712,N_1881);
or U5060 (N_5060,N_953,N_978);
or U5061 (N_5061,N_518,N_1489);
nor U5062 (N_5062,N_751,N_2657);
nand U5063 (N_5063,N_1063,N_2065);
nor U5064 (N_5064,N_100,N_1166);
or U5065 (N_5065,N_2664,N_1514);
nor U5066 (N_5066,N_289,N_2195);
and U5067 (N_5067,N_335,N_833);
nor U5068 (N_5068,N_420,N_2860);
nor U5069 (N_5069,N_1213,N_1924);
and U5070 (N_5070,N_324,N_2798);
nor U5071 (N_5071,N_2405,N_1618);
nor U5072 (N_5072,N_1143,N_1371);
and U5073 (N_5073,N_286,N_1662);
nand U5074 (N_5074,N_2451,N_2700);
nor U5075 (N_5075,N_593,N_1153);
nand U5076 (N_5076,N_1301,N_638);
and U5077 (N_5077,N_322,N_43);
nand U5078 (N_5078,N_1217,N_555);
and U5079 (N_5079,N_2999,N_1329);
and U5080 (N_5080,N_1549,N_2580);
nand U5081 (N_5081,N_2218,N_2577);
or U5082 (N_5082,N_1857,N_2792);
or U5083 (N_5083,N_1123,N_277);
nor U5084 (N_5084,N_738,N_2557);
nand U5085 (N_5085,N_271,N_2372);
nor U5086 (N_5086,N_2486,N_924);
or U5087 (N_5087,N_568,N_418);
nor U5088 (N_5088,N_1989,N_2565);
or U5089 (N_5089,N_2763,N_2706);
or U5090 (N_5090,N_279,N_1141);
or U5091 (N_5091,N_2306,N_2688);
nand U5092 (N_5092,N_495,N_2097);
or U5093 (N_5093,N_2180,N_1397);
nor U5094 (N_5094,N_2485,N_2537);
nand U5095 (N_5095,N_2563,N_2656);
nand U5096 (N_5096,N_1369,N_1558);
nor U5097 (N_5097,N_907,N_2386);
nand U5098 (N_5098,N_1772,N_1857);
nand U5099 (N_5099,N_2333,N_1481);
nand U5100 (N_5100,N_863,N_1695);
nand U5101 (N_5101,N_1489,N_2488);
nor U5102 (N_5102,N_778,N_2937);
xnor U5103 (N_5103,N_1181,N_2267);
and U5104 (N_5104,N_416,N_54);
nor U5105 (N_5105,N_106,N_1705);
nor U5106 (N_5106,N_1744,N_678);
or U5107 (N_5107,N_350,N_1923);
nand U5108 (N_5108,N_974,N_2320);
nand U5109 (N_5109,N_1875,N_2224);
or U5110 (N_5110,N_1491,N_2036);
nor U5111 (N_5111,N_708,N_2077);
or U5112 (N_5112,N_1523,N_1894);
nor U5113 (N_5113,N_795,N_235);
nand U5114 (N_5114,N_2621,N_185);
nand U5115 (N_5115,N_982,N_2710);
nand U5116 (N_5116,N_905,N_987);
or U5117 (N_5117,N_2725,N_15);
nand U5118 (N_5118,N_167,N_431);
or U5119 (N_5119,N_2346,N_670);
nor U5120 (N_5120,N_350,N_8);
nor U5121 (N_5121,N_1656,N_2369);
nor U5122 (N_5122,N_1148,N_2279);
nand U5123 (N_5123,N_1816,N_1513);
or U5124 (N_5124,N_1175,N_1683);
or U5125 (N_5125,N_183,N_1826);
and U5126 (N_5126,N_2590,N_2240);
nand U5127 (N_5127,N_471,N_605);
nor U5128 (N_5128,N_1785,N_1459);
and U5129 (N_5129,N_1605,N_1449);
nand U5130 (N_5130,N_2708,N_1494);
and U5131 (N_5131,N_2190,N_344);
or U5132 (N_5132,N_1262,N_2497);
nand U5133 (N_5133,N_146,N_436);
and U5134 (N_5134,N_268,N_933);
nand U5135 (N_5135,N_2989,N_1161);
nand U5136 (N_5136,N_2670,N_260);
or U5137 (N_5137,N_2372,N_2974);
or U5138 (N_5138,N_981,N_2684);
or U5139 (N_5139,N_2665,N_196);
or U5140 (N_5140,N_2944,N_7);
and U5141 (N_5141,N_2503,N_1789);
nor U5142 (N_5142,N_630,N_1534);
and U5143 (N_5143,N_481,N_1889);
and U5144 (N_5144,N_50,N_78);
and U5145 (N_5145,N_1638,N_2877);
nand U5146 (N_5146,N_2046,N_47);
and U5147 (N_5147,N_1243,N_2880);
nor U5148 (N_5148,N_2561,N_1594);
nor U5149 (N_5149,N_1068,N_481);
and U5150 (N_5150,N_45,N_2040);
or U5151 (N_5151,N_969,N_2128);
nand U5152 (N_5152,N_2227,N_2437);
or U5153 (N_5153,N_240,N_1009);
xor U5154 (N_5154,N_468,N_2671);
or U5155 (N_5155,N_732,N_544);
or U5156 (N_5156,N_1577,N_1295);
nor U5157 (N_5157,N_1330,N_738);
or U5158 (N_5158,N_591,N_1809);
nor U5159 (N_5159,N_2394,N_2889);
and U5160 (N_5160,N_238,N_1966);
nor U5161 (N_5161,N_380,N_87);
or U5162 (N_5162,N_1009,N_2474);
and U5163 (N_5163,N_367,N_925);
or U5164 (N_5164,N_887,N_1240);
or U5165 (N_5165,N_2434,N_269);
nor U5166 (N_5166,N_345,N_988);
and U5167 (N_5167,N_1704,N_390);
and U5168 (N_5168,N_2761,N_1306);
nor U5169 (N_5169,N_2344,N_2588);
or U5170 (N_5170,N_416,N_2485);
nand U5171 (N_5171,N_32,N_2663);
nor U5172 (N_5172,N_2593,N_2745);
and U5173 (N_5173,N_2335,N_968);
and U5174 (N_5174,N_279,N_664);
and U5175 (N_5175,N_1188,N_672);
nand U5176 (N_5176,N_2374,N_1390);
and U5177 (N_5177,N_659,N_2328);
nor U5178 (N_5178,N_1488,N_2146);
and U5179 (N_5179,N_823,N_638);
nor U5180 (N_5180,N_1741,N_1347);
or U5181 (N_5181,N_2260,N_149);
xnor U5182 (N_5182,N_1324,N_361);
or U5183 (N_5183,N_2804,N_870);
or U5184 (N_5184,N_1415,N_2409);
and U5185 (N_5185,N_1978,N_1817);
xnor U5186 (N_5186,N_2475,N_396);
and U5187 (N_5187,N_82,N_2848);
nand U5188 (N_5188,N_1587,N_2896);
nand U5189 (N_5189,N_1718,N_2870);
nor U5190 (N_5190,N_1897,N_26);
and U5191 (N_5191,N_1956,N_766);
and U5192 (N_5192,N_1788,N_1719);
nand U5193 (N_5193,N_460,N_361);
nand U5194 (N_5194,N_1223,N_2165);
nor U5195 (N_5195,N_984,N_2692);
nor U5196 (N_5196,N_1523,N_2786);
nand U5197 (N_5197,N_419,N_702);
and U5198 (N_5198,N_1184,N_687);
nor U5199 (N_5199,N_1584,N_2089);
and U5200 (N_5200,N_1074,N_1128);
nor U5201 (N_5201,N_1711,N_2639);
and U5202 (N_5202,N_1959,N_1978);
nand U5203 (N_5203,N_1751,N_1780);
nor U5204 (N_5204,N_1041,N_2768);
nand U5205 (N_5205,N_2344,N_2672);
nor U5206 (N_5206,N_1770,N_1589);
nor U5207 (N_5207,N_1628,N_2952);
nand U5208 (N_5208,N_784,N_538);
nand U5209 (N_5209,N_2262,N_1673);
nand U5210 (N_5210,N_2133,N_2886);
nor U5211 (N_5211,N_1453,N_2183);
and U5212 (N_5212,N_1229,N_539);
and U5213 (N_5213,N_1403,N_479);
and U5214 (N_5214,N_2962,N_2174);
or U5215 (N_5215,N_2267,N_147);
or U5216 (N_5216,N_1963,N_2284);
and U5217 (N_5217,N_819,N_2065);
and U5218 (N_5218,N_500,N_2995);
or U5219 (N_5219,N_583,N_1682);
nor U5220 (N_5220,N_2445,N_2974);
nor U5221 (N_5221,N_95,N_174);
xnor U5222 (N_5222,N_2269,N_2340);
and U5223 (N_5223,N_2477,N_2744);
nor U5224 (N_5224,N_1448,N_2456);
nand U5225 (N_5225,N_1200,N_350);
or U5226 (N_5226,N_942,N_2729);
or U5227 (N_5227,N_1342,N_2632);
nand U5228 (N_5228,N_1575,N_2443);
or U5229 (N_5229,N_595,N_811);
and U5230 (N_5230,N_1721,N_756);
nand U5231 (N_5231,N_1764,N_1458);
nor U5232 (N_5232,N_2286,N_1840);
or U5233 (N_5233,N_599,N_325);
or U5234 (N_5234,N_2806,N_1557);
or U5235 (N_5235,N_2591,N_2419);
or U5236 (N_5236,N_2348,N_293);
nor U5237 (N_5237,N_616,N_2965);
nor U5238 (N_5238,N_454,N_269);
or U5239 (N_5239,N_1417,N_1971);
nand U5240 (N_5240,N_1220,N_1818);
and U5241 (N_5241,N_2906,N_779);
and U5242 (N_5242,N_87,N_2335);
or U5243 (N_5243,N_1135,N_2448);
nor U5244 (N_5244,N_604,N_87);
nand U5245 (N_5245,N_1144,N_493);
or U5246 (N_5246,N_1495,N_39);
nor U5247 (N_5247,N_376,N_2870);
and U5248 (N_5248,N_2280,N_2784);
or U5249 (N_5249,N_774,N_994);
and U5250 (N_5250,N_1820,N_1033);
or U5251 (N_5251,N_764,N_531);
or U5252 (N_5252,N_1993,N_2486);
and U5253 (N_5253,N_2705,N_860);
nor U5254 (N_5254,N_2301,N_1778);
nor U5255 (N_5255,N_2677,N_661);
nand U5256 (N_5256,N_1883,N_812);
and U5257 (N_5257,N_553,N_1841);
nor U5258 (N_5258,N_2818,N_2456);
or U5259 (N_5259,N_41,N_1827);
or U5260 (N_5260,N_1704,N_1051);
nand U5261 (N_5261,N_1736,N_2110);
and U5262 (N_5262,N_2531,N_584);
nand U5263 (N_5263,N_1723,N_2873);
or U5264 (N_5264,N_1721,N_819);
and U5265 (N_5265,N_1524,N_2962);
nand U5266 (N_5266,N_1505,N_1426);
and U5267 (N_5267,N_1340,N_175);
nor U5268 (N_5268,N_1687,N_2723);
nor U5269 (N_5269,N_859,N_1287);
and U5270 (N_5270,N_828,N_2929);
or U5271 (N_5271,N_308,N_1872);
nand U5272 (N_5272,N_2140,N_2450);
nand U5273 (N_5273,N_2457,N_2765);
or U5274 (N_5274,N_703,N_2236);
nand U5275 (N_5275,N_404,N_571);
or U5276 (N_5276,N_2766,N_245);
nand U5277 (N_5277,N_47,N_2670);
nor U5278 (N_5278,N_2580,N_1773);
or U5279 (N_5279,N_696,N_1337);
and U5280 (N_5280,N_323,N_338);
nand U5281 (N_5281,N_995,N_2713);
and U5282 (N_5282,N_1469,N_634);
and U5283 (N_5283,N_1539,N_883);
nor U5284 (N_5284,N_172,N_924);
or U5285 (N_5285,N_2353,N_229);
nand U5286 (N_5286,N_1286,N_93);
nor U5287 (N_5287,N_25,N_50);
or U5288 (N_5288,N_427,N_23);
or U5289 (N_5289,N_2960,N_1867);
nand U5290 (N_5290,N_706,N_1467);
nand U5291 (N_5291,N_1176,N_930);
nand U5292 (N_5292,N_1786,N_1618);
or U5293 (N_5293,N_711,N_1974);
nor U5294 (N_5294,N_686,N_1728);
nand U5295 (N_5295,N_1710,N_199);
nand U5296 (N_5296,N_2137,N_2978);
and U5297 (N_5297,N_2499,N_2798);
nor U5298 (N_5298,N_1469,N_1125);
nand U5299 (N_5299,N_1667,N_2393);
or U5300 (N_5300,N_286,N_686);
or U5301 (N_5301,N_1549,N_1744);
nand U5302 (N_5302,N_2456,N_1908);
nor U5303 (N_5303,N_2068,N_1211);
and U5304 (N_5304,N_601,N_2094);
and U5305 (N_5305,N_2227,N_1215);
and U5306 (N_5306,N_495,N_1649);
nor U5307 (N_5307,N_35,N_114);
nand U5308 (N_5308,N_558,N_842);
nand U5309 (N_5309,N_2243,N_2115);
and U5310 (N_5310,N_47,N_740);
and U5311 (N_5311,N_2264,N_375);
or U5312 (N_5312,N_1416,N_1237);
and U5313 (N_5313,N_2428,N_2032);
or U5314 (N_5314,N_649,N_947);
nand U5315 (N_5315,N_481,N_1811);
nand U5316 (N_5316,N_419,N_627);
or U5317 (N_5317,N_1098,N_2263);
and U5318 (N_5318,N_242,N_1740);
and U5319 (N_5319,N_2828,N_1097);
and U5320 (N_5320,N_237,N_2884);
nor U5321 (N_5321,N_2081,N_1585);
nand U5322 (N_5322,N_2383,N_2550);
and U5323 (N_5323,N_1136,N_2385);
nor U5324 (N_5324,N_1171,N_1769);
and U5325 (N_5325,N_2866,N_2300);
and U5326 (N_5326,N_1880,N_584);
or U5327 (N_5327,N_238,N_2514);
and U5328 (N_5328,N_2521,N_477);
nand U5329 (N_5329,N_2048,N_190);
nor U5330 (N_5330,N_2155,N_1954);
or U5331 (N_5331,N_2704,N_733);
nand U5332 (N_5332,N_1648,N_985);
and U5333 (N_5333,N_2214,N_2866);
nor U5334 (N_5334,N_60,N_577);
and U5335 (N_5335,N_221,N_1970);
nor U5336 (N_5336,N_2131,N_1684);
nand U5337 (N_5337,N_910,N_2770);
or U5338 (N_5338,N_1864,N_104);
or U5339 (N_5339,N_275,N_1829);
xor U5340 (N_5340,N_838,N_326);
nand U5341 (N_5341,N_1198,N_393);
or U5342 (N_5342,N_336,N_2956);
nor U5343 (N_5343,N_2031,N_1999);
and U5344 (N_5344,N_1096,N_188);
and U5345 (N_5345,N_645,N_1268);
nand U5346 (N_5346,N_680,N_881);
nor U5347 (N_5347,N_386,N_592);
or U5348 (N_5348,N_1635,N_255);
nand U5349 (N_5349,N_2395,N_2019);
or U5350 (N_5350,N_1639,N_632);
and U5351 (N_5351,N_1461,N_1227);
nand U5352 (N_5352,N_1803,N_2124);
and U5353 (N_5353,N_273,N_2047);
and U5354 (N_5354,N_1143,N_2654);
and U5355 (N_5355,N_2049,N_940);
and U5356 (N_5356,N_2958,N_1813);
or U5357 (N_5357,N_1972,N_767);
nand U5358 (N_5358,N_601,N_874);
nor U5359 (N_5359,N_961,N_463);
and U5360 (N_5360,N_2892,N_72);
nand U5361 (N_5361,N_2688,N_764);
nor U5362 (N_5362,N_986,N_1513);
and U5363 (N_5363,N_2288,N_2366);
and U5364 (N_5364,N_2006,N_2650);
nand U5365 (N_5365,N_2234,N_944);
and U5366 (N_5366,N_1391,N_1992);
nor U5367 (N_5367,N_1370,N_1733);
nand U5368 (N_5368,N_1591,N_1570);
or U5369 (N_5369,N_1978,N_928);
xnor U5370 (N_5370,N_2631,N_2530);
and U5371 (N_5371,N_2006,N_1569);
and U5372 (N_5372,N_135,N_537);
nand U5373 (N_5373,N_2970,N_382);
nor U5374 (N_5374,N_1927,N_2174);
and U5375 (N_5375,N_1177,N_1536);
or U5376 (N_5376,N_801,N_2848);
nand U5377 (N_5377,N_219,N_1007);
or U5378 (N_5378,N_2084,N_1227);
nor U5379 (N_5379,N_2178,N_1207);
nor U5380 (N_5380,N_853,N_2913);
and U5381 (N_5381,N_520,N_637);
or U5382 (N_5382,N_616,N_627);
nor U5383 (N_5383,N_575,N_807);
and U5384 (N_5384,N_733,N_434);
and U5385 (N_5385,N_1546,N_2212);
and U5386 (N_5386,N_1634,N_1742);
and U5387 (N_5387,N_2236,N_897);
and U5388 (N_5388,N_2897,N_756);
or U5389 (N_5389,N_1838,N_1970);
and U5390 (N_5390,N_2886,N_704);
nand U5391 (N_5391,N_216,N_83);
or U5392 (N_5392,N_1839,N_2322);
and U5393 (N_5393,N_613,N_2313);
or U5394 (N_5394,N_2606,N_249);
or U5395 (N_5395,N_1093,N_1681);
or U5396 (N_5396,N_145,N_1771);
nor U5397 (N_5397,N_812,N_1727);
xor U5398 (N_5398,N_321,N_1051);
and U5399 (N_5399,N_207,N_683);
nor U5400 (N_5400,N_1331,N_233);
or U5401 (N_5401,N_2171,N_2773);
and U5402 (N_5402,N_2795,N_102);
and U5403 (N_5403,N_1463,N_626);
or U5404 (N_5404,N_2377,N_1704);
nor U5405 (N_5405,N_1390,N_602);
or U5406 (N_5406,N_775,N_348);
or U5407 (N_5407,N_2944,N_2463);
and U5408 (N_5408,N_299,N_735);
or U5409 (N_5409,N_1695,N_2726);
and U5410 (N_5410,N_2275,N_426);
or U5411 (N_5411,N_2913,N_1667);
and U5412 (N_5412,N_2620,N_1582);
and U5413 (N_5413,N_1186,N_2459);
or U5414 (N_5414,N_695,N_779);
and U5415 (N_5415,N_2153,N_2054);
and U5416 (N_5416,N_205,N_2304);
and U5417 (N_5417,N_2340,N_1857);
and U5418 (N_5418,N_588,N_1735);
and U5419 (N_5419,N_2395,N_1515);
and U5420 (N_5420,N_2001,N_1140);
and U5421 (N_5421,N_988,N_2496);
nand U5422 (N_5422,N_346,N_1584);
and U5423 (N_5423,N_1731,N_1596);
or U5424 (N_5424,N_85,N_2961);
nor U5425 (N_5425,N_2986,N_2939);
or U5426 (N_5426,N_1374,N_280);
or U5427 (N_5427,N_2599,N_2933);
or U5428 (N_5428,N_1947,N_2305);
nand U5429 (N_5429,N_939,N_892);
or U5430 (N_5430,N_551,N_2703);
nor U5431 (N_5431,N_1468,N_2740);
or U5432 (N_5432,N_2533,N_2263);
xor U5433 (N_5433,N_2025,N_767);
nand U5434 (N_5434,N_1225,N_1502);
xnor U5435 (N_5435,N_699,N_1947);
or U5436 (N_5436,N_33,N_2198);
and U5437 (N_5437,N_873,N_1366);
nand U5438 (N_5438,N_1517,N_910);
or U5439 (N_5439,N_1291,N_147);
or U5440 (N_5440,N_219,N_2667);
nand U5441 (N_5441,N_1647,N_2343);
or U5442 (N_5442,N_2609,N_440);
or U5443 (N_5443,N_832,N_1923);
and U5444 (N_5444,N_1805,N_2626);
or U5445 (N_5445,N_277,N_493);
nor U5446 (N_5446,N_1098,N_2885);
or U5447 (N_5447,N_2025,N_421);
nor U5448 (N_5448,N_1301,N_2452);
nand U5449 (N_5449,N_2944,N_1492);
nor U5450 (N_5450,N_1855,N_2045);
nand U5451 (N_5451,N_1143,N_413);
nor U5452 (N_5452,N_2216,N_510);
or U5453 (N_5453,N_321,N_785);
nand U5454 (N_5454,N_2543,N_827);
or U5455 (N_5455,N_1196,N_1528);
and U5456 (N_5456,N_1385,N_2423);
nand U5457 (N_5457,N_1916,N_2867);
nor U5458 (N_5458,N_2651,N_1210);
and U5459 (N_5459,N_2959,N_1671);
and U5460 (N_5460,N_174,N_1321);
nor U5461 (N_5461,N_2676,N_2312);
or U5462 (N_5462,N_556,N_1313);
nor U5463 (N_5463,N_1604,N_119);
nor U5464 (N_5464,N_1879,N_456);
nand U5465 (N_5465,N_2569,N_1165);
or U5466 (N_5466,N_2524,N_1464);
and U5467 (N_5467,N_1926,N_87);
nor U5468 (N_5468,N_1658,N_1810);
nand U5469 (N_5469,N_1689,N_1681);
and U5470 (N_5470,N_146,N_1390);
nand U5471 (N_5471,N_140,N_2836);
or U5472 (N_5472,N_105,N_2871);
nor U5473 (N_5473,N_2302,N_684);
nand U5474 (N_5474,N_515,N_821);
or U5475 (N_5475,N_2385,N_808);
and U5476 (N_5476,N_22,N_1961);
and U5477 (N_5477,N_1233,N_2450);
nand U5478 (N_5478,N_939,N_1182);
or U5479 (N_5479,N_276,N_1678);
nand U5480 (N_5480,N_2716,N_2258);
nand U5481 (N_5481,N_1347,N_1211);
nand U5482 (N_5482,N_2245,N_1087);
nand U5483 (N_5483,N_1632,N_1098);
nor U5484 (N_5484,N_1405,N_1116);
nand U5485 (N_5485,N_314,N_502);
and U5486 (N_5486,N_2126,N_1588);
and U5487 (N_5487,N_2447,N_809);
nand U5488 (N_5488,N_2364,N_301);
nand U5489 (N_5489,N_2767,N_8);
or U5490 (N_5490,N_2143,N_2876);
nand U5491 (N_5491,N_2815,N_362);
and U5492 (N_5492,N_1533,N_2374);
nand U5493 (N_5493,N_2496,N_1044);
and U5494 (N_5494,N_1070,N_1392);
or U5495 (N_5495,N_302,N_2208);
nand U5496 (N_5496,N_1346,N_652);
nand U5497 (N_5497,N_1374,N_1565);
and U5498 (N_5498,N_993,N_461);
and U5499 (N_5499,N_1320,N_614);
and U5500 (N_5500,N_764,N_1417);
nor U5501 (N_5501,N_1771,N_806);
or U5502 (N_5502,N_515,N_1312);
or U5503 (N_5503,N_2987,N_1580);
nand U5504 (N_5504,N_1574,N_174);
nand U5505 (N_5505,N_1390,N_1387);
and U5506 (N_5506,N_1206,N_1340);
nand U5507 (N_5507,N_2330,N_2704);
nand U5508 (N_5508,N_883,N_936);
nor U5509 (N_5509,N_468,N_2248);
nand U5510 (N_5510,N_2412,N_654);
or U5511 (N_5511,N_1383,N_467);
and U5512 (N_5512,N_2994,N_1082);
and U5513 (N_5513,N_790,N_1566);
nor U5514 (N_5514,N_253,N_1601);
nor U5515 (N_5515,N_2831,N_2502);
nand U5516 (N_5516,N_402,N_256);
nand U5517 (N_5517,N_2378,N_1599);
and U5518 (N_5518,N_2972,N_450);
and U5519 (N_5519,N_2405,N_2051);
or U5520 (N_5520,N_2129,N_1421);
nor U5521 (N_5521,N_2593,N_833);
or U5522 (N_5522,N_2327,N_1948);
nand U5523 (N_5523,N_2543,N_986);
nand U5524 (N_5524,N_2728,N_1358);
nand U5525 (N_5525,N_1517,N_946);
or U5526 (N_5526,N_2021,N_2936);
nand U5527 (N_5527,N_1116,N_2002);
nor U5528 (N_5528,N_45,N_1253);
or U5529 (N_5529,N_707,N_1375);
or U5530 (N_5530,N_2454,N_291);
nor U5531 (N_5531,N_599,N_824);
and U5532 (N_5532,N_943,N_667);
or U5533 (N_5533,N_478,N_235);
and U5534 (N_5534,N_1488,N_113);
nor U5535 (N_5535,N_823,N_730);
and U5536 (N_5536,N_2354,N_398);
nand U5537 (N_5537,N_1875,N_1838);
nor U5538 (N_5538,N_172,N_1809);
and U5539 (N_5539,N_2192,N_1731);
nor U5540 (N_5540,N_2705,N_2861);
nand U5541 (N_5541,N_778,N_1254);
or U5542 (N_5542,N_149,N_2392);
nor U5543 (N_5543,N_1500,N_1831);
or U5544 (N_5544,N_1721,N_2774);
and U5545 (N_5545,N_2875,N_1904);
nor U5546 (N_5546,N_914,N_51);
nor U5547 (N_5547,N_417,N_618);
nand U5548 (N_5548,N_2602,N_1434);
and U5549 (N_5549,N_2271,N_188);
nand U5550 (N_5550,N_935,N_2080);
nand U5551 (N_5551,N_2442,N_1122);
nor U5552 (N_5552,N_1490,N_239);
nand U5553 (N_5553,N_2392,N_2568);
and U5554 (N_5554,N_2372,N_811);
or U5555 (N_5555,N_214,N_1618);
and U5556 (N_5556,N_438,N_2093);
or U5557 (N_5557,N_551,N_247);
nand U5558 (N_5558,N_2384,N_2292);
nand U5559 (N_5559,N_700,N_2029);
or U5560 (N_5560,N_1794,N_6);
nor U5561 (N_5561,N_100,N_2163);
and U5562 (N_5562,N_669,N_636);
nand U5563 (N_5563,N_2137,N_2300);
xnor U5564 (N_5564,N_2274,N_2518);
nand U5565 (N_5565,N_433,N_46);
and U5566 (N_5566,N_1240,N_168);
nor U5567 (N_5567,N_1099,N_2620);
and U5568 (N_5568,N_970,N_420);
and U5569 (N_5569,N_652,N_416);
and U5570 (N_5570,N_788,N_1786);
or U5571 (N_5571,N_2974,N_2331);
nor U5572 (N_5572,N_2163,N_335);
or U5573 (N_5573,N_2545,N_799);
or U5574 (N_5574,N_745,N_980);
or U5575 (N_5575,N_857,N_231);
and U5576 (N_5576,N_136,N_2059);
nand U5577 (N_5577,N_2189,N_2337);
nor U5578 (N_5578,N_1357,N_1278);
nand U5579 (N_5579,N_975,N_824);
nand U5580 (N_5580,N_319,N_1228);
or U5581 (N_5581,N_1207,N_139);
nor U5582 (N_5582,N_1119,N_1000);
nor U5583 (N_5583,N_1003,N_1941);
nand U5584 (N_5584,N_2824,N_1105);
nand U5585 (N_5585,N_1578,N_280);
nor U5586 (N_5586,N_1614,N_273);
and U5587 (N_5587,N_274,N_1113);
nand U5588 (N_5588,N_538,N_720);
and U5589 (N_5589,N_266,N_1019);
and U5590 (N_5590,N_617,N_2882);
and U5591 (N_5591,N_2281,N_430);
nor U5592 (N_5592,N_354,N_157);
or U5593 (N_5593,N_146,N_1514);
or U5594 (N_5594,N_1555,N_2942);
nand U5595 (N_5595,N_1405,N_2267);
nand U5596 (N_5596,N_2458,N_1910);
nand U5597 (N_5597,N_1702,N_2997);
nand U5598 (N_5598,N_522,N_2834);
or U5599 (N_5599,N_2470,N_2800);
nand U5600 (N_5600,N_125,N_867);
and U5601 (N_5601,N_249,N_82);
and U5602 (N_5602,N_618,N_1352);
and U5603 (N_5603,N_4,N_236);
or U5604 (N_5604,N_1153,N_904);
nor U5605 (N_5605,N_160,N_2178);
and U5606 (N_5606,N_2683,N_2646);
or U5607 (N_5607,N_2713,N_339);
or U5608 (N_5608,N_2914,N_1132);
or U5609 (N_5609,N_199,N_2009);
nor U5610 (N_5610,N_2588,N_1155);
nand U5611 (N_5611,N_2630,N_2350);
nand U5612 (N_5612,N_458,N_1393);
nand U5613 (N_5613,N_2548,N_2777);
nand U5614 (N_5614,N_631,N_520);
nor U5615 (N_5615,N_1685,N_754);
or U5616 (N_5616,N_342,N_1992);
or U5617 (N_5617,N_2470,N_638);
nor U5618 (N_5618,N_1863,N_974);
and U5619 (N_5619,N_676,N_1638);
or U5620 (N_5620,N_2722,N_2949);
nor U5621 (N_5621,N_2315,N_2952);
and U5622 (N_5622,N_1015,N_1899);
nor U5623 (N_5623,N_352,N_1380);
or U5624 (N_5624,N_1212,N_1941);
or U5625 (N_5625,N_1495,N_67);
and U5626 (N_5626,N_1676,N_794);
or U5627 (N_5627,N_956,N_555);
nor U5628 (N_5628,N_2548,N_351);
nor U5629 (N_5629,N_2413,N_603);
nand U5630 (N_5630,N_821,N_158);
nor U5631 (N_5631,N_958,N_1505);
and U5632 (N_5632,N_460,N_2315);
nor U5633 (N_5633,N_2072,N_42);
or U5634 (N_5634,N_1581,N_2046);
nand U5635 (N_5635,N_1609,N_175);
nand U5636 (N_5636,N_1611,N_1959);
nor U5637 (N_5637,N_2119,N_752);
and U5638 (N_5638,N_1581,N_615);
nand U5639 (N_5639,N_520,N_669);
nand U5640 (N_5640,N_199,N_525);
nand U5641 (N_5641,N_2319,N_724);
or U5642 (N_5642,N_854,N_1878);
and U5643 (N_5643,N_2836,N_133);
nor U5644 (N_5644,N_2918,N_640);
nor U5645 (N_5645,N_51,N_2893);
and U5646 (N_5646,N_537,N_1915);
nor U5647 (N_5647,N_407,N_2692);
nor U5648 (N_5648,N_1577,N_815);
nor U5649 (N_5649,N_2636,N_1719);
nand U5650 (N_5650,N_1418,N_200);
nor U5651 (N_5651,N_1100,N_2156);
nand U5652 (N_5652,N_1749,N_2172);
or U5653 (N_5653,N_2011,N_1268);
nand U5654 (N_5654,N_865,N_527);
nor U5655 (N_5655,N_2350,N_1025);
nand U5656 (N_5656,N_2430,N_2074);
and U5657 (N_5657,N_1871,N_1517);
nor U5658 (N_5658,N_1984,N_1109);
nand U5659 (N_5659,N_2411,N_344);
nor U5660 (N_5660,N_1216,N_2827);
and U5661 (N_5661,N_670,N_826);
or U5662 (N_5662,N_971,N_673);
nand U5663 (N_5663,N_1127,N_1944);
or U5664 (N_5664,N_1409,N_2862);
or U5665 (N_5665,N_556,N_2044);
nand U5666 (N_5666,N_943,N_2711);
nor U5667 (N_5667,N_2780,N_2113);
nand U5668 (N_5668,N_490,N_1355);
or U5669 (N_5669,N_1080,N_1236);
and U5670 (N_5670,N_373,N_1952);
nand U5671 (N_5671,N_132,N_2790);
and U5672 (N_5672,N_217,N_2994);
or U5673 (N_5673,N_142,N_1805);
or U5674 (N_5674,N_2876,N_2665);
or U5675 (N_5675,N_2570,N_698);
nand U5676 (N_5676,N_2381,N_2781);
and U5677 (N_5677,N_641,N_154);
and U5678 (N_5678,N_1062,N_1765);
or U5679 (N_5679,N_1353,N_1049);
nand U5680 (N_5680,N_1870,N_894);
or U5681 (N_5681,N_393,N_2403);
or U5682 (N_5682,N_1598,N_521);
nand U5683 (N_5683,N_368,N_844);
or U5684 (N_5684,N_892,N_419);
nor U5685 (N_5685,N_844,N_1636);
nor U5686 (N_5686,N_1243,N_2383);
or U5687 (N_5687,N_1026,N_267);
or U5688 (N_5688,N_963,N_1218);
nor U5689 (N_5689,N_583,N_2167);
and U5690 (N_5690,N_1001,N_1840);
or U5691 (N_5691,N_2098,N_2231);
or U5692 (N_5692,N_2126,N_50);
or U5693 (N_5693,N_2996,N_1130);
nand U5694 (N_5694,N_729,N_1860);
or U5695 (N_5695,N_1057,N_609);
nor U5696 (N_5696,N_367,N_181);
nand U5697 (N_5697,N_2588,N_75);
nand U5698 (N_5698,N_860,N_286);
nand U5699 (N_5699,N_1761,N_2567);
or U5700 (N_5700,N_383,N_1723);
nand U5701 (N_5701,N_2335,N_510);
nor U5702 (N_5702,N_2052,N_2292);
or U5703 (N_5703,N_1705,N_516);
nand U5704 (N_5704,N_2707,N_2364);
nand U5705 (N_5705,N_983,N_931);
nand U5706 (N_5706,N_2822,N_2073);
and U5707 (N_5707,N_2515,N_1710);
or U5708 (N_5708,N_2780,N_2888);
and U5709 (N_5709,N_2598,N_2076);
or U5710 (N_5710,N_2232,N_2881);
nor U5711 (N_5711,N_2985,N_2347);
or U5712 (N_5712,N_1734,N_2869);
nor U5713 (N_5713,N_1595,N_1452);
or U5714 (N_5714,N_2767,N_2294);
or U5715 (N_5715,N_1294,N_1887);
and U5716 (N_5716,N_2565,N_2399);
nand U5717 (N_5717,N_2443,N_2743);
or U5718 (N_5718,N_1638,N_2966);
or U5719 (N_5719,N_1506,N_1615);
nor U5720 (N_5720,N_2670,N_778);
nor U5721 (N_5721,N_22,N_1175);
or U5722 (N_5722,N_1561,N_1248);
nor U5723 (N_5723,N_1188,N_1749);
nor U5724 (N_5724,N_2351,N_35);
nand U5725 (N_5725,N_960,N_1109);
nor U5726 (N_5726,N_1709,N_641);
nand U5727 (N_5727,N_461,N_713);
and U5728 (N_5728,N_99,N_764);
nand U5729 (N_5729,N_60,N_1255);
nor U5730 (N_5730,N_1988,N_1099);
nand U5731 (N_5731,N_791,N_2358);
nor U5732 (N_5732,N_1810,N_61);
nor U5733 (N_5733,N_548,N_2372);
nor U5734 (N_5734,N_740,N_1225);
or U5735 (N_5735,N_1094,N_1744);
and U5736 (N_5736,N_2468,N_352);
and U5737 (N_5737,N_1998,N_932);
nor U5738 (N_5738,N_2109,N_53);
nor U5739 (N_5739,N_1950,N_1847);
and U5740 (N_5740,N_2278,N_2170);
and U5741 (N_5741,N_1177,N_850);
and U5742 (N_5742,N_1972,N_746);
and U5743 (N_5743,N_2394,N_1224);
nor U5744 (N_5744,N_1807,N_700);
nand U5745 (N_5745,N_1970,N_749);
or U5746 (N_5746,N_579,N_1394);
nand U5747 (N_5747,N_2328,N_863);
or U5748 (N_5748,N_2954,N_397);
xor U5749 (N_5749,N_780,N_173);
nor U5750 (N_5750,N_1169,N_974);
nand U5751 (N_5751,N_691,N_499);
and U5752 (N_5752,N_1608,N_1171);
nand U5753 (N_5753,N_2024,N_2367);
or U5754 (N_5754,N_592,N_1043);
and U5755 (N_5755,N_1816,N_1045);
and U5756 (N_5756,N_2668,N_570);
or U5757 (N_5757,N_1210,N_2984);
nor U5758 (N_5758,N_2603,N_803);
nor U5759 (N_5759,N_613,N_1368);
or U5760 (N_5760,N_2722,N_2424);
nand U5761 (N_5761,N_2677,N_1219);
or U5762 (N_5762,N_2241,N_390);
and U5763 (N_5763,N_2966,N_1563);
and U5764 (N_5764,N_1947,N_923);
nor U5765 (N_5765,N_2302,N_2588);
nand U5766 (N_5766,N_2522,N_2109);
nand U5767 (N_5767,N_2819,N_344);
nor U5768 (N_5768,N_2406,N_1916);
nand U5769 (N_5769,N_706,N_1367);
nand U5770 (N_5770,N_53,N_2403);
or U5771 (N_5771,N_367,N_378);
or U5772 (N_5772,N_2262,N_1335);
nor U5773 (N_5773,N_1566,N_2450);
or U5774 (N_5774,N_959,N_1938);
and U5775 (N_5775,N_612,N_1181);
nor U5776 (N_5776,N_1623,N_2272);
nand U5777 (N_5777,N_1790,N_588);
nor U5778 (N_5778,N_1336,N_97);
nand U5779 (N_5779,N_2520,N_2793);
nor U5780 (N_5780,N_2824,N_2963);
nand U5781 (N_5781,N_1115,N_1066);
nor U5782 (N_5782,N_2266,N_1600);
nand U5783 (N_5783,N_1035,N_1656);
nor U5784 (N_5784,N_162,N_2284);
or U5785 (N_5785,N_879,N_2449);
nand U5786 (N_5786,N_2037,N_2702);
nor U5787 (N_5787,N_2162,N_67);
nand U5788 (N_5788,N_1614,N_2192);
nor U5789 (N_5789,N_870,N_1639);
or U5790 (N_5790,N_2545,N_675);
and U5791 (N_5791,N_941,N_418);
nand U5792 (N_5792,N_1604,N_1194);
nand U5793 (N_5793,N_2599,N_2630);
nand U5794 (N_5794,N_458,N_2346);
nand U5795 (N_5795,N_1194,N_2016);
and U5796 (N_5796,N_2647,N_2617);
nor U5797 (N_5797,N_408,N_1220);
nor U5798 (N_5798,N_2140,N_1299);
nor U5799 (N_5799,N_409,N_708);
nor U5800 (N_5800,N_783,N_123);
nor U5801 (N_5801,N_1946,N_1117);
nand U5802 (N_5802,N_1389,N_504);
nand U5803 (N_5803,N_1613,N_1954);
or U5804 (N_5804,N_2104,N_472);
nand U5805 (N_5805,N_2199,N_2504);
nor U5806 (N_5806,N_2888,N_574);
or U5807 (N_5807,N_1495,N_856);
nand U5808 (N_5808,N_2282,N_1033);
nor U5809 (N_5809,N_1821,N_209);
or U5810 (N_5810,N_850,N_23);
and U5811 (N_5811,N_861,N_781);
or U5812 (N_5812,N_1112,N_2389);
and U5813 (N_5813,N_456,N_2450);
nor U5814 (N_5814,N_2755,N_2180);
nand U5815 (N_5815,N_1482,N_2033);
and U5816 (N_5816,N_2417,N_558);
and U5817 (N_5817,N_453,N_465);
nor U5818 (N_5818,N_1789,N_2487);
or U5819 (N_5819,N_2347,N_2799);
nor U5820 (N_5820,N_1075,N_2533);
nand U5821 (N_5821,N_2804,N_651);
nor U5822 (N_5822,N_2640,N_1015);
nor U5823 (N_5823,N_1189,N_112);
nand U5824 (N_5824,N_586,N_2753);
and U5825 (N_5825,N_1944,N_1006);
nor U5826 (N_5826,N_183,N_536);
nand U5827 (N_5827,N_805,N_922);
or U5828 (N_5828,N_2947,N_1068);
nand U5829 (N_5829,N_1546,N_2838);
and U5830 (N_5830,N_2743,N_2351);
and U5831 (N_5831,N_2598,N_812);
and U5832 (N_5832,N_2379,N_680);
and U5833 (N_5833,N_511,N_912);
nor U5834 (N_5834,N_2865,N_2353);
or U5835 (N_5835,N_1153,N_1541);
or U5836 (N_5836,N_1101,N_1237);
nand U5837 (N_5837,N_341,N_2269);
nand U5838 (N_5838,N_476,N_1035);
xor U5839 (N_5839,N_2690,N_819);
and U5840 (N_5840,N_24,N_182);
and U5841 (N_5841,N_622,N_662);
nand U5842 (N_5842,N_282,N_524);
nand U5843 (N_5843,N_2733,N_228);
nand U5844 (N_5844,N_470,N_831);
nor U5845 (N_5845,N_553,N_910);
and U5846 (N_5846,N_1685,N_2396);
nor U5847 (N_5847,N_1799,N_2811);
nor U5848 (N_5848,N_564,N_1148);
nor U5849 (N_5849,N_841,N_568);
and U5850 (N_5850,N_1373,N_1622);
and U5851 (N_5851,N_521,N_2432);
or U5852 (N_5852,N_973,N_2651);
and U5853 (N_5853,N_1253,N_1254);
nor U5854 (N_5854,N_2234,N_1193);
nor U5855 (N_5855,N_2405,N_1668);
nand U5856 (N_5856,N_2424,N_238);
or U5857 (N_5857,N_1470,N_2503);
nand U5858 (N_5858,N_1611,N_2009);
and U5859 (N_5859,N_2582,N_1342);
or U5860 (N_5860,N_82,N_1823);
nand U5861 (N_5861,N_415,N_148);
and U5862 (N_5862,N_1007,N_2829);
nor U5863 (N_5863,N_211,N_1880);
and U5864 (N_5864,N_235,N_2168);
and U5865 (N_5865,N_2847,N_2739);
nor U5866 (N_5866,N_2831,N_461);
nor U5867 (N_5867,N_1220,N_1930);
nand U5868 (N_5868,N_2068,N_544);
nor U5869 (N_5869,N_751,N_220);
nor U5870 (N_5870,N_2138,N_360);
or U5871 (N_5871,N_2715,N_101);
nor U5872 (N_5872,N_2328,N_2001);
or U5873 (N_5873,N_360,N_2469);
nor U5874 (N_5874,N_1811,N_1751);
or U5875 (N_5875,N_2347,N_427);
nor U5876 (N_5876,N_18,N_2295);
nor U5877 (N_5877,N_1507,N_166);
or U5878 (N_5878,N_1629,N_1341);
or U5879 (N_5879,N_1652,N_148);
and U5880 (N_5880,N_1059,N_2243);
or U5881 (N_5881,N_1342,N_680);
nor U5882 (N_5882,N_2733,N_2830);
nand U5883 (N_5883,N_1143,N_2968);
or U5884 (N_5884,N_2849,N_2491);
nand U5885 (N_5885,N_471,N_2088);
nor U5886 (N_5886,N_1376,N_2919);
or U5887 (N_5887,N_194,N_2885);
or U5888 (N_5888,N_1518,N_1853);
and U5889 (N_5889,N_2759,N_262);
or U5890 (N_5890,N_2398,N_277);
and U5891 (N_5891,N_2578,N_133);
or U5892 (N_5892,N_408,N_2859);
or U5893 (N_5893,N_2787,N_2218);
nor U5894 (N_5894,N_2543,N_2430);
nand U5895 (N_5895,N_2275,N_126);
nand U5896 (N_5896,N_685,N_2618);
nand U5897 (N_5897,N_1271,N_2827);
nand U5898 (N_5898,N_206,N_1762);
xor U5899 (N_5899,N_2613,N_2506);
xor U5900 (N_5900,N_2844,N_430);
nand U5901 (N_5901,N_1454,N_357);
nor U5902 (N_5902,N_32,N_947);
and U5903 (N_5903,N_2928,N_1677);
or U5904 (N_5904,N_510,N_1216);
or U5905 (N_5905,N_1150,N_222);
nand U5906 (N_5906,N_1053,N_488);
and U5907 (N_5907,N_2533,N_2414);
nand U5908 (N_5908,N_2741,N_2803);
nor U5909 (N_5909,N_1836,N_2970);
and U5910 (N_5910,N_2241,N_805);
nor U5911 (N_5911,N_2404,N_1059);
nor U5912 (N_5912,N_1635,N_293);
nor U5913 (N_5913,N_696,N_795);
or U5914 (N_5914,N_2801,N_641);
and U5915 (N_5915,N_712,N_1399);
nor U5916 (N_5916,N_1636,N_231);
and U5917 (N_5917,N_2135,N_144);
nand U5918 (N_5918,N_2116,N_922);
nor U5919 (N_5919,N_2333,N_1699);
or U5920 (N_5920,N_2201,N_2343);
nor U5921 (N_5921,N_1726,N_481);
nand U5922 (N_5922,N_933,N_759);
nor U5923 (N_5923,N_2558,N_1765);
nand U5924 (N_5924,N_2582,N_2848);
or U5925 (N_5925,N_609,N_217);
or U5926 (N_5926,N_165,N_363);
nor U5927 (N_5927,N_1282,N_655);
nand U5928 (N_5928,N_2395,N_2828);
or U5929 (N_5929,N_1901,N_1090);
and U5930 (N_5930,N_584,N_2916);
nand U5931 (N_5931,N_1995,N_705);
and U5932 (N_5932,N_91,N_2855);
nor U5933 (N_5933,N_1957,N_1713);
or U5934 (N_5934,N_867,N_2559);
nor U5935 (N_5935,N_1787,N_417);
and U5936 (N_5936,N_850,N_1110);
nand U5937 (N_5937,N_624,N_2967);
or U5938 (N_5938,N_2895,N_2267);
or U5939 (N_5939,N_2816,N_128);
nor U5940 (N_5940,N_1678,N_2814);
nand U5941 (N_5941,N_1863,N_1731);
nor U5942 (N_5942,N_2291,N_1316);
or U5943 (N_5943,N_407,N_2255);
or U5944 (N_5944,N_1961,N_151);
or U5945 (N_5945,N_736,N_797);
or U5946 (N_5946,N_1628,N_2406);
or U5947 (N_5947,N_2481,N_2374);
or U5948 (N_5948,N_1838,N_2017);
and U5949 (N_5949,N_2288,N_2794);
and U5950 (N_5950,N_1436,N_1039);
or U5951 (N_5951,N_2113,N_1917);
nand U5952 (N_5952,N_2492,N_2196);
nand U5953 (N_5953,N_1220,N_1190);
nor U5954 (N_5954,N_1349,N_2919);
nor U5955 (N_5955,N_594,N_2688);
and U5956 (N_5956,N_917,N_1873);
or U5957 (N_5957,N_1789,N_2803);
nand U5958 (N_5958,N_1092,N_124);
and U5959 (N_5959,N_199,N_298);
nand U5960 (N_5960,N_1557,N_1714);
nor U5961 (N_5961,N_547,N_1214);
and U5962 (N_5962,N_403,N_2388);
and U5963 (N_5963,N_616,N_2194);
nand U5964 (N_5964,N_2213,N_2091);
or U5965 (N_5965,N_1795,N_1315);
and U5966 (N_5966,N_2490,N_1067);
nand U5967 (N_5967,N_985,N_1353);
nor U5968 (N_5968,N_454,N_1784);
nor U5969 (N_5969,N_1457,N_987);
and U5970 (N_5970,N_2134,N_416);
nor U5971 (N_5971,N_2983,N_1693);
nor U5972 (N_5972,N_1381,N_2954);
nor U5973 (N_5973,N_551,N_925);
or U5974 (N_5974,N_665,N_1797);
nand U5975 (N_5975,N_2048,N_986);
and U5976 (N_5976,N_1348,N_2579);
nand U5977 (N_5977,N_2497,N_2869);
or U5978 (N_5978,N_2077,N_194);
or U5979 (N_5979,N_887,N_1534);
or U5980 (N_5980,N_2266,N_2682);
or U5981 (N_5981,N_1555,N_2303);
nand U5982 (N_5982,N_661,N_465);
and U5983 (N_5983,N_1641,N_2333);
nor U5984 (N_5984,N_44,N_2240);
or U5985 (N_5985,N_1437,N_1075);
and U5986 (N_5986,N_1655,N_1943);
or U5987 (N_5987,N_1862,N_2638);
nor U5988 (N_5988,N_1102,N_757);
nor U5989 (N_5989,N_2974,N_2082);
and U5990 (N_5990,N_2376,N_1369);
or U5991 (N_5991,N_2675,N_2624);
nor U5992 (N_5992,N_1840,N_67);
and U5993 (N_5993,N_2991,N_584);
nor U5994 (N_5994,N_234,N_1025);
and U5995 (N_5995,N_1141,N_327);
or U5996 (N_5996,N_2569,N_910);
or U5997 (N_5997,N_2882,N_346);
nor U5998 (N_5998,N_2897,N_1219);
nand U5999 (N_5999,N_2414,N_797);
nand U6000 (N_6000,N_5764,N_3529);
and U6001 (N_6001,N_4087,N_5322);
nand U6002 (N_6002,N_4821,N_4398);
and U6003 (N_6003,N_4996,N_3411);
nand U6004 (N_6004,N_4740,N_5330);
nor U6005 (N_6005,N_5631,N_5678);
or U6006 (N_6006,N_3104,N_5347);
nor U6007 (N_6007,N_5189,N_3454);
and U6008 (N_6008,N_4635,N_4409);
and U6009 (N_6009,N_5407,N_4864);
and U6010 (N_6010,N_4437,N_3913);
and U6011 (N_6011,N_3910,N_5188);
nand U6012 (N_6012,N_4460,N_4036);
or U6013 (N_6013,N_4482,N_3685);
nor U6014 (N_6014,N_3260,N_4678);
nand U6015 (N_6015,N_3281,N_3124);
or U6016 (N_6016,N_5969,N_4534);
or U6017 (N_6017,N_4797,N_5450);
nor U6018 (N_6018,N_3163,N_3423);
nand U6019 (N_6019,N_3049,N_5873);
or U6020 (N_6020,N_3984,N_3036);
or U6021 (N_6021,N_5492,N_3594);
or U6022 (N_6022,N_3439,N_5504);
and U6023 (N_6023,N_3224,N_3363);
or U6024 (N_6024,N_5232,N_4410);
nor U6025 (N_6025,N_4074,N_3034);
and U6026 (N_6026,N_4549,N_4433);
or U6027 (N_6027,N_5650,N_5657);
nand U6028 (N_6028,N_3221,N_5518);
nor U6029 (N_6029,N_3120,N_3237);
nor U6030 (N_6030,N_3409,N_4747);
or U6031 (N_6031,N_4965,N_4824);
and U6032 (N_6032,N_3185,N_5253);
or U6033 (N_6033,N_5823,N_4538);
or U6034 (N_6034,N_3442,N_5173);
nor U6035 (N_6035,N_5515,N_5001);
nor U6036 (N_6036,N_5222,N_3259);
and U6037 (N_6037,N_5441,N_3089);
nand U6038 (N_6038,N_3231,N_4761);
nor U6039 (N_6039,N_4639,N_4187);
or U6040 (N_6040,N_3515,N_3177);
and U6041 (N_6041,N_5763,N_4464);
nand U6042 (N_6042,N_3417,N_5096);
and U6043 (N_6043,N_3256,N_3161);
or U6044 (N_6044,N_4853,N_3450);
or U6045 (N_6045,N_5342,N_5206);
nand U6046 (N_6046,N_3894,N_5185);
nand U6047 (N_6047,N_4512,N_3004);
and U6048 (N_6048,N_5731,N_3751);
or U6049 (N_6049,N_5896,N_4123);
or U6050 (N_6050,N_5017,N_4939);
nor U6051 (N_6051,N_3655,N_5652);
nor U6052 (N_6052,N_5385,N_4583);
or U6053 (N_6053,N_3262,N_5457);
or U6054 (N_6054,N_3844,N_5554);
or U6055 (N_6055,N_4271,N_3957);
or U6056 (N_6056,N_4387,N_5511);
nand U6057 (N_6057,N_3056,N_5961);
nand U6058 (N_6058,N_4714,N_5449);
nor U6059 (N_6059,N_5295,N_4364);
nand U6060 (N_6060,N_4155,N_5230);
or U6061 (N_6061,N_4990,N_3097);
nor U6062 (N_6062,N_4057,N_5806);
and U6063 (N_6063,N_4945,N_4816);
nor U6064 (N_6064,N_3550,N_3123);
nand U6065 (N_6065,N_3987,N_5828);
and U6066 (N_6066,N_4934,N_4967);
nand U6067 (N_6067,N_5054,N_4624);
and U6068 (N_6068,N_5890,N_4008);
nor U6069 (N_6069,N_5831,N_4120);
and U6070 (N_6070,N_3863,N_4017);
or U6071 (N_6071,N_4535,N_3369);
or U6072 (N_6072,N_4484,N_3634);
nand U6073 (N_6073,N_5036,N_3760);
or U6074 (N_6074,N_4633,N_3646);
nor U6075 (N_6075,N_4210,N_3179);
or U6076 (N_6076,N_4431,N_4694);
or U6077 (N_6077,N_5509,N_5061);
nor U6078 (N_6078,N_4589,N_3452);
nor U6079 (N_6079,N_4318,N_4357);
and U6080 (N_6080,N_3683,N_4901);
and U6081 (N_6081,N_4929,N_5703);
nand U6082 (N_6082,N_3448,N_3145);
and U6083 (N_6083,N_5181,N_5577);
nand U6084 (N_6084,N_3579,N_5746);
and U6085 (N_6085,N_4041,N_4831);
and U6086 (N_6086,N_4661,N_4006);
and U6087 (N_6087,N_3168,N_5847);
nor U6088 (N_6088,N_3003,N_5599);
nand U6089 (N_6089,N_5924,N_3821);
and U6090 (N_6090,N_4707,N_5335);
or U6091 (N_6091,N_4869,N_5947);
nand U6092 (N_6092,N_3695,N_5639);
nand U6093 (N_6093,N_5562,N_4013);
nand U6094 (N_6094,N_3122,N_5312);
nor U6095 (N_6095,N_5648,N_5462);
and U6096 (N_6096,N_5803,N_4923);
and U6097 (N_6097,N_5461,N_5986);
nand U6098 (N_6098,N_3756,N_4776);
or U6099 (N_6099,N_3228,N_5794);
nor U6100 (N_6100,N_4018,N_3016);
and U6101 (N_6101,N_3178,N_4362);
or U6102 (N_6102,N_3410,N_3412);
nand U6103 (N_6103,N_5760,N_3075);
xnor U6104 (N_6104,N_3549,N_5276);
nor U6105 (N_6105,N_4937,N_4973);
and U6106 (N_6106,N_4880,N_3284);
and U6107 (N_6107,N_3286,N_4803);
nor U6108 (N_6108,N_4345,N_4098);
and U6109 (N_6109,N_5358,N_5557);
nand U6110 (N_6110,N_3400,N_4446);
and U6111 (N_6111,N_5008,N_3767);
nor U6112 (N_6112,N_4314,N_5150);
nor U6113 (N_6113,N_4019,N_5713);
nand U6114 (N_6114,N_4257,N_5854);
nand U6115 (N_6115,N_3880,N_5762);
nand U6116 (N_6116,N_5796,N_4618);
nand U6117 (N_6117,N_5499,N_3545);
and U6118 (N_6118,N_5395,N_4039);
or U6119 (N_6119,N_3496,N_5184);
and U6120 (N_6120,N_5260,N_3017);
nand U6121 (N_6121,N_4420,N_5651);
nand U6122 (N_6122,N_5418,N_5507);
and U6123 (N_6123,N_4980,N_4605);
nor U6124 (N_6124,N_4672,N_4554);
nor U6125 (N_6125,N_4327,N_4266);
nor U6126 (N_6126,N_3297,N_5098);
nor U6127 (N_6127,N_5741,N_4978);
nand U6128 (N_6128,N_5003,N_4664);
nor U6129 (N_6129,N_3257,N_4994);
nor U6130 (N_6130,N_4473,N_3864);
or U6131 (N_6131,N_3473,N_5560);
nor U6132 (N_6132,N_3798,N_5078);
nor U6133 (N_6133,N_5567,N_5467);
or U6134 (N_6134,N_3506,N_4703);
and U6135 (N_6135,N_4432,N_4375);
or U6136 (N_6136,N_3861,N_4686);
nor U6137 (N_6137,N_4366,N_5367);
nor U6138 (N_6138,N_5275,N_3159);
or U6139 (N_6139,N_5235,N_5944);
nor U6140 (N_6140,N_5332,N_4692);
nand U6141 (N_6141,N_4843,N_3934);
nand U6142 (N_6142,N_4477,N_4156);
and U6143 (N_6143,N_4405,N_5549);
nor U6144 (N_6144,N_4680,N_5878);
or U6145 (N_6145,N_4283,N_5673);
and U6146 (N_6146,N_4290,N_4564);
or U6147 (N_6147,N_4877,N_3770);
or U6148 (N_6148,N_3765,N_3740);
or U6149 (N_6149,N_5965,N_3626);
nor U6150 (N_6150,N_5880,N_5616);
nor U6151 (N_6151,N_4977,N_4617);
nand U6152 (N_6152,N_5212,N_5959);
nand U6153 (N_6153,N_5815,N_4706);
or U6154 (N_6154,N_4365,N_3640);
nor U6155 (N_6155,N_3132,N_5900);
nand U6156 (N_6156,N_3951,N_4455);
and U6157 (N_6157,N_5442,N_5667);
or U6158 (N_6158,N_4891,N_4146);
or U6159 (N_6159,N_4374,N_3703);
nand U6160 (N_6160,N_3681,N_4842);
or U6161 (N_6161,N_3062,N_4778);
nor U6162 (N_6162,N_3952,N_5963);
and U6163 (N_6163,N_5301,N_5066);
or U6164 (N_6164,N_4817,N_3280);
and U6165 (N_6165,N_3437,N_3697);
and U6166 (N_6166,N_5836,N_4453);
or U6167 (N_6167,N_4768,N_3607);
nand U6168 (N_6168,N_4058,N_4599);
and U6169 (N_6169,N_5738,N_5294);
or U6170 (N_6170,N_3255,N_4563);
or U6171 (N_6171,N_3108,N_4259);
and U6172 (N_6172,N_4935,N_3873);
nor U6173 (N_6173,N_4157,N_3074);
and U6174 (N_6174,N_5566,N_4304);
or U6175 (N_6175,N_5151,N_3544);
nand U6176 (N_6176,N_5153,N_3380);
and U6177 (N_6177,N_5886,N_3464);
or U6178 (N_6178,N_3040,N_5257);
nand U6179 (N_6179,N_3782,N_3136);
nand U6180 (N_6180,N_4269,N_3253);
nor U6181 (N_6181,N_5174,N_5936);
and U6182 (N_6182,N_3193,N_5500);
nor U6183 (N_6183,N_4732,N_4721);
nand U6184 (N_6184,N_5808,N_3476);
nand U6185 (N_6185,N_4650,N_5086);
nor U6186 (N_6186,N_5272,N_3785);
and U6187 (N_6187,N_4083,N_3250);
nand U6188 (N_6188,N_4104,N_4527);
nor U6189 (N_6189,N_5106,N_3650);
and U6190 (N_6190,N_3725,N_5879);
nor U6191 (N_6191,N_3229,N_4284);
nor U6192 (N_6192,N_3384,N_4874);
nor U6193 (N_6193,N_4401,N_4506);
nand U6194 (N_6194,N_3541,N_5131);
nor U6195 (N_6195,N_5946,N_4625);
nand U6196 (N_6196,N_4117,N_3467);
nor U6197 (N_6197,N_4495,N_5339);
or U6198 (N_6198,N_3605,N_4829);
or U6199 (N_6199,N_4430,N_3086);
and U6200 (N_6200,N_4636,N_5705);
or U6201 (N_6201,N_5041,N_3942);
or U6202 (N_6202,N_5000,N_3451);
or U6203 (N_6203,N_3890,N_5708);
and U6204 (N_6204,N_3436,N_3668);
or U6205 (N_6205,N_3649,N_4794);
nor U6206 (N_6206,N_4666,N_3225);
or U6207 (N_6207,N_3245,N_4397);
or U6208 (N_6208,N_3326,N_4812);
or U6209 (N_6209,N_3938,N_3282);
or U6210 (N_6210,N_5446,N_4199);
nor U6211 (N_6211,N_3689,N_3706);
nand U6212 (N_6212,N_5026,N_5242);
nor U6213 (N_6213,N_3519,N_4790);
and U6214 (N_6214,N_5364,N_4807);
and U6215 (N_6215,N_4360,N_4815);
and U6216 (N_6216,N_4823,N_4465);
and U6217 (N_6217,N_5775,N_3446);
nand U6218 (N_6218,N_3335,N_5215);
nor U6219 (N_6219,N_5956,N_5812);
nand U6220 (N_6220,N_4010,N_4785);
nor U6221 (N_6221,N_5659,N_4548);
or U6222 (N_6222,N_5234,N_5618);
or U6223 (N_6223,N_5785,N_3666);
and U6224 (N_6224,N_5976,N_4808);
or U6225 (N_6225,N_4687,N_5470);
nor U6226 (N_6226,N_4338,N_4236);
or U6227 (N_6227,N_3109,N_3390);
nand U6228 (N_6228,N_3818,N_3370);
or U6229 (N_6229,N_4905,N_5454);
or U6230 (N_6230,N_5917,N_3311);
nor U6231 (N_6231,N_5998,N_3275);
and U6232 (N_6232,N_5758,N_3285);
and U6233 (N_6233,N_3994,N_5093);
nand U6234 (N_6234,N_3797,N_5541);
nor U6235 (N_6235,N_3386,N_4903);
or U6236 (N_6236,N_5084,N_4412);
and U6237 (N_6237,N_4863,N_4195);
nor U6238 (N_6238,N_5002,N_4134);
and U6239 (N_6239,N_4508,N_5702);
and U6240 (N_6240,N_5736,N_4885);
nor U6241 (N_6241,N_5837,N_5352);
and U6242 (N_6242,N_4591,N_3560);
nor U6243 (N_6243,N_4987,N_5570);
or U6244 (N_6244,N_4164,N_3927);
nor U6245 (N_6245,N_4066,N_4498);
nor U6246 (N_6246,N_3637,N_3199);
and U6247 (N_6247,N_5876,N_3632);
nor U6248 (N_6248,N_5020,N_4059);
or U6249 (N_6249,N_5075,N_3595);
nor U6250 (N_6250,N_3340,N_5074);
nor U6251 (N_6251,N_4470,N_5829);
nor U6252 (N_6252,N_3848,N_4644);
and U6253 (N_6253,N_3498,N_3043);
nor U6254 (N_6254,N_4281,N_4056);
nor U6255 (N_6255,N_3548,N_3585);
and U6256 (N_6256,N_3433,N_5588);
nand U6257 (N_6257,N_3947,N_4393);
or U6258 (N_6258,N_5038,N_5076);
and U6259 (N_6259,N_5997,N_5130);
or U6260 (N_6260,N_4648,N_4321);
or U6261 (N_6261,N_4168,N_5704);
nor U6262 (N_6262,N_5291,N_5505);
nand U6263 (N_6263,N_4674,N_4016);
nand U6264 (N_6264,N_3713,N_5196);
nand U6265 (N_6265,N_4716,N_5519);
nor U6266 (N_6266,N_5714,N_4485);
nor U6267 (N_6267,N_4069,N_4933);
and U6268 (N_6268,N_5843,N_3542);
nor U6269 (N_6269,N_5563,N_5568);
or U6270 (N_6270,N_4324,N_3916);
xor U6271 (N_6271,N_4627,N_5425);
and U6272 (N_6272,N_3966,N_3528);
nor U6273 (N_6273,N_3094,N_4161);
or U6274 (N_6274,N_5191,N_5887);
nor U6275 (N_6275,N_4913,N_5428);
nand U6276 (N_6276,N_4342,N_5412);
and U6277 (N_6277,N_5533,N_3879);
or U6278 (N_6278,N_5695,N_3222);
nand U6279 (N_6279,N_5574,N_5376);
nor U6280 (N_6280,N_5217,N_4029);
nand U6281 (N_6281,N_4334,N_3035);
or U6282 (N_6282,N_5220,N_4337);
and U6283 (N_6283,N_3232,N_5875);
and U6284 (N_6284,N_5902,N_3206);
nor U6285 (N_6285,N_4382,N_3757);
nor U6286 (N_6286,N_3847,N_4184);
or U6287 (N_6287,N_5360,N_5256);
nand U6288 (N_6288,N_4102,N_4297);
and U6289 (N_6289,N_5857,N_4385);
nor U6290 (N_6290,N_5553,N_3458);
or U6291 (N_6291,N_4407,N_4969);
nand U6292 (N_6292,N_4542,N_5872);
and U6293 (N_6293,N_5589,N_5045);
and U6294 (N_6294,N_4400,N_5643);
or U6295 (N_6295,N_3569,N_4784);
and U6296 (N_6296,N_3465,N_5813);
nand U6297 (N_6297,N_4094,N_4277);
nor U6298 (N_6298,N_5473,N_5298);
or U6299 (N_6299,N_3432,N_3126);
xor U6300 (N_6300,N_3708,N_5278);
and U6301 (N_6301,N_5409,N_4766);
nor U6302 (N_6302,N_5940,N_3376);
and U6303 (N_6303,N_5202,N_3647);
and U6304 (N_6304,N_5680,N_5400);
nand U6305 (N_6305,N_5124,N_5465);
or U6306 (N_6306,N_4704,N_3907);
nand U6307 (N_6307,N_5996,N_3096);
nor U6308 (N_6308,N_5942,N_5883);
nor U6309 (N_6309,N_3771,N_4368);
or U6310 (N_6310,N_4450,N_4001);
nand U6311 (N_6311,N_4504,N_5517);
nand U6312 (N_6312,N_5089,N_3902);
and U6313 (N_6313,N_5635,N_5907);
or U6314 (N_6314,N_3719,N_5158);
or U6315 (N_6315,N_5608,N_5377);
and U6316 (N_6316,N_3868,N_5314);
and U6317 (N_6317,N_4819,N_4752);
or U6318 (N_6318,N_5120,N_5968);
and U6319 (N_6319,N_3928,N_5555);
nor U6320 (N_6320,N_3213,N_4558);
nand U6321 (N_6321,N_5982,N_3616);
or U6322 (N_6322,N_4129,N_4964);
or U6323 (N_6323,N_4580,N_4662);
nor U6324 (N_6324,N_3012,N_3813);
or U6325 (N_6325,N_5417,N_5233);
and U6326 (N_6326,N_4909,N_3730);
nor U6327 (N_6327,N_4571,N_4352);
or U6328 (N_6328,N_4938,N_5934);
or U6329 (N_6329,N_5710,N_3825);
nand U6330 (N_6330,N_4839,N_4291);
or U6331 (N_6331,N_5595,N_5072);
or U6332 (N_6332,N_4501,N_5030);
and U6333 (N_6333,N_5779,N_4031);
nand U6334 (N_6334,N_4852,N_5179);
or U6335 (N_6335,N_4867,N_4331);
nor U6336 (N_6336,N_5083,N_3128);
and U6337 (N_6337,N_3332,N_4739);
nor U6338 (N_6338,N_5593,N_5814);
nor U6339 (N_6339,N_5810,N_3182);
or U6340 (N_6340,N_5022,N_3742);
and U6341 (N_6341,N_3835,N_3112);
and U6342 (N_6342,N_4030,N_4423);
nand U6343 (N_6343,N_4806,N_5707);
and U6344 (N_6344,N_3693,N_3053);
nand U6345 (N_6345,N_4649,N_5621);
and U6346 (N_6346,N_4045,N_4858);
nor U6347 (N_6347,N_3667,N_3329);
and U6348 (N_6348,N_5378,N_3396);
and U6349 (N_6349,N_4932,N_5929);
nand U6350 (N_6350,N_5670,N_3198);
nand U6351 (N_6351,N_3025,N_3597);
nand U6352 (N_6352,N_4562,N_5063);
nand U6353 (N_6353,N_4051,N_3032);
nor U6354 (N_6354,N_5157,N_4668);
and U6355 (N_6355,N_5954,N_4026);
nor U6356 (N_6356,N_5576,N_4724);
nor U6357 (N_6357,N_5204,N_3274);
or U6358 (N_6358,N_5899,N_4669);
and U6359 (N_6359,N_3731,N_5190);
and U6360 (N_6360,N_4521,N_5610);
and U6361 (N_6361,N_4457,N_3009);
and U6362 (N_6362,N_3155,N_3728);
nand U6363 (N_6363,N_4246,N_5308);
or U6364 (N_6364,N_3299,N_4526);
nand U6365 (N_6365,N_5712,N_4490);
or U6366 (N_6366,N_4065,N_3917);
nand U6367 (N_6367,N_4763,N_4388);
nor U6368 (N_6368,N_3866,N_5754);
and U6369 (N_6369,N_4596,N_5460);
or U6370 (N_6370,N_5405,N_3775);
and U6371 (N_6371,N_3642,N_3618);
or U6372 (N_6372,N_5751,N_4762);
xor U6373 (N_6373,N_4267,N_5060);
or U6374 (N_6374,N_3787,N_4751);
nand U6375 (N_6375,N_3055,N_3582);
or U6376 (N_6376,N_5723,N_5226);
nor U6377 (N_6377,N_3111,N_5481);
or U6378 (N_6378,N_5720,N_5326);
or U6379 (N_6379,N_3098,N_3978);
nor U6380 (N_6380,N_4151,N_3300);
and U6381 (N_6381,N_4536,N_4109);
and U6382 (N_6382,N_4944,N_5247);
nor U6383 (N_6383,N_4876,N_3022);
or U6384 (N_6384,N_4466,N_4590);
or U6385 (N_6385,N_4735,N_3461);
nand U6386 (N_6386,N_5102,N_5134);
nand U6387 (N_6387,N_3977,N_5172);
nor U6388 (N_6388,N_3258,N_4711);
nand U6389 (N_6389,N_5641,N_3580);
nand U6390 (N_6390,N_4875,N_4261);
and U6391 (N_6391,N_3444,N_4836);
nor U6392 (N_6392,N_5908,N_3871);
and U6393 (N_6393,N_3325,N_5118);
or U6394 (N_6394,N_3659,N_5937);
or U6395 (N_6395,N_4294,N_3462);
nor U6396 (N_6396,N_3744,N_3202);
and U6397 (N_6397,N_4174,N_3853);
nor U6398 (N_6398,N_3865,N_3276);
nand U6399 (N_6399,N_5099,N_4171);
nor U6400 (N_6400,N_5088,N_3147);
nor U6401 (N_6401,N_5085,N_5716);
or U6402 (N_6402,N_3870,N_5672);
nor U6403 (N_6403,N_3581,N_3944);
or U6404 (N_6404,N_4456,N_3242);
nand U6405 (N_6405,N_5208,N_5349);
and U6406 (N_6406,N_4856,N_4924);
nor U6407 (N_6407,N_4197,N_5456);
nand U6408 (N_6408,N_4308,N_5218);
or U6409 (N_6409,N_4982,N_3521);
or U6410 (N_6410,N_3324,N_3567);
and U6411 (N_6411,N_3427,N_5306);
nand U6412 (N_6412,N_5480,N_4500);
and U6413 (N_6413,N_3536,N_4336);
nand U6414 (N_6414,N_3323,N_3071);
and U6415 (N_6415,N_4434,N_4305);
or U6416 (N_6416,N_5299,N_4683);
and U6417 (N_6417,N_3188,N_5682);
nand U6418 (N_6418,N_5438,N_3261);
or U6419 (N_6419,N_3302,N_3008);
and U6420 (N_6420,N_5144,N_4774);
nand U6421 (N_6421,N_5095,N_4320);
nor U6422 (N_6422,N_4959,N_4299);
or U6423 (N_6423,N_5201,N_4767);
and U6424 (N_6424,N_4167,N_4855);
nand U6425 (N_6425,N_5628,N_4175);
or U6426 (N_6426,N_5444,N_4182);
nand U6427 (N_6427,N_4093,N_3013);
and U6428 (N_6428,N_3830,N_4073);
and U6429 (N_6429,N_3696,N_5973);
nor U6430 (N_6430,N_3244,N_3503);
or U6431 (N_6431,N_5279,N_4658);
and U6432 (N_6432,N_4404,N_4519);
nand U6433 (N_6433,N_4615,N_5477);
nor U6434 (N_6434,N_4573,N_4791);
nand U6435 (N_6435,N_5696,N_3172);
nand U6436 (N_6436,N_3252,N_4176);
nor U6437 (N_6437,N_5646,N_4894);
and U6438 (N_6438,N_4381,N_5503);
and U6439 (N_6439,N_3981,N_4077);
or U6440 (N_6440,N_3500,N_5155);
nand U6441 (N_6441,N_3677,N_4531);
nand U6442 (N_6442,N_3558,N_3230);
or U6443 (N_6443,N_4921,N_5065);
and U6444 (N_6444,N_3362,N_4274);
nand U6445 (N_6445,N_5726,N_5354);
or U6446 (N_6446,N_5080,N_5901);
nor U6447 (N_6447,N_4848,N_4022);
nand U6448 (N_6448,N_3010,N_4135);
or U6449 (N_6449,N_5512,N_5214);
nor U6450 (N_6450,N_3641,N_3754);
nor U6451 (N_6451,N_3307,N_4601);
nand U6452 (N_6452,N_3645,N_5992);
and U6453 (N_6453,N_4961,N_5437);
nand U6454 (N_6454,N_3078,N_5759);
or U6455 (N_6455,N_5647,N_4023);
or U6456 (N_6456,N_4701,N_5368);
and U6457 (N_6457,N_5203,N_3779);
or U6458 (N_6458,N_5501,N_5478);
or U6459 (N_6459,N_5104,N_5868);
or U6460 (N_6460,N_5849,N_4015);
and U6461 (N_6461,N_4753,N_3090);
nor U6462 (N_6462,N_5375,N_3290);
and U6463 (N_6463,N_5394,N_4421);
nand U6464 (N_6464,N_5655,N_4480);
nand U6465 (N_6465,N_4847,N_5320);
or U6466 (N_6466,N_4020,N_3812);
nor U6467 (N_6467,N_4966,N_4062);
and U6468 (N_6468,N_3915,N_3184);
nor U6469 (N_6469,N_3763,N_3234);
nand U6470 (N_6470,N_5977,N_3316);
nor U6471 (N_6471,N_4827,N_5784);
nand U6472 (N_6472,N_5420,N_4553);
and U6473 (N_6473,N_5129,N_5615);
or U6474 (N_6474,N_5127,N_4656);
xor U6475 (N_6475,N_3148,N_3463);
or U6476 (N_6476,N_4780,N_4238);
or U6477 (N_6477,N_5825,N_5141);
and U6478 (N_6478,N_4225,N_4377);
nand U6479 (N_6479,N_3872,N_5891);
and U6480 (N_6480,N_3627,N_4193);
nand U6481 (N_6481,N_5029,N_4286);
nor U6482 (N_6482,N_3425,N_3336);
or U6483 (N_6483,N_5472,N_4745);
nand U6484 (N_6484,N_4252,N_3709);
and U6485 (N_6485,N_3174,N_3313);
nor U6486 (N_6486,N_4702,N_4798);
nand U6487 (N_6487,N_5846,N_4042);
nand U6488 (N_6488,N_5033,N_3710);
nor U6489 (N_6489,N_3832,N_4516);
nand U6490 (N_6490,N_4585,N_5573);
and U6491 (N_6491,N_5734,N_5110);
nor U6492 (N_6492,N_4483,N_4219);
nor U6493 (N_6493,N_5152,N_4486);
nor U6494 (N_6494,N_4064,N_5448);
and U6495 (N_6495,N_5431,N_5550);
nand U6496 (N_6496,N_4429,N_5336);
or U6497 (N_6497,N_3557,N_4092);
nand U6498 (N_6498,N_5370,N_5858);
nand U6499 (N_6499,N_3364,N_4699);
nand U6500 (N_6500,N_5081,N_5869);
nand U6501 (N_6501,N_5371,N_5390);
nor U6502 (N_6502,N_5042,N_5459);
nand U6503 (N_6503,N_3941,N_5665);
or U6504 (N_6504,N_3974,N_5522);
or U6505 (N_6505,N_4781,N_3048);
and U6506 (N_6506,N_4414,N_5451);
and U6507 (N_6507,N_5693,N_3900);
nand U6508 (N_6508,N_4837,N_3073);
or U6509 (N_6509,N_4832,N_3110);
or U6510 (N_6510,N_4032,N_5258);
nand U6511 (N_6511,N_5778,N_5051);
and U6512 (N_6512,N_4640,N_3959);
nand U6513 (N_6513,N_3737,N_5458);
and U6514 (N_6514,N_4152,N_4142);
and U6515 (N_6515,N_4425,N_3602);
nand U6516 (N_6516,N_3125,N_3114);
or U6517 (N_6517,N_3615,N_3753);
or U6518 (N_6518,N_3998,N_3733);
nor U6519 (N_6519,N_5584,N_5388);
or U6520 (N_6520,N_3183,N_4068);
nand U6521 (N_6521,N_3217,N_3682);
nand U6522 (N_6522,N_3804,N_4502);
nor U6523 (N_6523,N_5197,N_4356);
and U6524 (N_6524,N_5591,N_4796);
nor U6525 (N_6525,N_4492,N_4116);
or U6526 (N_6526,N_4946,N_5408);
nor U6527 (N_6527,N_4612,N_4613);
nor U6528 (N_6528,N_3429,N_3546);
and U6529 (N_6529,N_5911,N_4777);
or U6530 (N_6530,N_3963,N_3639);
xor U6531 (N_6531,N_3064,N_3679);
or U6532 (N_6532,N_5495,N_3854);
nor U6533 (N_6533,N_3648,N_4424);
or U6534 (N_6534,N_3418,N_4954);
nand U6535 (N_6535,N_3317,N_3511);
or U6536 (N_6536,N_4124,N_5565);
nand U6537 (N_6537,N_5750,N_5935);
nor U6538 (N_6538,N_3227,N_3822);
or U6539 (N_6539,N_4879,N_3516);
and U6540 (N_6540,N_5090,N_5701);
nand U6541 (N_6541,N_4955,N_3819);
nand U6542 (N_6542,N_3748,N_3794);
or U6543 (N_6543,N_4113,N_4488);
and U6544 (N_6544,N_4750,N_4147);
or U6545 (N_6545,N_3065,N_3971);
nor U6546 (N_6546,N_4902,N_3901);
and U6547 (N_6547,N_4137,N_5819);
and U6548 (N_6548,N_4295,N_4332);
or U6549 (N_6549,N_5633,N_3115);
nor U6550 (N_6550,N_4629,N_5135);
nand U6551 (N_6551,N_4086,N_4481);
nand U6552 (N_6552,N_4908,N_3932);
nand U6553 (N_6553,N_5547,N_5592);
or U6554 (N_6554,N_3976,N_5874);
and U6555 (N_6555,N_3191,N_3475);
nand U6556 (N_6556,N_5387,N_3070);
nand U6557 (N_6557,N_5856,N_5993);
nand U6558 (N_6558,N_5194,N_4713);
or U6559 (N_6559,N_4850,N_4361);
and U6560 (N_6560,N_4244,N_4126);
and U6561 (N_6561,N_4559,N_5686);
or U6562 (N_6562,N_5816,N_3576);
and U6563 (N_6563,N_4606,N_4201);
and U6564 (N_6564,N_5548,N_3428);
or U6565 (N_6565,N_3956,N_5004);
nand U6566 (N_6566,N_5694,N_3216);
nor U6567 (N_6567,N_3711,N_4216);
and U6568 (N_6568,N_4520,N_4044);
nor U6569 (N_6569,N_3077,N_5386);
and U6570 (N_6570,N_4872,N_3834);
nor U6571 (N_6571,N_4415,N_3958);
nand U6572 (N_6572,N_3486,N_3360);
nand U6573 (N_6573,N_3377,N_4667);
and U6574 (N_6574,N_3195,N_3658);
and U6575 (N_6575,N_4103,N_5748);
or U6576 (N_6576,N_4577,N_3815);
or U6577 (N_6577,N_3330,N_5483);
nor U6578 (N_6578,N_4467,N_5266);
or U6579 (N_6579,N_5945,N_5424);
nor U6580 (N_6580,N_5912,N_5293);
or U6581 (N_6581,N_5538,N_4054);
or U6582 (N_6582,N_4826,N_4021);
nand U6583 (N_6583,N_3403,N_3273);
nor U6584 (N_6584,N_5398,N_4204);
or U6585 (N_6585,N_4632,N_5283);
and U6586 (N_6586,N_5043,N_4458);
nor U6587 (N_6587,N_4811,N_3718);
nand U6588 (N_6588,N_4943,N_4154);
nor U6589 (N_6589,N_3746,N_4474);
and U6590 (N_6590,N_5379,N_5116);
and U6591 (N_6591,N_4422,N_5485);
nor U6592 (N_6592,N_3887,N_4461);
xor U6593 (N_6593,N_4651,N_5073);
nand U6594 (N_6594,N_4048,N_4543);
xor U6595 (N_6595,N_3024,N_3395);
and U6596 (N_6596,N_3153,N_4951);
and U6597 (N_6597,N_3762,N_5287);
and U6598 (N_6598,N_5769,N_3026);
nor U6599 (N_6599,N_3678,N_3497);
or U6600 (N_6600,N_5684,N_4411);
and U6601 (N_6601,N_3367,N_5761);
or U6602 (N_6602,N_5537,N_3562);
or U6603 (N_6603,N_5572,N_3298);
or U6604 (N_6604,N_4545,N_4917);
nor U6605 (N_6605,N_3823,N_5310);
or U6606 (N_6606,N_5820,N_3383);
nor U6607 (N_6607,N_3249,N_4950);
or U6608 (N_6608,N_5801,N_4726);
or U6609 (N_6609,N_5315,N_3385);
nand U6610 (N_6610,N_4801,N_4084);
and U6611 (N_6611,N_5730,N_4028);
or U6612 (N_6612,N_3724,N_4660);
or U6613 (N_6613,N_3657,N_5559);
and U6614 (N_6614,N_5489,N_3263);
xor U6615 (N_6615,N_3800,N_3493);
nor U6616 (N_6616,N_5288,N_3768);
nor U6617 (N_6617,N_4111,N_5864);
nand U6618 (N_6618,N_5988,N_3365);
and U6619 (N_6619,N_5068,N_3449);
nand U6620 (N_6620,N_5679,N_4524);
or U6621 (N_6621,N_5575,N_3858);
or U6622 (N_6622,N_3144,N_5776);
xnor U6623 (N_6623,N_5343,N_4922);
and U6624 (N_6624,N_5049,N_3614);
nand U6625 (N_6625,N_3979,N_3989);
nor U6626 (N_6626,N_5248,N_4183);
and U6627 (N_6627,N_5318,N_4264);
nand U6628 (N_6628,N_3479,N_3272);
nand U6629 (N_6629,N_4024,N_5502);
or U6630 (N_6630,N_5596,N_5255);
or U6631 (N_6631,N_5105,N_4597);
and U6632 (N_6632,N_5161,N_3522);
and U6633 (N_6633,N_3653,N_5906);
nor U6634 (N_6634,N_4655,N_3993);
and U6635 (N_6635,N_3769,N_4000);
nor U6636 (N_6636,N_4251,N_4213);
and U6637 (N_6637,N_5263,N_3911);
or U6638 (N_6638,N_5848,N_4670);
nor U6639 (N_6639,N_5578,N_3714);
and U6640 (N_6640,N_4301,N_5156);
and U6641 (N_6641,N_3404,N_3780);
nand U6642 (N_6642,N_3573,N_4034);
nand U6643 (N_6643,N_5587,N_5966);
nor U6644 (N_6644,N_3431,N_4158);
nand U6645 (N_6645,N_3574,N_3398);
nor U6646 (N_6646,N_4828,N_4335);
nor U6647 (N_6647,N_4359,N_3914);
nor U6648 (N_6648,N_4047,N_3173);
or U6649 (N_6649,N_3707,N_4565);
nor U6650 (N_6650,N_5267,N_4800);
and U6651 (N_6651,N_4110,N_5822);
nand U6652 (N_6652,N_4638,N_3334);
and U6653 (N_6653,N_5254,N_4127);
nand U6654 (N_6654,N_4159,N_3063);
nand U6655 (N_6655,N_5677,N_4186);
or U6656 (N_6656,N_3793,N_3129);
and U6657 (N_6657,N_3208,N_5359);
or U6658 (N_6658,N_4718,N_3029);
nand U6659 (N_6659,N_5292,N_4859);
nand U6660 (N_6660,N_3867,N_5674);
nor U6661 (N_6661,N_4988,N_5178);
or U6662 (N_6662,N_4734,N_4416);
or U6663 (N_6663,N_3954,N_3200);
and U6664 (N_6664,N_5251,N_5926);
or U6665 (N_6665,N_3100,N_4475);
and U6666 (N_6666,N_5133,N_4581);
or U6667 (N_6667,N_4118,N_4514);
nor U6668 (N_6668,N_3061,N_4265);
and U6669 (N_6669,N_3106,N_4188);
nand U6670 (N_6670,N_4695,N_3160);
nor U6671 (N_6671,N_3338,N_4673);
and U6672 (N_6672,N_3883,N_3684);
nand U6673 (N_6673,N_5170,N_3068);
and U6674 (N_6674,N_5623,N_4802);
nor U6675 (N_6675,N_5097,N_3239);
nand U6676 (N_6676,N_5241,N_4203);
and U6677 (N_6677,N_5013,N_5689);
and U6678 (N_6678,N_4380,N_3388);
and U6679 (N_6679,N_5216,N_5432);
nand U6680 (N_6680,N_5752,N_4749);
nand U6681 (N_6681,N_3936,N_3885);
nor U6682 (N_6682,N_3505,N_3392);
nor U6683 (N_6683,N_3859,N_4786);
nor U6684 (N_6684,N_5951,N_3482);
or U6685 (N_6685,N_5122,N_4717);
or U6686 (N_6686,N_5316,N_3672);
and U6687 (N_6687,N_5307,N_4814);
nand U6688 (N_6688,N_4315,N_5916);
and U6689 (N_6689,N_3165,N_4106);
nor U6690 (N_6690,N_4497,N_5619);
or U6691 (N_6691,N_4227,N_4743);
nand U6692 (N_6692,N_5171,N_5077);
nand U6693 (N_6693,N_3831,N_5744);
or U6694 (N_6694,N_3824,N_3490);
and U6695 (N_6695,N_4956,N_3162);
nor U6696 (N_6696,N_5913,N_3350);
or U6697 (N_6697,N_3838,N_5540);
or U6698 (N_6698,N_5606,N_5137);
nor U6699 (N_6699,N_3922,N_5668);
nand U6700 (N_6700,N_4963,N_5669);
or U6701 (N_6701,N_3038,N_5627);
nor U6702 (N_6702,N_4510,N_4438);
or U6703 (N_6703,N_4268,N_4725);
and U6704 (N_6704,N_3196,N_5274);
nor U6705 (N_6705,N_4447,N_5757);
and U6706 (N_6706,N_3551,N_5035);
nand U6707 (N_6707,N_5632,N_3170);
nand U6708 (N_6708,N_5108,N_4080);
and U6709 (N_6709,N_3547,N_5807);
nor U6710 (N_6710,N_5938,N_4805);
and U6711 (N_6711,N_5798,N_5827);
nand U6712 (N_6712,N_3152,N_3149);
nor U6713 (N_6713,N_5115,N_3309);
nor U6714 (N_6714,N_5010,N_3306);
nor U6715 (N_6715,N_5044,N_3485);
or U6716 (N_6716,N_3139,N_3884);
or U6717 (N_6717,N_3248,N_5192);
nor U6718 (N_6718,N_4962,N_3201);
or U6719 (N_6719,N_3294,N_3720);
and U6720 (N_6720,N_3088,N_5867);
or U6721 (N_6721,N_5309,N_4288);
nand U6722 (N_6722,N_4348,N_5243);
nand U6723 (N_6723,N_3816,N_4392);
nand U6724 (N_6724,N_5357,N_3140);
nor U6725 (N_6725,N_4035,N_3553);
nor U6726 (N_6726,N_4253,N_5841);
or U6727 (N_6727,N_3606,N_3532);
nand U6728 (N_6728,N_4371,N_3583);
or U6729 (N_6729,N_3898,N_4505);
nor U6730 (N_6730,N_3665,N_5721);
nand U6731 (N_6731,N_5727,N_3680);
nor U6732 (N_6732,N_5019,N_3556);
or U6733 (N_6733,N_4960,N_4773);
and U6734 (N_6734,N_3572,N_3805);
or U6735 (N_6735,N_3537,N_4709);
nand U6736 (N_6736,N_5327,N_4046);
nand U6737 (N_6737,N_5296,N_5490);
or U6738 (N_6738,N_3726,N_5892);
nand U6739 (N_6739,N_5177,N_3087);
nand U6740 (N_6740,N_5011,N_3189);
nand U6741 (N_6741,N_5422,N_3354);
nand U6742 (N_6742,N_3836,N_4883);
nand U6743 (N_6743,N_3729,N_5666);
nand U6744 (N_6744,N_4897,N_4239);
nand U6745 (N_6745,N_3623,N_3596);
and U6746 (N_6746,N_3328,N_4372);
or U6747 (N_6747,N_3015,N_5884);
or U6748 (N_6748,N_3803,N_4736);
nand U6749 (N_6749,N_4999,N_3888);
nand U6750 (N_6750,N_3716,N_3158);
and U6751 (N_6751,N_3745,N_4089);
nor U6752 (N_6752,N_4630,N_3349);
or U6753 (N_6753,N_3631,N_4682);
nand U6754 (N_6754,N_4149,N_4478);
nor U6755 (N_6755,N_3381,N_5768);
and U6756 (N_6756,N_5284,N_5285);
or U6757 (N_6757,N_5183,N_3687);
or U6758 (N_6758,N_4487,N_3829);
nor U6759 (N_6759,N_4136,N_3796);
and U6760 (N_6760,N_5957,N_5475);
nand U6761 (N_6761,N_3571,N_5027);
nor U6762 (N_6762,N_5897,N_3212);
nor U6763 (N_6763,N_5372,N_5826);
or U6764 (N_6764,N_4925,N_4529);
xor U6765 (N_6765,N_3688,N_4712);
nor U6766 (N_6766,N_4544,N_5062);
or U6767 (N_6767,N_3622,N_4262);
or U6768 (N_6768,N_4256,N_3827);
nor U6769 (N_6769,N_4033,N_5268);
and U6770 (N_6770,N_3037,N_4866);
nand U6771 (N_6771,N_3291,N_3116);
or U6772 (N_6772,N_3283,N_4561);
and U6773 (N_6773,N_4081,N_5626);
nor U6774 (N_6774,N_4275,N_4681);
and U6775 (N_6775,N_3021,N_4489);
nor U6776 (N_6776,N_3082,N_4207);
nor U6777 (N_6777,N_5474,N_5649);
nand U6778 (N_6778,N_4025,N_3066);
and U6779 (N_6779,N_3712,N_5426);
and U6780 (N_6780,N_5792,N_5782);
or U6781 (N_6781,N_3480,N_3484);
nand U6782 (N_6782,N_5787,N_5863);
nand U6783 (N_6783,N_5305,N_5321);
nand U6784 (N_6784,N_3457,N_4250);
or U6785 (N_6785,N_3613,N_4340);
nor U6786 (N_6786,N_3491,N_3322);
nand U6787 (N_6787,N_5780,N_4957);
nand U6788 (N_6788,N_4205,N_4892);
nand U6789 (N_6789,N_4731,N_4906);
and U6790 (N_6790,N_3318,N_5497);
or U6791 (N_6791,N_3141,N_5922);
nand U6792 (N_6792,N_5877,N_5082);
nand U6793 (N_6793,N_5928,N_4936);
nand U6794 (N_6794,N_3817,N_4760);
nor U6795 (N_6795,N_5024,N_3430);
nor U6796 (N_6796,N_5910,N_3406);
and U6797 (N_6797,N_3058,N_3435);
or U6798 (N_6798,N_4326,N_3588);
nand U6799 (N_6799,N_4220,N_4513);
and U6800 (N_6800,N_5653,N_5015);
or U6801 (N_6801,N_5636,N_5087);
nand U6802 (N_6802,N_3346,N_4949);
and U6803 (N_6803,N_4190,N_4697);
and U6804 (N_6804,N_4121,N_3561);
nor U6805 (N_6805,N_5871,N_3243);
and U6806 (N_6806,N_5265,N_5498);
or U6807 (N_6807,N_3031,N_4998);
nand U6808 (N_6808,N_4696,N_3143);
nor U6809 (N_6809,N_5958,N_3166);
nor U6810 (N_6810,N_3564,N_4576);
or U6811 (N_6811,N_4744,N_5271);
nor U6812 (N_6812,N_3990,N_4099);
nand U6813 (N_6813,N_4143,N_3131);
and U6814 (N_6814,N_3138,N_3589);
nor U6815 (N_6815,N_5297,N_5675);
nor U6816 (N_6816,N_4878,N_5034);
or U6817 (N_6817,N_5154,N_5148);
nor U6818 (N_6818,N_3609,N_5923);
nor U6819 (N_6819,N_4748,N_3523);
nand U6820 (N_6820,N_5239,N_3690);
and U6821 (N_6821,N_4700,N_5579);
and U6822 (N_6822,N_4108,N_3265);
nand U6823 (N_6823,N_4011,N_4272);
nand U6824 (N_6824,N_5709,N_5365);
and U6825 (N_6825,N_4003,N_5581);
nand U6826 (N_6826,N_3154,N_4313);
and U6827 (N_6827,N_5551,N_3732);
nand U6828 (N_6828,N_4547,N_3414);
and U6829 (N_6829,N_4494,N_4830);
and U6830 (N_6830,N_3407,N_4402);
or U6831 (N_6831,N_3345,N_4222);
nor U6832 (N_6832,N_5382,N_4140);
nand U6833 (N_6833,N_5052,N_4862);
nor U6834 (N_6834,N_3176,N_4379);
nand U6835 (N_6835,N_5545,N_5661);
or U6836 (N_6836,N_4540,N_5569);
and U6837 (N_6837,N_3171,N_4310);
and U6838 (N_6838,N_5818,N_4471);
nand U6839 (N_6839,N_5246,N_3042);
and U6840 (N_6840,N_3489,N_5530);
nand U6841 (N_6841,N_4594,N_5949);
nand U6842 (N_6842,N_3194,N_4579);
or U6843 (N_6843,N_5149,N_4788);
nor U6844 (N_6844,N_3181,N_5656);
and U6845 (N_6845,N_4052,N_3897);
or U6846 (N_6846,N_3361,N_3534);
nand U6847 (N_6847,N_3007,N_5146);
or U6848 (N_6848,N_4620,N_3715);
nand U6849 (N_6849,N_3599,N_5040);
and U6850 (N_6850,N_3011,N_4834);
and U6851 (N_6851,N_5921,N_5605);
nand U6852 (N_6852,N_4793,N_3986);
and U6853 (N_6853,N_3474,N_5524);
nor U6854 (N_6854,N_4742,N_5223);
nand U6855 (N_6855,N_3638,N_4061);
nor U6856 (N_6856,N_5139,N_4979);
or U6857 (N_6857,N_5056,N_5273);
nor U6858 (N_6858,N_4900,N_3357);
nor U6859 (N_6859,N_3358,N_5427);
or U6860 (N_6860,N_3331,N_4442);
nor U6861 (N_6861,N_5770,N_3220);
and U6862 (N_6862,N_3929,N_5439);
and U6863 (N_6863,N_3531,N_5440);
and U6864 (N_6864,N_4173,N_4419);
or U6865 (N_6865,N_3759,N_5338);
and U6866 (N_6866,N_4063,N_3644);
or U6867 (N_6867,N_4150,N_5597);
nand U6868 (N_6868,N_4070,N_4038);
nand U6869 (N_6869,N_5198,N_3636);
nor U6870 (N_6870,N_4952,N_5603);
and U6871 (N_6871,N_5162,N_4728);
nor U6872 (N_6872,N_3675,N_4223);
nor U6873 (N_6873,N_4128,N_5870);
xnor U6874 (N_6874,N_3554,N_3214);
nor U6875 (N_6875,N_5362,N_3912);
nor U6876 (N_6876,N_5006,N_5739);
and U6877 (N_6877,N_4302,N_4889);
nand U6878 (N_6878,N_3920,N_4511);
nand U6879 (N_6879,N_3856,N_3002);
or U6880 (N_6880,N_3477,N_5882);
nand U6881 (N_6881,N_3875,N_3923);
nor U6882 (N_6882,N_3310,N_5277);
nand U6883 (N_6883,N_3530,N_5861);
and U6884 (N_6884,N_5205,N_4198);
nand U6885 (N_6885,N_4710,N_3686);
nand U6886 (N_6886,N_3508,N_3970);
nor U6887 (N_6887,N_4643,N_3933);
or U6888 (N_6888,N_5111,N_5311);
nand U6889 (N_6889,N_3799,N_3527);
nor U6890 (N_6890,N_4789,N_3151);
nand U6891 (N_6891,N_5334,N_5915);
nor U6892 (N_6892,N_3499,N_4330);
and U6893 (N_6893,N_4775,N_4860);
and U6894 (N_6894,N_3694,N_3470);
nor U6895 (N_6895,N_5729,N_4611);
nand U6896 (N_6896,N_3118,N_4984);
or U6897 (N_6897,N_4276,N_5421);
or U6898 (N_6898,N_5802,N_3266);
nand U6899 (N_6899,N_4014,N_3886);
and U6900 (N_6900,N_4248,N_3674);
nand U6901 (N_6901,N_3076,N_3937);
and U6902 (N_6902,N_5724,N_3670);
or U6903 (N_6903,N_3587,N_5488);
nor U6904 (N_6904,N_5025,N_4472);
or U6905 (N_6905,N_4947,N_5950);
nand U6906 (N_6906,N_3164,N_3254);
or U6907 (N_6907,N_3438,N_4515);
nor U6908 (N_6908,N_3584,N_5018);
nand U6909 (N_6909,N_5023,N_5850);
nand U6910 (N_6910,N_4208,N_4652);
nor U6911 (N_6911,N_4991,N_3918);
nor U6912 (N_6912,N_4804,N_4071);
nand U6913 (N_6913,N_3877,N_4316);
nor U6914 (N_6914,N_4112,N_5117);
and U6915 (N_6915,N_4844,N_3807);
and U6916 (N_6916,N_3849,N_5604);
nand U6917 (N_6917,N_3150,N_4072);
or U6918 (N_6918,N_3904,N_3791);
or U6919 (N_6919,N_4628,N_5114);
nor U6920 (N_6920,N_5353,N_5904);
and U6921 (N_6921,N_5700,N_5356);
nor U6922 (N_6922,N_5585,N_4067);
nor U6923 (N_6923,N_5423,N_3518);
nand U6924 (N_6924,N_4347,N_4343);
or U6925 (N_6925,N_3091,N_3455);
and U6926 (N_6926,N_5542,N_3027);
nor U6927 (N_6927,N_5732,N_5145);
and U6928 (N_6928,N_3691,N_4665);
and U6929 (N_6929,N_4351,N_4642);
xnor U6930 (N_6930,N_5070,N_3514);
and U6931 (N_6931,N_3218,N_5496);
nor U6932 (N_6932,N_3203,N_5905);
and U6933 (N_6933,N_3839,N_3215);
or U6934 (N_6934,N_5745,N_4539);
and U6935 (N_6935,N_4053,N_5634);
and U6936 (N_6936,N_5687,N_3397);
or U6937 (N_6937,N_4211,N_3965);
nand U6938 (N_6938,N_5381,N_5396);
and U6939 (N_6939,N_5953,N_3663);
nand U6940 (N_6940,N_3169,N_5920);
or U6941 (N_6941,N_5558,N_5979);
nor U6942 (N_6942,N_5718,N_3399);
and U6943 (N_6943,N_4141,N_4910);
nor U6944 (N_6944,N_3092,N_3047);
or U6945 (N_6945,N_4551,N_3676);
nand U6946 (N_6946,N_5249,N_3001);
nand U6947 (N_6947,N_3749,N_5374);
nor U6948 (N_6948,N_4145,N_4746);
and U6949 (N_6949,N_3656,N_4319);
nand U6950 (N_6950,N_4622,N_3960);
or U6951 (N_6951,N_3790,N_5366);
nand U6952 (N_6952,N_5799,N_5341);
or U6953 (N_6953,N_5793,N_3107);
nand U6954 (N_6954,N_4181,N_5984);
nand U6955 (N_6955,N_4180,N_3559);
nor U6956 (N_6956,N_3600,N_3940);
and U6957 (N_6957,N_4189,N_3833);
nand U6958 (N_6958,N_3999,N_4976);
and U6959 (N_6959,N_3992,N_4226);
and U6960 (N_6960,N_4503,N_4217);
and U6961 (N_6961,N_4582,N_4452);
nand U6962 (N_6962,N_4546,N_4296);
nand U6963 (N_6963,N_3654,N_3852);
or U6964 (N_6964,N_5941,N_4783);
nand U6965 (N_6965,N_4206,N_4228);
nand U6966 (N_6966,N_3054,N_4233);
nor U6967 (N_6967,N_3586,N_3483);
nor U6968 (N_6968,N_4975,N_3661);
nand U6969 (N_6969,N_4810,N_4413);
nand U6970 (N_6970,N_5598,N_3862);
nor U6971 (N_6971,N_3236,N_5692);
nor U6972 (N_6972,N_4755,N_3855);
nand U6973 (N_6973,N_4927,N_5329);
nand U6974 (N_6974,N_3983,N_4390);
and U6975 (N_6975,N_5795,N_3593);
and U6976 (N_6976,N_4845,N_5270);
and U6977 (N_6977,N_5416,N_5046);
and U6978 (N_6978,N_3896,N_3624);
nand U6979 (N_6979,N_3543,N_4439);
nor U6980 (N_6980,N_5391,N_5660);
nor U6981 (N_6981,N_4593,N_5471);
or U6982 (N_6982,N_4948,N_4723);
nand U6983 (N_6983,N_4787,N_3739);
nand U6984 (N_6984,N_4273,N_5536);
and U6985 (N_6985,N_3459,N_5698);
nor U6986 (N_6986,N_5888,N_5404);
nand U6987 (N_6987,N_5142,N_4241);
and U6988 (N_6988,N_5225,N_5280);
and U6989 (N_6989,N_3909,N_3603);
or U6990 (N_6990,N_4968,N_3752);
nor U6991 (N_6991,N_5350,N_5620);
or U6992 (N_6992,N_4122,N_4115);
nor U6993 (N_6993,N_4170,N_5531);
or U6994 (N_6994,N_3612,N_4552);
nor U6995 (N_6995,N_4004,N_3781);
and U6996 (N_6996,N_5991,N_5064);
nor U6997 (N_6997,N_5629,N_5389);
nor U6998 (N_6998,N_5164,N_3000);
and U6999 (N_6999,N_5556,N_3840);
and U7000 (N_7000,N_3857,N_3293);
nor U7001 (N_7001,N_3278,N_4224);
or U7002 (N_7002,N_4448,N_5859);
nor U7003 (N_7003,N_3943,N_4989);
and U7004 (N_7004,N_5414,N_3814);
nand U7005 (N_7005,N_5399,N_3786);
or U7006 (N_7006,N_5943,N_3421);
nand U7007 (N_7007,N_5637,N_3359);
or U7008 (N_7008,N_4572,N_5544);
or U7009 (N_7009,N_5676,N_3028);
nand U7010 (N_7010,N_3701,N_4882);
and U7011 (N_7011,N_4418,N_5031);
nand U7012 (N_7012,N_5948,N_3190);
or U7013 (N_7013,N_4260,N_3925);
nor U7014 (N_7014,N_4610,N_5109);
and U7015 (N_7015,N_5047,N_3669);
nor U7016 (N_7016,N_3980,N_3535);
or U7017 (N_7017,N_3080,N_4232);
nand U7018 (N_7018,N_3167,N_3773);
nand U7019 (N_7019,N_5981,N_4088);
and U7020 (N_7020,N_4584,N_3611);
nand U7021 (N_7021,N_5037,N_5021);
or U7022 (N_7022,N_3850,N_4857);
and U7023 (N_7023,N_3699,N_5325);
and U7024 (N_7024,N_4570,N_4384);
and U7025 (N_7025,N_3487,N_4598);
and U7026 (N_7026,N_3795,N_3368);
nor U7027 (N_7027,N_3723,N_3949);
or U7028 (N_7028,N_5434,N_4881);
or U7029 (N_7029,N_5264,N_4325);
and U7030 (N_7030,N_5397,N_4818);
nand U7031 (N_7031,N_5079,N_3424);
nand U7032 (N_7032,N_4646,N_4078);
nor U7033 (N_7033,N_4462,N_5160);
or U7034 (N_7034,N_4886,N_5237);
or U7035 (N_7035,N_4607,N_3356);
or U7036 (N_7036,N_3127,N_5304);
or U7037 (N_7037,N_3738,N_4311);
nor U7038 (N_7038,N_3372,N_4541);
and U7039 (N_7039,N_3565,N_3033);
and U7040 (N_7040,N_4907,N_4344);
nor U7041 (N_7041,N_4323,N_4055);
and U7042 (N_7042,N_5962,N_4653);
nor U7043 (N_7043,N_5430,N_4586);
nand U7044 (N_7044,N_3305,N_4730);
nand U7045 (N_7045,N_3344,N_5845);
or U7046 (N_7046,N_4899,N_5733);
and U7047 (N_7047,N_3389,N_4263);
xor U7048 (N_7048,N_3005,N_3134);
or U7049 (N_7049,N_3287,N_3478);
nor U7050 (N_7050,N_4085,N_3440);
nor U7051 (N_7051,N_3774,N_5756);
and U7052 (N_7052,N_4919,N_3764);
nand U7053 (N_7053,N_3402,N_5970);
nor U7054 (N_7054,N_3175,N_3946);
and U7055 (N_7055,N_5839,N_4049);
nand U7056 (N_7056,N_4231,N_4981);
nand U7057 (N_7057,N_4904,N_4782);
nand U7058 (N_7058,N_3240,N_5195);
nor U7059 (N_7059,N_4440,N_3279);
or U7060 (N_7060,N_5925,N_4970);
or U7061 (N_7061,N_3270,N_4166);
nand U7062 (N_7062,N_4012,N_5737);
and U7063 (N_7063,N_5753,N_5494);
nand U7064 (N_7064,N_3481,N_3113);
or U7065 (N_7065,N_4163,N_3692);
and U7066 (N_7066,N_5435,N_3419);
or U7067 (N_7067,N_3072,N_4575);
and U7068 (N_7068,N_5614,N_4427);
nor U7069 (N_7069,N_3903,N_5406);
nand U7070 (N_7070,N_3539,N_5486);
or U7071 (N_7071,N_5514,N_5715);
nor U7072 (N_7072,N_4720,N_3578);
nor U7073 (N_7073,N_4518,N_4202);
nand U7074 (N_7074,N_5419,N_3320);
or U7075 (N_7075,N_3722,N_5484);
and U7076 (N_7076,N_3930,N_5050);
and U7077 (N_7077,N_3044,N_3235);
nand U7078 (N_7078,N_4428,N_3292);
nand U7079 (N_7079,N_3955,N_5586);
xor U7080 (N_7080,N_4619,N_3219);
nor U7081 (N_7081,N_3629,N_5182);
and U7082 (N_7082,N_4992,N_5939);
nor U7083 (N_7083,N_4870,N_4258);
or U7084 (N_7084,N_4931,N_4328);
or U7085 (N_7085,N_4493,N_3837);
nand U7086 (N_7086,N_4119,N_5221);
and U7087 (N_7087,N_3146,N_3102);
nand U7088 (N_7088,N_4060,N_4209);
or U7089 (N_7089,N_3895,N_3869);
and U7090 (N_7090,N_3935,N_5528);
nand U7091 (N_7091,N_5804,N_5228);
nor U7092 (N_7092,N_5774,N_5101);
or U7093 (N_7093,N_5209,N_4890);
or U7094 (N_7094,N_5952,N_3085);
or U7095 (N_7095,N_4849,N_4691);
nand U7096 (N_7096,N_5071,N_5817);
or U7097 (N_7097,N_5805,N_3319);
and U7098 (N_7098,N_4574,N_5229);
or U7099 (N_7099,N_3772,N_3382);
nand U7100 (N_7100,N_3891,N_5771);
nor U7101 (N_7101,N_5683,N_4659);
and U7102 (N_7102,N_5931,N_5749);
or U7103 (N_7103,N_5967,N_3997);
and U7104 (N_7104,N_3460,N_3968);
nor U7105 (N_7105,N_3504,N_3882);
and U7106 (N_7106,N_3924,N_5681);
nand U7107 (N_7107,N_3985,N_5138);
or U7108 (N_7108,N_3982,N_3471);
nor U7109 (N_7109,N_5613,N_5747);
and U7110 (N_7110,N_3810,N_4459);
nand U7111 (N_7111,N_4096,N_5717);
nand U7112 (N_7112,N_3524,N_4771);
and U7113 (N_7113,N_3736,N_5240);
and U7114 (N_7114,N_3405,N_5380);
or U7115 (N_7115,N_4507,N_4679);
nand U7116 (N_7116,N_5781,N_3926);
nor U7117 (N_7117,N_3843,N_4395);
or U7118 (N_7118,N_5482,N_3628);
and U7119 (N_7119,N_4738,N_4690);
nand U7120 (N_7120,N_4298,N_3355);
nand U7121 (N_7121,N_3045,N_5889);
and U7122 (N_7122,N_5691,N_5213);
nand U7123 (N_7123,N_3295,N_4556);
and U7124 (N_7124,N_3525,N_4317);
nor U7125 (N_7125,N_5058,N_4138);
and U7126 (N_7126,N_5898,N_3512);
nor U7127 (N_7127,N_3466,N_4243);
nor U7128 (N_7128,N_3808,N_3333);
or U7129 (N_7129,N_3057,N_3778);
nand U7130 (N_7130,N_3393,N_3180);
nor U7131 (N_7131,N_4754,N_3717);
or U7132 (N_7132,N_4235,N_4708);
nand U7133 (N_7133,N_3051,N_4993);
or U7134 (N_7134,N_3761,N_5642);
nand U7135 (N_7135,N_5852,N_3828);
nand U7136 (N_7136,N_4285,N_4958);
nand U7137 (N_7137,N_3197,N_5281);
nand U7138 (N_7138,N_5978,N_5014);
and U7139 (N_7139,N_4349,N_4229);
nor U7140 (N_7140,N_3241,N_3083);
nand U7141 (N_7141,N_4378,N_5324);
and U7142 (N_7142,N_3735,N_5903);
or U7143 (N_7143,N_5169,N_3700);
and U7144 (N_7144,N_4043,N_5933);
and U7145 (N_7145,N_5797,N_5032);
nor U7146 (N_7146,N_3967,N_4868);
and U7147 (N_7147,N_3251,N_3101);
nor U7148 (N_7148,N_3777,N_4101);
and U7149 (N_7149,N_3264,N_4279);
nor U7150 (N_7150,N_3931,N_5227);
nand U7151 (N_7151,N_4757,N_5269);
nor U7152 (N_7152,N_4165,N_4595);
or U7153 (N_7153,N_5690,N_5012);
or U7154 (N_7154,N_3652,N_4426);
nand U7155 (N_7155,N_4443,N_4300);
nand U7156 (N_7156,N_4234,N_3741);
or U7157 (N_7157,N_5128,N_4496);
nor U7158 (N_7158,N_4916,N_3590);
nand U7159 (N_7159,N_5989,N_3269);
nor U7160 (N_7160,N_5250,N_3352);
and U7161 (N_7161,N_4675,N_4287);
and U7162 (N_7162,N_5583,N_3391);
nand U7163 (N_7163,N_5919,N_4671);
nor U7164 (N_7164,N_4912,N_3964);
nor U7165 (N_7165,N_3991,N_5403);
and U7166 (N_7166,N_5773,N_4192);
nor U7167 (N_7167,N_5838,N_4221);
nor U7168 (N_7168,N_4214,N_4095);
or U7169 (N_7169,N_5594,N_5625);
nand U7170 (N_7170,N_4603,N_4626);
nand U7171 (N_7171,N_3223,N_4758);
and U7172 (N_7172,N_3919,N_5107);
and U7173 (N_7173,N_3103,N_4169);
nand U7174 (N_7174,N_4009,N_5369);
and U7175 (N_7175,N_3495,N_4445);
or U7176 (N_7176,N_4282,N_5638);
or U7177 (N_7177,N_4533,N_4654);
and U7178 (N_7178,N_3303,N_4918);
and U7179 (N_7179,N_3373,N_4270);
nand U7180 (N_7180,N_3939,N_3747);
and U7181 (N_7181,N_4567,N_5259);
or U7182 (N_7182,N_4476,N_5800);
or U7183 (N_7183,N_5654,N_5658);
nand U7184 (N_7184,N_4050,N_5520);
or U7185 (N_7185,N_5136,N_3059);
nand U7186 (N_7186,N_4741,N_5664);
and U7187 (N_7187,N_3413,N_4306);
or U7188 (N_7188,N_5286,N_5914);
nand U7189 (N_7189,N_3117,N_4125);
and U7190 (N_7190,N_5645,N_5832);
nand U7191 (N_7191,N_4353,N_4971);
and U7192 (N_7192,N_3443,N_4444);
nand U7193 (N_7193,N_5411,N_3621);
nor U7194 (N_7194,N_5290,N_3314);
or U7195 (N_7195,N_3806,N_4200);
nand U7196 (N_7196,N_5123,N_5609);
nor U7197 (N_7197,N_4386,N_4698);
or U7198 (N_7198,N_4522,N_5885);
and U7199 (N_7199,N_4333,N_3604);
and U7200 (N_7200,N_4517,N_4737);
nand U7201 (N_7201,N_3018,N_4663);
nor U7202 (N_7202,N_3468,N_3826);
or U7203 (N_7203,N_4367,N_3973);
and U7204 (N_7204,N_4641,N_4838);
nand U7205 (N_7205,N_5479,N_4242);
nor U7206 (N_7206,N_3379,N_4893);
nor U7207 (N_7207,N_4408,N_4079);
and U7208 (N_7208,N_5466,N_3277);
nand U7209 (N_7209,N_5766,N_5862);
nor U7210 (N_7210,N_5328,N_5508);
nor U7211 (N_7211,N_3540,N_3337);
and U7212 (N_7212,N_3811,N_4040);
or U7213 (N_7213,N_4196,N_3598);
nor U7214 (N_7214,N_5103,N_5719);
and U7215 (N_7215,N_3157,N_4608);
or U7216 (N_7216,N_4363,N_3908);
nor U7217 (N_7217,N_4185,N_3378);
and U7218 (N_7218,N_5783,N_3635);
and U7219 (N_7219,N_3592,N_5811);
nor U7220 (N_7220,N_3575,N_5493);
nor U7221 (N_7221,N_5091,N_4634);
and U7222 (N_7222,N_5833,N_4841);
or U7223 (N_7223,N_4799,N_4469);
and U7224 (N_7224,N_4153,N_5513);
and U7225 (N_7225,N_3447,N_4090);
nand U7226 (N_7226,N_5355,N_5402);
and U7227 (N_7227,N_4530,N_5980);
or U7228 (N_7228,N_4191,N_5974);
xor U7229 (N_7229,N_5168,N_4896);
nor U7230 (N_7230,N_3698,N_4230);
nor U7231 (N_7231,N_3702,N_5455);
and U7232 (N_7232,N_5895,N_5119);
and U7233 (N_7233,N_4194,N_4940);
and U7234 (N_7234,N_5972,N_4369);
nand U7235 (N_7235,N_4354,N_3526);
and U7236 (N_7236,N_4920,N_5300);
nor U7237 (N_7237,N_5600,N_5436);
nor U7238 (N_7238,N_5893,N_5373);
nor U7239 (N_7239,N_3204,N_3906);
or U7240 (N_7240,N_3948,N_4846);
nand U7241 (N_7241,N_3453,N_5059);
nand U7242 (N_7242,N_4523,N_4609);
nand U7243 (N_7243,N_3563,N_3789);
nand U7244 (N_7244,N_3130,N_3662);
xnor U7245 (N_7245,N_5790,N_4985);
or U7246 (N_7246,N_3192,N_3878);
nor U7247 (N_7247,N_3643,N_4255);
nor U7248 (N_7248,N_3892,N_3039);
or U7249 (N_7249,N_4212,N_3416);
or U7250 (N_7250,N_3205,N_4491);
nand U7251 (N_7251,N_3023,N_5521);
nand U7252 (N_7252,N_4144,N_5506);
and U7253 (N_7253,N_5048,N_4550);
and U7254 (N_7254,N_4178,N_3456);
nand U7255 (N_7255,N_4237,N_5180);
nor U7256 (N_7256,N_4341,N_3660);
or U7257 (N_7257,N_4769,N_4148);
nor U7258 (N_7258,N_5231,N_4809);
or U7259 (N_7259,N_5163,N_3899);
nand U7260 (N_7260,N_3608,N_3353);
and U7261 (N_7261,N_5245,N_3792);
nor U7262 (N_7262,N_3133,N_5602);
nand U7263 (N_7263,N_4616,N_3348);
nand U7264 (N_7264,N_4528,N_3119);
and U7265 (N_7265,N_5345,N_5909);
and U7266 (N_7266,N_4688,N_5881);
nand U7267 (N_7267,N_3881,N_5644);
or U7268 (N_7268,N_5995,N_5955);
and U7269 (N_7269,N_4715,N_4733);
and U7270 (N_7270,N_4289,N_5348);
or U7271 (N_7271,N_5860,N_3766);
nor U7272 (N_7272,N_4403,N_3472);
nor U7273 (N_7273,N_3401,N_3961);
nand U7274 (N_7274,N_3619,N_4468);
or U7275 (N_7275,N_3953,N_5401);
xnor U7276 (N_7276,N_5262,N_4871);
or U7277 (N_7277,N_4854,N_3610);
nand U7278 (N_7278,N_4007,N_3591);
nand U7279 (N_7279,N_4568,N_5067);
or U7280 (N_7280,N_3802,N_3568);
nor U7281 (N_7281,N_4160,N_5219);
and U7282 (N_7282,N_5742,N_5788);
or U7283 (N_7283,N_3207,N_3788);
or U7284 (N_7284,N_3492,N_4600);
nand U7285 (N_7285,N_4179,N_4436);
nor U7286 (N_7286,N_4215,N_3538);
nand U7287 (N_7287,N_3502,N_5582);
nor U7288 (N_7288,N_3014,N_5842);
and U7289 (N_7289,N_3247,N_5452);
or U7290 (N_7290,N_3019,N_5865);
nand U7291 (N_7291,N_5463,N_4825);
nand U7292 (N_7292,N_4557,N_3095);
and U7293 (N_7293,N_5932,N_3801);
and U7294 (N_7294,N_3408,N_4974);
nand U7295 (N_7295,N_5743,N_4722);
nand U7296 (N_7296,N_3950,N_5186);
nor U7297 (N_7297,N_4637,N_4835);
nand U7298 (N_7298,N_4942,N_4614);
nor U7299 (N_7299,N_3041,N_5671);
nand U7300 (N_7300,N_4621,N_3727);
and U7301 (N_7301,N_5809,N_5009);
or U7302 (N_7302,N_4417,N_3633);
or U7303 (N_7303,N_5193,N_5640);
and U7304 (N_7304,N_5303,N_3962);
or U7305 (N_7305,N_5529,N_5055);
nor U7306 (N_7306,N_4764,N_5211);
and U7307 (N_7307,N_3577,N_4346);
nor U7308 (N_7308,N_3060,N_4449);
and U7309 (N_7309,N_5960,N_4911);
or U7310 (N_7310,N_4972,N_3555);
and U7311 (N_7311,N_4677,N_4100);
nand U7312 (N_7312,N_3420,N_5057);
nand U7313 (N_7313,N_4132,N_5344);
nor U7314 (N_7314,N_3121,N_5393);
and U7315 (N_7315,N_4604,N_4293);
or U7316 (N_7316,N_3469,N_3601);
and U7317 (N_7317,N_4002,N_3268);
nor U7318 (N_7318,N_3630,N_3434);
or U7319 (N_7319,N_5564,N_4705);
nand U7320 (N_7320,N_3342,N_3226);
nor U7321 (N_7321,N_5740,N_4303);
nor U7322 (N_7322,N_4647,N_5607);
nor U7323 (N_7323,N_3721,N_5166);
nor U7324 (N_7324,N_3347,N_5791);
and U7325 (N_7325,N_4309,N_4329);
and U7326 (N_7326,N_4884,N_4759);
or U7327 (N_7327,N_3366,N_3705);
or U7328 (N_7328,N_5126,N_4389);
nand U7329 (N_7329,N_3972,N_5685);
nand U7330 (N_7330,N_5363,N_5532);
nor U7331 (N_7331,N_5282,N_4729);
or U7332 (N_7332,N_5786,N_5930);
nor U7333 (N_7333,N_3820,N_5016);
nand U7334 (N_7334,N_4569,N_5313);
and U7335 (N_7335,N_5210,N_5175);
or U7336 (N_7336,N_3445,N_3374);
or U7337 (N_7337,N_5971,N_3052);
or U7338 (N_7338,N_5453,N_4915);
or U7339 (N_7339,N_4588,N_3415);
nor U7340 (N_7340,N_4779,N_3081);
or U7341 (N_7341,N_3422,N_3921);
nor U7342 (N_7342,N_5697,N_5443);
nand U7343 (N_7343,N_5445,N_5413);
or U7344 (N_7344,N_4406,N_5132);
nor U7345 (N_7345,N_5866,N_4435);
nand U7346 (N_7346,N_3570,N_3969);
nor U7347 (N_7347,N_4587,N_5244);
nand U7348 (N_7348,N_5236,N_4873);
nor U7349 (N_7349,N_5007,N_3507);
nand U7350 (N_7350,N_5147,N_5927);
nand U7351 (N_7351,N_4851,N_5323);
and U7352 (N_7352,N_4592,N_4928);
nand U7353 (N_7353,N_5894,N_3995);
nand U7354 (N_7354,N_3156,N_4394);
nor U7355 (N_7355,N_4645,N_4623);
nor U7356 (N_7356,N_4247,N_5663);
and U7357 (N_7357,N_4249,N_3210);
or U7358 (N_7358,N_4895,N_5383);
and U7359 (N_7359,N_5464,N_4941);
nor U7360 (N_7360,N_4532,N_4005);
nor U7361 (N_7361,N_4756,N_5340);
nand U7362 (N_7362,N_3375,N_3308);
or U7363 (N_7363,N_4898,N_3851);
nand U7364 (N_7364,N_5069,N_4888);
nor U7365 (N_7365,N_4114,N_5630);
or U7366 (N_7366,N_5546,N_4307);
nand U7367 (N_7367,N_5765,N_5415);
nor U7368 (N_7368,N_5789,N_5612);
nand U7369 (N_7369,N_5113,N_5361);
nand U7370 (N_7370,N_3651,N_3841);
nand U7371 (N_7371,N_3321,N_4139);
or U7372 (N_7372,N_3783,N_5964);
nor U7373 (N_7373,N_5844,N_3945);
or U7374 (N_7374,N_5125,N_5622);
nand U7375 (N_7375,N_4454,N_3186);
and U7376 (N_7376,N_5523,N_5527);
nand U7377 (N_7377,N_5447,N_3304);
nor U7378 (N_7378,N_4953,N_3704);
nand U7379 (N_7379,N_4555,N_4578);
and U7380 (N_7380,N_4130,N_3520);
nor U7381 (N_7381,N_5834,N_4986);
nor U7382 (N_7382,N_5510,N_4037);
or U7383 (N_7383,N_4076,N_5476);
nor U7384 (N_7384,N_5491,N_5410);
nand U7385 (N_7385,N_5392,N_3846);
nand U7386 (N_7386,N_4441,N_5767);
or U7387 (N_7387,N_3030,N_4770);
or U7388 (N_7388,N_3494,N_3664);
nor U7389 (N_7389,N_5571,N_3271);
and U7390 (N_7390,N_3750,N_3874);
nor U7391 (N_7391,N_4355,N_5688);
or U7392 (N_7392,N_5005,N_3312);
nor U7393 (N_7393,N_3673,N_5535);
and U7394 (N_7394,N_5261,N_3517);
nand U7395 (N_7395,N_4133,N_5824);
nand U7396 (N_7396,N_4373,N_4840);
and U7397 (N_7397,N_4097,N_4172);
or U7398 (N_7398,N_3876,N_5918);
or U7399 (N_7399,N_4396,N_5590);
nand U7400 (N_7400,N_4792,N_5601);
and U7401 (N_7401,N_5975,N_3509);
nand U7402 (N_7402,N_5987,N_4254);
nand U7403 (N_7403,N_5333,N_4689);
or U7404 (N_7404,N_3327,N_3441);
and U7405 (N_7405,N_5469,N_5094);
and U7406 (N_7406,N_4312,N_5028);
xnor U7407 (N_7407,N_5983,N_5351);
nor U7408 (N_7408,N_4370,N_4693);
or U7409 (N_7409,N_3351,N_3513);
nor U7410 (N_7410,N_5580,N_5159);
or U7411 (N_7411,N_5317,N_3067);
and U7412 (N_7412,N_5617,N_5200);
or U7413 (N_7413,N_3099,N_4685);
and U7414 (N_7414,N_5821,N_5985);
nor U7415 (N_7415,N_4765,N_4240);
nor U7416 (N_7416,N_3510,N_4537);
or U7417 (N_7417,N_5224,N_4105);
nor U7418 (N_7418,N_3975,N_4772);
nor U7419 (N_7419,N_4525,N_4813);
or U7420 (N_7420,N_5039,N_3860);
nand U7421 (N_7421,N_5611,N_5187);
nand U7422 (N_7422,N_4995,N_3006);
and U7423 (N_7423,N_4075,N_5207);
nor U7424 (N_7424,N_5165,N_4997);
nor U7425 (N_7425,N_3625,N_4027);
nand U7426 (N_7426,N_3566,N_3387);
and U7427 (N_7427,N_5772,N_5112);
or U7428 (N_7428,N_3315,N_5840);
and U7429 (N_7429,N_3046,N_5331);
or U7430 (N_7430,N_4657,N_3142);
nor U7431 (N_7431,N_3339,N_5777);
or U7432 (N_7432,N_4177,N_4082);
nand U7433 (N_7433,N_5143,N_5994);
or U7434 (N_7434,N_3755,N_4463);
nand U7435 (N_7435,N_3135,N_4292);
or U7436 (N_7436,N_3343,N_3238);
nor U7437 (N_7437,N_5429,N_4833);
and U7438 (N_7438,N_4376,N_4676);
nor U7439 (N_7439,N_3301,N_5346);
or U7440 (N_7440,N_5525,N_4926);
nand U7441 (N_7441,N_3394,N_3893);
nor U7442 (N_7442,N_4820,N_4278);
or U7443 (N_7443,N_3809,N_3137);
nor U7444 (N_7444,N_4391,N_3211);
or U7445 (N_7445,N_5302,N_5100);
nand U7446 (N_7446,N_5534,N_5289);
and U7447 (N_7447,N_3845,N_4358);
and U7448 (N_7448,N_4887,N_5728);
and U7449 (N_7449,N_4339,N_3671);
or U7450 (N_7450,N_4350,N_4684);
nor U7451 (N_7451,N_3093,N_5384);
and U7452 (N_7452,N_3842,N_4479);
or U7453 (N_7453,N_3734,N_3758);
nand U7454 (N_7454,N_5337,N_5725);
nand U7455 (N_7455,N_4930,N_3620);
or U7456 (N_7456,N_5711,N_3267);
and U7457 (N_7457,N_5543,N_3784);
and U7458 (N_7458,N_4566,N_3488);
nor U7459 (N_7459,N_3371,N_5662);
or U7460 (N_7460,N_4162,N_5199);
and U7461 (N_7461,N_3426,N_3079);
nor U7462 (N_7462,N_3289,N_5140);
nand U7463 (N_7463,N_3776,N_5722);
nor U7464 (N_7464,N_4861,N_5990);
or U7465 (N_7465,N_5487,N_5552);
nand U7466 (N_7466,N_3209,N_3288);
or U7467 (N_7467,N_3552,N_5830);
and U7468 (N_7468,N_5735,N_5433);
nand U7469 (N_7469,N_5167,N_4383);
nand U7470 (N_7470,N_4451,N_5092);
nand U7471 (N_7471,N_3341,N_5121);
nand U7472 (N_7472,N_3105,N_4399);
or U7473 (N_7473,N_3187,N_5468);
or U7474 (N_7474,N_5053,N_5539);
and U7475 (N_7475,N_5835,N_3501);
nor U7476 (N_7476,N_4245,N_4727);
nor U7477 (N_7477,N_5624,N_5526);
nor U7478 (N_7478,N_3084,N_5999);
or U7479 (N_7479,N_5699,N_4107);
and U7480 (N_7480,N_3905,N_5755);
nand U7481 (N_7481,N_5851,N_5855);
nor U7482 (N_7482,N_4602,N_3988);
and U7483 (N_7483,N_3996,N_3020);
nor U7484 (N_7484,N_4865,N_4560);
nor U7485 (N_7485,N_3050,N_5176);
nand U7486 (N_7486,N_5561,N_4280);
nand U7487 (N_7487,N_4719,N_3233);
and U7488 (N_7488,N_3069,N_4983);
nor U7489 (N_7489,N_4322,N_3743);
nand U7490 (N_7490,N_5706,N_3617);
nor U7491 (N_7491,N_4822,N_3889);
nor U7492 (N_7492,N_4091,N_4509);
or U7493 (N_7493,N_5319,N_3246);
or U7494 (N_7494,N_3296,N_5853);
nand U7495 (N_7495,N_4795,N_4218);
and U7496 (N_7496,N_4499,N_4631);
and U7497 (N_7497,N_5252,N_3533);
nand U7498 (N_7498,N_5238,N_4914);
nand U7499 (N_7499,N_4131,N_5516);
or U7500 (N_7500,N_3949,N_3961);
and U7501 (N_7501,N_4289,N_5293);
nor U7502 (N_7502,N_5369,N_3029);
and U7503 (N_7503,N_4849,N_5937);
nand U7504 (N_7504,N_5918,N_3429);
and U7505 (N_7505,N_3235,N_5382);
or U7506 (N_7506,N_5167,N_4496);
or U7507 (N_7507,N_3392,N_5904);
or U7508 (N_7508,N_5804,N_3154);
nor U7509 (N_7509,N_4262,N_3220);
nand U7510 (N_7510,N_4552,N_3747);
or U7511 (N_7511,N_4757,N_5470);
and U7512 (N_7512,N_4078,N_4754);
or U7513 (N_7513,N_5903,N_3713);
and U7514 (N_7514,N_5308,N_3134);
nand U7515 (N_7515,N_5086,N_4027);
nor U7516 (N_7516,N_3084,N_4566);
nor U7517 (N_7517,N_5913,N_4381);
and U7518 (N_7518,N_5514,N_5139);
and U7519 (N_7519,N_5598,N_4581);
nand U7520 (N_7520,N_4405,N_4164);
or U7521 (N_7521,N_4406,N_4240);
nor U7522 (N_7522,N_3493,N_5179);
and U7523 (N_7523,N_5537,N_5446);
nor U7524 (N_7524,N_3500,N_5145);
or U7525 (N_7525,N_5791,N_4560);
nand U7526 (N_7526,N_3069,N_5402);
nor U7527 (N_7527,N_3747,N_5591);
or U7528 (N_7528,N_4312,N_5287);
nor U7529 (N_7529,N_4022,N_5702);
nand U7530 (N_7530,N_5650,N_3594);
or U7531 (N_7531,N_5231,N_4067);
or U7532 (N_7532,N_3256,N_3731);
or U7533 (N_7533,N_4749,N_5834);
and U7534 (N_7534,N_4787,N_3367);
and U7535 (N_7535,N_5649,N_5309);
nor U7536 (N_7536,N_5561,N_4718);
nand U7537 (N_7537,N_3533,N_4403);
nand U7538 (N_7538,N_4875,N_3921);
and U7539 (N_7539,N_4705,N_3631);
nand U7540 (N_7540,N_5157,N_4020);
nor U7541 (N_7541,N_4335,N_3424);
and U7542 (N_7542,N_3107,N_5314);
nor U7543 (N_7543,N_4912,N_4339);
nand U7544 (N_7544,N_5314,N_5285);
nor U7545 (N_7545,N_4880,N_3229);
and U7546 (N_7546,N_5718,N_3937);
nor U7547 (N_7547,N_4636,N_5659);
nor U7548 (N_7548,N_3760,N_4539);
nor U7549 (N_7549,N_5738,N_5579);
and U7550 (N_7550,N_3614,N_4492);
and U7551 (N_7551,N_5530,N_4831);
or U7552 (N_7552,N_5166,N_5860);
and U7553 (N_7553,N_4503,N_5795);
and U7554 (N_7554,N_3159,N_3764);
and U7555 (N_7555,N_5231,N_3575);
nand U7556 (N_7556,N_3869,N_3400);
nand U7557 (N_7557,N_4624,N_5592);
nand U7558 (N_7558,N_4926,N_4352);
and U7559 (N_7559,N_5098,N_3422);
nand U7560 (N_7560,N_4016,N_5872);
or U7561 (N_7561,N_4145,N_3773);
or U7562 (N_7562,N_5927,N_3773);
and U7563 (N_7563,N_4472,N_5745);
and U7564 (N_7564,N_4818,N_4586);
or U7565 (N_7565,N_3699,N_3974);
nor U7566 (N_7566,N_3105,N_3925);
nor U7567 (N_7567,N_4587,N_5228);
and U7568 (N_7568,N_4279,N_4029);
nor U7569 (N_7569,N_3850,N_5155);
or U7570 (N_7570,N_5319,N_5462);
or U7571 (N_7571,N_4175,N_5560);
nand U7572 (N_7572,N_5031,N_3657);
or U7573 (N_7573,N_3645,N_4407);
and U7574 (N_7574,N_3434,N_4747);
nor U7575 (N_7575,N_3645,N_5173);
nand U7576 (N_7576,N_3281,N_5582);
or U7577 (N_7577,N_4608,N_5597);
or U7578 (N_7578,N_3882,N_5266);
or U7579 (N_7579,N_5465,N_3900);
or U7580 (N_7580,N_5805,N_4380);
nor U7581 (N_7581,N_4008,N_4616);
xor U7582 (N_7582,N_4227,N_5203);
nor U7583 (N_7583,N_4101,N_5498);
nand U7584 (N_7584,N_3011,N_5115);
or U7585 (N_7585,N_5818,N_4311);
nand U7586 (N_7586,N_3137,N_3830);
nor U7587 (N_7587,N_4615,N_3239);
or U7588 (N_7588,N_3988,N_3673);
nand U7589 (N_7589,N_4320,N_5303);
nand U7590 (N_7590,N_5837,N_4918);
or U7591 (N_7591,N_5869,N_5209);
and U7592 (N_7592,N_5950,N_3036);
or U7593 (N_7593,N_4984,N_4925);
and U7594 (N_7594,N_3932,N_4384);
nor U7595 (N_7595,N_4299,N_3712);
or U7596 (N_7596,N_4384,N_5978);
nor U7597 (N_7597,N_4411,N_4216);
and U7598 (N_7598,N_4743,N_3940);
or U7599 (N_7599,N_3199,N_4032);
nand U7600 (N_7600,N_5123,N_4337);
or U7601 (N_7601,N_4932,N_3466);
or U7602 (N_7602,N_5448,N_5868);
nand U7603 (N_7603,N_5460,N_3605);
and U7604 (N_7604,N_3534,N_5840);
nor U7605 (N_7605,N_5207,N_4385);
and U7606 (N_7606,N_4729,N_5788);
or U7607 (N_7607,N_5889,N_3863);
nand U7608 (N_7608,N_3886,N_5392);
nand U7609 (N_7609,N_5058,N_3607);
and U7610 (N_7610,N_3722,N_3337);
nand U7611 (N_7611,N_4997,N_4138);
or U7612 (N_7612,N_5578,N_3046);
nand U7613 (N_7613,N_5609,N_5888);
or U7614 (N_7614,N_5948,N_5223);
nand U7615 (N_7615,N_4437,N_3208);
or U7616 (N_7616,N_3014,N_5455);
nand U7617 (N_7617,N_5643,N_3395);
nor U7618 (N_7618,N_5111,N_4561);
and U7619 (N_7619,N_4401,N_4906);
nor U7620 (N_7620,N_3989,N_5494);
nor U7621 (N_7621,N_4479,N_4916);
nand U7622 (N_7622,N_4560,N_5225);
or U7623 (N_7623,N_4329,N_5704);
or U7624 (N_7624,N_5028,N_4178);
and U7625 (N_7625,N_3452,N_4903);
nand U7626 (N_7626,N_4523,N_4423);
and U7627 (N_7627,N_5281,N_3049);
nor U7628 (N_7628,N_3004,N_5710);
nand U7629 (N_7629,N_4126,N_5670);
and U7630 (N_7630,N_3978,N_4234);
and U7631 (N_7631,N_4278,N_3247);
nor U7632 (N_7632,N_5712,N_3617);
or U7633 (N_7633,N_4516,N_3984);
nand U7634 (N_7634,N_4768,N_3684);
nor U7635 (N_7635,N_4064,N_4040);
nor U7636 (N_7636,N_5628,N_3567);
or U7637 (N_7637,N_5730,N_3826);
and U7638 (N_7638,N_5246,N_3052);
or U7639 (N_7639,N_3521,N_4772);
nand U7640 (N_7640,N_4386,N_4510);
and U7641 (N_7641,N_3692,N_3175);
or U7642 (N_7642,N_4901,N_4301);
nand U7643 (N_7643,N_4842,N_3919);
and U7644 (N_7644,N_5140,N_5383);
nand U7645 (N_7645,N_5457,N_5624);
and U7646 (N_7646,N_4823,N_4613);
or U7647 (N_7647,N_5634,N_5585);
or U7648 (N_7648,N_3584,N_3880);
and U7649 (N_7649,N_3854,N_4466);
nor U7650 (N_7650,N_5891,N_5064);
or U7651 (N_7651,N_3545,N_5396);
nor U7652 (N_7652,N_5356,N_5790);
nand U7653 (N_7653,N_4953,N_3773);
nand U7654 (N_7654,N_5167,N_4711);
nor U7655 (N_7655,N_5365,N_3040);
or U7656 (N_7656,N_5028,N_4641);
nor U7657 (N_7657,N_4101,N_3467);
nor U7658 (N_7658,N_4298,N_4140);
and U7659 (N_7659,N_3981,N_4017);
and U7660 (N_7660,N_3738,N_5285);
and U7661 (N_7661,N_5432,N_3385);
or U7662 (N_7662,N_4666,N_5176);
or U7663 (N_7663,N_5904,N_3340);
or U7664 (N_7664,N_3102,N_5817);
nand U7665 (N_7665,N_3631,N_3941);
nand U7666 (N_7666,N_5882,N_3786);
or U7667 (N_7667,N_4848,N_3145);
or U7668 (N_7668,N_5010,N_4197);
nor U7669 (N_7669,N_4584,N_5774);
and U7670 (N_7670,N_3182,N_5837);
nand U7671 (N_7671,N_3612,N_3348);
and U7672 (N_7672,N_4073,N_3579);
nor U7673 (N_7673,N_4513,N_5425);
and U7674 (N_7674,N_5278,N_3073);
nand U7675 (N_7675,N_4444,N_5297);
nand U7676 (N_7676,N_4801,N_4580);
nor U7677 (N_7677,N_3683,N_3491);
nand U7678 (N_7678,N_3952,N_4951);
nand U7679 (N_7679,N_5809,N_3684);
or U7680 (N_7680,N_3487,N_4580);
or U7681 (N_7681,N_3807,N_5174);
nand U7682 (N_7682,N_5241,N_4537);
nand U7683 (N_7683,N_3629,N_5975);
or U7684 (N_7684,N_3561,N_4806);
xor U7685 (N_7685,N_4261,N_3243);
or U7686 (N_7686,N_5066,N_3109);
and U7687 (N_7687,N_3174,N_5073);
nor U7688 (N_7688,N_5356,N_3865);
xnor U7689 (N_7689,N_5930,N_4892);
nor U7690 (N_7690,N_3145,N_4535);
and U7691 (N_7691,N_4023,N_3726);
nor U7692 (N_7692,N_4793,N_4475);
and U7693 (N_7693,N_5835,N_4234);
and U7694 (N_7694,N_5900,N_3805);
or U7695 (N_7695,N_4463,N_5523);
and U7696 (N_7696,N_5958,N_4249);
nand U7697 (N_7697,N_5668,N_4491);
or U7698 (N_7698,N_3858,N_5579);
nand U7699 (N_7699,N_3020,N_4893);
or U7700 (N_7700,N_4023,N_3082);
and U7701 (N_7701,N_5644,N_5803);
nor U7702 (N_7702,N_5543,N_4961);
and U7703 (N_7703,N_4238,N_3244);
and U7704 (N_7704,N_5237,N_4377);
or U7705 (N_7705,N_5396,N_3644);
xnor U7706 (N_7706,N_3550,N_3389);
nand U7707 (N_7707,N_3746,N_4733);
and U7708 (N_7708,N_3990,N_5296);
nor U7709 (N_7709,N_4143,N_3470);
and U7710 (N_7710,N_3406,N_5629);
nor U7711 (N_7711,N_4258,N_5720);
nand U7712 (N_7712,N_5829,N_4924);
nand U7713 (N_7713,N_4163,N_3795);
or U7714 (N_7714,N_4403,N_5843);
or U7715 (N_7715,N_4417,N_4218);
nand U7716 (N_7716,N_3201,N_3540);
nor U7717 (N_7717,N_3996,N_5377);
or U7718 (N_7718,N_5696,N_5720);
and U7719 (N_7719,N_4790,N_5473);
nand U7720 (N_7720,N_5573,N_4590);
and U7721 (N_7721,N_3366,N_5401);
or U7722 (N_7722,N_4409,N_3413);
or U7723 (N_7723,N_5373,N_4097);
or U7724 (N_7724,N_3964,N_4861);
nor U7725 (N_7725,N_5986,N_3414);
nand U7726 (N_7726,N_5681,N_3495);
or U7727 (N_7727,N_5347,N_5357);
nor U7728 (N_7728,N_5314,N_3121);
and U7729 (N_7729,N_3515,N_5906);
or U7730 (N_7730,N_3676,N_3612);
nor U7731 (N_7731,N_5677,N_5595);
and U7732 (N_7732,N_5039,N_5626);
or U7733 (N_7733,N_3974,N_4806);
nand U7734 (N_7734,N_3698,N_5249);
or U7735 (N_7735,N_4853,N_3300);
nand U7736 (N_7736,N_3147,N_3020);
or U7737 (N_7737,N_3466,N_4562);
nand U7738 (N_7738,N_5123,N_4444);
nor U7739 (N_7739,N_3963,N_3445);
nand U7740 (N_7740,N_5834,N_4478);
or U7741 (N_7741,N_5976,N_4044);
nand U7742 (N_7742,N_4394,N_4403);
and U7743 (N_7743,N_3099,N_3360);
or U7744 (N_7744,N_3239,N_3819);
and U7745 (N_7745,N_3504,N_5918);
nor U7746 (N_7746,N_5438,N_5856);
nor U7747 (N_7747,N_4398,N_5124);
nor U7748 (N_7748,N_3551,N_3885);
xnor U7749 (N_7749,N_5576,N_4696);
nand U7750 (N_7750,N_3275,N_3348);
nand U7751 (N_7751,N_5761,N_5956);
nor U7752 (N_7752,N_3066,N_3080);
and U7753 (N_7753,N_4962,N_5598);
nor U7754 (N_7754,N_3331,N_5072);
and U7755 (N_7755,N_5899,N_5568);
and U7756 (N_7756,N_3608,N_4203);
and U7757 (N_7757,N_5260,N_4619);
nand U7758 (N_7758,N_5848,N_5511);
or U7759 (N_7759,N_4687,N_3865);
nor U7760 (N_7760,N_3368,N_4145);
or U7761 (N_7761,N_4230,N_5271);
nand U7762 (N_7762,N_4263,N_4799);
nor U7763 (N_7763,N_3972,N_3982);
xnor U7764 (N_7764,N_3425,N_5658);
or U7765 (N_7765,N_3376,N_3590);
nand U7766 (N_7766,N_5470,N_5514);
and U7767 (N_7767,N_5985,N_3565);
or U7768 (N_7768,N_3620,N_5342);
nand U7769 (N_7769,N_4092,N_5163);
nor U7770 (N_7770,N_3859,N_5055);
nand U7771 (N_7771,N_4519,N_5598);
nor U7772 (N_7772,N_5094,N_4496);
nand U7773 (N_7773,N_3077,N_5682);
nor U7774 (N_7774,N_4904,N_3856);
nand U7775 (N_7775,N_3277,N_5517);
or U7776 (N_7776,N_5078,N_3068);
nand U7777 (N_7777,N_4911,N_3822);
and U7778 (N_7778,N_4705,N_5549);
nor U7779 (N_7779,N_4311,N_5824);
nand U7780 (N_7780,N_5567,N_5658);
nand U7781 (N_7781,N_5328,N_5589);
and U7782 (N_7782,N_5704,N_4550);
nor U7783 (N_7783,N_5886,N_4002);
nand U7784 (N_7784,N_3882,N_3129);
and U7785 (N_7785,N_5033,N_3028);
nor U7786 (N_7786,N_4763,N_3369);
nor U7787 (N_7787,N_3496,N_5138);
and U7788 (N_7788,N_4133,N_5722);
and U7789 (N_7789,N_4336,N_5411);
nand U7790 (N_7790,N_4324,N_5806);
nor U7791 (N_7791,N_3844,N_3721);
and U7792 (N_7792,N_3940,N_3029);
nand U7793 (N_7793,N_3161,N_3542);
nand U7794 (N_7794,N_3532,N_4376);
nor U7795 (N_7795,N_5269,N_4376);
nand U7796 (N_7796,N_3789,N_5714);
nand U7797 (N_7797,N_4360,N_3847);
and U7798 (N_7798,N_5182,N_3551);
nor U7799 (N_7799,N_3168,N_4819);
xnor U7800 (N_7800,N_3190,N_4370);
and U7801 (N_7801,N_4851,N_3240);
and U7802 (N_7802,N_3693,N_4971);
and U7803 (N_7803,N_5759,N_4149);
and U7804 (N_7804,N_4756,N_3211);
nor U7805 (N_7805,N_5863,N_3149);
or U7806 (N_7806,N_5146,N_5717);
nand U7807 (N_7807,N_5081,N_4151);
nand U7808 (N_7808,N_5947,N_3535);
nand U7809 (N_7809,N_3305,N_3005);
nand U7810 (N_7810,N_3448,N_5322);
and U7811 (N_7811,N_4474,N_4060);
nand U7812 (N_7812,N_3476,N_4386);
and U7813 (N_7813,N_4127,N_3919);
or U7814 (N_7814,N_3316,N_3694);
or U7815 (N_7815,N_5543,N_4042);
or U7816 (N_7816,N_4156,N_5659);
and U7817 (N_7817,N_3196,N_4172);
nor U7818 (N_7818,N_4134,N_3495);
or U7819 (N_7819,N_5884,N_5132);
or U7820 (N_7820,N_4164,N_4298);
nand U7821 (N_7821,N_5707,N_4189);
or U7822 (N_7822,N_5325,N_3109);
nand U7823 (N_7823,N_4126,N_3375);
or U7824 (N_7824,N_4326,N_3393);
nor U7825 (N_7825,N_4696,N_5890);
nand U7826 (N_7826,N_5608,N_3811);
nand U7827 (N_7827,N_4670,N_4542);
nor U7828 (N_7828,N_3253,N_5181);
and U7829 (N_7829,N_5275,N_5870);
or U7830 (N_7830,N_5603,N_5056);
or U7831 (N_7831,N_4719,N_4948);
nand U7832 (N_7832,N_3442,N_3132);
and U7833 (N_7833,N_3978,N_4509);
and U7834 (N_7834,N_4566,N_5818);
nor U7835 (N_7835,N_5431,N_3594);
and U7836 (N_7836,N_4929,N_4789);
and U7837 (N_7837,N_5360,N_5050);
or U7838 (N_7838,N_3324,N_4630);
nor U7839 (N_7839,N_3768,N_5061);
nor U7840 (N_7840,N_4189,N_3076);
or U7841 (N_7841,N_5435,N_3282);
nand U7842 (N_7842,N_4788,N_4824);
nor U7843 (N_7843,N_5954,N_4599);
nand U7844 (N_7844,N_3309,N_4004);
nor U7845 (N_7845,N_5877,N_4302);
or U7846 (N_7846,N_3829,N_3274);
and U7847 (N_7847,N_4824,N_5363);
nand U7848 (N_7848,N_3580,N_3308);
or U7849 (N_7849,N_4380,N_5709);
and U7850 (N_7850,N_5161,N_5040);
nand U7851 (N_7851,N_3240,N_4108);
nand U7852 (N_7852,N_5602,N_4110);
or U7853 (N_7853,N_5801,N_4138);
or U7854 (N_7854,N_3602,N_4528);
nand U7855 (N_7855,N_5904,N_5080);
and U7856 (N_7856,N_4310,N_3741);
and U7857 (N_7857,N_3765,N_3554);
and U7858 (N_7858,N_4154,N_4479);
or U7859 (N_7859,N_3038,N_4184);
nor U7860 (N_7860,N_3260,N_4629);
or U7861 (N_7861,N_4678,N_5135);
nand U7862 (N_7862,N_5341,N_3218);
and U7863 (N_7863,N_3578,N_3306);
or U7864 (N_7864,N_3848,N_4143);
xnor U7865 (N_7865,N_3572,N_4190);
nand U7866 (N_7866,N_4231,N_5842);
or U7867 (N_7867,N_3661,N_5095);
nand U7868 (N_7868,N_5947,N_3374);
or U7869 (N_7869,N_4323,N_4063);
nor U7870 (N_7870,N_4084,N_3875);
xnor U7871 (N_7871,N_5772,N_4636);
nand U7872 (N_7872,N_3149,N_5730);
or U7873 (N_7873,N_3356,N_5831);
and U7874 (N_7874,N_5774,N_4270);
or U7875 (N_7875,N_5935,N_4241);
nand U7876 (N_7876,N_3799,N_4895);
or U7877 (N_7877,N_5538,N_5070);
and U7878 (N_7878,N_5383,N_5834);
nor U7879 (N_7879,N_4883,N_4553);
or U7880 (N_7880,N_3838,N_5180);
nand U7881 (N_7881,N_5436,N_3986);
nor U7882 (N_7882,N_4662,N_4931);
or U7883 (N_7883,N_3020,N_4915);
nor U7884 (N_7884,N_3160,N_3726);
and U7885 (N_7885,N_5080,N_5855);
and U7886 (N_7886,N_3220,N_5058);
and U7887 (N_7887,N_4992,N_3647);
nand U7888 (N_7888,N_5481,N_4782);
or U7889 (N_7889,N_5638,N_4387);
nand U7890 (N_7890,N_4553,N_4965);
nor U7891 (N_7891,N_3480,N_5718);
and U7892 (N_7892,N_5147,N_5819);
and U7893 (N_7893,N_4878,N_5762);
nor U7894 (N_7894,N_4466,N_4821);
nor U7895 (N_7895,N_3302,N_5866);
and U7896 (N_7896,N_5756,N_5854);
nand U7897 (N_7897,N_5713,N_3736);
nor U7898 (N_7898,N_3724,N_3132);
nor U7899 (N_7899,N_5430,N_4056);
or U7900 (N_7900,N_3170,N_4616);
or U7901 (N_7901,N_4784,N_4392);
nor U7902 (N_7902,N_4360,N_5414);
nand U7903 (N_7903,N_3882,N_4321);
nand U7904 (N_7904,N_4019,N_3729);
nand U7905 (N_7905,N_5026,N_4231);
nor U7906 (N_7906,N_5748,N_4121);
nand U7907 (N_7907,N_4071,N_3555);
nand U7908 (N_7908,N_5639,N_4263);
nand U7909 (N_7909,N_3380,N_4322);
nor U7910 (N_7910,N_5791,N_4647);
and U7911 (N_7911,N_4669,N_5434);
nor U7912 (N_7912,N_5653,N_3107);
and U7913 (N_7913,N_5533,N_4577);
or U7914 (N_7914,N_3642,N_4723);
and U7915 (N_7915,N_5257,N_4621);
nor U7916 (N_7916,N_5062,N_5489);
nor U7917 (N_7917,N_5841,N_3578);
nor U7918 (N_7918,N_5109,N_4943);
nand U7919 (N_7919,N_3285,N_5964);
nor U7920 (N_7920,N_5191,N_5568);
nand U7921 (N_7921,N_3637,N_3680);
or U7922 (N_7922,N_5599,N_5726);
nand U7923 (N_7923,N_5407,N_5644);
or U7924 (N_7924,N_3295,N_4371);
nand U7925 (N_7925,N_5220,N_5424);
xnor U7926 (N_7926,N_4451,N_4926);
or U7927 (N_7927,N_3806,N_3583);
nor U7928 (N_7928,N_3014,N_3485);
nor U7929 (N_7929,N_3814,N_3788);
and U7930 (N_7930,N_3176,N_4765);
nand U7931 (N_7931,N_5684,N_4374);
or U7932 (N_7932,N_5468,N_3835);
nand U7933 (N_7933,N_3673,N_3695);
nand U7934 (N_7934,N_5123,N_5060);
and U7935 (N_7935,N_3903,N_5975);
and U7936 (N_7936,N_4267,N_5686);
and U7937 (N_7937,N_4658,N_5951);
and U7938 (N_7938,N_4924,N_3062);
or U7939 (N_7939,N_3585,N_3388);
or U7940 (N_7940,N_5674,N_4915);
or U7941 (N_7941,N_3489,N_4160);
xnor U7942 (N_7942,N_5494,N_3609);
nand U7943 (N_7943,N_5330,N_5209);
nand U7944 (N_7944,N_4923,N_5852);
nand U7945 (N_7945,N_5038,N_3131);
nand U7946 (N_7946,N_3440,N_4178);
nor U7947 (N_7947,N_5688,N_5557);
and U7948 (N_7948,N_5597,N_4859);
nand U7949 (N_7949,N_5337,N_3903);
nand U7950 (N_7950,N_4103,N_3262);
or U7951 (N_7951,N_5377,N_3870);
and U7952 (N_7952,N_3687,N_4091);
and U7953 (N_7953,N_4756,N_3139);
nand U7954 (N_7954,N_3563,N_3273);
nor U7955 (N_7955,N_4585,N_5221);
nor U7956 (N_7956,N_3654,N_3651);
and U7957 (N_7957,N_5132,N_5552);
or U7958 (N_7958,N_3610,N_5856);
or U7959 (N_7959,N_4589,N_3491);
nor U7960 (N_7960,N_3244,N_4404);
or U7961 (N_7961,N_5492,N_4465);
nand U7962 (N_7962,N_3186,N_5992);
nand U7963 (N_7963,N_3392,N_5883);
nor U7964 (N_7964,N_5890,N_3063);
nor U7965 (N_7965,N_5620,N_3742);
nor U7966 (N_7966,N_4915,N_3667);
or U7967 (N_7967,N_4332,N_4150);
or U7968 (N_7968,N_5265,N_5386);
xnor U7969 (N_7969,N_4965,N_3453);
nand U7970 (N_7970,N_4005,N_5931);
nor U7971 (N_7971,N_4658,N_3024);
and U7972 (N_7972,N_4643,N_3366);
or U7973 (N_7973,N_4685,N_3242);
or U7974 (N_7974,N_4239,N_3299);
nand U7975 (N_7975,N_3803,N_4911);
or U7976 (N_7976,N_3699,N_3635);
and U7977 (N_7977,N_3892,N_3661);
and U7978 (N_7978,N_5985,N_5288);
nor U7979 (N_7979,N_5349,N_4512);
nor U7980 (N_7980,N_3127,N_3120);
nor U7981 (N_7981,N_4065,N_5628);
and U7982 (N_7982,N_5007,N_5279);
or U7983 (N_7983,N_4359,N_4459);
nor U7984 (N_7984,N_4133,N_3259);
nor U7985 (N_7985,N_5357,N_4929);
nand U7986 (N_7986,N_4140,N_3044);
nand U7987 (N_7987,N_5584,N_5705);
and U7988 (N_7988,N_4781,N_3397);
or U7989 (N_7989,N_3440,N_4308);
and U7990 (N_7990,N_3017,N_3801);
and U7991 (N_7991,N_5637,N_4280);
or U7992 (N_7992,N_5212,N_4764);
nand U7993 (N_7993,N_5500,N_5423);
and U7994 (N_7994,N_5143,N_3859);
nand U7995 (N_7995,N_4066,N_3713);
and U7996 (N_7996,N_3964,N_3255);
and U7997 (N_7997,N_3778,N_3407);
or U7998 (N_7998,N_4468,N_4373);
nor U7999 (N_7999,N_4437,N_5917);
nor U8000 (N_8000,N_3460,N_4262);
nand U8001 (N_8001,N_3176,N_5606);
nand U8002 (N_8002,N_4646,N_5496);
nor U8003 (N_8003,N_4602,N_5827);
nor U8004 (N_8004,N_4498,N_4481);
and U8005 (N_8005,N_5060,N_3030);
or U8006 (N_8006,N_4338,N_3207);
or U8007 (N_8007,N_3362,N_3820);
nor U8008 (N_8008,N_3068,N_5936);
and U8009 (N_8009,N_4315,N_5825);
nor U8010 (N_8010,N_3270,N_4459);
or U8011 (N_8011,N_3045,N_4582);
and U8012 (N_8012,N_4261,N_4442);
nand U8013 (N_8013,N_3868,N_3279);
and U8014 (N_8014,N_5296,N_5040);
nor U8015 (N_8015,N_5171,N_3790);
or U8016 (N_8016,N_3534,N_4410);
or U8017 (N_8017,N_3868,N_3913);
nor U8018 (N_8018,N_4294,N_4805);
or U8019 (N_8019,N_4966,N_5586);
and U8020 (N_8020,N_3302,N_4729);
nor U8021 (N_8021,N_3021,N_4697);
or U8022 (N_8022,N_4811,N_3157);
nand U8023 (N_8023,N_3248,N_5902);
and U8024 (N_8024,N_3965,N_5804);
nor U8025 (N_8025,N_4196,N_5006);
nor U8026 (N_8026,N_5020,N_4497);
nor U8027 (N_8027,N_4233,N_5353);
nand U8028 (N_8028,N_4613,N_5558);
nand U8029 (N_8029,N_4969,N_5380);
nor U8030 (N_8030,N_5608,N_5068);
and U8031 (N_8031,N_5185,N_4976);
nor U8032 (N_8032,N_4200,N_3717);
nor U8033 (N_8033,N_3621,N_4546);
or U8034 (N_8034,N_4897,N_4447);
nor U8035 (N_8035,N_4289,N_5584);
nand U8036 (N_8036,N_5943,N_4536);
nor U8037 (N_8037,N_3902,N_4735);
nor U8038 (N_8038,N_4238,N_4802);
xnor U8039 (N_8039,N_5171,N_3596);
or U8040 (N_8040,N_3506,N_3945);
nand U8041 (N_8041,N_5581,N_3684);
nand U8042 (N_8042,N_3176,N_3199);
and U8043 (N_8043,N_4375,N_3993);
nand U8044 (N_8044,N_4939,N_4957);
nor U8045 (N_8045,N_3201,N_5317);
nand U8046 (N_8046,N_4621,N_5834);
or U8047 (N_8047,N_4600,N_3007);
nand U8048 (N_8048,N_4408,N_3831);
or U8049 (N_8049,N_3546,N_5421);
nor U8050 (N_8050,N_3892,N_4270);
nand U8051 (N_8051,N_4074,N_5772);
nand U8052 (N_8052,N_5680,N_3656);
nand U8053 (N_8053,N_4628,N_4046);
nand U8054 (N_8054,N_4518,N_5706);
xor U8055 (N_8055,N_4237,N_4649);
nand U8056 (N_8056,N_3341,N_5234);
nand U8057 (N_8057,N_3800,N_4485);
and U8058 (N_8058,N_4102,N_5264);
nor U8059 (N_8059,N_3399,N_5054);
or U8060 (N_8060,N_3681,N_4111);
and U8061 (N_8061,N_3774,N_5311);
and U8062 (N_8062,N_5315,N_5390);
nor U8063 (N_8063,N_5917,N_3314);
nand U8064 (N_8064,N_5261,N_5946);
nor U8065 (N_8065,N_4022,N_4420);
nor U8066 (N_8066,N_4902,N_4129);
nor U8067 (N_8067,N_4710,N_4178);
xnor U8068 (N_8068,N_4694,N_3627);
or U8069 (N_8069,N_5891,N_5744);
nand U8070 (N_8070,N_3889,N_3445);
nor U8071 (N_8071,N_3286,N_4943);
or U8072 (N_8072,N_4434,N_5076);
and U8073 (N_8073,N_4553,N_5048);
and U8074 (N_8074,N_3124,N_3444);
and U8075 (N_8075,N_5256,N_4014);
or U8076 (N_8076,N_4418,N_3753);
nand U8077 (N_8077,N_4360,N_5131);
nor U8078 (N_8078,N_5702,N_5991);
and U8079 (N_8079,N_3879,N_3282);
nand U8080 (N_8080,N_4187,N_3158);
nand U8081 (N_8081,N_3590,N_4046);
nor U8082 (N_8082,N_4703,N_4574);
nand U8083 (N_8083,N_5998,N_5310);
and U8084 (N_8084,N_4740,N_4988);
nor U8085 (N_8085,N_4771,N_5913);
nand U8086 (N_8086,N_4324,N_5659);
nand U8087 (N_8087,N_3775,N_3974);
nand U8088 (N_8088,N_5860,N_3991);
nand U8089 (N_8089,N_4015,N_3411);
and U8090 (N_8090,N_5357,N_4676);
and U8091 (N_8091,N_4982,N_3300);
nor U8092 (N_8092,N_3843,N_3414);
nand U8093 (N_8093,N_4691,N_4312);
or U8094 (N_8094,N_5839,N_4005);
nor U8095 (N_8095,N_4087,N_5444);
or U8096 (N_8096,N_3389,N_3689);
nor U8097 (N_8097,N_4493,N_5702);
nor U8098 (N_8098,N_3515,N_5759);
or U8099 (N_8099,N_3694,N_4154);
nand U8100 (N_8100,N_3405,N_5927);
nor U8101 (N_8101,N_3795,N_5742);
nor U8102 (N_8102,N_3916,N_4677);
or U8103 (N_8103,N_4000,N_5462);
nand U8104 (N_8104,N_3407,N_4325);
nand U8105 (N_8105,N_5978,N_4205);
or U8106 (N_8106,N_4882,N_4257);
nor U8107 (N_8107,N_4296,N_4843);
and U8108 (N_8108,N_3533,N_3369);
nor U8109 (N_8109,N_5351,N_5559);
and U8110 (N_8110,N_4082,N_4578);
nand U8111 (N_8111,N_3901,N_4450);
and U8112 (N_8112,N_3435,N_5590);
nand U8113 (N_8113,N_4240,N_4219);
nand U8114 (N_8114,N_4780,N_4503);
nor U8115 (N_8115,N_4706,N_3771);
and U8116 (N_8116,N_4041,N_3213);
and U8117 (N_8117,N_4877,N_3133);
nand U8118 (N_8118,N_5081,N_3548);
nand U8119 (N_8119,N_5544,N_5888);
and U8120 (N_8120,N_5758,N_3268);
nand U8121 (N_8121,N_5755,N_4283);
or U8122 (N_8122,N_5990,N_5438);
nand U8123 (N_8123,N_5916,N_4501);
or U8124 (N_8124,N_5258,N_4608);
and U8125 (N_8125,N_4120,N_4651);
nand U8126 (N_8126,N_5693,N_5112);
nand U8127 (N_8127,N_5045,N_3754);
or U8128 (N_8128,N_4648,N_5924);
or U8129 (N_8129,N_3388,N_5808);
and U8130 (N_8130,N_5500,N_4310);
nor U8131 (N_8131,N_5824,N_5105);
and U8132 (N_8132,N_3018,N_5536);
xor U8133 (N_8133,N_3446,N_4575);
nor U8134 (N_8134,N_3419,N_3626);
and U8135 (N_8135,N_5287,N_5861);
or U8136 (N_8136,N_3325,N_3501);
and U8137 (N_8137,N_4784,N_4684);
or U8138 (N_8138,N_3378,N_5990);
nor U8139 (N_8139,N_5280,N_4594);
nor U8140 (N_8140,N_3423,N_3721);
and U8141 (N_8141,N_5961,N_5945);
and U8142 (N_8142,N_5516,N_4572);
and U8143 (N_8143,N_4999,N_3380);
or U8144 (N_8144,N_3534,N_3830);
nor U8145 (N_8145,N_5466,N_5257);
and U8146 (N_8146,N_3699,N_5827);
nor U8147 (N_8147,N_5517,N_5462);
nand U8148 (N_8148,N_4541,N_3265);
and U8149 (N_8149,N_4464,N_5094);
and U8150 (N_8150,N_3051,N_3462);
nand U8151 (N_8151,N_3298,N_5460);
and U8152 (N_8152,N_5774,N_4433);
nand U8153 (N_8153,N_3317,N_5240);
nor U8154 (N_8154,N_5574,N_5144);
and U8155 (N_8155,N_4079,N_3704);
and U8156 (N_8156,N_3043,N_5716);
or U8157 (N_8157,N_3019,N_5318);
nor U8158 (N_8158,N_3805,N_5236);
and U8159 (N_8159,N_3222,N_4778);
or U8160 (N_8160,N_4712,N_3655);
or U8161 (N_8161,N_3090,N_4966);
or U8162 (N_8162,N_5115,N_3657);
xor U8163 (N_8163,N_5920,N_3077);
and U8164 (N_8164,N_3924,N_4460);
nand U8165 (N_8165,N_3520,N_5569);
nor U8166 (N_8166,N_4466,N_4230);
nand U8167 (N_8167,N_4884,N_5205);
or U8168 (N_8168,N_5918,N_4590);
nor U8169 (N_8169,N_5457,N_4150);
or U8170 (N_8170,N_5225,N_4783);
nand U8171 (N_8171,N_3948,N_3270);
nand U8172 (N_8172,N_3569,N_3251);
nor U8173 (N_8173,N_3828,N_4890);
or U8174 (N_8174,N_5925,N_3923);
and U8175 (N_8175,N_4797,N_5164);
nor U8176 (N_8176,N_3346,N_4098);
or U8177 (N_8177,N_4431,N_5032);
or U8178 (N_8178,N_5231,N_4546);
and U8179 (N_8179,N_3345,N_5269);
and U8180 (N_8180,N_4838,N_3369);
nor U8181 (N_8181,N_4172,N_3080);
nor U8182 (N_8182,N_3316,N_5652);
nand U8183 (N_8183,N_3163,N_3334);
xor U8184 (N_8184,N_4270,N_4230);
nand U8185 (N_8185,N_4519,N_5074);
nand U8186 (N_8186,N_5205,N_4732);
nand U8187 (N_8187,N_5770,N_4178);
and U8188 (N_8188,N_3860,N_5585);
nand U8189 (N_8189,N_5775,N_4066);
and U8190 (N_8190,N_4251,N_3495);
and U8191 (N_8191,N_4456,N_4973);
nor U8192 (N_8192,N_3386,N_5103);
and U8193 (N_8193,N_3507,N_3310);
or U8194 (N_8194,N_5376,N_3693);
and U8195 (N_8195,N_5783,N_3435);
xor U8196 (N_8196,N_5166,N_5825);
or U8197 (N_8197,N_4272,N_3064);
nor U8198 (N_8198,N_3186,N_4982);
or U8199 (N_8199,N_4862,N_5801);
nand U8200 (N_8200,N_5709,N_3178);
and U8201 (N_8201,N_4773,N_5854);
nand U8202 (N_8202,N_4270,N_4767);
and U8203 (N_8203,N_4344,N_4996);
and U8204 (N_8204,N_3709,N_3908);
nand U8205 (N_8205,N_4579,N_5109);
nor U8206 (N_8206,N_3402,N_5982);
or U8207 (N_8207,N_5073,N_5192);
or U8208 (N_8208,N_5241,N_4389);
or U8209 (N_8209,N_4562,N_4709);
and U8210 (N_8210,N_5696,N_4276);
xnor U8211 (N_8211,N_3705,N_5486);
or U8212 (N_8212,N_4668,N_3210);
and U8213 (N_8213,N_4977,N_5373);
nand U8214 (N_8214,N_4669,N_3272);
and U8215 (N_8215,N_3328,N_4081);
or U8216 (N_8216,N_5234,N_3972);
or U8217 (N_8217,N_4900,N_3845);
or U8218 (N_8218,N_3221,N_4491);
nand U8219 (N_8219,N_5287,N_3516);
and U8220 (N_8220,N_3772,N_4248);
and U8221 (N_8221,N_4907,N_5630);
nand U8222 (N_8222,N_4865,N_3506);
and U8223 (N_8223,N_5834,N_5503);
nor U8224 (N_8224,N_3194,N_5772);
and U8225 (N_8225,N_5991,N_5905);
or U8226 (N_8226,N_5424,N_4202);
nand U8227 (N_8227,N_3728,N_3611);
and U8228 (N_8228,N_5289,N_3978);
or U8229 (N_8229,N_4074,N_4592);
nor U8230 (N_8230,N_4971,N_3888);
nand U8231 (N_8231,N_5164,N_4242);
xnor U8232 (N_8232,N_4294,N_5906);
and U8233 (N_8233,N_4289,N_4733);
nand U8234 (N_8234,N_3549,N_3375);
and U8235 (N_8235,N_4153,N_5366);
nor U8236 (N_8236,N_4694,N_3989);
and U8237 (N_8237,N_4431,N_4148);
and U8238 (N_8238,N_5755,N_4981);
nor U8239 (N_8239,N_4963,N_5002);
or U8240 (N_8240,N_5072,N_5536);
and U8241 (N_8241,N_3374,N_3888);
and U8242 (N_8242,N_3364,N_4136);
nor U8243 (N_8243,N_5975,N_4644);
or U8244 (N_8244,N_3633,N_3800);
nand U8245 (N_8245,N_5464,N_3301);
and U8246 (N_8246,N_5326,N_4791);
and U8247 (N_8247,N_5590,N_4715);
or U8248 (N_8248,N_3467,N_4525);
nor U8249 (N_8249,N_5028,N_4025);
nor U8250 (N_8250,N_4674,N_3556);
nand U8251 (N_8251,N_3137,N_4225);
nor U8252 (N_8252,N_4288,N_5524);
and U8253 (N_8253,N_4747,N_4198);
and U8254 (N_8254,N_4819,N_3746);
and U8255 (N_8255,N_4469,N_3485);
or U8256 (N_8256,N_3310,N_3148);
or U8257 (N_8257,N_5887,N_3802);
and U8258 (N_8258,N_3347,N_5739);
nand U8259 (N_8259,N_4673,N_4187);
and U8260 (N_8260,N_5107,N_5648);
or U8261 (N_8261,N_3807,N_4466);
nand U8262 (N_8262,N_4263,N_3198);
and U8263 (N_8263,N_4719,N_4349);
nor U8264 (N_8264,N_3696,N_4915);
or U8265 (N_8265,N_5065,N_3867);
and U8266 (N_8266,N_3846,N_3431);
and U8267 (N_8267,N_3363,N_4735);
or U8268 (N_8268,N_5631,N_5472);
and U8269 (N_8269,N_3253,N_5520);
or U8270 (N_8270,N_5499,N_4455);
nand U8271 (N_8271,N_5596,N_4736);
or U8272 (N_8272,N_5222,N_4491);
nor U8273 (N_8273,N_3977,N_3026);
or U8274 (N_8274,N_4790,N_3471);
nor U8275 (N_8275,N_3708,N_4308);
nor U8276 (N_8276,N_4490,N_4751);
or U8277 (N_8277,N_4520,N_4449);
nand U8278 (N_8278,N_5796,N_3160);
nor U8279 (N_8279,N_5733,N_4611);
xnor U8280 (N_8280,N_4587,N_3243);
nor U8281 (N_8281,N_3004,N_3737);
nor U8282 (N_8282,N_4273,N_4961);
or U8283 (N_8283,N_5900,N_3604);
and U8284 (N_8284,N_3431,N_5562);
or U8285 (N_8285,N_4076,N_4932);
or U8286 (N_8286,N_3908,N_5769);
and U8287 (N_8287,N_3409,N_4856);
nor U8288 (N_8288,N_4590,N_3770);
or U8289 (N_8289,N_4596,N_5446);
and U8290 (N_8290,N_3190,N_3957);
nor U8291 (N_8291,N_4409,N_3934);
nor U8292 (N_8292,N_4436,N_3185);
or U8293 (N_8293,N_3015,N_4001);
nand U8294 (N_8294,N_4288,N_4918);
and U8295 (N_8295,N_4619,N_5162);
nand U8296 (N_8296,N_5336,N_4980);
nand U8297 (N_8297,N_4852,N_5993);
and U8298 (N_8298,N_5334,N_4157);
nor U8299 (N_8299,N_5855,N_4961);
or U8300 (N_8300,N_5581,N_3857);
and U8301 (N_8301,N_4548,N_3612);
and U8302 (N_8302,N_5987,N_3871);
and U8303 (N_8303,N_5131,N_4666);
nand U8304 (N_8304,N_3612,N_4058);
nand U8305 (N_8305,N_4386,N_4975);
or U8306 (N_8306,N_4203,N_4185);
nor U8307 (N_8307,N_3580,N_5653);
nand U8308 (N_8308,N_5320,N_3726);
and U8309 (N_8309,N_3123,N_3437);
nand U8310 (N_8310,N_4824,N_4675);
nor U8311 (N_8311,N_3475,N_4773);
nor U8312 (N_8312,N_3047,N_3560);
nand U8313 (N_8313,N_4021,N_5521);
or U8314 (N_8314,N_5691,N_3668);
nor U8315 (N_8315,N_3638,N_5505);
nor U8316 (N_8316,N_3734,N_3345);
or U8317 (N_8317,N_3089,N_3274);
nor U8318 (N_8318,N_4839,N_5031);
nand U8319 (N_8319,N_5634,N_4713);
nor U8320 (N_8320,N_4759,N_5378);
nor U8321 (N_8321,N_3132,N_4107);
nor U8322 (N_8322,N_4554,N_3509);
nor U8323 (N_8323,N_5046,N_4945);
nand U8324 (N_8324,N_3641,N_5992);
nor U8325 (N_8325,N_4365,N_3317);
nor U8326 (N_8326,N_5121,N_3513);
or U8327 (N_8327,N_5658,N_4909);
and U8328 (N_8328,N_4675,N_4473);
and U8329 (N_8329,N_5507,N_5264);
and U8330 (N_8330,N_3561,N_4707);
nand U8331 (N_8331,N_3465,N_4322);
or U8332 (N_8332,N_5174,N_3974);
or U8333 (N_8333,N_5862,N_5735);
or U8334 (N_8334,N_3415,N_4218);
and U8335 (N_8335,N_4533,N_3404);
nor U8336 (N_8336,N_3566,N_3249);
and U8337 (N_8337,N_3003,N_5524);
and U8338 (N_8338,N_4751,N_4326);
or U8339 (N_8339,N_5535,N_4776);
or U8340 (N_8340,N_5476,N_4594);
or U8341 (N_8341,N_5006,N_4521);
and U8342 (N_8342,N_4520,N_5078);
nor U8343 (N_8343,N_5958,N_5159);
nor U8344 (N_8344,N_5482,N_5684);
nand U8345 (N_8345,N_4181,N_3428);
nor U8346 (N_8346,N_5230,N_3791);
or U8347 (N_8347,N_5446,N_3939);
nand U8348 (N_8348,N_4942,N_4959);
nand U8349 (N_8349,N_4116,N_4247);
nor U8350 (N_8350,N_5283,N_5434);
or U8351 (N_8351,N_3278,N_3338);
nand U8352 (N_8352,N_5070,N_3371);
nand U8353 (N_8353,N_3154,N_5072);
nor U8354 (N_8354,N_4005,N_4202);
or U8355 (N_8355,N_4633,N_4723);
nor U8356 (N_8356,N_5486,N_4181);
or U8357 (N_8357,N_3021,N_3605);
nor U8358 (N_8358,N_5794,N_4249);
nand U8359 (N_8359,N_5897,N_5269);
nand U8360 (N_8360,N_3457,N_3213);
or U8361 (N_8361,N_4718,N_3465);
or U8362 (N_8362,N_5347,N_4343);
and U8363 (N_8363,N_3265,N_4036);
and U8364 (N_8364,N_5517,N_3619);
and U8365 (N_8365,N_5442,N_4757);
and U8366 (N_8366,N_4863,N_3939);
nor U8367 (N_8367,N_4212,N_3152);
and U8368 (N_8368,N_5217,N_4744);
nand U8369 (N_8369,N_3731,N_3296);
nand U8370 (N_8370,N_5516,N_4302);
or U8371 (N_8371,N_5365,N_3461);
nor U8372 (N_8372,N_4180,N_3807);
nor U8373 (N_8373,N_4192,N_4228);
nand U8374 (N_8374,N_4804,N_4968);
and U8375 (N_8375,N_4262,N_4043);
nand U8376 (N_8376,N_4968,N_5601);
nand U8377 (N_8377,N_5616,N_3797);
nand U8378 (N_8378,N_4937,N_5818);
and U8379 (N_8379,N_3292,N_4217);
nor U8380 (N_8380,N_4142,N_3185);
or U8381 (N_8381,N_3958,N_3242);
and U8382 (N_8382,N_5629,N_5913);
nand U8383 (N_8383,N_5108,N_3690);
or U8384 (N_8384,N_5366,N_5239);
and U8385 (N_8385,N_3958,N_3496);
nand U8386 (N_8386,N_3000,N_4937);
nand U8387 (N_8387,N_5557,N_4840);
nand U8388 (N_8388,N_5232,N_4977);
nand U8389 (N_8389,N_4853,N_5721);
and U8390 (N_8390,N_3404,N_3108);
and U8391 (N_8391,N_3571,N_5014);
nand U8392 (N_8392,N_3713,N_4789);
nand U8393 (N_8393,N_3864,N_4112);
nand U8394 (N_8394,N_5985,N_5697);
nor U8395 (N_8395,N_5945,N_4605);
or U8396 (N_8396,N_5914,N_4543);
and U8397 (N_8397,N_3519,N_4137);
or U8398 (N_8398,N_3733,N_4973);
or U8399 (N_8399,N_4074,N_4644);
and U8400 (N_8400,N_3270,N_4973);
nor U8401 (N_8401,N_5223,N_4790);
nor U8402 (N_8402,N_4731,N_5156);
or U8403 (N_8403,N_4792,N_5982);
xnor U8404 (N_8404,N_4334,N_5563);
or U8405 (N_8405,N_4457,N_4822);
xnor U8406 (N_8406,N_3001,N_3721);
or U8407 (N_8407,N_3313,N_3942);
nand U8408 (N_8408,N_4412,N_4409);
nor U8409 (N_8409,N_5071,N_3779);
and U8410 (N_8410,N_4732,N_5409);
nand U8411 (N_8411,N_4847,N_3527);
nand U8412 (N_8412,N_4958,N_3720);
nand U8413 (N_8413,N_3826,N_4572);
nand U8414 (N_8414,N_4264,N_5285);
and U8415 (N_8415,N_5384,N_3301);
and U8416 (N_8416,N_5486,N_5844);
or U8417 (N_8417,N_5396,N_3798);
nor U8418 (N_8418,N_3071,N_4056);
nand U8419 (N_8419,N_5028,N_4519);
nand U8420 (N_8420,N_5182,N_3652);
nand U8421 (N_8421,N_3545,N_3690);
nor U8422 (N_8422,N_5160,N_3913);
nor U8423 (N_8423,N_4225,N_3639);
or U8424 (N_8424,N_4094,N_5961);
nand U8425 (N_8425,N_3449,N_4148);
nand U8426 (N_8426,N_5704,N_3171);
and U8427 (N_8427,N_3228,N_4502);
or U8428 (N_8428,N_5145,N_4323);
nand U8429 (N_8429,N_4939,N_5996);
nand U8430 (N_8430,N_3718,N_5970);
and U8431 (N_8431,N_3066,N_4496);
xnor U8432 (N_8432,N_3768,N_3693);
and U8433 (N_8433,N_4287,N_4742);
nor U8434 (N_8434,N_5926,N_5125);
nand U8435 (N_8435,N_4533,N_5819);
nand U8436 (N_8436,N_5492,N_3585);
or U8437 (N_8437,N_5795,N_4022);
and U8438 (N_8438,N_3282,N_5341);
or U8439 (N_8439,N_4555,N_4269);
nand U8440 (N_8440,N_4700,N_5655);
and U8441 (N_8441,N_4265,N_3195);
nor U8442 (N_8442,N_5619,N_3027);
and U8443 (N_8443,N_4674,N_3803);
nor U8444 (N_8444,N_5621,N_3290);
nor U8445 (N_8445,N_3095,N_4763);
nand U8446 (N_8446,N_5732,N_4249);
or U8447 (N_8447,N_5001,N_4109);
or U8448 (N_8448,N_3019,N_3929);
and U8449 (N_8449,N_3432,N_4977);
and U8450 (N_8450,N_4914,N_3223);
or U8451 (N_8451,N_5545,N_4498);
nor U8452 (N_8452,N_3570,N_5311);
nand U8453 (N_8453,N_4818,N_4353);
nor U8454 (N_8454,N_3761,N_5993);
or U8455 (N_8455,N_4449,N_4437);
or U8456 (N_8456,N_4242,N_5253);
nand U8457 (N_8457,N_5601,N_5285);
or U8458 (N_8458,N_3440,N_5975);
or U8459 (N_8459,N_3198,N_4802);
or U8460 (N_8460,N_3104,N_3997);
nand U8461 (N_8461,N_5805,N_4939);
nor U8462 (N_8462,N_3537,N_5216);
and U8463 (N_8463,N_5856,N_4612);
nor U8464 (N_8464,N_3456,N_5618);
nor U8465 (N_8465,N_4886,N_3267);
nor U8466 (N_8466,N_3071,N_3770);
nand U8467 (N_8467,N_4993,N_3785);
nand U8468 (N_8468,N_5146,N_4885);
nor U8469 (N_8469,N_4895,N_5698);
or U8470 (N_8470,N_4382,N_4095);
or U8471 (N_8471,N_5999,N_3557);
nor U8472 (N_8472,N_4434,N_3763);
nand U8473 (N_8473,N_5031,N_4792);
nor U8474 (N_8474,N_5596,N_5611);
nor U8475 (N_8475,N_3951,N_3356);
nor U8476 (N_8476,N_3411,N_5805);
nor U8477 (N_8477,N_5093,N_3481);
and U8478 (N_8478,N_5156,N_4003);
and U8479 (N_8479,N_3281,N_5409);
nand U8480 (N_8480,N_3294,N_4372);
nor U8481 (N_8481,N_4050,N_5120);
nand U8482 (N_8482,N_5207,N_4710);
nand U8483 (N_8483,N_3042,N_5342);
nand U8484 (N_8484,N_5003,N_3181);
and U8485 (N_8485,N_3039,N_3468);
or U8486 (N_8486,N_3324,N_3348);
nor U8487 (N_8487,N_5738,N_3572);
or U8488 (N_8488,N_3136,N_4452);
or U8489 (N_8489,N_5905,N_5493);
nor U8490 (N_8490,N_5356,N_3459);
nand U8491 (N_8491,N_3595,N_3298);
nor U8492 (N_8492,N_5250,N_3108);
and U8493 (N_8493,N_3643,N_5354);
or U8494 (N_8494,N_5638,N_4839);
and U8495 (N_8495,N_3347,N_4235);
or U8496 (N_8496,N_3166,N_4859);
or U8497 (N_8497,N_4302,N_3902);
and U8498 (N_8498,N_4078,N_4182);
nor U8499 (N_8499,N_5308,N_3927);
nand U8500 (N_8500,N_4390,N_4180);
nand U8501 (N_8501,N_4942,N_4601);
nor U8502 (N_8502,N_4736,N_3331);
nand U8503 (N_8503,N_5132,N_5989);
nand U8504 (N_8504,N_3765,N_3321);
and U8505 (N_8505,N_3192,N_3931);
nor U8506 (N_8506,N_3917,N_4417);
nor U8507 (N_8507,N_4631,N_5691);
nor U8508 (N_8508,N_3943,N_3015);
and U8509 (N_8509,N_4274,N_3202);
nand U8510 (N_8510,N_4087,N_4167);
and U8511 (N_8511,N_4313,N_5405);
and U8512 (N_8512,N_3879,N_4199);
nand U8513 (N_8513,N_4229,N_4361);
nor U8514 (N_8514,N_5244,N_4313);
or U8515 (N_8515,N_3603,N_3371);
or U8516 (N_8516,N_4953,N_3179);
nor U8517 (N_8517,N_4029,N_3376);
nand U8518 (N_8518,N_3564,N_3614);
or U8519 (N_8519,N_3249,N_3599);
nand U8520 (N_8520,N_3494,N_5698);
nand U8521 (N_8521,N_3107,N_4754);
nor U8522 (N_8522,N_4461,N_5606);
and U8523 (N_8523,N_4567,N_3957);
and U8524 (N_8524,N_4322,N_5544);
and U8525 (N_8525,N_4828,N_5598);
and U8526 (N_8526,N_5159,N_3471);
and U8527 (N_8527,N_5318,N_3801);
nand U8528 (N_8528,N_4171,N_4632);
or U8529 (N_8529,N_5949,N_5001);
or U8530 (N_8530,N_5506,N_3723);
or U8531 (N_8531,N_5933,N_5785);
or U8532 (N_8532,N_3251,N_5028);
and U8533 (N_8533,N_3956,N_4332);
or U8534 (N_8534,N_5229,N_3538);
nand U8535 (N_8535,N_3423,N_3791);
nor U8536 (N_8536,N_5590,N_3066);
and U8537 (N_8537,N_3810,N_5412);
or U8538 (N_8538,N_3985,N_5679);
and U8539 (N_8539,N_3575,N_4981);
nand U8540 (N_8540,N_4987,N_3678);
and U8541 (N_8541,N_4277,N_3529);
and U8542 (N_8542,N_3306,N_4435);
and U8543 (N_8543,N_4971,N_4174);
and U8544 (N_8544,N_5804,N_4664);
and U8545 (N_8545,N_4367,N_3220);
nand U8546 (N_8546,N_3373,N_4209);
and U8547 (N_8547,N_4081,N_5027);
nor U8548 (N_8548,N_3044,N_3640);
nor U8549 (N_8549,N_3517,N_3289);
and U8550 (N_8550,N_4089,N_5640);
nand U8551 (N_8551,N_5725,N_3506);
or U8552 (N_8552,N_3758,N_3692);
and U8553 (N_8553,N_4263,N_4518);
or U8554 (N_8554,N_5374,N_5507);
nand U8555 (N_8555,N_5319,N_3482);
nor U8556 (N_8556,N_3310,N_4657);
nand U8557 (N_8557,N_3027,N_5245);
or U8558 (N_8558,N_4191,N_5576);
nor U8559 (N_8559,N_4797,N_3038);
nand U8560 (N_8560,N_4220,N_4885);
nand U8561 (N_8561,N_3834,N_5437);
nand U8562 (N_8562,N_3773,N_3260);
and U8563 (N_8563,N_3556,N_5277);
nand U8564 (N_8564,N_4221,N_5155);
or U8565 (N_8565,N_4629,N_5448);
and U8566 (N_8566,N_4086,N_4397);
or U8567 (N_8567,N_3795,N_4237);
nor U8568 (N_8568,N_3860,N_3755);
xor U8569 (N_8569,N_4278,N_4897);
xnor U8570 (N_8570,N_3312,N_5220);
nand U8571 (N_8571,N_5473,N_3383);
and U8572 (N_8572,N_4670,N_5167);
or U8573 (N_8573,N_3527,N_5738);
or U8574 (N_8574,N_5716,N_5238);
or U8575 (N_8575,N_4508,N_4117);
or U8576 (N_8576,N_4377,N_4932);
and U8577 (N_8577,N_5848,N_4460);
and U8578 (N_8578,N_3018,N_5391);
and U8579 (N_8579,N_4716,N_5195);
nor U8580 (N_8580,N_3082,N_3973);
nor U8581 (N_8581,N_3954,N_3557);
nand U8582 (N_8582,N_5930,N_4238);
or U8583 (N_8583,N_3422,N_3293);
and U8584 (N_8584,N_4739,N_5273);
nand U8585 (N_8585,N_4659,N_3888);
or U8586 (N_8586,N_4460,N_4571);
or U8587 (N_8587,N_4219,N_3112);
or U8588 (N_8588,N_4593,N_4961);
and U8589 (N_8589,N_4442,N_3134);
or U8590 (N_8590,N_5853,N_3163);
nand U8591 (N_8591,N_5566,N_3696);
xnor U8592 (N_8592,N_3327,N_5846);
nand U8593 (N_8593,N_3972,N_4073);
and U8594 (N_8594,N_5097,N_3516);
nand U8595 (N_8595,N_5414,N_5652);
nand U8596 (N_8596,N_5322,N_3835);
nand U8597 (N_8597,N_5454,N_4774);
or U8598 (N_8598,N_3193,N_5495);
or U8599 (N_8599,N_5906,N_3410);
and U8600 (N_8600,N_3974,N_4947);
or U8601 (N_8601,N_3780,N_4907);
or U8602 (N_8602,N_4425,N_3697);
nor U8603 (N_8603,N_3072,N_3810);
nor U8604 (N_8604,N_3778,N_3907);
nand U8605 (N_8605,N_5516,N_5072);
and U8606 (N_8606,N_4194,N_3662);
nor U8607 (N_8607,N_4817,N_3212);
or U8608 (N_8608,N_5019,N_4283);
and U8609 (N_8609,N_4137,N_5567);
or U8610 (N_8610,N_4376,N_4107);
or U8611 (N_8611,N_5113,N_4307);
and U8612 (N_8612,N_4265,N_4477);
or U8613 (N_8613,N_4422,N_5477);
nor U8614 (N_8614,N_4025,N_4003);
nand U8615 (N_8615,N_4181,N_5871);
nand U8616 (N_8616,N_3017,N_5006);
and U8617 (N_8617,N_4176,N_4842);
nand U8618 (N_8618,N_4542,N_3421);
or U8619 (N_8619,N_3200,N_5668);
and U8620 (N_8620,N_3459,N_4440);
and U8621 (N_8621,N_5144,N_3601);
and U8622 (N_8622,N_5238,N_3581);
nand U8623 (N_8623,N_5680,N_4006);
and U8624 (N_8624,N_3948,N_4191);
nor U8625 (N_8625,N_3607,N_5076);
nor U8626 (N_8626,N_4349,N_3620);
and U8627 (N_8627,N_5746,N_4356);
or U8628 (N_8628,N_3954,N_4933);
nor U8629 (N_8629,N_3879,N_4556);
and U8630 (N_8630,N_5947,N_3112);
nand U8631 (N_8631,N_3619,N_4308);
nand U8632 (N_8632,N_3927,N_3675);
nor U8633 (N_8633,N_5696,N_3939);
or U8634 (N_8634,N_5975,N_3111);
nor U8635 (N_8635,N_3778,N_3570);
nor U8636 (N_8636,N_5811,N_3995);
and U8637 (N_8637,N_4887,N_5741);
nor U8638 (N_8638,N_4537,N_3728);
or U8639 (N_8639,N_5235,N_4266);
or U8640 (N_8640,N_4650,N_4143);
nor U8641 (N_8641,N_3624,N_3087);
nand U8642 (N_8642,N_3636,N_4902);
nor U8643 (N_8643,N_5923,N_4613);
and U8644 (N_8644,N_3440,N_5627);
and U8645 (N_8645,N_5910,N_5418);
and U8646 (N_8646,N_3867,N_4412);
and U8647 (N_8647,N_5602,N_4674);
nand U8648 (N_8648,N_5393,N_4699);
nor U8649 (N_8649,N_5533,N_3054);
or U8650 (N_8650,N_3651,N_4579);
nor U8651 (N_8651,N_4351,N_5655);
nand U8652 (N_8652,N_3501,N_3955);
nor U8653 (N_8653,N_4299,N_3958);
nand U8654 (N_8654,N_4135,N_4895);
or U8655 (N_8655,N_5524,N_5405);
nor U8656 (N_8656,N_3349,N_4142);
or U8657 (N_8657,N_4202,N_5755);
nand U8658 (N_8658,N_5784,N_3914);
or U8659 (N_8659,N_5755,N_3269);
nor U8660 (N_8660,N_4821,N_4783);
nor U8661 (N_8661,N_5491,N_4300);
and U8662 (N_8662,N_4644,N_3039);
nand U8663 (N_8663,N_4577,N_3075);
nor U8664 (N_8664,N_5950,N_5967);
or U8665 (N_8665,N_5605,N_3184);
nand U8666 (N_8666,N_3655,N_5003);
and U8667 (N_8667,N_5780,N_3138);
nand U8668 (N_8668,N_5267,N_4875);
and U8669 (N_8669,N_3022,N_3231);
nor U8670 (N_8670,N_4543,N_5846);
and U8671 (N_8671,N_4170,N_4879);
nand U8672 (N_8672,N_4632,N_5950);
or U8673 (N_8673,N_3392,N_3863);
and U8674 (N_8674,N_3108,N_3501);
nor U8675 (N_8675,N_5725,N_4708);
or U8676 (N_8676,N_4803,N_3111);
nand U8677 (N_8677,N_5545,N_3068);
nand U8678 (N_8678,N_3904,N_3917);
and U8679 (N_8679,N_3609,N_5139);
or U8680 (N_8680,N_5428,N_5192);
nor U8681 (N_8681,N_3852,N_5108);
or U8682 (N_8682,N_4054,N_3440);
or U8683 (N_8683,N_4581,N_3935);
or U8684 (N_8684,N_5083,N_3765);
and U8685 (N_8685,N_5903,N_4448);
nor U8686 (N_8686,N_4274,N_3026);
nor U8687 (N_8687,N_5092,N_4301);
nand U8688 (N_8688,N_4374,N_4161);
or U8689 (N_8689,N_3909,N_5793);
nand U8690 (N_8690,N_3909,N_3107);
nand U8691 (N_8691,N_4304,N_4868);
nor U8692 (N_8692,N_3458,N_3731);
and U8693 (N_8693,N_5361,N_3179);
nor U8694 (N_8694,N_5455,N_3090);
and U8695 (N_8695,N_5296,N_5080);
or U8696 (N_8696,N_5358,N_4942);
nor U8697 (N_8697,N_4253,N_5395);
nand U8698 (N_8698,N_4452,N_4077);
xnor U8699 (N_8699,N_4085,N_4606);
nand U8700 (N_8700,N_3882,N_4396);
nor U8701 (N_8701,N_4015,N_4321);
nand U8702 (N_8702,N_3809,N_3600);
or U8703 (N_8703,N_3843,N_4727);
nor U8704 (N_8704,N_3126,N_3445);
or U8705 (N_8705,N_4955,N_5452);
and U8706 (N_8706,N_5301,N_5532);
and U8707 (N_8707,N_3319,N_5942);
nand U8708 (N_8708,N_5741,N_5443);
nor U8709 (N_8709,N_4671,N_4906);
nor U8710 (N_8710,N_5240,N_4508);
nand U8711 (N_8711,N_5586,N_5440);
or U8712 (N_8712,N_4061,N_5111);
nand U8713 (N_8713,N_5029,N_4927);
and U8714 (N_8714,N_5851,N_3917);
and U8715 (N_8715,N_3327,N_4531);
or U8716 (N_8716,N_4476,N_5504);
or U8717 (N_8717,N_4224,N_5331);
nor U8718 (N_8718,N_3251,N_4877);
or U8719 (N_8719,N_4434,N_5100);
nor U8720 (N_8720,N_4763,N_3143);
nand U8721 (N_8721,N_4336,N_4722);
or U8722 (N_8722,N_4226,N_5210);
or U8723 (N_8723,N_4422,N_4263);
nor U8724 (N_8724,N_5890,N_3675);
nor U8725 (N_8725,N_5678,N_4104);
and U8726 (N_8726,N_5543,N_5069);
and U8727 (N_8727,N_3483,N_5324);
nand U8728 (N_8728,N_4932,N_5989);
or U8729 (N_8729,N_3186,N_5556);
nand U8730 (N_8730,N_3562,N_3534);
and U8731 (N_8731,N_4732,N_5733);
or U8732 (N_8732,N_4355,N_4830);
or U8733 (N_8733,N_3590,N_3971);
nor U8734 (N_8734,N_3624,N_5088);
nand U8735 (N_8735,N_4547,N_5777);
and U8736 (N_8736,N_4948,N_5522);
or U8737 (N_8737,N_5368,N_3980);
or U8738 (N_8738,N_4245,N_3670);
nor U8739 (N_8739,N_3902,N_3750);
and U8740 (N_8740,N_5191,N_3066);
nand U8741 (N_8741,N_5518,N_4995);
or U8742 (N_8742,N_3510,N_4754);
nand U8743 (N_8743,N_4201,N_5073);
nor U8744 (N_8744,N_5927,N_3814);
and U8745 (N_8745,N_4987,N_4206);
nand U8746 (N_8746,N_3499,N_4301);
nor U8747 (N_8747,N_4713,N_5147);
nand U8748 (N_8748,N_4722,N_5804);
and U8749 (N_8749,N_3433,N_3955);
nand U8750 (N_8750,N_3160,N_4097);
and U8751 (N_8751,N_3851,N_5873);
and U8752 (N_8752,N_5221,N_3738);
nor U8753 (N_8753,N_5814,N_3629);
nor U8754 (N_8754,N_3879,N_5306);
or U8755 (N_8755,N_5214,N_3310);
or U8756 (N_8756,N_3932,N_4326);
and U8757 (N_8757,N_4223,N_5577);
and U8758 (N_8758,N_4061,N_4152);
nand U8759 (N_8759,N_4692,N_4730);
nand U8760 (N_8760,N_3508,N_5982);
or U8761 (N_8761,N_5580,N_4164);
or U8762 (N_8762,N_4220,N_4748);
nand U8763 (N_8763,N_5568,N_3892);
and U8764 (N_8764,N_3668,N_5637);
or U8765 (N_8765,N_4329,N_5262);
and U8766 (N_8766,N_3440,N_3305);
or U8767 (N_8767,N_3385,N_5596);
and U8768 (N_8768,N_3701,N_3098);
and U8769 (N_8769,N_5891,N_4700);
nor U8770 (N_8770,N_5538,N_3812);
nand U8771 (N_8771,N_3739,N_5757);
and U8772 (N_8772,N_5394,N_4879);
nand U8773 (N_8773,N_3931,N_3521);
or U8774 (N_8774,N_3823,N_4807);
and U8775 (N_8775,N_4903,N_4921);
nand U8776 (N_8776,N_4920,N_3415);
nor U8777 (N_8777,N_4354,N_4215);
nor U8778 (N_8778,N_3922,N_4478);
nor U8779 (N_8779,N_3112,N_5931);
and U8780 (N_8780,N_4447,N_4988);
nor U8781 (N_8781,N_5541,N_4252);
nor U8782 (N_8782,N_3713,N_3566);
and U8783 (N_8783,N_4269,N_4120);
nor U8784 (N_8784,N_4082,N_4754);
or U8785 (N_8785,N_3566,N_4874);
and U8786 (N_8786,N_3742,N_5482);
nand U8787 (N_8787,N_3386,N_5973);
nand U8788 (N_8788,N_3958,N_4506);
nor U8789 (N_8789,N_4475,N_5710);
and U8790 (N_8790,N_5329,N_3556);
and U8791 (N_8791,N_3078,N_5647);
nor U8792 (N_8792,N_4157,N_4385);
or U8793 (N_8793,N_3693,N_3268);
or U8794 (N_8794,N_4314,N_5789);
nand U8795 (N_8795,N_3954,N_4499);
nor U8796 (N_8796,N_5227,N_3066);
and U8797 (N_8797,N_4960,N_4817);
nand U8798 (N_8798,N_5171,N_5829);
and U8799 (N_8799,N_3009,N_4319);
or U8800 (N_8800,N_5824,N_5342);
or U8801 (N_8801,N_5956,N_5033);
nand U8802 (N_8802,N_4715,N_3452);
or U8803 (N_8803,N_5955,N_4644);
nor U8804 (N_8804,N_3454,N_4589);
and U8805 (N_8805,N_5801,N_5487);
nor U8806 (N_8806,N_4688,N_5900);
nand U8807 (N_8807,N_4188,N_3502);
or U8808 (N_8808,N_4917,N_4644);
or U8809 (N_8809,N_3301,N_3103);
nor U8810 (N_8810,N_5029,N_4806);
and U8811 (N_8811,N_4702,N_4369);
and U8812 (N_8812,N_4078,N_3072);
nand U8813 (N_8813,N_4055,N_4040);
and U8814 (N_8814,N_3245,N_4545);
nor U8815 (N_8815,N_5344,N_4761);
nand U8816 (N_8816,N_3114,N_3194);
or U8817 (N_8817,N_4917,N_4765);
and U8818 (N_8818,N_4707,N_5873);
nand U8819 (N_8819,N_4764,N_5116);
nor U8820 (N_8820,N_5552,N_3612);
nand U8821 (N_8821,N_3984,N_3740);
or U8822 (N_8822,N_3506,N_3858);
nand U8823 (N_8823,N_3035,N_5416);
or U8824 (N_8824,N_4458,N_3315);
nand U8825 (N_8825,N_4663,N_4873);
and U8826 (N_8826,N_5270,N_4709);
or U8827 (N_8827,N_4265,N_4370);
nor U8828 (N_8828,N_5409,N_4675);
or U8829 (N_8829,N_5809,N_5831);
nand U8830 (N_8830,N_3354,N_4689);
nor U8831 (N_8831,N_5237,N_4300);
nor U8832 (N_8832,N_3469,N_4302);
or U8833 (N_8833,N_4308,N_3535);
xor U8834 (N_8834,N_4889,N_3666);
or U8835 (N_8835,N_3382,N_5827);
nand U8836 (N_8836,N_5217,N_5631);
nand U8837 (N_8837,N_3448,N_5584);
or U8838 (N_8838,N_4954,N_5515);
or U8839 (N_8839,N_5087,N_3996);
nor U8840 (N_8840,N_3546,N_5553);
nor U8841 (N_8841,N_3856,N_5391);
nor U8842 (N_8842,N_5512,N_4430);
nor U8843 (N_8843,N_4522,N_3432);
or U8844 (N_8844,N_4057,N_5178);
nor U8845 (N_8845,N_3670,N_4434);
and U8846 (N_8846,N_4086,N_5134);
or U8847 (N_8847,N_3959,N_4480);
nand U8848 (N_8848,N_3256,N_4902);
and U8849 (N_8849,N_4427,N_3936);
or U8850 (N_8850,N_4312,N_3792);
nand U8851 (N_8851,N_3449,N_5502);
nor U8852 (N_8852,N_3392,N_4448);
nor U8853 (N_8853,N_3376,N_3399);
nor U8854 (N_8854,N_3519,N_5978);
xor U8855 (N_8855,N_3502,N_5958);
nand U8856 (N_8856,N_4943,N_5566);
or U8857 (N_8857,N_4030,N_4276);
nand U8858 (N_8858,N_4151,N_5146);
nand U8859 (N_8859,N_3561,N_3912);
nor U8860 (N_8860,N_4379,N_4303);
and U8861 (N_8861,N_5526,N_5696);
nand U8862 (N_8862,N_3181,N_4284);
or U8863 (N_8863,N_5369,N_3901);
and U8864 (N_8864,N_3868,N_3022);
or U8865 (N_8865,N_4057,N_5792);
or U8866 (N_8866,N_5005,N_4139);
or U8867 (N_8867,N_4613,N_5471);
or U8868 (N_8868,N_5387,N_3030);
nor U8869 (N_8869,N_4824,N_4012);
and U8870 (N_8870,N_3486,N_5738);
nand U8871 (N_8871,N_3537,N_3507);
and U8872 (N_8872,N_3146,N_5695);
or U8873 (N_8873,N_4238,N_4974);
nand U8874 (N_8874,N_4057,N_4849);
and U8875 (N_8875,N_3926,N_5353);
or U8876 (N_8876,N_3185,N_4914);
nor U8877 (N_8877,N_5052,N_3504);
nand U8878 (N_8878,N_4997,N_4705);
and U8879 (N_8879,N_5623,N_3062);
and U8880 (N_8880,N_4838,N_3055);
and U8881 (N_8881,N_5942,N_5367);
nor U8882 (N_8882,N_5240,N_3732);
or U8883 (N_8883,N_4755,N_4383);
nor U8884 (N_8884,N_5403,N_4027);
nor U8885 (N_8885,N_4939,N_5807);
and U8886 (N_8886,N_4909,N_5184);
nor U8887 (N_8887,N_5398,N_4010);
or U8888 (N_8888,N_3976,N_5627);
or U8889 (N_8889,N_3547,N_4539);
and U8890 (N_8890,N_5481,N_3459);
nand U8891 (N_8891,N_3497,N_3745);
nand U8892 (N_8892,N_3387,N_3509);
or U8893 (N_8893,N_3217,N_3283);
and U8894 (N_8894,N_4652,N_5390);
nand U8895 (N_8895,N_3188,N_5415);
or U8896 (N_8896,N_3584,N_3878);
or U8897 (N_8897,N_5555,N_3367);
or U8898 (N_8898,N_3951,N_5220);
nor U8899 (N_8899,N_5642,N_4629);
nand U8900 (N_8900,N_4553,N_4997);
and U8901 (N_8901,N_4459,N_5297);
or U8902 (N_8902,N_5360,N_4850);
nand U8903 (N_8903,N_3652,N_5743);
nor U8904 (N_8904,N_4788,N_5256);
nand U8905 (N_8905,N_3111,N_5958);
nand U8906 (N_8906,N_4497,N_5139);
nand U8907 (N_8907,N_5988,N_4507);
or U8908 (N_8908,N_4972,N_4776);
nand U8909 (N_8909,N_5662,N_4597);
and U8910 (N_8910,N_4476,N_5047);
and U8911 (N_8911,N_3253,N_5301);
or U8912 (N_8912,N_5538,N_5218);
nand U8913 (N_8913,N_5361,N_3021);
and U8914 (N_8914,N_5885,N_4336);
nor U8915 (N_8915,N_3596,N_4121);
nor U8916 (N_8916,N_3978,N_5074);
nor U8917 (N_8917,N_4256,N_3614);
or U8918 (N_8918,N_5231,N_4748);
and U8919 (N_8919,N_4981,N_3370);
nor U8920 (N_8920,N_3456,N_5448);
nor U8921 (N_8921,N_4664,N_3880);
nor U8922 (N_8922,N_4482,N_5066);
nand U8923 (N_8923,N_5790,N_5566);
nand U8924 (N_8924,N_3936,N_4474);
and U8925 (N_8925,N_4323,N_3053);
or U8926 (N_8926,N_4580,N_4815);
nand U8927 (N_8927,N_3828,N_4542);
nor U8928 (N_8928,N_5315,N_3701);
and U8929 (N_8929,N_4610,N_5328);
nand U8930 (N_8930,N_5080,N_3510);
and U8931 (N_8931,N_4640,N_3391);
and U8932 (N_8932,N_4147,N_3047);
nor U8933 (N_8933,N_3783,N_5943);
and U8934 (N_8934,N_5994,N_4550);
nand U8935 (N_8935,N_3178,N_4559);
and U8936 (N_8936,N_3837,N_5666);
and U8937 (N_8937,N_4034,N_3981);
xor U8938 (N_8938,N_3874,N_5992);
and U8939 (N_8939,N_3075,N_4361);
nor U8940 (N_8940,N_4060,N_3744);
nor U8941 (N_8941,N_3315,N_4365);
and U8942 (N_8942,N_3041,N_3503);
nand U8943 (N_8943,N_3685,N_3250);
nor U8944 (N_8944,N_4506,N_4422);
nand U8945 (N_8945,N_5341,N_5615);
and U8946 (N_8946,N_5925,N_4241);
or U8947 (N_8947,N_3784,N_4071);
nand U8948 (N_8948,N_4646,N_3892);
and U8949 (N_8949,N_4141,N_5053);
nand U8950 (N_8950,N_4179,N_3480);
nand U8951 (N_8951,N_5315,N_3553);
and U8952 (N_8952,N_5630,N_5287);
or U8953 (N_8953,N_4547,N_3292);
and U8954 (N_8954,N_3872,N_5364);
or U8955 (N_8955,N_3574,N_4577);
nand U8956 (N_8956,N_3634,N_4362);
nand U8957 (N_8957,N_5650,N_3220);
or U8958 (N_8958,N_5037,N_5263);
nand U8959 (N_8959,N_3936,N_4267);
nor U8960 (N_8960,N_4955,N_5400);
nor U8961 (N_8961,N_4073,N_3282);
nor U8962 (N_8962,N_5652,N_5356);
and U8963 (N_8963,N_5204,N_4754);
nand U8964 (N_8964,N_4756,N_4388);
or U8965 (N_8965,N_3835,N_4874);
nand U8966 (N_8966,N_5053,N_5293);
nor U8967 (N_8967,N_3309,N_4353);
xor U8968 (N_8968,N_3974,N_5807);
and U8969 (N_8969,N_4136,N_3764);
or U8970 (N_8970,N_5962,N_3433);
nor U8971 (N_8971,N_4475,N_3334);
nand U8972 (N_8972,N_3482,N_3796);
nand U8973 (N_8973,N_5330,N_5964);
nand U8974 (N_8974,N_3543,N_3130);
nand U8975 (N_8975,N_3459,N_3068);
nand U8976 (N_8976,N_3588,N_5606);
nand U8977 (N_8977,N_3194,N_3441);
nor U8978 (N_8978,N_5594,N_3197);
nand U8979 (N_8979,N_4361,N_4332);
and U8980 (N_8980,N_4822,N_4814);
or U8981 (N_8981,N_3707,N_5826);
and U8982 (N_8982,N_4995,N_5304);
and U8983 (N_8983,N_4306,N_5497);
nor U8984 (N_8984,N_3282,N_4791);
nor U8985 (N_8985,N_4348,N_3279);
or U8986 (N_8986,N_4947,N_3829);
nor U8987 (N_8987,N_5229,N_5897);
and U8988 (N_8988,N_3935,N_5037);
nand U8989 (N_8989,N_4493,N_4785);
nor U8990 (N_8990,N_3094,N_4432);
nor U8991 (N_8991,N_3966,N_3085);
nand U8992 (N_8992,N_4251,N_3262);
and U8993 (N_8993,N_4771,N_4742);
nor U8994 (N_8994,N_4034,N_3811);
nor U8995 (N_8995,N_4690,N_3256);
nor U8996 (N_8996,N_5457,N_4109);
and U8997 (N_8997,N_3468,N_4707);
or U8998 (N_8998,N_4338,N_3273);
or U8999 (N_8999,N_3299,N_4280);
or U9000 (N_9000,N_8801,N_7906);
nor U9001 (N_9001,N_8494,N_7168);
nor U9002 (N_9002,N_8479,N_8847);
and U9003 (N_9003,N_8246,N_7037);
and U9004 (N_9004,N_6267,N_8364);
nand U9005 (N_9005,N_6674,N_7172);
and U9006 (N_9006,N_8231,N_7363);
nor U9007 (N_9007,N_8922,N_7779);
nand U9008 (N_9008,N_8728,N_6838);
and U9009 (N_9009,N_6625,N_8022);
nor U9010 (N_9010,N_8785,N_6233);
or U9011 (N_9011,N_6333,N_6847);
or U9012 (N_9012,N_6091,N_8314);
nor U9013 (N_9013,N_8724,N_6957);
nand U9014 (N_9014,N_6893,N_6307);
or U9015 (N_9015,N_6594,N_8032);
or U9016 (N_9016,N_7744,N_8476);
or U9017 (N_9017,N_7153,N_7200);
nand U9018 (N_9018,N_8576,N_8733);
and U9019 (N_9019,N_8600,N_8218);
nor U9020 (N_9020,N_7235,N_6071);
nand U9021 (N_9021,N_7760,N_8828);
and U9022 (N_9022,N_8668,N_7033);
or U9023 (N_9023,N_8968,N_6533);
or U9024 (N_9024,N_8791,N_6523);
nor U9025 (N_9025,N_6705,N_6548);
nor U9026 (N_9026,N_8481,N_8347);
or U9027 (N_9027,N_6166,N_7508);
and U9028 (N_9028,N_6664,N_8512);
nor U9029 (N_9029,N_8508,N_6709);
nor U9030 (N_9030,N_6308,N_6413);
nor U9031 (N_9031,N_8607,N_7680);
and U9032 (N_9032,N_7739,N_8831);
or U9033 (N_9033,N_6849,N_7403);
or U9034 (N_9034,N_6854,N_7872);
or U9035 (N_9035,N_8836,N_7888);
and U9036 (N_9036,N_7978,N_8123);
or U9037 (N_9037,N_7649,N_8956);
or U9038 (N_9038,N_8362,N_6571);
nand U9039 (N_9039,N_6846,N_8160);
nand U9040 (N_9040,N_7790,N_7691);
or U9041 (N_9041,N_6842,N_8626);
or U9042 (N_9042,N_8421,N_8878);
nor U9043 (N_9043,N_6287,N_8061);
nand U9044 (N_9044,N_6062,N_6836);
nor U9045 (N_9045,N_8647,N_7938);
or U9046 (N_9046,N_8114,N_8569);
nor U9047 (N_9047,N_6131,N_7438);
nor U9048 (N_9048,N_8480,N_7459);
nand U9049 (N_9049,N_6098,N_6367);
nand U9050 (N_9050,N_7187,N_8864);
nand U9051 (N_9051,N_8112,N_8935);
or U9052 (N_9052,N_7936,N_6115);
nor U9053 (N_9053,N_8797,N_8192);
nand U9054 (N_9054,N_7297,N_7345);
or U9055 (N_9055,N_8154,N_6868);
or U9056 (N_9056,N_7823,N_7251);
nand U9057 (N_9057,N_8553,N_8853);
nor U9058 (N_9058,N_6791,N_6941);
and U9059 (N_9059,N_8542,N_8683);
or U9060 (N_9060,N_6147,N_7287);
and U9061 (N_9061,N_7848,N_6279);
nor U9062 (N_9062,N_8136,N_6919);
nor U9063 (N_9063,N_7442,N_6624);
nand U9064 (N_9064,N_7968,N_8820);
nand U9065 (N_9065,N_7282,N_8838);
and U9066 (N_9066,N_6695,N_7934);
nor U9067 (N_9067,N_8285,N_7053);
nor U9068 (N_9068,N_8610,N_8526);
and U9069 (N_9069,N_6271,N_7441);
nand U9070 (N_9070,N_7504,N_8675);
nand U9071 (N_9071,N_6574,N_8059);
and U9072 (N_9072,N_6046,N_6990);
nand U9073 (N_9073,N_8748,N_7723);
nand U9074 (N_9074,N_8560,N_8570);
nor U9075 (N_9075,N_8143,N_7565);
nand U9076 (N_9076,N_8884,N_7068);
or U9077 (N_9077,N_8450,N_6778);
or U9078 (N_9078,N_6207,N_6770);
or U9079 (N_9079,N_7801,N_7218);
nand U9080 (N_9080,N_8999,N_6237);
nand U9081 (N_9081,N_6702,N_8240);
nor U9082 (N_9082,N_8590,N_8409);
and U9083 (N_9083,N_6741,N_8776);
nand U9084 (N_9084,N_6812,N_8313);
nor U9085 (N_9085,N_7277,N_8097);
or U9086 (N_9086,N_7498,N_6627);
nand U9087 (N_9087,N_7636,N_7897);
nand U9088 (N_9088,N_7810,N_8445);
and U9089 (N_9089,N_7969,N_6690);
nand U9090 (N_9090,N_7675,N_7700);
nor U9091 (N_9091,N_8958,N_7556);
nand U9092 (N_9092,N_7077,N_6833);
or U9093 (N_9093,N_6539,N_8721);
or U9094 (N_9094,N_6334,N_6987);
nor U9095 (N_9095,N_7358,N_8266);
nand U9096 (N_9096,N_8158,N_7065);
nand U9097 (N_9097,N_8507,N_7820);
or U9098 (N_9098,N_8622,N_7221);
nand U9099 (N_9099,N_7176,N_6878);
and U9100 (N_9100,N_8419,N_8068);
and U9101 (N_9101,N_7650,N_7450);
and U9102 (N_9102,N_7866,N_6542);
nand U9103 (N_9103,N_8593,N_7547);
and U9104 (N_9104,N_8008,N_8810);
nor U9105 (N_9105,N_6560,N_7245);
nand U9106 (N_9106,N_8462,N_6633);
xor U9107 (N_9107,N_8981,N_6465);
nand U9108 (N_9108,N_6301,N_6455);
nand U9109 (N_9109,N_6953,N_6628);
or U9110 (N_9110,N_7023,N_6830);
nor U9111 (N_9111,N_7155,N_7603);
nand U9112 (N_9112,N_7063,N_6154);
or U9113 (N_9113,N_6970,N_6840);
and U9114 (N_9114,N_8094,N_8066);
or U9115 (N_9115,N_6164,N_8581);
or U9116 (N_9116,N_6003,N_7757);
nor U9117 (N_9117,N_8245,N_6583);
nor U9118 (N_9118,N_8414,N_6156);
and U9119 (N_9119,N_8306,N_6779);
and U9120 (N_9120,N_8972,N_6075);
and U9121 (N_9121,N_6584,N_8416);
and U9122 (N_9122,N_7849,N_7387);
nor U9123 (N_9123,N_7036,N_8894);
and U9124 (N_9124,N_8187,N_8660);
nand U9125 (N_9125,N_8729,N_6685);
nor U9126 (N_9126,N_8255,N_6640);
and U9127 (N_9127,N_6315,N_8045);
nand U9128 (N_9128,N_8317,N_8238);
nor U9129 (N_9129,N_7350,N_6110);
or U9130 (N_9130,N_7107,N_6614);
nor U9131 (N_9131,N_8121,N_7139);
or U9132 (N_9132,N_7856,N_7943);
or U9133 (N_9133,N_8264,N_7079);
xnor U9134 (N_9134,N_6924,N_6587);
nor U9135 (N_9135,N_8321,N_6545);
nor U9136 (N_9136,N_7612,N_6610);
and U9137 (N_9137,N_8354,N_8657);
or U9138 (N_9138,N_8439,N_8635);
nand U9139 (N_9139,N_8713,N_6328);
nor U9140 (N_9140,N_8215,N_8407);
or U9141 (N_9141,N_7602,N_7770);
nand U9142 (N_9142,N_6401,N_6802);
nand U9143 (N_9143,N_6950,N_8665);
nor U9144 (N_9144,N_8868,N_8965);
nand U9145 (N_9145,N_7806,N_7325);
nand U9146 (N_9146,N_6662,N_6932);
nor U9147 (N_9147,N_7886,N_6861);
or U9148 (N_9148,N_8440,N_8769);
nand U9149 (N_9149,N_6656,N_8562);
nand U9150 (N_9150,N_7331,N_6290);
or U9151 (N_9151,N_7473,N_8423);
and U9152 (N_9152,N_7073,N_8153);
or U9153 (N_9153,N_7539,N_8992);
or U9154 (N_9154,N_7726,N_7526);
and U9155 (N_9155,N_6458,N_8372);
nor U9156 (N_9156,N_6208,N_8488);
nand U9157 (N_9157,N_7286,N_7613);
nor U9158 (N_9158,N_8361,N_7323);
nand U9159 (N_9159,N_6261,N_7844);
or U9160 (N_9160,N_8628,N_7243);
or U9161 (N_9161,N_8188,N_7792);
and U9162 (N_9162,N_7029,N_8203);
nand U9163 (N_9163,N_8537,N_8710);
nand U9164 (N_9164,N_6439,N_6923);
nor U9165 (N_9165,N_7554,N_6805);
nand U9166 (N_9166,N_8544,N_7316);
and U9167 (N_9167,N_6198,N_6556);
or U9168 (N_9168,N_7907,N_7558);
and U9169 (N_9169,N_7732,N_7617);
nor U9170 (N_9170,N_6194,N_8244);
or U9171 (N_9171,N_6193,N_8208);
nor U9172 (N_9172,N_6012,N_7851);
or U9173 (N_9173,N_7428,N_6379);
and U9174 (N_9174,N_7719,N_7877);
nor U9175 (N_9175,N_8391,N_7151);
or U9176 (N_9176,N_6885,N_6965);
and U9177 (N_9177,N_8516,N_8596);
nor U9178 (N_9178,N_7382,N_6577);
nand U9179 (N_9179,N_6349,N_7163);
or U9180 (N_9180,N_6515,N_7256);
nor U9181 (N_9181,N_6117,N_7673);
nand U9182 (N_9182,N_7294,N_6289);
or U9183 (N_9183,N_7089,N_6719);
nor U9184 (N_9184,N_7572,N_6736);
and U9185 (N_9185,N_8222,N_7633);
nand U9186 (N_9186,N_6155,N_8014);
nor U9187 (N_9187,N_8455,N_8169);
or U9188 (N_9188,N_6394,N_7947);
or U9189 (N_9189,N_6371,N_8976);
and U9190 (N_9190,N_7413,N_6351);
nand U9191 (N_9191,N_7360,N_7571);
nand U9192 (N_9192,N_7229,N_7987);
and U9193 (N_9193,N_6771,N_8195);
nor U9194 (N_9194,N_6845,N_6517);
nand U9195 (N_9195,N_7206,N_7445);
or U9196 (N_9196,N_6378,N_7889);
and U9197 (N_9197,N_8661,N_7359);
nor U9198 (N_9198,N_7753,N_7878);
or U9199 (N_9199,N_7748,N_7192);
nor U9200 (N_9200,N_8278,N_6353);
nor U9201 (N_9201,N_8987,N_7665);
and U9202 (N_9202,N_6330,N_6390);
nor U9203 (N_9203,N_6943,N_6966);
and U9204 (N_9204,N_7560,N_6151);
or U9205 (N_9205,N_6241,N_6227);
nor U9206 (N_9206,N_7483,N_7505);
or U9207 (N_9207,N_7304,N_6858);
nor U9208 (N_9208,N_8275,N_7480);
and U9209 (N_9209,N_8583,N_6036);
and U9210 (N_9210,N_6139,N_6590);
nor U9211 (N_9211,N_6900,N_8989);
and U9212 (N_9212,N_8950,N_7787);
nand U9213 (N_9213,N_6268,N_7536);
nor U9214 (N_9214,N_7653,N_7836);
or U9215 (N_9215,N_8429,N_7573);
nor U9216 (N_9216,N_7431,N_6368);
or U9217 (N_9217,N_6650,N_6444);
nand U9218 (N_9218,N_6199,N_6347);
and U9219 (N_9219,N_6471,N_7531);
and U9220 (N_9220,N_8289,N_6558);
and U9221 (N_9221,N_6914,N_7466);
nand U9222 (N_9222,N_6165,N_8337);
nand U9223 (N_9223,N_6944,N_8457);
nor U9224 (N_9224,N_7123,N_8131);
or U9225 (N_9225,N_7171,N_8146);
nor U9226 (N_9226,N_6647,N_6031);
nand U9227 (N_9227,N_6224,N_8885);
or U9228 (N_9228,N_6171,N_6596);
nand U9229 (N_9229,N_8890,N_8308);
nor U9230 (N_9230,N_8210,N_6781);
nor U9231 (N_9231,N_6374,N_8305);
and U9232 (N_9232,N_8165,N_8252);
or U9233 (N_9233,N_6875,N_8028);
nor U9234 (N_9234,N_6936,N_8110);
and U9235 (N_9235,N_8869,N_8900);
or U9236 (N_9236,N_8650,N_7561);
nor U9237 (N_9237,N_6190,N_7534);
and U9238 (N_9238,N_7310,N_6903);
nor U9239 (N_9239,N_6230,N_6430);
and U9240 (N_9240,N_7425,N_6697);
and U9241 (N_9241,N_8216,N_8076);
nor U9242 (N_9242,N_7958,N_8638);
or U9243 (N_9243,N_7657,N_6000);
xnor U9244 (N_9244,N_8898,N_8379);
nand U9245 (N_9245,N_7692,N_6454);
nor U9246 (N_9246,N_8684,N_6554);
and U9247 (N_9247,N_6426,N_7610);
or U9248 (N_9248,N_6566,N_7231);
nand U9249 (N_9249,N_8918,N_7880);
or U9250 (N_9250,N_8053,N_7755);
nor U9251 (N_9251,N_8789,N_6145);
or U9252 (N_9252,N_7800,N_7831);
and U9253 (N_9253,N_8062,N_6293);
nand U9254 (N_9254,N_8856,N_8469);
nand U9255 (N_9255,N_8304,N_7273);
nand U9256 (N_9256,N_6658,N_8237);
nand U9257 (N_9257,N_8793,N_8738);
and U9258 (N_9258,N_8659,N_7411);
nand U9259 (N_9259,N_8707,N_7905);
nor U9260 (N_9260,N_6569,N_8730);
or U9261 (N_9261,N_6911,N_7254);
or U9262 (N_9262,N_8921,N_7362);
or U9263 (N_9263,N_7099,N_6255);
nor U9264 (N_9264,N_7608,N_8568);
nor U9265 (N_9265,N_6005,N_6797);
and U9266 (N_9266,N_7717,N_7392);
nor U9267 (N_9267,N_8257,N_6500);
or U9268 (N_9268,N_8830,N_8527);
nand U9269 (N_9269,N_7220,N_6129);
nor U9270 (N_9270,N_6019,N_6035);
nand U9271 (N_9271,N_7887,N_7516);
and U9272 (N_9272,N_7408,N_8572);
nand U9273 (N_9273,N_8943,N_6088);
nor U9274 (N_9274,N_7313,N_6921);
nor U9275 (N_9275,N_8848,N_6252);
nand U9276 (N_9276,N_7899,N_7095);
nor U9277 (N_9277,N_8515,N_8223);
nor U9278 (N_9278,N_6082,N_7930);
nand U9279 (N_9279,N_7419,N_6727);
nand U9280 (N_9280,N_7103,N_8552);
or U9281 (N_9281,N_7056,N_6704);
and U9282 (N_9282,N_6128,N_8452);
nand U9283 (N_9283,N_7058,N_7060);
nor U9284 (N_9284,N_8551,N_7807);
nand U9285 (N_9285,N_7860,N_8937);
nor U9286 (N_9286,N_6711,N_7365);
nand U9287 (N_9287,N_8201,N_7890);
and U9288 (N_9288,N_6435,N_8456);
or U9289 (N_9289,N_6244,N_7775);
nand U9290 (N_9290,N_7398,N_7942);
or U9291 (N_9291,N_6095,N_6079);
nand U9292 (N_9292,N_8103,N_6002);
nor U9293 (N_9293,N_7822,N_8430);
or U9294 (N_9294,N_6322,N_8938);
nor U9295 (N_9295,N_7224,N_8718);
nor U9296 (N_9296,N_6856,N_8545);
and U9297 (N_9297,N_8164,N_6639);
nand U9298 (N_9298,N_8895,N_7637);
or U9299 (N_9299,N_7071,N_8186);
nor U9300 (N_9300,N_7314,N_7903);
or U9301 (N_9301,N_6636,N_8566);
nor U9302 (N_9302,N_6559,N_7332);
nand U9303 (N_9303,N_6683,N_7551);
or U9304 (N_9304,N_7012,N_8915);
nor U9305 (N_9305,N_8087,N_7169);
nand U9306 (N_9306,N_8183,N_8385);
or U9307 (N_9307,N_7133,N_7335);
nand U9308 (N_9308,N_7664,N_8157);
nor U9309 (N_9309,N_7193,N_6366);
nand U9310 (N_9310,N_8587,N_6247);
nor U9311 (N_9311,N_7240,N_6060);
or U9312 (N_9312,N_6819,N_6714);
xnor U9313 (N_9313,N_6934,N_8389);
and U9314 (N_9314,N_6185,N_6420);
nand U9315 (N_9315,N_7743,N_6484);
nand U9316 (N_9316,N_8316,N_7179);
nor U9317 (N_9317,N_8287,N_7972);
and U9318 (N_9318,N_6703,N_6300);
nor U9319 (N_9319,N_6740,N_6160);
nor U9320 (N_9320,N_8107,N_6928);
nand U9321 (N_9321,N_6913,N_6872);
nand U9322 (N_9322,N_8178,N_6265);
or U9323 (N_9323,N_8444,N_7566);
and U9324 (N_9324,N_8861,N_7524);
and U9325 (N_9325,N_7919,N_8592);
nor U9326 (N_9326,N_8254,N_7926);
nand U9327 (N_9327,N_6310,N_7328);
nor U9328 (N_9328,N_7105,N_6687);
nor U9329 (N_9329,N_8705,N_7047);
or U9330 (N_9330,N_7656,N_8877);
nor U9331 (N_9331,N_7988,N_8725);
and U9332 (N_9332,N_8623,N_8067);
nor U9333 (N_9333,N_7763,N_8658);
nand U9334 (N_9334,N_7946,N_7783);
and U9335 (N_9335,N_7475,N_7085);
xor U9336 (N_9336,N_7658,N_8630);
and U9337 (N_9337,N_6930,N_7118);
or U9338 (N_9338,N_8001,N_7385);
nor U9339 (N_9339,N_8700,N_8799);
nand U9340 (N_9340,N_7396,N_8672);
and U9341 (N_9341,N_8980,N_7334);
xnor U9342 (N_9342,N_6058,N_8825);
or U9343 (N_9343,N_8502,N_8086);
nand U9344 (N_9344,N_7570,N_7094);
or U9345 (N_9345,N_7710,N_7850);
and U9346 (N_9346,N_6857,N_8465);
or U9347 (N_9347,N_6306,N_6203);
and U9348 (N_9348,N_7490,N_7709);
or U9349 (N_9349,N_7864,N_8072);
or U9350 (N_9350,N_6634,N_7016);
xnor U9351 (N_9351,N_8594,N_6931);
nand U9352 (N_9352,N_6294,N_8887);
nor U9353 (N_9353,N_8525,N_6197);
nand U9354 (N_9354,N_7101,N_8805);
nand U9355 (N_9355,N_7030,N_7042);
nor U9356 (N_9356,N_6281,N_8866);
nor U9357 (N_9357,N_6391,N_7814);
nand U9358 (N_9358,N_7552,N_7941);
nor U9359 (N_9359,N_8052,N_7548);
nand U9360 (N_9360,N_6651,N_7985);
nor U9361 (N_9361,N_8139,N_6761);
nor U9362 (N_9362,N_8147,N_6832);
nor U9363 (N_9363,N_8332,N_8905);
and U9364 (N_9364,N_7213,N_6278);
and U9365 (N_9365,N_6620,N_8099);
and U9366 (N_9366,N_7980,N_6971);
and U9367 (N_9367,N_8954,N_8152);
nor U9368 (N_9368,N_8106,N_8678);
or U9369 (N_9369,N_7130,N_8913);
nor U9370 (N_9370,N_6946,N_8944);
nand U9371 (N_9371,N_7045,N_7795);
nand U9372 (N_9372,N_7870,N_8338);
and U9373 (N_9373,N_8388,N_7302);
and U9374 (N_9374,N_6916,N_6059);
or U9375 (N_9375,N_7590,N_6862);
nor U9376 (N_9376,N_6654,N_6790);
or U9377 (N_9377,N_6667,N_6852);
or U9378 (N_9378,N_8605,N_6382);
nand U9379 (N_9379,N_7682,N_8751);
and U9380 (N_9380,N_8268,N_6958);
nor U9381 (N_9381,N_7429,N_7594);
nor U9382 (N_9382,N_8955,N_7769);
nand U9383 (N_9383,N_8875,N_6266);
nand U9384 (N_9384,N_6425,N_7935);
or U9385 (N_9385,N_7846,N_6381);
nand U9386 (N_9386,N_8876,N_6576);
nor U9387 (N_9387,N_7311,N_7076);
and U9388 (N_9388,N_6410,N_8132);
and U9389 (N_9389,N_6112,N_7443);
nor U9390 (N_9390,N_6406,N_6666);
or U9391 (N_9391,N_8617,N_7525);
and U9392 (N_9392,N_6085,N_7735);
nor U9393 (N_9393,N_6557,N_6803);
nor U9394 (N_9394,N_6442,N_6001);
and U9395 (N_9395,N_7996,N_6764);
nor U9396 (N_9396,N_7412,N_6758);
nand U9397 (N_9397,N_6416,N_8150);
and U9398 (N_9398,N_7303,N_8677);
or U9399 (N_9399,N_8324,N_8901);
and U9400 (N_9400,N_6905,N_7768);
nand U9401 (N_9401,N_7638,N_6179);
or U9402 (N_9402,N_8206,N_8100);
nand U9403 (N_9403,N_7745,N_7901);
nor U9404 (N_9404,N_8970,N_8571);
or U9405 (N_9405,N_8229,N_7322);
nor U9406 (N_9406,N_8902,N_6478);
or U9407 (N_9407,N_8396,N_6615);
and U9408 (N_9408,N_8564,N_6121);
nand U9409 (N_9409,N_6074,N_6008);
or U9410 (N_9410,N_6876,N_7916);
and U9411 (N_9411,N_6744,N_7492);
nand U9412 (N_9412,N_8674,N_6520);
nor U9413 (N_9413,N_8997,N_6671);
or U9414 (N_9414,N_8381,N_6772);
nand U9415 (N_9415,N_8503,N_8673);
nand U9416 (N_9416,N_8862,N_7344);
or U9417 (N_9417,N_7891,N_7262);
nor U9418 (N_9418,N_6344,N_6997);
nand U9419 (N_9419,N_6908,N_8620);
nand U9420 (N_9420,N_8543,N_7862);
or U9421 (N_9421,N_7456,N_8294);
nor U9422 (N_9422,N_7640,N_6320);
nand U9423 (N_9423,N_8835,N_7281);
or U9424 (N_9424,N_7977,N_8529);
or U9425 (N_9425,N_8418,N_8957);
or U9426 (N_9426,N_8370,N_6429);
nand U9427 (N_9427,N_7271,N_6204);
nor U9428 (N_9428,N_6562,N_6360);
nor U9429 (N_9429,N_8311,N_7198);
or U9430 (N_9430,N_7485,N_7290);
nor U9431 (N_9431,N_7788,N_7914);
or U9432 (N_9432,N_6167,N_6956);
or U9433 (N_9433,N_7832,N_7040);
nor U9434 (N_9434,N_7376,N_7289);
nor U9435 (N_9435,N_8239,N_7057);
or U9436 (N_9436,N_6039,N_6612);
nand U9437 (N_9437,N_8353,N_6525);
or U9438 (N_9438,N_7244,N_7388);
nand U9439 (N_9439,N_8148,N_7993);
and U9440 (N_9440,N_6468,N_6143);
or U9441 (N_9441,N_7024,N_8563);
nand U9442 (N_9442,N_7593,N_8971);
nand U9443 (N_9443,N_7353,N_7730);
nor U9444 (N_9444,N_6509,N_7537);
or U9445 (N_9445,N_8604,N_7315);
or U9446 (N_9446,N_7336,N_7232);
nand U9447 (N_9447,N_8843,N_7586);
nand U9448 (N_9448,N_8760,N_8889);
and U9449 (N_9449,N_6815,N_6906);
nor U9450 (N_9450,N_8631,N_6326);
or U9451 (N_9451,N_7246,N_6926);
nand U9452 (N_9452,N_8113,N_7904);
nor U9453 (N_9453,N_7370,N_6456);
or U9454 (N_9454,N_8767,N_7015);
nor U9455 (N_9455,N_8704,N_6105);
nand U9456 (N_9456,N_6635,N_7614);
and U9457 (N_9457,N_7180,N_7146);
and U9458 (N_9458,N_6829,N_6595);
or U9459 (N_9459,N_8404,N_7265);
nand U9460 (N_9460,N_8436,N_8649);
nand U9461 (N_9461,N_6531,N_8055);
nand U9462 (N_9462,N_6752,N_6737);
or U9463 (N_9463,N_8470,N_6445);
and U9464 (N_9464,N_7211,N_6214);
and U9465 (N_9465,N_8757,N_6572);
nor U9466 (N_9466,N_7309,N_7338);
or U9467 (N_9467,N_8702,N_7970);
nor U9468 (N_9468,N_7070,N_6891);
and U9469 (N_9469,N_6902,N_6086);
nor U9470 (N_9470,N_7909,N_8804);
and U9471 (N_9471,N_8790,N_7378);
nand U9472 (N_9472,N_7585,N_6159);
nand U9473 (N_9473,N_6952,N_8449);
or U9474 (N_9474,N_7166,N_6400);
and U9475 (N_9475,N_6041,N_8307);
nand U9476 (N_9476,N_6713,N_7685);
nand U9477 (N_9477,N_7312,N_7503);
nand U9478 (N_9478,N_6245,N_8888);
or U9479 (N_9479,N_7589,N_7575);
nand U9480 (N_9480,N_7611,N_7954);
nor U9481 (N_9481,N_8454,N_6132);
nor U9482 (N_9482,N_7839,N_7994);
or U9483 (N_9483,N_6487,N_7219);
or U9484 (N_9484,N_7207,N_6222);
nand U9485 (N_9485,N_6696,N_7357);
nor U9486 (N_9486,N_7659,N_8598);
and U9487 (N_9487,N_8845,N_7371);
nand U9488 (N_9488,N_8994,N_8366);
nor U9489 (N_9489,N_8079,N_7932);
and U9490 (N_9490,N_8122,N_6994);
or U9491 (N_9491,N_8927,N_8290);
nor U9492 (N_9492,N_6678,N_6124);
or U9493 (N_9493,N_6865,N_7161);
or U9494 (N_9494,N_6188,N_6220);
and U9495 (N_9495,N_7976,N_7722);
nor U9496 (N_9496,N_8069,N_8536);
and U9497 (N_9497,N_7546,N_7119);
nor U9498 (N_9498,N_7959,N_7000);
nor U9499 (N_9499,N_6898,N_8814);
and U9500 (N_9500,N_7631,N_7197);
or U9501 (N_9501,N_7025,N_6275);
and U9502 (N_9502,N_6755,N_7815);
or U9503 (N_9503,N_7789,N_8236);
or U9504 (N_9504,N_6481,N_6592);
nand U9505 (N_9505,N_8162,N_6339);
nor U9506 (N_9506,N_6116,N_7167);
and U9507 (N_9507,N_7170,N_7196);
and U9508 (N_9508,N_6681,N_6939);
and U9509 (N_9509,N_7829,N_6680);
and U9510 (N_9510,N_7293,N_7448);
and U9511 (N_9511,N_6774,N_8253);
and U9512 (N_9512,N_8669,N_7830);
nand U9513 (N_9513,N_8211,N_6134);
or U9514 (N_9514,N_7737,N_6701);
nand U9515 (N_9515,N_7216,N_6679);
or U9516 (N_9516,N_7410,N_6818);
nand U9517 (N_9517,N_7173,N_8010);
nand U9518 (N_9518,N_6092,N_8111);
nor U9519 (N_9519,N_8063,N_8258);
nor U9520 (N_9520,N_6228,N_8948);
and U9521 (N_9521,N_8523,N_6324);
or U9522 (N_9522,N_6766,N_7278);
xnor U9523 (N_9523,N_7518,N_6653);
nand U9524 (N_9524,N_7960,N_8618);
or U9525 (N_9525,N_8044,N_6530);
nand U9526 (N_9526,N_8340,N_8003);
or U9527 (N_9527,N_6354,N_8248);
nand U9528 (N_9528,N_8363,N_6253);
nand U9529 (N_9529,N_6835,N_8993);
nand U9530 (N_9530,N_7533,N_6446);
and U9531 (N_9531,N_8168,N_7502);
nand U9532 (N_9532,N_8006,N_7718);
or U9533 (N_9533,N_6609,N_7416);
or U9534 (N_9534,N_7896,N_8312);
and U9535 (N_9535,N_6518,N_6492);
or U9536 (N_9536,N_7600,N_8217);
or U9537 (N_9537,N_8482,N_6922);
nor U9538 (N_9538,N_7997,N_6473);
nand U9539 (N_9539,N_7797,N_7427);
or U9540 (N_9540,N_7446,N_6968);
nand U9541 (N_9541,N_6751,N_7944);
and U9542 (N_9542,N_7284,N_7714);
and U9543 (N_9543,N_6133,N_6338);
or U9544 (N_9544,N_6927,N_6969);
and U9545 (N_9545,N_6963,N_7435);
nand U9546 (N_9546,N_6886,N_8792);
and U9547 (N_9547,N_7423,N_8750);
and U9548 (N_9548,N_6249,N_7108);
nor U9549 (N_9549,N_8945,N_6948);
or U9550 (N_9550,N_6995,N_8517);
or U9551 (N_9551,N_6070,N_8772);
or U9552 (N_9552,N_8916,N_7406);
or U9553 (N_9553,N_7707,N_7424);
nor U9554 (N_9554,N_6106,N_7203);
nand U9555 (N_9555,N_6483,N_6209);
and U9556 (N_9556,N_8951,N_6397);
nand U9557 (N_9557,N_7974,N_6629);
nor U9558 (N_9558,N_7497,N_7132);
or U9559 (N_9559,N_6547,N_6168);
nor U9560 (N_9560,N_6361,N_8387);
nor U9561 (N_9561,N_6448,N_6340);
and U9562 (N_9562,N_7181,N_6161);
nand U9563 (N_9563,N_6887,N_8329);
xnor U9564 (N_9564,N_6282,N_8426);
or U9565 (N_9565,N_8842,N_6816);
or U9566 (N_9566,N_7937,N_7237);
nand U9567 (N_9567,N_6028,N_6644);
nand U9568 (N_9568,N_6050,N_7451);
or U9569 (N_9569,N_6659,N_8588);
or U9570 (N_9570,N_8051,N_7606);
nand U9571 (N_9571,N_6144,N_7186);
or U9572 (N_9572,N_6527,N_8612);
or U9573 (N_9573,N_8874,N_6718);
or U9574 (N_9574,N_8689,N_7910);
nand U9575 (N_9575,N_8739,N_8764);
and U9576 (N_9576,N_7472,N_6200);
nand U9577 (N_9577,N_8054,N_7746);
or U9578 (N_9578,N_8189,N_7569);
nor U9579 (N_9579,N_7306,N_7765);
and U9580 (N_9580,N_8412,N_7230);
nand U9581 (N_9581,N_7655,N_6153);
or U9582 (N_9582,N_6053,N_8393);
or U9583 (N_9583,N_8075,N_7622);
and U9584 (N_9584,N_6677,N_8325);
and U9585 (N_9585,N_7583,N_7545);
or U9586 (N_9586,N_6402,N_8011);
or U9587 (N_9587,N_6513,N_8382);
nand U9588 (N_9588,N_7017,N_7477);
nand U9589 (N_9589,N_8497,N_7728);
or U9590 (N_9590,N_8297,N_6649);
nand U9591 (N_9591,N_8358,N_6765);
or U9592 (N_9592,N_7495,N_7599);
or U9593 (N_9593,N_8602,N_7778);
or U9594 (N_9594,N_8130,N_6493);
nand U9595 (N_9595,N_7720,N_6206);
and U9596 (N_9596,N_7283,N_8643);
or U9597 (N_9597,N_7404,N_6603);
or U9598 (N_9598,N_6123,N_6196);
and U9599 (N_9599,N_8025,N_8039);
and U9600 (N_9600,N_8555,N_8342);
nor U9601 (N_9601,N_7268,N_7457);
nor U9602 (N_9602,N_8924,N_8173);
nand U9603 (N_9603,N_8198,N_7038);
nor U9604 (N_9604,N_6585,N_8749);
nand U9605 (N_9605,N_6866,N_7066);
or U9606 (N_9606,N_7791,N_7333);
and U9607 (N_9607,N_8904,N_8284);
and U9608 (N_9608,N_6920,N_7628);
nor U9609 (N_9609,N_7461,N_6336);
or U9610 (N_9610,N_6173,N_7014);
xor U9611 (N_9611,N_7449,N_7067);
and U9612 (N_9612,N_7212,N_7786);
and U9613 (N_9613,N_8941,N_8632);
or U9614 (N_9614,N_6480,N_6327);
nor U9615 (N_9615,N_8532,N_8891);
or U9616 (N_9616,N_6461,N_8547);
nand U9617 (N_9617,N_7803,N_6951);
or U9618 (N_9618,N_8015,N_7771);
nand U9619 (N_9619,N_8663,N_8124);
and U9620 (N_9620,N_6551,N_6672);
and U9621 (N_9621,N_8920,N_6728);
or U9622 (N_9622,N_6080,N_8013);
or U9623 (N_9623,N_7973,N_7845);
and U9624 (N_9624,N_8400,N_6489);
or U9625 (N_9625,N_7364,N_7701);
nand U9626 (N_9626,N_8318,N_6611);
and U9627 (N_9627,N_6384,N_6789);
nand U9628 (N_9628,N_6383,N_8586);
and U9629 (N_9629,N_7092,N_8758);
or U9630 (N_9630,N_7462,N_7124);
nand U9631 (N_9631,N_8690,N_7592);
and U9632 (N_9632,N_8019,N_7184);
nand U9633 (N_9633,N_6018,N_8490);
or U9634 (N_9634,N_6158,N_7384);
nand U9635 (N_9635,N_6229,N_6332);
nand U9636 (N_9636,N_7027,N_7267);
or U9637 (N_9637,N_8794,N_8899);
and U9638 (N_9638,N_8930,N_7553);
nand U9639 (N_9639,N_6463,N_7623);
nor U9640 (N_9640,N_8004,N_8694);
nand U9641 (N_9641,N_6021,N_7729);
or U9642 (N_9642,N_8267,N_7270);
and U9643 (N_9643,N_7007,N_7654);
nand U9644 (N_9644,N_8809,N_8759);
nor U9645 (N_9645,N_6169,N_6541);
nor U9646 (N_9646,N_8521,N_6984);
nor U9647 (N_9647,N_7918,N_8291);
nor U9648 (N_9648,N_8155,N_6482);
nor U9649 (N_9649,N_6749,N_8170);
nand U9650 (N_9650,N_8535,N_8403);
and U9651 (N_9651,N_6884,N_8172);
and U9652 (N_9652,N_8691,N_7135);
nor U9653 (N_9653,N_6844,N_7463);
or U9654 (N_9654,N_6386,N_7920);
and U9655 (N_9655,N_7296,N_8939);
nand U9656 (N_9656,N_7750,N_8235);
or U9657 (N_9657,N_7183,N_8870);
nand U9658 (N_9658,N_7952,N_8974);
or U9659 (N_9659,N_8380,N_6598);
nand U9660 (N_9660,N_6869,N_6689);
nand U9661 (N_9661,N_7596,N_7965);
nand U9662 (N_9662,N_7233,N_8686);
and U9663 (N_9663,N_8681,N_8269);
nand U9664 (N_9664,N_8609,N_8486);
nor U9665 (N_9665,N_8175,N_6180);
nor U9666 (N_9666,N_6304,N_8367);
nor U9667 (N_9667,N_8048,N_7493);
or U9668 (N_9668,N_8161,N_7215);
and U9669 (N_9669,N_6045,N_7838);
and U9670 (N_9670,N_6645,N_7439);
and U9671 (N_9671,N_7120,N_8091);
or U9672 (N_9672,N_6859,N_6638);
nand U9673 (N_9673,N_8762,N_6127);
nor U9674 (N_9674,N_7069,N_7339);
nor U9675 (N_9675,N_6880,N_6623);
nand U9676 (N_9676,N_7062,N_7715);
nand U9677 (N_9677,N_7489,N_8624);
or U9678 (N_9678,N_6083,N_7616);
or U9679 (N_9679,N_7308,N_8815);
and U9680 (N_9680,N_7032,N_7627);
and U9681 (N_9681,N_7367,N_7043);
nor U9682 (N_9682,N_7080,N_8860);
nand U9683 (N_9683,N_8967,N_7641);
nand U9684 (N_9684,N_7913,N_8907);
nand U9685 (N_9685,N_7247,N_8349);
nand U9686 (N_9686,N_7098,N_8300);
nand U9687 (N_9687,N_6896,N_8743);
nor U9688 (N_9688,N_7532,N_8256);
nand U9689 (N_9689,N_6004,N_6724);
nand U9690 (N_9690,N_6219,N_8043);
and U9691 (N_9691,N_7195,N_8402);
nor U9692 (N_9692,N_8723,N_8190);
nand U9693 (N_9693,N_7051,N_6350);
nor U9694 (N_9694,N_8280,N_6537);
nand U9695 (N_9695,N_8034,N_6682);
and U9696 (N_9696,N_8844,N_6423);
nor U9697 (N_9697,N_7228,N_6412);
nor U9698 (N_9698,N_6486,N_8652);
and U9699 (N_9699,N_6767,N_8331);
or U9700 (N_9700,N_6061,N_8082);
nor U9701 (N_9701,N_6375,N_6023);
nand U9702 (N_9702,N_7347,N_6785);
nor U9703 (N_9703,N_6256,N_7356);
nor U9704 (N_9704,N_7496,N_8667);
or U9705 (N_9705,N_6146,N_8030);
and U9706 (N_9706,N_7824,N_6210);
and U9707 (N_9707,N_6863,N_8448);
nand U9708 (N_9708,N_7506,N_8012);
nand U9709 (N_9709,N_8356,N_7827);
or U9710 (N_9710,N_8806,N_6068);
nor U9711 (N_9711,N_6260,N_8141);
and U9712 (N_9712,N_7134,N_7468);
or U9713 (N_9713,N_6404,N_7348);
nor U9714 (N_9714,N_8591,N_7194);
or U9715 (N_9715,N_6824,N_6619);
nand U9716 (N_9716,N_6469,N_6706);
or U9717 (N_9717,N_6798,N_6591);
or U9718 (N_9718,N_7933,N_7776);
and U9719 (N_9719,N_8947,N_7660);
nand U9720 (N_9720,N_8133,N_6396);
and U9721 (N_9721,N_8765,N_7305);
or U9722 (N_9722,N_8640,N_7758);
nand U9723 (N_9723,N_6213,N_6020);
nor U9724 (N_9724,N_6038,N_8666);
nor U9725 (N_9725,N_8855,N_8425);
nand U9726 (N_9726,N_7136,N_7401);
or U9727 (N_9727,N_7879,N_7164);
xor U9728 (N_9728,N_7005,N_6759);
nor U9729 (N_9729,N_6479,N_8384);
nand U9730 (N_9730,N_7259,N_8398);
nand U9731 (N_9731,N_7121,N_6177);
or U9732 (N_9732,N_6524,N_6700);
or U9733 (N_9733,N_8220,N_6034);
nand U9734 (N_9734,N_8101,N_7528);
or U9735 (N_9735,N_8906,N_7674);
nor U9736 (N_9736,N_8397,N_7529);
and U9737 (N_9737,N_6459,N_7989);
nand U9738 (N_9738,N_7847,N_8633);
nand U9739 (N_9739,N_6373,N_8437);
or U9740 (N_9740,N_6910,N_6511);
or U9741 (N_9741,N_6405,N_8653);
nand U9742 (N_9742,N_7676,N_8309);
or U9743 (N_9743,N_8641,N_7568);
nand U9744 (N_9744,N_7106,N_7559);
nor U9745 (N_9745,N_7458,N_6152);
or U9746 (N_9746,N_8849,N_7921);
or U9747 (N_9747,N_7704,N_6553);
and U9748 (N_9748,N_6292,N_8166);
and U9749 (N_9749,N_6311,N_6385);
nor U9750 (N_9750,N_7821,N_7520);
and U9751 (N_9751,N_6403,N_8625);
nand U9752 (N_9752,N_6894,N_8334);
or U9753 (N_9753,N_6436,N_7409);
or U9754 (N_9754,N_8163,N_6399);
nand U9755 (N_9755,N_6933,N_7867);
nand U9756 (N_9756,N_8579,N_8035);
nor U9757 (N_9757,N_8471,N_8606);
nor U9758 (N_9758,N_8474,N_8138);
or U9759 (N_9759,N_6904,N_6699);
nand U9760 (N_9760,N_6961,N_8786);
nor U9761 (N_9761,N_6432,N_6813);
or U9762 (N_9762,N_8619,N_6499);
xor U9763 (N_9763,N_6114,N_8156);
nor U9764 (N_9764,N_8319,N_7059);
and U9765 (N_9765,N_6621,N_6992);
nand U9766 (N_9766,N_7962,N_8251);
nand U9767 (N_9767,N_7266,N_6794);
nor U9768 (N_9768,N_7871,N_8811);
nand U9769 (N_9769,N_6355,N_7644);
nor U9770 (N_9770,N_8093,N_7634);
or U9771 (N_9771,N_6312,N_8645);
and U9772 (N_9772,N_6871,N_6398);
nand U9773 (N_9773,N_6119,N_8833);
nand U9774 (N_9774,N_7924,N_6746);
nor U9775 (N_9775,N_7054,N_6954);
and U9776 (N_9776,N_6626,N_8817);
or U9777 (N_9777,N_6335,N_6212);
or U9778 (N_9778,N_8292,N_6722);
nand U9779 (N_9779,N_6652,N_6890);
or U9780 (N_9780,N_6387,N_8886);
nand U9781 (N_9781,N_7494,N_7917);
nand U9782 (N_9782,N_7205,N_8693);
nor U9783 (N_9783,N_6181,N_7394);
and U9784 (N_9784,N_7953,N_7956);
or U9785 (N_9785,N_8813,N_7764);
and U9786 (N_9786,N_6467,N_7160);
nor U9787 (N_9787,N_8942,N_7581);
or U9788 (N_9788,N_6163,N_8024);
or U9789 (N_9789,N_6150,N_7109);
nor U9790 (N_9790,N_7111,N_6174);
nor U9791 (N_9791,N_8234,N_8282);
nand U9792 (N_9792,N_7869,N_7693);
or U9793 (N_9793,N_8227,N_6052);
nor U9794 (N_9794,N_7981,N_8346);
or U9795 (N_9795,N_7513,N_7400);
and U9796 (N_9796,N_8492,N_6176);
nand U9797 (N_9797,N_7686,N_6226);
or U9798 (N_9798,N_7541,N_7342);
or U9799 (N_9799,N_6365,N_6462);
and U9800 (N_9800,N_7318,N_6864);
and U9801 (N_9801,N_8046,N_6084);
nand U9802 (N_9802,N_7687,N_6508);
nor U9803 (N_9803,N_8696,N_8796);
nand U9804 (N_9804,N_8177,N_6895);
or U9805 (N_9805,N_8089,N_8982);
and U9806 (N_9806,N_8451,N_7579);
or U9807 (N_9807,N_7696,N_8088);
and U9808 (N_9808,N_8616,N_7434);
xor U9809 (N_9809,N_8042,N_7003);
or U9810 (N_9810,N_7618,N_6316);
nor U9811 (N_9811,N_7711,N_8298);
and U9812 (N_9812,N_8135,N_8197);
or U9813 (N_9813,N_8914,N_8839);
and U9814 (N_9814,N_6826,N_7467);
nor U9815 (N_9815,N_7740,N_8824);
or U9816 (N_9816,N_6768,N_7125);
or U9817 (N_9817,N_7544,N_8199);
or U9818 (N_9818,N_6889,N_7291);
nor U9819 (N_9819,N_6305,N_7835);
or U9820 (N_9820,N_7234,N_6991);
nor U9821 (N_9821,N_7258,N_7873);
or U9822 (N_9822,N_6285,N_6983);
nor U9823 (N_9823,N_8473,N_7639);
nor U9824 (N_9824,N_8466,N_8685);
nand U9825 (N_9825,N_6597,N_8383);
nor U9826 (N_9826,N_6357,N_8714);
nand U9827 (N_9827,N_6246,N_6535);
or U9828 (N_9828,N_8109,N_8611);
or U9829 (N_9829,N_7708,N_6135);
nor U9830 (N_9830,N_7582,N_8330);
nand U9831 (N_9831,N_6631,N_6747);
or U9832 (N_9832,N_6352,N_6066);
nand U9833 (N_9833,N_6142,N_8533);
nor U9834 (N_9834,N_6618,N_8080);
or U9835 (N_9835,N_7747,N_7114);
and U9836 (N_9836,N_6236,N_8908);
nor U9837 (N_9837,N_8040,N_7390);
and U9838 (N_9838,N_8961,N_6337);
and U9839 (N_9839,N_8219,N_8023);
nor U9840 (N_9840,N_7074,N_6232);
or U9841 (N_9841,N_7813,N_6172);
and U9842 (N_9842,N_8375,N_6733);
nand U9843 (N_9843,N_6601,N_7482);
and U9844 (N_9844,N_6814,N_7399);
nand U9845 (N_9845,N_8697,N_7929);
and U9846 (N_9846,N_6775,N_8120);
or U9847 (N_9847,N_6641,N_8561);
nand U9848 (N_9848,N_7471,N_8374);
or U9849 (N_9849,N_8504,N_7684);
or U9850 (N_9850,N_7651,N_8424);
nor U9851 (N_9851,N_8732,N_8934);
nor U9852 (N_9852,N_7222,N_6417);
nand U9853 (N_9853,N_8766,N_6892);
nor U9854 (N_9854,N_8373,N_7478);
nand U9855 (N_9855,N_8687,N_8621);
xnor U9856 (N_9856,N_7971,N_8499);
or U9857 (N_9857,N_7995,N_8719);
or U9858 (N_9858,N_6122,N_8698);
nor U9859 (N_9859,N_7713,N_6715);
or U9860 (N_9860,N_8741,N_7979);
and U9861 (N_9861,N_7874,N_7165);
or U9862 (N_9862,N_6981,N_7951);
xor U9863 (N_9863,N_8873,N_8639);
or U9864 (N_9864,N_8446,N_6443);
and U9865 (N_9865,N_8514,N_7420);
or U9866 (N_9866,N_6613,N_8546);
nor U9867 (N_9867,N_8615,N_8731);
or U9868 (N_9868,N_6792,N_7090);
nor U9869 (N_9869,N_6769,N_6345);
or U9870 (N_9870,N_6502,N_7141);
or U9871 (N_9871,N_8129,N_7454);
or U9872 (N_9872,N_6422,N_7248);
or U9873 (N_9873,N_7191,N_8002);
and U9874 (N_9874,N_6661,N_7805);
and U9875 (N_9875,N_8522,N_6985);
nand U9876 (N_9876,N_8857,N_6642);
nand U9877 (N_9877,N_6975,N_6427);
nor U9878 (N_9878,N_6725,N_7563);
or U9879 (N_9879,N_8966,N_8798);
xnor U9880 (N_9880,N_8807,N_6238);
nand U9881 (N_9881,N_8787,N_6784);
and U9882 (N_9882,N_7009,N_8119);
nor U9883 (N_9883,N_8295,N_7761);
and U9884 (N_9884,N_8510,N_6250);
nor U9885 (N_9885,N_8962,N_8461);
nand U9886 (N_9886,N_6726,N_6907);
or U9887 (N_9887,N_6452,N_8940);
or U9888 (N_9888,N_8108,N_6186);
nand U9889 (N_9889,N_8281,N_8036);
nor U9890 (N_9890,N_8128,N_6408);
nor U9891 (N_9891,N_6325,N_8487);
nor U9892 (N_9892,N_6243,N_6750);
and U9893 (N_9893,N_8115,N_7039);
nor U9894 (N_9894,N_6959,N_7422);
nand U9895 (N_9895,N_6810,N_6182);
nand U9896 (N_9896,N_8453,N_7615);
nor U9897 (N_9897,N_7131,N_8232);
nand U9898 (N_9898,N_6940,N_6561);
nor U9899 (N_9899,N_8780,N_6321);
nor U9900 (N_9900,N_8167,N_6113);
and U9901 (N_9901,N_7741,N_6850);
nor U9902 (N_9902,N_8735,N_7578);
nand U9903 (N_9903,N_6096,N_6979);
and U9904 (N_9904,N_8742,N_6686);
or U9905 (N_9905,N_6808,N_6688);
nand U9906 (N_9906,N_8333,N_6549);
nor U9907 (N_9907,N_7190,N_7772);
nor U9908 (N_9908,N_6973,N_8975);
and U9909 (N_9909,N_8871,N_6094);
nor U9910 (N_9910,N_6716,N_8528);
nand U9911 (N_9911,N_8646,N_8781);
and U9912 (N_9912,N_6575,N_7368);
nand U9913 (N_9913,N_6949,N_7697);
nand U9914 (N_9914,N_8603,N_7698);
nor U9915 (N_9915,N_7031,N_6777);
or U9916 (N_9916,N_8485,N_7484);
and U9917 (N_9917,N_6100,N_6118);
nor U9918 (N_9918,N_6466,N_8753);
and U9919 (N_9919,N_6917,N_8447);
and U9920 (N_9920,N_8459,N_7361);
nand U9921 (N_9921,N_7393,N_7487);
nand U9922 (N_9922,N_8574,N_8554);
or U9923 (N_9923,N_7945,N_7208);
nor U9924 (N_9924,N_6972,N_8709);
nand U9925 (N_9925,N_6693,N_7470);
or U9926 (N_9926,N_6753,N_7178);
nand U9927 (N_9927,N_7253,N_7991);
nand U9928 (N_9928,N_8344,N_7320);
nor U9929 (N_9929,N_7605,N_6195);
or U9930 (N_9930,N_8060,N_7379);
nor U9931 (N_9931,N_7833,N_7966);
and U9932 (N_9932,N_7083,N_8812);
nand U9933 (N_9933,N_8933,N_8125);
nand U9934 (N_9934,N_6474,N_6729);
and U9935 (N_9935,N_8973,N_6453);
nand U9936 (N_9936,N_7690,N_6976);
and U9937 (N_9937,N_8026,N_7819);
nor U9938 (N_9938,N_8841,N_8498);
nand U9939 (N_9939,N_7469,N_7430);
nand U9940 (N_9940,N_8368,N_7837);
nor U9941 (N_9941,N_8573,N_8411);
nor U9942 (N_9942,N_6692,N_7794);
and U9943 (N_9943,N_6507,N_6056);
nand U9944 (N_9944,N_7100,N_8601);
nand U9945 (N_9945,N_6800,N_8969);
or U9946 (N_9946,N_8405,N_8464);
and U9947 (N_9947,N_6546,N_7892);
and U9948 (N_9948,N_8736,N_6839);
and U9949 (N_9949,N_8773,N_8070);
or U9950 (N_9950,N_8511,N_8274);
or U9951 (N_9951,N_7538,N_7648);
or U9952 (N_9952,N_8984,N_6187);
nand U9953 (N_9953,N_8442,N_8988);
xnor U9954 (N_9954,N_6825,N_7499);
nand U9955 (N_9955,N_8301,N_7088);
or U9956 (N_9956,N_7668,N_7626);
or U9957 (N_9957,N_8800,N_6415);
nor U9958 (N_9958,N_8518,N_6665);
and U9959 (N_9959,N_8286,N_7843);
nor U9960 (N_9960,N_7352,N_8524);
and U9961 (N_9961,N_8243,N_7731);
or U9962 (N_9962,N_6288,N_7984);
or U9963 (N_9963,N_6016,N_6707);
or U9964 (N_9964,N_8085,N_7488);
and U9965 (N_9965,N_7116,N_8925);
and U9966 (N_9966,N_8963,N_8491);
or U9967 (N_9967,N_7452,N_7250);
nor U9968 (N_9968,N_7260,N_8979);
nand U9969 (N_9969,N_7214,N_6434);
or U9970 (N_9970,N_7785,N_7035);
or U9971 (N_9971,N_6834,N_7093);
or U9972 (N_9972,N_6580,N_6754);
or U9973 (N_9973,N_8196,N_6717);
and U9974 (N_9974,N_8174,N_6024);
nor U9975 (N_9975,N_8648,N_7683);
and U9976 (N_9976,N_6449,N_6497);
or U9977 (N_9977,N_7724,N_6780);
or U9978 (N_9978,N_7671,N_7301);
nor U9979 (N_9979,N_7175,N_6258);
and U9980 (N_9980,N_7925,N_7774);
or U9981 (N_9981,N_6986,N_6490);
nand U9982 (N_9982,N_7595,N_7225);
or U9983 (N_9983,N_6730,N_6578);
and U9984 (N_9984,N_7117,N_8953);
nor U9985 (N_9985,N_6437,N_7908);
and U9986 (N_9986,N_6660,N_8567);
or U9987 (N_9987,N_8182,N_7185);
nor U9988 (N_9988,N_7543,N_6015);
and U9989 (N_9989,N_6945,N_6393);
nor U9990 (N_9990,N_7992,N_6782);
or U9991 (N_9991,N_8558,N_7209);
or U9992 (N_9992,N_6389,N_6235);
nand U9993 (N_9993,N_6491,N_7242);
nor U9994 (N_9994,N_6720,N_8692);
or U9995 (N_9995,N_7019,N_8854);
or U9996 (N_9996,N_8355,N_8501);
nor U9997 (N_9997,N_6822,N_8221);
and U9998 (N_9998,N_8837,N_7415);
and U9999 (N_9999,N_8302,N_6745);
nand U10000 (N_10000,N_8443,N_7652);
or U10001 (N_10001,N_7295,N_8483);
or U10002 (N_10002,N_6157,N_7804);
nor U10003 (N_10003,N_6588,N_6341);
or U10004 (N_10004,N_8991,N_6348);
and U10005 (N_10005,N_7756,N_6897);
nor U10006 (N_10006,N_6477,N_8530);
and U10007 (N_10007,N_8892,N_6698);
nor U10008 (N_10008,N_8303,N_6691);
nand U10009 (N_10009,N_7894,N_7307);
nor U10010 (N_10010,N_7050,N_6081);
nand U10011 (N_10011,N_7733,N_6216);
nand U10012 (N_10012,N_7630,N_8140);
nand U10013 (N_10013,N_6475,N_8983);
or U10014 (N_10014,N_6795,N_6570);
nand U10015 (N_10015,N_6419,N_8708);
nand U10016 (N_10016,N_7046,N_8744);
and U10017 (N_10017,N_7662,N_7857);
and U10018 (N_10018,N_6538,N_8642);
nor U10019 (N_10019,N_8335,N_8057);
nand U10020 (N_10020,N_7464,N_6519);
nand U10021 (N_10021,N_7075,N_8788);
or U10022 (N_10022,N_8209,N_8752);
and U10023 (N_10023,N_7091,N_8193);
nor U10024 (N_10024,N_6411,N_6942);
and U10025 (N_10025,N_7842,N_8180);
nand U10026 (N_10026,N_8712,N_6309);
nand U10027 (N_10027,N_6137,N_7299);
or U10028 (N_10028,N_6879,N_6723);
and U10029 (N_10029,N_8808,N_7624);
and U10030 (N_10030,N_6076,N_7026);
or U10031 (N_10031,N_6205,N_6793);
nand U10032 (N_10032,N_7112,N_8557);
or U10033 (N_10033,N_7274,N_7666);
and U10034 (N_10034,N_8952,N_8784);
or U10035 (N_10035,N_8323,N_7853);
or U10036 (N_10036,N_6988,N_8637);
nor U10037 (N_10037,N_6663,N_7201);
and U10038 (N_10038,N_6431,N_8415);
nor U10039 (N_10039,N_6630,N_8205);
or U10040 (N_10040,N_6370,N_6823);
nand U10041 (N_10041,N_6102,N_6786);
nand U10042 (N_10042,N_7773,N_8038);
nor U10043 (N_10043,N_6739,N_7975);
or U10044 (N_10044,N_6441,N_7238);
nor U10045 (N_10045,N_6078,N_6317);
nand U10046 (N_10046,N_7550,N_7643);
nand U10047 (N_10047,N_8816,N_6223);
or U10048 (N_10048,N_7354,N_8259);
and U10049 (N_10049,N_7255,N_6108);
nand U10050 (N_10050,N_7621,N_6817);
or U10051 (N_10051,N_6239,N_8484);
or U10052 (N_10052,N_8850,N_6140);
or U10053 (N_10053,N_6604,N_8613);
and U10054 (N_10054,N_8213,N_6999);
nand U10055 (N_10055,N_6450,N_7669);
or U10056 (N_10056,N_8360,N_7072);
or U10057 (N_10057,N_7329,N_8467);
xnor U10058 (N_10058,N_7557,N_8249);
and U10059 (N_10059,N_8577,N_6710);
nor U10060 (N_10060,N_6496,N_7374);
nor U10061 (N_10061,N_6599,N_6234);
nor U10062 (N_10062,N_6742,N_6464);
nand U10063 (N_10063,N_7189,N_8846);
and U10064 (N_10064,N_8782,N_8747);
nor U10065 (N_10065,N_7128,N_6675);
nand U10066 (N_10066,N_7584,N_7702);
nor U10067 (N_10067,N_8541,N_7923);
and U10068 (N_10068,N_7324,N_8929);
or U10069 (N_10069,N_7642,N_7369);
nand U10070 (N_10070,N_8016,N_8202);
nand U10071 (N_10071,N_6881,N_8191);
and U10072 (N_10072,N_8575,N_6064);
and U10073 (N_10073,N_6048,N_7511);
nor U10074 (N_10074,N_6820,N_8932);
nor U10075 (N_10075,N_8371,N_7127);
or U10076 (N_10076,N_7102,N_7034);
nor U10077 (N_10077,N_7455,N_7143);
or U10078 (N_10078,N_8608,N_7742);
nand U10079 (N_10079,N_6669,N_6356);
nand U10080 (N_10080,N_6148,N_6318);
nor U10081 (N_10081,N_6837,N_6586);
and U10082 (N_10082,N_7129,N_8505);
nor U10083 (N_10083,N_6298,N_6735);
nor U10084 (N_10084,N_8230,N_8458);
or U10085 (N_10085,N_6065,N_7681);
or U10086 (N_10086,N_8413,N_6853);
nand U10087 (N_10087,N_8595,N_7199);
nand U10088 (N_10088,N_6033,N_8320);
or U10089 (N_10089,N_6363,N_6831);
or U10090 (N_10090,N_7598,N_8580);
nor U10091 (N_10091,N_6392,N_6622);
nor U10092 (N_10092,N_6069,N_8655);
nor U10093 (N_10093,N_8027,N_8378);
and U10094 (N_10094,N_7236,N_6162);
and U10095 (N_10095,N_8500,N_6270);
or U10096 (N_10096,N_7863,N_7766);
or U10097 (N_10097,N_6346,N_7911);
nor U10098 (N_10098,N_8851,N_7647);
and U10099 (N_10099,N_8241,N_6470);
nor U10100 (N_10100,N_8556,N_6978);
nand U10101 (N_10101,N_6029,N_7840);
or U10102 (N_10102,N_8181,N_6221);
and U10103 (N_10103,N_8513,N_6130);
nand U10104 (N_10104,N_7510,N_8755);
nand U10105 (N_10105,N_7241,N_8293);
nor U10106 (N_10106,N_6329,N_8578);
nor U10107 (N_10107,N_7725,N_8328);
nor U10108 (N_10108,N_6676,N_7950);
and U10109 (N_10109,N_8348,N_8472);
nand U10110 (N_10110,N_6451,N_8392);
nor U10111 (N_10111,N_7816,N_8224);
nor U10112 (N_10112,N_7279,N_8936);
nor U10113 (N_10113,N_6564,N_7645);
and U10114 (N_10114,N_6299,N_7402);
nor U10115 (N_10115,N_7859,N_8852);
nand U10116 (N_10116,N_8726,N_8350);
and U10117 (N_10117,N_6089,N_8768);
or U10118 (N_10118,N_6888,N_6099);
nand U10119 (N_10119,N_6269,N_7694);
and U10120 (N_10120,N_6138,N_7261);
or U10121 (N_10121,N_6054,N_8401);
or U10122 (N_10122,N_8144,N_7986);
or U10123 (N_10123,N_6980,N_7011);
and U10124 (N_10124,N_8422,N_8417);
nor U10125 (N_10125,N_8928,N_6047);
or U10126 (N_10126,N_6030,N_7928);
nand U10127 (N_10127,N_7705,N_8585);
nand U10128 (N_10128,N_8194,N_7632);
and U10129 (N_10129,N_8538,N_8050);
nand U10130 (N_10130,N_7781,N_8433);
or U10131 (N_10131,N_6783,N_6175);
nor U10132 (N_10132,N_6362,N_8322);
and U10133 (N_10133,N_6855,N_7940);
or U10134 (N_10134,N_8549,N_8225);
or U10135 (N_10135,N_7142,N_6440);
and U10136 (N_10136,N_7481,N_7963);
nand U10137 (N_10137,N_6149,N_7521);
nor U10138 (N_10138,N_8978,N_7809);
nand U10139 (N_10139,N_6929,N_7252);
nand U10140 (N_10140,N_7982,N_8763);
nand U10141 (N_10141,N_7292,N_7939);
and U10142 (N_10142,N_6101,N_7780);
xor U10143 (N_10143,N_6799,N_7798);
nor U10144 (N_10144,N_7346,N_8000);
nor U10145 (N_10145,N_8386,N_8242);
nor U10146 (N_10146,N_6418,N_8064);
and U10147 (N_10147,N_7865,N_8018);
nor U10148 (N_10148,N_8310,N_6414);
and U10149 (N_10149,N_7808,N_6982);
nand U10150 (N_10150,N_7269,N_7177);
nand U10151 (N_10151,N_7501,N_7052);
nand U10152 (N_10152,N_7341,N_8351);
nand U10153 (N_10153,N_8540,N_8777);
or U10154 (N_10154,N_8200,N_8496);
nor U10155 (N_10155,N_8910,N_7257);
or U10156 (N_10156,N_6579,N_7587);
and U10157 (N_10157,N_6009,N_8880);
or U10158 (N_10158,N_6974,N_6501);
and U10159 (N_10159,N_8711,N_7875);
nor U10160 (N_10160,N_8959,N_8559);
nand U10161 (N_10161,N_7882,N_7096);
and U10162 (N_10162,N_7967,N_6202);
or U10163 (N_10163,N_6938,N_8682);
and U10164 (N_10164,N_6748,N_7044);
or U10165 (N_10165,N_6734,N_7433);
or U10166 (N_10166,N_7540,N_6694);
and U10167 (N_10167,N_7564,N_8031);
and U10168 (N_10168,N_6617,N_6607);
nor U10169 (N_10169,N_7597,N_6860);
or U10170 (N_10170,N_7876,N_8233);
nand U10171 (N_10171,N_8071,N_7391);
or U10172 (N_10172,N_6555,N_7317);
or U10173 (N_10173,N_6262,N_6136);
nor U10174 (N_10174,N_6057,N_7162);
nor U10175 (N_10175,N_8919,N_6516);
and U10176 (N_10176,N_6738,N_7706);
or U10177 (N_10177,N_8771,N_8614);
nand U10178 (N_10178,N_8315,N_7210);
and U10179 (N_10179,N_6602,N_6369);
nand U10180 (N_10180,N_7337,N_8737);
nand U10181 (N_10181,N_7223,N_8250);
xnor U10182 (N_10182,N_7022,N_7263);
nand U10183 (N_10183,N_6457,N_8463);
and U10184 (N_10184,N_7319,N_8212);
nand U10185 (N_10185,N_8654,N_7002);
nor U10186 (N_10186,N_8917,N_7949);
or U10187 (N_10187,N_7588,N_6874);
or U10188 (N_10188,N_6043,N_7113);
nand U10189 (N_10189,N_6543,N_8778);
or U10190 (N_10190,N_7460,N_8247);
or U10191 (N_10191,N_7372,N_8204);
nor U10192 (N_10192,N_6605,N_6273);
nand U10193 (N_10193,N_8065,N_7081);
or U10194 (N_10194,N_8074,N_7239);
and U10195 (N_10195,N_8434,N_8960);
or U10196 (N_10196,N_6286,N_7048);
nor U10197 (N_10197,N_6510,N_8911);
nor U10198 (N_10198,N_6567,N_8644);
nand U10199 (N_10199,N_7751,N_8343);
nor U10200 (N_10200,N_6225,N_6915);
and U10201 (N_10201,N_7150,N_6867);
or U10202 (N_10202,N_6447,N_6040);
or U10203 (N_10203,N_7159,N_6376);
and U10204 (N_10204,N_8098,N_6632);
and U10205 (N_10205,N_7414,N_6637);
nor U10206 (N_10206,N_8519,N_8695);
or U10207 (N_10207,N_7474,N_8795);
nand U10208 (N_10208,N_6668,N_7522);
nand U10209 (N_10209,N_7841,N_7140);
nand U10210 (N_10210,N_7767,N_7577);
nand U10211 (N_10211,N_6503,N_6183);
or U10212 (N_10212,N_8029,N_6806);
and U10213 (N_10213,N_6532,N_8803);
nand U10214 (N_10214,N_8056,N_6433);
and U10215 (N_10215,N_6178,N_7174);
nor U10216 (N_10216,N_7204,N_7912);
nand U10217 (N_10217,N_6297,N_7854);
or U10218 (N_10218,N_7802,N_7549);
nand U10219 (N_10219,N_7519,N_7154);
nand U10220 (N_10220,N_6788,N_8998);
and U10221 (N_10221,N_7272,N_6218);
nor U10222 (N_10222,N_8651,N_7355);
or U10223 (N_10223,N_7373,N_8288);
nand U10224 (N_10224,N_6712,N_7818);
and U10225 (N_10225,N_8550,N_7688);
or U10226 (N_10226,N_6721,N_6643);
or U10227 (N_10227,N_8964,N_8834);
and U10228 (N_10228,N_6673,N_7893);
or U10229 (N_10229,N_7340,N_6296);
and U10230 (N_10230,N_8408,N_7749);
and U10231 (N_10231,N_7138,N_8260);
and U10232 (N_10232,N_6582,N_8438);
and U10233 (N_10233,N_6955,N_6125);
nor U10234 (N_10234,N_6272,N_7782);
and U10235 (N_10235,N_8589,N_8703);
nand U10236 (N_10236,N_7397,N_8092);
nand U10237 (N_10237,N_7507,N_7407);
and U10238 (N_10238,N_7366,N_6851);
nor U10239 (N_10239,N_8565,N_6947);
nor U10240 (N_10240,N_8214,N_6072);
nor U10241 (N_10241,N_7264,N_6568);
nor U10242 (N_10242,N_6014,N_6242);
or U10243 (N_10243,N_7738,N_6600);
nor U10244 (N_10244,N_7110,N_6372);
xnor U10245 (N_10245,N_6912,N_8145);
or U10246 (N_10246,N_6007,N_6962);
nand U10247 (N_10247,N_6821,N_7432);
and U10248 (N_10248,N_8326,N_6319);
or U10249 (N_10249,N_7145,N_7855);
and U10250 (N_10250,N_8126,N_7883);
nor U10251 (N_10251,N_6536,N_8727);
and U10252 (N_10252,N_8858,N_7858);
nand U10253 (N_10253,N_7699,N_8105);
nand U10254 (N_10254,N_7010,N_6107);
xor U10255 (N_10255,N_8716,N_8283);
nand U10256 (N_10256,N_7275,N_6552);
nand U10257 (N_10257,N_7381,N_6438);
and U10258 (N_10258,N_8761,N_6989);
and U10259 (N_10259,N_8273,N_6388);
or U10260 (N_10260,N_8745,N_7383);
and U10261 (N_10261,N_6708,N_8706);
and U10262 (N_10262,N_8077,N_8882);
nand U10263 (N_10263,N_8184,N_6254);
and U10264 (N_10264,N_8020,N_7607);
nor U10265 (N_10265,N_6873,N_7013);
and U10266 (N_10266,N_7672,N_8084);
and U10267 (N_10267,N_8775,N_8599);
nor U10268 (N_10268,N_8047,N_6534);
and U10269 (N_10269,N_7001,N_7202);
nand U10270 (N_10270,N_8149,N_8636);
nand U10271 (N_10271,N_7343,N_7852);
and U10272 (N_10272,N_7512,N_8779);
nand U10273 (N_10273,N_6189,N_8985);
or U10274 (N_10274,N_8095,N_8428);
nand U10275 (N_10275,N_8365,N_6022);
and U10276 (N_10276,N_6240,N_7957);
nand U10277 (N_10277,N_7055,N_8903);
nand U10278 (N_10278,N_8083,N_8460);
nand U10279 (N_10279,N_6843,N_7523);
and U10280 (N_10280,N_7895,N_8754);
and U10281 (N_10281,N_8990,N_8104);
nor U10282 (N_10282,N_6248,N_7087);
or U10283 (N_10283,N_8134,N_7321);
and U10284 (N_10284,N_6760,N_8037);
and U10285 (N_10285,N_7479,N_8137);
nand U10286 (N_10286,N_7983,N_8531);
nor U10287 (N_10287,N_7084,N_6773);
or U10288 (N_10288,N_6935,N_8117);
or U10289 (N_10289,N_8715,N_7604);
nor U10290 (N_10290,N_8127,N_6796);
or U10291 (N_10291,N_6998,N_6918);
nand U10292 (N_10292,N_8859,N_8096);
nor U10293 (N_10293,N_8478,N_6409);
and U10294 (N_10294,N_7491,N_6049);
nand U10295 (N_10295,N_7670,N_6407);
and U10296 (N_10296,N_6037,N_7736);
and U10297 (N_10297,N_7826,N_7998);
xnor U10298 (N_10298,N_6017,N_8090);
and U10299 (N_10299,N_8931,N_7517);
or U10300 (N_10300,N_6848,N_6055);
and U10301 (N_10301,N_6528,N_8506);
nand U10302 (N_10302,N_7727,N_8520);
nor U10303 (N_10303,N_7922,N_8005);
nand U10304 (N_10304,N_6529,N_7931);
nand U10305 (N_10305,N_7447,N_7157);
nor U10306 (N_10306,N_8883,N_7152);
nand U10307 (N_10307,N_7812,N_7509);
nor U10308 (N_10308,N_6087,N_7349);
and U10309 (N_10309,N_6364,N_6323);
nor U10310 (N_10310,N_6514,N_8676);
nand U10311 (N_10311,N_6109,N_7667);
nand U10312 (N_10312,N_8116,N_6126);
nand U10313 (N_10313,N_7784,N_6264);
nand U10314 (N_10314,N_6472,N_8802);
and U10315 (N_10315,N_6901,N_8865);
and U10316 (N_10316,N_6428,N_6684);
nand U10317 (N_10317,N_6103,N_6756);
and U10318 (N_10318,N_8818,N_6573);
nand U10319 (N_10319,N_8410,N_7601);
and U10320 (N_10320,N_7591,N_6550);
nor U10321 (N_10321,N_8597,N_7288);
or U10322 (N_10322,N_8142,N_7915);
nand U10323 (N_10323,N_8584,N_7703);
and U10324 (N_10324,N_7326,N_8151);
and U10325 (N_10325,N_6809,N_8118);
and U10326 (N_10326,N_7082,N_6646);
and U10327 (N_10327,N_6763,N_8872);
or U10328 (N_10328,N_7754,N_7964);
nand U10329 (N_10329,N_7086,N_7440);
nor U10330 (N_10330,N_8722,N_8369);
and U10331 (N_10331,N_8477,N_7375);
nor U10332 (N_10332,N_8041,N_8279);
or U10333 (N_10333,N_7418,N_7514);
nand U10334 (N_10334,N_7625,N_8734);
and U10335 (N_10335,N_7663,N_7476);
and U10336 (N_10336,N_6882,N_6743);
nor U10337 (N_10337,N_6544,N_8509);
nand U10338 (N_10338,N_6925,N_6331);
or U10339 (N_10339,N_8276,N_6899);
and U10340 (N_10340,N_6042,N_8699);
nor U10341 (N_10341,N_7902,N_6964);
nand U10342 (N_10342,N_7515,N_7276);
and U10343 (N_10343,N_8271,N_7799);
nand U10344 (N_10344,N_7149,N_6909);
nor U10345 (N_10345,N_6977,N_6522);
or U10346 (N_10346,N_7156,N_7948);
nor U10347 (N_10347,N_8893,N_6526);
nor U10348 (N_10348,N_7330,N_7535);
or U10349 (N_10349,N_6606,N_6870);
or U10350 (N_10350,N_6141,N_8995);
or U10351 (N_10351,N_6762,N_7300);
and U10352 (N_10352,N_8345,N_7426);
nor U10353 (N_10353,N_6589,N_7661);
or U10354 (N_10354,N_8339,N_6073);
or U10355 (N_10355,N_8746,N_8717);
nand U10356 (N_10356,N_6343,N_6359);
or U10357 (N_10357,N_8688,N_7453);
nor U10358 (N_10358,N_7752,N_6215);
and U10359 (N_10359,N_6565,N_8399);
nand U10360 (N_10360,N_6488,N_8390);
nor U10361 (N_10361,N_6093,N_8341);
and U10362 (N_10362,N_6006,N_6421);
and U10363 (N_10363,N_7437,N_6120);
nand U10364 (N_10364,N_7327,N_8822);
or U10365 (N_10365,N_8262,N_6026);
nor U10366 (N_10366,N_8009,N_6211);
and U10367 (N_10367,N_8261,N_7061);
and U10368 (N_10368,N_8827,N_6170);
nor U10369 (N_10369,N_7695,N_6217);
and U10370 (N_10370,N_8826,N_8489);
nor U10371 (N_10371,N_8582,N_6883);
and U10372 (N_10372,N_6506,N_7555);
and U10373 (N_10373,N_6807,N_7955);
or U10374 (N_10374,N_6251,N_6877);
and U10375 (N_10375,N_7677,N_7389);
nand U10376 (N_10376,N_8946,N_6303);
nand U10377 (N_10377,N_8296,N_8832);
nand U10378 (N_10378,N_6811,N_6302);
nand U10379 (N_10379,N_6841,N_8299);
or U10380 (N_10380,N_6192,N_8435);
nor U10381 (N_10381,N_8909,N_6776);
or U10382 (N_10382,N_6063,N_6476);
nand U10383 (N_10383,N_6027,N_7885);
or U10384 (N_10384,N_7158,N_6011);
or U10385 (N_10385,N_8420,N_7064);
and U10386 (N_10386,N_7280,N_7421);
and U10387 (N_10387,N_8078,N_6067);
or U10388 (N_10388,N_7834,N_7527);
or U10389 (N_10389,N_7436,N_8377);
or U10390 (N_10390,N_6097,N_7104);
nand U10391 (N_10391,N_8171,N_7249);
nor U10392 (N_10392,N_6757,N_7188);
nand U10393 (N_10393,N_8441,N_6295);
or U10394 (N_10394,N_6801,N_6828);
or U10395 (N_10395,N_8376,N_6013);
nand U10396 (N_10396,N_6313,N_8432);
nand U10397 (N_10397,N_8539,N_7126);
nor U10398 (N_10398,N_8548,N_7148);
and U10399 (N_10399,N_7020,N_6201);
nand U10400 (N_10400,N_7115,N_8634);
nor U10401 (N_10401,N_6581,N_6731);
and U10402 (N_10402,N_6804,N_6259);
nand U10403 (N_10403,N_7927,N_8352);
and U10404 (N_10404,N_6358,N_6827);
nand U10405 (N_10405,N_6505,N_8774);
and U10406 (N_10406,N_8670,N_6967);
and U10407 (N_10407,N_7444,N_8671);
nand U10408 (N_10408,N_8996,N_6276);
or U10409 (N_10409,N_6191,N_7900);
nor U10410 (N_10410,N_8840,N_7530);
nor U10411 (N_10411,N_6342,N_7721);
and U10412 (N_10412,N_7018,N_8272);
or U10413 (N_10413,N_7811,N_6277);
nor U10414 (N_10414,N_6380,N_6540);
or U10415 (N_10415,N_7629,N_7868);
nor U10416 (N_10416,N_7041,N_6937);
nor U10417 (N_10417,N_7486,N_6996);
and U10418 (N_10418,N_6608,N_8179);
and U10419 (N_10419,N_8664,N_7646);
or U10420 (N_10420,N_7734,N_7097);
nand U10421 (N_10421,N_8986,N_8896);
nor U10422 (N_10422,N_7500,N_8863);
or U10423 (N_10423,N_6104,N_6077);
xor U10424 (N_10424,N_7793,N_8357);
nand U10425 (N_10425,N_7567,N_8102);
nor U10426 (N_10426,N_7609,N_8395);
and U10427 (N_10427,N_8468,N_7796);
nor U10428 (N_10428,N_8277,N_7226);
nor U10429 (N_10429,N_8073,N_8185);
nor U10430 (N_10430,N_7999,N_7712);
nor U10431 (N_10431,N_7562,N_7678);
or U10432 (N_10432,N_8495,N_6314);
or U10433 (N_10433,N_6494,N_7182);
and U10434 (N_10434,N_6274,N_8926);
nand U10435 (N_10435,N_7861,N_8629);
nor U10436 (N_10436,N_7576,N_7817);
and U10437 (N_10437,N_6732,N_7777);
or U10438 (N_10438,N_7417,N_8829);
nand U10439 (N_10439,N_8007,N_8017);
or U10440 (N_10440,N_8720,N_8867);
or U10441 (N_10441,N_8336,N_6044);
nor U10442 (N_10442,N_8879,N_8427);
and U10443 (N_10443,N_7386,N_6051);
nand U10444 (N_10444,N_8058,N_6291);
nor U10445 (N_10445,N_7144,N_8897);
nor U10446 (N_10446,N_6655,N_8265);
nand U10447 (N_10447,N_7122,N_8021);
or U10448 (N_10448,N_6283,N_7574);
or U10449 (N_10449,N_8327,N_7006);
nor U10450 (N_10450,N_7759,N_8821);
and U10451 (N_10451,N_7395,N_6960);
nand U10452 (N_10452,N_8033,N_7884);
nand U10453 (N_10453,N_6424,N_8226);
nand U10454 (N_10454,N_7898,N_6284);
nand U10455 (N_10455,N_7828,N_6090);
nor U10456 (N_10456,N_7716,N_6111);
or U10457 (N_10457,N_8977,N_8662);
and U10458 (N_10458,N_6616,N_8783);
or U10459 (N_10459,N_6521,N_7351);
nor U10460 (N_10460,N_7881,N_6593);
and U10461 (N_10461,N_7762,N_8176);
nor U10462 (N_10462,N_6495,N_8228);
or U10463 (N_10463,N_6787,N_8679);
or U10464 (N_10464,N_7679,N_7990);
nand U10465 (N_10465,N_7405,N_7298);
nor U10466 (N_10466,N_8770,N_7689);
or U10467 (N_10467,N_7377,N_8740);
and U10468 (N_10468,N_7285,N_8431);
and U10469 (N_10469,N_8394,N_7619);
and U10470 (N_10470,N_8493,N_8406);
nand U10471 (N_10471,N_6498,N_7008);
nor U10472 (N_10472,N_6025,N_8081);
nor U10473 (N_10473,N_6670,N_8912);
nand U10474 (N_10474,N_7028,N_8207);
nor U10475 (N_10475,N_6504,N_6395);
nor U10476 (N_10476,N_7049,N_6648);
or U10477 (N_10477,N_8923,N_6657);
nand U10478 (N_10478,N_6231,N_7620);
nand U10479 (N_10479,N_7147,N_7217);
or U10480 (N_10480,N_7635,N_7465);
nor U10481 (N_10481,N_8823,N_8049);
nor U10482 (N_10482,N_6563,N_8656);
nand U10483 (N_10483,N_7227,N_6010);
and U10484 (N_10484,N_6377,N_8534);
nor U10485 (N_10485,N_8475,N_7021);
or U10486 (N_10486,N_8159,N_8949);
nand U10487 (N_10487,N_8680,N_7580);
xor U10488 (N_10488,N_7078,N_7380);
and U10489 (N_10489,N_7542,N_6263);
nand U10490 (N_10490,N_6184,N_8359);
and U10491 (N_10491,N_8263,N_7961);
and U10492 (N_10492,N_6280,N_7004);
or U10493 (N_10493,N_8819,N_7137);
nand U10494 (N_10494,N_8701,N_6032);
or U10495 (N_10495,N_6485,N_8881);
and U10496 (N_10496,N_8756,N_8627);
nor U10497 (N_10497,N_6512,N_6460);
nand U10498 (N_10498,N_6993,N_6257);
nand U10499 (N_10499,N_7825,N_8270);
nand U10500 (N_10500,N_8916,N_8322);
or U10501 (N_10501,N_8898,N_7761);
nor U10502 (N_10502,N_7374,N_8087);
nor U10503 (N_10503,N_6110,N_7106);
and U10504 (N_10504,N_8925,N_7254);
nor U10505 (N_10505,N_8478,N_8158);
and U10506 (N_10506,N_6688,N_7296);
nor U10507 (N_10507,N_7986,N_6284);
and U10508 (N_10508,N_8652,N_8791);
and U10509 (N_10509,N_8436,N_6349);
xor U10510 (N_10510,N_7530,N_6040);
or U10511 (N_10511,N_6910,N_7755);
nand U10512 (N_10512,N_7993,N_6133);
nand U10513 (N_10513,N_7303,N_6136);
and U10514 (N_10514,N_8137,N_6148);
or U10515 (N_10515,N_6207,N_6309);
or U10516 (N_10516,N_7364,N_6397);
nor U10517 (N_10517,N_6330,N_8027);
nor U10518 (N_10518,N_6365,N_7710);
nor U10519 (N_10519,N_6515,N_6759);
or U10520 (N_10520,N_8872,N_6474);
nor U10521 (N_10521,N_8528,N_7335);
nand U10522 (N_10522,N_6237,N_8561);
nand U10523 (N_10523,N_7427,N_6390);
or U10524 (N_10524,N_6286,N_8079);
or U10525 (N_10525,N_7001,N_8162);
nand U10526 (N_10526,N_7859,N_7733);
nor U10527 (N_10527,N_7870,N_8245);
or U10528 (N_10528,N_6264,N_8272);
or U10529 (N_10529,N_6806,N_6529);
and U10530 (N_10530,N_8202,N_7772);
nand U10531 (N_10531,N_6123,N_7823);
nor U10532 (N_10532,N_8795,N_8040);
or U10533 (N_10533,N_7024,N_8181);
nor U10534 (N_10534,N_7283,N_8452);
nand U10535 (N_10535,N_8734,N_7827);
nand U10536 (N_10536,N_6528,N_6857);
and U10537 (N_10537,N_6241,N_6330);
nand U10538 (N_10538,N_8225,N_7995);
or U10539 (N_10539,N_8755,N_8501);
nor U10540 (N_10540,N_8926,N_7450);
and U10541 (N_10541,N_8689,N_8130);
nor U10542 (N_10542,N_6707,N_7566);
and U10543 (N_10543,N_6009,N_6582);
nand U10544 (N_10544,N_7161,N_7008);
or U10545 (N_10545,N_8275,N_7676);
nor U10546 (N_10546,N_6418,N_6778);
nand U10547 (N_10547,N_6522,N_7435);
or U10548 (N_10548,N_8235,N_8265);
nor U10549 (N_10549,N_8081,N_8764);
and U10550 (N_10550,N_7571,N_8852);
or U10551 (N_10551,N_7075,N_7878);
nand U10552 (N_10552,N_7802,N_8484);
nand U10553 (N_10553,N_8906,N_7002);
nand U10554 (N_10554,N_8936,N_6422);
nor U10555 (N_10555,N_7899,N_8954);
or U10556 (N_10556,N_7542,N_6385);
nand U10557 (N_10557,N_8885,N_7514);
or U10558 (N_10558,N_8947,N_6312);
and U10559 (N_10559,N_6416,N_8076);
nor U10560 (N_10560,N_8605,N_8467);
nor U10561 (N_10561,N_7310,N_8729);
nand U10562 (N_10562,N_8166,N_6659);
or U10563 (N_10563,N_7998,N_7350);
or U10564 (N_10564,N_6818,N_6152);
nand U10565 (N_10565,N_7330,N_8017);
and U10566 (N_10566,N_8678,N_6982);
or U10567 (N_10567,N_8689,N_7235);
and U10568 (N_10568,N_6028,N_7623);
nand U10569 (N_10569,N_6297,N_8946);
nor U10570 (N_10570,N_6913,N_7949);
or U10571 (N_10571,N_8637,N_8139);
or U10572 (N_10572,N_7639,N_6084);
or U10573 (N_10573,N_7918,N_7763);
nor U10574 (N_10574,N_8860,N_7612);
and U10575 (N_10575,N_8567,N_8602);
nand U10576 (N_10576,N_8761,N_8558);
nor U10577 (N_10577,N_8687,N_8227);
and U10578 (N_10578,N_6035,N_6130);
nand U10579 (N_10579,N_7372,N_6066);
or U10580 (N_10580,N_6468,N_7948);
or U10581 (N_10581,N_8508,N_8904);
or U10582 (N_10582,N_6541,N_8704);
nand U10583 (N_10583,N_8284,N_7961);
nand U10584 (N_10584,N_6875,N_6413);
nor U10585 (N_10585,N_7302,N_7091);
or U10586 (N_10586,N_6158,N_7092);
and U10587 (N_10587,N_8665,N_7247);
nand U10588 (N_10588,N_6059,N_6721);
or U10589 (N_10589,N_8947,N_7037);
nor U10590 (N_10590,N_7619,N_6948);
nand U10591 (N_10591,N_6471,N_8507);
or U10592 (N_10592,N_8091,N_6180);
and U10593 (N_10593,N_7815,N_8642);
or U10594 (N_10594,N_7914,N_8111);
and U10595 (N_10595,N_8058,N_6085);
or U10596 (N_10596,N_6186,N_7034);
and U10597 (N_10597,N_8931,N_8725);
nand U10598 (N_10598,N_8562,N_6778);
nor U10599 (N_10599,N_6828,N_8631);
nand U10600 (N_10600,N_7977,N_7169);
nor U10601 (N_10601,N_6687,N_6638);
nand U10602 (N_10602,N_6385,N_8895);
and U10603 (N_10603,N_6527,N_7182);
nand U10604 (N_10604,N_8079,N_7169);
and U10605 (N_10605,N_7219,N_6715);
or U10606 (N_10606,N_6871,N_8702);
or U10607 (N_10607,N_8793,N_8820);
nor U10608 (N_10608,N_8851,N_7354);
nor U10609 (N_10609,N_8090,N_8802);
and U10610 (N_10610,N_7761,N_6875);
nor U10611 (N_10611,N_7989,N_8208);
or U10612 (N_10612,N_7988,N_6435);
and U10613 (N_10613,N_8219,N_8256);
nand U10614 (N_10614,N_6313,N_7473);
nor U10615 (N_10615,N_6687,N_6256);
nand U10616 (N_10616,N_6533,N_7720);
or U10617 (N_10617,N_6474,N_8588);
and U10618 (N_10618,N_6988,N_8378);
nand U10619 (N_10619,N_7006,N_7893);
or U10620 (N_10620,N_7633,N_8408);
and U10621 (N_10621,N_6003,N_7631);
nand U10622 (N_10622,N_6458,N_6236);
nor U10623 (N_10623,N_7664,N_7086);
and U10624 (N_10624,N_7815,N_6137);
nand U10625 (N_10625,N_7967,N_8580);
nor U10626 (N_10626,N_7925,N_7551);
nand U10627 (N_10627,N_7097,N_7992);
and U10628 (N_10628,N_8734,N_8722);
and U10629 (N_10629,N_7117,N_6395);
or U10630 (N_10630,N_8825,N_7894);
or U10631 (N_10631,N_8456,N_6764);
nand U10632 (N_10632,N_6178,N_7874);
and U10633 (N_10633,N_8287,N_8738);
nand U10634 (N_10634,N_6859,N_7499);
nand U10635 (N_10635,N_7837,N_8836);
and U10636 (N_10636,N_6917,N_6489);
nor U10637 (N_10637,N_6213,N_6749);
nand U10638 (N_10638,N_8143,N_8292);
nor U10639 (N_10639,N_6535,N_7607);
nor U10640 (N_10640,N_7453,N_8157);
or U10641 (N_10641,N_7509,N_8456);
nand U10642 (N_10642,N_6952,N_8712);
and U10643 (N_10643,N_7815,N_8029);
and U10644 (N_10644,N_8062,N_7513);
and U10645 (N_10645,N_6332,N_6174);
and U10646 (N_10646,N_6663,N_6696);
nand U10647 (N_10647,N_8868,N_7240);
and U10648 (N_10648,N_6010,N_7848);
or U10649 (N_10649,N_8095,N_6453);
nor U10650 (N_10650,N_7344,N_6061);
nand U10651 (N_10651,N_6165,N_6784);
and U10652 (N_10652,N_6629,N_6146);
and U10653 (N_10653,N_8331,N_6975);
nand U10654 (N_10654,N_6410,N_7773);
and U10655 (N_10655,N_8537,N_7446);
nand U10656 (N_10656,N_6804,N_6255);
nor U10657 (N_10657,N_7719,N_6301);
nand U10658 (N_10658,N_7391,N_7982);
nor U10659 (N_10659,N_8575,N_7731);
and U10660 (N_10660,N_7610,N_7312);
and U10661 (N_10661,N_6516,N_6265);
and U10662 (N_10662,N_6790,N_7667);
or U10663 (N_10663,N_6771,N_7294);
and U10664 (N_10664,N_6939,N_6555);
nor U10665 (N_10665,N_8691,N_8979);
or U10666 (N_10666,N_7651,N_6271);
nand U10667 (N_10667,N_6698,N_6813);
nor U10668 (N_10668,N_6355,N_8239);
and U10669 (N_10669,N_6814,N_8327);
or U10670 (N_10670,N_8079,N_6581);
and U10671 (N_10671,N_8168,N_7258);
nand U10672 (N_10672,N_8290,N_8990);
or U10673 (N_10673,N_7940,N_8085);
nand U10674 (N_10674,N_6315,N_8043);
nor U10675 (N_10675,N_6424,N_8481);
nor U10676 (N_10676,N_7081,N_8942);
nand U10677 (N_10677,N_7368,N_7262);
nand U10678 (N_10678,N_8900,N_8849);
nor U10679 (N_10679,N_7601,N_8300);
nor U10680 (N_10680,N_8671,N_6346);
nor U10681 (N_10681,N_6894,N_7345);
or U10682 (N_10682,N_8216,N_6891);
xor U10683 (N_10683,N_7711,N_6652);
nand U10684 (N_10684,N_8202,N_8628);
nor U10685 (N_10685,N_8180,N_6150);
nand U10686 (N_10686,N_6667,N_7858);
nand U10687 (N_10687,N_7133,N_8024);
nor U10688 (N_10688,N_8617,N_6023);
nand U10689 (N_10689,N_6907,N_7292);
and U10690 (N_10690,N_6816,N_6630);
nand U10691 (N_10691,N_6005,N_8348);
nand U10692 (N_10692,N_7661,N_8322);
or U10693 (N_10693,N_6571,N_8098);
nand U10694 (N_10694,N_7872,N_7570);
nand U10695 (N_10695,N_8790,N_6627);
nand U10696 (N_10696,N_6286,N_8403);
nor U10697 (N_10697,N_7419,N_8164);
or U10698 (N_10698,N_8259,N_6216);
or U10699 (N_10699,N_7701,N_6141);
or U10700 (N_10700,N_6509,N_6943);
or U10701 (N_10701,N_6502,N_7445);
and U10702 (N_10702,N_8395,N_6637);
nand U10703 (N_10703,N_8264,N_8183);
nand U10704 (N_10704,N_7856,N_6761);
and U10705 (N_10705,N_6711,N_6780);
or U10706 (N_10706,N_6378,N_8848);
and U10707 (N_10707,N_6152,N_8371);
or U10708 (N_10708,N_8220,N_7466);
and U10709 (N_10709,N_6865,N_6141);
nor U10710 (N_10710,N_6229,N_7763);
nor U10711 (N_10711,N_7464,N_6658);
and U10712 (N_10712,N_6277,N_6003);
or U10713 (N_10713,N_7231,N_8429);
nor U10714 (N_10714,N_6904,N_8704);
nor U10715 (N_10715,N_6714,N_7248);
or U10716 (N_10716,N_6211,N_6189);
and U10717 (N_10717,N_6109,N_7358);
or U10718 (N_10718,N_8476,N_8787);
nand U10719 (N_10719,N_7563,N_6188);
nor U10720 (N_10720,N_8942,N_7439);
and U10721 (N_10721,N_6575,N_6615);
and U10722 (N_10722,N_6324,N_8377);
and U10723 (N_10723,N_7482,N_7796);
or U10724 (N_10724,N_7777,N_8671);
nor U10725 (N_10725,N_8701,N_8791);
nor U10726 (N_10726,N_6712,N_8329);
nand U10727 (N_10727,N_6047,N_7260);
or U10728 (N_10728,N_6569,N_8328);
and U10729 (N_10729,N_7055,N_6787);
and U10730 (N_10730,N_8638,N_7872);
or U10731 (N_10731,N_6804,N_7513);
or U10732 (N_10732,N_6160,N_6664);
nand U10733 (N_10733,N_8586,N_7121);
nand U10734 (N_10734,N_6232,N_7971);
xor U10735 (N_10735,N_7253,N_6560);
or U10736 (N_10736,N_8739,N_8388);
nand U10737 (N_10737,N_8834,N_8587);
nor U10738 (N_10738,N_7047,N_8321);
nand U10739 (N_10739,N_6268,N_8797);
or U10740 (N_10740,N_8818,N_8219);
nor U10741 (N_10741,N_8249,N_8682);
or U10742 (N_10742,N_7516,N_6950);
and U10743 (N_10743,N_7164,N_6046);
or U10744 (N_10744,N_6581,N_7201);
or U10745 (N_10745,N_6516,N_6703);
or U10746 (N_10746,N_8465,N_7721);
nand U10747 (N_10747,N_7714,N_6218);
or U10748 (N_10748,N_8572,N_8493);
nor U10749 (N_10749,N_6571,N_6209);
or U10750 (N_10750,N_6449,N_7792);
nor U10751 (N_10751,N_8763,N_8520);
nor U10752 (N_10752,N_8083,N_7819);
or U10753 (N_10753,N_6555,N_7735);
or U10754 (N_10754,N_7565,N_8295);
or U10755 (N_10755,N_8316,N_7981);
nand U10756 (N_10756,N_8284,N_6605);
and U10757 (N_10757,N_8428,N_7694);
nand U10758 (N_10758,N_6265,N_6434);
nor U10759 (N_10759,N_6747,N_7424);
and U10760 (N_10760,N_6426,N_7114);
or U10761 (N_10761,N_6405,N_8658);
nand U10762 (N_10762,N_6048,N_6287);
or U10763 (N_10763,N_6801,N_7369);
nor U10764 (N_10764,N_7854,N_8318);
nor U10765 (N_10765,N_6868,N_7850);
or U10766 (N_10766,N_6613,N_8292);
nand U10767 (N_10767,N_6807,N_8448);
nor U10768 (N_10768,N_7529,N_7816);
or U10769 (N_10769,N_7655,N_8115);
nand U10770 (N_10770,N_6909,N_8892);
or U10771 (N_10771,N_6981,N_8152);
nand U10772 (N_10772,N_6748,N_7632);
nand U10773 (N_10773,N_7006,N_7823);
nand U10774 (N_10774,N_8428,N_7101);
or U10775 (N_10775,N_8360,N_6306);
or U10776 (N_10776,N_6014,N_6429);
nand U10777 (N_10777,N_7074,N_6831);
and U10778 (N_10778,N_8673,N_8350);
nor U10779 (N_10779,N_6791,N_6084);
and U10780 (N_10780,N_8964,N_8606);
nor U10781 (N_10781,N_7185,N_6361);
nand U10782 (N_10782,N_8314,N_6508);
or U10783 (N_10783,N_7023,N_6780);
nor U10784 (N_10784,N_7992,N_7099);
or U10785 (N_10785,N_6948,N_6380);
nor U10786 (N_10786,N_7945,N_6538);
or U10787 (N_10787,N_8699,N_8775);
nand U10788 (N_10788,N_6889,N_8607);
nor U10789 (N_10789,N_7011,N_6886);
nor U10790 (N_10790,N_8216,N_6798);
or U10791 (N_10791,N_8579,N_6743);
or U10792 (N_10792,N_8882,N_7423);
and U10793 (N_10793,N_6623,N_7414);
nor U10794 (N_10794,N_6442,N_6693);
and U10795 (N_10795,N_6964,N_6117);
nand U10796 (N_10796,N_8517,N_7929);
or U10797 (N_10797,N_7157,N_7661);
or U10798 (N_10798,N_7857,N_7418);
and U10799 (N_10799,N_6338,N_7154);
or U10800 (N_10800,N_6801,N_8004);
nor U10801 (N_10801,N_8769,N_7817);
or U10802 (N_10802,N_6243,N_8469);
or U10803 (N_10803,N_6430,N_7240);
or U10804 (N_10804,N_7895,N_7219);
or U10805 (N_10805,N_8722,N_6353);
nor U10806 (N_10806,N_8949,N_8518);
and U10807 (N_10807,N_6548,N_6643);
xor U10808 (N_10808,N_6292,N_6474);
and U10809 (N_10809,N_6845,N_7694);
and U10810 (N_10810,N_6942,N_6925);
or U10811 (N_10811,N_7359,N_8294);
or U10812 (N_10812,N_8535,N_7773);
nor U10813 (N_10813,N_6640,N_6623);
or U10814 (N_10814,N_6752,N_7324);
or U10815 (N_10815,N_6510,N_7628);
nor U10816 (N_10816,N_8798,N_6770);
or U10817 (N_10817,N_7487,N_7686);
xor U10818 (N_10818,N_7426,N_6069);
nor U10819 (N_10819,N_8565,N_6344);
and U10820 (N_10820,N_6392,N_6440);
nor U10821 (N_10821,N_7469,N_7672);
nor U10822 (N_10822,N_8049,N_7666);
nand U10823 (N_10823,N_7125,N_8941);
or U10824 (N_10824,N_8097,N_8977);
or U10825 (N_10825,N_6517,N_6960);
and U10826 (N_10826,N_6097,N_7256);
or U10827 (N_10827,N_7448,N_8712);
nand U10828 (N_10828,N_7287,N_7350);
nor U10829 (N_10829,N_6499,N_7515);
nand U10830 (N_10830,N_6664,N_8328);
nor U10831 (N_10831,N_8565,N_6643);
nand U10832 (N_10832,N_6186,N_6534);
nand U10833 (N_10833,N_6830,N_8804);
nor U10834 (N_10834,N_7085,N_8581);
nor U10835 (N_10835,N_6607,N_7749);
nand U10836 (N_10836,N_8855,N_8539);
and U10837 (N_10837,N_8696,N_7603);
nand U10838 (N_10838,N_7186,N_8810);
or U10839 (N_10839,N_8928,N_8551);
nor U10840 (N_10840,N_7595,N_8931);
nand U10841 (N_10841,N_6522,N_7513);
nor U10842 (N_10842,N_6602,N_8640);
nor U10843 (N_10843,N_7712,N_6377);
and U10844 (N_10844,N_8572,N_8390);
nor U10845 (N_10845,N_6985,N_8093);
nor U10846 (N_10846,N_8946,N_7204);
nor U10847 (N_10847,N_8056,N_8775);
and U10848 (N_10848,N_6150,N_8103);
nor U10849 (N_10849,N_6694,N_6277);
nand U10850 (N_10850,N_6747,N_6918);
and U10851 (N_10851,N_7443,N_6419);
or U10852 (N_10852,N_6032,N_8004);
nand U10853 (N_10853,N_8147,N_6242);
nand U10854 (N_10854,N_6046,N_7841);
nand U10855 (N_10855,N_8110,N_8628);
and U10856 (N_10856,N_8922,N_7525);
nor U10857 (N_10857,N_8857,N_7951);
nand U10858 (N_10858,N_6359,N_8129);
nand U10859 (N_10859,N_6010,N_8112);
or U10860 (N_10860,N_7528,N_8702);
nor U10861 (N_10861,N_8777,N_8710);
nand U10862 (N_10862,N_6509,N_7901);
nand U10863 (N_10863,N_8859,N_8793);
nand U10864 (N_10864,N_6189,N_6215);
and U10865 (N_10865,N_7899,N_6509);
and U10866 (N_10866,N_7096,N_6078);
or U10867 (N_10867,N_6094,N_8890);
and U10868 (N_10868,N_6842,N_6405);
nand U10869 (N_10869,N_7709,N_8759);
or U10870 (N_10870,N_8075,N_7552);
or U10871 (N_10871,N_7579,N_8642);
or U10872 (N_10872,N_8529,N_6693);
nand U10873 (N_10873,N_8899,N_8292);
nor U10874 (N_10874,N_8307,N_8846);
nor U10875 (N_10875,N_8003,N_6541);
and U10876 (N_10876,N_8379,N_8714);
nand U10877 (N_10877,N_7603,N_8221);
nand U10878 (N_10878,N_8416,N_6348);
and U10879 (N_10879,N_8506,N_6223);
nand U10880 (N_10880,N_6618,N_6154);
nand U10881 (N_10881,N_8498,N_6048);
or U10882 (N_10882,N_8232,N_7936);
nor U10883 (N_10883,N_8958,N_6417);
nand U10884 (N_10884,N_6018,N_8274);
nand U10885 (N_10885,N_7506,N_8023);
or U10886 (N_10886,N_6851,N_6540);
nor U10887 (N_10887,N_7909,N_8153);
and U10888 (N_10888,N_8336,N_7719);
nor U10889 (N_10889,N_6627,N_8549);
nand U10890 (N_10890,N_7378,N_6196);
or U10891 (N_10891,N_6923,N_6355);
nand U10892 (N_10892,N_7295,N_8956);
or U10893 (N_10893,N_7995,N_7121);
nor U10894 (N_10894,N_7930,N_8423);
nor U10895 (N_10895,N_8077,N_8995);
nand U10896 (N_10896,N_7848,N_8212);
nand U10897 (N_10897,N_6188,N_6023);
or U10898 (N_10898,N_6051,N_7204);
or U10899 (N_10899,N_6990,N_8883);
and U10900 (N_10900,N_8174,N_8944);
nor U10901 (N_10901,N_8942,N_7977);
or U10902 (N_10902,N_8678,N_7505);
and U10903 (N_10903,N_8721,N_8455);
or U10904 (N_10904,N_7777,N_8910);
nand U10905 (N_10905,N_8604,N_6484);
nor U10906 (N_10906,N_8770,N_6315);
and U10907 (N_10907,N_8771,N_8769);
or U10908 (N_10908,N_6012,N_8320);
or U10909 (N_10909,N_7606,N_8389);
nor U10910 (N_10910,N_8147,N_8447);
and U10911 (N_10911,N_7258,N_8190);
or U10912 (N_10912,N_8802,N_7012);
nand U10913 (N_10913,N_6508,N_7433);
and U10914 (N_10914,N_8325,N_7950);
nand U10915 (N_10915,N_8093,N_7366);
or U10916 (N_10916,N_7954,N_7587);
nor U10917 (N_10917,N_8271,N_8840);
nor U10918 (N_10918,N_6585,N_8582);
nand U10919 (N_10919,N_6527,N_6061);
nor U10920 (N_10920,N_6081,N_7383);
or U10921 (N_10921,N_7052,N_6123);
nand U10922 (N_10922,N_6810,N_7794);
nand U10923 (N_10923,N_8480,N_6274);
and U10924 (N_10924,N_6725,N_6489);
and U10925 (N_10925,N_6557,N_8956);
and U10926 (N_10926,N_8460,N_7410);
nand U10927 (N_10927,N_7540,N_6815);
nand U10928 (N_10928,N_7239,N_7381);
nor U10929 (N_10929,N_7285,N_7406);
nand U10930 (N_10930,N_7125,N_8194);
nand U10931 (N_10931,N_7627,N_8746);
or U10932 (N_10932,N_7218,N_8183);
nor U10933 (N_10933,N_8453,N_6702);
nor U10934 (N_10934,N_8050,N_8972);
nor U10935 (N_10935,N_6842,N_8311);
or U10936 (N_10936,N_8390,N_7233);
nor U10937 (N_10937,N_8401,N_6192);
or U10938 (N_10938,N_6961,N_8936);
nor U10939 (N_10939,N_8414,N_6416);
and U10940 (N_10940,N_8468,N_6427);
nand U10941 (N_10941,N_6711,N_6179);
and U10942 (N_10942,N_8288,N_6852);
or U10943 (N_10943,N_8430,N_6111);
nor U10944 (N_10944,N_7853,N_7859);
or U10945 (N_10945,N_8696,N_7806);
or U10946 (N_10946,N_7046,N_7470);
nor U10947 (N_10947,N_6007,N_7419);
or U10948 (N_10948,N_8757,N_6544);
and U10949 (N_10949,N_7787,N_8286);
and U10950 (N_10950,N_7358,N_8650);
nor U10951 (N_10951,N_6553,N_8637);
and U10952 (N_10952,N_8044,N_8287);
and U10953 (N_10953,N_8897,N_7150);
nor U10954 (N_10954,N_6429,N_8427);
nor U10955 (N_10955,N_7470,N_7993);
and U10956 (N_10956,N_8885,N_7883);
or U10957 (N_10957,N_7448,N_8472);
nor U10958 (N_10958,N_8915,N_8022);
or U10959 (N_10959,N_7803,N_6993);
nor U10960 (N_10960,N_8621,N_8665);
nor U10961 (N_10961,N_7732,N_7353);
or U10962 (N_10962,N_7114,N_6920);
or U10963 (N_10963,N_7903,N_6422);
nand U10964 (N_10964,N_8340,N_7040);
nor U10965 (N_10965,N_6212,N_7683);
or U10966 (N_10966,N_7300,N_7549);
nor U10967 (N_10967,N_7144,N_7137);
nor U10968 (N_10968,N_7860,N_6908);
nand U10969 (N_10969,N_7192,N_8497);
nand U10970 (N_10970,N_6069,N_7045);
nor U10971 (N_10971,N_7625,N_8279);
nor U10972 (N_10972,N_8538,N_8896);
or U10973 (N_10973,N_8037,N_6642);
and U10974 (N_10974,N_7307,N_6167);
and U10975 (N_10975,N_8833,N_7382);
and U10976 (N_10976,N_7258,N_8317);
or U10977 (N_10977,N_8595,N_7664);
nor U10978 (N_10978,N_7775,N_6425);
and U10979 (N_10979,N_6585,N_6643);
and U10980 (N_10980,N_7545,N_6967);
and U10981 (N_10981,N_8045,N_7666);
nand U10982 (N_10982,N_6326,N_8083);
or U10983 (N_10983,N_8287,N_6959);
and U10984 (N_10984,N_8589,N_8859);
or U10985 (N_10985,N_7616,N_7641);
and U10986 (N_10986,N_8047,N_8940);
nand U10987 (N_10987,N_6704,N_7280);
and U10988 (N_10988,N_8802,N_6202);
nor U10989 (N_10989,N_6530,N_6969);
nand U10990 (N_10990,N_6687,N_7303);
and U10991 (N_10991,N_7055,N_8679);
nor U10992 (N_10992,N_6060,N_7374);
and U10993 (N_10993,N_8071,N_8038);
or U10994 (N_10994,N_7411,N_8365);
and U10995 (N_10995,N_6063,N_6883);
and U10996 (N_10996,N_6106,N_6528);
nand U10997 (N_10997,N_7539,N_6699);
and U10998 (N_10998,N_8010,N_7697);
nor U10999 (N_10999,N_8407,N_6333);
nand U11000 (N_11000,N_7884,N_7374);
nand U11001 (N_11001,N_6459,N_7427);
and U11002 (N_11002,N_6665,N_6960);
nor U11003 (N_11003,N_7568,N_7670);
nor U11004 (N_11004,N_7541,N_8006);
nor U11005 (N_11005,N_8018,N_7354);
nand U11006 (N_11006,N_7651,N_7805);
or U11007 (N_11007,N_6488,N_7734);
or U11008 (N_11008,N_6606,N_6003);
and U11009 (N_11009,N_6472,N_6550);
or U11010 (N_11010,N_8311,N_6930);
nor U11011 (N_11011,N_7181,N_8054);
nand U11012 (N_11012,N_7476,N_8500);
xor U11013 (N_11013,N_6063,N_7895);
nor U11014 (N_11014,N_7706,N_8812);
or U11015 (N_11015,N_8536,N_8801);
nor U11016 (N_11016,N_8696,N_8676);
and U11017 (N_11017,N_6219,N_7691);
nand U11018 (N_11018,N_8854,N_7405);
or U11019 (N_11019,N_8443,N_6667);
nor U11020 (N_11020,N_7470,N_6408);
or U11021 (N_11021,N_8611,N_8283);
nand U11022 (N_11022,N_7120,N_6243);
or U11023 (N_11023,N_7119,N_7242);
nand U11024 (N_11024,N_6806,N_8944);
nand U11025 (N_11025,N_8526,N_7669);
nand U11026 (N_11026,N_8527,N_7797);
nand U11027 (N_11027,N_8243,N_6993);
nand U11028 (N_11028,N_7102,N_7592);
and U11029 (N_11029,N_8753,N_8006);
and U11030 (N_11030,N_8332,N_7181);
nor U11031 (N_11031,N_6237,N_6378);
or U11032 (N_11032,N_8653,N_7646);
and U11033 (N_11033,N_8217,N_8020);
and U11034 (N_11034,N_8179,N_8960);
and U11035 (N_11035,N_7464,N_6737);
and U11036 (N_11036,N_6120,N_6959);
or U11037 (N_11037,N_7290,N_8448);
nand U11038 (N_11038,N_8872,N_7192);
and U11039 (N_11039,N_8539,N_7894);
or U11040 (N_11040,N_8283,N_8446);
and U11041 (N_11041,N_8103,N_6149);
and U11042 (N_11042,N_6777,N_6226);
and U11043 (N_11043,N_6575,N_7946);
and U11044 (N_11044,N_6117,N_6228);
nand U11045 (N_11045,N_7749,N_6688);
nor U11046 (N_11046,N_6531,N_7761);
nor U11047 (N_11047,N_6152,N_7979);
and U11048 (N_11048,N_7670,N_7775);
nor U11049 (N_11049,N_8470,N_7074);
nor U11050 (N_11050,N_7535,N_8925);
and U11051 (N_11051,N_7154,N_7117);
nand U11052 (N_11052,N_6913,N_6814);
or U11053 (N_11053,N_7027,N_8776);
nand U11054 (N_11054,N_7525,N_7473);
xor U11055 (N_11055,N_7049,N_7212);
or U11056 (N_11056,N_7806,N_8894);
nand U11057 (N_11057,N_6369,N_6460);
or U11058 (N_11058,N_6702,N_7366);
or U11059 (N_11059,N_8724,N_6274);
and U11060 (N_11060,N_7818,N_6583);
or U11061 (N_11061,N_7221,N_7981);
nand U11062 (N_11062,N_7443,N_8959);
nand U11063 (N_11063,N_7824,N_8136);
nand U11064 (N_11064,N_7071,N_6313);
nand U11065 (N_11065,N_7760,N_7172);
nor U11066 (N_11066,N_7545,N_8077);
nor U11067 (N_11067,N_8281,N_7478);
or U11068 (N_11068,N_6195,N_6273);
nand U11069 (N_11069,N_8227,N_6725);
or U11070 (N_11070,N_6123,N_8450);
nand U11071 (N_11071,N_7839,N_8618);
nor U11072 (N_11072,N_7007,N_8675);
or U11073 (N_11073,N_8829,N_8663);
nand U11074 (N_11074,N_8761,N_7248);
nand U11075 (N_11075,N_7729,N_6135);
and U11076 (N_11076,N_8638,N_7909);
nor U11077 (N_11077,N_6721,N_6807);
nand U11078 (N_11078,N_7884,N_8142);
or U11079 (N_11079,N_7554,N_8568);
nand U11080 (N_11080,N_8496,N_6915);
nor U11081 (N_11081,N_8862,N_8613);
and U11082 (N_11082,N_7617,N_7683);
or U11083 (N_11083,N_6036,N_6026);
nand U11084 (N_11084,N_7346,N_8418);
nand U11085 (N_11085,N_7523,N_6826);
nor U11086 (N_11086,N_6887,N_8148);
nand U11087 (N_11087,N_8183,N_8574);
nand U11088 (N_11088,N_6025,N_6150);
and U11089 (N_11089,N_8436,N_7065);
and U11090 (N_11090,N_7832,N_8141);
and U11091 (N_11091,N_7235,N_8614);
nor U11092 (N_11092,N_8337,N_8609);
and U11093 (N_11093,N_7510,N_6677);
nor U11094 (N_11094,N_8770,N_6150);
and U11095 (N_11095,N_8959,N_6095);
and U11096 (N_11096,N_8387,N_7696);
or U11097 (N_11097,N_8737,N_6221);
nor U11098 (N_11098,N_6098,N_7781);
nand U11099 (N_11099,N_7978,N_7617);
nor U11100 (N_11100,N_6436,N_7233);
nor U11101 (N_11101,N_8567,N_6682);
nor U11102 (N_11102,N_8276,N_8133);
xor U11103 (N_11103,N_6645,N_8742);
nand U11104 (N_11104,N_7153,N_7478);
and U11105 (N_11105,N_7720,N_7145);
and U11106 (N_11106,N_7678,N_6574);
nor U11107 (N_11107,N_7469,N_6698);
nor U11108 (N_11108,N_6716,N_7372);
xnor U11109 (N_11109,N_7462,N_6495);
and U11110 (N_11110,N_8047,N_8212);
nand U11111 (N_11111,N_8803,N_8621);
nor U11112 (N_11112,N_7155,N_6324);
nor U11113 (N_11113,N_7498,N_7387);
nor U11114 (N_11114,N_8851,N_6903);
nor U11115 (N_11115,N_7754,N_8419);
or U11116 (N_11116,N_7075,N_7463);
or U11117 (N_11117,N_8859,N_7065);
or U11118 (N_11118,N_8848,N_8396);
or U11119 (N_11119,N_6728,N_8823);
or U11120 (N_11120,N_6732,N_7488);
nand U11121 (N_11121,N_8467,N_7368);
nand U11122 (N_11122,N_7239,N_8333);
nand U11123 (N_11123,N_8644,N_8426);
nor U11124 (N_11124,N_7730,N_6646);
or U11125 (N_11125,N_7393,N_8146);
nand U11126 (N_11126,N_6468,N_6054);
nor U11127 (N_11127,N_6581,N_8216);
xnor U11128 (N_11128,N_8497,N_8500);
and U11129 (N_11129,N_7081,N_8135);
nand U11130 (N_11130,N_8799,N_8207);
nor U11131 (N_11131,N_8632,N_6193);
nand U11132 (N_11132,N_8025,N_6081);
and U11133 (N_11133,N_6692,N_6761);
or U11134 (N_11134,N_8299,N_6404);
nand U11135 (N_11135,N_7946,N_7342);
or U11136 (N_11136,N_7611,N_7532);
or U11137 (N_11137,N_6557,N_8687);
or U11138 (N_11138,N_8953,N_8241);
nand U11139 (N_11139,N_8858,N_8906);
nand U11140 (N_11140,N_8093,N_8288);
and U11141 (N_11141,N_7576,N_6419);
nand U11142 (N_11142,N_7412,N_8987);
nor U11143 (N_11143,N_8918,N_7999);
and U11144 (N_11144,N_6790,N_7051);
nand U11145 (N_11145,N_6452,N_7047);
nand U11146 (N_11146,N_6965,N_8563);
or U11147 (N_11147,N_6767,N_6974);
nor U11148 (N_11148,N_8359,N_8308);
or U11149 (N_11149,N_7810,N_7116);
or U11150 (N_11150,N_6332,N_6762);
nand U11151 (N_11151,N_7508,N_7641);
nand U11152 (N_11152,N_6219,N_6232);
nor U11153 (N_11153,N_6689,N_6011);
nand U11154 (N_11154,N_8518,N_7774);
nand U11155 (N_11155,N_8233,N_6902);
nand U11156 (N_11156,N_8084,N_8021);
nand U11157 (N_11157,N_7098,N_6087);
nor U11158 (N_11158,N_8247,N_8713);
nor U11159 (N_11159,N_7837,N_6290);
nor U11160 (N_11160,N_6202,N_7074);
or U11161 (N_11161,N_6629,N_7572);
nor U11162 (N_11162,N_8479,N_8740);
nand U11163 (N_11163,N_8627,N_8366);
and U11164 (N_11164,N_8576,N_8797);
nand U11165 (N_11165,N_8838,N_6232);
nand U11166 (N_11166,N_8972,N_6367);
and U11167 (N_11167,N_7204,N_8535);
xnor U11168 (N_11168,N_7305,N_6393);
and U11169 (N_11169,N_8877,N_8378);
nor U11170 (N_11170,N_8521,N_8789);
nand U11171 (N_11171,N_8793,N_7659);
nand U11172 (N_11172,N_6576,N_6743);
and U11173 (N_11173,N_8098,N_6844);
or U11174 (N_11174,N_6088,N_7680);
nor U11175 (N_11175,N_8930,N_8534);
and U11176 (N_11176,N_8218,N_6842);
or U11177 (N_11177,N_7376,N_8592);
and U11178 (N_11178,N_7253,N_6015);
nor U11179 (N_11179,N_7866,N_6104);
nor U11180 (N_11180,N_7484,N_6154);
or U11181 (N_11181,N_7469,N_8757);
or U11182 (N_11182,N_7339,N_7010);
and U11183 (N_11183,N_6815,N_7462);
and U11184 (N_11184,N_7514,N_8754);
nor U11185 (N_11185,N_7033,N_7998);
and U11186 (N_11186,N_8652,N_7924);
or U11187 (N_11187,N_6508,N_8814);
or U11188 (N_11188,N_7046,N_8189);
nand U11189 (N_11189,N_7292,N_8670);
nand U11190 (N_11190,N_8822,N_6946);
nand U11191 (N_11191,N_6643,N_6780);
nand U11192 (N_11192,N_6376,N_6970);
nand U11193 (N_11193,N_8340,N_8527);
nor U11194 (N_11194,N_8065,N_6665);
and U11195 (N_11195,N_6889,N_8001);
and U11196 (N_11196,N_8328,N_7379);
and U11197 (N_11197,N_6074,N_7219);
and U11198 (N_11198,N_6094,N_8594);
and U11199 (N_11199,N_8132,N_8795);
nand U11200 (N_11200,N_7709,N_6675);
or U11201 (N_11201,N_8112,N_6509);
or U11202 (N_11202,N_6385,N_8274);
nand U11203 (N_11203,N_6191,N_8822);
nand U11204 (N_11204,N_6273,N_7064);
and U11205 (N_11205,N_6299,N_7079);
nor U11206 (N_11206,N_6013,N_6582);
or U11207 (N_11207,N_7425,N_7794);
nor U11208 (N_11208,N_8119,N_6628);
nor U11209 (N_11209,N_7741,N_6577);
or U11210 (N_11210,N_7896,N_8258);
and U11211 (N_11211,N_8899,N_8471);
or U11212 (N_11212,N_8723,N_8683);
and U11213 (N_11213,N_8798,N_7734);
nor U11214 (N_11214,N_8223,N_8958);
and U11215 (N_11215,N_6720,N_7621);
and U11216 (N_11216,N_8053,N_7878);
nand U11217 (N_11217,N_6818,N_6501);
nor U11218 (N_11218,N_6456,N_7358);
nor U11219 (N_11219,N_8265,N_7603);
or U11220 (N_11220,N_7155,N_7212);
or U11221 (N_11221,N_8556,N_7327);
nor U11222 (N_11222,N_7579,N_7520);
nand U11223 (N_11223,N_7104,N_7303);
or U11224 (N_11224,N_7693,N_7429);
nor U11225 (N_11225,N_7187,N_8262);
nand U11226 (N_11226,N_7215,N_8563);
and U11227 (N_11227,N_6157,N_8477);
or U11228 (N_11228,N_6375,N_6168);
nor U11229 (N_11229,N_8474,N_7841);
nor U11230 (N_11230,N_7539,N_6140);
nand U11231 (N_11231,N_7569,N_7547);
nand U11232 (N_11232,N_8471,N_6915);
nor U11233 (N_11233,N_7051,N_6553);
nor U11234 (N_11234,N_8947,N_6517);
nor U11235 (N_11235,N_7578,N_8974);
nand U11236 (N_11236,N_6421,N_6402);
and U11237 (N_11237,N_7712,N_6628);
or U11238 (N_11238,N_8131,N_7196);
xnor U11239 (N_11239,N_8610,N_8511);
nor U11240 (N_11240,N_6603,N_8405);
and U11241 (N_11241,N_8128,N_6258);
and U11242 (N_11242,N_8994,N_8295);
or U11243 (N_11243,N_7047,N_7398);
nor U11244 (N_11244,N_8785,N_7428);
and U11245 (N_11245,N_8705,N_6269);
nor U11246 (N_11246,N_7305,N_6779);
and U11247 (N_11247,N_8827,N_7700);
nor U11248 (N_11248,N_7414,N_6905);
nand U11249 (N_11249,N_8234,N_6138);
and U11250 (N_11250,N_6890,N_6102);
and U11251 (N_11251,N_7277,N_6653);
or U11252 (N_11252,N_7459,N_7419);
or U11253 (N_11253,N_7001,N_7516);
nor U11254 (N_11254,N_8195,N_7419);
or U11255 (N_11255,N_6403,N_7597);
and U11256 (N_11256,N_6269,N_7375);
xnor U11257 (N_11257,N_7681,N_7176);
nand U11258 (N_11258,N_6521,N_7048);
and U11259 (N_11259,N_7238,N_7690);
nor U11260 (N_11260,N_8941,N_6040);
and U11261 (N_11261,N_7443,N_7936);
and U11262 (N_11262,N_6780,N_6220);
nor U11263 (N_11263,N_7650,N_8938);
nor U11264 (N_11264,N_6434,N_7849);
nor U11265 (N_11265,N_8756,N_8107);
xor U11266 (N_11266,N_6178,N_6133);
and U11267 (N_11267,N_7158,N_6421);
nor U11268 (N_11268,N_7913,N_8219);
and U11269 (N_11269,N_8063,N_6998);
nand U11270 (N_11270,N_8478,N_8022);
nand U11271 (N_11271,N_7612,N_8825);
nor U11272 (N_11272,N_6201,N_7491);
and U11273 (N_11273,N_8846,N_8811);
nor U11274 (N_11274,N_8587,N_6095);
nand U11275 (N_11275,N_6975,N_6414);
or U11276 (N_11276,N_7350,N_7792);
nand U11277 (N_11277,N_6622,N_7801);
or U11278 (N_11278,N_7142,N_8940);
nor U11279 (N_11279,N_6609,N_7022);
nor U11280 (N_11280,N_8452,N_6597);
nor U11281 (N_11281,N_6256,N_6341);
nor U11282 (N_11282,N_8303,N_8705);
nand U11283 (N_11283,N_6060,N_6617);
nor U11284 (N_11284,N_7372,N_7090);
nor U11285 (N_11285,N_8337,N_7531);
nand U11286 (N_11286,N_6604,N_8102);
nand U11287 (N_11287,N_8870,N_8008);
xor U11288 (N_11288,N_7760,N_6771);
nor U11289 (N_11289,N_6502,N_8024);
xor U11290 (N_11290,N_7146,N_7958);
and U11291 (N_11291,N_6414,N_6554);
and U11292 (N_11292,N_6267,N_7638);
nor U11293 (N_11293,N_7678,N_7051);
nand U11294 (N_11294,N_6060,N_7478);
nor U11295 (N_11295,N_7059,N_8941);
nor U11296 (N_11296,N_7065,N_7543);
or U11297 (N_11297,N_8968,N_7927);
and U11298 (N_11298,N_7433,N_7194);
nand U11299 (N_11299,N_8189,N_8130);
nand U11300 (N_11300,N_6777,N_7564);
and U11301 (N_11301,N_6118,N_6457);
nor U11302 (N_11302,N_7074,N_6603);
or U11303 (N_11303,N_8056,N_6256);
or U11304 (N_11304,N_8547,N_6589);
nand U11305 (N_11305,N_6269,N_7981);
and U11306 (N_11306,N_8481,N_6654);
nor U11307 (N_11307,N_6859,N_7670);
or U11308 (N_11308,N_7588,N_7505);
nor U11309 (N_11309,N_6559,N_8279);
or U11310 (N_11310,N_6617,N_7767);
nand U11311 (N_11311,N_7137,N_7609);
xor U11312 (N_11312,N_8152,N_8325);
nor U11313 (N_11313,N_6098,N_6296);
nand U11314 (N_11314,N_7077,N_7945);
nand U11315 (N_11315,N_6493,N_7733);
nand U11316 (N_11316,N_6945,N_6479);
or U11317 (N_11317,N_6312,N_8281);
or U11318 (N_11318,N_6713,N_7378);
nor U11319 (N_11319,N_7918,N_7857);
and U11320 (N_11320,N_7895,N_8912);
nand U11321 (N_11321,N_8754,N_6735);
nand U11322 (N_11322,N_8184,N_8582);
nand U11323 (N_11323,N_7599,N_7545);
nor U11324 (N_11324,N_8772,N_8885);
or U11325 (N_11325,N_6505,N_6571);
xor U11326 (N_11326,N_8403,N_6746);
or U11327 (N_11327,N_7282,N_7407);
and U11328 (N_11328,N_6328,N_8813);
nand U11329 (N_11329,N_6874,N_7259);
nor U11330 (N_11330,N_6528,N_7345);
nor U11331 (N_11331,N_6347,N_6345);
xnor U11332 (N_11332,N_8952,N_6270);
or U11333 (N_11333,N_6272,N_7315);
nand U11334 (N_11334,N_6653,N_6376);
and U11335 (N_11335,N_6989,N_6208);
nand U11336 (N_11336,N_8066,N_8222);
nand U11337 (N_11337,N_8754,N_7457);
nand U11338 (N_11338,N_7063,N_7617);
nand U11339 (N_11339,N_8636,N_7358);
and U11340 (N_11340,N_6775,N_6500);
nand U11341 (N_11341,N_8883,N_7079);
or U11342 (N_11342,N_7662,N_8232);
and U11343 (N_11343,N_6116,N_8098);
nor U11344 (N_11344,N_8349,N_7781);
nand U11345 (N_11345,N_8277,N_8876);
nor U11346 (N_11346,N_7467,N_8954);
nand U11347 (N_11347,N_7705,N_8200);
nor U11348 (N_11348,N_6565,N_8209);
nor U11349 (N_11349,N_8204,N_6580);
nand U11350 (N_11350,N_8702,N_7974);
or U11351 (N_11351,N_6452,N_7170);
or U11352 (N_11352,N_6875,N_7412);
and U11353 (N_11353,N_7655,N_7211);
or U11354 (N_11354,N_7264,N_6115);
and U11355 (N_11355,N_6695,N_6447);
nand U11356 (N_11356,N_7757,N_7169);
or U11357 (N_11357,N_6778,N_8608);
nor U11358 (N_11358,N_7735,N_8717);
and U11359 (N_11359,N_6721,N_7131);
nor U11360 (N_11360,N_6039,N_7460);
nor U11361 (N_11361,N_7624,N_8585);
nor U11362 (N_11362,N_6679,N_6825);
and U11363 (N_11363,N_7732,N_6311);
nor U11364 (N_11364,N_8731,N_6649);
nor U11365 (N_11365,N_6188,N_6031);
or U11366 (N_11366,N_7231,N_6407);
nor U11367 (N_11367,N_8680,N_7874);
nand U11368 (N_11368,N_8501,N_6282);
and U11369 (N_11369,N_8922,N_6578);
nand U11370 (N_11370,N_8393,N_8448);
or U11371 (N_11371,N_7290,N_6803);
nand U11372 (N_11372,N_6783,N_8184);
and U11373 (N_11373,N_8551,N_6147);
xor U11374 (N_11374,N_6523,N_6104);
or U11375 (N_11375,N_6460,N_8038);
and U11376 (N_11376,N_8585,N_6215);
and U11377 (N_11377,N_6958,N_7916);
or U11378 (N_11378,N_7426,N_8818);
nor U11379 (N_11379,N_7299,N_7724);
or U11380 (N_11380,N_7741,N_8467);
nand U11381 (N_11381,N_8820,N_6636);
nor U11382 (N_11382,N_8976,N_7908);
nor U11383 (N_11383,N_7186,N_8866);
nor U11384 (N_11384,N_7107,N_7344);
or U11385 (N_11385,N_8078,N_6333);
nor U11386 (N_11386,N_8117,N_8499);
nor U11387 (N_11387,N_8468,N_8319);
nor U11388 (N_11388,N_7838,N_7013);
and U11389 (N_11389,N_6294,N_6188);
nor U11390 (N_11390,N_6278,N_6059);
and U11391 (N_11391,N_6462,N_8552);
nor U11392 (N_11392,N_6659,N_8041);
nand U11393 (N_11393,N_6285,N_6491);
nand U11394 (N_11394,N_6287,N_7788);
nand U11395 (N_11395,N_8874,N_6481);
and U11396 (N_11396,N_6260,N_7618);
nor U11397 (N_11397,N_7994,N_7526);
nor U11398 (N_11398,N_6612,N_7820);
and U11399 (N_11399,N_6701,N_8740);
or U11400 (N_11400,N_7894,N_6778);
xor U11401 (N_11401,N_6021,N_8818);
nor U11402 (N_11402,N_7000,N_6075);
nor U11403 (N_11403,N_8055,N_6698);
nor U11404 (N_11404,N_6114,N_8365);
nand U11405 (N_11405,N_7966,N_8625);
and U11406 (N_11406,N_8761,N_6675);
and U11407 (N_11407,N_7813,N_8487);
nor U11408 (N_11408,N_8318,N_6755);
nor U11409 (N_11409,N_7265,N_8730);
and U11410 (N_11410,N_7058,N_8287);
and U11411 (N_11411,N_8681,N_8257);
nand U11412 (N_11412,N_8294,N_8792);
nor U11413 (N_11413,N_8209,N_7584);
or U11414 (N_11414,N_6790,N_6049);
or U11415 (N_11415,N_6769,N_6314);
nand U11416 (N_11416,N_8550,N_7646);
nand U11417 (N_11417,N_7960,N_8283);
or U11418 (N_11418,N_8044,N_7758);
xnor U11419 (N_11419,N_8597,N_8859);
nand U11420 (N_11420,N_7711,N_7533);
nor U11421 (N_11421,N_7610,N_7855);
and U11422 (N_11422,N_6475,N_8215);
or U11423 (N_11423,N_8871,N_6878);
nand U11424 (N_11424,N_6227,N_8850);
nor U11425 (N_11425,N_6509,N_8004);
or U11426 (N_11426,N_8200,N_6577);
or U11427 (N_11427,N_6784,N_7372);
nor U11428 (N_11428,N_6676,N_6185);
nor U11429 (N_11429,N_6786,N_6040);
or U11430 (N_11430,N_6277,N_7755);
or U11431 (N_11431,N_6378,N_8096);
or U11432 (N_11432,N_8639,N_8950);
or U11433 (N_11433,N_8674,N_8839);
nor U11434 (N_11434,N_8580,N_7190);
nor U11435 (N_11435,N_6257,N_8661);
and U11436 (N_11436,N_8728,N_8614);
and U11437 (N_11437,N_7965,N_6577);
nor U11438 (N_11438,N_8343,N_8470);
and U11439 (N_11439,N_7640,N_7325);
nand U11440 (N_11440,N_8641,N_6937);
nor U11441 (N_11441,N_8829,N_7389);
nand U11442 (N_11442,N_8368,N_8586);
and U11443 (N_11443,N_8625,N_6058);
or U11444 (N_11444,N_6417,N_7019);
or U11445 (N_11445,N_6472,N_7649);
and U11446 (N_11446,N_7162,N_8893);
nor U11447 (N_11447,N_7144,N_7204);
nand U11448 (N_11448,N_7572,N_6590);
nand U11449 (N_11449,N_8872,N_7470);
or U11450 (N_11450,N_7554,N_6154);
nor U11451 (N_11451,N_8588,N_6526);
nand U11452 (N_11452,N_7877,N_8340);
nand U11453 (N_11453,N_6657,N_8073);
and U11454 (N_11454,N_7599,N_6459);
and U11455 (N_11455,N_6520,N_6475);
or U11456 (N_11456,N_7567,N_7735);
nor U11457 (N_11457,N_7121,N_7019);
and U11458 (N_11458,N_7825,N_7054);
nor U11459 (N_11459,N_6227,N_6957);
nand U11460 (N_11460,N_7206,N_6689);
nor U11461 (N_11461,N_8484,N_7145);
and U11462 (N_11462,N_6044,N_8328);
nor U11463 (N_11463,N_8775,N_7027);
nand U11464 (N_11464,N_7172,N_8780);
and U11465 (N_11465,N_8875,N_7237);
or U11466 (N_11466,N_7365,N_7020);
or U11467 (N_11467,N_6838,N_8815);
and U11468 (N_11468,N_6420,N_8850);
nor U11469 (N_11469,N_8189,N_8299);
nand U11470 (N_11470,N_6222,N_7818);
and U11471 (N_11471,N_6306,N_6983);
or U11472 (N_11472,N_7491,N_8080);
or U11473 (N_11473,N_6148,N_8588);
nand U11474 (N_11474,N_8054,N_7355);
nor U11475 (N_11475,N_8871,N_7675);
nor U11476 (N_11476,N_6990,N_7850);
nor U11477 (N_11477,N_6618,N_7310);
nand U11478 (N_11478,N_7568,N_8103);
and U11479 (N_11479,N_7687,N_7871);
nand U11480 (N_11480,N_7500,N_7849);
or U11481 (N_11481,N_7880,N_6118);
nand U11482 (N_11482,N_8802,N_7787);
nand U11483 (N_11483,N_7804,N_6938);
or U11484 (N_11484,N_6217,N_8693);
and U11485 (N_11485,N_8248,N_6205);
and U11486 (N_11486,N_8480,N_8320);
or U11487 (N_11487,N_6217,N_6929);
or U11488 (N_11488,N_7807,N_6334);
nand U11489 (N_11489,N_8858,N_8983);
nor U11490 (N_11490,N_6350,N_8366);
or U11491 (N_11491,N_7354,N_7634);
and U11492 (N_11492,N_6047,N_7416);
nor U11493 (N_11493,N_8504,N_7389);
or U11494 (N_11494,N_8000,N_8597);
nor U11495 (N_11495,N_7168,N_8090);
xor U11496 (N_11496,N_6413,N_8221);
nand U11497 (N_11497,N_6028,N_6060);
or U11498 (N_11498,N_8603,N_7669);
nor U11499 (N_11499,N_7853,N_8028);
nand U11500 (N_11500,N_6125,N_6008);
or U11501 (N_11501,N_6747,N_8422);
or U11502 (N_11502,N_6323,N_7474);
or U11503 (N_11503,N_7105,N_7629);
or U11504 (N_11504,N_8274,N_6496);
or U11505 (N_11505,N_7314,N_6876);
nand U11506 (N_11506,N_8817,N_6711);
nand U11507 (N_11507,N_6473,N_7115);
or U11508 (N_11508,N_7626,N_7790);
and U11509 (N_11509,N_7887,N_7461);
nand U11510 (N_11510,N_8505,N_8964);
or U11511 (N_11511,N_8105,N_7144);
or U11512 (N_11512,N_8312,N_8402);
or U11513 (N_11513,N_6250,N_7668);
nand U11514 (N_11514,N_6015,N_7172);
xor U11515 (N_11515,N_7709,N_8606);
nand U11516 (N_11516,N_6452,N_7281);
nand U11517 (N_11517,N_7884,N_7655);
or U11518 (N_11518,N_6271,N_6269);
nor U11519 (N_11519,N_8891,N_7808);
nor U11520 (N_11520,N_7503,N_6373);
or U11521 (N_11521,N_6012,N_8603);
nand U11522 (N_11522,N_8461,N_6683);
and U11523 (N_11523,N_7902,N_8112);
or U11524 (N_11524,N_6862,N_8583);
nor U11525 (N_11525,N_8922,N_7882);
nand U11526 (N_11526,N_6536,N_8611);
nor U11527 (N_11527,N_6371,N_7533);
or U11528 (N_11528,N_8724,N_7570);
nor U11529 (N_11529,N_7661,N_8560);
and U11530 (N_11530,N_7505,N_7962);
or U11531 (N_11531,N_8347,N_8246);
or U11532 (N_11532,N_7203,N_6308);
and U11533 (N_11533,N_8099,N_8141);
nor U11534 (N_11534,N_6380,N_6780);
and U11535 (N_11535,N_8588,N_7593);
nand U11536 (N_11536,N_7304,N_8184);
and U11537 (N_11537,N_7890,N_8119);
or U11538 (N_11538,N_7676,N_8443);
nor U11539 (N_11539,N_6963,N_6816);
nor U11540 (N_11540,N_6465,N_7651);
or U11541 (N_11541,N_8051,N_7206);
nand U11542 (N_11542,N_8577,N_6217);
nor U11543 (N_11543,N_6746,N_6962);
nor U11544 (N_11544,N_6421,N_7925);
nor U11545 (N_11545,N_7234,N_8759);
and U11546 (N_11546,N_8611,N_7705);
nor U11547 (N_11547,N_8754,N_8627);
nor U11548 (N_11548,N_7574,N_6622);
and U11549 (N_11549,N_7385,N_7566);
nor U11550 (N_11550,N_7787,N_8291);
and U11551 (N_11551,N_6008,N_6260);
or U11552 (N_11552,N_7447,N_6916);
nor U11553 (N_11553,N_6619,N_6433);
and U11554 (N_11554,N_8737,N_8370);
or U11555 (N_11555,N_6617,N_7618);
and U11556 (N_11556,N_8921,N_6683);
or U11557 (N_11557,N_7430,N_7090);
and U11558 (N_11558,N_7205,N_8882);
and U11559 (N_11559,N_6482,N_8128);
or U11560 (N_11560,N_8253,N_6166);
and U11561 (N_11561,N_6362,N_7296);
or U11562 (N_11562,N_8291,N_6767);
nor U11563 (N_11563,N_7433,N_7712);
nand U11564 (N_11564,N_6376,N_8069);
nor U11565 (N_11565,N_7057,N_7619);
nor U11566 (N_11566,N_7723,N_7981);
and U11567 (N_11567,N_8236,N_6523);
nand U11568 (N_11568,N_8942,N_7865);
nor U11569 (N_11569,N_6276,N_6864);
nand U11570 (N_11570,N_7483,N_8638);
or U11571 (N_11571,N_8280,N_7499);
nor U11572 (N_11572,N_7679,N_6554);
nor U11573 (N_11573,N_7077,N_7701);
or U11574 (N_11574,N_8172,N_6374);
nand U11575 (N_11575,N_8443,N_7131);
and U11576 (N_11576,N_7659,N_6754);
nand U11577 (N_11577,N_8201,N_8770);
nand U11578 (N_11578,N_6903,N_6132);
and U11579 (N_11579,N_7504,N_7537);
and U11580 (N_11580,N_7818,N_7634);
or U11581 (N_11581,N_6828,N_7217);
nor U11582 (N_11582,N_6615,N_7023);
xnor U11583 (N_11583,N_6320,N_6810);
and U11584 (N_11584,N_7742,N_8089);
and U11585 (N_11585,N_7745,N_6406);
or U11586 (N_11586,N_8319,N_8858);
and U11587 (N_11587,N_6682,N_8983);
and U11588 (N_11588,N_6045,N_6915);
or U11589 (N_11589,N_6197,N_7432);
or U11590 (N_11590,N_6825,N_7664);
and U11591 (N_11591,N_6518,N_8531);
nand U11592 (N_11592,N_7129,N_7446);
or U11593 (N_11593,N_6114,N_6577);
nand U11594 (N_11594,N_8602,N_6156);
and U11595 (N_11595,N_6620,N_7066);
nor U11596 (N_11596,N_6980,N_8704);
and U11597 (N_11597,N_7018,N_8109);
and U11598 (N_11598,N_7607,N_6317);
or U11599 (N_11599,N_7643,N_8181);
or U11600 (N_11600,N_8767,N_8616);
nor U11601 (N_11601,N_7367,N_7300);
or U11602 (N_11602,N_7175,N_8077);
nor U11603 (N_11603,N_7571,N_6880);
nand U11604 (N_11604,N_7359,N_8914);
and U11605 (N_11605,N_6685,N_7459);
or U11606 (N_11606,N_6245,N_8095);
and U11607 (N_11607,N_8373,N_8294);
nand U11608 (N_11608,N_8092,N_6763);
and U11609 (N_11609,N_6940,N_6887);
nand U11610 (N_11610,N_6266,N_7179);
nand U11611 (N_11611,N_7507,N_8752);
and U11612 (N_11612,N_7580,N_6556);
and U11613 (N_11613,N_7398,N_8971);
or U11614 (N_11614,N_6542,N_7859);
or U11615 (N_11615,N_7620,N_8546);
xnor U11616 (N_11616,N_7480,N_7833);
and U11617 (N_11617,N_8878,N_7271);
nor U11618 (N_11618,N_6689,N_7674);
or U11619 (N_11619,N_6328,N_7535);
or U11620 (N_11620,N_8829,N_7860);
nand U11621 (N_11621,N_6611,N_7200);
nand U11622 (N_11622,N_7525,N_6630);
and U11623 (N_11623,N_7711,N_8780);
nand U11624 (N_11624,N_6882,N_6407);
and U11625 (N_11625,N_7321,N_6253);
nor U11626 (N_11626,N_6623,N_8022);
or U11627 (N_11627,N_7063,N_6727);
nor U11628 (N_11628,N_6649,N_7399);
nor U11629 (N_11629,N_6915,N_7078);
or U11630 (N_11630,N_6130,N_7523);
and U11631 (N_11631,N_7733,N_7324);
and U11632 (N_11632,N_7840,N_8658);
or U11633 (N_11633,N_6357,N_6469);
or U11634 (N_11634,N_6497,N_6427);
and U11635 (N_11635,N_7435,N_7261);
nor U11636 (N_11636,N_6726,N_6643);
and U11637 (N_11637,N_6081,N_6980);
and U11638 (N_11638,N_6951,N_6222);
or U11639 (N_11639,N_7034,N_7243);
nor U11640 (N_11640,N_8011,N_7215);
or U11641 (N_11641,N_6761,N_6292);
or U11642 (N_11642,N_6265,N_8106);
nand U11643 (N_11643,N_6871,N_6364);
nor U11644 (N_11644,N_7519,N_8633);
nand U11645 (N_11645,N_6170,N_7833);
or U11646 (N_11646,N_7800,N_6634);
or U11647 (N_11647,N_8618,N_7344);
and U11648 (N_11648,N_6794,N_6245);
and U11649 (N_11649,N_7791,N_7415);
nand U11650 (N_11650,N_7801,N_8389);
or U11651 (N_11651,N_6888,N_8496);
nand U11652 (N_11652,N_7510,N_7677);
nand U11653 (N_11653,N_7258,N_6585);
or U11654 (N_11654,N_8186,N_7580);
nor U11655 (N_11655,N_6071,N_8380);
and U11656 (N_11656,N_6937,N_6485);
nand U11657 (N_11657,N_7476,N_6146);
and U11658 (N_11658,N_7766,N_8613);
and U11659 (N_11659,N_6545,N_6152);
nor U11660 (N_11660,N_6368,N_8480);
nand U11661 (N_11661,N_8563,N_7087);
and U11662 (N_11662,N_6169,N_6492);
and U11663 (N_11663,N_6797,N_6387);
nor U11664 (N_11664,N_7655,N_8786);
or U11665 (N_11665,N_6066,N_7829);
and U11666 (N_11666,N_6007,N_6281);
nor U11667 (N_11667,N_8814,N_8615);
and U11668 (N_11668,N_8523,N_6506);
or U11669 (N_11669,N_6537,N_7093);
or U11670 (N_11670,N_7091,N_7858);
xnor U11671 (N_11671,N_8734,N_8281);
or U11672 (N_11672,N_8660,N_8979);
nor U11673 (N_11673,N_7368,N_8987);
or U11674 (N_11674,N_6298,N_7232);
or U11675 (N_11675,N_8661,N_7806);
and U11676 (N_11676,N_6933,N_6775);
or U11677 (N_11677,N_7766,N_8450);
nor U11678 (N_11678,N_7949,N_7896);
nand U11679 (N_11679,N_8514,N_7028);
nor U11680 (N_11680,N_8302,N_7662);
or U11681 (N_11681,N_8571,N_7540);
and U11682 (N_11682,N_6454,N_8806);
nor U11683 (N_11683,N_7654,N_8357);
and U11684 (N_11684,N_8691,N_7087);
and U11685 (N_11685,N_8078,N_8216);
nor U11686 (N_11686,N_8230,N_7471);
or U11687 (N_11687,N_8793,N_8017);
or U11688 (N_11688,N_8229,N_7167);
and U11689 (N_11689,N_6411,N_6145);
nand U11690 (N_11690,N_7456,N_7216);
or U11691 (N_11691,N_6863,N_8569);
or U11692 (N_11692,N_6418,N_8613);
or U11693 (N_11693,N_7046,N_8906);
nand U11694 (N_11694,N_8427,N_8024);
and U11695 (N_11695,N_6733,N_6515);
nor U11696 (N_11696,N_7161,N_8020);
and U11697 (N_11697,N_8202,N_7935);
and U11698 (N_11698,N_8057,N_7712);
or U11699 (N_11699,N_8783,N_7661);
or U11700 (N_11700,N_8096,N_8675);
nand U11701 (N_11701,N_8388,N_6907);
or U11702 (N_11702,N_7499,N_6183);
nand U11703 (N_11703,N_6122,N_8693);
nor U11704 (N_11704,N_7426,N_6419);
nand U11705 (N_11705,N_8198,N_7243);
or U11706 (N_11706,N_8120,N_7546);
or U11707 (N_11707,N_8577,N_7199);
nand U11708 (N_11708,N_6009,N_7617);
or U11709 (N_11709,N_8297,N_7241);
nor U11710 (N_11710,N_6202,N_6267);
and U11711 (N_11711,N_7925,N_7765);
nand U11712 (N_11712,N_6080,N_6544);
or U11713 (N_11713,N_7586,N_6107);
nor U11714 (N_11714,N_7857,N_7069);
and U11715 (N_11715,N_8053,N_7117);
nor U11716 (N_11716,N_8366,N_7906);
nor U11717 (N_11717,N_6044,N_6668);
nand U11718 (N_11718,N_8185,N_7968);
or U11719 (N_11719,N_6881,N_8628);
nor U11720 (N_11720,N_8534,N_6557);
or U11721 (N_11721,N_8873,N_8934);
nor U11722 (N_11722,N_8677,N_8481);
and U11723 (N_11723,N_8435,N_6952);
nor U11724 (N_11724,N_7990,N_8707);
nor U11725 (N_11725,N_6431,N_7281);
or U11726 (N_11726,N_6768,N_6321);
nand U11727 (N_11727,N_7395,N_8035);
or U11728 (N_11728,N_8360,N_8102);
nor U11729 (N_11729,N_8609,N_7273);
nor U11730 (N_11730,N_8312,N_7297);
nand U11731 (N_11731,N_6630,N_7933);
nand U11732 (N_11732,N_7273,N_8926);
nor U11733 (N_11733,N_8786,N_8756);
xnor U11734 (N_11734,N_7911,N_8873);
nor U11735 (N_11735,N_7295,N_7333);
nor U11736 (N_11736,N_8340,N_7682);
nand U11737 (N_11737,N_6497,N_6611);
nor U11738 (N_11738,N_8119,N_8672);
or U11739 (N_11739,N_6231,N_7018);
nand U11740 (N_11740,N_6669,N_6926);
or U11741 (N_11741,N_8340,N_7382);
or U11742 (N_11742,N_6535,N_8345);
and U11743 (N_11743,N_6407,N_8682);
nor U11744 (N_11744,N_6709,N_8220);
or U11745 (N_11745,N_6099,N_7045);
nand U11746 (N_11746,N_6195,N_8039);
nand U11747 (N_11747,N_6500,N_6148);
or U11748 (N_11748,N_8569,N_6549);
and U11749 (N_11749,N_6147,N_7642);
or U11750 (N_11750,N_6129,N_8314);
nor U11751 (N_11751,N_6538,N_7984);
nand U11752 (N_11752,N_7226,N_8920);
or U11753 (N_11753,N_6208,N_7590);
and U11754 (N_11754,N_7441,N_6604);
nor U11755 (N_11755,N_8958,N_7026);
or U11756 (N_11756,N_8919,N_6126);
or U11757 (N_11757,N_6793,N_7911);
nand U11758 (N_11758,N_8569,N_8895);
or U11759 (N_11759,N_6761,N_7056);
nand U11760 (N_11760,N_8402,N_6878);
and U11761 (N_11761,N_7142,N_6674);
nand U11762 (N_11762,N_6967,N_8822);
nand U11763 (N_11763,N_6759,N_8000);
and U11764 (N_11764,N_7183,N_8161);
nor U11765 (N_11765,N_7624,N_7941);
nor U11766 (N_11766,N_8038,N_7767);
or U11767 (N_11767,N_7626,N_8955);
nand U11768 (N_11768,N_8611,N_7954);
nor U11769 (N_11769,N_6228,N_8136);
nor U11770 (N_11770,N_6011,N_6817);
xnor U11771 (N_11771,N_6656,N_6820);
and U11772 (N_11772,N_6489,N_8898);
or U11773 (N_11773,N_7639,N_7180);
and U11774 (N_11774,N_7453,N_8993);
or U11775 (N_11775,N_8485,N_8493);
or U11776 (N_11776,N_7265,N_7797);
and U11777 (N_11777,N_7352,N_6984);
or U11778 (N_11778,N_7596,N_6676);
nor U11779 (N_11779,N_7200,N_8824);
or U11780 (N_11780,N_8332,N_6380);
nand U11781 (N_11781,N_8036,N_8718);
nand U11782 (N_11782,N_7131,N_6682);
nor U11783 (N_11783,N_7325,N_7898);
or U11784 (N_11784,N_7831,N_6265);
or U11785 (N_11785,N_6245,N_6761);
nand U11786 (N_11786,N_7928,N_8392);
nor U11787 (N_11787,N_7892,N_8698);
nor U11788 (N_11788,N_8197,N_8864);
and U11789 (N_11789,N_6872,N_8915);
or U11790 (N_11790,N_8272,N_7073);
or U11791 (N_11791,N_8144,N_8126);
and U11792 (N_11792,N_7094,N_6498);
nor U11793 (N_11793,N_8193,N_7073);
nand U11794 (N_11794,N_8671,N_7971);
nand U11795 (N_11795,N_6988,N_8095);
nor U11796 (N_11796,N_7759,N_6164);
nor U11797 (N_11797,N_8448,N_7098);
nor U11798 (N_11798,N_8281,N_6904);
and U11799 (N_11799,N_6338,N_8922);
or U11800 (N_11800,N_8951,N_8210);
nand U11801 (N_11801,N_6548,N_7195);
or U11802 (N_11802,N_8898,N_8606);
nor U11803 (N_11803,N_7332,N_7652);
and U11804 (N_11804,N_7871,N_7962);
and U11805 (N_11805,N_7211,N_6280);
and U11806 (N_11806,N_8855,N_6503);
or U11807 (N_11807,N_6909,N_8959);
or U11808 (N_11808,N_6541,N_7634);
nand U11809 (N_11809,N_6793,N_6220);
and U11810 (N_11810,N_6620,N_6198);
nor U11811 (N_11811,N_7235,N_6531);
and U11812 (N_11812,N_7386,N_8980);
nand U11813 (N_11813,N_8410,N_7196);
or U11814 (N_11814,N_7388,N_8914);
and U11815 (N_11815,N_7153,N_7680);
or U11816 (N_11816,N_7374,N_6863);
nand U11817 (N_11817,N_7103,N_8718);
nand U11818 (N_11818,N_7210,N_6859);
xnor U11819 (N_11819,N_8298,N_8698);
nor U11820 (N_11820,N_7242,N_8271);
or U11821 (N_11821,N_8443,N_7538);
or U11822 (N_11822,N_7917,N_6369);
and U11823 (N_11823,N_6742,N_7276);
or U11824 (N_11824,N_7933,N_7782);
and U11825 (N_11825,N_8194,N_6678);
or U11826 (N_11826,N_8679,N_7806);
and U11827 (N_11827,N_7298,N_8115);
and U11828 (N_11828,N_8994,N_7173);
nor U11829 (N_11829,N_6849,N_7606);
and U11830 (N_11830,N_8552,N_8840);
nor U11831 (N_11831,N_6974,N_6102);
nor U11832 (N_11832,N_7838,N_6200);
nor U11833 (N_11833,N_7592,N_6578);
nor U11834 (N_11834,N_8398,N_7674);
nor U11835 (N_11835,N_8781,N_7772);
nand U11836 (N_11836,N_8638,N_7039);
or U11837 (N_11837,N_6059,N_7039);
nand U11838 (N_11838,N_7414,N_6182);
nand U11839 (N_11839,N_6309,N_7155);
or U11840 (N_11840,N_6821,N_6196);
and U11841 (N_11841,N_6351,N_6671);
or U11842 (N_11842,N_7905,N_8514);
nor U11843 (N_11843,N_6001,N_6833);
or U11844 (N_11844,N_7630,N_6545);
or U11845 (N_11845,N_7230,N_7106);
nor U11846 (N_11846,N_7394,N_6501);
nand U11847 (N_11847,N_8416,N_7632);
nand U11848 (N_11848,N_6280,N_7365);
and U11849 (N_11849,N_7015,N_7629);
and U11850 (N_11850,N_8224,N_7051);
nor U11851 (N_11851,N_6074,N_6280);
nand U11852 (N_11852,N_8507,N_6556);
nor U11853 (N_11853,N_6153,N_7074);
nand U11854 (N_11854,N_8778,N_8216);
nand U11855 (N_11855,N_6942,N_7256);
and U11856 (N_11856,N_6133,N_7471);
or U11857 (N_11857,N_6257,N_7459);
nand U11858 (N_11858,N_7731,N_6969);
nor U11859 (N_11859,N_8541,N_7437);
nor U11860 (N_11860,N_6523,N_7120);
nor U11861 (N_11861,N_6496,N_7889);
nor U11862 (N_11862,N_6458,N_7445);
or U11863 (N_11863,N_6710,N_7079);
nand U11864 (N_11864,N_8803,N_8414);
and U11865 (N_11865,N_6113,N_7581);
nor U11866 (N_11866,N_7618,N_8779);
or U11867 (N_11867,N_7893,N_8119);
or U11868 (N_11868,N_6569,N_6535);
or U11869 (N_11869,N_7238,N_8397);
nand U11870 (N_11870,N_8585,N_8034);
or U11871 (N_11871,N_6300,N_6619);
nand U11872 (N_11872,N_6465,N_7476);
nand U11873 (N_11873,N_7490,N_8912);
nor U11874 (N_11874,N_8930,N_7990);
nor U11875 (N_11875,N_7500,N_6908);
and U11876 (N_11876,N_7618,N_6680);
nor U11877 (N_11877,N_6425,N_6561);
nand U11878 (N_11878,N_7916,N_8614);
nand U11879 (N_11879,N_8832,N_8705);
or U11880 (N_11880,N_6104,N_8164);
and U11881 (N_11881,N_6535,N_6194);
nor U11882 (N_11882,N_8936,N_8931);
nor U11883 (N_11883,N_8381,N_7435);
and U11884 (N_11884,N_7985,N_7286);
or U11885 (N_11885,N_6923,N_6752);
or U11886 (N_11886,N_6873,N_7421);
nand U11887 (N_11887,N_6135,N_7153);
nand U11888 (N_11888,N_8177,N_8818);
and U11889 (N_11889,N_7584,N_8509);
and U11890 (N_11890,N_7553,N_8136);
and U11891 (N_11891,N_7287,N_8256);
or U11892 (N_11892,N_7030,N_7645);
nor U11893 (N_11893,N_6902,N_8090);
or U11894 (N_11894,N_8815,N_6799);
or U11895 (N_11895,N_6061,N_8864);
nor U11896 (N_11896,N_8106,N_8320);
nand U11897 (N_11897,N_7839,N_7354);
nor U11898 (N_11898,N_7989,N_6941);
and U11899 (N_11899,N_8140,N_7809);
and U11900 (N_11900,N_7850,N_6619);
or U11901 (N_11901,N_7681,N_7510);
and U11902 (N_11902,N_8747,N_7724);
and U11903 (N_11903,N_8288,N_7663);
nor U11904 (N_11904,N_6981,N_7941);
nor U11905 (N_11905,N_8148,N_8672);
nand U11906 (N_11906,N_7553,N_6261);
nand U11907 (N_11907,N_8029,N_6804);
nand U11908 (N_11908,N_6793,N_6533);
nor U11909 (N_11909,N_8508,N_8712);
nand U11910 (N_11910,N_8431,N_6565);
and U11911 (N_11911,N_6071,N_6461);
and U11912 (N_11912,N_6459,N_7248);
and U11913 (N_11913,N_8705,N_8684);
nand U11914 (N_11914,N_8324,N_8992);
or U11915 (N_11915,N_8127,N_6300);
or U11916 (N_11916,N_8028,N_6409);
or U11917 (N_11917,N_8880,N_7666);
nor U11918 (N_11918,N_8162,N_8896);
nor U11919 (N_11919,N_8896,N_7990);
nor U11920 (N_11920,N_7168,N_8032);
and U11921 (N_11921,N_6280,N_8012);
or U11922 (N_11922,N_7974,N_8658);
nor U11923 (N_11923,N_6150,N_7763);
nand U11924 (N_11924,N_6648,N_8450);
nor U11925 (N_11925,N_8171,N_7611);
or U11926 (N_11926,N_8384,N_6415);
or U11927 (N_11927,N_7736,N_7804);
nor U11928 (N_11928,N_7804,N_8942);
or U11929 (N_11929,N_7729,N_6634);
and U11930 (N_11930,N_6125,N_6582);
or U11931 (N_11931,N_8492,N_6118);
and U11932 (N_11932,N_6111,N_7108);
or U11933 (N_11933,N_6469,N_8533);
or U11934 (N_11934,N_6023,N_6925);
nand U11935 (N_11935,N_8708,N_6217);
and U11936 (N_11936,N_7745,N_8724);
nor U11937 (N_11937,N_6809,N_6756);
nand U11938 (N_11938,N_6592,N_6285);
nor U11939 (N_11939,N_6800,N_7361);
nand U11940 (N_11940,N_7338,N_6160);
and U11941 (N_11941,N_6618,N_6122);
nand U11942 (N_11942,N_6965,N_7684);
nand U11943 (N_11943,N_8654,N_7857);
and U11944 (N_11944,N_7812,N_8631);
or U11945 (N_11945,N_8308,N_8107);
nand U11946 (N_11946,N_6291,N_7316);
nand U11947 (N_11947,N_8766,N_7103);
nor U11948 (N_11948,N_8120,N_8073);
or U11949 (N_11949,N_6870,N_7544);
or U11950 (N_11950,N_7962,N_6055);
nand U11951 (N_11951,N_6094,N_8732);
nand U11952 (N_11952,N_7809,N_6213);
and U11953 (N_11953,N_7503,N_8620);
nor U11954 (N_11954,N_8863,N_7935);
nor U11955 (N_11955,N_7946,N_6786);
nand U11956 (N_11956,N_7451,N_6863);
and U11957 (N_11957,N_6975,N_8917);
or U11958 (N_11958,N_6663,N_8350);
and U11959 (N_11959,N_8505,N_8301);
and U11960 (N_11960,N_7930,N_6227);
nor U11961 (N_11961,N_7312,N_7992);
nand U11962 (N_11962,N_7537,N_8418);
or U11963 (N_11963,N_7327,N_6792);
nand U11964 (N_11964,N_6686,N_6879);
nor U11965 (N_11965,N_8562,N_7523);
nand U11966 (N_11966,N_7553,N_6477);
and U11967 (N_11967,N_8809,N_7801);
nor U11968 (N_11968,N_6703,N_8741);
nor U11969 (N_11969,N_6608,N_6929);
or U11970 (N_11970,N_8654,N_8224);
nand U11971 (N_11971,N_8543,N_7944);
nor U11972 (N_11972,N_8117,N_7180);
and U11973 (N_11973,N_7829,N_7164);
nand U11974 (N_11974,N_7202,N_7886);
and U11975 (N_11975,N_7298,N_8457);
nor U11976 (N_11976,N_8404,N_6607);
nor U11977 (N_11977,N_6050,N_7134);
nor U11978 (N_11978,N_6319,N_6923);
nor U11979 (N_11979,N_7814,N_6804);
nand U11980 (N_11980,N_8116,N_8399);
and U11981 (N_11981,N_6861,N_6489);
and U11982 (N_11982,N_7393,N_6310);
nand U11983 (N_11983,N_8124,N_7775);
or U11984 (N_11984,N_8345,N_8549);
nand U11985 (N_11985,N_6674,N_7604);
xor U11986 (N_11986,N_6302,N_6625);
nand U11987 (N_11987,N_7742,N_8165);
and U11988 (N_11988,N_8063,N_8335);
or U11989 (N_11989,N_6329,N_6463);
or U11990 (N_11990,N_8251,N_8301);
nand U11991 (N_11991,N_6057,N_8254);
or U11992 (N_11992,N_8569,N_8343);
nand U11993 (N_11993,N_8424,N_7064);
and U11994 (N_11994,N_8844,N_8155);
nand U11995 (N_11995,N_7937,N_7587);
nor U11996 (N_11996,N_7530,N_8406);
and U11997 (N_11997,N_6342,N_6314);
or U11998 (N_11998,N_7498,N_8377);
nor U11999 (N_11999,N_6702,N_7371);
or U12000 (N_12000,N_11287,N_10868);
or U12001 (N_12001,N_10954,N_9763);
nand U12002 (N_12002,N_11486,N_11417);
nor U12003 (N_12003,N_11386,N_9092);
or U12004 (N_12004,N_11732,N_9071);
or U12005 (N_12005,N_10154,N_9030);
or U12006 (N_12006,N_11433,N_10688);
nor U12007 (N_12007,N_9863,N_10880);
nand U12008 (N_12008,N_11166,N_9335);
nor U12009 (N_12009,N_11826,N_10651);
nand U12010 (N_12010,N_10682,N_11883);
or U12011 (N_12011,N_11077,N_10603);
and U12012 (N_12012,N_11797,N_9223);
or U12013 (N_12013,N_11507,N_10250);
or U12014 (N_12014,N_9102,N_9679);
and U12015 (N_12015,N_10198,N_9962);
nand U12016 (N_12016,N_9861,N_10658);
nand U12017 (N_12017,N_9789,N_10014);
and U12018 (N_12018,N_11154,N_9381);
nand U12019 (N_12019,N_9519,N_9716);
or U12020 (N_12020,N_9426,N_9216);
and U12021 (N_12021,N_9493,N_11435);
nand U12022 (N_12022,N_10816,N_9196);
nand U12023 (N_12023,N_9210,N_9620);
nor U12024 (N_12024,N_11312,N_9555);
nand U12025 (N_12025,N_10417,N_9820);
and U12026 (N_12026,N_9469,N_9240);
nor U12027 (N_12027,N_9358,N_9841);
and U12028 (N_12028,N_11849,N_10360);
or U12029 (N_12029,N_10452,N_11127);
and U12030 (N_12030,N_10226,N_10233);
and U12031 (N_12031,N_9914,N_11001);
nand U12032 (N_12032,N_11093,N_11179);
nand U12033 (N_12033,N_11480,N_11453);
nor U12034 (N_12034,N_11342,N_11542);
and U12035 (N_12035,N_9815,N_11650);
or U12036 (N_12036,N_9554,N_10049);
or U12037 (N_12037,N_11096,N_11873);
nor U12038 (N_12038,N_10229,N_11256);
nor U12039 (N_12039,N_10748,N_10734);
or U12040 (N_12040,N_10533,N_10013);
and U12041 (N_12041,N_9155,N_10235);
and U12042 (N_12042,N_11066,N_10369);
or U12043 (N_12043,N_9560,N_9608);
and U12044 (N_12044,N_11982,N_9219);
or U12045 (N_12045,N_10705,N_10812);
and U12046 (N_12046,N_9018,N_11167);
nor U12047 (N_12047,N_10960,N_10988);
nor U12048 (N_12048,N_9316,N_11887);
or U12049 (N_12049,N_11484,N_10917);
or U12050 (N_12050,N_11905,N_9576);
and U12051 (N_12051,N_10204,N_9984);
nor U12052 (N_12052,N_10168,N_9677);
nand U12053 (N_12053,N_9482,N_9627);
nor U12054 (N_12054,N_9070,N_11189);
nor U12055 (N_12055,N_11035,N_11334);
nor U12056 (N_12056,N_9099,N_9230);
and U12057 (N_12057,N_9543,N_11637);
or U12058 (N_12058,N_9975,N_9854);
xor U12059 (N_12059,N_9141,N_10343);
nand U12060 (N_12060,N_9334,N_10207);
or U12061 (N_12061,N_11967,N_9242);
or U12062 (N_12062,N_11393,N_11051);
nor U12063 (N_12063,N_9981,N_11536);
and U12064 (N_12064,N_9855,N_9303);
nand U12065 (N_12065,N_10984,N_10117);
or U12066 (N_12066,N_10908,N_11466);
nand U12067 (N_12067,N_10569,N_10973);
xor U12068 (N_12068,N_9600,N_10499);
or U12069 (N_12069,N_10981,N_10624);
nor U12070 (N_12070,N_10773,N_9236);
and U12071 (N_12071,N_10610,N_9321);
or U12072 (N_12072,N_9960,N_11403);
or U12073 (N_12073,N_10110,N_11860);
nand U12074 (N_12074,N_11136,N_11894);
nand U12075 (N_12075,N_10719,N_9668);
nor U12076 (N_12076,N_9691,N_11700);
nand U12077 (N_12077,N_11789,N_9501);
and U12078 (N_12078,N_9940,N_9597);
nor U12079 (N_12079,N_10510,N_11881);
nand U12080 (N_12080,N_11812,N_11016);
nand U12081 (N_12081,N_9568,N_11384);
nand U12082 (N_12082,N_10239,N_10124);
and U12083 (N_12083,N_11512,N_9735);
nand U12084 (N_12084,N_9729,N_10428);
and U12085 (N_12085,N_9400,N_10629);
and U12086 (N_12086,N_10445,N_9059);
nand U12087 (N_12087,N_9969,N_10384);
or U12088 (N_12088,N_11104,N_9314);
and U12089 (N_12089,N_9605,N_10405);
nand U12090 (N_12090,N_11635,N_11914);
nor U12091 (N_12091,N_9607,N_10644);
nor U12092 (N_12092,N_11203,N_11500);
and U12093 (N_12093,N_10485,N_10365);
and U12094 (N_12094,N_9667,N_11559);
and U12095 (N_12095,N_9165,N_10115);
or U12096 (N_12096,N_11007,N_9653);
nor U12097 (N_12097,N_9121,N_11118);
and U12098 (N_12098,N_10306,N_11761);
or U12099 (N_12099,N_11970,N_10581);
nand U12100 (N_12100,N_10677,N_10671);
and U12101 (N_12101,N_11913,N_11207);
or U12102 (N_12102,N_10656,N_11543);
or U12103 (N_12103,N_9098,N_10106);
nand U12104 (N_12104,N_10768,N_11152);
nand U12105 (N_12105,N_11090,N_10806);
nor U12106 (N_12106,N_11200,N_9376);
or U12107 (N_12107,N_11120,N_11385);
or U12108 (N_12108,N_11345,N_9159);
or U12109 (N_12109,N_9739,N_9042);
and U12110 (N_12110,N_9534,N_10664);
nand U12111 (N_12111,N_10319,N_9332);
nand U12112 (N_12112,N_9412,N_11355);
nand U12113 (N_12113,N_11545,N_10274);
nor U12114 (N_12114,N_9857,N_9272);
nand U12115 (N_12115,N_11459,N_10006);
and U12116 (N_12116,N_10669,N_9682);
nor U12117 (N_12117,N_11722,N_10446);
nand U12118 (N_12118,N_11909,N_11956);
nand U12119 (N_12119,N_9634,N_9421);
nor U12120 (N_12120,N_9034,N_9109);
nand U12121 (N_12121,N_10018,N_11827);
nor U12122 (N_12122,N_9909,N_11828);
or U12123 (N_12123,N_10711,N_9282);
or U12124 (N_12124,N_10961,N_9952);
or U12125 (N_12125,N_11874,N_11380);
nand U12126 (N_12126,N_9302,N_11735);
nand U12127 (N_12127,N_11482,N_11966);
or U12128 (N_12128,N_10573,N_9978);
or U12129 (N_12129,N_11862,N_11309);
and U12130 (N_12130,N_9447,N_10566);
or U12131 (N_12131,N_10093,N_11803);
or U12132 (N_12132,N_9517,N_9982);
and U12133 (N_12133,N_11632,N_11596);
and U12134 (N_12134,N_9930,N_9450);
and U12135 (N_12135,N_9271,N_11494);
and U12136 (N_12136,N_9858,N_10488);
nor U12137 (N_12137,N_10477,N_9963);
or U12138 (N_12138,N_11228,N_10469);
or U12139 (N_12139,N_10679,N_10759);
nor U12140 (N_12140,N_11353,N_9423);
nor U12141 (N_12141,N_11755,N_9237);
and U12142 (N_12142,N_9614,N_11788);
or U12143 (N_12143,N_9441,N_9273);
xor U12144 (N_12144,N_11156,N_10302);
nor U12145 (N_12145,N_9351,N_9557);
and U12146 (N_12146,N_11566,N_11173);
and U12147 (N_12147,N_9428,N_10251);
or U12148 (N_12148,N_11902,N_10090);
nand U12149 (N_12149,N_10043,N_11239);
and U12150 (N_12150,N_11984,N_11290);
and U12151 (N_12151,N_11135,N_11029);
nor U12152 (N_12152,N_11658,N_10256);
nand U12153 (N_12153,N_11548,N_10259);
nand U12154 (N_12154,N_9043,N_11416);
nand U12155 (N_12155,N_10301,N_11039);
nor U12156 (N_12156,N_10193,N_10991);
nor U12157 (N_12157,N_11933,N_11681);
nor U12158 (N_12158,N_10993,N_9726);
nor U12159 (N_12159,N_10326,N_10392);
nor U12160 (N_12160,N_11534,N_11616);
nand U12161 (N_12161,N_10772,N_10338);
nand U12162 (N_12162,N_9523,N_10003);
nor U12163 (N_12163,N_9499,N_10038);
and U12164 (N_12164,N_9561,N_10197);
or U12165 (N_12165,N_10820,N_10285);
or U12166 (N_12166,N_9184,N_9214);
or U12167 (N_12167,N_11861,N_10942);
nand U12168 (N_12168,N_11723,N_11428);
nand U12169 (N_12169,N_11033,N_10749);
and U12170 (N_12170,N_10680,N_10330);
nand U12171 (N_12171,N_9527,N_10733);
nor U12172 (N_12172,N_11147,N_11615);
nand U12173 (N_12173,N_9538,N_10083);
nor U12174 (N_12174,N_11574,N_11015);
nand U12175 (N_12175,N_9491,N_11864);
or U12176 (N_12176,N_11799,N_10081);
nor U12177 (N_12177,N_11145,N_9361);
nor U12178 (N_12178,N_9200,N_10930);
or U12179 (N_12179,N_10551,N_10591);
or U12180 (N_12180,N_9563,N_10946);
or U12181 (N_12181,N_11139,N_10178);
nor U12182 (N_12182,N_10766,N_9365);
nor U12183 (N_12183,N_10904,N_10780);
nand U12184 (N_12184,N_10414,N_9669);
nor U12185 (N_12185,N_10924,N_9664);
xnor U12186 (N_12186,N_11934,N_10784);
or U12187 (N_12187,N_9826,N_10964);
and U12188 (N_12188,N_9097,N_10875);
nand U12189 (N_12189,N_10934,N_9280);
nand U12190 (N_12190,N_11262,N_10713);
nand U12191 (N_12191,N_9281,N_9322);
or U12192 (N_12192,N_9442,N_9965);
nor U12193 (N_12193,N_11868,N_10706);
or U12194 (N_12194,N_9564,N_10832);
or U12195 (N_12195,N_10724,N_11124);
or U12196 (N_12196,N_11629,N_11742);
and U12197 (N_12197,N_9830,N_10609);
nor U12198 (N_12198,N_9465,N_9625);
or U12199 (N_12199,N_9736,N_11328);
nor U12200 (N_12200,N_9518,N_11734);
nand U12201 (N_12201,N_10130,N_9532);
nor U12202 (N_12202,N_9052,N_10995);
or U12203 (N_12203,N_9203,N_10148);
and U12204 (N_12204,N_11303,N_10002);
or U12205 (N_12205,N_11441,N_10577);
or U12206 (N_12206,N_10097,N_10364);
nor U12207 (N_12207,N_11892,N_9136);
and U12208 (N_12208,N_11515,N_10427);
or U12209 (N_12209,N_10670,N_10269);
nand U12210 (N_12210,N_9142,N_11644);
nor U12211 (N_12211,N_9039,N_9082);
and U12212 (N_12212,N_10096,N_9587);
xor U12213 (N_12213,N_11651,N_9166);
and U12214 (N_12214,N_11751,N_11769);
nor U12215 (N_12215,N_9119,N_10466);
or U12216 (N_12216,N_11923,N_10348);
or U12217 (N_12217,N_11140,N_10622);
or U12218 (N_12218,N_11265,N_9784);
and U12219 (N_12219,N_9911,N_9060);
and U12220 (N_12220,N_11017,N_11946);
or U12221 (N_12221,N_9101,N_11866);
and U12222 (N_12222,N_11920,N_10015);
and U12223 (N_12223,N_9602,N_10541);
nand U12224 (N_12224,N_9396,N_11058);
nor U12225 (N_12225,N_10542,N_9050);
nand U12226 (N_12226,N_9270,N_11302);
and U12227 (N_12227,N_9689,N_11927);
nand U12228 (N_12228,N_9559,N_10567);
nor U12229 (N_12229,N_10737,N_11363);
nor U12230 (N_12230,N_10983,N_9908);
or U12231 (N_12231,N_10423,N_11041);
or U12232 (N_12232,N_11606,N_11204);
nand U12233 (N_12233,N_9445,N_10896);
nor U12234 (N_12234,N_10668,N_9385);
or U12235 (N_12235,N_11641,N_9019);
nor U12236 (N_12236,N_10376,N_11037);
nand U12237 (N_12237,N_9306,N_10634);
and U12238 (N_12238,N_10728,N_11052);
nand U12239 (N_12239,N_11520,N_9842);
nand U12240 (N_12240,N_11131,N_11447);
or U12241 (N_12241,N_11977,N_9413);
nor U12242 (N_12242,N_11336,N_9081);
and U12243 (N_12243,N_9867,N_9635);
and U12244 (N_12244,N_10033,N_9521);
and U12245 (N_12245,N_11357,N_9367);
or U12246 (N_12246,N_9181,N_11772);
nor U12247 (N_12247,N_9697,N_10518);
or U12248 (N_12248,N_9250,N_11533);
and U12249 (N_12249,N_11850,N_11941);
nor U12250 (N_12250,N_10108,N_11061);
nand U12251 (N_12251,N_9730,N_11820);
and U12252 (N_12252,N_10482,N_11027);
and U12253 (N_12253,N_10559,N_9533);
nand U12254 (N_12254,N_9632,N_11325);
nor U12255 (N_12255,N_9639,N_11506);
nand U12256 (N_12256,N_11284,N_9658);
or U12257 (N_12257,N_11388,N_9284);
nor U12258 (N_12258,N_10189,N_10429);
and U12259 (N_12259,N_11177,N_9176);
and U12260 (N_12260,N_10963,N_11880);
nor U12261 (N_12261,N_10592,N_11582);
and U12262 (N_12262,N_9901,N_11579);
and U12263 (N_12263,N_9228,N_10208);
and U12264 (N_12264,N_11720,N_10279);
xnor U12265 (N_12265,N_9838,N_9710);
nor U12266 (N_12266,N_10598,N_11591);
and U12267 (N_12267,N_11815,N_9487);
nand U12268 (N_12268,N_10502,N_10025);
and U12269 (N_12269,N_9932,N_10051);
or U12270 (N_12270,N_10094,N_11298);
and U12271 (N_12271,N_9336,N_9275);
or U12272 (N_12272,N_11490,N_10861);
nand U12273 (N_12273,N_11562,N_11434);
or U12274 (N_12274,N_10347,N_9590);
or U12275 (N_12275,N_11554,N_9623);
nand U12276 (N_12276,N_9528,N_11620);
nor U12277 (N_12277,N_11472,N_9990);
nor U12278 (N_12278,N_10925,N_10635);
nand U12279 (N_12279,N_11757,N_10666);
and U12280 (N_12280,N_9440,N_10078);
or U12281 (N_12281,N_11974,N_10213);
or U12282 (N_12282,N_11219,N_10444);
and U12283 (N_12283,N_10980,N_11630);
and U12284 (N_12284,N_10951,N_10240);
or U12285 (N_12285,N_9048,N_9833);
nor U12286 (N_12286,N_11921,N_9657);
nor U12287 (N_12287,N_9399,N_10389);
nor U12288 (N_12288,N_11275,N_9254);
nand U12289 (N_12289,N_9850,N_9749);
nand U12290 (N_12290,N_11699,N_10434);
or U12291 (N_12291,N_10829,N_10987);
nand U12292 (N_12292,N_10170,N_10163);
or U12293 (N_12293,N_9645,N_11790);
or U12294 (N_12294,N_11437,N_11647);
nor U12295 (N_12295,N_9430,N_11034);
nand U12296 (N_12296,N_10493,N_10222);
nand U12297 (N_12297,N_9622,N_9531);
nor U12298 (N_12298,N_11105,N_10617);
nand U12299 (N_12299,N_10409,N_11444);
nor U12300 (N_12300,N_11009,N_10692);
nand U12301 (N_12301,N_10362,N_9156);
xnor U12302 (N_12302,N_10468,N_9129);
or U12303 (N_12303,N_10448,N_10522);
nor U12304 (N_12304,N_10216,N_11254);
and U12305 (N_12305,N_9209,N_11882);
and U12306 (N_12306,N_10704,N_9943);
or U12307 (N_12307,N_9106,N_10926);
nor U12308 (N_12308,N_11753,N_10363);
and U12309 (N_12309,N_10291,N_10877);
and U12310 (N_12310,N_9086,N_10220);
nor U12311 (N_12311,N_10643,N_9472);
xnor U12312 (N_12312,N_9797,N_10982);
or U12313 (N_12313,N_9562,N_10212);
nand U12314 (N_12314,N_9709,N_9063);
nor U12315 (N_12315,N_9859,N_10640);
nand U12316 (N_12316,N_11622,N_11288);
and U12317 (N_12317,N_9693,N_9187);
nor U12318 (N_12318,N_9067,N_11580);
or U12319 (N_12319,N_10840,N_10582);
and U12320 (N_12320,N_11940,N_9006);
and U12321 (N_12321,N_11130,N_10568);
and U12322 (N_12322,N_11704,N_9471);
or U12323 (N_12323,N_9516,N_11694);
or U12324 (N_12324,N_10823,N_11168);
and U12325 (N_12325,N_9233,N_11505);
and U12326 (N_12326,N_11429,N_11232);
nor U12327 (N_12327,N_11830,N_11918);
nand U12328 (N_12328,N_9919,N_11999);
and U12329 (N_12329,N_9725,N_9581);
nor U12330 (N_12330,N_10818,N_10919);
or U12331 (N_12331,N_11181,N_11194);
or U12332 (N_12332,N_9504,N_11642);
or U12333 (N_12333,N_9931,N_11844);
and U12334 (N_12334,N_11917,N_11981);
nand U12335 (N_12335,N_10390,N_11401);
nor U12336 (N_12336,N_11833,N_11473);
nand U12337 (N_12337,N_11646,N_10227);
and U12338 (N_12338,N_9126,N_11423);
or U12339 (N_12339,N_11611,N_10754);
nor U12340 (N_12340,N_10415,N_11258);
and U12341 (N_12341,N_11710,N_11257);
nand U12342 (N_12342,N_9765,N_10021);
nand U12343 (N_12343,N_11227,N_11365);
or U12344 (N_12344,N_11837,N_10915);
nor U12345 (N_12345,N_11906,N_10378);
and U12346 (N_12346,N_9149,N_9937);
nor U12347 (N_12347,N_11221,N_9031);
nand U12348 (N_12348,N_10703,N_10506);
or U12349 (N_12349,N_9393,N_11690);
nand U12350 (N_12350,N_11310,N_11274);
nand U12351 (N_12351,N_10177,N_9347);
or U12352 (N_12352,N_10174,N_9408);
nand U12353 (N_12353,N_10865,N_11855);
nor U12354 (N_12354,N_9825,N_9912);
nand U12355 (N_12355,N_11577,N_11889);
and U12356 (N_12356,N_10464,N_11841);
nor U12357 (N_12357,N_9705,N_9197);
nor U12358 (N_12358,N_9012,N_10492);
and U12359 (N_12359,N_11019,N_11747);
or U12360 (N_12360,N_11321,N_11285);
and U12361 (N_12361,N_10244,N_11936);
nand U12362 (N_12362,N_9434,N_9737);
or U12363 (N_12363,N_10805,N_11064);
nor U12364 (N_12364,N_11004,N_9146);
nor U12365 (N_12365,N_9738,N_10308);
nand U12366 (N_12366,N_10505,N_9460);
and U12367 (N_12367,N_10789,N_10470);
nand U12368 (N_12368,N_11108,N_9417);
or U12369 (N_12369,N_11043,N_9390);
or U12370 (N_12370,N_10138,N_11835);
or U12371 (N_12371,N_10661,N_9954);
nand U12372 (N_12372,N_10804,N_10282);
nand U12373 (N_12373,N_9733,N_11779);
nor U12374 (N_12374,N_10753,N_11020);
nand U12375 (N_12375,N_9001,N_10870);
nand U12376 (N_12376,N_10683,N_9327);
nor U12377 (N_12377,N_9721,N_10790);
nand U12378 (N_12378,N_9339,N_11176);
or U12379 (N_12379,N_11663,N_11592);
nor U12380 (N_12380,N_10091,N_11983);
nor U12381 (N_12381,N_11610,N_10828);
nor U12382 (N_12382,N_11006,N_10215);
nand U12383 (N_12383,N_10400,N_11604);
nand U12384 (N_12384,N_9026,N_9256);
nand U12385 (N_12385,N_9824,N_10322);
or U12386 (N_12386,N_11749,N_9222);
nor U12387 (N_12387,N_10752,N_11485);
nand U12388 (N_12388,N_9289,N_11252);
or U12389 (N_12389,N_10486,N_9637);
or U12390 (N_12390,N_9202,N_9551);
nand U12391 (N_12391,N_10720,N_9800);
nor U12392 (N_12392,N_10794,N_9950);
nand U12393 (N_12393,N_9466,N_11042);
and U12394 (N_12394,N_11969,N_11947);
and U12395 (N_12395,N_9897,N_9169);
nor U12396 (N_12396,N_11465,N_9353);
nand U12397 (N_12397,N_10260,N_9700);
or U12398 (N_12398,N_9619,N_9054);
and U12399 (N_12399,N_9263,N_9961);
nor U12400 (N_12400,N_9666,N_9309);
or U12401 (N_12401,N_10825,N_11564);
nand U12402 (N_12402,N_9292,N_11369);
xor U12403 (N_12403,N_9565,N_10536);
and U12404 (N_12404,N_9642,N_10885);
nor U12405 (N_12405,N_10810,N_10709);
nand U12406 (N_12406,N_10257,N_11787);
or U12407 (N_12407,N_9744,N_9446);
nor U12408 (N_12408,N_10187,N_11224);
or U12409 (N_12409,N_10950,N_10897);
and U12410 (N_12410,N_9062,N_11930);
or U12411 (N_12411,N_11959,N_11074);
or U12412 (N_12412,N_11343,N_11950);
or U12413 (N_12413,N_10026,N_10298);
nor U12414 (N_12414,N_11404,N_10192);
nand U12415 (N_12415,N_11050,N_9189);
nor U12416 (N_12416,N_10320,N_10318);
nor U12417 (N_12417,N_10529,N_9448);
and U12418 (N_12418,N_9927,N_10342);
and U12419 (N_12419,N_9206,N_9132);
or U12420 (N_12420,N_10602,N_11625);
or U12421 (N_12421,N_10611,N_10316);
nand U12422 (N_12422,N_11171,N_9552);
and U12423 (N_12423,N_11497,N_11774);
nor U12424 (N_12424,N_11421,N_9016);
nor U12425 (N_12425,N_11689,N_11952);
nor U12426 (N_12426,N_9970,N_11366);
or U12427 (N_12427,N_11904,N_10909);
and U12428 (N_12428,N_11945,N_11323);
nand U12429 (N_12429,N_10201,N_11455);
nor U12430 (N_12430,N_10283,N_10345);
or U12431 (N_12431,N_10011,N_10627);
and U12432 (N_12432,N_9384,N_11476);
nor U12433 (N_12433,N_10133,N_10850);
nand U12434 (N_12434,N_10372,N_10143);
nor U12435 (N_12435,N_10461,N_10943);
or U12436 (N_12436,N_9652,N_10103);
nand U12437 (N_12437,N_10676,N_9175);
and U12438 (N_12438,N_11858,N_10150);
nor U12439 (N_12439,N_9180,N_10167);
and U12440 (N_12440,N_9572,N_10398);
or U12441 (N_12441,N_11474,N_11280);
or U12442 (N_12442,N_11549,N_9802);
nand U12443 (N_12443,N_9756,N_10763);
nor U12444 (N_12444,N_11481,N_11511);
nand U12445 (N_12445,N_9717,N_10128);
or U12446 (N_12446,N_10895,N_11313);
and U12447 (N_12447,N_10863,N_9659);
or U12448 (N_12448,N_9477,N_10152);
nand U12449 (N_12449,N_9285,N_10795);
or U12450 (N_12450,N_10561,N_9612);
nand U12451 (N_12451,N_9049,N_9025);
or U12452 (N_12452,N_10000,N_11391);
or U12453 (N_12453,N_9922,N_10767);
or U12454 (N_12454,N_11525,N_11079);
nor U12455 (N_12455,N_11062,N_10546);
or U12456 (N_12456,N_10487,N_9939);
nor U12457 (N_12457,N_9920,N_11169);
and U12458 (N_12458,N_9371,N_11259);
and U12459 (N_12459,N_11504,N_11438);
and U12460 (N_12460,N_11085,N_9215);
or U12461 (N_12461,N_10126,N_9145);
nand U12462 (N_12462,N_11141,N_10657);
or U12463 (N_12463,N_9526,N_9752);
and U12464 (N_12464,N_11249,N_10430);
and U12465 (N_12465,N_10537,N_9740);
nor U12466 (N_12466,N_9260,N_9718);
nor U12467 (N_12467,N_10304,N_9898);
or U12468 (N_12468,N_10041,N_10095);
nand U12469 (N_12469,N_9033,N_10268);
or U12470 (N_12470,N_10479,N_11502);
or U12471 (N_12471,N_11133,N_9849);
nand U12472 (N_12472,N_11432,N_10275);
nand U12473 (N_12473,N_11277,N_11198);
or U12474 (N_12474,N_9860,N_11306);
or U12475 (N_12475,N_10141,N_9311);
nor U12476 (N_12476,N_10501,N_10911);
nand U12477 (N_12477,N_9787,N_9734);
or U12478 (N_12478,N_9732,N_10990);
or U12479 (N_12479,N_9383,N_10969);
or U12480 (N_12480,N_9964,N_11659);
nand U12481 (N_12481,N_9195,N_10262);
or U12482 (N_12482,N_11684,N_10681);
nand U12483 (N_12483,N_9529,N_10156);
xor U12484 (N_12484,N_9483,N_11854);
nor U12485 (N_12485,N_10953,N_9712);
or U12486 (N_12486,N_9300,N_9056);
nand U12487 (N_12487,N_11910,N_9976);
nor U12488 (N_12488,N_11150,N_10565);
and U12489 (N_12489,N_11399,N_11091);
nand U12490 (N_12490,N_9934,N_9722);
nor U12491 (N_12491,N_10817,N_9817);
and U12492 (N_12492,N_10967,N_10601);
nor U12493 (N_12493,N_10712,N_10102);
nand U12494 (N_12494,N_11590,N_9217);
and U12495 (N_12495,N_9702,N_11420);
nor U12496 (N_12496,N_10920,N_10439);
or U12497 (N_12497,N_11005,N_9431);
or U12498 (N_12498,N_9929,N_11202);
or U12499 (N_12499,N_11273,N_9688);
nor U12500 (N_12500,N_9151,N_10292);
nand U12501 (N_12501,N_10787,N_11780);
and U12502 (N_12502,N_11764,N_9595);
nand U12503 (N_12503,N_10513,N_11375);
nor U12504 (N_12504,N_9072,N_10238);
or U12505 (N_12505,N_11018,N_10890);
nand U12506 (N_12506,N_9706,N_10310);
or U12507 (N_12507,N_11055,N_10181);
nand U12508 (N_12508,N_9836,N_11925);
nand U12509 (N_12509,N_11733,N_10571);
and U12510 (N_12510,N_11266,N_10425);
nand U12511 (N_12511,N_10028,N_9317);
or U12512 (N_12512,N_11382,N_9397);
and U12513 (N_12513,N_9753,N_9377);
nor U12514 (N_12514,N_9877,N_9388);
nand U12515 (N_12515,N_11535,N_11551);
and U12516 (N_12516,N_10745,N_9648);
or U12517 (N_12517,N_10129,N_9192);
nor U12518 (N_12518,N_11781,N_10431);
and U12519 (N_12519,N_11065,N_10008);
and U12520 (N_12520,N_11412,N_9182);
and U12521 (N_12521,N_11031,N_10067);
nor U12522 (N_12522,N_9544,N_11282);
nor U12523 (N_12523,N_9340,N_11514);
or U12524 (N_12524,N_11899,N_10523);
and U12525 (N_12525,N_9498,N_11829);
nor U12526 (N_12526,N_9556,N_9603);
nor U12527 (N_12527,N_11419,N_11737);
or U12528 (N_12528,N_9811,N_9345);
or U12529 (N_12529,N_9462,N_10394);
nand U12530 (N_12530,N_9878,N_11993);
nor U12531 (N_12531,N_11509,N_9299);
and U12532 (N_12532,N_10489,N_11075);
nor U12533 (N_12533,N_9373,N_9246);
and U12534 (N_12534,N_9968,N_10779);
nor U12535 (N_12535,N_11957,N_11996);
and U12536 (N_12536,N_11980,N_10938);
or U12537 (N_12537,N_9636,N_10637);
and U12538 (N_12538,N_10660,N_11901);
or U12539 (N_12539,N_9890,N_11253);
or U12540 (N_12540,N_9085,N_9571);
nand U12541 (N_12541,N_10907,N_11460);
nand U12542 (N_12542,N_9768,N_9007);
and U12543 (N_12543,N_9925,N_11247);
nor U12544 (N_12544,N_9401,N_9114);
nand U12545 (N_12545,N_11541,N_9750);
nand U12546 (N_12546,N_11197,N_10898);
and U12547 (N_12547,N_11350,N_9329);
nor U12548 (N_12548,N_10972,N_11839);
nand U12549 (N_12549,N_10889,N_10922);
nand U12550 (N_12550,N_11808,N_10517);
and U12551 (N_12551,N_10809,N_10300);
and U12552 (N_12552,N_9338,N_9205);
and U12553 (N_12553,N_9856,N_11307);
or U12554 (N_12554,N_10104,N_11750);
nand U12555 (N_12555,N_10999,N_10299);
nor U12556 (N_12556,N_11628,N_10135);
and U12557 (N_12557,N_11117,N_9091);
nand U12558 (N_12558,N_10965,N_11289);
nand U12559 (N_12559,N_9244,N_11475);
nand U12560 (N_12560,N_10814,N_11724);
nand U12561 (N_12561,N_11445,N_10386);
or U12562 (N_12562,N_11161,N_11794);
nor U12563 (N_12563,N_11121,N_11107);
nor U12564 (N_12564,N_10367,N_9809);
nor U12565 (N_12565,N_11607,N_9355);
nand U12566 (N_12566,N_11978,N_10408);
nand U12567 (N_12567,N_11354,N_9125);
or U12568 (N_12568,N_10272,N_9795);
nand U12569 (N_12569,N_9133,N_11032);
or U12570 (N_12570,N_11624,N_9360);
or U12571 (N_12571,N_9610,N_11928);
nand U12572 (N_12572,N_9424,N_9578);
nand U12573 (N_12573,N_11002,N_11778);
nor U12574 (N_12574,N_9375,N_10082);
nand U12575 (N_12575,N_11195,N_10701);
nand U12576 (N_12576,N_9907,N_10689);
nand U12577 (N_12577,N_9307,N_10887);
nand U12578 (N_12578,N_10847,N_9276);
nand U12579 (N_12579,N_10005,N_10290);
and U12580 (N_12580,N_10830,N_10387);
and U12581 (N_12581,N_10055,N_9261);
nand U12582 (N_12582,N_9695,N_11718);
and U12583 (N_12583,N_11633,N_11144);
and U12584 (N_12584,N_10037,N_11226);
and U12585 (N_12585,N_10871,N_11569);
and U12586 (N_12586,N_10746,N_11180);
and U12587 (N_12587,N_11488,N_11316);
nand U12588 (N_12588,N_10246,N_10309);
nor U12589 (N_12589,N_11396,N_11326);
and U12590 (N_12590,N_9349,N_11686);
nor U12591 (N_12591,N_9624,N_11332);
and U12592 (N_12592,N_11116,N_10088);
or U12593 (N_12593,N_9535,N_10520);
and U12594 (N_12594,N_10587,N_10080);
nor U12595 (N_12595,N_9616,N_11692);
or U12596 (N_12596,N_9579,N_10001);
or U12597 (N_12597,N_11463,N_10997);
or U12598 (N_12598,N_10048,N_11261);
nand U12599 (N_12599,N_11190,N_11711);
and U12600 (N_12600,N_11172,N_10113);
nand U12601 (N_12601,N_10280,N_10628);
nand U12602 (N_12602,N_11673,N_10985);
nor U12603 (N_12603,N_11370,N_10952);
nand U12604 (N_12604,N_9308,N_9113);
xor U12605 (N_12605,N_10750,N_11223);
or U12606 (N_12606,N_10855,N_10854);
nor U12607 (N_12607,N_11080,N_9028);
nor U12608 (N_12608,N_11600,N_11106);
or U12609 (N_12609,N_11199,N_11763);
nor U12610 (N_12610,N_10645,N_10620);
nand U12611 (N_12611,N_10525,N_9350);
and U12612 (N_12612,N_11300,N_9991);
nand U12613 (N_12613,N_9356,N_10905);
nand U12614 (N_12614,N_10757,N_11997);
and U12615 (N_12615,N_9812,N_11758);
nor U12616 (N_12616,N_10802,N_11267);
and U12617 (N_12617,N_9790,N_11318);
or U12618 (N_12618,N_10312,N_11745);
nand U12619 (N_12619,N_9185,N_10153);
nor U12620 (N_12620,N_9507,N_10380);
and U12621 (N_12621,N_10157,N_9479);
nor U12622 (N_12622,N_11122,N_11170);
or U12623 (N_12623,N_9268,N_9872);
nand U12624 (N_12624,N_10357,N_10182);
and U12625 (N_12625,N_10120,N_9999);
or U12626 (N_12626,N_11806,N_9433);
xnor U12627 (N_12627,N_10404,N_9198);
nor U12628 (N_12628,N_10714,N_11518);
or U12629 (N_12629,N_11123,N_11304);
or U12630 (N_12630,N_11440,N_9415);
nand U12631 (N_12631,N_11738,N_10483);
nand U12632 (N_12632,N_10807,N_11623);
nor U12633 (N_12633,N_11402,N_9486);
nand U12634 (N_12634,N_10844,N_11795);
and U12635 (N_12635,N_10721,N_11893);
or U12636 (N_12636,N_11553,N_11540);
nand U12637 (N_12637,N_10570,N_10421);
nor U12638 (N_12638,N_11852,N_9933);
nor U12639 (N_12639,N_10788,N_10183);
or U12640 (N_12640,N_10785,N_10532);
and U12641 (N_12641,N_9245,N_9541);
and U12642 (N_12642,N_11076,N_9032);
nand U12643 (N_12643,N_11094,N_10313);
and U12644 (N_12644,N_11400,N_9046);
nor U12645 (N_12645,N_9995,N_11163);
and U12646 (N_12646,N_11599,N_10248);
and U12647 (N_12647,N_9948,N_9851);
and U12648 (N_12648,N_9816,N_9870);
nand U12649 (N_12649,N_9495,N_9599);
nand U12650 (N_12650,N_10743,N_10254);
nor U12651 (N_12651,N_11426,N_10891);
nor U12652 (N_12652,N_11397,N_10155);
nor U12653 (N_12653,N_10914,N_9882);
or U12654 (N_12654,N_11613,N_9542);
or U12655 (N_12655,N_10866,N_10219);
nand U12656 (N_12656,N_11832,N_11184);
or U12657 (N_12657,N_9988,N_10626);
and U12658 (N_12658,N_11813,N_11110);
or U12659 (N_12659,N_10957,N_11814);
xnor U12660 (N_12660,N_11349,N_11557);
and U12661 (N_12661,N_11331,N_10968);
or U12662 (N_12662,N_10406,N_9760);
or U12663 (N_12663,N_9986,N_10261);
nand U12664 (N_12664,N_11736,N_10564);
nand U12665 (N_12665,N_10063,N_11519);
and U12666 (N_12666,N_11471,N_11220);
and U12667 (N_12667,N_9846,N_11817);
or U12668 (N_12668,N_9232,N_9297);
nor U12669 (N_12669,N_10112,N_10191);
nand U12670 (N_12670,N_10879,N_9685);
and U12671 (N_12671,N_11943,N_10707);
or U12672 (N_12672,N_9264,N_11965);
nor U12673 (N_12673,N_11367,N_11584);
or U12674 (N_12674,N_9207,N_11593);
nor U12675 (N_12675,N_10744,N_9036);
or U12676 (N_12676,N_11527,N_10294);
nor U12677 (N_12677,N_10132,N_10726);
or U12678 (N_12678,N_11424,N_11594);
or U12679 (N_12679,N_10190,N_11523);
and U12680 (N_12680,N_9294,N_10563);
or U12681 (N_12681,N_10179,N_9896);
or U12682 (N_12682,N_9804,N_9628);
and U12683 (N_12683,N_11225,N_11986);
or U12684 (N_12684,N_11470,N_10481);
and U12685 (N_12685,N_11614,N_11081);
nor U12686 (N_12686,N_11821,N_9631);
nor U12687 (N_12687,N_9414,N_11218);
and U12688 (N_12688,N_9138,N_10846);
or U12689 (N_12689,N_11919,N_11452);
nand U12690 (N_12690,N_10395,N_10194);
or U12691 (N_12691,N_9985,N_9286);
or U12692 (N_12692,N_9936,N_11895);
or U12693 (N_12693,N_10822,N_9662);
nand U12694 (N_12694,N_9678,N_10834);
or U12695 (N_12695,N_10010,N_11271);
and U12696 (N_12696,N_11561,N_10864);
or U12697 (N_12697,N_9253,N_11696);
nor U12698 (N_12698,N_11612,N_11293);
nor U12699 (N_12699,N_9435,N_10131);
nor U12700 (N_12700,N_10060,N_10122);
or U12701 (N_12701,N_9781,N_11665);
nand U12702 (N_12702,N_11372,N_11241);
nand U12703 (N_12703,N_10783,N_10791);
nor U12704 (N_12704,N_9906,N_9758);
and U12705 (N_12705,N_10996,N_9630);
nand U12706 (N_12706,N_11054,N_11348);
nand U12707 (N_12707,N_9152,N_10710);
or U12708 (N_12708,N_9913,N_9757);
or U12709 (N_12709,N_9037,N_11183);
and U12710 (N_12710,N_9341,N_10455);
nand U12711 (N_12711,N_9819,N_9799);
and U12712 (N_12712,N_9530,N_11602);
nand U12713 (N_12713,N_9769,N_10385);
nand U12714 (N_12714,N_10808,N_11896);
nor U12715 (N_12715,N_10619,N_10199);
nor U12716 (N_12716,N_11989,N_9591);
and U12717 (N_12717,N_9675,N_11073);
nor U12718 (N_12718,N_9550,N_11211);
or U12719 (N_12719,N_10388,N_9267);
nand U12720 (N_12720,N_11479,N_11677);
or U12721 (N_12721,N_11530,N_10184);
nand U12722 (N_12722,N_11030,N_10058);
nand U12723 (N_12723,N_9193,N_9105);
or U12724 (N_12724,N_10554,N_9893);
xnor U12725 (N_12725,N_9835,N_10327);
nor U12726 (N_12726,N_11731,N_10059);
nor U12727 (N_12727,N_11234,N_10590);
nor U12728 (N_12728,N_10447,N_9728);
and U12729 (N_12729,N_11605,N_9500);
nor U12730 (N_12730,N_10118,N_9391);
or U12731 (N_12731,N_11759,N_10084);
nor U12732 (N_12732,N_9069,N_10747);
and U12733 (N_12733,N_11299,N_11070);
nand U12734 (N_12734,N_11754,N_10399);
and U12735 (N_12735,N_11544,N_11728);
and U12736 (N_12736,N_11092,N_10371);
nor U12737 (N_12737,N_9997,N_11703);
or U12738 (N_12738,N_10729,N_10484);
and U12739 (N_12739,N_11570,N_10498);
nor U12740 (N_12740,N_10545,N_9456);
nor U12741 (N_12741,N_9582,N_9892);
and U12742 (N_12742,N_10210,N_11674);
nor U12743 (N_12743,N_9324,N_11209);
nand U12744 (N_12744,N_9298,N_11903);
nor U12745 (N_12745,N_10307,N_11801);
nand U12746 (N_12746,N_10450,N_10069);
nor U12747 (N_12747,N_11347,N_10778);
or U12748 (N_12748,N_10442,N_9161);
nand U12749 (N_12749,N_10776,N_9604);
or U12750 (N_12750,N_10228,N_9122);
or U12751 (N_12751,N_9177,N_9676);
or U12752 (N_12752,N_10243,N_11643);
and U12753 (N_12753,N_9905,N_11951);
nand U12754 (N_12754,N_11847,N_9157);
or U12755 (N_12755,N_9503,N_11645);
nand U12756 (N_12756,N_10368,N_9843);
or U12757 (N_12757,N_9000,N_11667);
and U12758 (N_12758,N_9536,N_10774);
and U12759 (N_12759,N_10979,N_10762);
or U12760 (N_12760,N_9038,N_9095);
nor U12761 (N_12761,N_10036,N_9382);
nor U12762 (N_12762,N_11119,N_9051);
nand U12763 (N_12763,N_9899,N_11912);
or U12764 (N_12764,N_11245,N_10860);
nor U12765 (N_12765,N_10443,N_9370);
and U12766 (N_12766,N_11908,N_11389);
nor U12767 (N_12767,N_9780,N_10621);
and U12768 (N_12768,N_9403,N_11890);
and U12769 (N_12769,N_10373,N_9163);
and U12770 (N_12770,N_10284,N_11182);
nor U12771 (N_12771,N_10214,N_10526);
or U12772 (N_12772,N_10151,N_10730);
or U12773 (N_12773,N_11376,N_11014);
nor U12774 (N_12774,N_10277,N_9093);
nor U12775 (N_12775,N_11657,N_10515);
nand U12776 (N_12776,N_11149,N_11201);
nor U12777 (N_12777,N_11816,N_11205);
nand U12778 (N_12778,N_10391,N_11430);
or U12779 (N_12779,N_11413,N_11068);
nor U12780 (N_12780,N_10349,N_9596);
nor U12781 (N_12781,N_9425,N_9116);
nand U12782 (N_12782,N_9333,N_11462);
nor U12783 (N_12783,N_11291,N_11766);
nor U12784 (N_12784,N_11049,N_9437);
or U12785 (N_12785,N_10584,N_11454);
or U12786 (N_12786,N_10457,N_10358);
nor U12787 (N_12787,N_10267,N_9337);
and U12788 (N_12788,N_10782,N_9941);
nor U12789 (N_12789,N_11021,N_11053);
nor U12790 (N_12790,N_10883,N_9655);
nand U12791 (N_12791,N_10087,N_10699);
nor U12792 (N_12792,N_10792,N_10196);
or U12793 (N_12793,N_11589,N_11478);
xnor U12794 (N_12794,N_11922,N_9123);
and U12795 (N_12795,N_9731,N_10494);
or U12796 (N_12796,N_11114,N_10056);
or U12797 (N_12797,N_11340,N_11408);
and U12798 (N_12798,N_10076,N_10146);
nor U12799 (N_12799,N_9621,N_10786);
or U12800 (N_12800,N_10659,N_11898);
or U12801 (N_12801,N_10716,N_10588);
or U12802 (N_12802,N_10977,N_9617);
nand U12803 (N_12803,N_9801,N_10116);
or U12804 (N_12804,N_9609,N_11063);
and U12805 (N_12805,N_11825,N_10857);
and U12806 (N_12806,N_11938,N_10068);
or U12807 (N_12807,N_11924,N_11811);
nor U12808 (N_12808,N_11409,N_10927);
and U12809 (N_12809,N_11818,N_11730);
and U12810 (N_12810,N_10615,N_11859);
nor U12811 (N_12811,N_9372,N_10004);
and U12812 (N_12812,N_9974,N_9323);
nor U12813 (N_12813,N_10323,N_9368);
nand U12814 (N_12814,N_11744,N_10955);
or U12815 (N_12815,N_11468,N_10020);
nand U12816 (N_12816,N_10739,N_11508);
or U12817 (N_12817,N_10641,N_10824);
or U12818 (N_12818,N_11339,N_10723);
or U12819 (N_12819,N_9088,N_10725);
nand U12820 (N_12820,N_11676,N_11567);
nor U12821 (N_12821,N_10606,N_9357);
nor U12822 (N_12822,N_10630,N_10558);
nand U12823 (N_12823,N_9320,N_10508);
nor U12824 (N_12824,N_10100,N_11891);
and U12825 (N_12825,N_11320,N_10831);
nand U12826 (N_12826,N_10948,N_9484);
nand U12827 (N_12827,N_11770,N_10173);
nor U12828 (N_12828,N_9650,N_10509);
nand U12829 (N_12829,N_9058,N_11588);
nand U12830 (N_12830,N_10793,N_9045);
nand U12831 (N_12831,N_9777,N_10175);
nor U12832 (N_12832,N_11425,N_11501);
or U12833 (N_12833,N_11990,N_10140);
nand U12834 (N_12834,N_9742,N_11191);
nand U12835 (N_12835,N_10030,N_11359);
xnor U12836 (N_12836,N_11648,N_9135);
nor U12837 (N_12837,N_11973,N_9147);
or U12838 (N_12838,N_11160,N_11087);
and U12839 (N_12839,N_11159,N_9453);
or U12840 (N_12840,N_11598,N_10632);
nand U12841 (N_12841,N_10211,N_10560);
nand U12842 (N_12842,N_9793,N_11371);
nand U12843 (N_12843,N_9255,N_10352);
nand U12844 (N_12844,N_11351,N_9696);
nand U12845 (N_12845,N_11538,N_9476);
or U12846 (N_12846,N_11011,N_9522);
nor U12847 (N_12847,N_11546,N_10833);
nand U12848 (N_12848,N_9586,N_11875);
nand U12849 (N_12849,N_9179,N_10631);
nand U12850 (N_12850,N_9389,N_11264);
and U12851 (N_12851,N_9884,N_10158);
nor U12852 (N_12852,N_10742,N_11877);
nand U12853 (N_12853,N_10543,N_9084);
or U12854 (N_12854,N_10451,N_9296);
nor U12855 (N_12855,N_11655,N_11856);
and U12856 (N_12856,N_10945,N_10370);
nor U12857 (N_12857,N_11477,N_10939);
and U12858 (N_12858,N_9674,N_10503);
nand U12859 (N_12859,N_9553,N_10045);
nor U12860 (N_12860,N_10162,N_10265);
or U12861 (N_12861,N_10105,N_9873);
or U12862 (N_12862,N_11581,N_10418);
and U12863 (N_12863,N_11448,N_11863);
or U12864 (N_12864,N_11573,N_10098);
nand U12865 (N_12865,N_9352,N_9497);
and U12866 (N_12866,N_9754,N_10655);
nor U12867 (N_12867,N_9828,N_9510);
and U12868 (N_12868,N_9153,N_9199);
nor U12869 (N_12869,N_9017,N_11586);
and U12870 (N_12870,N_9079,N_10449);
or U12871 (N_12871,N_9762,N_11222);
nand U12872 (N_12872,N_10022,N_9673);
nor U12873 (N_12873,N_10366,N_9569);
and U12874 (N_12874,N_9035,N_10407);
or U12875 (N_12875,N_10397,N_11666);
and U12876 (N_12876,N_9485,N_9212);
and U12877 (N_12877,N_10899,N_11188);
and U12878 (N_12878,N_11146,N_11129);
nand U12879 (N_12879,N_11158,N_11186);
nor U12880 (N_12880,N_10396,N_9183);
or U12881 (N_12881,N_9839,N_11560);
nor U12882 (N_12882,N_10777,N_10234);
nand U12883 (N_12883,N_11867,N_9363);
nand U12884 (N_12884,N_11709,N_11522);
nand U12885 (N_12885,N_9847,N_9916);
and U12886 (N_12886,N_11503,N_9840);
nor U12887 (N_12887,N_10586,N_9935);
nand U12888 (N_12888,N_11132,N_11212);
nand U12889 (N_12889,N_10413,N_11756);
nand U12890 (N_12890,N_10195,N_9162);
and U12891 (N_12891,N_9748,N_11804);
nor U12892 (N_12892,N_10217,N_10218);
or U12893 (N_12893,N_11848,N_9108);
or U12894 (N_12894,N_9513,N_10209);
and U12895 (N_12895,N_10359,N_9714);
or U12896 (N_12896,N_9348,N_9204);
and U12897 (N_12897,N_9703,N_10221);
nand U12898 (N_12898,N_11047,N_9670);
nor U12899 (N_12899,N_9137,N_11360);
nor U12900 (N_12900,N_10928,N_11702);
nand U12901 (N_12901,N_9290,N_9547);
or U12902 (N_12902,N_9759,N_10463);
or U12903 (N_12903,N_10781,N_9994);
nand U12904 (N_12904,N_9004,N_11157);
and U12905 (N_12905,N_9014,N_9761);
nand U12906 (N_12906,N_11872,N_11491);
nor U12907 (N_12907,N_9248,N_9707);
nor U12908 (N_12908,N_10862,N_11418);
or U12909 (N_12909,N_10065,N_11879);
or U12910 (N_12910,N_10801,N_11851);
nor U12911 (N_12911,N_11255,N_10356);
and U12912 (N_12912,N_9305,N_9537);
or U12913 (N_12913,N_9418,N_10636);
nor U12914 (N_12914,N_9525,N_10975);
nor U12915 (N_12915,N_11843,N_11805);
nor U12916 (N_12916,N_10333,N_9713);
or U12917 (N_12917,N_9686,N_10684);
nand U12918 (N_12918,N_9902,N_10974);
nor U12919 (N_12919,N_9224,N_10305);
nand U12920 (N_12920,N_11857,N_11729);
nand U12921 (N_12921,N_11869,N_9549);
and U12922 (N_12922,N_9459,N_9265);
nor U12923 (N_12923,N_11796,N_10769);
nand U12924 (N_12924,N_9889,N_11968);
nand U12925 (N_12925,N_11654,N_10402);
and U12926 (N_12926,N_10403,N_10944);
and U12927 (N_12927,N_10496,N_11115);
nor U12928 (N_12928,N_11457,N_10346);
nand U12929 (N_12929,N_10511,N_11143);
nand U12930 (N_12930,N_10161,N_9633);
nand U12931 (N_12931,N_10478,N_11498);
nor U12932 (N_12932,N_9387,N_10166);
nand U12933 (N_12933,N_11846,N_10740);
nor U12934 (N_12934,N_10616,N_9720);
or U12935 (N_12935,N_11489,N_9154);
and U12936 (N_12936,N_10738,N_9926);
and U12937 (N_12937,N_9987,N_10976);
nand U12938 (N_12938,N_11840,N_9269);
or U12939 (N_12939,N_11682,N_9671);
and U12940 (N_12940,N_10796,N_10881);
nand U12941 (N_12941,N_9747,N_11492);
and U12942 (N_12942,N_11760,N_9594);
or U12943 (N_12943,N_10539,N_11192);
nand U12944 (N_12944,N_9638,N_9947);
or U12945 (N_12945,N_10736,N_9888);
or U12946 (N_12946,N_11636,N_10023);
nand U12947 (N_12947,N_9680,N_9956);
or U12948 (N_12948,N_9900,N_9951);
nor U12949 (N_12949,N_11662,N_10295);
nor U12950 (N_12950,N_9301,N_11352);
nand U12951 (N_12951,N_11603,N_10476);
and U12952 (N_12952,N_9651,N_9227);
nor U12953 (N_12953,N_11374,N_9331);
and U12954 (N_12954,N_9128,N_9871);
and U12955 (N_12955,N_9715,N_9251);
nor U12956 (N_12956,N_10604,N_9078);
or U12957 (N_12957,N_10072,N_9989);
and U12958 (N_12958,N_11762,N_10555);
and U12959 (N_12959,N_10755,N_9213);
and U12960 (N_12960,N_9130,N_10200);
nand U12961 (N_12961,N_9310,N_9003);
nor U12962 (N_12962,N_9201,N_11785);
nand U12963 (N_12963,N_10382,N_11044);
nand U12964 (N_12964,N_10230,N_9661);
and U12965 (N_12965,N_11295,N_11845);
nand U12966 (N_12966,N_11008,N_11948);
or U12967 (N_12967,N_11521,N_9110);
or U12968 (N_12968,N_10495,N_10061);
or U12969 (N_12969,N_11060,N_11415);
or U12970 (N_12970,N_10293,N_10989);
and U12971 (N_12971,N_9029,N_10838);
nand U12972 (N_12972,N_11669,N_11467);
or U12973 (N_12973,N_10962,N_10270);
nand U12974 (N_12974,N_10435,N_10702);
nor U12975 (N_12975,N_11954,N_9366);
or U12976 (N_12976,N_10472,N_9681);
nor U12977 (N_12977,N_10321,N_9208);
and U12978 (N_12978,N_11410,N_10936);
nor U12979 (N_12979,N_9111,N_10614);
nand U12980 (N_12980,N_11791,N_10827);
or U12981 (N_12981,N_11853,N_10538);
or U12982 (N_12982,N_10903,N_9083);
or U12983 (N_12983,N_9803,N_9767);
and U12984 (N_12984,N_9794,N_10741);
or U12985 (N_12985,N_10514,N_9776);
nand U12986 (N_12986,N_10437,N_10432);
nand U12987 (N_12987,N_10203,N_9010);
nor U12988 (N_12988,N_9618,N_10797);
nor U12989 (N_12989,N_9822,N_10935);
and U12990 (N_12990,N_9574,N_10583);
and U12991 (N_12991,N_10147,N_11317);
or U12992 (N_12992,N_10521,N_11619);
or U12993 (N_12993,N_9649,N_10328);
nand U12994 (N_12994,N_9727,N_10311);
and U12995 (N_12995,N_11056,N_9378);
nor U12996 (N_12996,N_9883,N_9328);
nor U12997 (N_12997,N_10186,N_9998);
nor U12998 (N_12998,N_9313,N_10245);
xor U12999 (N_12999,N_11800,N_10553);
or U13000 (N_13000,N_11991,N_10596);
and U13001 (N_13001,N_10959,N_9771);
nand U13002 (N_13002,N_11134,N_10458);
nand U13003 (N_13003,N_11379,N_11783);
nor U13004 (N_13004,N_9235,N_11206);
or U13005 (N_13005,N_10420,N_9779);
nand U13006 (N_13006,N_9944,N_10241);
nor U13007 (N_13007,N_10504,N_9993);
nand U13008 (N_13008,N_9027,N_10869);
or U13009 (N_13009,N_9745,N_10035);
nor U13010 (N_13010,N_9823,N_11911);
xor U13011 (N_13011,N_10901,N_11405);
nand U13012 (N_13012,N_11653,N_11026);
or U13013 (N_13013,N_10892,N_9786);
nor U13014 (N_13014,N_10467,N_11268);
nand U13015 (N_13015,N_9090,N_9711);
nand U13016 (N_13016,N_9160,N_10460);
and U13017 (N_13017,N_9548,N_10516);
or U13018 (N_13018,N_9539,N_11422);
nand U13019 (N_13019,N_10441,N_11270);
nor U13020 (N_13020,N_10205,N_11798);
or U13021 (N_13021,N_9788,N_10764);
nand U13022 (N_13022,N_10252,N_11656);
or U13023 (N_13023,N_10708,N_10296);
nor U13024 (N_13024,N_9315,N_11939);
nor U13025 (N_13025,N_10929,N_10281);
nand U13026 (N_13026,N_9796,N_10599);
nand U13027 (N_13027,N_9848,N_11337);
and U13028 (N_13028,N_9342,N_9044);
nor U13029 (N_13029,N_10412,N_10685);
nand U13030 (N_13030,N_11069,N_10263);
or U13031 (N_13031,N_9798,N_9024);
or U13032 (N_13032,N_11528,N_11040);
and U13033 (N_13033,N_10572,N_9959);
or U13034 (N_13034,N_11784,N_9467);
nor U13035 (N_13035,N_11165,N_9394);
or U13036 (N_13036,N_10039,N_11025);
nor U13037 (N_13037,N_11344,N_10071);
xnor U13038 (N_13038,N_10528,N_10169);
nor U13039 (N_13039,N_11012,N_9875);
or U13040 (N_13040,N_11618,N_11398);
or U13041 (N_13041,N_11153,N_10044);
nand U13042 (N_13042,N_9087,N_11082);
nand U13043 (N_13043,N_10852,N_10297);
nand U13044 (N_13044,N_10337,N_9567);
and U13045 (N_13045,N_10401,N_9461);
nand U13046 (N_13046,N_11524,N_11208);
and U13047 (N_13047,N_11358,N_10998);
nor U13048 (N_13048,N_11944,N_9546);
and U13049 (N_13049,N_10480,N_11953);
nor U13050 (N_13050,N_11443,N_11450);
nand U13051 (N_13051,N_9065,N_11793);
or U13052 (N_13052,N_10841,N_10512);
nor U13053 (N_13053,N_11083,N_9047);
nor U13054 (N_13054,N_10978,N_11038);
nand U13055 (N_13055,N_10949,N_9886);
nor U13056 (N_13056,N_10639,N_11960);
and U13057 (N_13057,N_10377,N_9474);
and U13058 (N_13058,N_10206,N_10436);
or U13059 (N_13059,N_9231,N_10638);
and U13060 (N_13060,N_10700,N_10137);
nand U13061 (N_13061,N_11496,N_9915);
and U13062 (N_13062,N_11935,N_11407);
and U13063 (N_13063,N_11000,N_10597);
or U13064 (N_13064,N_9392,N_9701);
or U13065 (N_13065,N_10687,N_11022);
nand U13066 (N_13066,N_10009,N_10771);
nand U13067 (N_13067,N_9723,N_11128);
or U13068 (N_13068,N_9891,N_11719);
nor U13069 (N_13069,N_11048,N_11531);
nor U13070 (N_13070,N_11727,N_9115);
nand U13071 (N_13071,N_9188,N_11368);
and U13072 (N_13072,N_11721,N_11431);
or U13073 (N_13073,N_10941,N_10149);
or U13074 (N_13074,N_11716,N_10562);
nor U13075 (N_13075,N_11338,N_9778);
nor U13076 (N_13076,N_11237,N_11698);
and U13077 (N_13077,N_10966,N_9626);
or U13078 (N_13078,N_10017,N_10109);
and U13079 (N_13079,N_10077,N_9427);
nand U13080 (N_13080,N_9764,N_10276);
nand U13081 (N_13081,N_9983,N_10475);
nand U13082 (N_13082,N_9743,N_9672);
nor U13083 (N_13083,N_9194,N_10821);
and U13084 (N_13084,N_11138,N_10970);
and U13085 (N_13085,N_10459,N_11768);
and U13086 (N_13086,N_11876,N_9663);
nand U13087 (N_13087,N_10690,N_11926);
nor U13088 (N_13088,N_11964,N_9173);
nand U13089 (N_13089,N_9008,N_11652);
nand U13090 (N_13090,N_9443,N_11971);
nor U13091 (N_13091,N_11529,N_9545);
nor U13092 (N_13092,N_11552,N_11446);
or U13093 (N_13093,N_10139,N_11771);
and U13094 (N_13094,N_9992,N_9359);
or U13095 (N_13095,N_9076,N_10314);
nand U13096 (N_13096,N_11701,N_11885);
nor U13097 (N_13097,N_10303,N_11691);
nor U13098 (N_13098,N_11824,N_9810);
xnor U13099 (N_13099,N_11707,N_11998);
nor U13100 (N_13100,N_10101,N_10819);
nor U13101 (N_13101,N_9277,N_9226);
and U13102 (N_13102,N_10674,N_11550);
and U13103 (N_13103,N_9326,N_11609);
nor U13104 (N_13104,N_10253,N_10856);
and U13105 (N_13105,N_11929,N_9494);
or U13106 (N_13106,N_11617,N_11361);
and U13107 (N_13107,N_11726,N_9312);
or U13108 (N_13108,N_9924,N_10057);
or U13109 (N_13109,N_11099,N_11276);
nor U13110 (N_13110,N_9089,N_9118);
nand U13111 (N_13111,N_11963,N_9805);
and U13112 (N_13112,N_9640,N_9243);
and U13113 (N_13113,N_9945,N_10923);
or U13114 (N_13114,N_9444,N_9917);
or U13115 (N_13115,N_11251,N_11126);
and U13116 (N_13116,N_9894,N_10527);
and U13117 (N_13117,N_9724,N_11301);
nor U13118 (N_13118,N_11961,N_10064);
nor U13119 (N_13119,N_9644,N_9020);
or U13120 (N_13120,N_10416,N_11378);
nor U13121 (N_13121,N_10732,N_10994);
xnor U13122 (N_13122,N_10232,N_10715);
or U13123 (N_13123,N_11109,N_10837);
xnor U13124 (N_13124,N_10695,N_10836);
nor U13125 (N_13125,N_10086,N_9139);
nor U13126 (N_13126,N_9420,N_11333);
and U13127 (N_13127,N_9061,N_10910);
and U13128 (N_13128,N_11327,N_9481);
nand U13129 (N_13129,N_9478,N_9021);
nor U13130 (N_13130,N_10958,N_10134);
nand U13131 (N_13131,N_9150,N_9174);
nand U13132 (N_13132,N_9573,N_11807);
or U13133 (N_13133,N_9073,N_11907);
nand U13134 (N_13134,N_11151,N_10535);
nand U13135 (N_13135,N_11248,N_10574);
and U13136 (N_13136,N_11558,N_10507);
or U13137 (N_13137,N_11634,N_11672);
or U13138 (N_13138,N_10160,N_11842);
nor U13139 (N_13139,N_11695,N_11499);
or U13140 (N_13140,N_10381,N_11230);
and U13141 (N_13141,N_11987,N_9015);
nor U13142 (N_13142,N_10172,N_9879);
and U13143 (N_13143,N_11886,N_9834);
or U13144 (N_13144,N_11937,N_10760);
and U13145 (N_13145,N_10646,N_10099);
nor U13146 (N_13146,N_9880,N_11112);
nand U13147 (N_13147,N_11244,N_11955);
and U13148 (N_13148,N_9492,N_9953);
nand U13149 (N_13149,N_10440,N_10649);
nand U13150 (N_13150,N_10756,N_9665);
or U13151 (N_13151,N_9234,N_9966);
and U13152 (N_13152,N_9910,N_10092);
and U13153 (N_13153,N_9134,N_11746);
or U13154 (N_13154,N_9598,N_9946);
nor U13155 (N_13155,N_9170,N_9488);
nor U13156 (N_13156,N_11516,N_9996);
nor U13157 (N_13157,N_11281,N_10815);
nor U13158 (N_13158,N_9009,N_9746);
and U13159 (N_13159,N_11513,N_11314);
or U13160 (N_13160,N_10647,N_11279);
or U13161 (N_13161,N_11028,N_10317);
and U13162 (N_13162,N_10433,N_9104);
xnor U13163 (N_13163,N_9257,N_10419);
and U13164 (N_13164,N_9096,N_11324);
and U13165 (N_13165,N_9895,N_10070);
nor U13166 (N_13166,N_11098,N_11210);
and U13167 (N_13167,N_10931,N_10422);
nand U13168 (N_13168,N_11985,N_9818);
nand U13169 (N_13169,N_11162,N_11583);
or U13170 (N_13170,N_11660,N_9470);
or U13171 (N_13171,N_10940,N_10007);
and U13172 (N_13172,N_11175,N_9164);
nand U13173 (N_13173,N_11383,N_11537);
or U13174 (N_13174,N_9143,N_10286);
or U13175 (N_13175,N_11888,N_9511);
nand U13176 (N_13176,N_11627,N_9451);
or U13177 (N_13177,N_10971,N_10225);
nand U13178 (N_13178,N_10351,N_11975);
and U13179 (N_13179,N_11979,N_9279);
and U13180 (N_13180,N_10697,N_9386);
and U13181 (N_13181,N_9520,N_9611);
and U13182 (N_13182,N_10355,N_10612);
or U13183 (N_13183,N_11193,N_11568);
nand U13184 (N_13184,N_10332,N_10249);
nand U13185 (N_13185,N_11587,N_11740);
nand U13186 (N_13186,N_10544,N_9874);
nor U13187 (N_13187,N_10913,N_11078);
nand U13188 (N_13188,N_10867,N_9100);
nand U13189 (N_13189,N_9374,N_11387);
nor U13190 (N_13190,N_11680,N_10340);
and U13191 (N_13191,N_9692,N_11792);
or U13192 (N_13192,N_10344,N_11992);
and U13193 (N_13193,N_10171,N_9881);
nor U13194 (N_13194,N_11495,N_11414);
or U13195 (N_13195,N_10202,N_11319);
or U13196 (N_13196,N_10605,N_10765);
and U13197 (N_13197,N_9239,N_10811);
or U13198 (N_13198,N_9266,N_9575);
xor U13199 (N_13199,N_9958,N_11451);
nand U13200 (N_13200,N_10956,N_10916);
and U13201 (N_13201,N_11296,N_11097);
nand U13202 (N_13202,N_9274,N_9186);
nor U13203 (N_13203,N_10698,N_10751);
nand U13204 (N_13204,N_10845,N_11767);
and U13205 (N_13205,N_11532,N_9719);
nor U13206 (N_13206,N_9077,N_9829);
nor U13207 (N_13207,N_11526,N_11113);
nand U13208 (N_13208,N_10937,N_10266);
and U13209 (N_13209,N_10694,N_11838);
nand U13210 (N_13210,N_9585,N_10652);
nand U13211 (N_13211,N_10032,N_11900);
xnor U13212 (N_13212,N_11743,N_11216);
and U13213 (N_13213,N_10851,N_10575);
nand U13214 (N_13214,N_11003,N_11449);
nand U13215 (N_13215,N_10608,N_11931);
and U13216 (N_13216,N_11972,N_9684);
or U13217 (N_13217,N_11229,N_10888);
or U13218 (N_13218,N_11571,N_9053);
nand U13219 (N_13219,N_11988,N_11563);
and U13220 (N_13220,N_10594,N_11263);
nor U13221 (N_13221,N_9791,N_11362);
and U13222 (N_13222,N_9429,N_9362);
nand U13223 (N_13223,N_10933,N_9354);
nand U13224 (N_13224,N_9304,N_10237);
or U13225 (N_13225,N_11576,N_11715);
or U13226 (N_13226,N_11067,N_11390);
nor U13227 (N_13227,N_11297,N_11059);
nand U13228 (N_13228,N_10085,N_11329);
or U13229 (N_13229,N_10231,N_11897);
nor U13230 (N_13230,N_9409,N_10799);
xnor U13231 (N_13231,N_9364,N_11010);
nand U13232 (N_13232,N_9057,N_9404);
and U13233 (N_13233,N_9458,N_9775);
nor U13234 (N_13234,N_11311,N_9865);
or U13235 (N_13235,N_9783,N_11777);
nor U13236 (N_13236,N_11394,N_11238);
nand U13237 (N_13237,N_10633,N_10136);
nor U13238 (N_13238,N_10549,N_10034);
or U13239 (N_13239,N_9406,N_10900);
and U13240 (N_13240,N_10111,N_9422);
or U13241 (N_13241,N_11250,N_9864);
nand U13242 (N_13242,N_10653,N_10672);
nor U13243 (N_13243,N_9124,N_10165);
nand U13244 (N_13244,N_11565,N_9704);
or U13245 (N_13245,N_9094,N_11556);
nand U13246 (N_13246,N_10379,N_9040);
or U13247 (N_13247,N_11765,N_11725);
nand U13248 (N_13248,N_9463,N_10107);
and U13249 (N_13249,N_9770,N_11517);
or U13250 (N_13250,N_10424,N_11802);
nand U13251 (N_13251,N_10607,N_9080);
or U13252 (N_13252,N_9751,N_9853);
or U13253 (N_13253,N_9660,N_11621);
nor U13254 (N_13254,N_9887,N_10329);
or U13255 (N_13255,N_11292,N_9013);
nor U13256 (N_13256,N_11510,N_9808);
nand U13257 (N_13257,N_11575,N_9694);
and U13258 (N_13258,N_10053,N_9772);
nand U13259 (N_13259,N_11706,N_9514);
nand U13260 (N_13260,N_11687,N_9687);
nor U13261 (N_13261,N_11377,N_10717);
or U13262 (N_13262,N_9741,N_9869);
and U13263 (N_13263,N_11214,N_9319);
nor U13264 (N_13264,N_9593,N_10079);
and U13265 (N_13265,N_11236,N_10471);
nor U13266 (N_13266,N_9171,N_9904);
nor U13267 (N_13267,N_11294,N_11278);
nand U13268 (N_13268,N_9827,N_10027);
or U13269 (N_13269,N_11315,N_9515);
nand U13270 (N_13270,N_9439,N_11341);
nor U13271 (N_13271,N_9158,N_11217);
nand U13272 (N_13272,N_11608,N_10224);
nor U13273 (N_13273,N_9613,N_11916);
or U13274 (N_13274,N_11155,N_9923);
and U13275 (N_13275,N_11103,N_11102);
nand U13276 (N_13276,N_10341,N_10593);
and U13277 (N_13277,N_11693,N_10273);
nor U13278 (N_13278,N_9220,N_11994);
nor U13279 (N_13279,N_10315,N_11639);
or U13280 (N_13280,N_10336,N_10663);
or U13281 (N_13281,N_11024,N_10223);
and U13282 (N_13282,N_11712,N_9127);
nor U13283 (N_13283,N_10531,N_11773);
and U13284 (N_13284,N_9457,N_9773);
nand U13285 (N_13285,N_11240,N_9821);
and U13286 (N_13286,N_9416,N_10918);
nand U13287 (N_13287,N_11539,N_11752);
nand U13288 (N_13288,N_9577,N_10678);
nand U13289 (N_13289,N_9957,N_10046);
nand U13290 (N_13290,N_10287,N_10271);
nand U13291 (N_13291,N_10803,N_9938);
nor U13292 (N_13292,N_9464,N_10718);
or U13293 (N_13293,N_9508,N_11461);
and U13294 (N_13294,N_11649,N_11269);
nor U13295 (N_13295,N_11322,N_11776);
and U13296 (N_13296,N_10770,N_10411);
nand U13297 (N_13297,N_9238,N_9967);
nor U13298 (N_13298,N_9490,N_11878);
nor U13299 (N_13299,N_11668,N_9112);
nand U13300 (N_13300,N_10731,N_11585);
nand U13301 (N_13301,N_11045,N_10012);
nand U13302 (N_13302,N_11685,N_9468);
nor U13303 (N_13303,N_10872,N_9583);
nor U13304 (N_13304,N_10665,N_9407);
or U13305 (N_13305,N_11932,N_9844);
nor U13306 (N_13306,N_9792,N_11411);
nor U13307 (N_13307,N_10453,N_10454);
nor U13308 (N_13308,N_10874,N_10324);
nand U13309 (N_13309,N_9288,N_10547);
nor U13310 (N_13310,N_9903,N_11483);
nor U13311 (N_13311,N_9131,N_11640);
or U13312 (N_13312,N_9641,N_9190);
and U13313 (N_13313,N_10188,N_9168);
nor U13314 (N_13314,N_11095,N_9977);
or U13315 (N_13315,N_9140,N_10335);
nor U13316 (N_13316,N_10947,N_11865);
or U13317 (N_13317,N_10331,N_11439);
and U13318 (N_13318,N_10722,N_9318);
and U13319 (N_13319,N_11638,N_9055);
nand U13320 (N_13320,N_9438,N_9814);
nor U13321 (N_13321,N_11679,N_10066);
nor U13322 (N_13322,N_10278,N_11714);
nand U13323 (N_13323,N_11683,N_11137);
and U13324 (N_13324,N_9524,N_11675);
and U13325 (N_13325,N_9287,N_11142);
nor U13326 (N_13326,N_9785,N_9068);
nand U13327 (N_13327,N_9064,N_11260);
or U13328 (N_13328,N_10775,N_11708);
nor U13329 (N_13329,N_9011,N_9584);
nor U13330 (N_13330,N_10350,N_9005);
nand U13331 (N_13331,N_10073,N_11286);
nor U13332 (N_13332,N_9346,N_11100);
nand U13333 (N_13333,N_10473,N_10438);
or U13334 (N_13334,N_9831,N_9432);
nor U13335 (N_13335,N_11595,N_10842);
or U13336 (N_13336,N_10761,N_9592);
or U13337 (N_13337,N_9566,N_11089);
nor U13338 (N_13338,N_11242,N_9410);
nor U13339 (N_13339,N_11213,N_11631);
or U13340 (N_13340,N_9211,N_11976);
nand U13341 (N_13341,N_10289,N_11356);
nand U13342 (N_13342,N_10024,N_11057);
nor U13343 (N_13343,N_10029,N_10912);
and U13344 (N_13344,N_11547,N_11046);
or U13345 (N_13345,N_11819,N_10727);
nor U13346 (N_13346,N_9656,N_9225);
nor U13347 (N_13347,N_9698,N_11111);
or U13348 (N_13348,N_10491,N_9708);
or U13349 (N_13349,N_10578,N_11775);
or U13350 (N_13350,N_10119,N_9398);
nand U13351 (N_13351,N_11555,N_10902);
or U13352 (N_13352,N_11381,N_10848);
and U13353 (N_13353,N_11072,N_9402);
nor U13354 (N_13354,N_10835,N_9540);
or U13355 (N_13355,N_10456,N_9928);
and U13356 (N_13356,N_11915,N_9229);
nand U13357 (N_13357,N_10247,N_11748);
or U13358 (N_13358,N_11148,N_9395);
or U13359 (N_13359,N_11884,N_9647);
nor U13360 (N_13360,N_10667,N_11572);
or U13361 (N_13361,N_11809,N_9580);
nor U13362 (N_13362,N_9489,N_9606);
or U13363 (N_13363,N_9343,N_10534);
nand U13364 (N_13364,N_9570,N_9259);
nor U13365 (N_13365,N_9480,N_9654);
or U13366 (N_13366,N_9022,N_11187);
nand U13367 (N_13367,N_11330,N_10185);
nand U13368 (N_13368,N_9885,N_10654);
and U13369 (N_13369,N_9558,N_10579);
or U13370 (N_13370,N_9344,N_9949);
or U13371 (N_13371,N_11071,N_10921);
nor U13372 (N_13372,N_9971,N_9601);
nor U13373 (N_13373,N_10374,N_10236);
xnor U13374 (N_13374,N_10696,N_9837);
nor U13375 (N_13375,N_11101,N_9436);
or U13376 (N_13376,N_10242,N_10176);
and U13377 (N_13377,N_9191,N_10932);
or U13378 (N_13378,N_10642,N_9074);
and U13379 (N_13379,N_9862,N_10500);
nand U13380 (N_13380,N_9502,N_9629);
and U13381 (N_13381,N_10648,N_10550);
and U13382 (N_13382,N_11185,N_11741);
or U13383 (N_13383,N_9120,N_10074);
and U13384 (N_13384,N_11664,N_10595);
nor U13385 (N_13385,N_11713,N_11373);
or U13386 (N_13386,N_11836,N_9615);
or U13387 (N_13387,N_9325,N_9588);
nand U13388 (N_13388,N_10992,N_10530);
nand U13389 (N_13389,N_10758,N_10843);
nor U13390 (N_13390,N_10042,N_10465);
and U13391 (N_13391,N_10800,N_9806);
and U13392 (N_13392,N_9178,N_10589);
or U13393 (N_13393,N_10121,N_11671);
or U13394 (N_13394,N_10125,N_9379);
nor U13395 (N_13395,N_10339,N_11036);
and U13396 (N_13396,N_10123,N_10145);
nor U13397 (N_13397,N_9252,N_10040);
xnor U13398 (N_13398,N_10613,N_11678);
nor U13399 (N_13399,N_10548,N_11164);
nor U13400 (N_13400,N_9144,N_9921);
and U13401 (N_13401,N_11246,N_9646);
nand U13402 (N_13402,N_10576,N_11233);
or U13403 (N_13403,N_11243,N_11487);
and U13404 (N_13404,N_11084,N_9107);
and U13405 (N_13405,N_10882,N_10839);
nor U13406 (N_13406,N_9813,N_11597);
nor U13407 (N_13407,N_9868,N_9103);
nand U13408 (N_13408,N_9258,N_9589);
nand U13409 (N_13409,N_10325,N_10859);
nor U13410 (N_13410,N_10142,N_11283);
nand U13411 (N_13411,N_9002,N_10625);
and U13412 (N_13412,N_10075,N_11871);
nor U13413 (N_13413,N_10849,N_10159);
nand U13414 (N_13414,N_9241,N_9117);
nand U13415 (N_13415,N_9866,N_9295);
nor U13416 (N_13416,N_10047,N_10884);
and U13417 (N_13417,N_9918,N_9972);
xnor U13418 (N_13418,N_11697,N_9278);
and U13419 (N_13419,N_11346,N_9452);
and U13420 (N_13420,N_10906,N_10375);
and U13421 (N_13421,N_10853,N_11464);
nand U13422 (N_13422,N_11493,N_10691);
or U13423 (N_13423,N_11308,N_10524);
and U13424 (N_13424,N_10353,N_9876);
or U13425 (N_13425,N_9023,N_10426);
and U13426 (N_13426,N_9782,N_10585);
or U13427 (N_13427,N_10334,N_10623);
nand U13428 (N_13428,N_10873,N_9330);
xor U13429 (N_13429,N_11215,N_9041);
or U13430 (N_13430,N_9832,N_10255);
nor U13431 (N_13431,N_9643,N_11436);
and U13432 (N_13432,N_10735,N_9980);
nand U13433 (N_13433,N_11810,N_11705);
or U13434 (N_13434,N_10673,N_11823);
nor U13435 (N_13435,N_10361,N_11406);
nor U13436 (N_13436,N_11670,N_11717);
nor U13437 (N_13437,N_9262,N_11196);
and U13438 (N_13438,N_9979,N_10693);
or U13439 (N_13439,N_10054,N_11231);
nand U13440 (N_13440,N_11469,N_11272);
nand U13441 (N_13441,N_10052,N_11786);
nand U13442 (N_13442,N_11086,N_11831);
nor U13443 (N_13443,N_9066,N_11364);
and U13444 (N_13444,N_9512,N_9683);
nand U13445 (N_13445,N_9699,N_10164);
nand U13446 (N_13446,N_11235,N_11834);
nor U13447 (N_13447,N_10354,N_10264);
nor U13448 (N_13448,N_11870,N_10490);
or U13449 (N_13449,N_10886,N_11305);
or U13450 (N_13450,N_10089,N_11942);
nor U13451 (N_13451,N_11949,N_10127);
or U13452 (N_13452,N_11822,N_10826);
nand U13453 (N_13453,N_9852,N_10031);
nand U13454 (N_13454,N_9774,N_10019);
nor U13455 (N_13455,N_9955,N_10288);
or U13456 (N_13456,N_11458,N_10410);
nand U13457 (N_13457,N_10893,N_9505);
nor U13458 (N_13458,N_10813,N_10858);
nor U13459 (N_13459,N_9766,N_10686);
nand U13460 (N_13460,N_11335,N_10144);
or U13461 (N_13461,N_9075,N_10580);
xor U13462 (N_13462,N_11578,N_9506);
nor U13463 (N_13463,N_11626,N_11427);
or U13464 (N_13464,N_9405,N_9172);
or U13465 (N_13465,N_9454,N_9369);
nand U13466 (N_13466,N_11013,N_9247);
nor U13467 (N_13467,N_9845,N_11442);
nor U13468 (N_13468,N_10383,N_9167);
and U13469 (N_13469,N_9690,N_9293);
and U13470 (N_13470,N_10258,N_10462);
nor U13471 (N_13471,N_10798,N_11456);
or U13472 (N_13472,N_11782,N_11601);
nor U13473 (N_13473,N_11125,N_10393);
and U13474 (N_13474,N_10474,N_10650);
or U13475 (N_13475,N_9455,N_10618);
and U13476 (N_13476,N_10675,N_10519);
nor U13477 (N_13477,N_9283,N_10062);
nor U13478 (N_13478,N_10662,N_10016);
nand U13479 (N_13479,N_10180,N_9473);
nand U13480 (N_13480,N_10114,N_9419);
and U13481 (N_13481,N_10600,N_9496);
nand U13482 (N_13482,N_11962,N_11023);
nand U13483 (N_13483,N_9475,N_10556);
xnor U13484 (N_13484,N_11178,N_10552);
nor U13485 (N_13485,N_9291,N_11088);
nor U13486 (N_13486,N_11395,N_9148);
and U13487 (N_13487,N_9973,N_9411);
xnor U13488 (N_13488,N_11995,N_9221);
nor U13489 (N_13489,N_10878,N_11688);
nor U13490 (N_13490,N_10557,N_10986);
nor U13491 (N_13491,N_9249,N_9380);
nor U13492 (N_13492,N_9449,N_11661);
nor U13493 (N_13493,N_9755,N_10050);
nor U13494 (N_13494,N_11958,N_9942);
or U13495 (N_13495,N_9218,N_9807);
or U13496 (N_13496,N_9509,N_11174);
nand U13497 (N_13497,N_10876,N_10540);
nand U13498 (N_13498,N_10894,N_11739);
and U13499 (N_13499,N_10497,N_11392);
and U13500 (N_13500,N_9338,N_9459);
or U13501 (N_13501,N_11607,N_11438);
and U13502 (N_13502,N_10818,N_11147);
and U13503 (N_13503,N_11296,N_10363);
nor U13504 (N_13504,N_11546,N_9994);
nor U13505 (N_13505,N_10277,N_11786);
and U13506 (N_13506,N_9755,N_9510);
nor U13507 (N_13507,N_10061,N_10117);
and U13508 (N_13508,N_10484,N_10640);
xnor U13509 (N_13509,N_10501,N_11949);
or U13510 (N_13510,N_11807,N_10493);
nand U13511 (N_13511,N_10493,N_11970);
or U13512 (N_13512,N_9589,N_10400);
or U13513 (N_13513,N_9561,N_10272);
or U13514 (N_13514,N_9458,N_11246);
or U13515 (N_13515,N_11929,N_10079);
nor U13516 (N_13516,N_11975,N_11465);
or U13517 (N_13517,N_11132,N_9323);
nand U13518 (N_13518,N_9201,N_11360);
and U13519 (N_13519,N_11938,N_9936);
xor U13520 (N_13520,N_11820,N_9794);
nor U13521 (N_13521,N_11144,N_10860);
and U13522 (N_13522,N_10440,N_11988);
or U13523 (N_13523,N_11243,N_11655);
nand U13524 (N_13524,N_10301,N_9041);
nand U13525 (N_13525,N_10131,N_11760);
nor U13526 (N_13526,N_9105,N_9448);
and U13527 (N_13527,N_10921,N_11866);
and U13528 (N_13528,N_9719,N_11026);
and U13529 (N_13529,N_9464,N_9717);
or U13530 (N_13530,N_11897,N_11493);
and U13531 (N_13531,N_9531,N_11023);
or U13532 (N_13532,N_11309,N_9776);
and U13533 (N_13533,N_10652,N_10749);
xnor U13534 (N_13534,N_10036,N_11706);
nor U13535 (N_13535,N_10728,N_10815);
or U13536 (N_13536,N_9542,N_11549);
nand U13537 (N_13537,N_11981,N_11638);
nor U13538 (N_13538,N_10002,N_10844);
nand U13539 (N_13539,N_10029,N_9288);
nor U13540 (N_13540,N_10895,N_11927);
or U13541 (N_13541,N_11709,N_10962);
and U13542 (N_13542,N_10511,N_10569);
nand U13543 (N_13543,N_9677,N_11287);
and U13544 (N_13544,N_11362,N_9484);
and U13545 (N_13545,N_11022,N_9998);
or U13546 (N_13546,N_10639,N_9610);
or U13547 (N_13547,N_9886,N_11383);
or U13548 (N_13548,N_11704,N_11815);
and U13549 (N_13549,N_9296,N_9821);
or U13550 (N_13550,N_11779,N_10806);
or U13551 (N_13551,N_10905,N_10311);
or U13552 (N_13552,N_10840,N_10115);
nor U13553 (N_13553,N_10725,N_9419);
nand U13554 (N_13554,N_10359,N_9239);
nor U13555 (N_13555,N_10054,N_10985);
nor U13556 (N_13556,N_10701,N_11499);
or U13557 (N_13557,N_10789,N_9733);
nand U13558 (N_13558,N_10212,N_11073);
nor U13559 (N_13559,N_11912,N_10250);
and U13560 (N_13560,N_11978,N_11961);
nor U13561 (N_13561,N_11105,N_10434);
and U13562 (N_13562,N_9427,N_11607);
and U13563 (N_13563,N_9450,N_9762);
nor U13564 (N_13564,N_10324,N_10151);
and U13565 (N_13565,N_10831,N_10662);
nand U13566 (N_13566,N_10166,N_10804);
and U13567 (N_13567,N_9353,N_10251);
nor U13568 (N_13568,N_9692,N_11997);
or U13569 (N_13569,N_10531,N_11818);
nor U13570 (N_13570,N_11958,N_9787);
nor U13571 (N_13571,N_9427,N_10733);
nand U13572 (N_13572,N_10984,N_11738);
or U13573 (N_13573,N_11913,N_10713);
nor U13574 (N_13574,N_10397,N_9939);
nand U13575 (N_13575,N_9615,N_9539);
nand U13576 (N_13576,N_10204,N_9010);
or U13577 (N_13577,N_10251,N_10395);
and U13578 (N_13578,N_10996,N_11842);
and U13579 (N_13579,N_11451,N_10476);
nor U13580 (N_13580,N_10122,N_10206);
and U13581 (N_13581,N_10834,N_9422);
nand U13582 (N_13582,N_9665,N_10836);
nor U13583 (N_13583,N_11544,N_9038);
nand U13584 (N_13584,N_9677,N_10690);
and U13585 (N_13585,N_9828,N_11225);
and U13586 (N_13586,N_11992,N_11018);
or U13587 (N_13587,N_9955,N_11197);
and U13588 (N_13588,N_9673,N_9061);
nor U13589 (N_13589,N_9550,N_10908);
or U13590 (N_13590,N_10168,N_9997);
and U13591 (N_13591,N_9286,N_9922);
nand U13592 (N_13592,N_10045,N_11576);
and U13593 (N_13593,N_9284,N_10971);
or U13594 (N_13594,N_9106,N_10359);
or U13595 (N_13595,N_10650,N_9452);
or U13596 (N_13596,N_11131,N_11145);
or U13597 (N_13597,N_10455,N_10807);
or U13598 (N_13598,N_9669,N_9635);
or U13599 (N_13599,N_10148,N_9299);
and U13600 (N_13600,N_9334,N_11893);
or U13601 (N_13601,N_11543,N_9636);
nand U13602 (N_13602,N_10578,N_9711);
nor U13603 (N_13603,N_9863,N_9430);
or U13604 (N_13604,N_11160,N_9945);
and U13605 (N_13605,N_10674,N_9382);
or U13606 (N_13606,N_10560,N_10859);
nand U13607 (N_13607,N_11937,N_10057);
nor U13608 (N_13608,N_10403,N_10946);
nand U13609 (N_13609,N_10051,N_9168);
nor U13610 (N_13610,N_11520,N_10490);
nand U13611 (N_13611,N_11429,N_10116);
or U13612 (N_13612,N_10291,N_11728);
or U13613 (N_13613,N_10230,N_10485);
and U13614 (N_13614,N_9722,N_9768);
and U13615 (N_13615,N_10878,N_11714);
nand U13616 (N_13616,N_10634,N_10461);
and U13617 (N_13617,N_10679,N_9730);
nor U13618 (N_13618,N_9432,N_9374);
or U13619 (N_13619,N_9814,N_9790);
or U13620 (N_13620,N_10800,N_9772);
or U13621 (N_13621,N_9012,N_10475);
nand U13622 (N_13622,N_9424,N_11117);
and U13623 (N_13623,N_10798,N_10439);
nor U13624 (N_13624,N_10296,N_9209);
or U13625 (N_13625,N_10889,N_11802);
and U13626 (N_13626,N_11918,N_10734);
nand U13627 (N_13627,N_9403,N_9584);
or U13628 (N_13628,N_10553,N_9621);
nor U13629 (N_13629,N_11223,N_9624);
nor U13630 (N_13630,N_10158,N_11791);
nand U13631 (N_13631,N_10310,N_9877);
nand U13632 (N_13632,N_10178,N_11927);
nor U13633 (N_13633,N_11471,N_9857);
and U13634 (N_13634,N_9561,N_10621);
nor U13635 (N_13635,N_11198,N_9604);
nor U13636 (N_13636,N_10438,N_11681);
nor U13637 (N_13637,N_11024,N_9994);
nand U13638 (N_13638,N_10725,N_9509);
and U13639 (N_13639,N_10434,N_10964);
and U13640 (N_13640,N_9942,N_11732);
and U13641 (N_13641,N_9182,N_11375);
nor U13642 (N_13642,N_10873,N_10951);
and U13643 (N_13643,N_11377,N_10990);
nor U13644 (N_13644,N_11558,N_9866);
or U13645 (N_13645,N_10860,N_11482);
and U13646 (N_13646,N_9355,N_10513);
or U13647 (N_13647,N_10442,N_9711);
nand U13648 (N_13648,N_9556,N_10000);
or U13649 (N_13649,N_10179,N_9779);
nor U13650 (N_13650,N_11250,N_11458);
nand U13651 (N_13651,N_10335,N_11792);
nand U13652 (N_13652,N_10507,N_9641);
nor U13653 (N_13653,N_9992,N_9573);
and U13654 (N_13654,N_10906,N_11917);
or U13655 (N_13655,N_9437,N_10081);
and U13656 (N_13656,N_11507,N_10836);
nor U13657 (N_13657,N_10149,N_11265);
and U13658 (N_13658,N_9529,N_10436);
or U13659 (N_13659,N_9710,N_10720);
and U13660 (N_13660,N_11165,N_10708);
or U13661 (N_13661,N_10112,N_10782);
and U13662 (N_13662,N_9674,N_9228);
and U13663 (N_13663,N_10947,N_9051);
or U13664 (N_13664,N_11818,N_10084);
nor U13665 (N_13665,N_11243,N_9665);
nor U13666 (N_13666,N_11823,N_9586);
nor U13667 (N_13667,N_11760,N_10818);
or U13668 (N_13668,N_10956,N_9063);
and U13669 (N_13669,N_10895,N_10677);
nor U13670 (N_13670,N_9613,N_11184);
and U13671 (N_13671,N_9478,N_11239);
nor U13672 (N_13672,N_11774,N_11354);
nor U13673 (N_13673,N_11669,N_9605);
and U13674 (N_13674,N_9252,N_10001);
or U13675 (N_13675,N_10632,N_11134);
or U13676 (N_13676,N_10780,N_10005);
or U13677 (N_13677,N_9008,N_9893);
nor U13678 (N_13678,N_9251,N_11197);
or U13679 (N_13679,N_9345,N_10003);
nor U13680 (N_13680,N_9011,N_9459);
and U13681 (N_13681,N_11413,N_11352);
nor U13682 (N_13682,N_9507,N_10462);
nand U13683 (N_13683,N_11368,N_10822);
nor U13684 (N_13684,N_9704,N_11563);
nor U13685 (N_13685,N_9310,N_10805);
nor U13686 (N_13686,N_10520,N_9171);
nand U13687 (N_13687,N_9817,N_11570);
nor U13688 (N_13688,N_9406,N_11310);
or U13689 (N_13689,N_9605,N_11202);
and U13690 (N_13690,N_9138,N_9805);
nand U13691 (N_13691,N_9508,N_11209);
nand U13692 (N_13692,N_9197,N_10206);
or U13693 (N_13693,N_10948,N_9851);
nand U13694 (N_13694,N_9175,N_10907);
or U13695 (N_13695,N_11659,N_11930);
nand U13696 (N_13696,N_9425,N_10039);
and U13697 (N_13697,N_9346,N_9388);
nor U13698 (N_13698,N_10513,N_9891);
nor U13699 (N_13699,N_10063,N_9898);
and U13700 (N_13700,N_11303,N_9577);
nor U13701 (N_13701,N_10538,N_10492);
and U13702 (N_13702,N_11889,N_9092);
nor U13703 (N_13703,N_10117,N_10526);
nor U13704 (N_13704,N_11213,N_9943);
nand U13705 (N_13705,N_10475,N_10512);
nor U13706 (N_13706,N_11523,N_11736);
nand U13707 (N_13707,N_10969,N_11226);
nor U13708 (N_13708,N_10857,N_9610);
nand U13709 (N_13709,N_9089,N_9796);
nor U13710 (N_13710,N_11187,N_10145);
nand U13711 (N_13711,N_9267,N_9522);
or U13712 (N_13712,N_10208,N_11208);
or U13713 (N_13713,N_10605,N_11305);
nand U13714 (N_13714,N_9043,N_10810);
nand U13715 (N_13715,N_11638,N_11444);
or U13716 (N_13716,N_11708,N_10416);
and U13717 (N_13717,N_10177,N_11620);
nand U13718 (N_13718,N_9940,N_9788);
or U13719 (N_13719,N_9499,N_11052);
nor U13720 (N_13720,N_11449,N_9092);
nor U13721 (N_13721,N_9646,N_10658);
nand U13722 (N_13722,N_10420,N_11239);
nor U13723 (N_13723,N_9914,N_11276);
nor U13724 (N_13724,N_11494,N_9747);
and U13725 (N_13725,N_11785,N_11501);
nor U13726 (N_13726,N_10183,N_10205);
or U13727 (N_13727,N_10449,N_9816);
or U13728 (N_13728,N_10668,N_10611);
xnor U13729 (N_13729,N_9139,N_11729);
nand U13730 (N_13730,N_10727,N_9043);
nor U13731 (N_13731,N_9286,N_10672);
or U13732 (N_13732,N_10122,N_9043);
nand U13733 (N_13733,N_10095,N_9143);
or U13734 (N_13734,N_9811,N_9620);
nand U13735 (N_13735,N_11637,N_9330);
nand U13736 (N_13736,N_9015,N_9088);
or U13737 (N_13737,N_11209,N_9451);
or U13738 (N_13738,N_11122,N_11605);
nor U13739 (N_13739,N_11879,N_11158);
nor U13740 (N_13740,N_11260,N_9883);
and U13741 (N_13741,N_11173,N_9262);
nor U13742 (N_13742,N_9346,N_10304);
or U13743 (N_13743,N_10418,N_9791);
and U13744 (N_13744,N_11459,N_9801);
nor U13745 (N_13745,N_11924,N_11267);
nand U13746 (N_13746,N_11052,N_9630);
and U13747 (N_13747,N_10028,N_11692);
or U13748 (N_13748,N_9085,N_10417);
nand U13749 (N_13749,N_11041,N_9138);
nor U13750 (N_13750,N_11663,N_9475);
or U13751 (N_13751,N_10751,N_9378);
or U13752 (N_13752,N_10433,N_9856);
or U13753 (N_13753,N_10796,N_11429);
nor U13754 (N_13754,N_10256,N_10536);
nand U13755 (N_13755,N_10350,N_10512);
or U13756 (N_13756,N_11188,N_10658);
and U13757 (N_13757,N_11079,N_9352);
nor U13758 (N_13758,N_11723,N_11189);
or U13759 (N_13759,N_11570,N_9239);
or U13760 (N_13760,N_9046,N_10200);
nor U13761 (N_13761,N_9663,N_9708);
nand U13762 (N_13762,N_11140,N_10190);
nand U13763 (N_13763,N_9877,N_11808);
nor U13764 (N_13764,N_11906,N_10026);
and U13765 (N_13765,N_9282,N_11606);
and U13766 (N_13766,N_9040,N_9271);
nand U13767 (N_13767,N_10565,N_11262);
and U13768 (N_13768,N_9180,N_11020);
and U13769 (N_13769,N_10696,N_11666);
nand U13770 (N_13770,N_9708,N_10942);
nand U13771 (N_13771,N_10988,N_10821);
and U13772 (N_13772,N_10799,N_10484);
and U13773 (N_13773,N_11497,N_9489);
nand U13774 (N_13774,N_11045,N_11672);
and U13775 (N_13775,N_11484,N_9144);
nand U13776 (N_13776,N_9437,N_9696);
and U13777 (N_13777,N_11909,N_10542);
nor U13778 (N_13778,N_9100,N_11298);
nor U13779 (N_13779,N_10716,N_9140);
nor U13780 (N_13780,N_9979,N_9465);
or U13781 (N_13781,N_9465,N_9681);
nand U13782 (N_13782,N_11462,N_11889);
or U13783 (N_13783,N_10166,N_10198);
nor U13784 (N_13784,N_9088,N_9553);
nand U13785 (N_13785,N_11258,N_11682);
and U13786 (N_13786,N_9114,N_11097);
nand U13787 (N_13787,N_11124,N_9540);
nand U13788 (N_13788,N_11221,N_9265);
or U13789 (N_13789,N_10028,N_10978);
nand U13790 (N_13790,N_11213,N_9501);
and U13791 (N_13791,N_10090,N_11938);
and U13792 (N_13792,N_10783,N_10941);
and U13793 (N_13793,N_11675,N_9672);
nand U13794 (N_13794,N_9016,N_9101);
or U13795 (N_13795,N_9028,N_9545);
and U13796 (N_13796,N_9860,N_10772);
and U13797 (N_13797,N_10724,N_11263);
or U13798 (N_13798,N_10206,N_10819);
or U13799 (N_13799,N_9641,N_9991);
and U13800 (N_13800,N_11715,N_9366);
and U13801 (N_13801,N_9185,N_11345);
or U13802 (N_13802,N_9925,N_9106);
nand U13803 (N_13803,N_10388,N_11184);
nand U13804 (N_13804,N_9111,N_9146);
or U13805 (N_13805,N_9378,N_9619);
nor U13806 (N_13806,N_11014,N_11474);
nand U13807 (N_13807,N_10553,N_10434);
or U13808 (N_13808,N_9140,N_9346);
and U13809 (N_13809,N_9915,N_11128);
or U13810 (N_13810,N_10340,N_11507);
nor U13811 (N_13811,N_10924,N_9420);
and U13812 (N_13812,N_11384,N_11121);
nor U13813 (N_13813,N_10491,N_11263);
nor U13814 (N_13814,N_11248,N_9498);
or U13815 (N_13815,N_11425,N_11693);
and U13816 (N_13816,N_11749,N_9545);
nor U13817 (N_13817,N_9543,N_10584);
nand U13818 (N_13818,N_11222,N_10904);
nor U13819 (N_13819,N_10470,N_10609);
nor U13820 (N_13820,N_10009,N_9807);
xnor U13821 (N_13821,N_9071,N_11631);
and U13822 (N_13822,N_10554,N_11483);
and U13823 (N_13823,N_10566,N_9842);
and U13824 (N_13824,N_11652,N_10833);
nand U13825 (N_13825,N_11594,N_9585);
and U13826 (N_13826,N_9044,N_10733);
and U13827 (N_13827,N_9815,N_11892);
nor U13828 (N_13828,N_10123,N_11704);
xor U13829 (N_13829,N_10474,N_9976);
nand U13830 (N_13830,N_11050,N_11945);
nand U13831 (N_13831,N_11681,N_9179);
nand U13832 (N_13832,N_11794,N_11225);
nor U13833 (N_13833,N_11200,N_11345);
and U13834 (N_13834,N_10235,N_9479);
or U13835 (N_13835,N_9266,N_11532);
nor U13836 (N_13836,N_11564,N_11481);
or U13837 (N_13837,N_10555,N_10260);
nor U13838 (N_13838,N_10636,N_10898);
or U13839 (N_13839,N_9479,N_11954);
nor U13840 (N_13840,N_11468,N_11965);
and U13841 (N_13841,N_10995,N_9775);
nor U13842 (N_13842,N_10347,N_10701);
or U13843 (N_13843,N_9454,N_9449);
nand U13844 (N_13844,N_9674,N_9085);
or U13845 (N_13845,N_11784,N_11682);
nor U13846 (N_13846,N_11991,N_9197);
or U13847 (N_13847,N_9813,N_9050);
or U13848 (N_13848,N_9877,N_10965);
nor U13849 (N_13849,N_10300,N_9805);
nand U13850 (N_13850,N_10664,N_9880);
nor U13851 (N_13851,N_10512,N_10532);
nand U13852 (N_13852,N_9104,N_9576);
nor U13853 (N_13853,N_9612,N_10564);
or U13854 (N_13854,N_10891,N_10069);
and U13855 (N_13855,N_9587,N_11989);
and U13856 (N_13856,N_10055,N_11178);
nand U13857 (N_13857,N_10120,N_9677);
or U13858 (N_13858,N_11022,N_11271);
nand U13859 (N_13859,N_9309,N_11832);
nand U13860 (N_13860,N_10458,N_9634);
or U13861 (N_13861,N_11984,N_9036);
nand U13862 (N_13862,N_9670,N_10607);
or U13863 (N_13863,N_10927,N_9274);
nor U13864 (N_13864,N_10091,N_10614);
nor U13865 (N_13865,N_9558,N_11359);
and U13866 (N_13866,N_10371,N_9693);
and U13867 (N_13867,N_9073,N_11580);
nand U13868 (N_13868,N_11198,N_11855);
and U13869 (N_13869,N_9403,N_10123);
nand U13870 (N_13870,N_10288,N_9718);
or U13871 (N_13871,N_10395,N_10870);
and U13872 (N_13872,N_9859,N_9380);
or U13873 (N_13873,N_10566,N_9419);
or U13874 (N_13874,N_11416,N_10530);
and U13875 (N_13875,N_9221,N_11735);
and U13876 (N_13876,N_9759,N_11933);
and U13877 (N_13877,N_9871,N_9164);
and U13878 (N_13878,N_11989,N_9981);
nand U13879 (N_13879,N_11843,N_10848);
and U13880 (N_13880,N_9305,N_9708);
nor U13881 (N_13881,N_10658,N_11247);
nand U13882 (N_13882,N_10133,N_11040);
or U13883 (N_13883,N_9824,N_10640);
nor U13884 (N_13884,N_11824,N_11332);
and U13885 (N_13885,N_10689,N_10435);
and U13886 (N_13886,N_10471,N_11756);
or U13887 (N_13887,N_11913,N_11133);
and U13888 (N_13888,N_9061,N_10048);
or U13889 (N_13889,N_9142,N_11928);
or U13890 (N_13890,N_10561,N_10815);
or U13891 (N_13891,N_11624,N_10543);
and U13892 (N_13892,N_9727,N_9029);
nand U13893 (N_13893,N_10612,N_10176);
or U13894 (N_13894,N_9675,N_10779);
nand U13895 (N_13895,N_9118,N_11789);
nand U13896 (N_13896,N_11926,N_10916);
nor U13897 (N_13897,N_9968,N_9533);
nand U13898 (N_13898,N_11868,N_10956);
nand U13899 (N_13899,N_11977,N_10551);
nand U13900 (N_13900,N_9657,N_10644);
and U13901 (N_13901,N_9592,N_10064);
nand U13902 (N_13902,N_11899,N_11818);
or U13903 (N_13903,N_10284,N_10209);
and U13904 (N_13904,N_10226,N_9343);
nor U13905 (N_13905,N_11765,N_11800);
nand U13906 (N_13906,N_9243,N_9637);
or U13907 (N_13907,N_11333,N_11227);
or U13908 (N_13908,N_11083,N_10027);
nand U13909 (N_13909,N_10981,N_11065);
xor U13910 (N_13910,N_10179,N_11652);
or U13911 (N_13911,N_11500,N_11739);
nor U13912 (N_13912,N_9361,N_10097);
nand U13913 (N_13913,N_11954,N_11010);
or U13914 (N_13914,N_11301,N_11788);
or U13915 (N_13915,N_9043,N_9331);
nand U13916 (N_13916,N_9678,N_10462);
nor U13917 (N_13917,N_11393,N_11529);
nand U13918 (N_13918,N_11012,N_11987);
nand U13919 (N_13919,N_10698,N_9220);
nor U13920 (N_13920,N_9027,N_9263);
and U13921 (N_13921,N_10707,N_9077);
nand U13922 (N_13922,N_10076,N_9512);
nand U13923 (N_13923,N_9091,N_9075);
or U13924 (N_13924,N_10072,N_11878);
nor U13925 (N_13925,N_11538,N_11039);
and U13926 (N_13926,N_9714,N_10654);
nand U13927 (N_13927,N_10828,N_11860);
and U13928 (N_13928,N_9778,N_11209);
nand U13929 (N_13929,N_9551,N_11889);
and U13930 (N_13930,N_9772,N_10848);
nand U13931 (N_13931,N_9642,N_9031);
nand U13932 (N_13932,N_11233,N_11593);
or U13933 (N_13933,N_11347,N_9051);
or U13934 (N_13934,N_9468,N_11197);
nor U13935 (N_13935,N_10450,N_9177);
or U13936 (N_13936,N_11345,N_11623);
nor U13937 (N_13937,N_9130,N_9176);
and U13938 (N_13938,N_10749,N_10743);
and U13939 (N_13939,N_10855,N_9248);
or U13940 (N_13940,N_11019,N_9796);
and U13941 (N_13941,N_11047,N_11946);
nand U13942 (N_13942,N_10610,N_11374);
and U13943 (N_13943,N_9585,N_9464);
nor U13944 (N_13944,N_9447,N_10779);
or U13945 (N_13945,N_9460,N_10124);
or U13946 (N_13946,N_11185,N_11237);
nor U13947 (N_13947,N_9024,N_10876);
or U13948 (N_13948,N_9112,N_10392);
nor U13949 (N_13949,N_11559,N_10835);
and U13950 (N_13950,N_9390,N_11946);
and U13951 (N_13951,N_10338,N_10334);
or U13952 (N_13952,N_10735,N_11518);
or U13953 (N_13953,N_10984,N_9762);
nor U13954 (N_13954,N_9308,N_10609);
or U13955 (N_13955,N_10993,N_11174);
and U13956 (N_13956,N_11902,N_11288);
nand U13957 (N_13957,N_10347,N_11739);
or U13958 (N_13958,N_9606,N_9771);
nand U13959 (N_13959,N_10800,N_9105);
nand U13960 (N_13960,N_9326,N_11235);
or U13961 (N_13961,N_9969,N_9065);
nor U13962 (N_13962,N_9439,N_9675);
nor U13963 (N_13963,N_10200,N_9876);
nor U13964 (N_13964,N_10033,N_9193);
nor U13965 (N_13965,N_11126,N_11487);
nand U13966 (N_13966,N_11309,N_11928);
or U13967 (N_13967,N_10807,N_9210);
and U13968 (N_13968,N_9561,N_10495);
or U13969 (N_13969,N_11695,N_11316);
nor U13970 (N_13970,N_11864,N_10478);
nand U13971 (N_13971,N_11907,N_9200);
and U13972 (N_13972,N_9802,N_10693);
or U13973 (N_13973,N_9920,N_9321);
or U13974 (N_13974,N_9724,N_10467);
nand U13975 (N_13975,N_11465,N_9228);
nand U13976 (N_13976,N_10133,N_9691);
and U13977 (N_13977,N_10349,N_10739);
or U13978 (N_13978,N_10071,N_10269);
or U13979 (N_13979,N_11653,N_10395);
or U13980 (N_13980,N_11969,N_9969);
or U13981 (N_13981,N_9441,N_10203);
and U13982 (N_13982,N_11483,N_9738);
and U13983 (N_13983,N_10252,N_10409);
nand U13984 (N_13984,N_10637,N_9375);
and U13985 (N_13985,N_10227,N_11725);
nor U13986 (N_13986,N_11640,N_10886);
nand U13987 (N_13987,N_10581,N_9602);
xor U13988 (N_13988,N_9373,N_11914);
and U13989 (N_13989,N_11348,N_11016);
and U13990 (N_13990,N_9326,N_9054);
nand U13991 (N_13991,N_9672,N_11812);
nor U13992 (N_13992,N_11735,N_11407);
nand U13993 (N_13993,N_11245,N_10029);
nor U13994 (N_13994,N_11317,N_9335);
nor U13995 (N_13995,N_9866,N_9436);
nor U13996 (N_13996,N_9949,N_10535);
xnor U13997 (N_13997,N_11266,N_11891);
and U13998 (N_13998,N_11004,N_9289);
or U13999 (N_13999,N_10138,N_10690);
nor U14000 (N_14000,N_11473,N_9529);
nand U14001 (N_14001,N_9451,N_10780);
or U14002 (N_14002,N_11855,N_9997);
nor U14003 (N_14003,N_9164,N_11592);
nor U14004 (N_14004,N_11027,N_9783);
nor U14005 (N_14005,N_11643,N_9507);
and U14006 (N_14006,N_9793,N_9454);
nor U14007 (N_14007,N_11461,N_10884);
nand U14008 (N_14008,N_9777,N_10472);
nor U14009 (N_14009,N_11953,N_11880);
nand U14010 (N_14010,N_10197,N_9229);
nor U14011 (N_14011,N_11300,N_9496);
nand U14012 (N_14012,N_10066,N_11905);
nand U14013 (N_14013,N_10924,N_9365);
nand U14014 (N_14014,N_11438,N_10000);
or U14015 (N_14015,N_9092,N_9638);
or U14016 (N_14016,N_10889,N_11024);
nand U14017 (N_14017,N_10040,N_10743);
nand U14018 (N_14018,N_11165,N_9665);
nor U14019 (N_14019,N_9391,N_11446);
xor U14020 (N_14020,N_11338,N_11536);
or U14021 (N_14021,N_9324,N_9049);
nor U14022 (N_14022,N_9345,N_9233);
nor U14023 (N_14023,N_10804,N_11546);
or U14024 (N_14024,N_11248,N_9579);
and U14025 (N_14025,N_11480,N_10827);
and U14026 (N_14026,N_10112,N_9817);
nor U14027 (N_14027,N_9362,N_10597);
nor U14028 (N_14028,N_11604,N_11102);
and U14029 (N_14029,N_9272,N_9182);
and U14030 (N_14030,N_11293,N_11494);
nand U14031 (N_14031,N_9516,N_10098);
and U14032 (N_14032,N_10835,N_9683);
nand U14033 (N_14033,N_11420,N_11462);
and U14034 (N_14034,N_11295,N_9021);
and U14035 (N_14035,N_9329,N_9837);
xnor U14036 (N_14036,N_10409,N_10934);
and U14037 (N_14037,N_9275,N_9667);
xnor U14038 (N_14038,N_9191,N_9884);
nor U14039 (N_14039,N_11996,N_11272);
nand U14040 (N_14040,N_10239,N_11818);
and U14041 (N_14041,N_10529,N_10974);
nand U14042 (N_14042,N_9196,N_9157);
or U14043 (N_14043,N_11585,N_9972);
nand U14044 (N_14044,N_10833,N_9553);
nor U14045 (N_14045,N_10667,N_9886);
xnor U14046 (N_14046,N_9106,N_9627);
and U14047 (N_14047,N_9499,N_9460);
and U14048 (N_14048,N_9371,N_9785);
nor U14049 (N_14049,N_10075,N_10425);
and U14050 (N_14050,N_9887,N_9096);
or U14051 (N_14051,N_9123,N_11049);
nand U14052 (N_14052,N_9397,N_10645);
or U14053 (N_14053,N_9099,N_11089);
nor U14054 (N_14054,N_10020,N_11289);
and U14055 (N_14055,N_10449,N_10551);
xnor U14056 (N_14056,N_11579,N_11570);
nor U14057 (N_14057,N_9587,N_11225);
nand U14058 (N_14058,N_10589,N_11801);
and U14059 (N_14059,N_11832,N_11596);
nand U14060 (N_14060,N_11459,N_11384);
or U14061 (N_14061,N_9543,N_10931);
nand U14062 (N_14062,N_10927,N_10835);
or U14063 (N_14063,N_11498,N_10903);
nor U14064 (N_14064,N_10624,N_11062);
nor U14065 (N_14065,N_10478,N_10933);
nor U14066 (N_14066,N_10202,N_9302);
and U14067 (N_14067,N_10013,N_9950);
nand U14068 (N_14068,N_9746,N_9732);
nor U14069 (N_14069,N_9253,N_11715);
or U14070 (N_14070,N_11898,N_9644);
nand U14071 (N_14071,N_10032,N_9981);
nand U14072 (N_14072,N_9051,N_9571);
nor U14073 (N_14073,N_10932,N_10643);
nand U14074 (N_14074,N_11412,N_9922);
or U14075 (N_14075,N_11266,N_9097);
nor U14076 (N_14076,N_10604,N_11242);
and U14077 (N_14077,N_10580,N_9548);
and U14078 (N_14078,N_10524,N_11418);
nor U14079 (N_14079,N_11895,N_10321);
and U14080 (N_14080,N_10288,N_11015);
and U14081 (N_14081,N_9199,N_10508);
nor U14082 (N_14082,N_11610,N_10845);
or U14083 (N_14083,N_10795,N_9681);
nand U14084 (N_14084,N_9918,N_11130);
and U14085 (N_14085,N_10820,N_10330);
or U14086 (N_14086,N_11023,N_9535);
nand U14087 (N_14087,N_9570,N_10128);
and U14088 (N_14088,N_11223,N_9910);
nor U14089 (N_14089,N_9461,N_10160);
or U14090 (N_14090,N_11378,N_11475);
nand U14091 (N_14091,N_9462,N_11226);
nand U14092 (N_14092,N_11254,N_9244);
or U14093 (N_14093,N_10384,N_9916);
nor U14094 (N_14094,N_10635,N_10800);
or U14095 (N_14095,N_11171,N_10823);
nand U14096 (N_14096,N_10437,N_11551);
and U14097 (N_14097,N_11221,N_11669);
or U14098 (N_14098,N_11466,N_11153);
and U14099 (N_14099,N_10126,N_11736);
nor U14100 (N_14100,N_9243,N_10888);
and U14101 (N_14101,N_11633,N_9655);
nor U14102 (N_14102,N_11256,N_9281);
nand U14103 (N_14103,N_11231,N_9405);
or U14104 (N_14104,N_9102,N_9423);
nor U14105 (N_14105,N_11172,N_11413);
or U14106 (N_14106,N_11217,N_11999);
or U14107 (N_14107,N_9983,N_9183);
nand U14108 (N_14108,N_11085,N_9216);
nand U14109 (N_14109,N_11975,N_11372);
nand U14110 (N_14110,N_10939,N_10456);
nand U14111 (N_14111,N_10816,N_10101);
nor U14112 (N_14112,N_9669,N_9947);
nor U14113 (N_14113,N_10735,N_11223);
or U14114 (N_14114,N_11425,N_11702);
nand U14115 (N_14115,N_11256,N_11458);
nand U14116 (N_14116,N_11818,N_11343);
nand U14117 (N_14117,N_10654,N_9723);
or U14118 (N_14118,N_10779,N_10418);
nand U14119 (N_14119,N_11405,N_11808);
nand U14120 (N_14120,N_10564,N_11541);
nor U14121 (N_14121,N_9884,N_11854);
nand U14122 (N_14122,N_9510,N_11488);
nand U14123 (N_14123,N_10298,N_11538);
or U14124 (N_14124,N_10441,N_9096);
nand U14125 (N_14125,N_10820,N_9465);
nand U14126 (N_14126,N_9796,N_11716);
and U14127 (N_14127,N_10520,N_11275);
nand U14128 (N_14128,N_11343,N_11693);
or U14129 (N_14129,N_10500,N_9311);
nor U14130 (N_14130,N_9815,N_9418);
and U14131 (N_14131,N_9728,N_10951);
nand U14132 (N_14132,N_10870,N_9146);
nor U14133 (N_14133,N_10835,N_10071);
and U14134 (N_14134,N_10750,N_11308);
nor U14135 (N_14135,N_11809,N_10373);
nor U14136 (N_14136,N_9990,N_9637);
nor U14137 (N_14137,N_11318,N_9423);
xnor U14138 (N_14138,N_11346,N_10354);
and U14139 (N_14139,N_10692,N_10266);
nand U14140 (N_14140,N_10286,N_9788);
and U14141 (N_14141,N_10977,N_10035);
nand U14142 (N_14142,N_10870,N_9582);
xor U14143 (N_14143,N_9335,N_11433);
nor U14144 (N_14144,N_10361,N_9506);
nor U14145 (N_14145,N_10264,N_9165);
nand U14146 (N_14146,N_11121,N_9679);
nand U14147 (N_14147,N_11450,N_11025);
or U14148 (N_14148,N_9448,N_9240);
nand U14149 (N_14149,N_10330,N_11779);
nor U14150 (N_14150,N_11943,N_10280);
nand U14151 (N_14151,N_10654,N_11432);
nor U14152 (N_14152,N_9811,N_11438);
nand U14153 (N_14153,N_10231,N_11821);
or U14154 (N_14154,N_11275,N_9133);
and U14155 (N_14155,N_11489,N_10626);
and U14156 (N_14156,N_11136,N_10256);
and U14157 (N_14157,N_10847,N_11684);
nor U14158 (N_14158,N_10275,N_9252);
nand U14159 (N_14159,N_9767,N_11864);
nand U14160 (N_14160,N_10731,N_9809);
or U14161 (N_14161,N_9067,N_10304);
nand U14162 (N_14162,N_10727,N_11603);
nor U14163 (N_14163,N_11540,N_10992);
or U14164 (N_14164,N_9153,N_10627);
nor U14165 (N_14165,N_11106,N_11633);
nand U14166 (N_14166,N_11573,N_11403);
nor U14167 (N_14167,N_10536,N_11563);
and U14168 (N_14168,N_9513,N_11540);
or U14169 (N_14169,N_10210,N_9215);
and U14170 (N_14170,N_9530,N_11616);
nor U14171 (N_14171,N_11385,N_10558);
or U14172 (N_14172,N_10649,N_10573);
or U14173 (N_14173,N_9611,N_11169);
or U14174 (N_14174,N_9218,N_11213);
nand U14175 (N_14175,N_9043,N_11485);
or U14176 (N_14176,N_10850,N_9422);
nand U14177 (N_14177,N_10966,N_11009);
nand U14178 (N_14178,N_11591,N_10400);
nand U14179 (N_14179,N_10330,N_11459);
or U14180 (N_14180,N_10749,N_9747);
nand U14181 (N_14181,N_11355,N_11622);
and U14182 (N_14182,N_9299,N_9561);
and U14183 (N_14183,N_11883,N_11715);
and U14184 (N_14184,N_10610,N_9163);
or U14185 (N_14185,N_11698,N_11041);
nor U14186 (N_14186,N_9489,N_11707);
nand U14187 (N_14187,N_11615,N_9305);
nor U14188 (N_14188,N_9191,N_10907);
nand U14189 (N_14189,N_10628,N_10050);
and U14190 (N_14190,N_11391,N_11629);
or U14191 (N_14191,N_10500,N_9487);
or U14192 (N_14192,N_10473,N_9363);
and U14193 (N_14193,N_11520,N_10604);
or U14194 (N_14194,N_9363,N_9095);
nor U14195 (N_14195,N_9829,N_10585);
nand U14196 (N_14196,N_10871,N_11414);
nand U14197 (N_14197,N_11948,N_9758);
or U14198 (N_14198,N_11022,N_11868);
nor U14199 (N_14199,N_10897,N_9199);
and U14200 (N_14200,N_11733,N_10287);
or U14201 (N_14201,N_10157,N_10768);
and U14202 (N_14202,N_11560,N_10794);
or U14203 (N_14203,N_11302,N_11929);
or U14204 (N_14204,N_11061,N_10247);
and U14205 (N_14205,N_10116,N_9830);
nand U14206 (N_14206,N_11594,N_11650);
nor U14207 (N_14207,N_10244,N_11289);
and U14208 (N_14208,N_11154,N_11347);
nand U14209 (N_14209,N_10397,N_11404);
nand U14210 (N_14210,N_9199,N_9491);
or U14211 (N_14211,N_11735,N_11420);
nor U14212 (N_14212,N_9458,N_9065);
nand U14213 (N_14213,N_10900,N_10842);
nor U14214 (N_14214,N_11873,N_10099);
nand U14215 (N_14215,N_11195,N_11260);
nor U14216 (N_14216,N_11551,N_9165);
nand U14217 (N_14217,N_11293,N_11158);
nor U14218 (N_14218,N_9170,N_9744);
or U14219 (N_14219,N_11878,N_9582);
and U14220 (N_14220,N_9837,N_11626);
nor U14221 (N_14221,N_11309,N_11207);
or U14222 (N_14222,N_9334,N_9873);
and U14223 (N_14223,N_11827,N_10940);
nand U14224 (N_14224,N_10789,N_11875);
nand U14225 (N_14225,N_11271,N_11386);
and U14226 (N_14226,N_10379,N_11682);
nor U14227 (N_14227,N_11689,N_11784);
nor U14228 (N_14228,N_10046,N_10060);
nand U14229 (N_14229,N_11994,N_9281);
nand U14230 (N_14230,N_11581,N_11348);
or U14231 (N_14231,N_9047,N_10332);
nor U14232 (N_14232,N_11893,N_9386);
or U14233 (N_14233,N_9971,N_9650);
or U14234 (N_14234,N_9732,N_9844);
and U14235 (N_14235,N_10589,N_11399);
and U14236 (N_14236,N_9164,N_11804);
nand U14237 (N_14237,N_11233,N_11087);
nor U14238 (N_14238,N_10313,N_10844);
nand U14239 (N_14239,N_11495,N_10420);
nand U14240 (N_14240,N_11420,N_10205);
nand U14241 (N_14241,N_10611,N_9236);
nor U14242 (N_14242,N_10471,N_9004);
and U14243 (N_14243,N_9153,N_11772);
nor U14244 (N_14244,N_11204,N_9445);
and U14245 (N_14245,N_10014,N_9026);
nor U14246 (N_14246,N_10426,N_9148);
or U14247 (N_14247,N_9484,N_9035);
and U14248 (N_14248,N_10985,N_9114);
and U14249 (N_14249,N_9790,N_10686);
or U14250 (N_14250,N_9031,N_10508);
and U14251 (N_14251,N_11078,N_9795);
nand U14252 (N_14252,N_10428,N_10271);
and U14253 (N_14253,N_10253,N_9100);
or U14254 (N_14254,N_9504,N_10388);
nor U14255 (N_14255,N_10603,N_10041);
nand U14256 (N_14256,N_11563,N_10648);
nor U14257 (N_14257,N_10499,N_11696);
nor U14258 (N_14258,N_9855,N_10405);
nand U14259 (N_14259,N_9197,N_9450);
or U14260 (N_14260,N_11044,N_9490);
or U14261 (N_14261,N_10409,N_9889);
and U14262 (N_14262,N_10397,N_9035);
and U14263 (N_14263,N_9759,N_10622);
and U14264 (N_14264,N_10194,N_9843);
nor U14265 (N_14265,N_10210,N_10495);
or U14266 (N_14266,N_11515,N_11383);
nor U14267 (N_14267,N_10548,N_11064);
or U14268 (N_14268,N_9761,N_9735);
nor U14269 (N_14269,N_10808,N_11252);
and U14270 (N_14270,N_11541,N_11220);
and U14271 (N_14271,N_11333,N_9548);
or U14272 (N_14272,N_9653,N_11689);
nor U14273 (N_14273,N_10445,N_10147);
nand U14274 (N_14274,N_11974,N_10885);
nand U14275 (N_14275,N_11615,N_9795);
nor U14276 (N_14276,N_10086,N_10402);
nor U14277 (N_14277,N_9906,N_11406);
nor U14278 (N_14278,N_10209,N_9429);
nor U14279 (N_14279,N_9935,N_10871);
nor U14280 (N_14280,N_9605,N_11068);
nand U14281 (N_14281,N_9639,N_10973);
xor U14282 (N_14282,N_9093,N_10209);
or U14283 (N_14283,N_11861,N_9527);
nor U14284 (N_14284,N_9459,N_11937);
or U14285 (N_14285,N_10727,N_9259);
nand U14286 (N_14286,N_11986,N_10140);
nand U14287 (N_14287,N_11979,N_10329);
nand U14288 (N_14288,N_9138,N_10009);
and U14289 (N_14289,N_10945,N_9332);
or U14290 (N_14290,N_10925,N_11691);
nand U14291 (N_14291,N_10974,N_9981);
or U14292 (N_14292,N_10396,N_9862);
nand U14293 (N_14293,N_11625,N_10230);
nor U14294 (N_14294,N_10131,N_9775);
and U14295 (N_14295,N_11745,N_11332);
nand U14296 (N_14296,N_10044,N_11449);
and U14297 (N_14297,N_10985,N_9654);
and U14298 (N_14298,N_9960,N_10427);
and U14299 (N_14299,N_9800,N_9940);
and U14300 (N_14300,N_9631,N_10477);
and U14301 (N_14301,N_11675,N_10319);
nor U14302 (N_14302,N_9208,N_9753);
nand U14303 (N_14303,N_11291,N_11582);
nand U14304 (N_14304,N_10500,N_9058);
or U14305 (N_14305,N_10713,N_10202);
nor U14306 (N_14306,N_9424,N_9096);
nand U14307 (N_14307,N_11708,N_11309);
nor U14308 (N_14308,N_9786,N_10224);
and U14309 (N_14309,N_10639,N_9153);
and U14310 (N_14310,N_9613,N_11157);
or U14311 (N_14311,N_9924,N_11509);
or U14312 (N_14312,N_9510,N_11262);
nor U14313 (N_14313,N_9634,N_11548);
or U14314 (N_14314,N_10500,N_9108);
and U14315 (N_14315,N_11040,N_9544);
nand U14316 (N_14316,N_10524,N_9796);
nor U14317 (N_14317,N_9775,N_9951);
nor U14318 (N_14318,N_9697,N_11665);
nand U14319 (N_14319,N_9089,N_11534);
and U14320 (N_14320,N_11861,N_10215);
and U14321 (N_14321,N_10227,N_9906);
and U14322 (N_14322,N_11320,N_11913);
nor U14323 (N_14323,N_10019,N_10383);
nor U14324 (N_14324,N_11590,N_11496);
nand U14325 (N_14325,N_11766,N_9425);
nand U14326 (N_14326,N_10500,N_10604);
nand U14327 (N_14327,N_11615,N_11787);
or U14328 (N_14328,N_10444,N_11372);
or U14329 (N_14329,N_11606,N_9325);
and U14330 (N_14330,N_10660,N_10160);
nand U14331 (N_14331,N_11985,N_11520);
nor U14332 (N_14332,N_9862,N_10231);
or U14333 (N_14333,N_10515,N_10277);
nand U14334 (N_14334,N_9244,N_10545);
nor U14335 (N_14335,N_9907,N_9413);
or U14336 (N_14336,N_9953,N_11663);
nand U14337 (N_14337,N_10611,N_9378);
nor U14338 (N_14338,N_10808,N_11696);
nand U14339 (N_14339,N_9160,N_9710);
nand U14340 (N_14340,N_10598,N_10875);
nor U14341 (N_14341,N_9637,N_11131);
and U14342 (N_14342,N_11101,N_11674);
nor U14343 (N_14343,N_10674,N_9530);
or U14344 (N_14344,N_9366,N_9000);
or U14345 (N_14345,N_9741,N_11160);
nand U14346 (N_14346,N_9624,N_10192);
or U14347 (N_14347,N_9989,N_9909);
or U14348 (N_14348,N_10057,N_11035);
nor U14349 (N_14349,N_9088,N_11696);
nor U14350 (N_14350,N_9226,N_11486);
xor U14351 (N_14351,N_10803,N_10207);
and U14352 (N_14352,N_10974,N_11366);
or U14353 (N_14353,N_10285,N_11075);
nor U14354 (N_14354,N_9476,N_10625);
and U14355 (N_14355,N_11184,N_9399);
nor U14356 (N_14356,N_10673,N_11883);
nand U14357 (N_14357,N_9058,N_10239);
and U14358 (N_14358,N_9603,N_9195);
or U14359 (N_14359,N_10378,N_10505);
or U14360 (N_14360,N_11861,N_11738);
nand U14361 (N_14361,N_10560,N_10162);
nor U14362 (N_14362,N_10125,N_9758);
and U14363 (N_14363,N_9304,N_9819);
nor U14364 (N_14364,N_11790,N_10556);
nand U14365 (N_14365,N_9475,N_9362);
nor U14366 (N_14366,N_11811,N_9985);
and U14367 (N_14367,N_11972,N_10446);
or U14368 (N_14368,N_10940,N_11319);
nor U14369 (N_14369,N_11112,N_10751);
nand U14370 (N_14370,N_11979,N_10192);
and U14371 (N_14371,N_11756,N_11884);
and U14372 (N_14372,N_10156,N_10900);
nand U14373 (N_14373,N_11735,N_9575);
nand U14374 (N_14374,N_9668,N_11341);
and U14375 (N_14375,N_9307,N_11407);
nor U14376 (N_14376,N_11769,N_9747);
and U14377 (N_14377,N_11004,N_10312);
or U14378 (N_14378,N_9966,N_10613);
nor U14379 (N_14379,N_9061,N_11331);
nor U14380 (N_14380,N_11926,N_11129);
nand U14381 (N_14381,N_9686,N_9819);
and U14382 (N_14382,N_11994,N_10717);
or U14383 (N_14383,N_9198,N_9330);
nand U14384 (N_14384,N_11425,N_11203);
nor U14385 (N_14385,N_10724,N_10273);
nor U14386 (N_14386,N_10439,N_11382);
and U14387 (N_14387,N_11687,N_9987);
nor U14388 (N_14388,N_10853,N_9825);
nor U14389 (N_14389,N_10998,N_10452);
nor U14390 (N_14390,N_9004,N_11646);
or U14391 (N_14391,N_10163,N_11890);
nand U14392 (N_14392,N_9486,N_10124);
or U14393 (N_14393,N_11767,N_11004);
nor U14394 (N_14394,N_11553,N_11169);
nand U14395 (N_14395,N_10336,N_10192);
nand U14396 (N_14396,N_10457,N_10467);
nor U14397 (N_14397,N_9731,N_11426);
or U14398 (N_14398,N_9069,N_11367);
and U14399 (N_14399,N_11886,N_10225);
nand U14400 (N_14400,N_10835,N_10983);
and U14401 (N_14401,N_9021,N_10555);
nand U14402 (N_14402,N_10765,N_10317);
nor U14403 (N_14403,N_10380,N_9594);
and U14404 (N_14404,N_11614,N_11147);
and U14405 (N_14405,N_10928,N_9914);
and U14406 (N_14406,N_11458,N_11915);
and U14407 (N_14407,N_10484,N_10457);
and U14408 (N_14408,N_11824,N_9991);
nand U14409 (N_14409,N_10564,N_10307);
nor U14410 (N_14410,N_9578,N_11701);
nor U14411 (N_14411,N_11025,N_11462);
nor U14412 (N_14412,N_11098,N_10884);
and U14413 (N_14413,N_10575,N_10970);
nor U14414 (N_14414,N_11790,N_10086);
nor U14415 (N_14415,N_11903,N_11624);
or U14416 (N_14416,N_11571,N_11530);
nor U14417 (N_14417,N_9999,N_10918);
and U14418 (N_14418,N_11530,N_11127);
and U14419 (N_14419,N_11233,N_9045);
nand U14420 (N_14420,N_10364,N_10305);
nor U14421 (N_14421,N_9385,N_10130);
nor U14422 (N_14422,N_9287,N_9241);
and U14423 (N_14423,N_10955,N_10792);
or U14424 (N_14424,N_9170,N_10490);
nor U14425 (N_14425,N_11288,N_10721);
and U14426 (N_14426,N_11137,N_9358);
or U14427 (N_14427,N_9598,N_10233);
or U14428 (N_14428,N_11354,N_11284);
and U14429 (N_14429,N_11861,N_9908);
and U14430 (N_14430,N_11545,N_9636);
or U14431 (N_14431,N_9082,N_11782);
or U14432 (N_14432,N_9124,N_11884);
or U14433 (N_14433,N_9980,N_9499);
or U14434 (N_14434,N_9339,N_10818);
and U14435 (N_14435,N_9500,N_9707);
or U14436 (N_14436,N_11516,N_11076);
nor U14437 (N_14437,N_11868,N_10460);
and U14438 (N_14438,N_11892,N_9819);
and U14439 (N_14439,N_9179,N_10040);
and U14440 (N_14440,N_9405,N_10066);
or U14441 (N_14441,N_10109,N_10995);
nand U14442 (N_14442,N_10760,N_10862);
nor U14443 (N_14443,N_11279,N_11297);
nand U14444 (N_14444,N_10665,N_10020);
or U14445 (N_14445,N_11338,N_9877);
and U14446 (N_14446,N_10344,N_10107);
nand U14447 (N_14447,N_9659,N_9515);
and U14448 (N_14448,N_11474,N_10967);
and U14449 (N_14449,N_11593,N_11057);
and U14450 (N_14450,N_9181,N_9771);
nor U14451 (N_14451,N_10281,N_9777);
nor U14452 (N_14452,N_10636,N_9312);
or U14453 (N_14453,N_11117,N_10429);
and U14454 (N_14454,N_10004,N_11611);
and U14455 (N_14455,N_10946,N_9458);
nor U14456 (N_14456,N_11688,N_11074);
nand U14457 (N_14457,N_10886,N_9429);
nor U14458 (N_14458,N_9928,N_9058);
nor U14459 (N_14459,N_11116,N_9425);
nor U14460 (N_14460,N_9969,N_9277);
or U14461 (N_14461,N_10047,N_10678);
nor U14462 (N_14462,N_9703,N_11417);
nand U14463 (N_14463,N_11997,N_10721);
nand U14464 (N_14464,N_11941,N_11564);
and U14465 (N_14465,N_10549,N_11966);
nand U14466 (N_14466,N_11256,N_9036);
nand U14467 (N_14467,N_11789,N_11461);
or U14468 (N_14468,N_9719,N_10175);
nand U14469 (N_14469,N_11020,N_11918);
nor U14470 (N_14470,N_10262,N_10858);
and U14471 (N_14471,N_11333,N_11663);
nor U14472 (N_14472,N_11969,N_10759);
or U14473 (N_14473,N_11850,N_10164);
nor U14474 (N_14474,N_10547,N_11730);
or U14475 (N_14475,N_9911,N_11680);
and U14476 (N_14476,N_10642,N_11819);
nor U14477 (N_14477,N_9243,N_10133);
and U14478 (N_14478,N_9619,N_10174);
nand U14479 (N_14479,N_10125,N_11036);
nand U14480 (N_14480,N_9297,N_10043);
nand U14481 (N_14481,N_9589,N_11768);
nor U14482 (N_14482,N_9101,N_11841);
and U14483 (N_14483,N_9900,N_10240);
nor U14484 (N_14484,N_10184,N_10360);
nor U14485 (N_14485,N_10453,N_11349);
and U14486 (N_14486,N_11564,N_9029);
and U14487 (N_14487,N_10481,N_10140);
or U14488 (N_14488,N_10911,N_9651);
or U14489 (N_14489,N_11312,N_11424);
or U14490 (N_14490,N_9827,N_10404);
nand U14491 (N_14491,N_11446,N_11761);
nand U14492 (N_14492,N_10483,N_11517);
nand U14493 (N_14493,N_10273,N_9128);
nor U14494 (N_14494,N_11587,N_9725);
nand U14495 (N_14495,N_11053,N_11144);
or U14496 (N_14496,N_11863,N_9704);
or U14497 (N_14497,N_11746,N_10821);
and U14498 (N_14498,N_9234,N_10045);
nand U14499 (N_14499,N_11475,N_11839);
nand U14500 (N_14500,N_10135,N_9231);
nor U14501 (N_14501,N_10064,N_11896);
nor U14502 (N_14502,N_10683,N_11711);
and U14503 (N_14503,N_9404,N_10916);
or U14504 (N_14504,N_11991,N_10230);
nand U14505 (N_14505,N_9032,N_11119);
or U14506 (N_14506,N_11588,N_9684);
nor U14507 (N_14507,N_10860,N_9345);
nand U14508 (N_14508,N_11369,N_9830);
or U14509 (N_14509,N_10787,N_11589);
or U14510 (N_14510,N_9703,N_10697);
nand U14511 (N_14511,N_9829,N_10258);
and U14512 (N_14512,N_10803,N_11300);
nand U14513 (N_14513,N_10061,N_11936);
nor U14514 (N_14514,N_11478,N_9509);
and U14515 (N_14515,N_9427,N_9486);
and U14516 (N_14516,N_11468,N_11935);
xnor U14517 (N_14517,N_9834,N_9022);
or U14518 (N_14518,N_9022,N_9545);
nor U14519 (N_14519,N_11676,N_11274);
or U14520 (N_14520,N_10825,N_10550);
nor U14521 (N_14521,N_9898,N_11572);
or U14522 (N_14522,N_11091,N_9763);
nor U14523 (N_14523,N_10702,N_9795);
nor U14524 (N_14524,N_11863,N_10425);
and U14525 (N_14525,N_9290,N_11529);
nand U14526 (N_14526,N_10028,N_11634);
nor U14527 (N_14527,N_9470,N_9917);
or U14528 (N_14528,N_9240,N_9493);
or U14529 (N_14529,N_10137,N_10596);
nor U14530 (N_14530,N_10671,N_9062);
and U14531 (N_14531,N_10136,N_9626);
or U14532 (N_14532,N_11331,N_10191);
nand U14533 (N_14533,N_9806,N_11092);
nand U14534 (N_14534,N_9671,N_9838);
and U14535 (N_14535,N_11410,N_9093);
nor U14536 (N_14536,N_11199,N_10208);
or U14537 (N_14537,N_10947,N_10112);
or U14538 (N_14538,N_9790,N_9907);
nor U14539 (N_14539,N_11742,N_10356);
or U14540 (N_14540,N_10134,N_9386);
nand U14541 (N_14541,N_11674,N_10197);
or U14542 (N_14542,N_9503,N_11602);
and U14543 (N_14543,N_9614,N_10563);
nand U14544 (N_14544,N_10758,N_11920);
and U14545 (N_14545,N_11147,N_9548);
and U14546 (N_14546,N_11567,N_10002);
and U14547 (N_14547,N_10733,N_10410);
nand U14548 (N_14548,N_10420,N_11679);
and U14549 (N_14549,N_10493,N_11426);
or U14550 (N_14550,N_9204,N_10656);
and U14551 (N_14551,N_11160,N_10012);
nand U14552 (N_14552,N_11802,N_10753);
or U14553 (N_14553,N_9461,N_9083);
and U14554 (N_14554,N_11238,N_11936);
nand U14555 (N_14555,N_11673,N_10947);
or U14556 (N_14556,N_10354,N_10613);
nand U14557 (N_14557,N_10958,N_11645);
and U14558 (N_14558,N_10407,N_9817);
and U14559 (N_14559,N_11278,N_9612);
or U14560 (N_14560,N_9602,N_9370);
nand U14561 (N_14561,N_9196,N_9573);
nand U14562 (N_14562,N_10928,N_10606);
and U14563 (N_14563,N_9572,N_10057);
nand U14564 (N_14564,N_10664,N_10997);
nand U14565 (N_14565,N_9469,N_11064);
and U14566 (N_14566,N_11045,N_11072);
and U14567 (N_14567,N_10845,N_10998);
nor U14568 (N_14568,N_9992,N_11738);
nand U14569 (N_14569,N_10975,N_11610);
nor U14570 (N_14570,N_10035,N_10020);
or U14571 (N_14571,N_10902,N_9540);
and U14572 (N_14572,N_11938,N_9027);
or U14573 (N_14573,N_11686,N_11717);
nor U14574 (N_14574,N_10446,N_10867);
nor U14575 (N_14575,N_9543,N_9014);
and U14576 (N_14576,N_9058,N_10808);
or U14577 (N_14577,N_10458,N_9141);
nand U14578 (N_14578,N_10337,N_9410);
and U14579 (N_14579,N_10790,N_10609);
nand U14580 (N_14580,N_10787,N_11224);
and U14581 (N_14581,N_10858,N_11059);
and U14582 (N_14582,N_9417,N_9144);
nor U14583 (N_14583,N_10726,N_10764);
nor U14584 (N_14584,N_10890,N_11102);
nand U14585 (N_14585,N_11198,N_10214);
nor U14586 (N_14586,N_10188,N_9055);
nand U14587 (N_14587,N_10406,N_9503);
nor U14588 (N_14588,N_11220,N_11752);
or U14589 (N_14589,N_10164,N_10074);
or U14590 (N_14590,N_11117,N_9280);
or U14591 (N_14591,N_10055,N_9992);
nor U14592 (N_14592,N_10585,N_10235);
nor U14593 (N_14593,N_9711,N_11984);
or U14594 (N_14594,N_9512,N_10962);
or U14595 (N_14595,N_10267,N_9417);
or U14596 (N_14596,N_10233,N_9207);
nand U14597 (N_14597,N_10987,N_9032);
nand U14598 (N_14598,N_11736,N_11827);
and U14599 (N_14599,N_11871,N_11409);
nand U14600 (N_14600,N_11993,N_9297);
or U14601 (N_14601,N_10224,N_9491);
nand U14602 (N_14602,N_9224,N_11626);
and U14603 (N_14603,N_10781,N_10641);
nor U14604 (N_14604,N_9907,N_11649);
nand U14605 (N_14605,N_10975,N_10480);
and U14606 (N_14606,N_11425,N_9142);
nand U14607 (N_14607,N_10657,N_11342);
and U14608 (N_14608,N_9275,N_11991);
nand U14609 (N_14609,N_11075,N_9252);
nand U14610 (N_14610,N_9334,N_10955);
and U14611 (N_14611,N_11178,N_10648);
and U14612 (N_14612,N_9723,N_10661);
and U14613 (N_14613,N_10872,N_11582);
or U14614 (N_14614,N_11015,N_10648);
nand U14615 (N_14615,N_11116,N_9669);
nor U14616 (N_14616,N_10623,N_10085);
and U14617 (N_14617,N_9658,N_11661);
and U14618 (N_14618,N_9864,N_11380);
and U14619 (N_14619,N_10959,N_11724);
nor U14620 (N_14620,N_10574,N_9081);
and U14621 (N_14621,N_9478,N_11126);
nand U14622 (N_14622,N_9625,N_9183);
and U14623 (N_14623,N_11667,N_10204);
or U14624 (N_14624,N_10043,N_11343);
or U14625 (N_14625,N_9944,N_10537);
or U14626 (N_14626,N_11777,N_10390);
nand U14627 (N_14627,N_9611,N_9726);
nor U14628 (N_14628,N_10805,N_11317);
nand U14629 (N_14629,N_11037,N_9195);
nor U14630 (N_14630,N_11957,N_9771);
nand U14631 (N_14631,N_10921,N_11570);
and U14632 (N_14632,N_10924,N_9692);
and U14633 (N_14633,N_9429,N_9129);
nand U14634 (N_14634,N_10398,N_11100);
nand U14635 (N_14635,N_11777,N_11149);
nor U14636 (N_14636,N_10366,N_9496);
or U14637 (N_14637,N_11169,N_10740);
nor U14638 (N_14638,N_10423,N_9226);
nand U14639 (N_14639,N_10540,N_10478);
or U14640 (N_14640,N_9896,N_10756);
and U14641 (N_14641,N_10414,N_10780);
or U14642 (N_14642,N_9512,N_10500);
nor U14643 (N_14643,N_10421,N_9456);
and U14644 (N_14644,N_11615,N_9140);
or U14645 (N_14645,N_9734,N_11343);
nand U14646 (N_14646,N_11747,N_9031);
or U14647 (N_14647,N_10506,N_9858);
nand U14648 (N_14648,N_10992,N_9502);
nand U14649 (N_14649,N_9140,N_10322);
or U14650 (N_14650,N_10437,N_10532);
nor U14651 (N_14651,N_10429,N_9548);
and U14652 (N_14652,N_9978,N_9025);
nand U14653 (N_14653,N_10177,N_9196);
and U14654 (N_14654,N_9223,N_10920);
nand U14655 (N_14655,N_9507,N_10473);
and U14656 (N_14656,N_10488,N_9297);
nand U14657 (N_14657,N_9782,N_10605);
or U14658 (N_14658,N_10554,N_10698);
nor U14659 (N_14659,N_9701,N_10240);
nor U14660 (N_14660,N_11932,N_11413);
or U14661 (N_14661,N_11944,N_11591);
or U14662 (N_14662,N_11186,N_11639);
or U14663 (N_14663,N_9610,N_11777);
nor U14664 (N_14664,N_9903,N_9879);
nand U14665 (N_14665,N_11689,N_9762);
nor U14666 (N_14666,N_11667,N_10091);
and U14667 (N_14667,N_11464,N_10659);
nand U14668 (N_14668,N_9399,N_11630);
nand U14669 (N_14669,N_11030,N_10330);
or U14670 (N_14670,N_9088,N_9222);
and U14671 (N_14671,N_10429,N_9250);
or U14672 (N_14672,N_9474,N_11937);
and U14673 (N_14673,N_9013,N_9215);
and U14674 (N_14674,N_9262,N_10997);
or U14675 (N_14675,N_10147,N_11056);
or U14676 (N_14676,N_11823,N_11925);
or U14677 (N_14677,N_9540,N_11229);
nor U14678 (N_14678,N_10024,N_11226);
nand U14679 (N_14679,N_10762,N_9399);
and U14680 (N_14680,N_10254,N_11764);
and U14681 (N_14681,N_11766,N_10661);
nor U14682 (N_14682,N_10456,N_9509);
and U14683 (N_14683,N_11078,N_10956);
or U14684 (N_14684,N_11873,N_11951);
nor U14685 (N_14685,N_9318,N_10133);
and U14686 (N_14686,N_11334,N_10809);
or U14687 (N_14687,N_11685,N_9427);
and U14688 (N_14688,N_11524,N_9960);
and U14689 (N_14689,N_11995,N_10174);
or U14690 (N_14690,N_11680,N_10874);
nor U14691 (N_14691,N_11924,N_9969);
or U14692 (N_14692,N_9326,N_9004);
nand U14693 (N_14693,N_10600,N_9006);
or U14694 (N_14694,N_11742,N_10970);
nor U14695 (N_14695,N_9916,N_10865);
nor U14696 (N_14696,N_11993,N_10202);
and U14697 (N_14697,N_10374,N_10127);
and U14698 (N_14698,N_9006,N_11159);
nand U14699 (N_14699,N_10233,N_11255);
or U14700 (N_14700,N_10899,N_9461);
and U14701 (N_14701,N_11135,N_9909);
nor U14702 (N_14702,N_9631,N_9201);
or U14703 (N_14703,N_10475,N_10623);
nor U14704 (N_14704,N_11446,N_10140);
and U14705 (N_14705,N_10745,N_11704);
nor U14706 (N_14706,N_11824,N_10712);
and U14707 (N_14707,N_9015,N_9645);
or U14708 (N_14708,N_10857,N_11388);
and U14709 (N_14709,N_11298,N_10190);
nor U14710 (N_14710,N_11175,N_10637);
nand U14711 (N_14711,N_10725,N_10495);
nand U14712 (N_14712,N_10569,N_11259);
nand U14713 (N_14713,N_11255,N_11597);
or U14714 (N_14714,N_9478,N_11322);
nor U14715 (N_14715,N_10705,N_11259);
and U14716 (N_14716,N_11581,N_11980);
nand U14717 (N_14717,N_10275,N_9574);
or U14718 (N_14718,N_9972,N_11025);
or U14719 (N_14719,N_11725,N_11622);
or U14720 (N_14720,N_10383,N_11939);
or U14721 (N_14721,N_9306,N_11049);
nor U14722 (N_14722,N_10171,N_11685);
nor U14723 (N_14723,N_10431,N_10805);
and U14724 (N_14724,N_11146,N_9206);
nor U14725 (N_14725,N_10842,N_9045);
and U14726 (N_14726,N_9143,N_11962);
nor U14727 (N_14727,N_10810,N_10668);
and U14728 (N_14728,N_9879,N_11533);
and U14729 (N_14729,N_11153,N_11989);
nand U14730 (N_14730,N_9190,N_9182);
or U14731 (N_14731,N_10289,N_11494);
or U14732 (N_14732,N_9227,N_9751);
and U14733 (N_14733,N_9857,N_11038);
nor U14734 (N_14734,N_10349,N_10834);
and U14735 (N_14735,N_9046,N_10893);
xnor U14736 (N_14736,N_10586,N_9011);
nand U14737 (N_14737,N_11716,N_10169);
and U14738 (N_14738,N_10285,N_10138);
and U14739 (N_14739,N_10805,N_10950);
or U14740 (N_14740,N_11768,N_11154);
and U14741 (N_14741,N_10431,N_9655);
or U14742 (N_14742,N_11078,N_10896);
nand U14743 (N_14743,N_9253,N_10156);
nor U14744 (N_14744,N_11929,N_9412);
nand U14745 (N_14745,N_10299,N_10147);
and U14746 (N_14746,N_10014,N_11704);
nand U14747 (N_14747,N_9898,N_10430);
nor U14748 (N_14748,N_9879,N_10442);
and U14749 (N_14749,N_10062,N_11858);
nor U14750 (N_14750,N_11745,N_11215);
or U14751 (N_14751,N_11187,N_9005);
and U14752 (N_14752,N_11993,N_11836);
or U14753 (N_14753,N_10173,N_9597);
nor U14754 (N_14754,N_9629,N_10621);
nor U14755 (N_14755,N_10402,N_10644);
or U14756 (N_14756,N_9763,N_11625);
nor U14757 (N_14757,N_10800,N_11273);
nor U14758 (N_14758,N_9143,N_9390);
nor U14759 (N_14759,N_11606,N_10798);
and U14760 (N_14760,N_11474,N_9255);
or U14761 (N_14761,N_11186,N_9891);
nand U14762 (N_14762,N_10064,N_11341);
or U14763 (N_14763,N_10584,N_11887);
and U14764 (N_14764,N_11951,N_10128);
or U14765 (N_14765,N_9075,N_11775);
nor U14766 (N_14766,N_9045,N_10021);
and U14767 (N_14767,N_11481,N_11546);
nand U14768 (N_14768,N_9055,N_10098);
and U14769 (N_14769,N_9648,N_10989);
or U14770 (N_14770,N_10253,N_11522);
nor U14771 (N_14771,N_10132,N_9353);
and U14772 (N_14772,N_10892,N_11217);
nand U14773 (N_14773,N_10427,N_10375);
nor U14774 (N_14774,N_10497,N_10116);
xor U14775 (N_14775,N_9411,N_9466);
or U14776 (N_14776,N_11752,N_9094);
nor U14777 (N_14777,N_10241,N_11078);
nand U14778 (N_14778,N_10190,N_10592);
nand U14779 (N_14779,N_9268,N_10986);
and U14780 (N_14780,N_11390,N_10454);
nand U14781 (N_14781,N_9947,N_10812);
or U14782 (N_14782,N_11740,N_10180);
nor U14783 (N_14783,N_10398,N_10344);
or U14784 (N_14784,N_10466,N_9203);
nor U14785 (N_14785,N_11895,N_11888);
and U14786 (N_14786,N_10537,N_10309);
nand U14787 (N_14787,N_9750,N_11758);
nor U14788 (N_14788,N_10398,N_10636);
nor U14789 (N_14789,N_9101,N_10992);
nand U14790 (N_14790,N_10269,N_10286);
nor U14791 (N_14791,N_11199,N_9463);
nor U14792 (N_14792,N_10765,N_10777);
nor U14793 (N_14793,N_11797,N_11687);
nand U14794 (N_14794,N_11753,N_10765);
nand U14795 (N_14795,N_10937,N_10833);
nand U14796 (N_14796,N_11720,N_10802);
and U14797 (N_14797,N_10014,N_9816);
and U14798 (N_14798,N_11921,N_10310);
nand U14799 (N_14799,N_10960,N_10531);
or U14800 (N_14800,N_10125,N_11032);
or U14801 (N_14801,N_10217,N_11288);
nand U14802 (N_14802,N_10565,N_11978);
or U14803 (N_14803,N_11745,N_9117);
or U14804 (N_14804,N_10834,N_9782);
nand U14805 (N_14805,N_11158,N_10379);
or U14806 (N_14806,N_9164,N_10221);
or U14807 (N_14807,N_10411,N_11555);
nand U14808 (N_14808,N_11658,N_10593);
or U14809 (N_14809,N_9708,N_10050);
and U14810 (N_14810,N_10558,N_11411);
nand U14811 (N_14811,N_11198,N_9311);
and U14812 (N_14812,N_10623,N_9404);
xor U14813 (N_14813,N_11539,N_11260);
nor U14814 (N_14814,N_10103,N_9484);
or U14815 (N_14815,N_10911,N_9024);
nor U14816 (N_14816,N_11690,N_10265);
nor U14817 (N_14817,N_11943,N_9835);
or U14818 (N_14818,N_10572,N_9755);
or U14819 (N_14819,N_11162,N_11826);
nor U14820 (N_14820,N_9253,N_11250);
and U14821 (N_14821,N_9767,N_9375);
nand U14822 (N_14822,N_9019,N_11409);
nor U14823 (N_14823,N_11809,N_10131);
nand U14824 (N_14824,N_9823,N_9117);
nand U14825 (N_14825,N_10597,N_9969);
and U14826 (N_14826,N_10970,N_9129);
and U14827 (N_14827,N_10302,N_11928);
xor U14828 (N_14828,N_9468,N_10743);
nor U14829 (N_14829,N_9506,N_11940);
or U14830 (N_14830,N_11862,N_10224);
nor U14831 (N_14831,N_9179,N_10086);
or U14832 (N_14832,N_11076,N_11799);
or U14833 (N_14833,N_11056,N_9389);
and U14834 (N_14834,N_10369,N_10299);
nand U14835 (N_14835,N_11740,N_9253);
nand U14836 (N_14836,N_11934,N_10139);
or U14837 (N_14837,N_11303,N_9388);
nor U14838 (N_14838,N_10937,N_9869);
nor U14839 (N_14839,N_10000,N_11684);
nand U14840 (N_14840,N_10774,N_11396);
nand U14841 (N_14841,N_11913,N_11278);
nand U14842 (N_14842,N_9058,N_9244);
nor U14843 (N_14843,N_10882,N_10047);
or U14844 (N_14844,N_10767,N_11751);
nor U14845 (N_14845,N_11341,N_9366);
nor U14846 (N_14846,N_10326,N_9316);
nand U14847 (N_14847,N_9727,N_11185);
nand U14848 (N_14848,N_11028,N_11622);
and U14849 (N_14849,N_10939,N_9698);
xor U14850 (N_14850,N_11449,N_10022);
or U14851 (N_14851,N_11610,N_10346);
nand U14852 (N_14852,N_10239,N_11023);
nand U14853 (N_14853,N_11758,N_10541);
and U14854 (N_14854,N_9431,N_11220);
nor U14855 (N_14855,N_9024,N_11927);
or U14856 (N_14856,N_10231,N_9406);
nand U14857 (N_14857,N_11524,N_9646);
nor U14858 (N_14858,N_9771,N_11738);
nand U14859 (N_14859,N_11623,N_11606);
or U14860 (N_14860,N_9947,N_10918);
or U14861 (N_14861,N_10184,N_11081);
nor U14862 (N_14862,N_10492,N_11818);
nand U14863 (N_14863,N_10360,N_11527);
and U14864 (N_14864,N_10812,N_9552);
nor U14865 (N_14865,N_11907,N_11970);
nand U14866 (N_14866,N_10567,N_11903);
nand U14867 (N_14867,N_10902,N_9587);
nor U14868 (N_14868,N_11508,N_10827);
and U14869 (N_14869,N_11883,N_11383);
nand U14870 (N_14870,N_10923,N_10196);
or U14871 (N_14871,N_9161,N_10353);
nand U14872 (N_14872,N_11008,N_11899);
and U14873 (N_14873,N_10802,N_10366);
nand U14874 (N_14874,N_9979,N_11679);
nand U14875 (N_14875,N_10409,N_11481);
and U14876 (N_14876,N_11960,N_9937);
and U14877 (N_14877,N_9949,N_10574);
nor U14878 (N_14878,N_9099,N_9865);
nand U14879 (N_14879,N_10833,N_10331);
nand U14880 (N_14880,N_10447,N_10090);
or U14881 (N_14881,N_9633,N_9302);
or U14882 (N_14882,N_9489,N_10298);
or U14883 (N_14883,N_11993,N_10276);
or U14884 (N_14884,N_9989,N_9628);
and U14885 (N_14885,N_9386,N_11646);
nand U14886 (N_14886,N_10709,N_9822);
nand U14887 (N_14887,N_10291,N_9817);
nand U14888 (N_14888,N_11984,N_10389);
nor U14889 (N_14889,N_11677,N_9855);
or U14890 (N_14890,N_10317,N_11801);
nor U14891 (N_14891,N_10045,N_10410);
or U14892 (N_14892,N_10779,N_11355);
and U14893 (N_14893,N_10298,N_9504);
or U14894 (N_14894,N_11234,N_10930);
nand U14895 (N_14895,N_10863,N_11713);
and U14896 (N_14896,N_9816,N_10740);
or U14897 (N_14897,N_10444,N_11146);
nor U14898 (N_14898,N_9299,N_11752);
or U14899 (N_14899,N_10363,N_9920);
and U14900 (N_14900,N_9039,N_11776);
nand U14901 (N_14901,N_9251,N_9460);
nand U14902 (N_14902,N_11780,N_9613);
nand U14903 (N_14903,N_11606,N_9733);
xnor U14904 (N_14904,N_11196,N_9785);
nor U14905 (N_14905,N_11576,N_9433);
or U14906 (N_14906,N_11887,N_10909);
or U14907 (N_14907,N_11358,N_11668);
nor U14908 (N_14908,N_11619,N_11942);
and U14909 (N_14909,N_9548,N_9990);
nand U14910 (N_14910,N_11727,N_11796);
xnor U14911 (N_14911,N_11259,N_9390);
or U14912 (N_14912,N_10067,N_11739);
and U14913 (N_14913,N_11494,N_9860);
nor U14914 (N_14914,N_9984,N_9156);
nand U14915 (N_14915,N_9467,N_9741);
or U14916 (N_14916,N_9429,N_9750);
nand U14917 (N_14917,N_11381,N_11679);
and U14918 (N_14918,N_10137,N_10015);
nand U14919 (N_14919,N_10048,N_11203);
or U14920 (N_14920,N_9621,N_11348);
and U14921 (N_14921,N_10538,N_10812);
or U14922 (N_14922,N_9580,N_11769);
and U14923 (N_14923,N_10886,N_9353);
or U14924 (N_14924,N_10823,N_10984);
or U14925 (N_14925,N_11993,N_10128);
nor U14926 (N_14926,N_9814,N_9777);
nand U14927 (N_14927,N_9483,N_11283);
or U14928 (N_14928,N_11010,N_11293);
and U14929 (N_14929,N_10216,N_10940);
and U14930 (N_14930,N_11863,N_9003);
nor U14931 (N_14931,N_9510,N_10817);
nor U14932 (N_14932,N_11276,N_10155);
or U14933 (N_14933,N_11931,N_11192);
nor U14934 (N_14934,N_10454,N_10461);
nand U14935 (N_14935,N_11619,N_9027);
nand U14936 (N_14936,N_11790,N_11663);
nand U14937 (N_14937,N_11296,N_9454);
and U14938 (N_14938,N_9119,N_11601);
and U14939 (N_14939,N_9248,N_9030);
xor U14940 (N_14940,N_9837,N_10700);
or U14941 (N_14941,N_11622,N_11196);
nor U14942 (N_14942,N_11902,N_9279);
nor U14943 (N_14943,N_9980,N_11219);
nor U14944 (N_14944,N_9777,N_10321);
nor U14945 (N_14945,N_11033,N_10353);
nor U14946 (N_14946,N_10988,N_11845);
and U14947 (N_14947,N_9525,N_9411);
nor U14948 (N_14948,N_9397,N_11014);
nor U14949 (N_14949,N_11860,N_9957);
nor U14950 (N_14950,N_11293,N_11586);
or U14951 (N_14951,N_11198,N_10608);
or U14952 (N_14952,N_9808,N_10691);
nor U14953 (N_14953,N_11004,N_10151);
nor U14954 (N_14954,N_11423,N_10133);
nand U14955 (N_14955,N_11984,N_10318);
or U14956 (N_14956,N_9108,N_11338);
and U14957 (N_14957,N_10112,N_11964);
and U14958 (N_14958,N_9765,N_9944);
nor U14959 (N_14959,N_10458,N_9546);
and U14960 (N_14960,N_9908,N_11227);
or U14961 (N_14961,N_11533,N_9551);
or U14962 (N_14962,N_11685,N_9330);
nand U14963 (N_14963,N_9356,N_10585);
and U14964 (N_14964,N_10593,N_10150);
or U14965 (N_14965,N_10625,N_9502);
nand U14966 (N_14966,N_11419,N_10020);
nand U14967 (N_14967,N_9730,N_10336);
nor U14968 (N_14968,N_9816,N_10555);
nor U14969 (N_14969,N_9542,N_9788);
nor U14970 (N_14970,N_11115,N_11962);
and U14971 (N_14971,N_9616,N_10046);
nor U14972 (N_14972,N_9445,N_10866);
or U14973 (N_14973,N_11763,N_9695);
and U14974 (N_14974,N_10451,N_9661);
or U14975 (N_14975,N_10120,N_11604);
or U14976 (N_14976,N_10877,N_11197);
and U14977 (N_14977,N_10021,N_9874);
or U14978 (N_14978,N_10214,N_10578);
or U14979 (N_14979,N_11102,N_10639);
nor U14980 (N_14980,N_10833,N_9386);
and U14981 (N_14981,N_10380,N_10365);
nand U14982 (N_14982,N_9398,N_9464);
and U14983 (N_14983,N_10844,N_11075);
nor U14984 (N_14984,N_9937,N_10052);
or U14985 (N_14985,N_10958,N_10528);
nor U14986 (N_14986,N_9642,N_9526);
and U14987 (N_14987,N_11580,N_9476);
nor U14988 (N_14988,N_11336,N_10557);
nand U14989 (N_14989,N_10506,N_11591);
or U14990 (N_14990,N_11944,N_10681);
or U14991 (N_14991,N_11138,N_9067);
nor U14992 (N_14992,N_9216,N_9583);
nor U14993 (N_14993,N_11612,N_10559);
nand U14994 (N_14994,N_9695,N_10336);
or U14995 (N_14995,N_10028,N_11434);
nor U14996 (N_14996,N_9865,N_11589);
and U14997 (N_14997,N_10312,N_10401);
nand U14998 (N_14998,N_9180,N_9512);
and U14999 (N_14999,N_10459,N_9474);
nand UO_0 (O_0,N_13445,N_14385);
or UO_1 (O_1,N_13659,N_14071);
or UO_2 (O_2,N_14397,N_12166);
nand UO_3 (O_3,N_14223,N_13069);
and UO_4 (O_4,N_13023,N_12497);
and UO_5 (O_5,N_12786,N_13720);
nand UO_6 (O_6,N_14208,N_12840);
nand UO_7 (O_7,N_12267,N_13314);
and UO_8 (O_8,N_12665,N_14265);
or UO_9 (O_9,N_12318,N_13722);
and UO_10 (O_10,N_12337,N_13505);
nand UO_11 (O_11,N_14360,N_12382);
and UO_12 (O_12,N_13498,N_12137);
nor UO_13 (O_13,N_13506,N_14312);
and UO_14 (O_14,N_13852,N_14988);
or UO_15 (O_15,N_14139,N_12702);
or UO_16 (O_16,N_12364,N_13988);
nor UO_17 (O_17,N_13904,N_14827);
and UO_18 (O_18,N_14779,N_14732);
and UO_19 (O_19,N_14088,N_13052);
and UO_20 (O_20,N_12269,N_13782);
and UO_21 (O_21,N_12075,N_12353);
and UO_22 (O_22,N_12213,N_14233);
nand UO_23 (O_23,N_13715,N_13593);
nor UO_24 (O_24,N_13510,N_12654);
nand UO_25 (O_25,N_14555,N_13084);
xor UO_26 (O_26,N_13848,N_13316);
or UO_27 (O_27,N_13628,N_13135);
or UO_28 (O_28,N_14703,N_13345);
nor UO_29 (O_29,N_13875,N_14965);
nand UO_30 (O_30,N_13858,N_12719);
nand UO_31 (O_31,N_14632,N_13353);
nor UO_32 (O_32,N_13101,N_14776);
nand UO_33 (O_33,N_14638,N_12707);
or UO_34 (O_34,N_13789,N_13265);
and UO_35 (O_35,N_12495,N_12234);
nor UO_36 (O_36,N_13572,N_14782);
nor UO_37 (O_37,N_14103,N_12192);
nand UO_38 (O_38,N_12329,N_13427);
or UO_39 (O_39,N_14468,N_14963);
or UO_40 (O_40,N_14339,N_13838);
nand UO_41 (O_41,N_13251,N_12303);
and UO_42 (O_42,N_14157,N_12549);
or UO_43 (O_43,N_14852,N_14459);
nand UO_44 (O_44,N_12024,N_13692);
nand UO_45 (O_45,N_14443,N_13480);
nand UO_46 (O_46,N_14004,N_14876);
nor UO_47 (O_47,N_14238,N_12165);
or UO_48 (O_48,N_14277,N_13563);
and UO_49 (O_49,N_14712,N_12806);
nor UO_50 (O_50,N_13965,N_12920);
nand UO_51 (O_51,N_14814,N_12120);
nand UO_52 (O_52,N_13654,N_14102);
nand UO_53 (O_53,N_12961,N_12930);
and UO_54 (O_54,N_13341,N_13677);
and UO_55 (O_55,N_12035,N_12476);
and UO_56 (O_56,N_12051,N_14906);
nand UO_57 (O_57,N_12407,N_12564);
nor UO_58 (O_58,N_12756,N_14597);
nor UO_59 (O_59,N_14544,N_13291);
and UO_60 (O_60,N_12862,N_14493);
nor UO_61 (O_61,N_13079,N_12972);
nor UO_62 (O_62,N_13211,N_14126);
nor UO_63 (O_63,N_13496,N_14993);
and UO_64 (O_64,N_13526,N_14047);
or UO_65 (O_65,N_14474,N_13614);
or UO_66 (O_66,N_14106,N_12133);
or UO_67 (O_67,N_12985,N_14550);
and UO_68 (O_68,N_12945,N_13119);
or UO_69 (O_69,N_14013,N_14887);
or UO_70 (O_70,N_14028,N_12567);
nor UO_71 (O_71,N_12760,N_14200);
or UO_72 (O_72,N_14596,N_13944);
and UO_73 (O_73,N_14051,N_14345);
or UO_74 (O_74,N_12538,N_12134);
or UO_75 (O_75,N_13636,N_12406);
nand UO_76 (O_76,N_13343,N_13707);
and UO_77 (O_77,N_12630,N_14284);
nand UO_78 (O_78,N_12742,N_14000);
nand UO_79 (O_79,N_12206,N_12148);
nor UO_80 (O_80,N_13869,N_13716);
or UO_81 (O_81,N_12129,N_13169);
nor UO_82 (O_82,N_14784,N_13287);
or UO_83 (O_83,N_12127,N_13357);
and UO_84 (O_84,N_12621,N_12219);
nor UO_85 (O_85,N_14214,N_13093);
nand UO_86 (O_86,N_14984,N_12601);
nand UO_87 (O_87,N_14749,N_13954);
and UO_88 (O_88,N_12019,N_14371);
or UO_89 (O_89,N_13958,N_12596);
nand UO_90 (O_90,N_13232,N_12233);
or UO_91 (O_91,N_14029,N_12284);
and UO_92 (O_92,N_14383,N_13723);
nor UO_93 (O_93,N_13840,N_12465);
or UO_94 (O_94,N_14183,N_13532);
nand UO_95 (O_95,N_14772,N_12734);
nand UO_96 (O_96,N_14046,N_12259);
nand UO_97 (O_97,N_13292,N_14883);
or UO_98 (O_98,N_14444,N_13969);
or UO_99 (O_99,N_12777,N_13043);
nor UO_100 (O_100,N_13805,N_13365);
and UO_101 (O_101,N_13772,N_14836);
nor UO_102 (O_102,N_12677,N_13398);
nor UO_103 (O_103,N_12510,N_14871);
nor UO_104 (O_104,N_13786,N_12074);
and UO_105 (O_105,N_14042,N_12241);
or UO_106 (O_106,N_12060,N_14018);
nor UO_107 (O_107,N_14636,N_14558);
nor UO_108 (O_108,N_13679,N_12713);
or UO_109 (O_109,N_12471,N_12688);
or UO_110 (O_110,N_12907,N_12705);
nand UO_111 (O_111,N_12433,N_12584);
and UO_112 (O_112,N_12229,N_12285);
and UO_113 (O_113,N_12451,N_13968);
and UO_114 (O_114,N_14881,N_13906);
nor UO_115 (O_115,N_13459,N_13437);
nand UO_116 (O_116,N_12992,N_14930);
nor UO_117 (O_117,N_14671,N_12845);
nand UO_118 (O_118,N_13305,N_14367);
or UO_119 (O_119,N_14982,N_14378);
or UO_120 (O_120,N_13433,N_12888);
and UO_121 (O_121,N_14389,N_14594);
and UO_122 (O_122,N_14975,N_12748);
and UO_123 (O_123,N_12894,N_14464);
nand UO_124 (O_124,N_13037,N_14972);
and UO_125 (O_125,N_13661,N_13820);
and UO_126 (O_126,N_13829,N_14281);
nor UO_127 (O_127,N_13774,N_12694);
and UO_128 (O_128,N_13957,N_14868);
and UO_129 (O_129,N_13313,N_13465);
nor UO_130 (O_130,N_14395,N_12076);
nand UO_131 (O_131,N_14408,N_14798);
and UO_132 (O_132,N_14897,N_14672);
or UO_133 (O_133,N_12294,N_13222);
nor UO_134 (O_134,N_13367,N_12668);
or UO_135 (O_135,N_14878,N_12373);
or UO_136 (O_136,N_14316,N_14174);
nand UO_137 (O_137,N_12249,N_13229);
or UO_138 (O_138,N_12614,N_14471);
and UO_139 (O_139,N_14918,N_13897);
nand UO_140 (O_140,N_12362,N_12185);
or UO_141 (O_141,N_13718,N_13434);
nor UO_142 (O_142,N_14295,N_14437);
nand UO_143 (O_143,N_12325,N_13430);
xnor UO_144 (O_144,N_13389,N_14329);
nand UO_145 (O_145,N_14832,N_12718);
nand UO_146 (O_146,N_13947,N_13502);
and UO_147 (O_147,N_14677,N_14384);
nand UO_148 (O_148,N_14967,N_14318);
or UO_149 (O_149,N_14762,N_13472);
nand UO_150 (O_150,N_14181,N_13545);
and UO_151 (O_151,N_14510,N_14856);
nor UO_152 (O_152,N_13142,N_12048);
nand UO_153 (O_153,N_13621,N_13562);
and UO_154 (O_154,N_12121,N_12996);
nand UO_155 (O_155,N_12480,N_14716);
nand UO_156 (O_156,N_14870,N_14575);
nor UO_157 (O_157,N_12741,N_13187);
or UO_158 (O_158,N_13531,N_14956);
nand UO_159 (O_159,N_12975,N_14723);
or UO_160 (O_160,N_12319,N_13997);
nand UO_161 (O_161,N_12624,N_14830);
and UO_162 (O_162,N_13773,N_13635);
nor UO_163 (O_163,N_13310,N_13426);
nor UO_164 (O_164,N_14623,N_14450);
nor UO_165 (O_165,N_14645,N_14566);
xor UO_166 (O_166,N_14504,N_12589);
and UO_167 (O_167,N_12757,N_13309);
nand UO_168 (O_168,N_13412,N_12272);
nand UO_169 (O_169,N_12336,N_14076);
xor UO_170 (O_170,N_14118,N_13216);
nor UO_171 (O_171,N_12411,N_12289);
and UO_172 (O_172,N_12556,N_14280);
nand UO_173 (O_173,N_13095,N_13380);
or UO_174 (O_174,N_14552,N_14934);
and UO_175 (O_175,N_14753,N_14251);
nor UO_176 (O_176,N_13181,N_14182);
nand UO_177 (O_177,N_12004,N_14586);
nand UO_178 (O_178,N_13073,N_12735);
nor UO_179 (O_179,N_14922,N_12101);
nand UO_180 (O_180,N_13753,N_13613);
and UO_181 (O_181,N_14700,N_12118);
nor UO_182 (O_182,N_12717,N_12415);
nor UO_183 (O_183,N_12568,N_14678);
nor UO_184 (O_184,N_13001,N_14068);
and UO_185 (O_185,N_14080,N_14439);
nand UO_186 (O_186,N_14415,N_14646);
or UO_187 (O_187,N_12933,N_13642);
and UO_188 (O_188,N_13517,N_13620);
nand UO_189 (O_189,N_13485,N_14452);
nor UO_190 (O_190,N_14040,N_13457);
nor UO_191 (O_191,N_13020,N_14518);
or UO_192 (O_192,N_14971,N_14061);
nor UO_193 (O_193,N_12498,N_12901);
and UO_194 (O_194,N_14795,N_13451);
nand UO_195 (O_195,N_13790,N_14551);
nand UO_196 (O_196,N_13070,N_14660);
or UO_197 (O_197,N_14232,N_14224);
nor UO_198 (O_198,N_14885,N_12546);
nand UO_199 (O_199,N_12256,N_14170);
and UO_200 (O_200,N_12205,N_13118);
and UO_201 (O_201,N_13177,N_14990);
or UO_202 (O_202,N_12924,N_13959);
nand UO_203 (O_203,N_12053,N_14563);
or UO_204 (O_204,N_13974,N_14215);
and UO_205 (O_205,N_13903,N_12248);
nor UO_206 (O_206,N_13901,N_13928);
nand UO_207 (O_207,N_12847,N_12044);
or UO_208 (O_208,N_14941,N_12386);
or UO_209 (O_209,N_13622,N_13623);
nand UO_210 (O_210,N_12291,N_12902);
nand UO_211 (O_211,N_14011,N_14760);
or UO_212 (O_212,N_13193,N_13551);
and UO_213 (O_213,N_14469,N_12349);
or UO_214 (O_214,N_14599,N_12739);
nand UO_215 (O_215,N_13694,N_14433);
nor UO_216 (O_216,N_13166,N_14486);
nor UO_217 (O_217,N_13953,N_13985);
nand UO_218 (O_218,N_12409,N_12089);
and UO_219 (O_219,N_12798,N_12957);
and UO_220 (O_220,N_14565,N_14419);
nor UO_221 (O_221,N_13534,N_13618);
nand UO_222 (O_222,N_13120,N_13911);
or UO_223 (O_223,N_12460,N_12037);
nand UO_224 (O_224,N_12014,N_12785);
or UO_225 (O_225,N_12102,N_12892);
nand UO_226 (O_226,N_13397,N_13317);
nand UO_227 (O_227,N_14012,N_14884);
xnor UO_228 (O_228,N_14403,N_14615);
or UO_229 (O_229,N_12991,N_14557);
nand UO_230 (O_230,N_14966,N_12764);
nor UO_231 (O_231,N_12203,N_13704);
nand UO_232 (O_232,N_13438,N_12028);
nor UO_233 (O_233,N_13784,N_13266);
or UO_234 (O_234,N_14767,N_13049);
and UO_235 (O_235,N_13246,N_14719);
or UO_236 (O_236,N_14304,N_12054);
or UO_237 (O_237,N_13776,N_13569);
nor UO_238 (O_238,N_14263,N_13989);
nor UO_239 (O_239,N_13812,N_12853);
nor UO_240 (O_240,N_14705,N_12091);
nand UO_241 (O_241,N_13197,N_12725);
and UO_242 (O_242,N_13797,N_13910);
nor UO_243 (O_243,N_14788,N_14659);
nand UO_244 (O_244,N_13796,N_14041);
nor UO_245 (O_245,N_14497,N_13148);
nor UO_246 (O_246,N_13515,N_14577);
or UO_247 (O_247,N_12381,N_12968);
or UO_248 (O_248,N_13567,N_14944);
nand UO_249 (O_249,N_13711,N_12855);
or UO_250 (O_250,N_12598,N_12640);
nor UO_251 (O_251,N_12354,N_12058);
nand UO_252 (O_252,N_13799,N_13298);
or UO_253 (O_253,N_13355,N_13421);
or UO_254 (O_254,N_12002,N_14877);
or UO_255 (O_255,N_12009,N_14454);
or UO_256 (O_256,N_13386,N_14016);
and UO_257 (O_257,N_12155,N_12246);
nor UO_258 (O_258,N_14188,N_12854);
and UO_259 (O_259,N_14920,N_13497);
nor UO_260 (O_260,N_12330,N_14356);
nor UO_261 (O_261,N_12056,N_14568);
xnor UO_262 (O_262,N_13979,N_12818);
nand UO_263 (O_263,N_12485,N_12343);
xnor UO_264 (O_264,N_12222,N_13670);
or UO_265 (O_265,N_13547,N_14642);
xor UO_266 (O_266,N_12508,N_14255);
nand UO_267 (O_267,N_14620,N_14205);
and UO_268 (O_268,N_12721,N_12743);
or UO_269 (O_269,N_12999,N_13557);
xnor UO_270 (O_270,N_12979,N_12466);
nand UO_271 (O_271,N_14848,N_14134);
and UO_272 (O_272,N_14905,N_14766);
nor UO_273 (O_273,N_12324,N_14413);
nand UO_274 (O_274,N_14485,N_14748);
and UO_275 (O_275,N_14618,N_13383);
nor UO_276 (O_276,N_12196,N_12410);
and UO_277 (O_277,N_12475,N_13596);
nand UO_278 (O_278,N_12365,N_12951);
or UO_279 (O_279,N_13468,N_12569);
nand UO_280 (O_280,N_12681,N_12971);
nor UO_281 (O_281,N_12852,N_12963);
or UO_282 (O_282,N_12450,N_13334);
nor UO_283 (O_283,N_14372,N_12690);
or UO_284 (O_284,N_12808,N_13484);
and UO_285 (O_285,N_13111,N_14527);
nor UO_286 (O_286,N_14229,N_14128);
and UO_287 (O_287,N_13295,N_12701);
and UO_288 (O_288,N_12011,N_14349);
and UO_289 (O_289,N_12426,N_13164);
nor UO_290 (O_290,N_13764,N_13059);
nand UO_291 (O_291,N_12385,N_13931);
or UO_292 (O_292,N_12886,N_14697);
nor UO_293 (O_293,N_14501,N_13132);
or UO_294 (O_294,N_14838,N_13755);
and UO_295 (O_295,N_14608,N_13205);
nand UO_296 (O_296,N_13420,N_12472);
nor UO_297 (O_297,N_14479,N_14178);
or UO_298 (O_298,N_14010,N_12268);
or UO_299 (O_299,N_14526,N_12882);
or UO_300 (O_300,N_12714,N_13208);
nand UO_301 (O_301,N_13739,N_13999);
nand UO_302 (O_302,N_12526,N_14352);
nor UO_303 (O_303,N_12428,N_12116);
and UO_304 (O_304,N_13004,N_12006);
nor UO_305 (O_305,N_12750,N_12063);
nor UO_306 (O_306,N_12417,N_14421);
or UO_307 (O_307,N_14744,N_12533);
nor UO_308 (O_308,N_13824,N_13323);
and UO_309 (O_309,N_13582,N_14017);
and UO_310 (O_310,N_13743,N_13051);
and UO_311 (O_311,N_12611,N_14512);
nor UO_312 (O_312,N_14804,N_12391);
or UO_313 (O_313,N_12594,N_14507);
nor UO_314 (O_314,N_14136,N_14588);
nor UO_315 (O_315,N_14542,N_14974);
nor UO_316 (O_316,N_12919,N_12858);
nand UO_317 (O_317,N_13807,N_13105);
nor UO_318 (O_318,N_14726,N_12224);
nor UO_319 (O_319,N_14092,N_12610);
nand UO_320 (O_320,N_12293,N_14931);
or UO_321 (O_321,N_14015,N_13311);
or UO_322 (O_322,N_14926,N_14811);
nand UO_323 (O_323,N_14082,N_12987);
and UO_324 (O_324,N_13814,N_12142);
nor UO_325 (O_325,N_14923,N_13778);
nor UO_326 (O_326,N_13519,N_14258);
or UO_327 (O_327,N_14770,N_14708);
and UO_328 (O_328,N_14430,N_13149);
nor UO_329 (O_329,N_14725,N_12299);
or UO_330 (O_330,N_12307,N_13245);
and UO_331 (O_331,N_14520,N_13733);
or UO_332 (O_332,N_13100,N_12017);
nand UO_333 (O_333,N_12592,N_14969);
and UO_334 (O_334,N_12140,N_12516);
nand UO_335 (O_335,N_14573,N_14275);
and UO_336 (O_336,N_12023,N_12470);
nand UO_337 (O_337,N_12615,N_14562);
nor UO_338 (O_338,N_12228,N_13206);
nor UO_339 (O_339,N_14289,N_13214);
or UO_340 (O_340,N_14976,N_13153);
nand UO_341 (O_341,N_12295,N_14517);
and UO_342 (O_342,N_13372,N_14406);
or UO_343 (O_343,N_13634,N_12966);
or UO_344 (O_344,N_13631,N_13709);
and UO_345 (O_345,N_14494,N_13746);
or UO_346 (O_346,N_12696,N_13455);
or UO_347 (O_347,N_12168,N_13826);
nand UO_348 (O_348,N_12125,N_14824);
or UO_349 (O_349,N_14682,N_13996);
nand UO_350 (O_350,N_14322,N_14955);
or UO_351 (O_351,N_14704,N_12593);
and UO_352 (O_352,N_14394,N_12745);
and UO_353 (O_353,N_13032,N_14211);
nor UO_354 (O_354,N_12207,N_13751);
nor UO_355 (O_355,N_12445,N_13587);
or UO_356 (O_356,N_12368,N_12164);
nand UO_357 (O_357,N_13012,N_13603);
xnor UO_358 (O_358,N_12488,N_12704);
and UO_359 (O_359,N_12220,N_12573);
nor UO_360 (O_360,N_14083,N_13090);
nor UO_361 (O_361,N_14301,N_12988);
nand UO_362 (O_362,N_12575,N_12595);
nor UO_363 (O_363,N_14366,N_12970);
nand UO_364 (O_364,N_14900,N_14822);
or UO_365 (O_365,N_13609,N_14303);
nor UO_366 (O_366,N_13410,N_14655);
nor UO_367 (O_367,N_14609,N_13019);
and UO_368 (O_368,N_14351,N_14968);
and UO_369 (O_369,N_12317,N_14353);
nor UO_370 (O_370,N_14821,N_13611);
nand UO_371 (O_371,N_13008,N_12637);
nand UO_372 (O_372,N_12899,N_13044);
nor UO_373 (O_373,N_13456,N_14579);
or UO_374 (O_374,N_14809,N_14225);
and UO_375 (O_375,N_13393,N_13471);
nand UO_376 (O_376,N_13218,N_12332);
or UO_377 (O_377,N_14359,N_12962);
nand UO_378 (O_378,N_13580,N_14543);
nand UO_379 (O_379,N_13228,N_12603);
nor UO_380 (O_380,N_13320,N_14161);
or UO_381 (O_381,N_12941,N_12715);
nor UO_382 (O_382,N_14325,N_14034);
nor UO_383 (O_383,N_12320,N_14751);
nor UO_384 (O_384,N_14635,N_13136);
nand UO_385 (O_385,N_13712,N_12327);
and UO_386 (O_386,N_13527,N_13225);
and UO_387 (O_387,N_14940,N_13146);
and UO_388 (O_388,N_12523,N_14243);
nand UO_389 (O_389,N_12550,N_12012);
or UO_390 (O_390,N_14833,N_14539);
and UO_391 (O_391,N_14120,N_12350);
nand UO_392 (O_392,N_12642,N_12553);
nor UO_393 (O_393,N_13913,N_13074);
and UO_394 (O_394,N_12298,N_13689);
and UO_395 (O_395,N_13941,N_14368);
nand UO_396 (O_396,N_12109,N_13007);
nor UO_397 (O_397,N_12186,N_14077);
and UO_398 (O_398,N_13554,N_14457);
or UO_399 (O_399,N_12238,N_12374);
and UO_400 (O_400,N_14591,N_13740);
nor UO_401 (O_401,N_14999,N_14624);
nand UO_402 (O_402,N_13573,N_14778);
nor UO_403 (O_403,N_12657,N_13277);
nor UO_404 (O_404,N_14230,N_12995);
nor UO_405 (O_405,N_14484,N_12499);
and UO_406 (O_406,N_14172,N_13737);
nor UO_407 (O_407,N_13354,N_12571);
or UO_408 (O_408,N_13196,N_14310);
or UO_409 (O_409,N_12982,N_13518);
nand UO_410 (O_410,N_13939,N_12181);
or UO_411 (O_411,N_13752,N_14006);
or UO_412 (O_412,N_13972,N_13512);
and UO_413 (O_413,N_12736,N_12096);
nor UO_414 (O_414,N_12939,N_13775);
nand UO_415 (O_415,N_12221,N_14619);
nand UO_416 (O_416,N_13945,N_14515);
or UO_417 (O_417,N_13422,N_13942);
or UO_418 (O_418,N_14180,N_13040);
nand UO_419 (O_419,N_12449,N_12521);
nand UO_420 (O_420,N_14582,N_14741);
or UO_421 (O_421,N_12931,N_12561);
nand UO_422 (O_422,N_12505,N_12340);
nand UO_423 (O_423,N_12956,N_12938);
nand UO_424 (O_424,N_12395,N_14717);
nor UO_425 (O_425,N_12693,N_13442);
nand UO_426 (O_426,N_13483,N_14994);
nor UO_427 (O_427,N_14513,N_12747);
nand UO_428 (O_428,N_12789,N_12986);
and UO_429 (O_429,N_14869,N_12280);
nor UO_430 (O_430,N_13666,N_14585);
and UO_431 (O_431,N_14189,N_13467);
and UO_432 (O_432,N_12240,N_13283);
and UO_433 (O_433,N_13263,N_12829);
or UO_434 (O_434,N_13331,N_12940);
and UO_435 (O_435,N_14052,N_14154);
nor UO_436 (O_436,N_13699,N_14216);
nor UO_437 (O_437,N_13543,N_14595);
nand UO_438 (O_438,N_13564,N_14673);
and UO_439 (O_439,N_13322,N_12699);
and UO_440 (O_440,N_14979,N_12176);
and UO_441 (O_441,N_14613,N_14584);
nor UO_442 (O_442,N_13702,N_12126);
nand UO_443 (O_443,N_12960,N_14733);
nand UO_444 (O_444,N_12998,N_12288);
nand UO_445 (O_445,N_12698,N_14909);
and UO_446 (O_446,N_14724,N_14813);
or UO_447 (O_447,N_14675,N_12586);
or UO_448 (O_448,N_12309,N_13171);
and UO_449 (O_449,N_14683,N_12762);
and UO_450 (O_450,N_13630,N_14657);
nand UO_451 (O_451,N_13038,N_12375);
or UO_452 (O_452,N_13203,N_14589);
and UO_453 (O_453,N_12923,N_14007);
nor UO_454 (O_454,N_14107,N_14122);
nand UO_455 (O_455,N_13750,N_13676);
nand UO_456 (O_456,N_12169,N_13960);
and UO_457 (O_457,N_13473,N_13139);
nand UO_458 (O_458,N_14773,N_12903);
nand UO_459 (O_459,N_12257,N_12787);
and UO_460 (O_460,N_14625,N_12652);
nor UO_461 (O_461,N_13159,N_13185);
nand UO_462 (O_462,N_13065,N_13102);
and UO_463 (O_463,N_12469,N_12345);
nor UO_464 (O_464,N_14451,N_13934);
or UO_465 (O_465,N_13655,N_13030);
or UO_466 (O_466,N_13128,N_14808);
nor UO_467 (O_467,N_13907,N_14110);
and UO_468 (O_468,N_12039,N_14818);
nor UO_469 (O_469,N_12579,N_12083);
nand UO_470 (O_470,N_14872,N_13429);
or UO_471 (O_471,N_12994,N_13385);
or UO_472 (O_472,N_13470,N_14458);
and UO_473 (O_473,N_13542,N_14307);
nor UO_474 (O_474,N_12638,N_14765);
and UO_475 (O_475,N_13035,N_13841);
nor UO_476 (O_476,N_13871,N_13207);
nor UO_477 (O_477,N_12323,N_13652);
or UO_478 (O_478,N_13346,N_13057);
and UO_479 (O_479,N_12837,N_12119);
nand UO_480 (O_480,N_13419,N_13478);
nor UO_481 (O_481,N_13920,N_12467);
and UO_482 (O_482,N_14522,N_12531);
nor UO_483 (O_483,N_12388,N_12195);
and UO_484 (O_484,N_13441,N_12772);
nand UO_485 (O_485,N_12669,N_13358);
or UO_486 (O_486,N_14864,N_13282);
nor UO_487 (O_487,N_12174,N_12007);
or UO_488 (O_488,N_14025,N_13949);
nor UO_489 (O_489,N_13813,N_14849);
and UO_490 (O_490,N_14123,N_14094);
or UO_491 (O_491,N_12749,N_14268);
nand UO_492 (O_492,N_13150,N_13077);
and UO_493 (O_493,N_12380,N_13501);
or UO_494 (O_494,N_13474,N_13765);
or UO_495 (O_495,N_12997,N_13938);
and UO_496 (O_496,N_14490,N_12722);
or UO_497 (O_497,N_12043,N_14875);
or UO_498 (O_498,N_14311,N_12200);
or UO_499 (O_499,N_14722,N_12653);
or UO_500 (O_500,N_14343,N_14100);
and UO_501 (O_501,N_14912,N_13568);
or UO_502 (O_502,N_12636,N_13986);
and UO_503 (O_503,N_13094,N_14924);
nand UO_504 (O_504,N_12904,N_14855);
and UO_505 (O_505,N_12369,N_12834);
nand UO_506 (O_506,N_12447,N_13637);
nor UO_507 (O_507,N_12030,N_12239);
and UO_508 (O_508,N_13791,N_12384);
nor UO_509 (O_509,N_13238,N_14980);
or UO_510 (O_510,N_14226,N_13318);
nand UO_511 (O_511,N_12535,N_14160);
nand UO_512 (O_512,N_13391,N_12444);
nor UO_513 (O_513,N_12077,N_13462);
nor UO_514 (O_514,N_12755,N_12848);
or UO_515 (O_515,N_14294,N_13415);
or UO_516 (O_516,N_12989,N_13589);
nand UO_517 (O_517,N_12439,N_14105);
nor UO_518 (O_518,N_14534,N_13464);
nand UO_519 (O_519,N_12790,N_12159);
nor UO_520 (O_520,N_12860,N_14323);
or UO_521 (O_521,N_12070,N_12131);
or UO_522 (O_522,N_13300,N_12477);
and UO_523 (O_523,N_14005,N_13809);
or UO_524 (O_524,N_14209,N_12231);
or UO_525 (O_525,N_13680,N_12519);
or UO_526 (O_526,N_14684,N_14932);
and UO_527 (O_527,N_14404,N_13847);
and UO_528 (O_528,N_14387,N_13883);
nor UO_529 (O_529,N_13449,N_12607);
nor UO_530 (O_530,N_12171,N_14826);
or UO_531 (O_531,N_13215,N_12128);
and UO_532 (O_532,N_13034,N_14587);
and UO_533 (O_533,N_12390,N_12646);
and UO_534 (O_534,N_14828,N_12738);
nor UO_535 (O_535,N_13632,N_14089);
nor UO_536 (O_536,N_13308,N_13602);
and UO_537 (O_537,N_14482,N_13486);
or UO_538 (O_538,N_14044,N_13581);
and UO_539 (O_539,N_12916,N_12953);
nand UO_540 (O_540,N_13022,N_14401);
nor UO_541 (O_541,N_14531,N_13705);
or UO_542 (O_542,N_13792,N_12286);
or UO_543 (O_543,N_14373,N_14942);
nor UO_544 (O_544,N_13031,N_13304);
nor UO_545 (O_545,N_12292,N_13520);
and UO_546 (O_546,N_14293,N_12032);
or UO_547 (O_547,N_12955,N_12297);
nand UO_548 (O_548,N_13117,N_12360);
nor UO_549 (O_549,N_14097,N_14037);
and UO_550 (O_550,N_14521,N_12013);
nor UO_551 (O_551,N_12424,N_14348);
nand UO_552 (O_552,N_14962,N_13588);
nand UO_553 (O_553,N_14141,N_12328);
nor UO_554 (O_554,N_13717,N_14781);
nor UO_555 (O_555,N_12082,N_14651);
and UO_556 (O_556,N_13366,N_14422);
or UO_557 (O_557,N_14472,N_14880);
nand UO_558 (O_558,N_12874,N_12663);
nor UO_559 (O_559,N_13066,N_13431);
or UO_560 (O_560,N_12394,N_12697);
or UO_561 (O_561,N_12045,N_13072);
and UO_562 (O_562,N_14145,N_13339);
nor UO_563 (O_563,N_12978,N_12691);
and UO_564 (O_564,N_13747,N_13167);
nand UO_565 (O_565,N_14560,N_12588);
and UO_566 (O_566,N_13600,N_12236);
nand UO_567 (O_567,N_13446,N_14896);
and UO_568 (O_568,N_13157,N_14685);
nor UO_569 (O_569,N_14278,N_13761);
or UO_570 (O_570,N_13112,N_12421);
nor UO_571 (O_571,N_14184,N_13605);
nor UO_572 (O_572,N_14393,N_13578);
xnor UO_573 (O_573,N_14545,N_14259);
nor UO_574 (O_574,N_12115,N_14567);
and UO_575 (O_575,N_12838,N_14132);
nor UO_576 (O_576,N_13644,N_14417);
or UO_577 (O_577,N_13818,N_12344);
and UO_578 (O_578,N_14297,N_14541);
and UO_579 (O_579,N_13698,N_13481);
nor UO_580 (O_580,N_13980,N_14863);
and UO_581 (O_581,N_13143,N_14498);
nand UO_582 (O_582,N_13289,N_13244);
and UO_583 (O_583,N_13533,N_12566);
and UO_584 (O_584,N_12878,N_12453);
nand UO_585 (O_585,N_13595,N_14888);
and UO_586 (O_586,N_14927,N_12841);
nand UO_587 (O_587,N_14317,N_14516);
or UO_588 (O_588,N_14424,N_12130);
and UO_589 (O_589,N_12342,N_12509);
and UO_590 (O_590,N_13373,N_12720);
nor UO_591 (O_591,N_14928,N_13884);
xnor UO_592 (O_592,N_14977,N_12026);
nand UO_593 (O_593,N_12676,N_12093);
nand UO_594 (O_594,N_14252,N_14890);
nor UO_595 (O_595,N_13352,N_14279);
nand UO_596 (O_596,N_14369,N_12372);
nand UO_597 (O_597,N_12487,N_13350);
or UO_598 (O_598,N_14747,N_14274);
nor UO_599 (O_599,N_12915,N_12018);
nand UO_600 (O_600,N_13490,N_14027);
and UO_601 (O_601,N_13330,N_13256);
or UO_602 (O_602,N_12396,N_13200);
nand UO_603 (O_603,N_12666,N_13845);
and UO_604 (O_604,N_14266,N_12047);
nor UO_605 (O_605,N_12478,N_12572);
or UO_606 (O_606,N_12791,N_12254);
nand UO_607 (O_607,N_14559,N_13971);
nor UO_608 (O_608,N_13819,N_14202);
or UO_609 (O_609,N_14674,N_14287);
and UO_610 (O_610,N_14561,N_14381);
or UO_611 (O_611,N_14283,N_12208);
or UO_612 (O_612,N_14391,N_13671);
or UO_613 (O_613,N_12574,N_13141);
and UO_614 (O_614,N_13900,N_13932);
or UO_615 (O_615,N_14961,N_12435);
or UO_616 (O_616,N_12275,N_13912);
nor UO_617 (O_617,N_14173,N_12484);
or UO_618 (O_618,N_13180,N_13681);
nor UO_619 (O_619,N_13536,N_13836);
or UO_620 (O_620,N_12823,N_13016);
or UO_621 (O_621,N_14981,N_14665);
nor UO_622 (O_622,N_14769,N_14340);
or UO_623 (O_623,N_14739,N_13210);
or UO_624 (O_624,N_14639,N_14300);
nor UO_625 (O_625,N_14039,N_13125);
nor UO_626 (O_626,N_13230,N_13168);
nor UO_627 (O_627,N_14874,N_14954);
or UO_628 (O_628,N_13538,N_12245);
and UO_629 (O_629,N_14109,N_13163);
nor UO_630 (O_630,N_13458,N_12212);
nand UO_631 (O_631,N_12483,N_12529);
and UO_632 (O_632,N_14669,N_12746);
or UO_633 (O_633,N_14187,N_14461);
nand UO_634 (O_634,N_12105,N_14143);
nor UO_635 (O_635,N_12819,N_12178);
or UO_636 (O_636,N_13650,N_14862);
or UO_637 (O_637,N_13048,N_12976);
and UO_638 (O_638,N_13264,N_13586);
nand UO_639 (O_639,N_14299,N_13929);
nor UO_640 (O_640,N_12943,N_14218);
nor UO_641 (O_641,N_13788,N_13290);
and UO_642 (O_642,N_13565,N_12106);
and UO_643 (O_643,N_12527,N_12189);
nor UO_644 (O_644,N_13662,N_12990);
nand UO_645 (O_645,N_13639,N_13624);
nor UO_646 (O_646,N_13378,N_13610);
nor UO_647 (O_647,N_12909,N_12656);
nor UO_648 (O_648,N_12402,N_14432);
and UO_649 (O_649,N_12664,N_14911);
and UO_650 (O_650,N_14400,N_13891);
or UO_651 (O_651,N_14341,N_12709);
nand UO_652 (O_652,N_13835,N_12766);
or UO_653 (O_653,N_14668,N_12507);
and UO_654 (O_654,N_14652,N_12815);
nand UO_655 (O_655,N_13424,N_12455);
and UO_656 (O_656,N_13983,N_13759);
nand UO_657 (O_657,N_12883,N_14072);
nor UO_658 (O_658,N_14714,N_14576);
and UO_659 (O_659,N_13905,N_14194);
and UO_660 (O_660,N_13013,N_12072);
or UO_661 (O_661,N_13085,N_14819);
or UO_662 (O_662,N_12264,N_14057);
nor UO_663 (O_663,N_12528,N_12773);
nor UO_664 (O_664,N_14812,N_14666);
nand UO_665 (O_665,N_13503,N_13665);
nand UO_666 (O_666,N_12461,N_13219);
nor UO_667 (O_667,N_12504,N_14946);
or UO_668 (O_668,N_13147,N_13769);
nand UO_669 (O_669,N_12025,N_14785);
or UO_670 (O_670,N_13925,N_13529);
nor UO_671 (O_671,N_14150,N_13626);
nor UO_672 (O_672,N_14203,N_14488);
nor UO_673 (O_673,N_13050,N_14321);
and UO_674 (O_674,N_12587,N_13110);
nand UO_675 (O_675,N_13227,N_13492);
nand UO_676 (O_676,N_12333,N_13302);
nor UO_677 (O_677,N_13880,N_13260);
or UO_678 (O_678,N_14514,N_12684);
or UO_679 (O_679,N_13444,N_13212);
or UO_680 (O_680,N_12005,N_14771);
nand UO_681 (O_681,N_12261,N_14315);
and UO_682 (O_682,N_13815,N_13499);
and UO_683 (O_683,N_12474,N_14950);
nand UO_684 (O_684,N_12767,N_14462);
nor UO_685 (O_685,N_14556,N_14073);
nand UO_686 (O_686,N_14399,N_14392);
or UO_687 (O_687,N_12172,N_14442);
and UO_688 (O_688,N_14217,N_13922);
or UO_689 (O_689,N_12708,N_13673);
or UO_690 (O_690,N_13594,N_14163);
nor UO_691 (O_691,N_14374,N_13332);
or UO_692 (O_692,N_13493,N_13384);
or UO_693 (O_693,N_13109,N_12993);
nand UO_694 (O_694,N_14460,N_14879);
or UO_695 (O_695,N_13097,N_12080);
nand UO_696 (O_696,N_12754,N_12627);
nor UO_697 (O_697,N_14346,N_14569);
or UO_698 (O_698,N_14538,N_12558);
nor UO_699 (O_699,N_12167,N_12367);
and UO_700 (O_700,N_13017,N_13521);
nor UO_701 (O_701,N_13627,N_12255);
or UO_702 (O_702,N_12310,N_14113);
and UO_703 (O_703,N_13686,N_12670);
nand UO_704 (O_704,N_12434,N_12225);
nand UO_705 (O_705,N_12230,N_13239);
and UO_706 (O_706,N_13406,N_12440);
or UO_707 (O_707,N_12918,N_13982);
nand UO_708 (O_708,N_12250,N_14446);
nand UO_709 (O_709,N_12896,N_12263);
and UO_710 (O_710,N_13337,N_13114);
or UO_711 (O_711,N_14519,N_12795);
nor UO_712 (O_712,N_13364,N_14129);
nor UO_713 (O_713,N_12582,N_12689);
or UO_714 (O_714,N_12399,N_14158);
nand UO_715 (O_715,N_14108,N_14604);
nand UO_716 (O_716,N_13326,N_14362);
nand UO_717 (O_717,N_13608,N_13152);
or UO_718 (O_718,N_14583,N_12864);
and UO_719 (O_719,N_14285,N_13234);
nand UO_720 (O_720,N_14465,N_14344);
nand UO_721 (O_721,N_14730,N_13952);
nand UO_722 (O_722,N_14691,N_12613);
and UO_723 (O_723,N_12605,N_12379);
nand UO_724 (O_724,N_13560,N_12473);
or UO_725 (O_725,N_13909,N_12276);
and UO_726 (O_726,N_14694,N_12431);
nor UO_727 (O_727,N_12926,N_13061);
nor UO_728 (O_728,N_13992,N_13082);
nand UO_729 (O_729,N_13404,N_13160);
nor UO_730 (O_730,N_13436,N_12422);
and UO_731 (O_731,N_13226,N_13401);
or UO_732 (O_732,N_12163,N_14440);
nor UO_733 (O_733,N_14790,N_14030);
nand UO_734 (O_734,N_14125,N_12577);
nand UO_735 (O_735,N_13098,N_12948);
nor UO_736 (O_736,N_12464,N_13162);
or UO_737 (O_737,N_13028,N_14581);
nand UO_738 (O_738,N_14264,N_12825);
or UO_739 (O_739,N_14445,N_13523);
or UO_740 (O_740,N_13943,N_14503);
nor UO_741 (O_741,N_12880,N_12778);
and UO_742 (O_742,N_12813,N_13377);
nor UO_743 (O_743,N_12723,N_14436);
nand UO_744 (O_744,N_14104,N_14358);
and UO_745 (O_745,N_12929,N_14650);
nor UO_746 (O_746,N_13832,N_13915);
nor UO_747 (O_747,N_14960,N_14754);
or UO_748 (O_748,N_14331,N_13916);
nand UO_749 (O_749,N_14347,N_13862);
nor UO_750 (O_750,N_13987,N_13221);
and UO_751 (O_751,N_14810,N_14130);
and UO_752 (O_752,N_14166,N_13269);
or UO_753 (O_753,N_12242,N_14069);
nor UO_754 (O_754,N_12824,N_14533);
and UO_755 (O_755,N_14026,N_14792);
or UO_756 (O_756,N_12769,N_13191);
and UO_757 (O_757,N_14670,N_13042);
and UO_758 (O_758,N_13803,N_13047);
and UO_759 (O_759,N_12253,N_14320);
nand UO_760 (O_760,N_12581,N_14611);
xor UO_761 (O_761,N_13176,N_13889);
nor UO_762 (O_762,N_14742,N_12351);
nand UO_763 (O_763,N_13541,N_12525);
or UO_764 (O_764,N_13394,N_12835);
and UO_765 (O_765,N_13967,N_12917);
and UO_766 (O_766,N_14729,N_12491);
nor UO_767 (O_767,N_13830,N_14043);
and UO_768 (O_768,N_13325,N_14418);
and UO_769 (O_769,N_12761,N_12644);
or UO_770 (O_770,N_12489,N_12898);
nor UO_771 (O_771,N_13617,N_14382);
and UO_772 (O_772,N_13041,N_12316);
nor UO_773 (O_773,N_14429,N_14692);
or UO_774 (O_774,N_12021,N_13351);
nor UO_775 (O_775,N_13846,N_13223);
nand UO_776 (O_776,N_12104,N_12403);
and UO_777 (O_777,N_13293,N_13508);
nor UO_778 (O_778,N_13550,N_13927);
nand UO_779 (O_779,N_12758,N_12251);
nand UO_780 (O_780,N_12606,N_12383);
and UO_781 (O_781,N_14438,N_12188);
and UO_782 (O_782,N_13220,N_14087);
and UO_783 (O_783,N_12859,N_13616);
nor UO_784 (O_784,N_12802,N_13336);
and UO_785 (O_785,N_12563,N_13804);
nor UO_786 (O_786,N_12097,N_13333);
nand UO_787 (O_787,N_12937,N_13270);
nand UO_788 (O_788,N_13381,N_13950);
nor UO_789 (O_789,N_13831,N_12557);
or UO_790 (O_790,N_13933,N_14718);
nand UO_791 (O_791,N_13408,N_14179);
nor UO_792 (O_792,N_12346,N_14840);
and UO_793 (O_793,N_14254,N_13280);
and UO_794 (O_794,N_14098,N_12768);
and UO_795 (O_795,N_14333,N_12123);
nand UO_796 (O_796,N_12729,N_13876);
and UO_797 (O_797,N_13865,N_12392);
nor UO_798 (O_798,N_14327,N_12441);
or UO_799 (O_799,N_14755,N_13647);
nand UO_800 (O_800,N_13249,N_14605);
nand UO_801 (O_801,N_13204,N_14571);
nor UO_802 (O_802,N_14447,N_13514);
and UO_803 (O_803,N_14910,N_14267);
nor UO_804 (O_804,N_12545,N_14630);
nand UO_805 (O_805,N_12635,N_13756);
and UO_806 (O_806,N_12179,N_12108);
or UO_807 (O_807,N_14509,N_12895);
and UO_808 (O_808,N_14593,N_12518);
nor UO_809 (O_809,N_14986,N_13409);
nor UO_810 (O_810,N_14420,N_12486);
nand UO_811 (O_811,N_13978,N_13556);
and UO_812 (O_812,N_13414,N_13088);
or UO_813 (O_813,N_13863,N_14020);
and UO_814 (O_814,N_12107,N_13338);
nand UO_815 (O_815,N_13535,N_13861);
nor UO_816 (O_816,N_14641,N_13528);
or UO_817 (O_817,N_12110,N_12287);
and UO_818 (O_818,N_12580,N_12357);
and UO_819 (O_819,N_12260,N_12194);
or UO_820 (O_820,N_12190,N_13802);
nor UO_821 (O_821,N_12059,N_12087);
or UO_822 (O_822,N_14066,N_12315);
or UO_823 (O_823,N_13873,N_14835);
nor UO_824 (O_824,N_14631,N_14337);
nor UO_825 (O_825,N_13259,N_14480);
nand UO_826 (O_826,N_14002,N_14892);
nor UO_827 (O_827,N_13513,N_13656);
nor UO_828 (O_828,N_12984,N_13288);
nand UO_829 (O_829,N_14662,N_12067);
nand UO_830 (O_830,N_14449,N_13801);
and UO_831 (O_831,N_12532,N_12675);
nor UO_832 (O_832,N_12038,N_13425);
or UO_833 (O_833,N_12981,N_12068);
nor UO_834 (O_834,N_14342,N_14153);
and UO_835 (O_835,N_14843,N_13688);
nand UO_836 (O_836,N_12055,N_12891);
or UO_837 (O_837,N_14667,N_14647);
or UO_838 (O_838,N_14750,N_13576);
nand UO_839 (O_839,N_13810,N_12265);
or UO_840 (O_840,N_13254,N_12826);
and UO_841 (O_841,N_13975,N_14978);
and UO_842 (O_842,N_12794,N_12081);
or UO_843 (O_843,N_14416,N_12153);
or UO_844 (O_844,N_14156,N_14114);
nor UO_845 (O_845,N_13548,N_14621);
and UO_846 (O_846,N_12913,N_14959);
and UO_847 (O_847,N_13156,N_13145);
and UO_848 (O_848,N_12020,N_14249);
nor UO_849 (O_849,N_13976,N_12626);
and UO_850 (O_850,N_13137,N_13476);
nor UO_851 (O_851,N_14219,N_14093);
nor UO_852 (O_852,N_13089,N_12326);
or UO_853 (O_853,N_12530,N_14434);
or UO_854 (O_854,N_13175,N_13417);
and UO_855 (O_855,N_13347,N_14698);
and UO_856 (O_856,N_14481,N_13549);
nor UO_857 (O_857,N_14768,N_14314);
nor UO_858 (O_858,N_14628,N_14914);
and UO_859 (O_859,N_14477,N_13006);
or UO_860 (O_860,N_12517,N_13870);
nor UO_861 (O_861,N_14038,N_12010);
nand UO_862 (O_862,N_13713,N_12779);
or UO_863 (O_863,N_12865,N_13837);
and UO_864 (O_864,N_13400,N_12313);
and UO_865 (O_865,N_13463,N_14177);
nor UO_866 (O_866,N_13500,N_12832);
and UO_867 (O_867,N_12784,N_14834);
nor UO_868 (O_868,N_12400,N_12565);
and UO_869 (O_869,N_12634,N_13081);
nand UO_870 (O_870,N_12703,N_12731);
nor UO_871 (O_871,N_14137,N_14328);
nand UO_872 (O_872,N_13495,N_14273);
and UO_873 (O_873,N_14540,N_14248);
nor UO_874 (O_874,N_12482,N_13399);
or UO_875 (O_875,N_14302,N_13768);
or UO_876 (O_876,N_12057,N_14825);
nand UO_877 (O_877,N_12100,N_13991);
nor UO_878 (O_878,N_12321,N_14851);
nor UO_879 (O_879,N_12456,N_14529);
nand UO_880 (O_880,N_13695,N_13633);
nor UO_881 (O_881,N_12496,N_12609);
and UO_882 (O_882,N_13946,N_12420);
or UO_883 (O_883,N_12866,N_14925);
xnor UO_884 (O_884,N_12551,N_13107);
nand UO_885 (O_885,N_12314,N_12423);
and UO_886 (O_886,N_12876,N_12524);
nand UO_887 (O_887,N_13658,N_14805);
nand UO_888 (O_888,N_12911,N_13063);
nor UO_889 (O_889,N_12775,N_14633);
and UO_890 (O_890,N_14846,N_12554);
or UO_891 (O_891,N_13839,N_14734);
and UO_892 (O_892,N_13667,N_14916);
and UO_893 (O_893,N_13075,N_13811);
xnor UO_894 (O_894,N_14135,N_13546);
nand UO_895 (O_895,N_14065,N_13108);
nand UO_896 (O_896,N_14146,N_14475);
nand UO_897 (O_897,N_14525,N_14793);
nor UO_898 (O_898,N_12836,N_13885);
nor UO_899 (O_899,N_14661,N_14523);
nand UO_900 (O_900,N_13606,N_12252);
nand UO_901 (O_901,N_12204,N_13127);
and UO_902 (O_902,N_12647,N_13684);
nor UO_903 (O_903,N_14164,N_14687);
nand UO_904 (O_904,N_13071,N_14131);
or UO_905 (O_905,N_13902,N_14735);
nor UO_906 (O_906,N_14998,N_13970);
nand UO_907 (O_907,N_13736,N_12370);
or UO_908 (O_908,N_13887,N_12036);
and UO_909 (O_909,N_13590,N_14271);
nor UO_910 (O_910,N_12099,N_14865);
nor UO_911 (O_911,N_14502,N_14787);
nand UO_912 (O_912,N_13237,N_13312);
nor UO_913 (O_913,N_12912,N_13653);
nand UO_914 (O_914,N_13247,N_13015);
or UO_915 (O_915,N_13416,N_13273);
nor UO_916 (O_916,N_13703,N_12842);
nor UO_917 (O_917,N_14973,N_12559);
nand UO_918 (O_918,N_12897,N_13443);
nor UO_919 (O_919,N_14090,N_13243);
and UO_920 (O_920,N_12187,N_13140);
or UO_921 (O_921,N_13482,N_12712);
nand UO_922 (O_922,N_12576,N_13303);
or UO_923 (O_923,N_14149,N_13779);
nor UO_924 (O_924,N_14626,N_14364);
or UO_925 (O_925,N_14210,N_13780);
or UO_926 (O_926,N_12830,N_12143);
nor UO_927 (O_927,N_13896,N_12135);
and UO_928 (O_928,N_12001,N_12583);
nor UO_929 (O_929,N_12687,N_13583);
and UO_930 (O_930,N_12648,N_12889);
or UO_931 (O_931,N_13571,N_14951);
or UO_932 (O_932,N_12311,N_12443);
nor UO_933 (O_933,N_14060,N_12942);
or UO_934 (O_934,N_13823,N_12201);
nand UO_935 (O_935,N_14062,N_13361);
and UO_936 (O_936,N_12958,N_14898);
nor UO_937 (O_937,N_14261,N_12732);
or UO_938 (O_938,N_14055,N_13301);
or UO_939 (O_939,N_12740,N_13857);
nor UO_940 (O_940,N_13794,N_13977);
nand UO_941 (O_941,N_13448,N_14162);
nand UO_942 (O_942,N_14899,N_14257);
xor UO_943 (O_943,N_14336,N_12969);
nand UO_944 (O_944,N_12944,N_14913);
nor UO_945 (O_945,N_14711,N_14171);
nand UO_946 (O_946,N_12278,N_12658);
nor UO_947 (O_947,N_14117,N_13324);
or UO_948 (O_948,N_14144,N_13579);
or UO_949 (O_949,N_12849,N_12674);
nand UO_950 (O_950,N_12405,N_14802);
or UO_951 (O_951,N_14075,N_14854);
and UO_952 (O_952,N_12661,N_14236);
and UO_953 (O_953,N_13405,N_12906);
or UO_954 (O_954,N_12049,N_13584);
and UO_955 (O_955,N_13319,N_12662);
nand UO_956 (O_956,N_13064,N_14487);
nor UO_957 (O_957,N_12446,N_12872);
nor UO_958 (O_958,N_12437,N_14791);
and UO_959 (O_959,N_14536,N_14653);
and UO_960 (O_960,N_12811,N_12429);
and UO_961 (O_961,N_14680,N_13450);
and UO_962 (O_962,N_13440,N_14572);
and UO_963 (O_963,N_14693,N_12515);
or UO_964 (O_964,N_12900,N_13202);
or UO_965 (O_965,N_12744,N_14196);
nor UO_966 (O_966,N_14806,N_13382);
and UO_967 (O_967,N_14262,N_14204);
and UO_968 (O_968,N_14794,N_13956);
nor UO_969 (O_969,N_12856,N_13682);
or UO_970 (O_970,N_13240,N_14201);
nand UO_971 (O_971,N_13675,N_14410);
or UO_972 (O_972,N_14033,N_12522);
or UO_973 (O_973,N_14921,N_12218);
nand UO_974 (O_974,N_12710,N_14334);
nor UO_975 (O_975,N_14376,N_14695);
or UO_976 (O_976,N_13315,N_14032);
or UO_977 (O_977,N_13258,N_13138);
nand UO_978 (O_978,N_13144,N_12695);
nand UO_979 (O_979,N_14866,N_14478);
nand UO_980 (O_980,N_13899,N_12863);
nand UO_981 (O_981,N_14165,N_12112);
and UO_982 (O_982,N_12821,N_12809);
nor UO_983 (O_983,N_12355,N_13898);
and UO_984 (O_984,N_12781,N_12799);
and UO_985 (O_985,N_13106,N_13461);
or UO_986 (O_986,N_13834,N_14859);
or UO_987 (O_987,N_13890,N_12033);
and UO_988 (O_988,N_12932,N_14815);
or UO_989 (O_989,N_13452,N_12064);
nor UO_990 (O_990,N_12921,N_12805);
or UO_991 (O_991,N_14796,N_14411);
and UO_992 (O_992,N_12397,N_14602);
nand UO_993 (O_993,N_13558,N_13951);
nand UO_994 (O_994,N_13592,N_14338);
or UO_995 (O_995,N_14549,N_14829);
nand UO_996 (O_996,N_13279,N_12146);
and UO_997 (O_997,N_12602,N_13363);
and UO_998 (O_998,N_14721,N_12659);
or UO_999 (O_999,N_13195,N_14388);
nor UO_1000 (O_1000,N_14081,N_13842);
xor UO_1001 (O_1001,N_13990,N_14841);
and UO_1002 (O_1002,N_12534,N_14198);
or UO_1003 (O_1003,N_13402,N_13881);
nor UO_1004 (O_1004,N_12416,N_13570);
and UO_1005 (O_1005,N_14903,N_14453);
xor UO_1006 (O_1006,N_13843,N_13504);
or UO_1007 (O_1007,N_13370,N_13721);
nor UO_1008 (O_1008,N_12079,N_14528);
nand UO_1009 (O_1009,N_14952,N_12839);
and UO_1010 (O_1010,N_14101,N_14600);
or UO_1011 (O_1011,N_13648,N_14363);
nand UO_1012 (O_1012,N_14763,N_13172);
nand UO_1013 (O_1013,N_12193,N_13151);
or UO_1014 (O_1014,N_12827,N_13165);
nor UO_1015 (O_1015,N_12377,N_13018);
nand UO_1016 (O_1016,N_13116,N_12879);
or UO_1017 (O_1017,N_13730,N_13272);
or UO_1018 (O_1018,N_12459,N_14379);
or UO_1019 (O_1019,N_14738,N_12503);
nor UO_1020 (O_1020,N_14783,N_13199);
nand UO_1021 (O_1021,N_14500,N_13344);
nor UO_1022 (O_1022,N_13917,N_12641);
and UO_1023 (O_1023,N_13327,N_13777);
and UO_1024 (O_1024,N_13561,N_14059);
nand UO_1025 (O_1025,N_14001,N_14050);
nand UO_1026 (O_1026,N_13494,N_12138);
nand UO_1027 (O_1027,N_12922,N_14524);
nand UO_1028 (O_1028,N_12273,N_12339);
nor UO_1029 (O_1029,N_12807,N_13795);
nand UO_1030 (O_1030,N_13687,N_13130);
or UO_1031 (O_1031,N_13281,N_14159);
and UO_1032 (O_1032,N_14079,N_12347);
xnor UO_1033 (O_1033,N_12266,N_12031);
nand UO_1034 (O_1034,N_12442,N_12156);
nor UO_1035 (O_1035,N_14643,N_12639);
or UO_1036 (O_1036,N_12016,N_12000);
nor UO_1037 (O_1037,N_12800,N_13348);
nand UO_1038 (O_1038,N_13706,N_12810);
or UO_1039 (O_1039,N_14853,N_12893);
and UO_1040 (O_1040,N_12468,N_12404);
nand UO_1041 (O_1041,N_13725,N_12774);
nand UO_1042 (O_1042,N_14191,N_13821);
and UO_1043 (O_1043,N_13993,N_14823);
or UO_1044 (O_1044,N_12022,N_14710);
nor UO_1045 (O_1045,N_13024,N_14350);
nor UO_1046 (O_1046,N_14409,N_13696);
or UO_1047 (O_1047,N_12149,N_12335);
or UO_1048 (O_1048,N_12217,N_12162);
and UO_1049 (O_1049,N_14483,N_12540);
nand UO_1050 (O_1050,N_14736,N_14407);
nor UO_1051 (O_1051,N_14476,N_14957);
and UO_1052 (O_1052,N_13174,N_12454);
or UO_1053 (O_1053,N_12934,N_13963);
nor UO_1054 (O_1054,N_12358,N_14992);
and UO_1055 (O_1055,N_12296,N_14844);
nand UO_1056 (O_1056,N_14111,N_14644);
or UO_1057 (O_1057,N_14291,N_14861);
or UO_1058 (O_1058,N_13710,N_14470);
nor UO_1059 (O_1059,N_12844,N_13224);
nand UO_1060 (O_1060,N_14435,N_12620);
and UO_1061 (O_1061,N_14288,N_14195);
and UO_1062 (O_1062,N_12881,N_12672);
nor UO_1063 (O_1063,N_13555,N_13418);
or UO_1064 (O_1064,N_12765,N_14801);
or UO_1065 (O_1065,N_12502,N_13161);
nand UO_1066 (O_1066,N_12875,N_13577);
or UO_1067 (O_1067,N_12616,N_14554);
and UO_1068 (O_1068,N_12954,N_13371);
nor UO_1069 (O_1069,N_12494,N_12928);
and UO_1070 (O_1070,N_14256,N_12692);
nor UO_1071 (O_1071,N_12008,N_13255);
nor UO_1072 (O_1072,N_13055,N_12649);
and UO_1073 (O_1073,N_12631,N_14614);
or UO_1074 (O_1074,N_13754,N_13099);
or UO_1075 (O_1075,N_12686,N_12034);
or UO_1076 (O_1076,N_12432,N_12094);
nor UO_1077 (O_1077,N_13198,N_13749);
nor UO_1078 (O_1078,N_14332,N_12727);
or UO_1079 (O_1079,N_13054,N_14237);
nand UO_1080 (O_1080,N_12959,N_12144);
nor UO_1081 (O_1081,N_13182,N_14759);
and UO_1082 (O_1082,N_14121,N_14116);
nor UO_1083 (O_1083,N_13056,N_14022);
nor UO_1084 (O_1084,N_12730,N_14706);
and UO_1085 (O_1085,N_13439,N_13021);
or UO_1086 (O_1086,N_14764,N_12271);
or UO_1087 (O_1087,N_12822,N_14290);
and UO_1088 (O_1088,N_13131,N_13825);
and UO_1089 (O_1089,N_12925,N_12542);
nor UO_1090 (O_1090,N_13104,N_14190);
nor UO_1091 (O_1091,N_13731,N_13252);
and UO_1092 (O_1092,N_14175,N_13806);
nand UO_1093 (O_1093,N_13553,N_13651);
nand UO_1094 (O_1094,N_13882,N_14816);
nor UO_1095 (O_1095,N_13566,N_13888);
nor UO_1096 (O_1096,N_13188,N_13894);
or UO_1097 (O_1097,N_14127,N_13770);
nand UO_1098 (O_1098,N_14412,N_13643);
and UO_1099 (O_1099,N_12861,N_12209);
or UO_1100 (O_1100,N_14390,N_14629);
nand UO_1101 (O_1101,N_12262,N_14690);
nor UO_1102 (O_1102,N_12632,N_12578);
and UO_1103 (O_1103,N_13619,N_14292);
or UO_1104 (O_1104,N_12438,N_14370);
or UO_1105 (O_1105,N_12816,N_13124);
or UO_1106 (O_1106,N_13014,N_14867);
or UO_1107 (O_1107,N_12061,N_14019);
nand UO_1108 (O_1108,N_13060,N_12555);
or UO_1109 (O_1109,N_13604,N_13591);
nor UO_1110 (O_1110,N_12132,N_12831);
nand UO_1111 (O_1111,N_14414,N_12562);
nand UO_1112 (O_1112,N_13886,N_12560);
or UO_1113 (O_1113,N_12243,N_13995);
nand UO_1114 (O_1114,N_13329,N_14985);
nor UO_1115 (O_1115,N_13306,N_12628);
nand UO_1116 (O_1116,N_13734,N_13115);
nand UO_1117 (O_1117,N_14607,N_14799);
or UO_1118 (O_1118,N_14777,N_12803);
and UO_1119 (O_1119,N_13924,N_14260);
or UO_1120 (O_1120,N_12599,N_13411);
nor UO_1121 (O_1121,N_14901,N_12052);
nor UO_1122 (O_1122,N_14610,N_13923);
or UO_1123 (O_1123,N_12199,N_12655);
or UO_1124 (O_1124,N_14063,N_12770);
nand UO_1125 (O_1125,N_13250,N_14996);
and UO_1126 (O_1126,N_14152,N_12160);
and UO_1127 (O_1127,N_12706,N_13257);
nand UO_1128 (O_1128,N_14246,N_13793);
nand UO_1129 (O_1129,N_13342,N_13937);
nor UO_1130 (O_1130,N_13294,N_13080);
nand UO_1131 (O_1131,N_14186,N_14720);
nor UO_1132 (O_1132,N_13241,N_13918);
and UO_1133 (O_1133,N_14473,N_13597);
nor UO_1134 (O_1134,N_12980,N_14176);
nand UO_1135 (O_1135,N_14713,N_13189);
or UO_1136 (O_1136,N_12182,N_12436);
nand UO_1137 (O_1137,N_12425,N_12338);
and UO_1138 (O_1138,N_13068,N_14857);
nand UO_1139 (O_1139,N_14664,N_12398);
and UO_1140 (O_1140,N_13930,N_14850);
nand UO_1141 (O_1141,N_14070,N_12520);
or UO_1142 (O_1142,N_14496,N_12877);
nand UO_1143 (O_1143,N_12506,N_12782);
or UO_1144 (O_1144,N_12544,N_14938);
nor UO_1145 (O_1145,N_14466,N_14686);
and UO_1146 (O_1146,N_13209,N_13827);
nand UO_1147 (O_1147,N_14789,N_14084);
nor UO_1148 (O_1148,N_12936,N_12629);
or UO_1149 (O_1149,N_12237,N_14564);
nor UO_1150 (O_1150,N_13738,N_14396);
and UO_1151 (O_1151,N_12300,N_14728);
and UO_1152 (O_1152,N_13748,N_12884);
nor UO_1153 (O_1153,N_12413,N_14091);
and UO_1154 (O_1154,N_14058,N_14298);
and UO_1155 (O_1155,N_13360,N_13192);
and UO_1156 (O_1156,N_12175,N_13036);
and UO_1157 (O_1157,N_13724,N_14380);
or UO_1158 (O_1158,N_13158,N_13155);
and UO_1159 (O_1159,N_13005,N_14688);
and UO_1160 (O_1160,N_12548,N_14991);
nor UO_1161 (O_1161,N_13552,N_14286);
nand UO_1162 (O_1162,N_13867,N_12235);
nand UO_1163 (O_1163,N_14702,N_14847);
and UO_1164 (O_1164,N_13062,N_12801);
nor UO_1165 (O_1165,N_14580,N_13735);
nor UO_1166 (O_1166,N_12124,N_12585);
and UO_1167 (O_1167,N_12184,N_13261);
nand UO_1168 (O_1168,N_13091,N_13083);
or UO_1169 (O_1169,N_13700,N_12780);
and UO_1170 (O_1170,N_13798,N_12870);
and UO_1171 (O_1171,N_12737,N_12590);
nand UO_1172 (O_1172,N_12660,N_12645);
and UO_1173 (O_1173,N_14995,N_13375);
nor UO_1174 (O_1174,N_14948,N_13544);
nand UO_1175 (O_1175,N_13369,N_12050);
or UO_1176 (O_1176,N_14099,N_14839);
nor UO_1177 (O_1177,N_12733,N_14601);
or UO_1178 (O_1178,N_14679,N_12103);
and UO_1179 (O_1179,N_14235,N_14048);
or UO_1180 (O_1180,N_12570,N_13190);
and UO_1181 (O_1181,N_12095,N_14904);
nor UO_1182 (O_1182,N_12914,N_13800);
and UO_1183 (O_1183,N_12935,N_12258);
nor UO_1184 (O_1184,N_14306,N_14035);
nand UO_1185 (O_1185,N_13000,N_13864);
nand UO_1186 (O_1186,N_14147,N_13286);
nand UO_1187 (O_1187,N_14276,N_14689);
and UO_1188 (O_1188,N_12868,N_13488);
and UO_1189 (O_1189,N_13491,N_12114);
nand UO_1190 (O_1190,N_14895,N_13126);
nand UO_1191 (O_1191,N_14499,N_12700);
and UO_1192 (O_1192,N_14423,N_12152);
nor UO_1193 (O_1193,N_12873,N_14820);
nor UO_1194 (O_1194,N_12857,N_13742);
nor UO_1195 (O_1195,N_13540,N_12817);
nand UO_1196 (O_1196,N_12910,N_14220);
nor UO_1197 (O_1197,N_12150,N_12147);
and UO_1198 (O_1198,N_14064,N_13866);
nand UO_1199 (O_1199,N_12071,N_13690);
nand UO_1200 (O_1200,N_13374,N_13242);
nor UO_1201 (O_1201,N_12843,N_13262);
and UO_1202 (O_1202,N_14578,N_13278);
or UO_1203 (O_1203,N_13691,N_14142);
and UO_1204 (O_1204,N_12457,N_14731);
nor UO_1205 (O_1205,N_13914,N_12890);
nor UO_1206 (O_1206,N_14780,N_14699);
and UO_1207 (O_1207,N_12065,N_12753);
nor UO_1208 (O_1208,N_14009,N_12401);
or UO_1209 (O_1209,N_13787,N_13766);
or UO_1210 (O_1210,N_13307,N_14537);
nand UO_1211 (O_1211,N_13396,N_14319);
nand UO_1212 (O_1212,N_13516,N_14656);
nor UO_1213 (O_1213,N_14676,N_14752);
or UO_1214 (O_1214,N_14612,N_13878);
nand UO_1215 (O_1215,N_14197,N_12161);
or UO_1216 (O_1216,N_12393,N_12927);
nand UO_1217 (O_1217,N_12493,N_13601);
nor UO_1218 (O_1218,N_13299,N_14654);
and UO_1219 (O_1219,N_12967,N_12232);
nor UO_1220 (O_1220,N_13133,N_12685);
and UO_1221 (O_1221,N_14947,N_12177);
nor UO_1222 (O_1222,N_12359,N_12796);
nor UO_1223 (O_1223,N_12462,N_13432);
nor UO_1224 (O_1224,N_13248,N_14800);
nand UO_1225 (O_1225,N_12887,N_13413);
and UO_1226 (O_1226,N_13321,N_13388);
or UO_1227 (O_1227,N_13392,N_12227);
or UO_1228 (O_1228,N_14192,N_13086);
or UO_1229 (O_1229,N_12214,N_12305);
or UO_1230 (O_1230,N_13379,N_14361);
nand UO_1231 (O_1231,N_12122,N_12069);
and UO_1232 (O_1232,N_13693,N_13509);
nor UO_1233 (O_1233,N_12797,N_13874);
or UO_1234 (O_1234,N_13729,N_13660);
nand UO_1235 (O_1235,N_13178,N_13539);
and UO_1236 (O_1236,N_13076,N_14908);
nor UO_1237 (O_1237,N_14547,N_12117);
and UO_1238 (O_1238,N_13423,N_14945);
nand UO_1239 (O_1239,N_14199,N_14053);
nor UO_1240 (O_1240,N_14707,N_12946);
nor UO_1241 (O_1241,N_14386,N_13122);
nor UO_1242 (O_1242,N_13026,N_13783);
and UO_1243 (O_1243,N_12412,N_13657);
nand UO_1244 (O_1244,N_14140,N_12041);
nand UO_1245 (O_1245,N_13387,N_14045);
nand UO_1246 (O_1246,N_14112,N_13649);
nor UO_1247 (O_1247,N_13892,N_13640);
nor UO_1248 (O_1248,N_13103,N_12759);
or UO_1249 (O_1249,N_13668,N_12793);
nor UO_1250 (O_1250,N_14495,N_12173);
or UO_1251 (O_1251,N_13599,N_13359);
nand UO_1252 (O_1252,N_13253,N_13678);
nor UO_1253 (O_1253,N_12078,N_12027);
or UO_1254 (O_1254,N_14031,N_12086);
and UO_1255 (O_1255,N_13559,N_13530);
nand UO_1256 (O_1256,N_14757,N_13879);
nor UO_1257 (O_1257,N_12430,N_12716);
or UO_1258 (O_1258,N_12752,N_14727);
nor UO_1259 (O_1259,N_12965,N_13921);
nand UO_1260 (O_1260,N_14402,N_14489);
nand UO_1261 (O_1261,N_13407,N_14427);
and UO_1262 (O_1262,N_13368,N_13173);
and UO_1263 (O_1263,N_14860,N_12092);
or UO_1264 (O_1264,N_13027,N_12619);
nand UO_1265 (O_1265,N_14003,N_13981);
nor UO_1266 (O_1266,N_13489,N_14592);
nor UO_1267 (O_1267,N_14425,N_13641);
and UO_1268 (O_1268,N_14505,N_14014);
and UO_1269 (O_1269,N_14943,N_13087);
nand UO_1270 (O_1270,N_12270,N_13274);
nor UO_1271 (O_1271,N_13868,N_13908);
nand UO_1272 (O_1272,N_12136,N_12783);
and UO_1273 (O_1273,N_14270,N_12667);
and UO_1274 (O_1274,N_13763,N_12608);
nor UO_1275 (O_1275,N_14096,N_12949);
and UO_1276 (O_1276,N_12378,N_12408);
nand UO_1277 (O_1277,N_12977,N_14663);
or UO_1278 (O_1278,N_14696,N_13469);
nand UO_1279 (O_1279,N_14148,N_13340);
and UO_1280 (O_1280,N_12198,N_14756);
nand UO_1281 (O_1281,N_14933,N_13955);
or UO_1282 (O_1282,N_14964,N_13113);
nand UO_1283 (O_1283,N_13962,N_14511);
or UO_1284 (O_1284,N_12964,N_12151);
and UO_1285 (O_1285,N_14119,N_12541);
and UO_1286 (O_1286,N_14250,N_14598);
nor UO_1287 (O_1287,N_13612,N_14873);
nand UO_1288 (O_1288,N_12947,N_12427);
or UO_1289 (O_1289,N_13235,N_12846);
or UO_1290 (O_1290,N_14169,N_12042);
nor UO_1291 (O_1291,N_13860,N_12481);
and UO_1292 (O_1292,N_14937,N_13522);
or UO_1293 (O_1293,N_12145,N_14936);
nor UO_1294 (O_1294,N_14054,N_13460);
and UO_1295 (O_1295,N_13926,N_12537);
and UO_1296 (O_1296,N_13893,N_12331);
or UO_1297 (O_1297,N_13822,N_14456);
and UO_1298 (O_1298,N_12226,N_13453);
or UO_1299 (O_1299,N_13183,N_13935);
and UO_1300 (O_1300,N_14907,N_13744);
nand UO_1301 (O_1301,N_13849,N_12084);
nor UO_1302 (O_1302,N_13877,N_12625);
nand UO_1303 (O_1303,N_12290,N_14168);
and UO_1304 (O_1304,N_13771,N_14817);
nor UO_1305 (O_1305,N_12776,N_14431);
nand UO_1306 (O_1306,N_12154,N_12389);
and UO_1307 (O_1307,N_12304,N_13477);
nand UO_1308 (O_1308,N_13854,N_14606);
nor UO_1309 (O_1309,N_12090,N_13123);
nand UO_1310 (O_1310,N_14917,N_12302);
nand UO_1311 (O_1311,N_12334,N_13025);
nor UO_1312 (O_1312,N_12850,N_13356);
and UO_1313 (O_1313,N_12650,N_13762);
nor UO_1314 (O_1314,N_14151,N_12711);
or UO_1315 (O_1315,N_13466,N_13201);
nand UO_1316 (O_1316,N_13267,N_12348);
nor UO_1317 (O_1317,N_12210,N_13058);
and UO_1318 (O_1318,N_13645,N_13781);
and UO_1319 (O_1319,N_12612,N_13011);
nor UO_1320 (O_1320,N_14241,N_13760);
nand UO_1321 (O_1321,N_13585,N_12788);
or UO_1322 (O_1322,N_14193,N_12490);
nor UO_1323 (O_1323,N_12974,N_14894);
nand UO_1324 (O_1324,N_14240,N_14296);
nor UO_1325 (O_1325,N_12308,N_12046);
or UO_1326 (O_1326,N_12418,N_14335);
and UO_1327 (O_1327,N_13697,N_12352);
nand UO_1328 (O_1328,N_12514,N_12312);
and UO_1329 (O_1329,N_13895,N_13851);
nand UO_1330 (O_1330,N_14658,N_14234);
nand UO_1331 (O_1331,N_13625,N_12170);
and UO_1332 (O_1332,N_14463,N_14138);
and UO_1333 (O_1333,N_14987,N_14919);
and UO_1334 (O_1334,N_12812,N_14737);
or UO_1335 (O_1335,N_14634,N_14842);
or UO_1336 (O_1336,N_13674,N_12139);
or UO_1337 (O_1337,N_12180,N_14206);
nand UO_1338 (O_1338,N_13029,N_14242);
and UO_1339 (O_1339,N_13390,N_13537);
nor UO_1340 (O_1340,N_12617,N_14858);
nand UO_1341 (O_1341,N_14036,N_12501);
nand UO_1342 (O_1342,N_14324,N_14882);
or UO_1343 (O_1343,N_12073,N_12098);
and UO_1344 (O_1344,N_14648,N_13607);
nor UO_1345 (O_1345,N_14056,N_14622);
nor UO_1346 (O_1346,N_12885,N_14893);
nand UO_1347 (O_1347,N_14929,N_13134);
nand UO_1348 (O_1348,N_13998,N_14709);
nand UO_1349 (O_1349,N_14239,N_13129);
or UO_1350 (O_1350,N_13757,N_12283);
nor UO_1351 (O_1351,N_13435,N_13184);
and UO_1352 (O_1352,N_14155,N_12591);
and UO_1353 (O_1353,N_14309,N_14085);
nor UO_1354 (O_1354,N_14935,N_12277);
and UO_1355 (O_1355,N_14492,N_12157);
nor UO_1356 (O_1356,N_12600,N_14949);
or UO_1357 (O_1357,N_14590,N_14746);
or UO_1358 (O_1358,N_12671,N_13708);
nor UO_1359 (O_1359,N_14640,N_14891);
and UO_1360 (O_1360,N_12414,N_14958);
or UO_1361 (O_1361,N_13714,N_12952);
or UO_1362 (O_1362,N_14701,N_14603);
nand UO_1363 (O_1363,N_12804,N_12202);
nand UO_1364 (O_1364,N_12726,N_13067);
nor UO_1365 (O_1365,N_12724,N_12183);
xor UO_1366 (O_1366,N_13395,N_13732);
and UO_1367 (O_1367,N_14775,N_13727);
and UO_1368 (O_1368,N_12604,N_14247);
nand UO_1369 (O_1369,N_12552,N_12452);
nor UO_1370 (O_1370,N_12216,N_13817);
nand UO_1371 (O_1371,N_13475,N_13816);
or UO_1372 (O_1372,N_12622,N_14989);
or UO_1373 (O_1373,N_12751,N_13403);
nand UO_1374 (O_1374,N_12950,N_12322);
nand UO_1375 (O_1375,N_14441,N_14574);
and UO_1376 (O_1376,N_14023,N_13853);
nand UO_1377 (O_1377,N_13638,N_12792);
nand UO_1378 (O_1378,N_14078,N_14627);
nor UO_1379 (O_1379,N_12682,N_12279);
nand UO_1380 (O_1380,N_14222,N_14357);
or UO_1381 (O_1381,N_12366,N_13574);
and UO_1382 (O_1382,N_13767,N_12908);
or UO_1383 (O_1383,N_14269,N_13053);
and UO_1384 (O_1384,N_12458,N_14570);
and UO_1385 (O_1385,N_13728,N_12833);
or UO_1386 (O_1386,N_13236,N_12113);
nand UO_1387 (O_1387,N_13349,N_13479);
and UO_1388 (O_1388,N_12158,N_13701);
nand UO_1389 (O_1389,N_12511,N_12973);
or UO_1390 (O_1390,N_13994,N_12111);
nand UO_1391 (O_1391,N_13487,N_14889);
nor UO_1392 (O_1392,N_14024,N_14715);
or UO_1393 (O_1393,N_14467,N_13231);
or UO_1394 (O_1394,N_13092,N_13683);
and UO_1395 (O_1395,N_14455,N_13121);
nor UO_1396 (O_1396,N_13672,N_13855);
nor UO_1397 (O_1397,N_12597,N_12301);
nand UO_1398 (O_1398,N_13511,N_13598);
or UO_1399 (O_1399,N_13039,N_12244);
or UO_1400 (O_1400,N_13575,N_12062);
nor UO_1401 (O_1401,N_13186,N_13276);
or UO_1402 (O_1402,N_14970,N_13454);
nor UO_1403 (O_1403,N_14185,N_13758);
or UO_1404 (O_1404,N_13872,N_12448);
or UO_1405 (O_1405,N_13615,N_12029);
nor UO_1406 (O_1406,N_14221,N_13828);
and UO_1407 (O_1407,N_14398,N_12820);
or UO_1408 (O_1408,N_12361,N_12678);
nor UO_1409 (O_1409,N_12387,N_13376);
nor UO_1410 (O_1410,N_13940,N_12683);
nand UO_1411 (O_1411,N_12828,N_14831);
nor UO_1412 (O_1412,N_13284,N_14902);
nor UO_1413 (O_1413,N_12513,N_13010);
or UO_1414 (O_1414,N_12680,N_12643);
and UO_1415 (O_1415,N_12419,N_13664);
and UO_1416 (O_1416,N_14939,N_13447);
nor UO_1417 (O_1417,N_13833,N_13170);
nand UO_1418 (O_1418,N_12763,N_13268);
nor UO_1419 (O_1419,N_14008,N_14405);
or UO_1420 (O_1420,N_12223,N_12867);
or UO_1421 (O_1421,N_12673,N_14115);
or UO_1422 (O_1422,N_13154,N_13002);
and UO_1423 (O_1423,N_14546,N_13217);
and UO_1424 (O_1424,N_14428,N_12306);
nand UO_1425 (O_1425,N_13096,N_13362);
and UO_1426 (O_1426,N_14548,N_14786);
or UO_1427 (O_1427,N_14448,N_14803);
and UO_1428 (O_1428,N_12479,N_12633);
or UO_1429 (O_1429,N_12463,N_14213);
or UO_1430 (O_1430,N_13856,N_14074);
and UO_1431 (O_1431,N_12651,N_13179);
or UO_1432 (O_1432,N_13919,N_14681);
nor UO_1433 (O_1433,N_12341,N_13525);
or UO_1434 (O_1434,N_12191,N_12539);
or UO_1435 (O_1435,N_14506,N_14228);
and UO_1436 (O_1436,N_13936,N_12623);
nand UO_1437 (O_1437,N_12211,N_13009);
nor UO_1438 (O_1438,N_14375,N_13669);
nor UO_1439 (O_1439,N_14997,N_12376);
nand UO_1440 (O_1440,N_14086,N_12771);
nor UO_1441 (O_1441,N_13328,N_13297);
nor UO_1442 (O_1442,N_14212,N_12015);
or UO_1443 (O_1443,N_14227,N_13961);
nor UO_1444 (O_1444,N_13719,N_13948);
or UO_1445 (O_1445,N_14532,N_14837);
nand UO_1446 (O_1446,N_13213,N_14167);
nand UO_1447 (O_1447,N_13296,N_12905);
nor UO_1448 (O_1448,N_14797,N_13859);
nand UO_1449 (O_1449,N_14365,N_13964);
nor UO_1450 (O_1450,N_12371,N_13726);
nand UO_1451 (O_1451,N_14272,N_12492);
nand UO_1452 (O_1452,N_14244,N_14253);
nand UO_1453 (O_1453,N_13194,N_12363);
nand UO_1454 (O_1454,N_14508,N_14886);
nor UO_1455 (O_1455,N_13663,N_13850);
and UO_1456 (O_1456,N_12141,N_13233);
nand UO_1457 (O_1457,N_14983,N_12066);
and UO_1458 (O_1458,N_13275,N_12215);
and UO_1459 (O_1459,N_14067,N_14535);
nor UO_1460 (O_1460,N_14745,N_13046);
nand UO_1461 (O_1461,N_14637,N_14617);
and UO_1462 (O_1462,N_13335,N_12679);
nand UO_1463 (O_1463,N_13745,N_14021);
or UO_1464 (O_1464,N_13524,N_13966);
nand UO_1465 (O_1465,N_12247,N_13033);
or UO_1466 (O_1466,N_14326,N_12282);
xnor UO_1467 (O_1467,N_12814,N_12088);
nand UO_1468 (O_1468,N_13844,N_13629);
or UO_1469 (O_1469,N_12851,N_14491);
nor UO_1470 (O_1470,N_12543,N_14758);
nand UO_1471 (O_1471,N_13271,N_12281);
nand UO_1472 (O_1472,N_13003,N_14377);
nand UO_1473 (O_1473,N_12728,N_14649);
and UO_1474 (O_1474,N_12040,N_12003);
or UO_1475 (O_1475,N_14282,N_14095);
or UO_1476 (O_1476,N_14553,N_14313);
nand UO_1477 (O_1477,N_14354,N_14245);
and UO_1478 (O_1478,N_14953,N_14330);
nor UO_1479 (O_1479,N_12869,N_13685);
and UO_1480 (O_1480,N_14231,N_12197);
and UO_1481 (O_1481,N_12356,N_14305);
and UO_1482 (O_1482,N_14308,N_12871);
or UO_1483 (O_1483,N_13285,N_14207);
nand UO_1484 (O_1484,N_13428,N_14426);
or UO_1485 (O_1485,N_14774,N_12618);
nor UO_1486 (O_1486,N_13646,N_12512);
nor UO_1487 (O_1487,N_12085,N_13741);
or UO_1488 (O_1488,N_14049,N_13984);
or UO_1489 (O_1489,N_13785,N_13507);
or UO_1490 (O_1490,N_13808,N_14355);
nor UO_1491 (O_1491,N_14915,N_14845);
nand UO_1492 (O_1492,N_13078,N_14124);
nand UO_1493 (O_1493,N_14761,N_12500);
or UO_1494 (O_1494,N_12536,N_14807);
and UO_1495 (O_1495,N_12274,N_14616);
and UO_1496 (O_1496,N_14743,N_12983);
or UO_1497 (O_1497,N_12547,N_13045);
nor UO_1498 (O_1498,N_14740,N_14133);
nor UO_1499 (O_1499,N_13973,N_14530);
nand UO_1500 (O_1500,N_14968,N_12224);
nand UO_1501 (O_1501,N_13689,N_13397);
or UO_1502 (O_1502,N_14337,N_12749);
nor UO_1503 (O_1503,N_13236,N_13050);
and UO_1504 (O_1504,N_13661,N_13513);
and UO_1505 (O_1505,N_13690,N_14958);
nand UO_1506 (O_1506,N_13824,N_13183);
or UO_1507 (O_1507,N_12178,N_14255);
nand UO_1508 (O_1508,N_12402,N_13006);
nor UO_1509 (O_1509,N_13771,N_14737);
and UO_1510 (O_1510,N_13293,N_13773);
or UO_1511 (O_1511,N_12767,N_13371);
or UO_1512 (O_1512,N_14699,N_14832);
and UO_1513 (O_1513,N_12643,N_13108);
nor UO_1514 (O_1514,N_14565,N_13340);
nor UO_1515 (O_1515,N_13650,N_13271);
or UO_1516 (O_1516,N_14770,N_14225);
nor UO_1517 (O_1517,N_12680,N_14041);
and UO_1518 (O_1518,N_12257,N_12264);
and UO_1519 (O_1519,N_12818,N_14129);
and UO_1520 (O_1520,N_12464,N_14830);
nor UO_1521 (O_1521,N_12998,N_14358);
or UO_1522 (O_1522,N_12132,N_12313);
nor UO_1523 (O_1523,N_12369,N_12575);
nand UO_1524 (O_1524,N_14181,N_12928);
nor UO_1525 (O_1525,N_12850,N_13256);
and UO_1526 (O_1526,N_12421,N_12339);
nor UO_1527 (O_1527,N_12960,N_14775);
nor UO_1528 (O_1528,N_13099,N_13608);
nor UO_1529 (O_1529,N_12303,N_12449);
nor UO_1530 (O_1530,N_12473,N_12683);
and UO_1531 (O_1531,N_14783,N_13216);
xnor UO_1532 (O_1532,N_14804,N_13074);
and UO_1533 (O_1533,N_14661,N_12327);
nor UO_1534 (O_1534,N_13461,N_12765);
nor UO_1535 (O_1535,N_14349,N_12784);
and UO_1536 (O_1536,N_14273,N_12298);
or UO_1537 (O_1537,N_14034,N_14760);
nor UO_1538 (O_1538,N_14380,N_13461);
or UO_1539 (O_1539,N_12117,N_14581);
or UO_1540 (O_1540,N_13167,N_12634);
and UO_1541 (O_1541,N_13512,N_13907);
nand UO_1542 (O_1542,N_13448,N_13311);
nand UO_1543 (O_1543,N_12684,N_14545);
nor UO_1544 (O_1544,N_13480,N_13997);
or UO_1545 (O_1545,N_14263,N_12829);
and UO_1546 (O_1546,N_14822,N_14740);
or UO_1547 (O_1547,N_13470,N_13703);
or UO_1548 (O_1548,N_12374,N_13937);
nor UO_1549 (O_1549,N_13994,N_13763);
and UO_1550 (O_1550,N_12245,N_14943);
nor UO_1551 (O_1551,N_12215,N_14083);
nor UO_1552 (O_1552,N_12508,N_14683);
nor UO_1553 (O_1553,N_14677,N_14937);
or UO_1554 (O_1554,N_12129,N_12014);
nor UO_1555 (O_1555,N_13966,N_12933);
nor UO_1556 (O_1556,N_13229,N_12913);
and UO_1557 (O_1557,N_13262,N_14336);
and UO_1558 (O_1558,N_14110,N_12775);
and UO_1559 (O_1559,N_13740,N_14251);
nand UO_1560 (O_1560,N_12650,N_14792);
and UO_1561 (O_1561,N_12066,N_14780);
nand UO_1562 (O_1562,N_14827,N_13576);
nand UO_1563 (O_1563,N_13371,N_12513);
nor UO_1564 (O_1564,N_13022,N_14743);
nand UO_1565 (O_1565,N_13242,N_13066);
xnor UO_1566 (O_1566,N_13660,N_12884);
and UO_1567 (O_1567,N_14386,N_12306);
and UO_1568 (O_1568,N_14638,N_14635);
nand UO_1569 (O_1569,N_12261,N_13776);
nand UO_1570 (O_1570,N_13376,N_14469);
or UO_1571 (O_1571,N_14588,N_12970);
nand UO_1572 (O_1572,N_13537,N_12511);
nand UO_1573 (O_1573,N_13537,N_12875);
and UO_1574 (O_1574,N_12937,N_12622);
or UO_1575 (O_1575,N_13865,N_13491);
or UO_1576 (O_1576,N_14826,N_14960);
and UO_1577 (O_1577,N_13339,N_13841);
or UO_1578 (O_1578,N_12632,N_12766);
nand UO_1579 (O_1579,N_14781,N_13464);
or UO_1580 (O_1580,N_13587,N_12137);
nand UO_1581 (O_1581,N_13902,N_14293);
nand UO_1582 (O_1582,N_12406,N_13548);
nand UO_1583 (O_1583,N_13424,N_13086);
xor UO_1584 (O_1584,N_13074,N_14381);
nand UO_1585 (O_1585,N_14260,N_13017);
nor UO_1586 (O_1586,N_13320,N_14491);
and UO_1587 (O_1587,N_14273,N_14485);
nand UO_1588 (O_1588,N_14510,N_14605);
nand UO_1589 (O_1589,N_13306,N_13013);
or UO_1590 (O_1590,N_14587,N_13844);
or UO_1591 (O_1591,N_14359,N_13424);
or UO_1592 (O_1592,N_14897,N_12303);
and UO_1593 (O_1593,N_13486,N_13072);
nand UO_1594 (O_1594,N_12782,N_13133);
or UO_1595 (O_1595,N_12620,N_14697);
xor UO_1596 (O_1596,N_13102,N_12175);
nor UO_1597 (O_1597,N_14607,N_12324);
nand UO_1598 (O_1598,N_12320,N_13246);
or UO_1599 (O_1599,N_14934,N_12799);
or UO_1600 (O_1600,N_13270,N_12715);
nor UO_1601 (O_1601,N_12846,N_14676);
and UO_1602 (O_1602,N_12100,N_14003);
or UO_1603 (O_1603,N_14935,N_14844);
nor UO_1604 (O_1604,N_14207,N_13278);
and UO_1605 (O_1605,N_12423,N_13674);
nand UO_1606 (O_1606,N_12192,N_14643);
xor UO_1607 (O_1607,N_13241,N_12437);
and UO_1608 (O_1608,N_14509,N_12871);
and UO_1609 (O_1609,N_12342,N_14560);
and UO_1610 (O_1610,N_12586,N_12544);
or UO_1611 (O_1611,N_14861,N_13739);
nand UO_1612 (O_1612,N_14451,N_14099);
nand UO_1613 (O_1613,N_14903,N_12755);
nor UO_1614 (O_1614,N_14676,N_13651);
or UO_1615 (O_1615,N_14422,N_13654);
and UO_1616 (O_1616,N_13203,N_14355);
and UO_1617 (O_1617,N_13041,N_14416);
nand UO_1618 (O_1618,N_12495,N_12226);
or UO_1619 (O_1619,N_12152,N_12188);
or UO_1620 (O_1620,N_12993,N_14258);
nor UO_1621 (O_1621,N_14366,N_14938);
nor UO_1622 (O_1622,N_12356,N_14194);
or UO_1623 (O_1623,N_14583,N_12205);
nor UO_1624 (O_1624,N_14067,N_12265);
nand UO_1625 (O_1625,N_14125,N_12370);
or UO_1626 (O_1626,N_14845,N_14072);
nand UO_1627 (O_1627,N_13501,N_14400);
or UO_1628 (O_1628,N_13825,N_12966);
or UO_1629 (O_1629,N_13498,N_14064);
and UO_1630 (O_1630,N_13113,N_14037);
nand UO_1631 (O_1631,N_14531,N_12887);
nor UO_1632 (O_1632,N_14641,N_14360);
and UO_1633 (O_1633,N_14989,N_14918);
nor UO_1634 (O_1634,N_14405,N_14143);
nor UO_1635 (O_1635,N_13850,N_12405);
or UO_1636 (O_1636,N_13628,N_14435);
or UO_1637 (O_1637,N_14182,N_14364);
nand UO_1638 (O_1638,N_12561,N_12572);
nand UO_1639 (O_1639,N_12214,N_14988);
or UO_1640 (O_1640,N_12654,N_12779);
nand UO_1641 (O_1641,N_12642,N_12211);
nor UO_1642 (O_1642,N_14170,N_14101);
xor UO_1643 (O_1643,N_12679,N_14463);
nand UO_1644 (O_1644,N_14460,N_13570);
nor UO_1645 (O_1645,N_12540,N_14326);
or UO_1646 (O_1646,N_12936,N_13559);
nor UO_1647 (O_1647,N_12679,N_13849);
nand UO_1648 (O_1648,N_13290,N_12475);
or UO_1649 (O_1649,N_12683,N_14420);
nor UO_1650 (O_1650,N_13590,N_12894);
nand UO_1651 (O_1651,N_13098,N_14019);
nor UO_1652 (O_1652,N_12012,N_14110);
nor UO_1653 (O_1653,N_13594,N_13307);
and UO_1654 (O_1654,N_13495,N_14917);
or UO_1655 (O_1655,N_13834,N_13365);
nand UO_1656 (O_1656,N_12701,N_13745);
xnor UO_1657 (O_1657,N_14384,N_13869);
and UO_1658 (O_1658,N_14754,N_12282);
and UO_1659 (O_1659,N_13143,N_12699);
or UO_1660 (O_1660,N_12985,N_13979);
and UO_1661 (O_1661,N_13113,N_14247);
and UO_1662 (O_1662,N_13880,N_13710);
or UO_1663 (O_1663,N_12869,N_12591);
nor UO_1664 (O_1664,N_12323,N_14813);
nor UO_1665 (O_1665,N_12125,N_12950);
and UO_1666 (O_1666,N_12348,N_12781);
nor UO_1667 (O_1667,N_13699,N_14267);
nor UO_1668 (O_1668,N_14408,N_13488);
xnor UO_1669 (O_1669,N_14556,N_14537);
or UO_1670 (O_1670,N_13335,N_14844);
nand UO_1671 (O_1671,N_13230,N_14475);
nand UO_1672 (O_1672,N_14786,N_14991);
nor UO_1673 (O_1673,N_12364,N_12503);
and UO_1674 (O_1674,N_13168,N_12275);
nand UO_1675 (O_1675,N_14123,N_12586);
nor UO_1676 (O_1676,N_12672,N_14666);
and UO_1677 (O_1677,N_12474,N_13842);
nor UO_1678 (O_1678,N_13285,N_13816);
nor UO_1679 (O_1679,N_13482,N_12555);
nor UO_1680 (O_1680,N_13125,N_13695);
nor UO_1681 (O_1681,N_14539,N_14892);
or UO_1682 (O_1682,N_14521,N_12617);
nand UO_1683 (O_1683,N_14390,N_12920);
nor UO_1684 (O_1684,N_13432,N_12727);
nor UO_1685 (O_1685,N_13741,N_14570);
nand UO_1686 (O_1686,N_14726,N_14387);
nor UO_1687 (O_1687,N_13614,N_13653);
and UO_1688 (O_1688,N_14825,N_14501);
and UO_1689 (O_1689,N_13431,N_12092);
or UO_1690 (O_1690,N_13020,N_13534);
nor UO_1691 (O_1691,N_14950,N_14351);
nor UO_1692 (O_1692,N_13970,N_12647);
nor UO_1693 (O_1693,N_13705,N_14407);
nand UO_1694 (O_1694,N_12274,N_13639);
and UO_1695 (O_1695,N_14119,N_14522);
nand UO_1696 (O_1696,N_13263,N_13023);
or UO_1697 (O_1697,N_13106,N_13843);
or UO_1698 (O_1698,N_12801,N_13552);
nor UO_1699 (O_1699,N_14296,N_14124);
nor UO_1700 (O_1700,N_14011,N_12991);
or UO_1701 (O_1701,N_13373,N_12322);
and UO_1702 (O_1702,N_12237,N_12671);
nor UO_1703 (O_1703,N_13908,N_13687);
xnor UO_1704 (O_1704,N_14902,N_12822);
or UO_1705 (O_1705,N_13581,N_13658);
nand UO_1706 (O_1706,N_14700,N_13043);
nor UO_1707 (O_1707,N_13701,N_12554);
and UO_1708 (O_1708,N_13061,N_12751);
and UO_1709 (O_1709,N_14814,N_12597);
or UO_1710 (O_1710,N_14261,N_12932);
and UO_1711 (O_1711,N_14575,N_13678);
or UO_1712 (O_1712,N_13714,N_12683);
or UO_1713 (O_1713,N_14300,N_13670);
and UO_1714 (O_1714,N_13380,N_12574);
or UO_1715 (O_1715,N_14611,N_12404);
or UO_1716 (O_1716,N_14687,N_14046);
nor UO_1717 (O_1717,N_13477,N_14807);
or UO_1718 (O_1718,N_14295,N_13244);
or UO_1719 (O_1719,N_13275,N_13558);
nand UO_1720 (O_1720,N_12910,N_14312);
nand UO_1721 (O_1721,N_14872,N_13291);
and UO_1722 (O_1722,N_12969,N_14818);
nand UO_1723 (O_1723,N_12376,N_13092);
nand UO_1724 (O_1724,N_12594,N_12118);
or UO_1725 (O_1725,N_13030,N_12503);
or UO_1726 (O_1726,N_12424,N_13678);
nand UO_1727 (O_1727,N_14669,N_12193);
and UO_1728 (O_1728,N_12265,N_14485);
nor UO_1729 (O_1729,N_12880,N_12183);
nand UO_1730 (O_1730,N_14172,N_12741);
or UO_1731 (O_1731,N_14149,N_13686);
and UO_1732 (O_1732,N_14233,N_12256);
or UO_1733 (O_1733,N_14953,N_12356);
and UO_1734 (O_1734,N_14083,N_14860);
nor UO_1735 (O_1735,N_13598,N_13463);
and UO_1736 (O_1736,N_14094,N_13464);
nor UO_1737 (O_1737,N_14145,N_13624);
and UO_1738 (O_1738,N_13402,N_13408);
and UO_1739 (O_1739,N_13479,N_12469);
or UO_1740 (O_1740,N_13591,N_13957);
nand UO_1741 (O_1741,N_14305,N_14716);
and UO_1742 (O_1742,N_12252,N_14911);
or UO_1743 (O_1743,N_12196,N_14559);
nor UO_1744 (O_1744,N_12988,N_14557);
nand UO_1745 (O_1745,N_13777,N_13013);
and UO_1746 (O_1746,N_13658,N_14905);
nand UO_1747 (O_1747,N_13859,N_14347);
nand UO_1748 (O_1748,N_14887,N_13930);
nand UO_1749 (O_1749,N_14832,N_13895);
nor UO_1750 (O_1750,N_14651,N_13372);
or UO_1751 (O_1751,N_12402,N_12416);
nor UO_1752 (O_1752,N_13783,N_13761);
or UO_1753 (O_1753,N_13466,N_14468);
or UO_1754 (O_1754,N_12347,N_14592);
and UO_1755 (O_1755,N_12679,N_13742);
or UO_1756 (O_1756,N_13389,N_14500);
nand UO_1757 (O_1757,N_12602,N_14760);
or UO_1758 (O_1758,N_12482,N_14711);
and UO_1759 (O_1759,N_13929,N_12651);
nor UO_1760 (O_1760,N_13328,N_12084);
or UO_1761 (O_1761,N_13862,N_13185);
xor UO_1762 (O_1762,N_13603,N_13723);
nand UO_1763 (O_1763,N_12295,N_12374);
nand UO_1764 (O_1764,N_14605,N_14665);
and UO_1765 (O_1765,N_13413,N_13416);
nand UO_1766 (O_1766,N_14509,N_13386);
nor UO_1767 (O_1767,N_13299,N_12971);
nor UO_1768 (O_1768,N_14501,N_12226);
nor UO_1769 (O_1769,N_14809,N_12821);
nor UO_1770 (O_1770,N_13897,N_12675);
nor UO_1771 (O_1771,N_14273,N_13523);
or UO_1772 (O_1772,N_13531,N_13250);
or UO_1773 (O_1773,N_13749,N_12794);
nand UO_1774 (O_1774,N_13455,N_13103);
nand UO_1775 (O_1775,N_12497,N_14401);
nand UO_1776 (O_1776,N_12418,N_12757);
or UO_1777 (O_1777,N_12445,N_14366);
nor UO_1778 (O_1778,N_13674,N_12376);
nor UO_1779 (O_1779,N_14099,N_13307);
or UO_1780 (O_1780,N_14047,N_12946);
nor UO_1781 (O_1781,N_14958,N_13377);
nand UO_1782 (O_1782,N_14574,N_13592);
or UO_1783 (O_1783,N_14647,N_13328);
nor UO_1784 (O_1784,N_13225,N_12900);
nor UO_1785 (O_1785,N_14390,N_13904);
or UO_1786 (O_1786,N_12006,N_12860);
and UO_1787 (O_1787,N_12542,N_14562);
nor UO_1788 (O_1788,N_13145,N_12038);
or UO_1789 (O_1789,N_14779,N_12942);
or UO_1790 (O_1790,N_13268,N_14384);
and UO_1791 (O_1791,N_14400,N_14691);
and UO_1792 (O_1792,N_13115,N_13633);
or UO_1793 (O_1793,N_12849,N_12241);
and UO_1794 (O_1794,N_13430,N_13917);
and UO_1795 (O_1795,N_14384,N_12931);
nand UO_1796 (O_1796,N_12279,N_14894);
and UO_1797 (O_1797,N_13977,N_12802);
nand UO_1798 (O_1798,N_13150,N_12620);
or UO_1799 (O_1799,N_13427,N_14149);
or UO_1800 (O_1800,N_13762,N_14487);
or UO_1801 (O_1801,N_13235,N_14575);
or UO_1802 (O_1802,N_12154,N_13532);
or UO_1803 (O_1803,N_13412,N_12311);
or UO_1804 (O_1804,N_14227,N_12773);
or UO_1805 (O_1805,N_12759,N_14326);
nor UO_1806 (O_1806,N_13473,N_14799);
and UO_1807 (O_1807,N_12494,N_12451);
nor UO_1808 (O_1808,N_12835,N_14290);
and UO_1809 (O_1809,N_14507,N_13000);
nand UO_1810 (O_1810,N_12908,N_14761);
nor UO_1811 (O_1811,N_12594,N_14642);
nor UO_1812 (O_1812,N_12070,N_14441);
nand UO_1813 (O_1813,N_14696,N_12808);
and UO_1814 (O_1814,N_14301,N_13302);
nand UO_1815 (O_1815,N_14783,N_13328);
nor UO_1816 (O_1816,N_12995,N_13232);
nand UO_1817 (O_1817,N_14052,N_12876);
nor UO_1818 (O_1818,N_14139,N_13472);
or UO_1819 (O_1819,N_12694,N_13200);
nor UO_1820 (O_1820,N_12954,N_13323);
nand UO_1821 (O_1821,N_14710,N_12880);
and UO_1822 (O_1822,N_12350,N_13886);
or UO_1823 (O_1823,N_13352,N_13598);
and UO_1824 (O_1824,N_12018,N_14084);
or UO_1825 (O_1825,N_14003,N_14255);
nand UO_1826 (O_1826,N_14304,N_12362);
or UO_1827 (O_1827,N_13080,N_12150);
nand UO_1828 (O_1828,N_14352,N_13046);
and UO_1829 (O_1829,N_13485,N_13992);
or UO_1830 (O_1830,N_14864,N_13667);
and UO_1831 (O_1831,N_12606,N_13518);
or UO_1832 (O_1832,N_13434,N_12438);
and UO_1833 (O_1833,N_14950,N_13636);
and UO_1834 (O_1834,N_13695,N_13173);
nand UO_1835 (O_1835,N_14764,N_13678);
or UO_1836 (O_1836,N_12945,N_12701);
or UO_1837 (O_1837,N_13964,N_12204);
and UO_1838 (O_1838,N_13534,N_12416);
and UO_1839 (O_1839,N_14325,N_13856);
nand UO_1840 (O_1840,N_12828,N_12772);
and UO_1841 (O_1841,N_14954,N_13709);
or UO_1842 (O_1842,N_12785,N_12904);
nand UO_1843 (O_1843,N_12973,N_12709);
nand UO_1844 (O_1844,N_14991,N_12841);
or UO_1845 (O_1845,N_14748,N_14430);
or UO_1846 (O_1846,N_13241,N_12263);
and UO_1847 (O_1847,N_13978,N_14059);
nor UO_1848 (O_1848,N_14311,N_13209);
and UO_1849 (O_1849,N_13432,N_13554);
or UO_1850 (O_1850,N_12659,N_14243);
or UO_1851 (O_1851,N_12387,N_12807);
and UO_1852 (O_1852,N_14017,N_12984);
and UO_1853 (O_1853,N_13147,N_13500);
nand UO_1854 (O_1854,N_13758,N_14928);
nand UO_1855 (O_1855,N_13693,N_13299);
nor UO_1856 (O_1856,N_13866,N_14515);
and UO_1857 (O_1857,N_12666,N_12855);
and UO_1858 (O_1858,N_12171,N_12666);
nand UO_1859 (O_1859,N_14223,N_12384);
or UO_1860 (O_1860,N_13994,N_13098);
or UO_1861 (O_1861,N_12422,N_13575);
or UO_1862 (O_1862,N_14032,N_13714);
and UO_1863 (O_1863,N_12252,N_14841);
and UO_1864 (O_1864,N_13649,N_12756);
and UO_1865 (O_1865,N_14841,N_13941);
or UO_1866 (O_1866,N_12592,N_12747);
nand UO_1867 (O_1867,N_13530,N_14451);
nand UO_1868 (O_1868,N_13683,N_12509);
or UO_1869 (O_1869,N_13620,N_14301);
and UO_1870 (O_1870,N_13966,N_14809);
nor UO_1871 (O_1871,N_14328,N_13375);
or UO_1872 (O_1872,N_12099,N_14891);
nand UO_1873 (O_1873,N_12675,N_13132);
or UO_1874 (O_1874,N_12368,N_13883);
nor UO_1875 (O_1875,N_13499,N_13847);
or UO_1876 (O_1876,N_12146,N_14426);
and UO_1877 (O_1877,N_13386,N_12985);
nor UO_1878 (O_1878,N_12991,N_14907);
nor UO_1879 (O_1879,N_13758,N_14971);
nor UO_1880 (O_1880,N_12869,N_14933);
and UO_1881 (O_1881,N_13540,N_13426);
nand UO_1882 (O_1882,N_14010,N_12559);
nand UO_1883 (O_1883,N_13664,N_14033);
nand UO_1884 (O_1884,N_14268,N_13371);
nor UO_1885 (O_1885,N_12261,N_14109);
nand UO_1886 (O_1886,N_13325,N_14279);
nand UO_1887 (O_1887,N_14169,N_13411);
and UO_1888 (O_1888,N_14767,N_14884);
or UO_1889 (O_1889,N_12765,N_12524);
nand UO_1890 (O_1890,N_12315,N_12195);
nand UO_1891 (O_1891,N_14298,N_14044);
xor UO_1892 (O_1892,N_13081,N_12960);
or UO_1893 (O_1893,N_13715,N_13821);
or UO_1894 (O_1894,N_14914,N_14515);
nand UO_1895 (O_1895,N_14195,N_14772);
nand UO_1896 (O_1896,N_12913,N_13785);
or UO_1897 (O_1897,N_14723,N_12717);
nor UO_1898 (O_1898,N_13022,N_14798);
nor UO_1899 (O_1899,N_13422,N_12929);
and UO_1900 (O_1900,N_12733,N_13874);
or UO_1901 (O_1901,N_13106,N_12059);
nand UO_1902 (O_1902,N_12355,N_12349);
or UO_1903 (O_1903,N_12922,N_14103);
and UO_1904 (O_1904,N_12525,N_12254);
and UO_1905 (O_1905,N_13751,N_12336);
or UO_1906 (O_1906,N_14156,N_12998);
and UO_1907 (O_1907,N_14567,N_14001);
or UO_1908 (O_1908,N_13337,N_14651);
and UO_1909 (O_1909,N_13926,N_12737);
nand UO_1910 (O_1910,N_14783,N_13947);
nor UO_1911 (O_1911,N_14842,N_13430);
nand UO_1912 (O_1912,N_12939,N_12081);
nand UO_1913 (O_1913,N_13037,N_12358);
or UO_1914 (O_1914,N_12773,N_14989);
nor UO_1915 (O_1915,N_12547,N_14028);
nand UO_1916 (O_1916,N_12266,N_14586);
nand UO_1917 (O_1917,N_14308,N_12603);
and UO_1918 (O_1918,N_14126,N_12098);
nor UO_1919 (O_1919,N_12827,N_14210);
nand UO_1920 (O_1920,N_12245,N_14411);
nor UO_1921 (O_1921,N_14624,N_12141);
nor UO_1922 (O_1922,N_13303,N_12292);
and UO_1923 (O_1923,N_12304,N_12601);
or UO_1924 (O_1924,N_12982,N_12588);
nor UO_1925 (O_1925,N_12874,N_14352);
nand UO_1926 (O_1926,N_14120,N_12500);
and UO_1927 (O_1927,N_12735,N_12179);
nand UO_1928 (O_1928,N_12544,N_12505);
or UO_1929 (O_1929,N_12597,N_13519);
or UO_1930 (O_1930,N_12675,N_13347);
and UO_1931 (O_1931,N_13743,N_14518);
and UO_1932 (O_1932,N_12052,N_14817);
nor UO_1933 (O_1933,N_14996,N_12619);
nand UO_1934 (O_1934,N_13339,N_14308);
nand UO_1935 (O_1935,N_13988,N_13195);
or UO_1936 (O_1936,N_14292,N_13887);
nor UO_1937 (O_1937,N_13834,N_12288);
or UO_1938 (O_1938,N_14525,N_14596);
or UO_1939 (O_1939,N_14261,N_13379);
and UO_1940 (O_1940,N_13612,N_12607);
and UO_1941 (O_1941,N_13422,N_13014);
nand UO_1942 (O_1942,N_13900,N_14870);
or UO_1943 (O_1943,N_14268,N_12619);
nand UO_1944 (O_1944,N_13875,N_13151);
nand UO_1945 (O_1945,N_14605,N_12122);
nand UO_1946 (O_1946,N_14479,N_13303);
or UO_1947 (O_1947,N_13630,N_13332);
and UO_1948 (O_1948,N_14023,N_13444);
or UO_1949 (O_1949,N_12035,N_14436);
nand UO_1950 (O_1950,N_13719,N_13123);
xnor UO_1951 (O_1951,N_14108,N_13505);
or UO_1952 (O_1952,N_13104,N_14174);
or UO_1953 (O_1953,N_13447,N_14984);
or UO_1954 (O_1954,N_13278,N_12150);
nor UO_1955 (O_1955,N_13469,N_14065);
or UO_1956 (O_1956,N_14342,N_14344);
and UO_1957 (O_1957,N_14738,N_13440);
and UO_1958 (O_1958,N_14756,N_13794);
nand UO_1959 (O_1959,N_13758,N_14157);
nand UO_1960 (O_1960,N_14584,N_14927);
nand UO_1961 (O_1961,N_13116,N_13821);
or UO_1962 (O_1962,N_12123,N_12426);
or UO_1963 (O_1963,N_13935,N_12575);
nor UO_1964 (O_1964,N_13526,N_13737);
and UO_1965 (O_1965,N_13406,N_12011);
and UO_1966 (O_1966,N_13640,N_12061);
or UO_1967 (O_1967,N_13406,N_13766);
and UO_1968 (O_1968,N_13658,N_13278);
nor UO_1969 (O_1969,N_13106,N_12663);
or UO_1970 (O_1970,N_12139,N_14390);
nand UO_1971 (O_1971,N_12974,N_13973);
or UO_1972 (O_1972,N_12579,N_14709);
nand UO_1973 (O_1973,N_14810,N_12141);
or UO_1974 (O_1974,N_12513,N_12254);
nand UO_1975 (O_1975,N_13630,N_13337);
nand UO_1976 (O_1976,N_14286,N_12055);
nor UO_1977 (O_1977,N_14219,N_14471);
nor UO_1978 (O_1978,N_13517,N_14612);
nor UO_1979 (O_1979,N_12350,N_12145);
nor UO_1980 (O_1980,N_12769,N_13627);
and UO_1981 (O_1981,N_13836,N_13839);
nand UO_1982 (O_1982,N_13282,N_13012);
nor UO_1983 (O_1983,N_13932,N_14248);
nand UO_1984 (O_1984,N_12149,N_12866);
nand UO_1985 (O_1985,N_14232,N_13334);
and UO_1986 (O_1986,N_12673,N_12730);
or UO_1987 (O_1987,N_14498,N_12893);
or UO_1988 (O_1988,N_12673,N_13454);
and UO_1989 (O_1989,N_13710,N_13613);
and UO_1990 (O_1990,N_12891,N_13884);
or UO_1991 (O_1991,N_14737,N_13390);
nand UO_1992 (O_1992,N_13757,N_12204);
nor UO_1993 (O_1993,N_12874,N_12792);
nor UO_1994 (O_1994,N_14688,N_13680);
nand UO_1995 (O_1995,N_12146,N_14234);
or UO_1996 (O_1996,N_13020,N_14767);
nor UO_1997 (O_1997,N_12555,N_14137);
and UO_1998 (O_1998,N_13185,N_14446);
and UO_1999 (O_1999,N_13104,N_13592);
endmodule