module basic_2500_25000_3000_8_levels_10xor_3(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999;
or U0 (N_0,In_1758,In_1764);
xnor U1 (N_1,In_565,In_1237);
xnor U2 (N_2,In_2461,In_722);
xnor U3 (N_3,In_801,In_422);
or U4 (N_4,In_1609,In_2449);
or U5 (N_5,In_1083,In_1020);
and U6 (N_6,In_1577,In_1504);
nor U7 (N_7,In_1870,In_2391);
xnor U8 (N_8,In_151,In_2473);
nand U9 (N_9,In_1395,In_517);
nand U10 (N_10,In_1131,In_1709);
xnor U11 (N_11,In_655,In_351);
and U12 (N_12,In_83,In_1613);
nor U13 (N_13,In_222,In_1645);
or U14 (N_14,In_1800,In_2260);
xnor U15 (N_15,In_1972,In_1897);
or U16 (N_16,In_2059,In_868);
or U17 (N_17,In_343,In_1430);
xor U18 (N_18,In_2344,In_39);
nor U19 (N_19,In_496,In_587);
or U20 (N_20,In_1635,In_695);
xnor U21 (N_21,In_2167,In_1572);
nand U22 (N_22,In_1673,In_2380);
or U23 (N_23,In_1832,In_1655);
and U24 (N_24,In_1871,In_2371);
nand U25 (N_25,In_2427,In_683);
or U26 (N_26,In_1711,In_440);
nor U27 (N_27,In_2193,In_1601);
xor U28 (N_28,In_844,In_2441);
xor U29 (N_29,In_955,In_312);
nor U30 (N_30,In_84,In_945);
xor U31 (N_31,In_956,In_1850);
xor U32 (N_32,In_1428,In_2030);
nor U33 (N_33,In_2021,In_1337);
nor U34 (N_34,In_1630,In_598);
nand U35 (N_35,In_1167,In_898);
or U36 (N_36,In_597,In_368);
and U37 (N_37,In_247,In_981);
nand U38 (N_38,In_1819,In_145);
nand U39 (N_39,In_917,In_2336);
and U40 (N_40,In_2346,In_1688);
nor U41 (N_41,In_309,In_1029);
and U42 (N_42,In_2240,In_2335);
nor U43 (N_43,In_1436,In_1672);
and U44 (N_44,In_1461,In_1889);
and U45 (N_45,In_2278,In_111);
or U46 (N_46,In_1175,In_458);
and U47 (N_47,In_553,In_761);
nand U48 (N_48,In_822,In_676);
nor U49 (N_49,In_2482,In_206);
or U50 (N_50,In_1761,In_2175);
nor U51 (N_51,In_1702,In_168);
nor U52 (N_52,In_578,In_279);
nand U53 (N_53,In_2189,In_1420);
xor U54 (N_54,In_1248,In_1352);
nand U55 (N_55,In_803,In_2141);
nand U56 (N_56,In_1391,In_256);
nor U57 (N_57,In_1447,In_2154);
nor U58 (N_58,In_1334,In_905);
xnor U59 (N_59,In_393,In_1346);
nor U60 (N_60,In_2147,In_1778);
xor U61 (N_61,In_2173,In_18);
nand U62 (N_62,In_1340,In_735);
xor U63 (N_63,In_1802,In_1);
xnor U64 (N_64,In_102,In_194);
nand U65 (N_65,In_1591,In_1215);
or U66 (N_66,In_1139,In_1569);
or U67 (N_67,In_579,In_1474);
and U68 (N_68,In_437,In_2137);
xnor U69 (N_69,In_1914,In_1234);
xnor U70 (N_70,In_2050,In_324);
nor U71 (N_71,In_1470,In_1756);
and U72 (N_72,In_3,In_1306);
and U73 (N_73,In_472,In_402);
or U74 (N_74,In_133,In_2263);
and U75 (N_75,In_1358,In_1922);
and U76 (N_76,In_1226,In_1230);
and U77 (N_77,In_2166,In_1479);
xor U78 (N_78,In_1191,In_130);
or U79 (N_79,In_120,In_1534);
xor U80 (N_80,In_2426,In_1085);
and U81 (N_81,In_667,In_662);
and U82 (N_82,In_119,In_2311);
or U83 (N_83,In_1211,In_2010);
nor U84 (N_84,In_221,In_2304);
nand U85 (N_85,In_1032,In_1098);
and U86 (N_86,In_1909,In_2483);
nor U87 (N_87,In_1462,In_240);
nand U88 (N_88,In_2377,In_1665);
nor U89 (N_89,In_1882,In_382);
and U90 (N_90,In_1667,In_937);
xor U91 (N_91,In_1294,In_428);
xnor U92 (N_92,In_1633,In_1296);
nand U93 (N_93,In_337,In_977);
nand U94 (N_94,In_1573,In_2396);
nand U95 (N_95,In_2381,In_1855);
and U96 (N_96,In_786,In_180);
or U97 (N_97,In_962,In_1096);
or U98 (N_98,In_2325,In_1051);
and U99 (N_99,In_74,In_816);
nor U100 (N_100,In_1349,In_314);
xor U101 (N_101,In_1152,In_892);
or U102 (N_102,In_227,In_1729);
nor U103 (N_103,In_336,In_327);
nand U104 (N_104,In_535,In_2215);
or U105 (N_105,In_2216,In_310);
and U106 (N_106,In_1977,In_1606);
nand U107 (N_107,In_620,In_27);
or U108 (N_108,In_1045,In_1144);
nor U109 (N_109,In_277,In_1901);
nor U110 (N_110,In_1722,In_56);
xnor U111 (N_111,In_1176,In_1915);
or U112 (N_112,In_2289,In_1203);
xor U113 (N_113,In_518,In_1811);
and U114 (N_114,In_1654,In_853);
nor U115 (N_115,In_797,In_665);
xnor U116 (N_116,In_13,In_1799);
or U117 (N_117,In_751,In_2379);
nor U118 (N_118,In_1787,In_295);
xnor U119 (N_119,In_2080,In_452);
and U120 (N_120,In_2122,In_420);
and U121 (N_121,In_1442,In_497);
or U122 (N_122,In_1602,In_2169);
nand U123 (N_123,In_2355,In_454);
and U124 (N_124,In_2358,In_873);
xor U125 (N_125,In_457,In_1755);
nor U126 (N_126,In_1035,In_1603);
nand U127 (N_127,In_2227,In_413);
nand U128 (N_128,In_2094,In_1331);
xor U129 (N_129,In_1836,In_2290);
or U130 (N_130,In_320,In_747);
xor U131 (N_131,In_2228,In_1412);
or U132 (N_132,In_1537,In_41);
or U133 (N_133,In_547,In_1379);
or U134 (N_134,In_1285,In_1048);
xor U135 (N_135,In_1245,In_2284);
and U136 (N_136,In_16,In_1851);
or U137 (N_137,In_651,In_1734);
nand U138 (N_138,In_1720,In_1130);
nor U139 (N_139,In_1402,In_765);
xnor U140 (N_140,In_2019,In_1934);
and U141 (N_141,In_213,In_2012);
xor U142 (N_142,In_1797,In_2330);
or U143 (N_143,In_1015,In_795);
and U144 (N_144,In_1894,In_411);
nor U145 (N_145,In_1413,In_789);
xnor U146 (N_146,In_19,In_170);
xor U147 (N_147,In_2130,In_303);
nor U148 (N_148,In_901,In_1794);
nor U149 (N_149,In_2034,In_2083);
nand U150 (N_150,In_608,In_1718);
and U151 (N_151,In_273,In_34);
nand U152 (N_152,In_1730,In_2115);
nand U153 (N_153,In_1699,In_2339);
and U154 (N_154,In_2170,In_628);
or U155 (N_155,In_2451,In_1313);
xor U156 (N_156,In_1372,In_763);
and U157 (N_157,In_467,In_1344);
xnor U158 (N_158,In_2453,In_2383);
and U159 (N_159,In_1866,In_2282);
nor U160 (N_160,In_1375,In_1565);
and U161 (N_161,In_2053,In_1993);
nand U162 (N_162,In_776,In_825);
xor U163 (N_163,In_2084,In_131);
nand U164 (N_164,In_2331,In_1779);
and U165 (N_165,In_1124,In_686);
nand U166 (N_166,In_289,In_882);
nor U167 (N_167,In_1437,In_2245);
and U168 (N_168,In_160,In_1692);
xnor U169 (N_169,In_2002,In_72);
or U170 (N_170,In_669,In_904);
nand U171 (N_171,In_1243,In_2210);
and U172 (N_172,In_2418,In_571);
nand U173 (N_173,In_2131,In_1286);
or U174 (N_174,In_1184,In_1129);
or U175 (N_175,In_921,In_2196);
nand U176 (N_176,In_1959,In_1874);
nand U177 (N_177,In_401,In_970);
xor U178 (N_178,In_1445,In_1450);
nor U179 (N_179,In_2499,In_828);
and U180 (N_180,In_895,In_191);
xor U181 (N_181,In_2270,In_2265);
and U182 (N_182,In_788,In_899);
xnor U183 (N_183,In_1491,In_2160);
nor U184 (N_184,In_2203,In_643);
and U185 (N_185,In_610,In_967);
nand U186 (N_186,In_2042,In_135);
and U187 (N_187,In_400,In_2001);
nand U188 (N_188,In_2433,In_1626);
nor U189 (N_189,In_1345,In_1305);
xnor U190 (N_190,In_2490,In_1468);
nand U191 (N_191,In_217,In_1276);
nand U192 (N_192,In_95,In_348);
nor U193 (N_193,In_2026,In_491);
xor U194 (N_194,In_1656,In_1596);
or U195 (N_195,In_1653,In_1679);
xnor U196 (N_196,In_614,In_434);
and U197 (N_197,In_1624,In_2345);
xnor U198 (N_198,In_724,In_1055);
and U199 (N_199,In_926,In_1767);
nor U200 (N_200,In_304,In_1456);
and U201 (N_201,In_1947,In_1806);
nor U202 (N_202,In_2123,In_1488);
nand U203 (N_203,In_1762,In_511);
nor U204 (N_204,In_2231,In_1001);
or U205 (N_205,In_1765,In_1381);
nand U206 (N_206,In_582,In_1900);
nor U207 (N_207,In_648,In_2457);
xnor U208 (N_208,In_177,In_2187);
nand U209 (N_209,In_1424,In_2370);
or U210 (N_210,In_684,In_605);
xor U211 (N_211,In_2181,In_826);
or U212 (N_212,In_592,In_1684);
or U213 (N_213,In_1404,In_1531);
xor U214 (N_214,In_2182,In_2204);
and U215 (N_215,In_1731,In_2314);
nand U216 (N_216,In_2129,In_1365);
xor U217 (N_217,In_1440,In_617);
and U218 (N_218,In_451,In_1739);
or U219 (N_219,In_299,In_373);
xor U220 (N_220,In_798,In_595);
nor U221 (N_221,In_306,In_2120);
nand U222 (N_222,In_1223,In_1078);
or U223 (N_223,In_819,In_2388);
and U224 (N_224,In_2430,In_1747);
xnor U225 (N_225,In_68,In_680);
or U226 (N_226,In_737,In_2484);
and U227 (N_227,In_297,In_378);
nor U228 (N_228,In_1007,In_2243);
xor U229 (N_229,In_1677,In_1273);
nor U230 (N_230,In_950,In_70);
and U231 (N_231,In_1817,In_1100);
nand U232 (N_232,In_2485,In_2403);
xor U233 (N_233,In_1809,In_510);
nor U234 (N_234,In_2163,In_2017);
and U235 (N_235,In_81,In_1022);
and U236 (N_236,In_2274,In_2275);
and U237 (N_237,In_1043,In_644);
nor U238 (N_238,In_1054,In_252);
nand U239 (N_239,In_563,In_1760);
nand U240 (N_240,In_1198,In_1540);
nor U241 (N_241,In_857,In_647);
nor U242 (N_242,In_673,In_840);
xnor U243 (N_243,In_118,In_1733);
nor U244 (N_244,In_2423,In_1695);
nand U245 (N_245,In_1042,In_415);
nand U246 (N_246,In_1978,In_2277);
xnor U247 (N_247,In_1328,In_2271);
and U248 (N_248,In_2164,In_228);
and U249 (N_249,In_558,In_1693);
and U250 (N_250,In_784,In_2434);
nor U251 (N_251,In_507,In_66);
nor U252 (N_252,In_1158,In_633);
or U253 (N_253,In_2224,In_762);
nor U254 (N_254,In_2481,In_2238);
and U255 (N_255,In_1946,In_1342);
and U256 (N_256,In_1524,In_2234);
nor U257 (N_257,In_865,In_2410);
nor U258 (N_258,In_2027,In_2152);
xor U259 (N_259,In_2319,In_909);
or U260 (N_260,In_1843,In_626);
xor U261 (N_261,In_1103,In_1782);
or U262 (N_262,In_696,In_1608);
nor U263 (N_263,In_1427,In_697);
and U264 (N_264,In_1827,In_1005);
and U265 (N_265,In_1854,In_802);
xnor U266 (N_266,In_1526,In_739);
xor U267 (N_267,In_2471,In_2014);
nand U268 (N_268,In_494,In_906);
xnor U269 (N_269,In_530,In_2202);
nor U270 (N_270,In_1196,In_77);
or U271 (N_271,In_1881,In_1320);
nor U272 (N_272,In_2463,In_2250);
nor U273 (N_273,In_1156,In_1019);
and U274 (N_274,In_1807,In_1600);
xnor U275 (N_275,In_1954,In_1724);
xor U276 (N_276,In_2397,In_1357);
or U277 (N_277,In_2015,In_1539);
nand U278 (N_278,In_1324,In_1682);
nand U279 (N_279,In_144,In_65);
nor U280 (N_280,In_782,In_2249);
and U281 (N_281,In_2322,In_448);
xnor U282 (N_282,In_1683,In_2393);
xnor U283 (N_283,In_2348,In_1240);
nand U284 (N_284,In_716,In_2256);
nor U285 (N_285,In_1271,In_968);
xnor U286 (N_286,In_2267,In_2382);
and U287 (N_287,In_1091,In_1239);
and U288 (N_288,In_288,In_860);
nand U289 (N_289,In_1443,In_1457);
nand U290 (N_290,In_1251,In_710);
nor U291 (N_291,In_1114,In_276);
and U292 (N_292,In_1815,In_55);
or U293 (N_293,In_2088,In_1578);
and U294 (N_294,In_108,In_2413);
nand U295 (N_295,In_874,In_640);
or U296 (N_296,In_999,In_278);
xnor U297 (N_297,In_1314,In_1986);
nand U298 (N_298,In_2352,In_934);
xor U299 (N_299,In_636,In_978);
and U300 (N_300,In_2007,In_158);
or U301 (N_301,In_199,In_1181);
and U302 (N_302,In_728,In_2035);
and U303 (N_303,In_2436,In_1745);
xnor U304 (N_304,In_1199,In_1566);
or U305 (N_305,In_1587,In_830);
or U306 (N_306,In_1192,In_1581);
nand U307 (N_307,In_263,In_1502);
nor U308 (N_308,In_1771,In_426);
nand U309 (N_309,In_2031,In_359);
and U310 (N_310,In_224,In_1991);
nand U311 (N_311,In_1675,In_2389);
nor U312 (N_312,In_560,In_1725);
and U313 (N_313,In_1805,In_1140);
nor U314 (N_314,In_539,In_780);
nand U315 (N_315,In_2110,In_1970);
xnor U316 (N_316,In_1902,In_886);
nand U317 (N_317,In_984,In_1589);
nor U318 (N_318,In_685,In_30);
xor U319 (N_319,In_2168,In_1723);
xor U320 (N_320,In_1023,In_664);
and U321 (N_321,In_1218,In_759);
nor U322 (N_322,In_1736,In_2048);
nand U323 (N_323,In_1863,In_61);
and U324 (N_324,In_62,In_1047);
nor U325 (N_325,In_1607,In_340);
nor U326 (N_326,In_1967,In_2401);
xor U327 (N_327,In_701,In_1172);
xor U328 (N_328,In_1353,In_202);
or U329 (N_329,In_1485,In_2272);
nand U330 (N_330,In_1859,In_1829);
and U331 (N_331,In_2340,In_2113);
nor U332 (N_332,In_646,In_2404);
or U333 (N_333,In_2440,In_281);
nor U334 (N_334,In_867,In_1400);
and U335 (N_335,In_1757,In_714);
or U336 (N_336,In_1965,In_637);
nand U337 (N_337,In_345,In_972);
nor U338 (N_338,In_2004,In_1772);
nand U339 (N_339,In_769,In_2038);
nor U340 (N_340,In_1280,In_2237);
or U341 (N_341,In_155,In_2140);
and U342 (N_342,In_961,In_1403);
or U343 (N_343,In_33,In_1551);
or U344 (N_344,In_1503,In_2065);
or U345 (N_345,In_98,In_2420);
nor U346 (N_346,In_1750,In_671);
nand U347 (N_347,In_933,In_848);
and U348 (N_348,In_76,In_1107);
or U349 (N_349,In_2468,In_2387);
nand U350 (N_350,In_556,In_2261);
xor U351 (N_351,In_2063,In_2324);
and U352 (N_352,In_2241,In_187);
and U353 (N_353,In_1522,In_2054);
nor U354 (N_354,In_588,In_1516);
or U355 (N_355,In_835,In_1744);
and U356 (N_356,In_139,In_2142);
nand U357 (N_357,In_1017,In_1363);
nor U358 (N_358,In_1826,In_89);
nor U359 (N_359,In_1561,In_150);
or U360 (N_360,In_2206,In_2003);
xnor U361 (N_361,In_1792,In_2244);
nand U362 (N_362,In_715,In_1359);
or U363 (N_363,In_196,In_1721);
or U364 (N_364,In_25,In_1899);
and U365 (N_365,In_302,In_1640);
nor U366 (N_366,In_441,In_301);
or U367 (N_367,In_1134,In_522);
or U368 (N_368,In_1360,In_2354);
nor U369 (N_369,In_1707,In_391);
and U370 (N_370,In_35,In_1006);
and U371 (N_371,In_2096,In_635);
and U372 (N_372,In_1303,In_707);
xor U373 (N_373,In_1691,In_2158);
or U374 (N_374,In_814,In_2246);
nand U375 (N_375,In_1696,In_1170);
and U376 (N_376,In_894,In_1451);
and U377 (N_377,In_1932,In_501);
xnor U378 (N_378,In_533,In_371);
nor U379 (N_379,In_1669,In_1680);
and U380 (N_380,In_653,In_757);
and U381 (N_381,In_2363,In_1030);
and U382 (N_382,In_2104,In_167);
nand U383 (N_383,In_1579,In_741);
nor U384 (N_384,In_2006,In_1446);
and U385 (N_385,In_1997,In_137);
xor U386 (N_386,In_425,In_1620);
and U387 (N_387,In_1396,In_210);
and U388 (N_388,In_1664,In_2082);
xnor U389 (N_389,In_123,In_1458);
or U390 (N_390,In_1088,In_675);
nor U391 (N_391,In_14,In_607);
or U392 (N_392,In_2293,In_1728);
xor U393 (N_393,In_201,In_2195);
xor U394 (N_394,In_8,In_36);
and U395 (N_395,In_1279,In_358);
nand U396 (N_396,In_1368,In_2254);
xnor U397 (N_397,In_2108,In_534);
xor U398 (N_398,In_1037,In_980);
or U399 (N_399,In_75,In_63);
nor U400 (N_400,In_418,In_296);
and U401 (N_401,In_212,In_1935);
nor U402 (N_402,In_758,In_1299);
or U403 (N_403,In_513,In_23);
xnor U404 (N_404,In_1394,In_1418);
nand U405 (N_405,In_1868,In_1873);
xor U406 (N_406,In_1186,In_1482);
or U407 (N_407,In_220,In_2298);
or U408 (N_408,In_1890,In_1956);
and U409 (N_409,In_2091,In_2302);
nor U410 (N_410,In_586,In_1763);
and U411 (N_411,In_1949,In_1117);
and U412 (N_412,In_1486,In_260);
nand U413 (N_413,In_2125,In_328);
xor U414 (N_414,In_271,In_1647);
nand U415 (N_415,In_113,In_2255);
nor U416 (N_416,In_1676,In_880);
xnor U417 (N_417,In_1464,In_1382);
nor U418 (N_418,In_1657,In_2116);
nand U419 (N_419,In_604,In_2446);
or U420 (N_420,In_1149,In_2315);
nand U421 (N_421,In_2497,In_1962);
or U422 (N_422,In_1270,In_568);
and U423 (N_423,In_1109,In_1634);
nor U424 (N_424,In_2185,In_2155);
or U425 (N_425,In_2151,In_430);
nand U426 (N_426,In_185,In_1594);
nand U427 (N_427,In_613,In_912);
nand U428 (N_428,In_2459,In_1431);
or U429 (N_429,In_1735,In_632);
and U430 (N_430,In_1580,In_1530);
nor U431 (N_431,In_785,In_845);
nor U432 (N_432,In_923,In_723);
nand U433 (N_433,In_2087,In_544);
nor U434 (N_434,In_421,In_1077);
nor U435 (N_435,In_564,In_2341);
xor U436 (N_436,In_733,In_1104);
nor U437 (N_437,In_1238,In_2398);
and U438 (N_438,In_1097,In_1236);
nor U439 (N_439,In_2157,In_2013);
or U440 (N_440,In_1974,In_96);
and U441 (N_441,In_708,In_363);
xnor U442 (N_442,In_1080,In_813);
and U443 (N_443,In_1495,In_954);
nor U444 (N_444,In_2402,In_1060);
nor U445 (N_445,In_639,In_2144);
xnor U446 (N_446,In_1904,In_251);
nor U447 (N_447,In_79,In_521);
or U448 (N_448,In_1034,In_367);
nand U449 (N_449,In_1411,In_162);
nand U450 (N_450,In_1810,In_1518);
nand U451 (N_451,In_520,In_2068);
xor U452 (N_452,In_1912,In_2297);
and U453 (N_453,In_2374,In_85);
xnor U454 (N_454,In_877,In_1075);
nor U455 (N_455,In_270,In_1574);
nand U456 (N_456,In_603,In_2495);
and U457 (N_457,In_2089,In_1074);
xnor U458 (N_458,In_1081,In_460);
nor U459 (N_459,In_456,In_1089);
or U460 (N_460,In_584,In_2476);
nand U461 (N_461,In_1769,In_1940);
xor U462 (N_462,In_858,In_2036);
nand U463 (N_463,In_576,In_862);
xnor U464 (N_464,In_1062,In_1113);
xnor U465 (N_465,In_1259,In_1708);
nor U466 (N_466,In_734,In_660);
xor U467 (N_467,In_837,In_172);
nand U468 (N_468,In_488,In_2056);
nor U469 (N_469,In_1025,In_2121);
xor U470 (N_470,In_2496,In_2086);
and U471 (N_471,In_1189,In_1801);
or U472 (N_472,In_807,In_104);
xnor U473 (N_473,In_1247,In_670);
or U474 (N_474,In_1244,In_188);
nand U475 (N_475,In_129,In_342);
xnor U476 (N_476,In_2266,In_864);
or U477 (N_477,In_285,In_709);
and U478 (N_478,In_1862,In_2342);
xor U479 (N_479,In_700,In_1738);
nor U480 (N_480,In_2074,In_1204);
xor U481 (N_481,In_1924,In_127);
xor U482 (N_482,In_1166,In_2111);
nand U483 (N_483,In_1713,In_1715);
and U484 (N_484,In_2070,In_1714);
or U485 (N_485,In_1785,In_939);
xnor U486 (N_486,In_52,In_919);
or U487 (N_487,In_1876,In_1793);
xor U488 (N_488,In_2409,In_1347);
nor U489 (N_489,In_887,In_1498);
xnor U490 (N_490,In_1028,In_993);
or U491 (N_491,In_2448,In_1849);
or U492 (N_492,In_1490,In_107);
xnor U493 (N_493,In_1466,In_2055);
and U494 (N_494,In_1858,In_717);
nor U495 (N_495,In_775,In_2317);
or U496 (N_496,In_743,In_1880);
and U497 (N_497,In_1407,In_204);
or U498 (N_498,In_122,In_376);
nand U499 (N_499,In_2022,In_1329);
xnor U500 (N_500,In_768,In_1508);
nor U501 (N_501,In_1842,In_2498);
xnor U502 (N_502,In_627,In_712);
or U503 (N_503,In_1895,In_115);
nand U504 (N_504,In_1183,In_1241);
xor U505 (N_505,In_112,In_753);
or U506 (N_506,In_100,In_190);
nor U507 (N_507,In_1312,In_2361);
nand U508 (N_508,In_2360,In_856);
and U509 (N_509,In_1825,In_504);
xnor U510 (N_510,In_1092,In_1926);
xnor U511 (N_511,In_793,In_136);
nand U512 (N_512,In_1681,In_506);
nor U513 (N_513,In_891,In_1388);
xor U514 (N_514,In_1687,In_1333);
and U515 (N_515,In_668,In_2437);
xnor U516 (N_516,In_2332,In_609);
and U517 (N_517,In_1153,In_31);
or U518 (N_518,In_152,In_834);
xor U519 (N_519,In_752,In_1289);
xnor U520 (N_520,In_1629,In_2207);
xor U521 (N_521,In_9,In_731);
nand U522 (N_522,In_2474,In_106);
nor U523 (N_523,In_1541,In_2323);
xor U524 (N_524,In_2259,In_1533);
nand U525 (N_525,In_738,In_1076);
xnor U526 (N_526,In_1136,In_2309);
and U527 (N_527,In_53,In_979);
nor U528 (N_528,In_1093,In_2286);
xor U529 (N_529,In_169,In_964);
xor U530 (N_530,In_408,In_1930);
xnor U531 (N_531,In_1105,In_963);
and U532 (N_532,In_2394,In_1497);
or U533 (N_533,In_1275,In_445);
nand U534 (N_534,In_580,In_965);
nand U535 (N_535,In_2146,In_1698);
and U536 (N_536,In_935,In_1867);
nand U537 (N_537,In_760,In_2225);
nor U538 (N_538,In_1435,In_259);
nor U539 (N_539,In_287,In_889);
xor U540 (N_540,In_91,In_879);
nor U541 (N_541,In_207,In_2180);
nand U542 (N_542,In_661,In_1976);
nor U543 (N_543,In_1291,In_799);
or U544 (N_544,In_2222,In_142);
nand U545 (N_545,In_267,In_1383);
nor U546 (N_546,In_1258,In_2431);
nor U547 (N_547,In_1187,In_897);
or U548 (N_548,In_2092,In_1548);
xor U549 (N_549,In_2177,In_985);
nand U550 (N_550,In_90,In_1178);
nand U551 (N_551,In_1550,In_2321);
nor U552 (N_552,In_2062,In_1410);
or U553 (N_553,In_57,In_1386);
nor U554 (N_554,In_357,In_313);
xnor U555 (N_555,In_2310,In_621);
or U556 (N_556,In_975,In_1896);
xor U557 (N_557,In_1101,In_2090);
nand U558 (N_558,In_1128,In_69);
nor U559 (N_559,In_516,In_1401);
nor U560 (N_560,In_1951,In_951);
and U561 (N_561,In_1549,In_1478);
xnor U562 (N_562,In_827,In_1563);
xnor U563 (N_563,In_941,In_2174);
nor U564 (N_564,In_146,In_1072);
xnor U565 (N_565,In_156,In_2051);
or U566 (N_566,In_2269,In_2390);
and U567 (N_567,In_907,In_2183);
and U568 (N_568,In_7,In_602);
xnor U569 (N_569,In_1473,In_773);
and U570 (N_570,In_2287,In_1616);
or U571 (N_571,In_1250,In_2029);
xor U572 (N_572,In_255,In_1833);
nor U573 (N_573,In_149,In_1119);
or U574 (N_574,In_2165,In_248);
or U575 (N_575,In_361,In_1952);
nor U576 (N_576,In_1791,In_1197);
nand U577 (N_577,In_1919,In_1126);
nand U578 (N_578,In_232,In_2220);
or U579 (N_579,In_164,In_1666);
and U580 (N_580,In_1472,In_1348);
or U581 (N_581,In_1903,In_1505);
xor U582 (N_582,In_2467,In_1267);
nand U583 (N_583,In_2201,In_1063);
xnor U584 (N_584,In_2159,In_932);
xnor U585 (N_585,In_5,In_101);
nand U586 (N_586,In_659,In_1169);
nor U587 (N_587,In_1837,In_1228);
and U588 (N_588,In_15,In_2456);
nor U589 (N_589,In_766,In_2306);
nor U590 (N_590,In_1011,In_927);
or U591 (N_591,In_2205,In_1040);
nor U592 (N_592,In_1564,In_1878);
nand U593 (N_593,In_1844,In_1393);
nand U594 (N_594,In_2452,In_410);
nand U595 (N_595,In_754,In_550);
nor U596 (N_596,In_464,In_184);
xor U597 (N_597,In_353,In_729);
or U598 (N_598,In_1036,In_1148);
and U599 (N_599,In_332,In_815);
or U600 (N_600,In_679,In_1031);
nand U601 (N_601,In_1309,In_1282);
xor U602 (N_602,In_1283,In_960);
or U603 (N_603,In_2258,In_480);
nor U604 (N_604,In_1527,In_1409);
and U605 (N_605,In_424,In_2044);
or U606 (N_606,In_638,In_334);
nor U607 (N_607,In_1749,In_2079);
and U608 (N_608,In_2049,In_1038);
xnor U609 (N_609,In_1082,In_2356);
xnor U610 (N_610,In_1067,In_721);
nand U611 (N_611,In_976,In_268);
or U612 (N_612,In_503,In_1115);
xnor U613 (N_613,In_615,In_974);
and U614 (N_614,In_931,In_1803);
xnor U615 (N_615,In_2276,In_1775);
or U616 (N_616,In_1253,In_869);
and U617 (N_617,In_1016,In_1483);
nand U618 (N_618,In_1918,In_2313);
nor U619 (N_619,In_1726,In_475);
or U620 (N_620,In_2248,In_515);
nand U621 (N_621,In_274,In_269);
or U622 (N_622,In_1262,In_1532);
and U623 (N_623,In_1597,In_525);
or U624 (N_624,In_377,In_258);
and U625 (N_625,In_1071,In_616);
nand U626 (N_626,In_554,In_861);
nand U627 (N_627,In_138,In_1557);
nor U628 (N_628,In_1086,In_2488);
nor U629 (N_629,In_1448,In_2232);
xor U630 (N_630,In_1496,In_2303);
nand U631 (N_631,In_349,In_1911);
nand U632 (N_632,In_246,In_1828);
and U633 (N_633,In_1399,In_311);
nand U634 (N_634,In_1717,In_1116);
xnor U635 (N_635,In_2218,In_1392);
nand U636 (N_636,In_2136,In_1585);
nand U637 (N_637,In_126,In_2307);
nor U638 (N_638,In_2296,In_284);
nor U639 (N_639,In_1122,In_1719);
or U640 (N_640,In_1773,In_1231);
nand U641 (N_641,In_1517,In_2188);
nand U642 (N_642,In_462,In_1453);
xnor U643 (N_643,In_1795,In_2107);
nand U644 (N_644,In_957,In_1936);
nand U645 (N_645,In_1958,In_1233);
or U646 (N_646,In_1026,In_344);
or U647 (N_647,In_2000,In_2235);
nor U648 (N_648,In_1180,In_2127);
nor U649 (N_649,In_1642,In_756);
xnor U650 (N_650,In_1018,In_1087);
nor U651 (N_651,In_1905,In_2494);
and U652 (N_652,In_1257,In_2285);
xor U653 (N_653,In_1658,In_208);
xnor U654 (N_654,In_1678,In_315);
and U655 (N_655,In_552,In_1406);
nand U656 (N_656,In_1390,In_1944);
and U657 (N_657,In_1263,In_2073);
or U658 (N_658,In_1157,In_1553);
xor U659 (N_659,In_47,In_186);
nand U660 (N_660,In_567,In_2209);
nand U661 (N_661,In_2411,In_1293);
nand U662 (N_662,In_2291,In_1766);
or U663 (N_663,In_2172,In_409);
xnor U664 (N_664,In_755,In_42);
nor U665 (N_665,In_404,In_1370);
or U666 (N_666,In_971,In_322);
nor U667 (N_667,In_374,In_1511);
nor U668 (N_668,In_1214,In_529);
and U669 (N_669,In_774,In_1434);
and U670 (N_670,In_677,In_1983);
nand U671 (N_671,In_989,In_2262);
xor U672 (N_672,In_1605,In_347);
nor U673 (N_673,In_1408,In_817);
and U674 (N_674,In_654,In_2133);
and U675 (N_675,In_1592,In_1992);
and U676 (N_676,In_116,In_1741);
xnor U677 (N_677,In_1351,In_2333);
nor U678 (N_678,In_1552,In_2095);
nor U679 (N_679,In_82,In_611);
and U680 (N_680,In_1099,In_1307);
nor U681 (N_681,In_2138,In_778);
and U682 (N_682,In_742,In_2162);
or U683 (N_683,In_555,In_2493);
nor U684 (N_684,In_470,In_1892);
and U685 (N_685,In_244,In_966);
nor U686 (N_686,In_720,In_1477);
nand U687 (N_687,In_385,In_183);
or U688 (N_688,In_2008,In_1910);
and U689 (N_689,In_1266,In_1740);
nor U690 (N_690,In_2114,In_688);
and U691 (N_691,In_1260,In_1102);
nand U692 (N_692,In_631,In_173);
and U693 (N_693,In_1604,In_117);
xnor U694 (N_694,In_2465,In_2406);
or U695 (N_695,In_1599,In_2033);
xnor U696 (N_696,In_1480,In_2489);
xnor U697 (N_697,In_1513,In_22);
and U698 (N_698,In_1012,In_262);
nor U699 (N_699,In_403,In_2040);
and U700 (N_700,In_1120,In_1225);
nor U701 (N_701,In_215,In_2462);
nor U702 (N_702,In_2472,In_1421);
nand U703 (N_703,In_1917,In_2045);
xor U704 (N_704,In_711,In_2149);
and U705 (N_705,In_45,In_1056);
or U706 (N_706,In_1948,In_450);
and U707 (N_707,In_1162,In_2150);
xnor U708 (N_708,In_405,In_1308);
nand U709 (N_709,In_1830,In_1737);
or U710 (N_710,In_839,In_652);
nor U711 (N_711,In_1582,In_2226);
and U712 (N_712,In_2349,In_1746);
nand U713 (N_713,In_852,In_478);
and U714 (N_714,In_2052,In_996);
or U715 (N_715,In_562,In_211);
xor U716 (N_716,In_2194,In_1341);
nand U717 (N_717,In_1476,In_1510);
xor U718 (N_718,In_1638,In_1321);
or U719 (N_719,In_1628,In_831);
xor U720 (N_720,In_1290,In_1145);
or U721 (N_721,In_719,In_1188);
and U722 (N_722,In_692,In_809);
nor U723 (N_723,In_1027,In_2320);
and U724 (N_724,In_2435,In_986);
or U725 (N_725,In_1110,In_1998);
and U726 (N_726,In_1378,In_226);
and U727 (N_727,In_1242,In_1697);
nor U728 (N_728,In_1950,In_2105);
xor U729 (N_729,In_1405,In_1945);
or U730 (N_730,In_189,In_338);
nand U731 (N_731,In_257,In_2305);
nor U732 (N_732,In_940,In_6);
and U733 (N_733,In_678,In_1615);
and U734 (N_734,In_1786,In_1506);
or U735 (N_735,In_952,In_1219);
nand U736 (N_736,In_463,In_854);
nand U737 (N_737,In_706,In_1990);
or U738 (N_738,In_1452,In_911);
or U739 (N_739,In_2148,In_1942);
nor U740 (N_740,In_1033,In_71);
or U741 (N_741,In_219,In_1254);
or U742 (N_742,In_988,In_2061);
xor U743 (N_743,In_205,In_1493);
nor U744 (N_744,In_481,In_147);
and U745 (N_745,In_2212,In_21);
or U746 (N_746,In_1367,In_1222);
xor U747 (N_747,In_1535,In_1908);
nor U748 (N_748,In_1643,In_2190);
nand U749 (N_749,In_447,In_2386);
nor U750 (N_750,In_423,In_1179);
nor U751 (N_751,In_1487,In_878);
nor U752 (N_752,In_674,In_1095);
xnor U753 (N_753,In_849,In_589);
nor U754 (N_754,In_1514,In_2373);
or U755 (N_755,In_265,In_1332);
and U756 (N_756,In_2392,In_157);
nand U757 (N_757,In_1920,In_1155);
nand U758 (N_758,In_490,In_820);
or U759 (N_759,In_335,In_58);
or U760 (N_760,In_872,In_165);
or U761 (N_761,In_1860,In_1570);
nor U762 (N_762,In_1748,In_159);
xor U763 (N_763,In_319,In_1710);
nand U764 (N_764,In_2171,In_166);
or U765 (N_765,In_379,In_2491);
and U766 (N_766,In_1700,In_1053);
and U767 (N_767,In_1789,In_1065);
and U768 (N_768,In_380,In_1509);
or U769 (N_769,In_1875,In_1938);
nor U770 (N_770,In_705,In_1512);
nand U771 (N_771,In_1742,In_1142);
xnor U772 (N_772,In_1287,In_1112);
nand U773 (N_773,In_471,In_1907);
nand U774 (N_774,In_1925,In_1070);
or U775 (N_775,In_241,In_1439);
nor U776 (N_776,In_1323,In_953);
xnor U777 (N_777,In_339,In_2312);
or U778 (N_778,In_499,In_1220);
and U779 (N_779,In_704,In_2071);
or U780 (N_780,In_1499,In_1554);
xnor U781 (N_781,In_537,In_855);
and U782 (N_782,In_2251,In_2428);
nor U783 (N_783,In_439,In_1834);
or U784 (N_784,In_540,In_1884);
and U785 (N_785,In_687,In_298);
and U786 (N_786,In_233,In_0);
and U787 (N_787,In_2334,In_2458);
or U788 (N_788,In_2362,In_1190);
xnor U789 (N_789,In_859,In_2058);
or U790 (N_790,In_969,In_573);
and U791 (N_791,In_2421,In_1988);
nor U792 (N_792,In_1467,In_740);
nor U793 (N_793,In_787,In_1614);
and U794 (N_794,In_198,In_767);
xnor U795 (N_795,In_1193,In_1235);
xnor U796 (N_796,In_1143,In_2124);
nor U797 (N_797,In_1090,In_1355);
or U798 (N_798,In_67,In_2217);
or U799 (N_799,In_1460,In_482);
xor U800 (N_800,In_1753,In_1135);
or U801 (N_801,In_2128,In_1471);
or U802 (N_802,In_477,In_1743);
and U803 (N_803,In_1160,In_1229);
nor U804 (N_804,In_197,In_1373);
xor U805 (N_805,In_280,In_699);
and U806 (N_806,In_1955,In_1292);
nor U807 (N_807,In_1545,In_1611);
and U808 (N_808,In_1438,In_804);
xnor U809 (N_809,In_60,In_1132);
or U810 (N_810,In_235,In_1674);
xor U811 (N_811,In_292,In_2064);
or U812 (N_812,In_148,In_908);
or U813 (N_813,In_948,In_333);
and U814 (N_814,In_1371,In_2078);
nand U815 (N_815,In_703,In_1975);
and U816 (N_816,In_1732,In_469);
xor U817 (N_817,In_2415,In_38);
xnor U818 (N_818,In_792,In_991);
xor U819 (N_819,In_618,In_2432);
nor U820 (N_820,In_174,In_736);
nor U821 (N_821,In_959,In_2);
nor U822 (N_822,In_997,In_230);
xnor U823 (N_823,In_1891,In_307);
and U824 (N_824,In_557,In_1376);
or U825 (N_825,In_468,In_1576);
or U826 (N_826,In_1350,In_1841);
nand U827 (N_827,In_1584,In_2318);
or U828 (N_828,In_200,In_548);
nand U829 (N_829,In_2300,In_983);
or U830 (N_830,In_1221,In_26);
or U831 (N_831,In_924,In_86);
nand U832 (N_832,In_1252,In_1455);
or U833 (N_833,In_1694,In_1963);
nor U834 (N_834,In_583,In_561);
xor U835 (N_835,In_1780,In_888);
or U836 (N_836,In_161,In_50);
nor U837 (N_837,In_2455,In_1893);
xor U838 (N_838,In_1979,In_245);
and U839 (N_839,In_1861,In_811);
xnor U840 (N_840,In_2365,In_681);
nand U841 (N_841,In_1644,In_253);
xor U842 (N_842,In_316,In_1432);
nand U843 (N_843,In_1706,In_225);
nor U844 (N_844,In_730,In_641);
and U845 (N_845,In_432,In_1426);
or U846 (N_846,In_1519,In_78);
nor U847 (N_847,In_843,In_1856);
and U848 (N_848,In_2252,In_153);
xor U849 (N_849,In_1982,In_1449);
and U850 (N_850,In_2347,In_2037);
nand U851 (N_851,In_1325,In_326);
nor U852 (N_852,In_486,In_375);
and U853 (N_853,In_1507,In_390);
and U854 (N_854,In_163,In_360);
or U855 (N_855,In_1014,In_2257);
or U856 (N_856,In_2242,In_1300);
nand U857 (N_857,In_1840,In_2076);
xnor U858 (N_858,In_1173,In_1433);
xor U859 (N_859,In_914,In_1212);
or U860 (N_860,In_2109,In_1898);
xor U861 (N_861,In_435,In_622);
nor U862 (N_862,In_356,In_1610);
and U863 (N_863,In_2081,In_2378);
or U864 (N_864,In_625,In_2097);
or U865 (N_865,In_195,In_2041);
or U866 (N_866,In_594,In_1354);
nor U867 (N_867,In_1168,In_1877);
xnor U868 (N_868,In_2425,In_443);
nor U869 (N_869,In_1796,In_2283);
nand U870 (N_870,In_493,In_829);
or U871 (N_871,In_2134,In_179);
xnor U872 (N_872,In_523,In_1598);
or U873 (N_873,In_1317,In_203);
nor U874 (N_874,In_1906,In_1668);
nor U875 (N_875,In_1374,In_841);
nand U876 (N_876,In_2301,In_1009);
nor U877 (N_877,In_370,In_1398);
nor U878 (N_878,In_1278,In_1073);
or U879 (N_879,In_691,In_1777);
nor U880 (N_880,In_2400,In_431);
and U881 (N_881,In_125,In_1704);
nor U882 (N_882,In_2414,In_43);
xor U883 (N_883,In_399,In_2279);
nor U884 (N_884,In_702,In_1649);
or U885 (N_885,In_871,In_663);
or U886 (N_886,In_1058,In_805);
nor U887 (N_887,In_1937,In_466);
xor U888 (N_888,In_1319,In_890);
nor U889 (N_889,In_17,In_512);
and U890 (N_890,In_690,In_1525);
and U891 (N_891,In_1567,In_1246);
nand U892 (N_892,In_396,In_1397);
and U893 (N_893,In_796,In_214);
and U894 (N_894,In_1049,In_870);
and U895 (N_895,In_1685,In_2020);
or U896 (N_896,In_243,In_2117);
or U897 (N_897,In_291,In_538);
and U898 (N_898,In_1923,In_87);
or U899 (N_899,In_2178,In_254);
and U900 (N_900,In_1586,In_250);
or U901 (N_901,In_474,In_325);
nand U902 (N_902,In_593,In_1364);
nor U903 (N_903,In_2419,In_1820);
and U904 (N_904,In_110,In_944);
nor U905 (N_905,In_1641,In_2197);
nand U906 (N_906,In_601,In_836);
and U907 (N_907,In_417,In_1444);
nand U908 (N_908,In_1297,In_1010);
nand U909 (N_909,In_1185,In_1121);
or U910 (N_910,In_2447,In_1489);
and U911 (N_911,In_581,In_2214);
and U912 (N_912,In_505,In_2395);
nor U913 (N_913,In_2417,In_656);
xnor U914 (N_914,In_2445,In_929);
xnor U915 (N_915,In_1465,In_1205);
and U916 (N_916,In_2408,In_1652);
and U917 (N_917,In_290,In_2039);
nor U918 (N_918,In_2253,In_294);
nor U919 (N_919,In_2364,In_1546);
nor U920 (N_920,In_2191,In_4);
or U921 (N_921,In_2099,In_1916);
or U922 (N_922,In_1933,In_175);
and U923 (N_923,In_851,In_1454);
nor U924 (N_924,In_1627,In_1384);
and U925 (N_925,In_1475,In_223);
or U926 (N_926,In_1052,In_1659);
xnor U927 (N_927,In_808,In_750);
xnor U928 (N_928,In_1969,In_444);
or U929 (N_929,In_2264,In_305);
nor U930 (N_930,In_1064,In_987);
nor U931 (N_931,In_1759,In_577);
or U932 (N_932,In_93,In_181);
or U933 (N_933,In_1318,In_99);
nand U934 (N_934,In_1768,In_1865);
xor U935 (N_935,In_2139,In_1301);
or U936 (N_936,In_794,In_1492);
xor U937 (N_937,In_317,In_1500);
or U938 (N_938,In_1147,In_1118);
nand U939 (N_939,In_600,In_2156);
xor U940 (N_940,In_29,In_489);
or U941 (N_941,In_1165,In_727);
and U942 (N_942,In_1387,In_2486);
xor U943 (N_943,In_2229,In_657);
xnor U944 (N_944,In_1798,In_1928);
nand U945 (N_945,In_381,In_1159);
xor U946 (N_946,In_2469,In_2211);
nor U947 (N_947,In_389,In_2057);
nand U948 (N_948,In_218,In_1835);
or U949 (N_949,In_1003,In_1057);
and U950 (N_950,In_994,In_479);
or U951 (N_951,In_746,In_1989);
and U952 (N_952,In_876,In_772);
nor U953 (N_953,In_487,In_73);
nor U954 (N_954,In_2359,In_2230);
xnor U955 (N_955,In_1133,In_943);
xor U956 (N_956,In_427,In_355);
xor U957 (N_957,In_569,In_2085);
xor U958 (N_958,In_103,In_2025);
and U959 (N_959,In_543,In_216);
and U960 (N_960,In_1316,In_1264);
nand U961 (N_961,In_623,In_745);
nand U962 (N_962,In_823,In_485);
or U963 (N_963,In_2308,In_2069);
or U964 (N_964,In_1913,In_1163);
nor U965 (N_965,In_526,In_1636);
xnor U966 (N_966,In_1154,In_1138);
nand U967 (N_967,In_1703,In_713);
and U968 (N_968,In_2233,In_1712);
nand U969 (N_969,In_1024,In_1061);
or U970 (N_970,In_1068,In_2376);
nor U971 (N_971,In_1417,In_1151);
and U972 (N_972,In_930,In_1562);
or U973 (N_973,In_1622,In_777);
xor U974 (N_974,In_1966,In_672);
and U975 (N_975,In_881,In_275);
or U976 (N_976,In_958,In_449);
xor U977 (N_977,In_1869,In_1174);
nor U978 (N_978,In_2422,In_1380);
xor U979 (N_979,In_599,In_1879);
xor U980 (N_980,In_1808,In_2075);
nor U981 (N_981,In_321,In_2464);
nand U982 (N_982,In_238,In_1927);
xnor U983 (N_983,In_2438,In_1021);
nand U984 (N_984,In_920,In_154);
and U985 (N_985,In_1853,In_1568);
xor U986 (N_986,In_1823,In_1008);
nand U987 (N_987,In_114,In_2337);
nand U988 (N_988,In_1377,In_838);
or U989 (N_989,In_893,In_846);
and U990 (N_990,In_2442,In_483);
nor U991 (N_991,In_236,In_764);
nor U992 (N_992,In_1217,In_1845);
or U993 (N_993,In_1754,In_1249);
xnor U994 (N_994,In_412,In_885);
nor U995 (N_995,In_416,In_1150);
or U996 (N_996,In_1846,In_946);
nand U997 (N_997,In_2219,In_134);
nand U998 (N_998,In_1984,In_476);
nor U999 (N_999,In_1816,In_771);
or U1000 (N_1000,In_1004,In_790);
xor U1001 (N_1001,In_1651,In_1315);
and U1002 (N_1002,In_810,In_936);
xnor U1003 (N_1003,In_407,In_11);
nor U1004 (N_1004,In_1961,In_2375);
and U1005 (N_1005,In_566,In_694);
or U1006 (N_1006,In_1814,In_2454);
nand U1007 (N_1007,In_1547,In_2024);
or U1008 (N_1008,In_2385,In_397);
and U1009 (N_1009,In_645,In_1481);
or U1010 (N_1010,In_141,In_973);
or U1011 (N_1011,In_97,In_1662);
and U1012 (N_1012,In_1423,In_2475);
and U1013 (N_1013,In_884,In_1330);
or U1014 (N_1014,In_2100,In_1069);
nor U1015 (N_1015,In_1752,In_171);
nor U1016 (N_1016,In_330,In_2199);
and U1017 (N_1017,In_1575,In_1171);
or U1018 (N_1018,In_2236,In_387);
xnor U1019 (N_1019,In_2366,In_619);
xnor U1020 (N_1020,In_2161,In_1194);
or U1021 (N_1021,In_1705,In_2368);
or U1022 (N_1022,In_947,In_1690);
xor U1023 (N_1023,In_352,In_1559);
or U1024 (N_1024,In_630,In_105);
and U1025 (N_1025,In_918,In_2112);
xnor U1026 (N_1026,In_2072,In_2213);
or U1027 (N_1027,In_1084,In_1288);
nor U1028 (N_1028,In_1277,In_2186);
and U1029 (N_1029,In_1361,In_922);
or U1030 (N_1030,In_2018,In_1528);
nor U1031 (N_1031,In_1041,In_1994);
nor U1032 (N_1032,In_2009,In_2119);
nor U1033 (N_1033,In_1195,In_1885);
and U1034 (N_1034,In_1123,In_1177);
xnor U1035 (N_1035,In_536,In_1788);
xnor U1036 (N_1036,In_1716,In_2338);
or U1037 (N_1037,In_1646,In_2153);
xor U1038 (N_1038,In_398,In_1232);
and U1039 (N_1039,In_1872,In_1216);
and U1040 (N_1040,In_1311,In_473);
or U1041 (N_1041,In_1971,In_1414);
and U1042 (N_1042,In_1106,In_2046);
or U1043 (N_1043,In_866,In_1625);
or U1044 (N_1044,In_49,In_575);
or U1045 (N_1045,In_546,In_1921);
nor U1046 (N_1046,In_1689,In_833);
and U1047 (N_1047,In_266,In_1366);
nor U1048 (N_1048,In_509,In_354);
nor U1049 (N_1049,In_1425,In_1059);
xnor U1050 (N_1050,In_1941,In_779);
or U1051 (N_1051,In_1108,In_1207);
and U1052 (N_1052,In_392,In_732);
or U1053 (N_1053,In_2060,In_541);
or U1054 (N_1054,In_770,In_239);
nor U1055 (N_1055,In_524,In_2176);
nor U1056 (N_1056,In_386,In_438);
nand U1057 (N_1057,In_1542,In_2032);
nor U1058 (N_1058,In_1339,In_2143);
and U1059 (N_1059,In_748,In_698);
or U1060 (N_1060,In_44,In_1650);
nor U1061 (N_1061,In_1957,In_143);
and U1062 (N_1062,In_590,In_624);
nor U1063 (N_1063,In_433,In_92);
or U1064 (N_1064,In_1558,In_1939);
nand U1065 (N_1065,In_1821,In_942);
or U1066 (N_1066,In_394,In_346);
or U1067 (N_1067,In_928,In_237);
and U1068 (N_1068,In_1310,In_800);
xor U1069 (N_1069,In_725,In_1046);
nand U1070 (N_1070,In_2316,In_508);
nand U1071 (N_1071,In_2405,In_1501);
nand U1072 (N_1072,In_1864,In_2328);
nor U1073 (N_1073,In_1623,In_916);
or U1074 (N_1074,In_40,In_1094);
and U1075 (N_1075,In_64,In_2118);
nor U1076 (N_1076,In_1544,In_1304);
xnor U1077 (N_1077,In_689,In_2295);
nor U1078 (N_1078,In_446,In_2479);
nand U1079 (N_1079,In_1776,In_37);
nand U1080 (N_1080,In_229,In_1039);
and U1081 (N_1081,In_128,In_572);
and U1082 (N_1082,In_818,In_1343);
or U1083 (N_1083,In_1987,In_492);
and U1084 (N_1084,In_1838,In_1079);
and U1085 (N_1085,In_384,In_1818);
nand U1086 (N_1086,In_1770,In_1000);
nand U1087 (N_1087,In_925,In_1201);
xor U1088 (N_1088,In_1617,In_2443);
and U1089 (N_1089,In_2135,In_2416);
nand U1090 (N_1090,In_124,In_498);
and U1091 (N_1091,In_2047,In_1822);
or U1092 (N_1092,In_1556,In_806);
and U1093 (N_1093,In_821,In_234);
nor U1094 (N_1094,In_2350,In_121);
or U1095 (N_1095,In_1050,In_1686);
nor U1096 (N_1096,In_182,In_383);
and U1097 (N_1097,In_1415,In_2439);
nand U1098 (N_1098,In_2280,In_1463);
and U1099 (N_1099,In_2288,In_1648);
xnor U1100 (N_1100,In_2028,In_2093);
xnor U1101 (N_1101,In_1044,In_2067);
and U1102 (N_1102,In_1981,In_2239);
xnor U1103 (N_1103,In_1125,In_1336);
nor U1104 (N_1104,In_1416,In_2329);
and U1105 (N_1105,In_1284,In_455);
nor U1106 (N_1106,In_2221,In_178);
and U1107 (N_1107,In_242,In_559);
xor U1108 (N_1108,In_2066,In_1161);
or U1109 (N_1109,In_1385,In_1389);
and U1110 (N_1110,In_249,In_995);
xor U1111 (N_1111,In_372,In_2184);
xor U1112 (N_1112,In_32,In_992);
xnor U1113 (N_1113,In_1663,In_551);
and U1114 (N_1114,In_51,In_1326);
nor U1115 (N_1115,In_2327,In_1202);
xor U1116 (N_1116,In_545,In_1631);
nor U1117 (N_1117,In_272,In_902);
nand U1118 (N_1118,In_1621,In_88);
and U1119 (N_1119,In_1960,In_1999);
xor U1120 (N_1120,In_1298,In_1583);
or U1121 (N_1121,In_1356,In_2179);
or U1122 (N_1122,In_48,In_1595);
or U1123 (N_1123,In_2208,In_442);
or U1124 (N_1124,In_329,In_1670);
xor U1125 (N_1125,In_1338,In_2273);
or U1126 (N_1126,In_140,In_1887);
nor U1127 (N_1127,In_2103,In_2077);
or U1128 (N_1128,In_193,In_591);
xnor U1129 (N_1129,In_1784,In_2247);
and U1130 (N_1130,In_1268,In_2005);
or U1131 (N_1131,In_1781,In_1459);
nor U1132 (N_1132,In_2292,In_1127);
xor U1133 (N_1133,In_1852,In_461);
nor U1134 (N_1134,In_791,In_453);
xor U1135 (N_1135,In_364,In_863);
nand U1136 (N_1136,In_2477,In_1612);
nand U1137 (N_1137,In_2098,In_1210);
and U1138 (N_1138,In_484,In_658);
nand U1139 (N_1139,In_94,In_1943);
nor U1140 (N_1140,In_1980,In_331);
nor U1141 (N_1141,In_2126,In_1295);
nand U1142 (N_1142,In_500,In_495);
or U1143 (N_1143,In_2043,In_1265);
or U1144 (N_1144,In_1327,In_2367);
nand U1145 (N_1145,In_2351,In_24);
nand U1146 (N_1146,In_596,In_12);
xnor U1147 (N_1147,In_1929,In_1521);
and U1148 (N_1148,In_1529,In_59);
nand U1149 (N_1149,In_990,In_2198);
nand U1150 (N_1150,In_1515,In_350);
and U1151 (N_1151,In_1281,In_842);
or U1152 (N_1152,In_2478,In_1206);
and U1153 (N_1153,In_2223,In_1520);
xnor U1154 (N_1154,In_847,In_2294);
nand U1155 (N_1155,In_1931,In_1639);
and U1156 (N_1156,In_1632,In_1783);
nor U1157 (N_1157,In_1182,In_1269);
or U1158 (N_1158,In_1227,In_406);
and U1159 (N_1159,In_726,In_938);
and U1160 (N_1160,In_2399,In_1774);
xor U1161 (N_1161,In_650,In_910);
or U1162 (N_1162,In_2450,In_900);
nor U1163 (N_1163,In_419,In_465);
xor U1164 (N_1164,In_781,In_1619);
or U1165 (N_1165,In_666,In_1888);
nand U1166 (N_1166,In_286,In_2132);
and U1167 (N_1167,In_2192,In_2412);
xor U1168 (N_1168,In_1274,In_1973);
nor U1169 (N_1169,In_1335,In_46);
and U1170 (N_1170,In_2357,In_1571);
nand U1171 (N_1171,In_1419,In_2480);
nand U1172 (N_1172,In_896,In_1804);
nor U1173 (N_1173,In_812,In_1111);
xnor U1174 (N_1174,In_2268,In_1369);
or U1175 (N_1175,In_1200,In_2016);
nand U1176 (N_1176,In_1701,In_2384);
xnor U1177 (N_1177,In_1146,In_365);
nor U1178 (N_1178,In_915,In_2011);
nand U1179 (N_1179,In_80,In_1813);
nor U1180 (N_1180,In_2326,In_414);
nor U1181 (N_1181,In_282,In_209);
and U1182 (N_1182,In_1256,In_528);
or U1183 (N_1183,In_2343,In_1671);
xor U1184 (N_1184,In_1002,In_850);
or U1185 (N_1185,In_1164,In_1362);
and U1186 (N_1186,In_2281,In_824);
nand U1187 (N_1187,In_532,In_388);
or U1188 (N_1188,In_264,In_531);
and U1189 (N_1189,In_2353,In_283);
and U1190 (N_1190,In_2101,In_1847);
nand U1191 (N_1191,In_2407,In_2299);
xor U1192 (N_1192,In_1523,In_132);
nor U1193 (N_1193,In_1886,In_261);
nand U1194 (N_1194,In_2372,In_832);
or U1195 (N_1195,In_718,In_459);
nor U1196 (N_1196,In_1790,In_629);
nand U1197 (N_1197,In_744,In_341);
xnor U1198 (N_1198,In_1964,In_2023);
or U1199 (N_1199,In_1995,In_913);
or U1200 (N_1200,In_1538,In_570);
nand U1201 (N_1201,In_542,In_1429);
nor U1202 (N_1202,In_949,In_2102);
nand U1203 (N_1203,In_54,In_519);
or U1204 (N_1204,In_1013,In_28);
and U1205 (N_1205,In_1484,In_1261);
nand U1206 (N_1206,In_682,In_634);
xnor U1207 (N_1207,In_2369,In_308);
and U1208 (N_1208,In_2470,In_982);
nand U1209 (N_1209,In_436,In_642);
xnor U1210 (N_1210,In_300,In_293);
or U1211 (N_1211,In_1661,In_1560);
nor U1212 (N_1212,In_1751,In_1824);
xor U1213 (N_1213,In_1224,In_1588);
xor U1214 (N_1214,In_1141,In_2145);
nand U1215 (N_1215,In_649,In_585);
xnor U1216 (N_1216,In_1590,In_1272);
xor U1217 (N_1217,In_1209,In_2200);
xnor U1218 (N_1218,In_231,In_693);
xnor U1219 (N_1219,In_176,In_1302);
and U1220 (N_1220,In_1727,In_1831);
nor U1221 (N_1221,In_1839,In_875);
or U1222 (N_1222,In_1322,In_2466);
and U1223 (N_1223,In_1968,In_749);
and U1224 (N_1224,In_323,In_606);
nor U1225 (N_1225,In_783,In_1208);
and U1226 (N_1226,In_1422,In_1066);
nor U1227 (N_1227,In_527,In_366);
or U1228 (N_1228,In_1441,In_1213);
xnor U1229 (N_1229,In_2444,In_1137);
nor U1230 (N_1230,In_2487,In_369);
xor U1231 (N_1231,In_549,In_362);
nor U1232 (N_1232,In_1660,In_1618);
or U1233 (N_1233,In_903,In_1883);
nor U1234 (N_1234,In_1812,In_883);
nor U1235 (N_1235,In_1494,In_318);
nor U1236 (N_1236,In_2429,In_998);
and U1237 (N_1237,In_2424,In_612);
or U1238 (N_1238,In_20,In_192);
and U1239 (N_1239,In_2492,In_1469);
xnor U1240 (N_1240,In_1857,In_502);
and U1241 (N_1241,In_1985,In_2106);
nand U1242 (N_1242,In_1996,In_1543);
xor U1243 (N_1243,In_1555,In_1637);
nand U1244 (N_1244,In_1536,In_574);
nor U1245 (N_1245,In_395,In_1953);
nand U1246 (N_1246,In_429,In_109);
and U1247 (N_1247,In_1255,In_1593);
or U1248 (N_1248,In_514,In_1848);
nor U1249 (N_1249,In_2460,In_10);
nand U1250 (N_1250,In_1132,In_1017);
nor U1251 (N_1251,In_381,In_810);
or U1252 (N_1252,In_2286,In_882);
or U1253 (N_1253,In_2337,In_2356);
xor U1254 (N_1254,In_1065,In_49);
xnor U1255 (N_1255,In_530,In_276);
or U1256 (N_1256,In_1844,In_1648);
nand U1257 (N_1257,In_1608,In_770);
nand U1258 (N_1258,In_1724,In_1008);
and U1259 (N_1259,In_972,In_2089);
nor U1260 (N_1260,In_452,In_1890);
and U1261 (N_1261,In_426,In_2297);
nand U1262 (N_1262,In_1932,In_500);
and U1263 (N_1263,In_1526,In_1360);
and U1264 (N_1264,In_13,In_1425);
and U1265 (N_1265,In_623,In_6);
nand U1266 (N_1266,In_2430,In_1005);
xnor U1267 (N_1267,In_438,In_1103);
nor U1268 (N_1268,In_76,In_1239);
nand U1269 (N_1269,In_270,In_2492);
nand U1270 (N_1270,In_824,In_737);
nor U1271 (N_1271,In_1598,In_1359);
nor U1272 (N_1272,In_819,In_1422);
and U1273 (N_1273,In_2100,In_99);
or U1274 (N_1274,In_2219,In_2309);
and U1275 (N_1275,In_926,In_2139);
or U1276 (N_1276,In_594,In_2427);
nor U1277 (N_1277,In_1348,In_122);
and U1278 (N_1278,In_444,In_1247);
or U1279 (N_1279,In_931,In_360);
nor U1280 (N_1280,In_58,In_187);
or U1281 (N_1281,In_355,In_1218);
xor U1282 (N_1282,In_1513,In_322);
nor U1283 (N_1283,In_1087,In_718);
nand U1284 (N_1284,In_2087,In_354);
or U1285 (N_1285,In_2380,In_296);
nor U1286 (N_1286,In_236,In_2175);
nor U1287 (N_1287,In_1092,In_261);
or U1288 (N_1288,In_102,In_531);
nand U1289 (N_1289,In_2129,In_102);
xor U1290 (N_1290,In_1890,In_1052);
xnor U1291 (N_1291,In_1924,In_2068);
or U1292 (N_1292,In_906,In_32);
xnor U1293 (N_1293,In_296,In_2237);
and U1294 (N_1294,In_1181,In_442);
or U1295 (N_1295,In_1404,In_428);
and U1296 (N_1296,In_1508,In_1561);
nor U1297 (N_1297,In_73,In_35);
nand U1298 (N_1298,In_1785,In_2275);
nand U1299 (N_1299,In_2151,In_1296);
xnor U1300 (N_1300,In_43,In_2281);
or U1301 (N_1301,In_2291,In_2304);
nor U1302 (N_1302,In_135,In_2079);
nor U1303 (N_1303,In_1174,In_212);
or U1304 (N_1304,In_562,In_2388);
nor U1305 (N_1305,In_2261,In_2183);
nand U1306 (N_1306,In_2484,In_1761);
or U1307 (N_1307,In_2049,In_2239);
xor U1308 (N_1308,In_686,In_1330);
xor U1309 (N_1309,In_1754,In_1080);
or U1310 (N_1310,In_1059,In_288);
nand U1311 (N_1311,In_419,In_2345);
nor U1312 (N_1312,In_2259,In_671);
and U1313 (N_1313,In_2421,In_1038);
xnor U1314 (N_1314,In_2423,In_895);
nor U1315 (N_1315,In_2263,In_1134);
or U1316 (N_1316,In_2323,In_1906);
or U1317 (N_1317,In_1144,In_2019);
nand U1318 (N_1318,In_539,In_605);
nor U1319 (N_1319,In_1592,In_49);
and U1320 (N_1320,In_161,In_1846);
nand U1321 (N_1321,In_670,In_258);
xnor U1322 (N_1322,In_1655,In_1522);
xnor U1323 (N_1323,In_695,In_1699);
xor U1324 (N_1324,In_1014,In_1734);
and U1325 (N_1325,In_1518,In_638);
or U1326 (N_1326,In_2071,In_2118);
and U1327 (N_1327,In_2390,In_1901);
or U1328 (N_1328,In_634,In_2146);
nor U1329 (N_1329,In_1353,In_283);
and U1330 (N_1330,In_1384,In_1989);
nor U1331 (N_1331,In_915,In_2459);
and U1332 (N_1332,In_2421,In_1787);
nor U1333 (N_1333,In_1885,In_1044);
or U1334 (N_1334,In_1410,In_480);
xnor U1335 (N_1335,In_558,In_928);
and U1336 (N_1336,In_158,In_938);
nand U1337 (N_1337,In_1974,In_1635);
and U1338 (N_1338,In_1170,In_1173);
nor U1339 (N_1339,In_676,In_1185);
xnor U1340 (N_1340,In_1149,In_2290);
and U1341 (N_1341,In_839,In_1548);
nand U1342 (N_1342,In_1123,In_336);
xor U1343 (N_1343,In_1443,In_1425);
nor U1344 (N_1344,In_1641,In_362);
nand U1345 (N_1345,In_711,In_2213);
and U1346 (N_1346,In_2360,In_2301);
nor U1347 (N_1347,In_418,In_375);
or U1348 (N_1348,In_1965,In_1987);
xor U1349 (N_1349,In_702,In_966);
and U1350 (N_1350,In_2203,In_2044);
xor U1351 (N_1351,In_434,In_1897);
nand U1352 (N_1352,In_371,In_210);
xnor U1353 (N_1353,In_55,In_1857);
or U1354 (N_1354,In_1117,In_660);
xor U1355 (N_1355,In_469,In_380);
and U1356 (N_1356,In_1332,In_1950);
xnor U1357 (N_1357,In_112,In_2079);
nand U1358 (N_1358,In_340,In_2055);
or U1359 (N_1359,In_1712,In_509);
nand U1360 (N_1360,In_2347,In_651);
or U1361 (N_1361,In_499,In_818);
or U1362 (N_1362,In_1593,In_2225);
nand U1363 (N_1363,In_98,In_1134);
nor U1364 (N_1364,In_157,In_1411);
or U1365 (N_1365,In_2022,In_232);
or U1366 (N_1366,In_2202,In_2163);
nand U1367 (N_1367,In_1657,In_238);
xor U1368 (N_1368,In_884,In_600);
xor U1369 (N_1369,In_84,In_1603);
nand U1370 (N_1370,In_1300,In_1946);
or U1371 (N_1371,In_1559,In_79);
xnor U1372 (N_1372,In_1368,In_2169);
or U1373 (N_1373,In_155,In_1883);
and U1374 (N_1374,In_2074,In_2148);
and U1375 (N_1375,In_2446,In_1068);
nand U1376 (N_1376,In_806,In_1930);
nand U1377 (N_1377,In_1794,In_1429);
or U1378 (N_1378,In_1427,In_223);
nand U1379 (N_1379,In_521,In_132);
nand U1380 (N_1380,In_20,In_2284);
or U1381 (N_1381,In_1309,In_1041);
and U1382 (N_1382,In_2280,In_277);
nand U1383 (N_1383,In_2485,In_1244);
and U1384 (N_1384,In_1491,In_2014);
xor U1385 (N_1385,In_1945,In_1080);
or U1386 (N_1386,In_2040,In_1015);
nand U1387 (N_1387,In_47,In_553);
nand U1388 (N_1388,In_1984,In_1916);
nor U1389 (N_1389,In_697,In_206);
nor U1390 (N_1390,In_245,In_302);
nor U1391 (N_1391,In_656,In_2034);
nand U1392 (N_1392,In_1995,In_623);
nor U1393 (N_1393,In_1389,In_1454);
nor U1394 (N_1394,In_722,In_2108);
nand U1395 (N_1395,In_949,In_749);
nand U1396 (N_1396,In_254,In_2485);
nor U1397 (N_1397,In_1030,In_1004);
or U1398 (N_1398,In_1992,In_1860);
nor U1399 (N_1399,In_1114,In_1306);
or U1400 (N_1400,In_676,In_881);
and U1401 (N_1401,In_1070,In_1701);
nor U1402 (N_1402,In_1708,In_762);
and U1403 (N_1403,In_2035,In_256);
and U1404 (N_1404,In_957,In_678);
xor U1405 (N_1405,In_1735,In_895);
and U1406 (N_1406,In_2204,In_389);
and U1407 (N_1407,In_1858,In_318);
nor U1408 (N_1408,In_863,In_902);
nor U1409 (N_1409,In_208,In_2304);
nor U1410 (N_1410,In_2109,In_500);
nor U1411 (N_1411,In_1510,In_1506);
nor U1412 (N_1412,In_2193,In_2060);
nor U1413 (N_1413,In_2010,In_2044);
or U1414 (N_1414,In_2452,In_1166);
and U1415 (N_1415,In_1116,In_943);
and U1416 (N_1416,In_1634,In_820);
nand U1417 (N_1417,In_1933,In_2115);
nand U1418 (N_1418,In_508,In_2454);
nor U1419 (N_1419,In_835,In_1091);
xor U1420 (N_1420,In_1514,In_1612);
and U1421 (N_1421,In_1961,In_919);
xor U1422 (N_1422,In_1346,In_168);
and U1423 (N_1423,In_904,In_305);
nand U1424 (N_1424,In_1868,In_639);
nand U1425 (N_1425,In_1418,In_2132);
or U1426 (N_1426,In_58,In_1593);
nand U1427 (N_1427,In_1670,In_1214);
nand U1428 (N_1428,In_1089,In_2381);
nor U1429 (N_1429,In_23,In_1436);
nand U1430 (N_1430,In_1873,In_1877);
nor U1431 (N_1431,In_31,In_531);
and U1432 (N_1432,In_1619,In_9);
or U1433 (N_1433,In_1436,In_1036);
xor U1434 (N_1434,In_1022,In_400);
xor U1435 (N_1435,In_177,In_67);
and U1436 (N_1436,In_1709,In_2298);
nor U1437 (N_1437,In_1277,In_2393);
nor U1438 (N_1438,In_1914,In_537);
or U1439 (N_1439,In_182,In_1500);
nand U1440 (N_1440,In_711,In_373);
nor U1441 (N_1441,In_1259,In_320);
or U1442 (N_1442,In_1074,In_2152);
xnor U1443 (N_1443,In_1628,In_108);
nand U1444 (N_1444,In_262,In_1389);
nor U1445 (N_1445,In_570,In_2267);
or U1446 (N_1446,In_163,In_1033);
and U1447 (N_1447,In_758,In_2318);
xor U1448 (N_1448,In_1735,In_785);
nor U1449 (N_1449,In_1376,In_52);
or U1450 (N_1450,In_2488,In_2448);
and U1451 (N_1451,In_2403,In_1103);
nand U1452 (N_1452,In_1107,In_1526);
or U1453 (N_1453,In_2191,In_1693);
nand U1454 (N_1454,In_670,In_1565);
nor U1455 (N_1455,In_1741,In_104);
and U1456 (N_1456,In_564,In_2386);
nand U1457 (N_1457,In_316,In_2221);
xor U1458 (N_1458,In_1391,In_882);
nand U1459 (N_1459,In_1421,In_1588);
xor U1460 (N_1460,In_426,In_1390);
or U1461 (N_1461,In_1404,In_1470);
or U1462 (N_1462,In_1436,In_1454);
or U1463 (N_1463,In_1683,In_2378);
or U1464 (N_1464,In_125,In_1367);
and U1465 (N_1465,In_2157,In_1005);
nand U1466 (N_1466,In_1553,In_2240);
and U1467 (N_1467,In_160,In_917);
xnor U1468 (N_1468,In_1350,In_264);
and U1469 (N_1469,In_969,In_1536);
nand U1470 (N_1470,In_1648,In_1537);
or U1471 (N_1471,In_1771,In_480);
xnor U1472 (N_1472,In_2146,In_2006);
nor U1473 (N_1473,In_1389,In_1487);
nand U1474 (N_1474,In_648,In_1908);
nor U1475 (N_1475,In_964,In_1631);
and U1476 (N_1476,In_296,In_1186);
nand U1477 (N_1477,In_1615,In_1693);
or U1478 (N_1478,In_1883,In_1368);
and U1479 (N_1479,In_2209,In_939);
xor U1480 (N_1480,In_2353,In_1351);
and U1481 (N_1481,In_1769,In_2426);
xor U1482 (N_1482,In_617,In_557);
nor U1483 (N_1483,In_1796,In_2313);
and U1484 (N_1484,In_1454,In_580);
xor U1485 (N_1485,In_515,In_1042);
xnor U1486 (N_1486,In_1731,In_780);
nand U1487 (N_1487,In_1017,In_1635);
or U1488 (N_1488,In_542,In_1683);
or U1489 (N_1489,In_244,In_1072);
and U1490 (N_1490,In_2068,In_366);
xnor U1491 (N_1491,In_1823,In_1653);
nor U1492 (N_1492,In_2497,In_2083);
and U1493 (N_1493,In_773,In_404);
nand U1494 (N_1494,In_2299,In_2231);
nor U1495 (N_1495,In_406,In_2001);
xor U1496 (N_1496,In_2291,In_911);
and U1497 (N_1497,In_1690,In_1524);
xor U1498 (N_1498,In_1221,In_1523);
nand U1499 (N_1499,In_1204,In_1066);
xnor U1500 (N_1500,In_1037,In_1307);
or U1501 (N_1501,In_1089,In_104);
and U1502 (N_1502,In_604,In_20);
or U1503 (N_1503,In_805,In_1000);
xor U1504 (N_1504,In_1763,In_761);
nor U1505 (N_1505,In_1179,In_1845);
nor U1506 (N_1506,In_1721,In_2146);
and U1507 (N_1507,In_2040,In_1492);
or U1508 (N_1508,In_1765,In_1209);
xor U1509 (N_1509,In_690,In_154);
nand U1510 (N_1510,In_495,In_2186);
or U1511 (N_1511,In_84,In_1282);
nor U1512 (N_1512,In_1278,In_1354);
and U1513 (N_1513,In_706,In_80);
nand U1514 (N_1514,In_1347,In_1680);
and U1515 (N_1515,In_2183,In_1009);
xnor U1516 (N_1516,In_1384,In_284);
nor U1517 (N_1517,In_142,In_2347);
or U1518 (N_1518,In_1310,In_1403);
nor U1519 (N_1519,In_2392,In_809);
nor U1520 (N_1520,In_183,In_252);
nand U1521 (N_1521,In_862,In_54);
xnor U1522 (N_1522,In_504,In_1392);
or U1523 (N_1523,In_750,In_960);
or U1524 (N_1524,In_1731,In_235);
nor U1525 (N_1525,In_2342,In_94);
nor U1526 (N_1526,In_853,In_1760);
or U1527 (N_1527,In_1479,In_2210);
and U1528 (N_1528,In_1578,In_518);
nor U1529 (N_1529,In_1950,In_905);
xnor U1530 (N_1530,In_389,In_149);
nand U1531 (N_1531,In_1998,In_379);
nor U1532 (N_1532,In_2387,In_2460);
nand U1533 (N_1533,In_1293,In_2398);
xnor U1534 (N_1534,In_2122,In_449);
or U1535 (N_1535,In_2075,In_179);
nor U1536 (N_1536,In_2453,In_1465);
or U1537 (N_1537,In_2119,In_2174);
xnor U1538 (N_1538,In_1069,In_2059);
xor U1539 (N_1539,In_694,In_1785);
nand U1540 (N_1540,In_458,In_726);
or U1541 (N_1541,In_464,In_1074);
nand U1542 (N_1542,In_901,In_966);
and U1543 (N_1543,In_2483,In_2170);
or U1544 (N_1544,In_1036,In_774);
or U1545 (N_1545,In_1526,In_1660);
or U1546 (N_1546,In_96,In_169);
nor U1547 (N_1547,In_348,In_1064);
nand U1548 (N_1548,In_1945,In_1717);
or U1549 (N_1549,In_1812,In_1242);
and U1550 (N_1550,In_772,In_1468);
or U1551 (N_1551,In_1146,In_2484);
xor U1552 (N_1552,In_511,In_1687);
xnor U1553 (N_1553,In_1398,In_1115);
nand U1554 (N_1554,In_707,In_507);
nor U1555 (N_1555,In_371,In_2015);
or U1556 (N_1556,In_1375,In_665);
and U1557 (N_1557,In_643,In_821);
nand U1558 (N_1558,In_900,In_1290);
nor U1559 (N_1559,In_2129,In_1347);
or U1560 (N_1560,In_2235,In_1274);
and U1561 (N_1561,In_2323,In_1201);
or U1562 (N_1562,In_1843,In_2082);
nor U1563 (N_1563,In_254,In_101);
xnor U1564 (N_1564,In_1110,In_2344);
nor U1565 (N_1565,In_1439,In_973);
nand U1566 (N_1566,In_2321,In_957);
nand U1567 (N_1567,In_378,In_548);
nor U1568 (N_1568,In_899,In_1060);
xor U1569 (N_1569,In_2466,In_2013);
nand U1570 (N_1570,In_938,In_234);
or U1571 (N_1571,In_2278,In_307);
xnor U1572 (N_1572,In_1706,In_1878);
or U1573 (N_1573,In_1041,In_178);
or U1574 (N_1574,In_2165,In_854);
nor U1575 (N_1575,In_146,In_2158);
nand U1576 (N_1576,In_464,In_2237);
or U1577 (N_1577,In_1056,In_248);
or U1578 (N_1578,In_927,In_1685);
and U1579 (N_1579,In_2380,In_362);
and U1580 (N_1580,In_376,In_662);
nor U1581 (N_1581,In_2406,In_428);
xnor U1582 (N_1582,In_1412,In_388);
xnor U1583 (N_1583,In_1750,In_2232);
nand U1584 (N_1584,In_1705,In_213);
nand U1585 (N_1585,In_190,In_1481);
nor U1586 (N_1586,In_1369,In_1103);
nor U1587 (N_1587,In_2319,In_1778);
xnor U1588 (N_1588,In_2244,In_44);
nand U1589 (N_1589,In_1144,In_836);
xnor U1590 (N_1590,In_1080,In_546);
and U1591 (N_1591,In_1688,In_1503);
and U1592 (N_1592,In_248,In_218);
nor U1593 (N_1593,In_722,In_2355);
xor U1594 (N_1594,In_1076,In_140);
or U1595 (N_1595,In_1635,In_1911);
and U1596 (N_1596,In_1495,In_1280);
xnor U1597 (N_1597,In_859,In_806);
and U1598 (N_1598,In_49,In_1514);
xor U1599 (N_1599,In_868,In_2332);
and U1600 (N_1600,In_839,In_393);
nor U1601 (N_1601,In_459,In_378);
and U1602 (N_1602,In_653,In_722);
xnor U1603 (N_1603,In_938,In_2325);
and U1604 (N_1604,In_1911,In_1285);
nor U1605 (N_1605,In_42,In_1124);
or U1606 (N_1606,In_290,In_1386);
xnor U1607 (N_1607,In_1435,In_1369);
and U1608 (N_1608,In_2032,In_1616);
xor U1609 (N_1609,In_1143,In_1845);
and U1610 (N_1610,In_382,In_1933);
nor U1611 (N_1611,In_2179,In_784);
nor U1612 (N_1612,In_2126,In_551);
nor U1613 (N_1613,In_644,In_1922);
nand U1614 (N_1614,In_962,In_683);
or U1615 (N_1615,In_1524,In_216);
nor U1616 (N_1616,In_1257,In_2272);
nor U1617 (N_1617,In_2299,In_800);
or U1618 (N_1618,In_1508,In_1878);
nand U1619 (N_1619,In_1247,In_1774);
nor U1620 (N_1620,In_212,In_1983);
and U1621 (N_1621,In_382,In_174);
nor U1622 (N_1622,In_1680,In_913);
or U1623 (N_1623,In_687,In_1187);
nor U1624 (N_1624,In_1636,In_1483);
or U1625 (N_1625,In_1239,In_2135);
nor U1626 (N_1626,In_1076,In_1978);
nand U1627 (N_1627,In_1271,In_1915);
nor U1628 (N_1628,In_1475,In_2460);
nand U1629 (N_1629,In_1708,In_309);
xnor U1630 (N_1630,In_1100,In_474);
nand U1631 (N_1631,In_1771,In_1950);
nor U1632 (N_1632,In_1208,In_531);
or U1633 (N_1633,In_1236,In_1034);
nand U1634 (N_1634,In_2120,In_1189);
nand U1635 (N_1635,In_930,In_2368);
nor U1636 (N_1636,In_2164,In_30);
nand U1637 (N_1637,In_1092,In_1546);
nand U1638 (N_1638,In_17,In_372);
xnor U1639 (N_1639,In_1088,In_1302);
xor U1640 (N_1640,In_271,In_997);
or U1641 (N_1641,In_2030,In_1595);
xor U1642 (N_1642,In_655,In_1274);
nor U1643 (N_1643,In_304,In_2425);
nor U1644 (N_1644,In_1519,In_2413);
and U1645 (N_1645,In_261,In_436);
or U1646 (N_1646,In_425,In_633);
xor U1647 (N_1647,In_1850,In_371);
or U1648 (N_1648,In_62,In_533);
nor U1649 (N_1649,In_1259,In_722);
and U1650 (N_1650,In_2473,In_1573);
and U1651 (N_1651,In_1066,In_1401);
nand U1652 (N_1652,In_476,In_2290);
or U1653 (N_1653,In_155,In_145);
nand U1654 (N_1654,In_269,In_1576);
and U1655 (N_1655,In_2397,In_665);
or U1656 (N_1656,In_1906,In_2199);
nand U1657 (N_1657,In_1130,In_1406);
xnor U1658 (N_1658,In_202,In_2145);
nor U1659 (N_1659,In_694,In_1998);
and U1660 (N_1660,In_1924,In_723);
xnor U1661 (N_1661,In_1015,In_1452);
nor U1662 (N_1662,In_230,In_2261);
and U1663 (N_1663,In_651,In_2093);
and U1664 (N_1664,In_1864,In_621);
and U1665 (N_1665,In_904,In_1666);
and U1666 (N_1666,In_330,In_1161);
xnor U1667 (N_1667,In_137,In_2030);
and U1668 (N_1668,In_2109,In_1868);
xor U1669 (N_1669,In_1272,In_1064);
xnor U1670 (N_1670,In_2459,In_291);
and U1671 (N_1671,In_2100,In_1468);
or U1672 (N_1672,In_1333,In_2462);
nand U1673 (N_1673,In_607,In_1936);
or U1674 (N_1674,In_381,In_440);
xnor U1675 (N_1675,In_345,In_490);
and U1676 (N_1676,In_2154,In_2438);
or U1677 (N_1677,In_2349,In_2085);
and U1678 (N_1678,In_1517,In_134);
nor U1679 (N_1679,In_1847,In_1114);
and U1680 (N_1680,In_545,In_1940);
or U1681 (N_1681,In_2244,In_1668);
nor U1682 (N_1682,In_135,In_1869);
nor U1683 (N_1683,In_390,In_252);
nor U1684 (N_1684,In_1004,In_1734);
and U1685 (N_1685,In_2307,In_565);
nand U1686 (N_1686,In_1222,In_1202);
nor U1687 (N_1687,In_1319,In_1557);
xor U1688 (N_1688,In_815,In_2294);
nor U1689 (N_1689,In_618,In_1998);
xor U1690 (N_1690,In_1264,In_1793);
nand U1691 (N_1691,In_1561,In_1985);
nand U1692 (N_1692,In_915,In_1345);
nor U1693 (N_1693,In_1991,In_327);
nand U1694 (N_1694,In_996,In_2431);
nand U1695 (N_1695,In_1362,In_889);
xor U1696 (N_1696,In_718,In_369);
nand U1697 (N_1697,In_1041,In_468);
xnor U1698 (N_1698,In_859,In_1887);
and U1699 (N_1699,In_1929,In_409);
nand U1700 (N_1700,In_586,In_1535);
xor U1701 (N_1701,In_790,In_2008);
nand U1702 (N_1702,In_992,In_1242);
or U1703 (N_1703,In_683,In_142);
and U1704 (N_1704,In_2014,In_593);
nor U1705 (N_1705,In_1555,In_887);
nand U1706 (N_1706,In_1561,In_224);
or U1707 (N_1707,In_1740,In_2276);
nor U1708 (N_1708,In_802,In_2403);
xnor U1709 (N_1709,In_729,In_1947);
and U1710 (N_1710,In_869,In_1331);
and U1711 (N_1711,In_2468,In_323);
and U1712 (N_1712,In_1539,In_275);
nor U1713 (N_1713,In_1724,In_533);
nor U1714 (N_1714,In_2409,In_1388);
or U1715 (N_1715,In_2408,In_334);
nand U1716 (N_1716,In_2100,In_563);
and U1717 (N_1717,In_1116,In_1226);
nor U1718 (N_1718,In_1934,In_1319);
nor U1719 (N_1719,In_1409,In_1588);
or U1720 (N_1720,In_1104,In_327);
nand U1721 (N_1721,In_474,In_2361);
and U1722 (N_1722,In_283,In_328);
or U1723 (N_1723,In_95,In_2352);
or U1724 (N_1724,In_1675,In_886);
nand U1725 (N_1725,In_542,In_1233);
xor U1726 (N_1726,In_586,In_380);
nand U1727 (N_1727,In_1623,In_157);
and U1728 (N_1728,In_1186,In_885);
nand U1729 (N_1729,In_2358,In_1348);
nor U1730 (N_1730,In_566,In_1886);
nor U1731 (N_1731,In_53,In_1216);
nor U1732 (N_1732,In_1679,In_1366);
nand U1733 (N_1733,In_937,In_603);
and U1734 (N_1734,In_2489,In_226);
and U1735 (N_1735,In_1327,In_1725);
or U1736 (N_1736,In_1180,In_1504);
or U1737 (N_1737,In_1898,In_1911);
xor U1738 (N_1738,In_2330,In_332);
or U1739 (N_1739,In_1390,In_51);
nor U1740 (N_1740,In_658,In_2448);
and U1741 (N_1741,In_2261,In_298);
or U1742 (N_1742,In_2256,In_861);
and U1743 (N_1743,In_615,In_1693);
or U1744 (N_1744,In_1676,In_1874);
xor U1745 (N_1745,In_571,In_1305);
and U1746 (N_1746,In_1722,In_476);
nor U1747 (N_1747,In_2473,In_1541);
and U1748 (N_1748,In_228,In_1529);
or U1749 (N_1749,In_966,In_416);
or U1750 (N_1750,In_2373,In_1585);
nor U1751 (N_1751,In_2134,In_1464);
nor U1752 (N_1752,In_2037,In_1140);
and U1753 (N_1753,In_2063,In_2270);
and U1754 (N_1754,In_2482,In_778);
and U1755 (N_1755,In_1611,In_462);
or U1756 (N_1756,In_1964,In_1592);
and U1757 (N_1757,In_465,In_1488);
xnor U1758 (N_1758,In_1327,In_1996);
xor U1759 (N_1759,In_2137,In_766);
nor U1760 (N_1760,In_1911,In_823);
and U1761 (N_1761,In_1069,In_1248);
and U1762 (N_1762,In_1942,In_1745);
or U1763 (N_1763,In_1588,In_1363);
nand U1764 (N_1764,In_1643,In_1111);
and U1765 (N_1765,In_816,In_2166);
nor U1766 (N_1766,In_389,In_816);
or U1767 (N_1767,In_228,In_764);
xor U1768 (N_1768,In_1022,In_1007);
or U1769 (N_1769,In_1494,In_191);
nor U1770 (N_1770,In_192,In_1813);
nand U1771 (N_1771,In_1921,In_1331);
and U1772 (N_1772,In_277,In_513);
or U1773 (N_1773,In_2098,In_1245);
nor U1774 (N_1774,In_83,In_740);
nor U1775 (N_1775,In_671,In_251);
xnor U1776 (N_1776,In_2269,In_1281);
nand U1777 (N_1777,In_882,In_794);
xor U1778 (N_1778,In_1398,In_1755);
or U1779 (N_1779,In_1674,In_456);
nand U1780 (N_1780,In_1867,In_681);
nor U1781 (N_1781,In_1405,In_707);
nand U1782 (N_1782,In_1226,In_1650);
or U1783 (N_1783,In_410,In_1017);
or U1784 (N_1784,In_523,In_1130);
xor U1785 (N_1785,In_977,In_2110);
nand U1786 (N_1786,In_116,In_1212);
nand U1787 (N_1787,In_429,In_2433);
and U1788 (N_1788,In_2202,In_1765);
nand U1789 (N_1789,In_663,In_1062);
and U1790 (N_1790,In_34,In_1653);
xor U1791 (N_1791,In_1335,In_591);
nor U1792 (N_1792,In_1548,In_2108);
and U1793 (N_1793,In_846,In_1912);
nand U1794 (N_1794,In_273,In_1903);
or U1795 (N_1795,In_367,In_1246);
or U1796 (N_1796,In_2138,In_743);
xnor U1797 (N_1797,In_628,In_831);
or U1798 (N_1798,In_1168,In_1774);
or U1799 (N_1799,In_1612,In_1873);
nor U1800 (N_1800,In_725,In_828);
and U1801 (N_1801,In_1767,In_1072);
nor U1802 (N_1802,In_2228,In_2233);
and U1803 (N_1803,In_910,In_919);
and U1804 (N_1804,In_2078,In_906);
xnor U1805 (N_1805,In_543,In_1125);
nand U1806 (N_1806,In_80,In_1728);
xor U1807 (N_1807,In_2134,In_2036);
and U1808 (N_1808,In_1304,In_908);
nand U1809 (N_1809,In_883,In_1777);
and U1810 (N_1810,In_1440,In_441);
nand U1811 (N_1811,In_1825,In_651);
nand U1812 (N_1812,In_2419,In_724);
nor U1813 (N_1813,In_2265,In_1801);
nor U1814 (N_1814,In_1112,In_96);
nand U1815 (N_1815,In_500,In_65);
and U1816 (N_1816,In_1504,In_348);
xnor U1817 (N_1817,In_944,In_2108);
xor U1818 (N_1818,In_1187,In_227);
and U1819 (N_1819,In_1817,In_1646);
nand U1820 (N_1820,In_2449,In_1694);
nor U1821 (N_1821,In_2305,In_1358);
or U1822 (N_1822,In_136,In_2447);
and U1823 (N_1823,In_1048,In_405);
and U1824 (N_1824,In_786,In_820);
nor U1825 (N_1825,In_1803,In_1085);
and U1826 (N_1826,In_70,In_808);
nor U1827 (N_1827,In_2003,In_1248);
nor U1828 (N_1828,In_1583,In_2347);
xnor U1829 (N_1829,In_2183,In_1969);
or U1830 (N_1830,In_1775,In_964);
nor U1831 (N_1831,In_533,In_1700);
or U1832 (N_1832,In_1711,In_1043);
nand U1833 (N_1833,In_2146,In_13);
nand U1834 (N_1834,In_318,In_1568);
or U1835 (N_1835,In_142,In_1124);
and U1836 (N_1836,In_1814,In_2439);
nand U1837 (N_1837,In_635,In_502);
xor U1838 (N_1838,In_761,In_2034);
nor U1839 (N_1839,In_637,In_284);
or U1840 (N_1840,In_2149,In_2481);
nand U1841 (N_1841,In_864,In_265);
and U1842 (N_1842,In_2139,In_1692);
or U1843 (N_1843,In_1391,In_1036);
nand U1844 (N_1844,In_646,In_1166);
nor U1845 (N_1845,In_752,In_12);
nand U1846 (N_1846,In_1666,In_1964);
or U1847 (N_1847,In_1970,In_1721);
or U1848 (N_1848,In_648,In_1993);
and U1849 (N_1849,In_435,In_1221);
xnor U1850 (N_1850,In_2488,In_911);
and U1851 (N_1851,In_2322,In_1996);
xor U1852 (N_1852,In_641,In_348);
or U1853 (N_1853,In_2002,In_372);
nor U1854 (N_1854,In_1600,In_1145);
nand U1855 (N_1855,In_1509,In_1046);
nand U1856 (N_1856,In_63,In_1201);
nor U1857 (N_1857,In_1110,In_1385);
or U1858 (N_1858,In_363,In_199);
xnor U1859 (N_1859,In_650,In_673);
nor U1860 (N_1860,In_420,In_545);
xnor U1861 (N_1861,In_1538,In_1764);
nor U1862 (N_1862,In_1171,In_118);
nor U1863 (N_1863,In_2103,In_2081);
nor U1864 (N_1864,In_171,In_2155);
and U1865 (N_1865,In_2214,In_2266);
nand U1866 (N_1866,In_1517,In_1862);
xnor U1867 (N_1867,In_1186,In_217);
and U1868 (N_1868,In_2157,In_972);
and U1869 (N_1869,In_2253,In_2018);
nand U1870 (N_1870,In_2124,In_1273);
nor U1871 (N_1871,In_1513,In_2414);
xnor U1872 (N_1872,In_2000,In_1877);
nand U1873 (N_1873,In_258,In_361);
nand U1874 (N_1874,In_1848,In_238);
nand U1875 (N_1875,In_255,In_1236);
and U1876 (N_1876,In_1817,In_2293);
xor U1877 (N_1877,In_886,In_265);
and U1878 (N_1878,In_934,In_1953);
and U1879 (N_1879,In_166,In_1092);
or U1880 (N_1880,In_2379,In_1825);
and U1881 (N_1881,In_1732,In_1674);
nor U1882 (N_1882,In_1014,In_742);
xor U1883 (N_1883,In_2056,In_2396);
nand U1884 (N_1884,In_2008,In_597);
xor U1885 (N_1885,In_2214,In_1927);
and U1886 (N_1886,In_1460,In_1686);
nand U1887 (N_1887,In_782,In_1162);
nand U1888 (N_1888,In_1602,In_622);
nand U1889 (N_1889,In_747,In_342);
nand U1890 (N_1890,In_884,In_2076);
xor U1891 (N_1891,In_2358,In_49);
nor U1892 (N_1892,In_205,In_207);
nand U1893 (N_1893,In_82,In_517);
nor U1894 (N_1894,In_211,In_939);
xnor U1895 (N_1895,In_883,In_437);
or U1896 (N_1896,In_1481,In_1932);
or U1897 (N_1897,In_147,In_2456);
and U1898 (N_1898,In_1835,In_2486);
or U1899 (N_1899,In_846,In_1501);
xor U1900 (N_1900,In_2214,In_1778);
nand U1901 (N_1901,In_318,In_8);
or U1902 (N_1902,In_890,In_186);
nor U1903 (N_1903,In_432,In_1050);
xnor U1904 (N_1904,In_1812,In_467);
or U1905 (N_1905,In_2127,In_202);
and U1906 (N_1906,In_948,In_1648);
nor U1907 (N_1907,In_1474,In_1585);
xnor U1908 (N_1908,In_73,In_1934);
and U1909 (N_1909,In_331,In_2279);
xnor U1910 (N_1910,In_451,In_1518);
nor U1911 (N_1911,In_2301,In_2329);
xnor U1912 (N_1912,In_1934,In_343);
xor U1913 (N_1913,In_1756,In_1328);
nor U1914 (N_1914,In_1451,In_347);
or U1915 (N_1915,In_2369,In_424);
nand U1916 (N_1916,In_1608,In_341);
nand U1917 (N_1917,In_1940,In_2374);
nand U1918 (N_1918,In_1486,In_2471);
or U1919 (N_1919,In_1379,In_2074);
or U1920 (N_1920,In_6,In_144);
and U1921 (N_1921,In_828,In_771);
nand U1922 (N_1922,In_2398,In_1457);
nor U1923 (N_1923,In_2099,In_2111);
or U1924 (N_1924,In_457,In_1344);
xnor U1925 (N_1925,In_1039,In_1671);
xnor U1926 (N_1926,In_2491,In_615);
and U1927 (N_1927,In_116,In_1294);
xor U1928 (N_1928,In_853,In_828);
and U1929 (N_1929,In_570,In_273);
nand U1930 (N_1930,In_475,In_1893);
xnor U1931 (N_1931,In_2344,In_946);
and U1932 (N_1932,In_52,In_996);
and U1933 (N_1933,In_633,In_1572);
and U1934 (N_1934,In_1843,In_1046);
xor U1935 (N_1935,In_1696,In_1841);
nor U1936 (N_1936,In_1382,In_2088);
xor U1937 (N_1937,In_827,In_472);
nand U1938 (N_1938,In_20,In_1151);
nor U1939 (N_1939,In_1341,In_2294);
nor U1940 (N_1940,In_1165,In_1838);
and U1941 (N_1941,In_1589,In_767);
nand U1942 (N_1942,In_1681,In_1655);
or U1943 (N_1943,In_420,In_2385);
or U1944 (N_1944,In_1770,In_1916);
nand U1945 (N_1945,In_2124,In_355);
nor U1946 (N_1946,In_1383,In_196);
and U1947 (N_1947,In_1214,In_2192);
and U1948 (N_1948,In_2431,In_500);
or U1949 (N_1949,In_2226,In_870);
and U1950 (N_1950,In_1969,In_1585);
nor U1951 (N_1951,In_379,In_237);
nor U1952 (N_1952,In_42,In_1068);
or U1953 (N_1953,In_2273,In_1828);
and U1954 (N_1954,In_13,In_1769);
nand U1955 (N_1955,In_768,In_108);
nor U1956 (N_1956,In_1336,In_260);
nor U1957 (N_1957,In_1188,In_1814);
nand U1958 (N_1958,In_1802,In_1626);
and U1959 (N_1959,In_420,In_648);
and U1960 (N_1960,In_1780,In_1322);
nor U1961 (N_1961,In_2292,In_1282);
xor U1962 (N_1962,In_1349,In_839);
nor U1963 (N_1963,In_539,In_2118);
and U1964 (N_1964,In_455,In_887);
and U1965 (N_1965,In_1267,In_1086);
nor U1966 (N_1966,In_407,In_1285);
nor U1967 (N_1967,In_784,In_1248);
or U1968 (N_1968,In_1681,In_590);
or U1969 (N_1969,In_1488,In_642);
or U1970 (N_1970,In_1612,In_1875);
nand U1971 (N_1971,In_1107,In_988);
or U1972 (N_1972,In_2380,In_133);
or U1973 (N_1973,In_451,In_96);
or U1974 (N_1974,In_368,In_1269);
xnor U1975 (N_1975,In_1077,In_654);
or U1976 (N_1976,In_1197,In_2312);
nand U1977 (N_1977,In_1025,In_522);
or U1978 (N_1978,In_956,In_429);
and U1979 (N_1979,In_2285,In_622);
nor U1980 (N_1980,In_1955,In_1180);
xnor U1981 (N_1981,In_997,In_290);
or U1982 (N_1982,In_2217,In_1594);
and U1983 (N_1983,In_1537,In_693);
nor U1984 (N_1984,In_1613,In_1747);
xor U1985 (N_1985,In_1041,In_2074);
nand U1986 (N_1986,In_213,In_1817);
or U1987 (N_1987,In_410,In_291);
or U1988 (N_1988,In_29,In_2358);
xnor U1989 (N_1989,In_504,In_44);
xnor U1990 (N_1990,In_2383,In_1991);
nand U1991 (N_1991,In_1724,In_340);
xnor U1992 (N_1992,In_186,In_1017);
nand U1993 (N_1993,In_236,In_1435);
nand U1994 (N_1994,In_2476,In_1198);
or U1995 (N_1995,In_605,In_448);
nand U1996 (N_1996,In_220,In_2251);
or U1997 (N_1997,In_223,In_503);
nand U1998 (N_1998,In_608,In_2102);
xor U1999 (N_1999,In_71,In_335);
and U2000 (N_2000,In_79,In_544);
or U2001 (N_2001,In_2103,In_415);
and U2002 (N_2002,In_1410,In_1513);
nand U2003 (N_2003,In_322,In_875);
or U2004 (N_2004,In_1511,In_1986);
and U2005 (N_2005,In_322,In_781);
xnor U2006 (N_2006,In_796,In_2037);
and U2007 (N_2007,In_2307,In_2182);
or U2008 (N_2008,In_270,In_1164);
nand U2009 (N_2009,In_2273,In_1185);
or U2010 (N_2010,In_215,In_775);
and U2011 (N_2011,In_727,In_1353);
and U2012 (N_2012,In_1353,In_1754);
nand U2013 (N_2013,In_640,In_1424);
and U2014 (N_2014,In_1432,In_1408);
nand U2015 (N_2015,In_1444,In_1990);
and U2016 (N_2016,In_1929,In_2100);
nand U2017 (N_2017,In_2452,In_332);
and U2018 (N_2018,In_1565,In_1241);
nor U2019 (N_2019,In_2311,In_307);
and U2020 (N_2020,In_1991,In_1689);
nand U2021 (N_2021,In_194,In_1050);
and U2022 (N_2022,In_1296,In_1712);
and U2023 (N_2023,In_943,In_1495);
and U2024 (N_2024,In_774,In_1109);
xor U2025 (N_2025,In_2460,In_1854);
nor U2026 (N_2026,In_447,In_426);
nor U2027 (N_2027,In_278,In_555);
nor U2028 (N_2028,In_932,In_239);
nor U2029 (N_2029,In_2251,In_785);
nor U2030 (N_2030,In_568,In_498);
or U2031 (N_2031,In_1850,In_1846);
nor U2032 (N_2032,In_1335,In_641);
or U2033 (N_2033,In_1212,In_677);
or U2034 (N_2034,In_1806,In_408);
or U2035 (N_2035,In_1221,In_1463);
or U2036 (N_2036,In_541,In_214);
xnor U2037 (N_2037,In_2219,In_1676);
or U2038 (N_2038,In_1058,In_1757);
nor U2039 (N_2039,In_2292,In_135);
and U2040 (N_2040,In_1508,In_1885);
and U2041 (N_2041,In_1131,In_842);
nor U2042 (N_2042,In_1064,In_1063);
and U2043 (N_2043,In_1708,In_637);
nor U2044 (N_2044,In_982,In_1070);
xnor U2045 (N_2045,In_1720,In_2053);
or U2046 (N_2046,In_1424,In_486);
nand U2047 (N_2047,In_286,In_1300);
or U2048 (N_2048,In_256,In_358);
or U2049 (N_2049,In_2199,In_1719);
xnor U2050 (N_2050,In_353,In_1938);
nand U2051 (N_2051,In_858,In_28);
and U2052 (N_2052,In_2350,In_971);
nand U2053 (N_2053,In_392,In_2175);
and U2054 (N_2054,In_227,In_1504);
xnor U2055 (N_2055,In_132,In_429);
nor U2056 (N_2056,In_175,In_689);
xnor U2057 (N_2057,In_1482,In_2326);
or U2058 (N_2058,In_1503,In_989);
and U2059 (N_2059,In_436,In_2311);
nor U2060 (N_2060,In_1103,In_716);
and U2061 (N_2061,In_540,In_932);
or U2062 (N_2062,In_254,In_577);
and U2063 (N_2063,In_1321,In_1255);
and U2064 (N_2064,In_1684,In_968);
xnor U2065 (N_2065,In_62,In_2145);
or U2066 (N_2066,In_479,In_96);
nor U2067 (N_2067,In_1898,In_1692);
or U2068 (N_2068,In_2382,In_832);
nand U2069 (N_2069,In_1354,In_1309);
nor U2070 (N_2070,In_1483,In_556);
or U2071 (N_2071,In_1492,In_1890);
xor U2072 (N_2072,In_725,In_2088);
nor U2073 (N_2073,In_466,In_1095);
or U2074 (N_2074,In_743,In_1515);
xor U2075 (N_2075,In_2323,In_2004);
nand U2076 (N_2076,In_663,In_220);
or U2077 (N_2077,In_895,In_1376);
or U2078 (N_2078,In_790,In_2019);
or U2079 (N_2079,In_1007,In_219);
and U2080 (N_2080,In_572,In_558);
or U2081 (N_2081,In_1660,In_260);
or U2082 (N_2082,In_1147,In_1329);
and U2083 (N_2083,In_741,In_2170);
nand U2084 (N_2084,In_2184,In_2131);
xor U2085 (N_2085,In_886,In_1585);
nor U2086 (N_2086,In_2106,In_2119);
and U2087 (N_2087,In_2043,In_271);
or U2088 (N_2088,In_2301,In_2255);
and U2089 (N_2089,In_682,In_2395);
and U2090 (N_2090,In_2462,In_1727);
or U2091 (N_2091,In_1363,In_1239);
or U2092 (N_2092,In_1932,In_560);
and U2093 (N_2093,In_851,In_2140);
and U2094 (N_2094,In_1417,In_1770);
and U2095 (N_2095,In_2166,In_1457);
and U2096 (N_2096,In_1463,In_2);
xor U2097 (N_2097,In_190,In_781);
nand U2098 (N_2098,In_1154,In_1242);
nand U2099 (N_2099,In_2247,In_2004);
xor U2100 (N_2100,In_1768,In_589);
and U2101 (N_2101,In_1259,In_1334);
nor U2102 (N_2102,In_2498,In_817);
and U2103 (N_2103,In_1244,In_1207);
and U2104 (N_2104,In_2032,In_1021);
xor U2105 (N_2105,In_2046,In_552);
and U2106 (N_2106,In_1772,In_252);
nand U2107 (N_2107,In_756,In_797);
or U2108 (N_2108,In_1269,In_880);
nor U2109 (N_2109,In_1847,In_1517);
or U2110 (N_2110,In_189,In_79);
or U2111 (N_2111,In_312,In_402);
or U2112 (N_2112,In_1222,In_599);
or U2113 (N_2113,In_1125,In_1603);
and U2114 (N_2114,In_560,In_1707);
nor U2115 (N_2115,In_1441,In_134);
nor U2116 (N_2116,In_1006,In_1110);
xor U2117 (N_2117,In_2306,In_2416);
nand U2118 (N_2118,In_1651,In_1636);
or U2119 (N_2119,In_780,In_2279);
nand U2120 (N_2120,In_1784,In_352);
nand U2121 (N_2121,In_1252,In_2194);
nor U2122 (N_2122,In_1725,In_313);
or U2123 (N_2123,In_1773,In_2265);
nand U2124 (N_2124,In_1931,In_1743);
nor U2125 (N_2125,In_545,In_1031);
and U2126 (N_2126,In_2376,In_1039);
nor U2127 (N_2127,In_2075,In_1550);
xor U2128 (N_2128,In_583,In_731);
nand U2129 (N_2129,In_1734,In_1638);
and U2130 (N_2130,In_1486,In_927);
and U2131 (N_2131,In_2459,In_181);
xnor U2132 (N_2132,In_2375,In_1392);
and U2133 (N_2133,In_646,In_721);
nor U2134 (N_2134,In_2086,In_720);
or U2135 (N_2135,In_86,In_1130);
nor U2136 (N_2136,In_2206,In_301);
xnor U2137 (N_2137,In_221,In_1001);
xor U2138 (N_2138,In_748,In_1487);
and U2139 (N_2139,In_1392,In_508);
and U2140 (N_2140,In_425,In_1505);
nand U2141 (N_2141,In_2019,In_71);
nor U2142 (N_2142,In_2280,In_1732);
and U2143 (N_2143,In_1263,In_857);
nand U2144 (N_2144,In_1236,In_903);
nand U2145 (N_2145,In_1537,In_139);
or U2146 (N_2146,In_2437,In_1491);
and U2147 (N_2147,In_1774,In_1323);
and U2148 (N_2148,In_1992,In_312);
nand U2149 (N_2149,In_1575,In_1472);
xor U2150 (N_2150,In_1995,In_953);
and U2151 (N_2151,In_477,In_923);
xnor U2152 (N_2152,In_1686,In_2367);
or U2153 (N_2153,In_1856,In_1153);
or U2154 (N_2154,In_1007,In_202);
nand U2155 (N_2155,In_1960,In_1530);
xnor U2156 (N_2156,In_109,In_838);
xnor U2157 (N_2157,In_2400,In_1411);
or U2158 (N_2158,In_2486,In_1650);
xnor U2159 (N_2159,In_788,In_1208);
xor U2160 (N_2160,In_1235,In_179);
or U2161 (N_2161,In_805,In_519);
or U2162 (N_2162,In_877,In_1651);
nand U2163 (N_2163,In_2061,In_405);
xor U2164 (N_2164,In_2168,In_851);
nor U2165 (N_2165,In_272,In_1274);
or U2166 (N_2166,In_98,In_544);
nand U2167 (N_2167,In_1635,In_412);
and U2168 (N_2168,In_1154,In_105);
xnor U2169 (N_2169,In_1945,In_707);
xor U2170 (N_2170,In_1141,In_1604);
nor U2171 (N_2171,In_1248,In_1290);
xor U2172 (N_2172,In_1048,In_2425);
nand U2173 (N_2173,In_17,In_157);
or U2174 (N_2174,In_1538,In_1557);
nor U2175 (N_2175,In_1927,In_2258);
and U2176 (N_2176,In_397,In_337);
nand U2177 (N_2177,In_1028,In_150);
or U2178 (N_2178,In_2272,In_1179);
nor U2179 (N_2179,In_1726,In_2221);
nor U2180 (N_2180,In_982,In_2342);
xor U2181 (N_2181,In_2396,In_283);
and U2182 (N_2182,In_892,In_408);
or U2183 (N_2183,In_2429,In_209);
xor U2184 (N_2184,In_2091,In_556);
nor U2185 (N_2185,In_21,In_1593);
and U2186 (N_2186,In_1340,In_2135);
or U2187 (N_2187,In_1361,In_569);
nor U2188 (N_2188,In_2323,In_164);
or U2189 (N_2189,In_873,In_2163);
nor U2190 (N_2190,In_952,In_1826);
and U2191 (N_2191,In_1228,In_2459);
nor U2192 (N_2192,In_713,In_1964);
and U2193 (N_2193,In_460,In_1992);
or U2194 (N_2194,In_1539,In_2026);
nor U2195 (N_2195,In_871,In_1191);
nor U2196 (N_2196,In_52,In_676);
nor U2197 (N_2197,In_45,In_187);
or U2198 (N_2198,In_2221,In_2125);
xor U2199 (N_2199,In_282,In_212);
nand U2200 (N_2200,In_1417,In_1138);
xnor U2201 (N_2201,In_881,In_582);
or U2202 (N_2202,In_2107,In_1668);
nand U2203 (N_2203,In_1852,In_515);
nor U2204 (N_2204,In_983,In_2);
nand U2205 (N_2205,In_2187,In_2418);
and U2206 (N_2206,In_990,In_519);
nor U2207 (N_2207,In_2335,In_2368);
xor U2208 (N_2208,In_378,In_2422);
nand U2209 (N_2209,In_1790,In_161);
xnor U2210 (N_2210,In_2486,In_217);
and U2211 (N_2211,In_544,In_719);
and U2212 (N_2212,In_77,In_275);
nor U2213 (N_2213,In_1923,In_1354);
nand U2214 (N_2214,In_434,In_1904);
nor U2215 (N_2215,In_2327,In_909);
nand U2216 (N_2216,In_2403,In_1961);
or U2217 (N_2217,In_743,In_1376);
xnor U2218 (N_2218,In_2476,In_1411);
and U2219 (N_2219,In_1833,In_1310);
nand U2220 (N_2220,In_321,In_945);
or U2221 (N_2221,In_376,In_1485);
or U2222 (N_2222,In_1869,In_1626);
or U2223 (N_2223,In_118,In_1873);
nand U2224 (N_2224,In_190,In_181);
xor U2225 (N_2225,In_1338,In_2453);
and U2226 (N_2226,In_1927,In_1986);
and U2227 (N_2227,In_642,In_806);
nand U2228 (N_2228,In_2044,In_1944);
nor U2229 (N_2229,In_1328,In_1035);
nor U2230 (N_2230,In_2348,In_1514);
nor U2231 (N_2231,In_137,In_738);
or U2232 (N_2232,In_210,In_1452);
or U2233 (N_2233,In_2296,In_134);
xnor U2234 (N_2234,In_459,In_848);
nor U2235 (N_2235,In_1158,In_1013);
and U2236 (N_2236,In_726,In_1532);
nor U2237 (N_2237,In_1199,In_828);
and U2238 (N_2238,In_1394,In_1532);
or U2239 (N_2239,In_576,In_1072);
and U2240 (N_2240,In_1605,In_1011);
xor U2241 (N_2241,In_984,In_1389);
nor U2242 (N_2242,In_1247,In_2123);
nor U2243 (N_2243,In_124,In_121);
nand U2244 (N_2244,In_961,In_365);
and U2245 (N_2245,In_1930,In_1675);
nor U2246 (N_2246,In_0,In_2397);
xnor U2247 (N_2247,In_1341,In_1853);
nor U2248 (N_2248,In_18,In_611);
xnor U2249 (N_2249,In_957,In_382);
nor U2250 (N_2250,In_1252,In_1857);
nand U2251 (N_2251,In_1496,In_1846);
xnor U2252 (N_2252,In_1282,In_2122);
or U2253 (N_2253,In_2119,In_463);
or U2254 (N_2254,In_294,In_2202);
or U2255 (N_2255,In_1558,In_1303);
or U2256 (N_2256,In_1289,In_450);
nor U2257 (N_2257,In_1139,In_1757);
xnor U2258 (N_2258,In_523,In_1928);
xnor U2259 (N_2259,In_1715,In_2234);
or U2260 (N_2260,In_1662,In_1434);
and U2261 (N_2261,In_719,In_1464);
and U2262 (N_2262,In_1651,In_1751);
nand U2263 (N_2263,In_2145,In_956);
nor U2264 (N_2264,In_1017,In_1880);
xnor U2265 (N_2265,In_760,In_699);
nor U2266 (N_2266,In_1174,In_1436);
xor U2267 (N_2267,In_2478,In_1702);
nand U2268 (N_2268,In_1351,In_2373);
nand U2269 (N_2269,In_1614,In_1076);
and U2270 (N_2270,In_2098,In_1697);
nand U2271 (N_2271,In_977,In_2320);
nand U2272 (N_2272,In_1480,In_80);
xnor U2273 (N_2273,In_1523,In_81);
nand U2274 (N_2274,In_1676,In_749);
nor U2275 (N_2275,In_316,In_1647);
or U2276 (N_2276,In_843,In_904);
and U2277 (N_2277,In_1133,In_230);
nor U2278 (N_2278,In_1695,In_2445);
nand U2279 (N_2279,In_1362,In_1287);
nand U2280 (N_2280,In_126,In_300);
or U2281 (N_2281,In_57,In_1994);
xor U2282 (N_2282,In_1122,In_2304);
or U2283 (N_2283,In_2184,In_944);
nor U2284 (N_2284,In_1078,In_1164);
nand U2285 (N_2285,In_1899,In_804);
and U2286 (N_2286,In_2443,In_1151);
nand U2287 (N_2287,In_760,In_278);
nor U2288 (N_2288,In_152,In_1689);
nor U2289 (N_2289,In_2236,In_2399);
nor U2290 (N_2290,In_38,In_1756);
nor U2291 (N_2291,In_1188,In_1400);
nand U2292 (N_2292,In_2154,In_371);
xor U2293 (N_2293,In_1977,In_1540);
xnor U2294 (N_2294,In_2414,In_1448);
and U2295 (N_2295,In_2353,In_1258);
nand U2296 (N_2296,In_2034,In_341);
nand U2297 (N_2297,In_268,In_965);
xnor U2298 (N_2298,In_1197,In_626);
xor U2299 (N_2299,In_1874,In_2434);
or U2300 (N_2300,In_424,In_1955);
nand U2301 (N_2301,In_2229,In_97);
nor U2302 (N_2302,In_504,In_1345);
or U2303 (N_2303,In_1968,In_1780);
nand U2304 (N_2304,In_2460,In_1843);
or U2305 (N_2305,In_2220,In_537);
and U2306 (N_2306,In_784,In_702);
and U2307 (N_2307,In_672,In_1159);
nor U2308 (N_2308,In_1920,In_458);
or U2309 (N_2309,In_573,In_603);
xor U2310 (N_2310,In_639,In_29);
nand U2311 (N_2311,In_2455,In_1342);
or U2312 (N_2312,In_262,In_701);
nand U2313 (N_2313,In_2087,In_401);
nor U2314 (N_2314,In_455,In_569);
or U2315 (N_2315,In_2124,In_1282);
and U2316 (N_2316,In_431,In_1965);
and U2317 (N_2317,In_204,In_2047);
or U2318 (N_2318,In_1384,In_652);
nand U2319 (N_2319,In_1545,In_2482);
xor U2320 (N_2320,In_1519,In_1840);
nor U2321 (N_2321,In_627,In_2023);
or U2322 (N_2322,In_390,In_282);
and U2323 (N_2323,In_1400,In_1410);
nand U2324 (N_2324,In_2244,In_710);
xnor U2325 (N_2325,In_1252,In_1253);
nor U2326 (N_2326,In_231,In_2378);
or U2327 (N_2327,In_2399,In_885);
or U2328 (N_2328,In_1663,In_784);
nor U2329 (N_2329,In_1852,In_1635);
or U2330 (N_2330,In_1807,In_1604);
nand U2331 (N_2331,In_424,In_2444);
nand U2332 (N_2332,In_1814,In_1018);
or U2333 (N_2333,In_2356,In_1365);
xnor U2334 (N_2334,In_1065,In_1584);
or U2335 (N_2335,In_511,In_1563);
nor U2336 (N_2336,In_359,In_1229);
nor U2337 (N_2337,In_1523,In_1321);
nor U2338 (N_2338,In_1686,In_32);
nand U2339 (N_2339,In_25,In_144);
nand U2340 (N_2340,In_1097,In_1093);
or U2341 (N_2341,In_607,In_936);
nor U2342 (N_2342,In_1632,In_1559);
and U2343 (N_2343,In_2099,In_1789);
nor U2344 (N_2344,In_1774,In_1317);
and U2345 (N_2345,In_1884,In_2226);
nor U2346 (N_2346,In_2482,In_90);
xnor U2347 (N_2347,In_1505,In_1600);
nor U2348 (N_2348,In_125,In_374);
and U2349 (N_2349,In_2063,In_1091);
and U2350 (N_2350,In_1345,In_1448);
or U2351 (N_2351,In_954,In_685);
xor U2352 (N_2352,In_773,In_221);
nor U2353 (N_2353,In_1478,In_338);
xnor U2354 (N_2354,In_1081,In_1335);
and U2355 (N_2355,In_1207,In_1687);
or U2356 (N_2356,In_1013,In_461);
or U2357 (N_2357,In_1310,In_543);
nand U2358 (N_2358,In_925,In_1078);
or U2359 (N_2359,In_292,In_1201);
xnor U2360 (N_2360,In_407,In_12);
nand U2361 (N_2361,In_526,In_518);
and U2362 (N_2362,In_1441,In_1903);
nor U2363 (N_2363,In_1633,In_404);
nor U2364 (N_2364,In_365,In_2476);
nand U2365 (N_2365,In_572,In_1766);
xor U2366 (N_2366,In_1428,In_2035);
xor U2367 (N_2367,In_1319,In_1839);
nand U2368 (N_2368,In_1178,In_476);
xnor U2369 (N_2369,In_2291,In_1280);
nor U2370 (N_2370,In_2057,In_1193);
xnor U2371 (N_2371,In_534,In_842);
xor U2372 (N_2372,In_215,In_2400);
nand U2373 (N_2373,In_1573,In_429);
nand U2374 (N_2374,In_1982,In_2253);
nor U2375 (N_2375,In_447,In_2358);
nand U2376 (N_2376,In_938,In_558);
xnor U2377 (N_2377,In_2438,In_2092);
xor U2378 (N_2378,In_853,In_388);
nand U2379 (N_2379,In_247,In_1364);
xnor U2380 (N_2380,In_1374,In_1052);
nand U2381 (N_2381,In_2367,In_538);
and U2382 (N_2382,In_703,In_54);
or U2383 (N_2383,In_215,In_886);
or U2384 (N_2384,In_1512,In_563);
and U2385 (N_2385,In_1856,In_2064);
nand U2386 (N_2386,In_1622,In_484);
xor U2387 (N_2387,In_1968,In_2129);
and U2388 (N_2388,In_425,In_1816);
nor U2389 (N_2389,In_2150,In_1253);
and U2390 (N_2390,In_2131,In_1832);
and U2391 (N_2391,In_1268,In_1810);
or U2392 (N_2392,In_628,In_1889);
and U2393 (N_2393,In_1762,In_1070);
xor U2394 (N_2394,In_1977,In_2399);
and U2395 (N_2395,In_1784,In_1537);
or U2396 (N_2396,In_1185,In_2165);
xnor U2397 (N_2397,In_890,In_715);
nand U2398 (N_2398,In_437,In_1394);
xnor U2399 (N_2399,In_2310,In_1676);
and U2400 (N_2400,In_511,In_89);
and U2401 (N_2401,In_585,In_605);
and U2402 (N_2402,In_890,In_1973);
nand U2403 (N_2403,In_493,In_2271);
xnor U2404 (N_2404,In_781,In_1489);
xor U2405 (N_2405,In_0,In_363);
or U2406 (N_2406,In_2300,In_2471);
nand U2407 (N_2407,In_605,In_362);
nand U2408 (N_2408,In_1102,In_1064);
and U2409 (N_2409,In_910,In_1434);
and U2410 (N_2410,In_78,In_1179);
and U2411 (N_2411,In_2324,In_1184);
xor U2412 (N_2412,In_920,In_996);
nor U2413 (N_2413,In_1925,In_512);
and U2414 (N_2414,In_1897,In_1300);
xnor U2415 (N_2415,In_221,In_138);
xnor U2416 (N_2416,In_872,In_248);
nor U2417 (N_2417,In_347,In_459);
nand U2418 (N_2418,In_314,In_68);
and U2419 (N_2419,In_1460,In_1108);
nor U2420 (N_2420,In_1281,In_2194);
or U2421 (N_2421,In_1055,In_708);
or U2422 (N_2422,In_2440,In_2286);
xor U2423 (N_2423,In_2025,In_1281);
nand U2424 (N_2424,In_472,In_1553);
nand U2425 (N_2425,In_1162,In_1392);
xor U2426 (N_2426,In_184,In_1209);
nor U2427 (N_2427,In_2184,In_1728);
xor U2428 (N_2428,In_755,In_2171);
xnor U2429 (N_2429,In_1751,In_1772);
or U2430 (N_2430,In_1027,In_901);
and U2431 (N_2431,In_73,In_959);
xnor U2432 (N_2432,In_2304,In_655);
xnor U2433 (N_2433,In_2202,In_2463);
nor U2434 (N_2434,In_2269,In_171);
nand U2435 (N_2435,In_1304,In_647);
and U2436 (N_2436,In_636,In_1387);
or U2437 (N_2437,In_318,In_1677);
or U2438 (N_2438,In_1116,In_2353);
nor U2439 (N_2439,In_769,In_951);
nand U2440 (N_2440,In_975,In_1936);
and U2441 (N_2441,In_73,In_577);
xnor U2442 (N_2442,In_283,In_479);
xnor U2443 (N_2443,In_1736,In_42);
nand U2444 (N_2444,In_2246,In_796);
xnor U2445 (N_2445,In_1189,In_1383);
nand U2446 (N_2446,In_1243,In_1233);
nor U2447 (N_2447,In_357,In_4);
nand U2448 (N_2448,In_117,In_669);
nor U2449 (N_2449,In_1233,In_717);
and U2450 (N_2450,In_2193,In_560);
nand U2451 (N_2451,In_470,In_62);
xor U2452 (N_2452,In_2219,In_2403);
or U2453 (N_2453,In_643,In_2175);
xor U2454 (N_2454,In_1394,In_1326);
nand U2455 (N_2455,In_1329,In_1448);
or U2456 (N_2456,In_574,In_1242);
and U2457 (N_2457,In_2019,In_2313);
nand U2458 (N_2458,In_1699,In_2390);
xor U2459 (N_2459,In_713,In_1012);
and U2460 (N_2460,In_1128,In_1082);
nand U2461 (N_2461,In_1436,In_36);
nor U2462 (N_2462,In_334,In_1796);
nor U2463 (N_2463,In_1404,In_205);
xnor U2464 (N_2464,In_42,In_1240);
nand U2465 (N_2465,In_985,In_1641);
nor U2466 (N_2466,In_926,In_2090);
nand U2467 (N_2467,In_378,In_610);
and U2468 (N_2468,In_84,In_1973);
xor U2469 (N_2469,In_320,In_5);
xnor U2470 (N_2470,In_2,In_541);
or U2471 (N_2471,In_749,In_896);
or U2472 (N_2472,In_913,In_229);
nor U2473 (N_2473,In_305,In_1337);
nor U2474 (N_2474,In_1090,In_2175);
or U2475 (N_2475,In_2329,In_1527);
or U2476 (N_2476,In_2353,In_858);
xor U2477 (N_2477,In_234,In_1269);
nor U2478 (N_2478,In_14,In_1140);
or U2479 (N_2479,In_878,In_398);
nand U2480 (N_2480,In_1377,In_1090);
and U2481 (N_2481,In_157,In_1362);
nand U2482 (N_2482,In_686,In_533);
or U2483 (N_2483,In_1346,In_2048);
nand U2484 (N_2484,In_862,In_918);
nor U2485 (N_2485,In_1764,In_1275);
nand U2486 (N_2486,In_193,In_1116);
or U2487 (N_2487,In_1742,In_2346);
and U2488 (N_2488,In_2015,In_1305);
nor U2489 (N_2489,In_2426,In_1317);
nor U2490 (N_2490,In_1590,In_561);
nand U2491 (N_2491,In_2241,In_771);
nand U2492 (N_2492,In_1218,In_2050);
or U2493 (N_2493,In_1582,In_1863);
xor U2494 (N_2494,In_22,In_1334);
xor U2495 (N_2495,In_2485,In_1917);
xnor U2496 (N_2496,In_1877,In_1141);
nor U2497 (N_2497,In_1757,In_889);
xor U2498 (N_2498,In_990,In_364);
nand U2499 (N_2499,In_820,In_81);
nand U2500 (N_2500,In_289,In_2080);
nor U2501 (N_2501,In_1165,In_2299);
xnor U2502 (N_2502,In_804,In_1673);
nor U2503 (N_2503,In_2251,In_293);
nor U2504 (N_2504,In_404,In_1128);
nor U2505 (N_2505,In_307,In_1083);
or U2506 (N_2506,In_1942,In_1948);
xnor U2507 (N_2507,In_1264,In_1533);
xnor U2508 (N_2508,In_2046,In_1422);
nor U2509 (N_2509,In_1579,In_1559);
or U2510 (N_2510,In_1026,In_2394);
nand U2511 (N_2511,In_1205,In_842);
nand U2512 (N_2512,In_2212,In_39);
or U2513 (N_2513,In_1158,In_173);
nor U2514 (N_2514,In_620,In_776);
nand U2515 (N_2515,In_1828,In_904);
xor U2516 (N_2516,In_834,In_262);
or U2517 (N_2517,In_619,In_2345);
nand U2518 (N_2518,In_64,In_1933);
and U2519 (N_2519,In_1270,In_1709);
or U2520 (N_2520,In_1848,In_1784);
nor U2521 (N_2521,In_1480,In_112);
xnor U2522 (N_2522,In_1371,In_657);
xnor U2523 (N_2523,In_1666,In_1369);
and U2524 (N_2524,In_2365,In_1387);
nand U2525 (N_2525,In_486,In_91);
nor U2526 (N_2526,In_1407,In_1637);
or U2527 (N_2527,In_1360,In_1652);
and U2528 (N_2528,In_2111,In_871);
xnor U2529 (N_2529,In_1231,In_2483);
nor U2530 (N_2530,In_1079,In_2372);
nor U2531 (N_2531,In_1077,In_756);
or U2532 (N_2532,In_2338,In_863);
and U2533 (N_2533,In_2000,In_2349);
or U2534 (N_2534,In_2444,In_1408);
or U2535 (N_2535,In_2325,In_463);
and U2536 (N_2536,In_183,In_2133);
nor U2537 (N_2537,In_925,In_1732);
xor U2538 (N_2538,In_1770,In_249);
xor U2539 (N_2539,In_1057,In_1779);
nand U2540 (N_2540,In_189,In_1005);
nand U2541 (N_2541,In_1997,In_222);
and U2542 (N_2542,In_1278,In_209);
nor U2543 (N_2543,In_1570,In_2280);
and U2544 (N_2544,In_1598,In_1100);
nand U2545 (N_2545,In_190,In_74);
or U2546 (N_2546,In_512,In_1418);
or U2547 (N_2547,In_2365,In_910);
nor U2548 (N_2548,In_1692,In_1607);
and U2549 (N_2549,In_2064,In_569);
xor U2550 (N_2550,In_240,In_1006);
or U2551 (N_2551,In_1290,In_554);
or U2552 (N_2552,In_2447,In_1662);
or U2553 (N_2553,In_1369,In_249);
nor U2554 (N_2554,In_1492,In_2455);
nand U2555 (N_2555,In_50,In_1914);
or U2556 (N_2556,In_1635,In_2168);
xnor U2557 (N_2557,In_1278,In_110);
or U2558 (N_2558,In_1240,In_1955);
xnor U2559 (N_2559,In_34,In_1456);
nand U2560 (N_2560,In_868,In_2370);
and U2561 (N_2561,In_2498,In_1173);
nand U2562 (N_2562,In_1817,In_1731);
nand U2563 (N_2563,In_142,In_930);
nand U2564 (N_2564,In_2272,In_2251);
and U2565 (N_2565,In_2492,In_1571);
and U2566 (N_2566,In_2464,In_915);
and U2567 (N_2567,In_1169,In_399);
nand U2568 (N_2568,In_186,In_1627);
or U2569 (N_2569,In_2262,In_1377);
nor U2570 (N_2570,In_694,In_1608);
or U2571 (N_2571,In_1011,In_519);
nor U2572 (N_2572,In_1938,In_212);
and U2573 (N_2573,In_1567,In_1587);
nor U2574 (N_2574,In_141,In_2301);
or U2575 (N_2575,In_1567,In_1001);
or U2576 (N_2576,In_370,In_1200);
nor U2577 (N_2577,In_447,In_1445);
xnor U2578 (N_2578,In_1239,In_1672);
and U2579 (N_2579,In_2116,In_2220);
or U2580 (N_2580,In_2037,In_838);
nand U2581 (N_2581,In_261,In_1196);
and U2582 (N_2582,In_582,In_1059);
or U2583 (N_2583,In_625,In_802);
xnor U2584 (N_2584,In_910,In_664);
nor U2585 (N_2585,In_345,In_810);
nor U2586 (N_2586,In_1011,In_1012);
and U2587 (N_2587,In_1672,In_136);
or U2588 (N_2588,In_1698,In_1119);
nand U2589 (N_2589,In_633,In_1772);
xnor U2590 (N_2590,In_1748,In_2079);
or U2591 (N_2591,In_698,In_829);
nor U2592 (N_2592,In_1642,In_1449);
or U2593 (N_2593,In_1169,In_2100);
nor U2594 (N_2594,In_959,In_100);
nor U2595 (N_2595,In_2124,In_1188);
xnor U2596 (N_2596,In_770,In_2110);
nand U2597 (N_2597,In_1546,In_273);
nand U2598 (N_2598,In_1680,In_63);
nand U2599 (N_2599,In_2191,In_828);
nand U2600 (N_2600,In_2155,In_626);
and U2601 (N_2601,In_2426,In_1984);
nand U2602 (N_2602,In_2065,In_630);
xnor U2603 (N_2603,In_634,In_1730);
nand U2604 (N_2604,In_1475,In_58);
nor U2605 (N_2605,In_379,In_3);
nor U2606 (N_2606,In_722,In_2059);
and U2607 (N_2607,In_1752,In_1016);
nand U2608 (N_2608,In_2305,In_580);
xnor U2609 (N_2609,In_797,In_993);
or U2610 (N_2610,In_408,In_2415);
nand U2611 (N_2611,In_1535,In_1370);
xnor U2612 (N_2612,In_2228,In_2046);
nand U2613 (N_2613,In_2065,In_1808);
and U2614 (N_2614,In_2482,In_863);
nor U2615 (N_2615,In_2339,In_2149);
or U2616 (N_2616,In_1382,In_832);
or U2617 (N_2617,In_2083,In_1341);
xnor U2618 (N_2618,In_2423,In_1098);
or U2619 (N_2619,In_2127,In_36);
or U2620 (N_2620,In_201,In_2447);
nor U2621 (N_2621,In_318,In_1502);
or U2622 (N_2622,In_1698,In_152);
nand U2623 (N_2623,In_346,In_331);
xnor U2624 (N_2624,In_206,In_2390);
xnor U2625 (N_2625,In_19,In_1667);
or U2626 (N_2626,In_2092,In_225);
and U2627 (N_2627,In_1506,In_616);
or U2628 (N_2628,In_467,In_1710);
or U2629 (N_2629,In_2424,In_1137);
nor U2630 (N_2630,In_2174,In_529);
nand U2631 (N_2631,In_1221,In_1858);
and U2632 (N_2632,In_1402,In_1083);
nand U2633 (N_2633,In_552,In_2376);
xor U2634 (N_2634,In_2429,In_1814);
nand U2635 (N_2635,In_562,In_338);
nand U2636 (N_2636,In_2268,In_126);
or U2637 (N_2637,In_846,In_1653);
nand U2638 (N_2638,In_1593,In_2230);
nor U2639 (N_2639,In_601,In_555);
xnor U2640 (N_2640,In_314,In_431);
nor U2641 (N_2641,In_1994,In_766);
nor U2642 (N_2642,In_159,In_1297);
and U2643 (N_2643,In_1805,In_2280);
nand U2644 (N_2644,In_1384,In_1310);
and U2645 (N_2645,In_873,In_2371);
nor U2646 (N_2646,In_1655,In_651);
or U2647 (N_2647,In_1123,In_2366);
or U2648 (N_2648,In_1719,In_2461);
and U2649 (N_2649,In_649,In_2300);
nor U2650 (N_2650,In_2251,In_2405);
or U2651 (N_2651,In_2038,In_645);
xor U2652 (N_2652,In_2079,In_1199);
xor U2653 (N_2653,In_477,In_1357);
nor U2654 (N_2654,In_795,In_402);
or U2655 (N_2655,In_2221,In_704);
xor U2656 (N_2656,In_139,In_1648);
and U2657 (N_2657,In_1885,In_1546);
and U2658 (N_2658,In_866,In_1034);
nor U2659 (N_2659,In_1309,In_519);
xnor U2660 (N_2660,In_2209,In_778);
or U2661 (N_2661,In_339,In_1088);
or U2662 (N_2662,In_986,In_337);
nor U2663 (N_2663,In_1031,In_1624);
nor U2664 (N_2664,In_1188,In_440);
and U2665 (N_2665,In_2266,In_103);
and U2666 (N_2666,In_750,In_1197);
nand U2667 (N_2667,In_2194,In_311);
xor U2668 (N_2668,In_583,In_431);
or U2669 (N_2669,In_1364,In_336);
nor U2670 (N_2670,In_524,In_1179);
and U2671 (N_2671,In_1927,In_1346);
and U2672 (N_2672,In_510,In_1159);
xor U2673 (N_2673,In_2118,In_758);
and U2674 (N_2674,In_1873,In_72);
or U2675 (N_2675,In_614,In_178);
and U2676 (N_2676,In_323,In_1349);
and U2677 (N_2677,In_2407,In_1312);
nand U2678 (N_2678,In_1002,In_1591);
and U2679 (N_2679,In_2084,In_671);
xnor U2680 (N_2680,In_1275,In_2125);
and U2681 (N_2681,In_845,In_323);
and U2682 (N_2682,In_1870,In_1137);
and U2683 (N_2683,In_269,In_1662);
nand U2684 (N_2684,In_1744,In_588);
and U2685 (N_2685,In_2313,In_2178);
xnor U2686 (N_2686,In_2248,In_1489);
nor U2687 (N_2687,In_351,In_731);
or U2688 (N_2688,In_681,In_1394);
nand U2689 (N_2689,In_1632,In_1715);
and U2690 (N_2690,In_1311,In_2390);
nor U2691 (N_2691,In_782,In_1325);
nand U2692 (N_2692,In_2234,In_1030);
and U2693 (N_2693,In_315,In_1495);
or U2694 (N_2694,In_253,In_1055);
nand U2695 (N_2695,In_1951,In_1760);
nand U2696 (N_2696,In_985,In_1342);
xnor U2697 (N_2697,In_723,In_317);
and U2698 (N_2698,In_1497,In_1393);
nand U2699 (N_2699,In_2368,In_53);
nor U2700 (N_2700,In_391,In_964);
nand U2701 (N_2701,In_966,In_360);
nand U2702 (N_2702,In_2016,In_83);
xor U2703 (N_2703,In_1884,In_2314);
and U2704 (N_2704,In_2126,In_1738);
nand U2705 (N_2705,In_10,In_2005);
xnor U2706 (N_2706,In_2029,In_1114);
and U2707 (N_2707,In_59,In_2358);
and U2708 (N_2708,In_1063,In_2180);
or U2709 (N_2709,In_1219,In_1454);
nand U2710 (N_2710,In_183,In_256);
xor U2711 (N_2711,In_2235,In_1760);
xor U2712 (N_2712,In_708,In_1854);
nand U2713 (N_2713,In_1403,In_2210);
nor U2714 (N_2714,In_1145,In_684);
and U2715 (N_2715,In_1082,In_2419);
xnor U2716 (N_2716,In_1653,In_1616);
or U2717 (N_2717,In_911,In_2187);
xnor U2718 (N_2718,In_2124,In_2183);
nor U2719 (N_2719,In_820,In_1);
nor U2720 (N_2720,In_1572,In_61);
or U2721 (N_2721,In_2011,In_1230);
or U2722 (N_2722,In_1864,In_1832);
nand U2723 (N_2723,In_1705,In_1962);
and U2724 (N_2724,In_1202,In_511);
xnor U2725 (N_2725,In_1312,In_23);
xnor U2726 (N_2726,In_1767,In_725);
and U2727 (N_2727,In_2143,In_1902);
and U2728 (N_2728,In_2331,In_2375);
or U2729 (N_2729,In_2322,In_207);
xnor U2730 (N_2730,In_1726,In_1915);
nand U2731 (N_2731,In_1454,In_1779);
and U2732 (N_2732,In_1793,In_79);
nor U2733 (N_2733,In_564,In_2419);
nand U2734 (N_2734,In_1007,In_1255);
nand U2735 (N_2735,In_2409,In_87);
or U2736 (N_2736,In_1473,In_2024);
or U2737 (N_2737,In_2401,In_396);
and U2738 (N_2738,In_1316,In_691);
nor U2739 (N_2739,In_2401,In_1814);
or U2740 (N_2740,In_919,In_1419);
nand U2741 (N_2741,In_818,In_2357);
or U2742 (N_2742,In_1104,In_1715);
nand U2743 (N_2743,In_1943,In_1952);
xnor U2744 (N_2744,In_984,In_2416);
xnor U2745 (N_2745,In_2213,In_2102);
nor U2746 (N_2746,In_200,In_1221);
or U2747 (N_2747,In_1838,In_116);
nor U2748 (N_2748,In_1609,In_840);
nor U2749 (N_2749,In_1489,In_239);
nor U2750 (N_2750,In_495,In_1495);
xor U2751 (N_2751,In_356,In_1222);
nor U2752 (N_2752,In_38,In_28);
nand U2753 (N_2753,In_1544,In_1422);
nand U2754 (N_2754,In_1959,In_1102);
or U2755 (N_2755,In_1521,In_1738);
or U2756 (N_2756,In_1457,In_730);
and U2757 (N_2757,In_6,In_285);
nand U2758 (N_2758,In_907,In_1068);
xor U2759 (N_2759,In_801,In_2416);
and U2760 (N_2760,In_307,In_2161);
xnor U2761 (N_2761,In_196,In_1506);
or U2762 (N_2762,In_1241,In_2301);
or U2763 (N_2763,In_1353,In_1372);
or U2764 (N_2764,In_1086,In_1053);
xor U2765 (N_2765,In_1632,In_2297);
xor U2766 (N_2766,In_247,In_207);
xnor U2767 (N_2767,In_2092,In_787);
or U2768 (N_2768,In_978,In_1624);
nand U2769 (N_2769,In_1597,In_1508);
or U2770 (N_2770,In_1789,In_1480);
nand U2771 (N_2771,In_473,In_1806);
and U2772 (N_2772,In_2428,In_382);
or U2773 (N_2773,In_634,In_1183);
nand U2774 (N_2774,In_607,In_299);
nor U2775 (N_2775,In_2146,In_949);
and U2776 (N_2776,In_995,In_803);
xnor U2777 (N_2777,In_970,In_1319);
nor U2778 (N_2778,In_444,In_1419);
or U2779 (N_2779,In_653,In_1303);
xor U2780 (N_2780,In_1591,In_386);
or U2781 (N_2781,In_2326,In_57);
xnor U2782 (N_2782,In_284,In_1241);
nor U2783 (N_2783,In_2438,In_1842);
or U2784 (N_2784,In_567,In_930);
nor U2785 (N_2785,In_1773,In_1173);
nand U2786 (N_2786,In_1049,In_392);
and U2787 (N_2787,In_688,In_2135);
nor U2788 (N_2788,In_1930,In_2099);
xnor U2789 (N_2789,In_305,In_1420);
or U2790 (N_2790,In_1716,In_1861);
nor U2791 (N_2791,In_811,In_1371);
nand U2792 (N_2792,In_605,In_1768);
and U2793 (N_2793,In_325,In_1017);
and U2794 (N_2794,In_505,In_42);
nand U2795 (N_2795,In_2023,In_1234);
xor U2796 (N_2796,In_1433,In_465);
xnor U2797 (N_2797,In_2389,In_356);
xor U2798 (N_2798,In_1890,In_393);
or U2799 (N_2799,In_1329,In_693);
and U2800 (N_2800,In_2348,In_2251);
nor U2801 (N_2801,In_2482,In_2409);
or U2802 (N_2802,In_504,In_129);
nor U2803 (N_2803,In_334,In_229);
or U2804 (N_2804,In_1183,In_2342);
or U2805 (N_2805,In_898,In_526);
xor U2806 (N_2806,In_252,In_2140);
nand U2807 (N_2807,In_712,In_1390);
xnor U2808 (N_2808,In_907,In_1144);
nand U2809 (N_2809,In_800,In_1480);
nand U2810 (N_2810,In_2492,In_2058);
or U2811 (N_2811,In_2040,In_2094);
nand U2812 (N_2812,In_2371,In_140);
xnor U2813 (N_2813,In_903,In_206);
nor U2814 (N_2814,In_2488,In_2387);
or U2815 (N_2815,In_2036,In_469);
nand U2816 (N_2816,In_2129,In_2382);
nand U2817 (N_2817,In_330,In_698);
xor U2818 (N_2818,In_1007,In_1518);
or U2819 (N_2819,In_890,In_897);
nor U2820 (N_2820,In_211,In_1339);
nor U2821 (N_2821,In_2461,In_901);
nand U2822 (N_2822,In_708,In_2317);
nand U2823 (N_2823,In_1316,In_25);
and U2824 (N_2824,In_1564,In_1166);
xnor U2825 (N_2825,In_2050,In_2270);
or U2826 (N_2826,In_1030,In_937);
nor U2827 (N_2827,In_1550,In_503);
xor U2828 (N_2828,In_2380,In_440);
nor U2829 (N_2829,In_1385,In_1140);
nor U2830 (N_2830,In_1297,In_15);
xnor U2831 (N_2831,In_1934,In_1534);
xnor U2832 (N_2832,In_1144,In_1261);
or U2833 (N_2833,In_2250,In_432);
nor U2834 (N_2834,In_2356,In_104);
nand U2835 (N_2835,In_2414,In_1378);
xnor U2836 (N_2836,In_590,In_498);
or U2837 (N_2837,In_1009,In_2244);
nand U2838 (N_2838,In_1372,In_1564);
nand U2839 (N_2839,In_1684,In_1891);
and U2840 (N_2840,In_344,In_1343);
or U2841 (N_2841,In_934,In_1491);
nand U2842 (N_2842,In_1999,In_1197);
and U2843 (N_2843,In_2148,In_762);
nor U2844 (N_2844,In_570,In_1808);
or U2845 (N_2845,In_2366,In_392);
xor U2846 (N_2846,In_80,In_2362);
or U2847 (N_2847,In_1720,In_246);
nor U2848 (N_2848,In_987,In_371);
nor U2849 (N_2849,In_229,In_1993);
and U2850 (N_2850,In_2479,In_2156);
nor U2851 (N_2851,In_433,In_1810);
xnor U2852 (N_2852,In_76,In_16);
nor U2853 (N_2853,In_1206,In_540);
and U2854 (N_2854,In_165,In_2371);
nor U2855 (N_2855,In_1754,In_322);
xor U2856 (N_2856,In_488,In_594);
and U2857 (N_2857,In_1276,In_807);
xor U2858 (N_2858,In_1264,In_2389);
nand U2859 (N_2859,In_1176,In_2380);
or U2860 (N_2860,In_1341,In_668);
and U2861 (N_2861,In_1559,In_624);
nor U2862 (N_2862,In_359,In_28);
nor U2863 (N_2863,In_178,In_892);
nand U2864 (N_2864,In_533,In_24);
or U2865 (N_2865,In_679,In_2498);
xor U2866 (N_2866,In_433,In_1117);
xnor U2867 (N_2867,In_948,In_47);
and U2868 (N_2868,In_534,In_1955);
nor U2869 (N_2869,In_170,In_2247);
nor U2870 (N_2870,In_988,In_820);
xnor U2871 (N_2871,In_226,In_2283);
nor U2872 (N_2872,In_926,In_2480);
nor U2873 (N_2873,In_1379,In_458);
or U2874 (N_2874,In_937,In_1747);
or U2875 (N_2875,In_2127,In_1190);
and U2876 (N_2876,In_179,In_1663);
xor U2877 (N_2877,In_486,In_1506);
and U2878 (N_2878,In_1956,In_1677);
and U2879 (N_2879,In_2414,In_793);
nand U2880 (N_2880,In_2213,In_825);
nor U2881 (N_2881,In_639,In_897);
nand U2882 (N_2882,In_1309,In_1444);
xor U2883 (N_2883,In_1318,In_1494);
xor U2884 (N_2884,In_639,In_128);
nand U2885 (N_2885,In_744,In_119);
or U2886 (N_2886,In_131,In_1277);
nor U2887 (N_2887,In_183,In_2443);
xor U2888 (N_2888,In_669,In_1705);
xor U2889 (N_2889,In_290,In_1460);
or U2890 (N_2890,In_692,In_456);
xor U2891 (N_2891,In_1122,In_1557);
or U2892 (N_2892,In_1703,In_1429);
or U2893 (N_2893,In_1886,In_1230);
xor U2894 (N_2894,In_322,In_248);
nor U2895 (N_2895,In_1499,In_1657);
nor U2896 (N_2896,In_1656,In_1403);
or U2897 (N_2897,In_462,In_1542);
nor U2898 (N_2898,In_281,In_1834);
nand U2899 (N_2899,In_2111,In_169);
or U2900 (N_2900,In_1337,In_2160);
nand U2901 (N_2901,In_2262,In_1214);
xor U2902 (N_2902,In_1631,In_2285);
nor U2903 (N_2903,In_1020,In_1856);
and U2904 (N_2904,In_731,In_2316);
nand U2905 (N_2905,In_974,In_1364);
or U2906 (N_2906,In_2118,In_1335);
nor U2907 (N_2907,In_239,In_888);
xor U2908 (N_2908,In_778,In_1979);
or U2909 (N_2909,In_664,In_2392);
nand U2910 (N_2910,In_73,In_1461);
xor U2911 (N_2911,In_1575,In_225);
xor U2912 (N_2912,In_1133,In_1950);
and U2913 (N_2913,In_1362,In_826);
nor U2914 (N_2914,In_1007,In_2157);
and U2915 (N_2915,In_1604,In_318);
nand U2916 (N_2916,In_1489,In_1082);
nor U2917 (N_2917,In_1394,In_2308);
and U2918 (N_2918,In_374,In_650);
nor U2919 (N_2919,In_1280,In_164);
nor U2920 (N_2920,In_746,In_905);
and U2921 (N_2921,In_544,In_1298);
or U2922 (N_2922,In_2428,In_355);
xor U2923 (N_2923,In_1294,In_1084);
nand U2924 (N_2924,In_835,In_2082);
nor U2925 (N_2925,In_1421,In_2214);
nor U2926 (N_2926,In_1502,In_574);
or U2927 (N_2927,In_1634,In_179);
nor U2928 (N_2928,In_660,In_129);
nand U2929 (N_2929,In_1482,In_1193);
and U2930 (N_2930,In_1349,In_2320);
nor U2931 (N_2931,In_888,In_762);
xnor U2932 (N_2932,In_2082,In_1939);
nand U2933 (N_2933,In_1157,In_1072);
and U2934 (N_2934,In_2344,In_214);
nand U2935 (N_2935,In_2220,In_21);
or U2936 (N_2936,In_1201,In_90);
xor U2937 (N_2937,In_790,In_1144);
and U2938 (N_2938,In_2146,In_135);
nand U2939 (N_2939,In_797,In_2128);
xor U2940 (N_2940,In_815,In_991);
nand U2941 (N_2941,In_344,In_107);
xor U2942 (N_2942,In_2076,In_1051);
or U2943 (N_2943,In_1015,In_2052);
and U2944 (N_2944,In_989,In_1340);
nor U2945 (N_2945,In_1908,In_1613);
nand U2946 (N_2946,In_58,In_1613);
xnor U2947 (N_2947,In_1292,In_553);
and U2948 (N_2948,In_1061,In_363);
xnor U2949 (N_2949,In_1454,In_494);
xor U2950 (N_2950,In_2110,In_254);
nand U2951 (N_2951,In_536,In_276);
and U2952 (N_2952,In_603,In_617);
nand U2953 (N_2953,In_523,In_2343);
xnor U2954 (N_2954,In_1281,In_2100);
and U2955 (N_2955,In_2219,In_726);
or U2956 (N_2956,In_1332,In_2281);
xor U2957 (N_2957,In_1087,In_732);
and U2958 (N_2958,In_451,In_35);
xor U2959 (N_2959,In_82,In_984);
or U2960 (N_2960,In_818,In_532);
and U2961 (N_2961,In_1942,In_865);
or U2962 (N_2962,In_2264,In_2233);
and U2963 (N_2963,In_293,In_2355);
nor U2964 (N_2964,In_270,In_837);
nor U2965 (N_2965,In_1932,In_1931);
nand U2966 (N_2966,In_345,In_125);
and U2967 (N_2967,In_2052,In_862);
nand U2968 (N_2968,In_1649,In_564);
xor U2969 (N_2969,In_672,In_1531);
or U2970 (N_2970,In_1519,In_1780);
or U2971 (N_2971,In_348,In_61);
or U2972 (N_2972,In_2011,In_1763);
or U2973 (N_2973,In_835,In_2177);
or U2974 (N_2974,In_881,In_889);
or U2975 (N_2975,In_194,In_1680);
or U2976 (N_2976,In_1472,In_1728);
xor U2977 (N_2977,In_70,In_2088);
or U2978 (N_2978,In_1617,In_937);
nor U2979 (N_2979,In_513,In_1666);
xor U2980 (N_2980,In_1737,In_2339);
nor U2981 (N_2981,In_2343,In_1334);
or U2982 (N_2982,In_2138,In_749);
nor U2983 (N_2983,In_2343,In_604);
nand U2984 (N_2984,In_1100,In_803);
nor U2985 (N_2985,In_433,In_1683);
and U2986 (N_2986,In_1443,In_2035);
nor U2987 (N_2987,In_1438,In_141);
nand U2988 (N_2988,In_211,In_1116);
and U2989 (N_2989,In_8,In_2447);
nand U2990 (N_2990,In_626,In_1752);
xnor U2991 (N_2991,In_1681,In_366);
xnor U2992 (N_2992,In_1027,In_602);
and U2993 (N_2993,In_2090,In_1106);
nor U2994 (N_2994,In_1977,In_1899);
or U2995 (N_2995,In_430,In_1938);
and U2996 (N_2996,In_1216,In_657);
and U2997 (N_2997,In_2497,In_2197);
and U2998 (N_2998,In_125,In_2236);
nor U2999 (N_2999,In_527,In_506);
and U3000 (N_3000,In_2320,In_2358);
nor U3001 (N_3001,In_1043,In_2091);
nand U3002 (N_3002,In_1460,In_1743);
xnor U3003 (N_3003,In_746,In_1545);
or U3004 (N_3004,In_1293,In_80);
xnor U3005 (N_3005,In_1106,In_1059);
xnor U3006 (N_3006,In_730,In_299);
and U3007 (N_3007,In_1020,In_185);
nand U3008 (N_3008,In_1561,In_426);
xor U3009 (N_3009,In_1575,In_2116);
or U3010 (N_3010,In_2350,In_170);
nand U3011 (N_3011,In_1905,In_1278);
nand U3012 (N_3012,In_426,In_481);
and U3013 (N_3013,In_1818,In_1231);
xor U3014 (N_3014,In_501,In_1339);
nor U3015 (N_3015,In_1697,In_1853);
and U3016 (N_3016,In_204,In_986);
nand U3017 (N_3017,In_1795,In_1650);
and U3018 (N_3018,In_1491,In_1291);
and U3019 (N_3019,In_316,In_1264);
or U3020 (N_3020,In_1626,In_763);
or U3021 (N_3021,In_1836,In_1478);
nand U3022 (N_3022,In_1583,In_181);
and U3023 (N_3023,In_577,In_1541);
or U3024 (N_3024,In_204,In_1385);
nand U3025 (N_3025,In_2087,In_1264);
and U3026 (N_3026,In_2350,In_485);
xor U3027 (N_3027,In_1440,In_588);
xor U3028 (N_3028,In_2125,In_283);
or U3029 (N_3029,In_2169,In_1606);
or U3030 (N_3030,In_1541,In_1832);
and U3031 (N_3031,In_1171,In_1082);
or U3032 (N_3032,In_1029,In_657);
nor U3033 (N_3033,In_1184,In_1761);
nand U3034 (N_3034,In_1887,In_1660);
nor U3035 (N_3035,In_1426,In_1949);
and U3036 (N_3036,In_1545,In_668);
nor U3037 (N_3037,In_1558,In_2051);
and U3038 (N_3038,In_1954,In_2295);
nor U3039 (N_3039,In_327,In_257);
nand U3040 (N_3040,In_1275,In_1898);
and U3041 (N_3041,In_2051,In_1803);
and U3042 (N_3042,In_422,In_785);
xnor U3043 (N_3043,In_2401,In_1702);
or U3044 (N_3044,In_439,In_2435);
and U3045 (N_3045,In_367,In_1393);
xnor U3046 (N_3046,In_859,In_487);
or U3047 (N_3047,In_733,In_1932);
xor U3048 (N_3048,In_1089,In_1264);
nand U3049 (N_3049,In_836,In_2391);
and U3050 (N_3050,In_2338,In_894);
nand U3051 (N_3051,In_1568,In_1431);
xor U3052 (N_3052,In_2042,In_1365);
xnor U3053 (N_3053,In_142,In_1957);
nand U3054 (N_3054,In_543,In_1155);
or U3055 (N_3055,In_1000,In_1926);
xor U3056 (N_3056,In_1127,In_1748);
nor U3057 (N_3057,In_1296,In_1607);
or U3058 (N_3058,In_2329,In_2303);
nand U3059 (N_3059,In_329,In_2149);
or U3060 (N_3060,In_1410,In_663);
nor U3061 (N_3061,In_74,In_243);
nand U3062 (N_3062,In_657,In_231);
xnor U3063 (N_3063,In_518,In_271);
and U3064 (N_3064,In_2099,In_1587);
xnor U3065 (N_3065,In_2163,In_1711);
nor U3066 (N_3066,In_1012,In_1103);
or U3067 (N_3067,In_1073,In_1634);
and U3068 (N_3068,In_736,In_672);
xnor U3069 (N_3069,In_896,In_810);
nor U3070 (N_3070,In_602,In_1083);
or U3071 (N_3071,In_1320,In_2338);
or U3072 (N_3072,In_502,In_138);
xnor U3073 (N_3073,In_2210,In_456);
nand U3074 (N_3074,In_218,In_1885);
xnor U3075 (N_3075,In_292,In_1593);
or U3076 (N_3076,In_59,In_768);
and U3077 (N_3077,In_299,In_368);
xor U3078 (N_3078,In_1362,In_1871);
or U3079 (N_3079,In_2025,In_715);
nor U3080 (N_3080,In_2242,In_1745);
or U3081 (N_3081,In_338,In_2359);
xor U3082 (N_3082,In_1781,In_1675);
nor U3083 (N_3083,In_562,In_2372);
nor U3084 (N_3084,In_36,In_1380);
nand U3085 (N_3085,In_2038,In_2010);
nor U3086 (N_3086,In_1314,In_360);
xnor U3087 (N_3087,In_441,In_622);
or U3088 (N_3088,In_2236,In_1355);
nand U3089 (N_3089,In_1555,In_865);
nor U3090 (N_3090,In_378,In_2053);
and U3091 (N_3091,In_146,In_752);
and U3092 (N_3092,In_1682,In_138);
xnor U3093 (N_3093,In_414,In_564);
or U3094 (N_3094,In_1760,In_715);
and U3095 (N_3095,In_839,In_1898);
and U3096 (N_3096,In_2482,In_692);
and U3097 (N_3097,In_368,In_1113);
xnor U3098 (N_3098,In_768,In_361);
xnor U3099 (N_3099,In_1118,In_499);
and U3100 (N_3100,In_1588,In_1214);
or U3101 (N_3101,In_69,In_200);
or U3102 (N_3102,In_1926,In_1265);
xor U3103 (N_3103,In_1152,In_1844);
and U3104 (N_3104,In_1120,In_647);
or U3105 (N_3105,In_1838,In_1203);
xor U3106 (N_3106,In_356,In_962);
nor U3107 (N_3107,In_2055,In_1055);
or U3108 (N_3108,In_2177,In_2136);
or U3109 (N_3109,In_1663,In_2132);
nand U3110 (N_3110,In_143,In_1540);
nand U3111 (N_3111,In_2371,In_1910);
or U3112 (N_3112,In_1287,In_496);
nor U3113 (N_3113,In_512,In_1896);
nor U3114 (N_3114,In_2451,In_1798);
xor U3115 (N_3115,In_650,In_2422);
nand U3116 (N_3116,In_1257,In_1397);
or U3117 (N_3117,In_1459,In_627);
xor U3118 (N_3118,In_46,In_960);
or U3119 (N_3119,In_225,In_2422);
nand U3120 (N_3120,In_1039,In_206);
nand U3121 (N_3121,In_831,In_1270);
or U3122 (N_3122,In_2370,In_1311);
or U3123 (N_3123,In_1468,In_1196);
nand U3124 (N_3124,In_1251,In_1659);
xnor U3125 (N_3125,N_648,N_1029);
and U3126 (N_3126,N_2191,N_446);
and U3127 (N_3127,N_2112,N_2229);
and U3128 (N_3128,N_2896,N_2254);
or U3129 (N_3129,N_1284,N_1514);
or U3130 (N_3130,N_2716,N_2830);
and U3131 (N_3131,N_1585,N_2682);
or U3132 (N_3132,N_2624,N_2765);
and U3133 (N_3133,N_1248,N_325);
and U3134 (N_3134,N_2945,N_518);
and U3135 (N_3135,N_803,N_813);
nor U3136 (N_3136,N_1535,N_1543);
nand U3137 (N_3137,N_2573,N_2657);
nand U3138 (N_3138,N_1783,N_2640);
xnor U3139 (N_3139,N_658,N_1249);
nor U3140 (N_3140,N_2637,N_1297);
and U3141 (N_3141,N_2193,N_3043);
xor U3142 (N_3142,N_1207,N_2662);
and U3143 (N_3143,N_2769,N_958);
and U3144 (N_3144,N_2136,N_1409);
nor U3145 (N_3145,N_163,N_2722);
nor U3146 (N_3146,N_2151,N_370);
nand U3147 (N_3147,N_1961,N_72);
nand U3148 (N_3148,N_2788,N_2702);
or U3149 (N_3149,N_2060,N_1092);
and U3150 (N_3150,N_1583,N_1548);
and U3151 (N_3151,N_1194,N_988);
nand U3152 (N_3152,N_38,N_391);
or U3153 (N_3153,N_295,N_1550);
or U3154 (N_3154,N_206,N_2620);
nor U3155 (N_3155,N_1105,N_2921);
xnor U3156 (N_3156,N_1059,N_2403);
and U3157 (N_3157,N_866,N_79);
nor U3158 (N_3158,N_2417,N_2705);
or U3159 (N_3159,N_2839,N_2787);
or U3160 (N_3160,N_146,N_92);
nor U3161 (N_3161,N_1598,N_1016);
xnor U3162 (N_3162,N_2103,N_2764);
and U3163 (N_3163,N_1214,N_465);
nor U3164 (N_3164,N_45,N_1623);
and U3165 (N_3165,N_2426,N_1336);
and U3166 (N_3166,N_1710,N_1854);
and U3167 (N_3167,N_1526,N_2363);
nand U3168 (N_3168,N_2972,N_697);
nand U3169 (N_3169,N_1838,N_2026);
nor U3170 (N_3170,N_748,N_440);
nand U3171 (N_3171,N_1947,N_2899);
xor U3172 (N_3172,N_727,N_1458);
nor U3173 (N_3173,N_1397,N_739);
nor U3174 (N_3174,N_2671,N_2385);
or U3175 (N_3175,N_3089,N_1952);
nor U3176 (N_3176,N_2485,N_423);
xnor U3177 (N_3177,N_750,N_1371);
xnor U3178 (N_3178,N_2725,N_1689);
xor U3179 (N_3179,N_1880,N_531);
nor U3180 (N_3180,N_898,N_1109);
and U3181 (N_3181,N_2840,N_1825);
or U3182 (N_3182,N_2737,N_897);
xnor U3183 (N_3183,N_1309,N_1918);
xnor U3184 (N_3184,N_1324,N_2467);
and U3185 (N_3185,N_2249,N_1255);
nor U3186 (N_3186,N_2983,N_2668);
nand U3187 (N_3187,N_1075,N_3093);
and U3188 (N_3188,N_2789,N_1787);
nand U3189 (N_3189,N_2586,N_1945);
xnor U3190 (N_3190,N_2137,N_1086);
or U3191 (N_3191,N_2939,N_2172);
nand U3192 (N_3192,N_2852,N_2567);
nand U3193 (N_3193,N_1799,N_277);
and U3194 (N_3194,N_7,N_1250);
nand U3195 (N_3195,N_2578,N_563);
xor U3196 (N_3196,N_1957,N_728);
and U3197 (N_3197,N_784,N_2038);
nand U3198 (N_3198,N_2121,N_2978);
xnor U3199 (N_3199,N_3012,N_3091);
xnor U3200 (N_3200,N_461,N_2314);
or U3201 (N_3201,N_2773,N_1404);
xor U3202 (N_3202,N_2376,N_2425);
nor U3203 (N_3203,N_687,N_837);
xor U3204 (N_3204,N_1399,N_1418);
nor U3205 (N_3205,N_3019,N_2591);
and U3206 (N_3206,N_2453,N_2642);
and U3207 (N_3207,N_194,N_2751);
or U3208 (N_3208,N_1089,N_1036);
nand U3209 (N_3209,N_1939,N_1822);
nand U3210 (N_3210,N_1402,N_1911);
xnor U3211 (N_3211,N_1031,N_178);
and U3212 (N_3212,N_1857,N_1979);
nor U3213 (N_3213,N_1684,N_2760);
xor U3214 (N_3214,N_183,N_1746);
xor U3215 (N_3215,N_699,N_1283);
and U3216 (N_3216,N_1410,N_1888);
nand U3217 (N_3217,N_2289,N_1739);
nor U3218 (N_3218,N_413,N_3000);
or U3219 (N_3219,N_2888,N_2890);
nand U3220 (N_3220,N_2298,N_1352);
or U3221 (N_3221,N_2218,N_2023);
nand U3222 (N_3222,N_2373,N_2280);
and U3223 (N_3223,N_224,N_611);
xnor U3224 (N_3224,N_2655,N_592);
nand U3225 (N_3225,N_3057,N_1424);
nor U3226 (N_3226,N_404,N_1836);
nor U3227 (N_3227,N_3095,N_457);
xnor U3228 (N_3228,N_2987,N_294);
xnor U3229 (N_3229,N_2597,N_1847);
xor U3230 (N_3230,N_225,N_2950);
nand U3231 (N_3231,N_1403,N_1515);
and U3232 (N_3232,N_706,N_1319);
or U3233 (N_3233,N_1197,N_3058);
or U3234 (N_3234,N_2680,N_2006);
nor U3235 (N_3235,N_68,N_1563);
and U3236 (N_3236,N_1198,N_2113);
xor U3237 (N_3237,N_334,N_908);
and U3238 (N_3238,N_2362,N_948);
xnor U3239 (N_3239,N_2246,N_2643);
and U3240 (N_3240,N_2964,N_2577);
and U3241 (N_3241,N_54,N_176);
or U3242 (N_3242,N_267,N_1124);
or U3243 (N_3243,N_2822,N_1940);
or U3244 (N_3244,N_107,N_2458);
xor U3245 (N_3245,N_3022,N_1891);
nand U3246 (N_3246,N_2412,N_1706);
nand U3247 (N_3247,N_712,N_1693);
or U3248 (N_3248,N_1375,N_2953);
nor U3249 (N_3249,N_828,N_2776);
nor U3250 (N_3250,N_280,N_1362);
nor U3251 (N_3251,N_1208,N_756);
or U3252 (N_3252,N_1976,N_1987);
and U3253 (N_3253,N_2534,N_2792);
nor U3254 (N_3254,N_1131,N_3001);
xnor U3255 (N_3255,N_676,N_688);
xor U3256 (N_3256,N_2438,N_1020);
xnor U3257 (N_3257,N_84,N_2117);
xnor U3258 (N_3258,N_1005,N_2482);
nor U3259 (N_3259,N_537,N_1567);
or U3260 (N_3260,N_259,N_2866);
or U3261 (N_3261,N_418,N_1367);
xnor U3262 (N_3262,N_600,N_2456);
xnor U3263 (N_3263,N_529,N_2454);
or U3264 (N_3264,N_2302,N_448);
nand U3265 (N_3265,N_268,N_202);
or U3266 (N_3266,N_1586,N_3099);
or U3267 (N_3267,N_2092,N_65);
xor U3268 (N_3268,N_516,N_165);
or U3269 (N_3269,N_2673,N_1938);
or U3270 (N_3270,N_1396,N_2460);
or U3271 (N_3271,N_2605,N_984);
nand U3272 (N_3272,N_2204,N_1926);
nand U3273 (N_3273,N_911,N_2768);
nand U3274 (N_3274,N_1553,N_1033);
or U3275 (N_3275,N_401,N_1675);
or U3276 (N_3276,N_1641,N_2982);
or U3277 (N_3277,N_2261,N_468);
nor U3278 (N_3278,N_2336,N_2728);
xor U3279 (N_3279,N_1747,N_3034);
or U3280 (N_3280,N_2423,N_1099);
or U3281 (N_3281,N_308,N_3031);
and U3282 (N_3282,N_715,N_1039);
xor U3283 (N_3283,N_2594,N_2979);
nor U3284 (N_3284,N_546,N_2918);
or U3285 (N_3285,N_1671,N_1286);
xor U3286 (N_3286,N_2312,N_2075);
and U3287 (N_3287,N_2540,N_2750);
nand U3288 (N_3288,N_222,N_2128);
nor U3289 (N_3289,N_685,N_1719);
nor U3290 (N_3290,N_2942,N_3060);
xor U3291 (N_3291,N_2390,N_463);
xor U3292 (N_3292,N_105,N_320);
nor U3293 (N_3293,N_1308,N_1784);
and U3294 (N_3294,N_232,N_1179);
nor U3295 (N_3295,N_1216,N_223);
xor U3296 (N_3296,N_2645,N_1451);
xor U3297 (N_3297,N_2459,N_1018);
xnor U3298 (N_3298,N_2993,N_2366);
nor U3299 (N_3299,N_1392,N_883);
and U3300 (N_3300,N_2991,N_1999);
nor U3301 (N_3301,N_554,N_339);
nand U3302 (N_3302,N_3106,N_4);
and U3303 (N_3303,N_1146,N_2646);
nor U3304 (N_3304,N_949,N_1380);
xor U3305 (N_3305,N_2757,N_2473);
or U3306 (N_3306,N_1774,N_1660);
nand U3307 (N_3307,N_1186,N_1815);
nor U3308 (N_3308,N_3039,N_2013);
xnor U3309 (N_3309,N_264,N_597);
and U3310 (N_3310,N_125,N_2324);
xnor U3311 (N_3311,N_1287,N_1254);
xnor U3312 (N_3312,N_1870,N_1436);
nor U3313 (N_3313,N_2420,N_735);
and U3314 (N_3314,N_381,N_1264);
and U3315 (N_3315,N_786,N_1485);
or U3316 (N_3316,N_3070,N_2095);
nor U3317 (N_3317,N_241,N_1128);
nand U3318 (N_3318,N_1628,N_1541);
xor U3319 (N_3319,N_3059,N_2464);
or U3320 (N_3320,N_2190,N_1317);
nor U3321 (N_3321,N_919,N_1795);
and U3322 (N_3322,N_2205,N_1730);
or U3323 (N_3323,N_483,N_2549);
nor U3324 (N_3324,N_1607,N_1382);
and U3325 (N_3325,N_2533,N_3086);
nand U3326 (N_3326,N_50,N_1465);
xnor U3327 (N_3327,N_141,N_1653);
nor U3328 (N_3328,N_953,N_1801);
and U3329 (N_3329,N_1225,N_1683);
and U3330 (N_3330,N_2746,N_742);
xor U3331 (N_3331,N_618,N_1236);
and U3332 (N_3332,N_573,N_1142);
nand U3333 (N_3333,N_1085,N_700);
nor U3334 (N_3334,N_1476,N_2271);
or U3335 (N_3335,N_686,N_604);
and U3336 (N_3336,N_2322,N_1276);
or U3337 (N_3337,N_796,N_926);
nand U3338 (N_3338,N_2518,N_104);
nor U3339 (N_3339,N_1949,N_605);
and U3340 (N_3340,N_207,N_918);
nand U3341 (N_3341,N_1323,N_2844);
or U3342 (N_3342,N_1391,N_1440);
nor U3343 (N_3343,N_2435,N_598);
nand U3344 (N_3344,N_255,N_1521);
and U3345 (N_3345,N_3047,N_2869);
and U3346 (N_3346,N_2730,N_2186);
xnor U3347 (N_3347,N_1630,N_1528);
or U3348 (N_3348,N_1723,N_2210);
nand U3349 (N_3349,N_1077,N_2321);
or U3350 (N_3350,N_507,N_374);
xor U3351 (N_3351,N_1067,N_359);
and U3352 (N_3352,N_3042,N_2628);
xnor U3353 (N_3353,N_1055,N_2816);
nand U3354 (N_3354,N_972,N_2735);
and U3355 (N_3355,N_32,N_798);
nor U3356 (N_3356,N_1707,N_2875);
nor U3357 (N_3357,N_3108,N_2073);
and U3358 (N_3358,N_2238,N_342);
xor U3359 (N_3359,N_2841,N_2080);
or U3360 (N_3360,N_1708,N_2359);
and U3361 (N_3361,N_1613,N_3037);
nand U3362 (N_3362,N_2732,N_43);
and U3363 (N_3363,N_624,N_2040);
xor U3364 (N_3364,N_635,N_1224);
and U3365 (N_3365,N_1296,N_2074);
or U3366 (N_3366,N_2820,N_2328);
or U3367 (N_3367,N_1429,N_430);
xnor U3368 (N_3368,N_1183,N_2440);
nor U3369 (N_3369,N_134,N_416);
nor U3370 (N_3370,N_469,N_375);
xnor U3371 (N_3371,N_724,N_1281);
and U3372 (N_3372,N_2585,N_421);
and U3373 (N_3373,N_2995,N_383);
or U3374 (N_3374,N_890,N_188);
or U3375 (N_3375,N_3124,N_1472);
or U3376 (N_3376,N_1412,N_2853);
and U3377 (N_3377,N_2468,N_2546);
nand U3378 (N_3378,N_1602,N_405);
nor U3379 (N_3379,N_2589,N_2743);
or U3380 (N_3380,N_754,N_818);
nor U3381 (N_3381,N_876,N_2339);
xnor U3382 (N_3382,N_2267,N_3103);
or U3383 (N_3383,N_662,N_2353);
nand U3384 (N_3384,N_903,N_3122);
or U3385 (N_3385,N_213,N_1346);
nor U3386 (N_3386,N_626,N_212);
and U3387 (N_3387,N_2529,N_127);
and U3388 (N_3388,N_1265,N_2696);
xor U3389 (N_3389,N_1393,N_1017);
xnor U3390 (N_3390,N_200,N_978);
and U3391 (N_3391,N_1824,N_2164);
or U3392 (N_3392,N_2824,N_1912);
and U3393 (N_3393,N_1975,N_2602);
and U3394 (N_3394,N_298,N_1758);
nor U3395 (N_3395,N_1956,N_517);
and U3396 (N_3396,N_1648,N_807);
or U3397 (N_3397,N_1864,N_1073);
xnor U3398 (N_3398,N_426,N_508);
nor U3399 (N_3399,N_2452,N_1100);
and U3400 (N_3400,N_2631,N_1994);
nor U3401 (N_3401,N_1921,N_2576);
or U3402 (N_3402,N_1027,N_1043);
nor U3403 (N_3403,N_2803,N_2632);
nor U3404 (N_3404,N_2244,N_774);
or U3405 (N_3405,N_2650,N_2392);
and U3406 (N_3406,N_2545,N_1449);
and U3407 (N_3407,N_2356,N_872);
xnor U3408 (N_3408,N_714,N_425);
or U3409 (N_3409,N_2493,N_2588);
and U3410 (N_3410,N_1428,N_2414);
xor U3411 (N_3411,N_377,N_2036);
xor U3412 (N_3412,N_870,N_603);
nand U3413 (N_3413,N_695,N_2063);
nor U3414 (N_3414,N_1,N_1698);
nor U3415 (N_3415,N_1877,N_386);
xnor U3416 (N_3416,N_2834,N_1047);
nor U3417 (N_3417,N_2019,N_1509);
and U3418 (N_3418,N_2887,N_2706);
nand U3419 (N_3419,N_338,N_356);
and U3420 (N_3420,N_454,N_99);
and U3421 (N_3421,N_2835,N_2329);
nand U3422 (N_3422,N_2962,N_3082);
xnor U3423 (N_3423,N_2913,N_3046);
nor U3424 (N_3424,N_2278,N_1669);
xor U3425 (N_3425,N_2144,N_1469);
and U3426 (N_3426,N_2603,N_2695);
xor U3427 (N_3427,N_1110,N_1327);
and U3428 (N_3428,N_2487,N_2946);
and U3429 (N_3429,N_1019,N_2090);
xor U3430 (N_3430,N_1483,N_913);
or U3431 (N_3431,N_2821,N_22);
xnor U3432 (N_3432,N_1614,N_616);
nand U3433 (N_3433,N_1106,N_2192);
nand U3434 (N_3434,N_435,N_378);
xnor U3435 (N_3435,N_594,N_856);
or U3436 (N_3436,N_891,N_1066);
nor U3437 (N_3437,N_1720,N_1721);
xnor U3438 (N_3438,N_2431,N_799);
or U3439 (N_3439,N_2120,N_1965);
nand U3440 (N_3440,N_596,N_229);
or U3441 (N_3441,N_2608,N_253);
nand U3442 (N_3442,N_1692,N_1775);
nand U3443 (N_3443,N_2031,N_2763);
nand U3444 (N_3444,N_1522,N_1411);
and U3445 (N_3445,N_1232,N_874);
or U3446 (N_3446,N_1656,N_2521);
nor U3447 (N_3447,N_1892,N_1427);
nand U3448 (N_3448,N_2729,N_653);
nor U3449 (N_3449,N_836,N_1572);
and U3450 (N_3450,N_2806,N_2927);
nand U3451 (N_3451,N_942,N_1839);
and U3452 (N_3452,N_1491,N_2842);
and U3453 (N_3453,N_1667,N_2227);
or U3454 (N_3454,N_2916,N_1329);
nand U3455 (N_3455,N_1811,N_15);
nand U3456 (N_3456,N_449,N_2288);
nand U3457 (N_3457,N_3007,N_2401);
xor U3458 (N_3458,N_337,N_94);
and U3459 (N_3459,N_1702,N_1445);
and U3460 (N_3460,N_195,N_2086);
xnor U3461 (N_3461,N_484,N_452);
or U3462 (N_3462,N_2669,N_655);
and U3463 (N_3463,N_1941,N_2797);
nor U3464 (N_3464,N_1907,N_2156);
and U3465 (N_3465,N_1853,N_2130);
or U3466 (N_3466,N_2097,N_1727);
or U3467 (N_3467,N_1805,N_2268);
xor U3468 (N_3468,N_2538,N_1158);
and U3469 (N_3469,N_3068,N_1405);
xnor U3470 (N_3470,N_740,N_1148);
and U3471 (N_3471,N_800,N_2727);
nor U3472 (N_3472,N_2644,N_5);
or U3473 (N_3473,N_2457,N_620);
and U3474 (N_3474,N_1307,N_665);
xor U3475 (N_3475,N_1685,N_649);
or U3476 (N_3476,N_1544,N_2739);
and U3477 (N_3477,N_902,N_589);
nor U3478 (N_3478,N_3079,N_539);
and U3479 (N_3479,N_2004,N_820);
nand U3480 (N_3480,N_2397,N_34);
or U3481 (N_3481,N_276,N_2110);
nor U3482 (N_3482,N_1722,N_861);
nor U3483 (N_3483,N_845,N_1591);
nor U3484 (N_3484,N_450,N_2761);
xor U3485 (N_3485,N_1454,N_868);
nor U3486 (N_3486,N_1149,N_887);
nor U3487 (N_3487,N_1792,N_710);
xor U3488 (N_3488,N_2614,N_744);
nand U3489 (N_3489,N_191,N_490);
or U3490 (N_3490,N_2886,N_2948);
or U3491 (N_3491,N_37,N_2997);
nor U3492 (N_3492,N_963,N_2832);
and U3493 (N_3493,N_1873,N_2548);
or U3494 (N_3494,N_1417,N_392);
nor U3495 (N_3495,N_2871,N_1088);
or U3496 (N_3496,N_393,N_2749);
nor U3497 (N_3497,N_844,N_1355);
xor U3498 (N_3498,N_2779,N_2300);
and U3499 (N_3499,N_543,N_1866);
xor U3500 (N_3500,N_506,N_236);
nor U3501 (N_3501,N_1426,N_265);
nand U3502 (N_3502,N_1026,N_2836);
or U3503 (N_3503,N_2230,N_1756);
nor U3504 (N_3504,N_2936,N_2909);
and U3505 (N_3505,N_228,N_2035);
and U3506 (N_3506,N_2348,N_346);
and U3507 (N_3507,N_2703,N_2216);
or U3508 (N_3508,N_3113,N_2648);
and U3509 (N_3509,N_2952,N_451);
or U3510 (N_3510,N_3078,N_2537);
and U3511 (N_3511,N_2947,N_2303);
nand U3512 (N_3512,N_1884,N_436);
xnor U3513 (N_3513,N_2301,N_2162);
xnor U3514 (N_3514,N_522,N_2045);
or U3515 (N_3515,N_525,N_210);
and U3516 (N_3516,N_2744,N_345);
and U3517 (N_3517,N_2506,N_167);
and U3518 (N_3518,N_1090,N_1447);
nor U3519 (N_3519,N_58,N_208);
or U3520 (N_3520,N_924,N_1215);
nor U3521 (N_3521,N_2174,N_2880);
nor U3522 (N_3522,N_2653,N_2220);
or U3523 (N_3523,N_3123,N_1434);
or U3524 (N_3524,N_2494,N_1676);
and U3525 (N_3525,N_2513,N_62);
nand U3526 (N_3526,N_788,N_2782);
xnor U3527 (N_3527,N_643,N_1933);
nand U3528 (N_3528,N_896,N_2897);
or U3529 (N_3529,N_1072,N_149);
nor U3530 (N_3530,N_1903,N_1978);
xor U3531 (N_3531,N_2147,N_3044);
and U3532 (N_3532,N_2652,N_36);
xor U3533 (N_3533,N_2829,N_2185);
or U3534 (N_3534,N_2087,N_1495);
xnor U3535 (N_3535,N_1849,N_3120);
xor U3536 (N_3536,N_2396,N_1369);
nand U3537 (N_3537,N_2505,N_1477);
or U3538 (N_3538,N_502,N_3014);
and U3539 (N_3539,N_2181,N_809);
nand U3540 (N_3540,N_2477,N_1637);
nor U3541 (N_3541,N_1136,N_2251);
or U3542 (N_3542,N_3041,N_2106);
and U3543 (N_3543,N_1237,N_1318);
nand U3544 (N_3544,N_561,N_2149);
and U3545 (N_3545,N_1876,N_91);
or U3546 (N_3546,N_2837,N_711);
nor U3547 (N_3547,N_2944,N_419);
nor U3548 (N_3548,N_279,N_1137);
xnor U3549 (N_3549,N_1456,N_2781);
nor U3550 (N_3550,N_869,N_2222);
nor U3551 (N_3551,N_503,N_467);
nand U3552 (N_3552,N_1627,N_936);
xnor U3553 (N_3553,N_1230,N_126);
xnor U3554 (N_3554,N_1504,N_933);
or U3555 (N_3555,N_1222,N_785);
or U3556 (N_3556,N_2299,N_990);
xnor U3557 (N_3557,N_329,N_1359);
nand U3558 (N_3558,N_646,N_460);
nand U3559 (N_3559,N_1852,N_238);
or U3560 (N_3560,N_437,N_2057);
or U3561 (N_3561,N_2072,N_2187);
or U3562 (N_3562,N_397,N_2058);
and U3563 (N_3563,N_1626,N_1642);
nor U3564 (N_3564,N_1790,N_1345);
nand U3565 (N_3565,N_3081,N_833);
xor U3566 (N_3566,N_233,N_67);
nor U3567 (N_3567,N_3008,N_1924);
and U3568 (N_3568,N_1791,N_1647);
or U3569 (N_3569,N_1244,N_1299);
and U3570 (N_3570,N_2524,N_90);
nor U3571 (N_3571,N_474,N_341);
nand U3572 (N_3572,N_1499,N_1135);
and U3573 (N_3573,N_2209,N_1753);
xor U3574 (N_3574,N_1761,N_633);
xor U3575 (N_3575,N_1322,N_3032);
or U3576 (N_3576,N_350,N_197);
xnor U3577 (N_3577,N_639,N_1154);
or U3578 (N_3578,N_2260,N_1837);
or U3579 (N_3579,N_3100,N_2122);
or U3580 (N_3580,N_825,N_1430);
and U3581 (N_3581,N_854,N_2433);
nor U3582 (N_3582,N_2818,N_1431);
or U3583 (N_3583,N_400,N_1512);
or U3584 (N_3584,N_2912,N_2255);
nand U3585 (N_3585,N_145,N_941);
nand U3586 (N_3586,N_583,N_1780);
nand U3587 (N_3587,N_551,N_2126);
or U3588 (N_3588,N_2527,N_231);
xnor U3589 (N_3589,N_2201,N_1718);
and U3590 (N_3590,N_1769,N_2002);
nor U3591 (N_3591,N_945,N_975);
nor U3592 (N_3592,N_3105,N_619);
nor U3593 (N_3593,N_2618,N_863);
and U3594 (N_3594,N_691,N_1115);
and U3595 (N_3595,N_888,N_2692);
nand U3596 (N_3596,N_2168,N_2253);
nand U3597 (N_3597,N_808,N_925);
xor U3598 (N_3598,N_3110,N_441);
nand U3599 (N_3599,N_2461,N_2713);
and U3600 (N_3600,N_301,N_2902);
nand U3601 (N_3601,N_3006,N_1717);
nor U3602 (N_3602,N_1724,N_1481);
nand U3603 (N_3603,N_480,N_545);
xnor U3604 (N_3604,N_2091,N_1119);
or U3605 (N_3605,N_970,N_2340);
nand U3606 (N_3606,N_2639,N_2647);
xnor U3607 (N_3607,N_76,N_1079);
nand U3608 (N_3608,N_2306,N_2171);
or U3609 (N_3609,N_1246,N_1779);
nand U3610 (N_3610,N_2582,N_139);
nand U3611 (N_3611,N_599,N_1661);
and U3612 (N_3612,N_932,N_1599);
xor U3613 (N_3613,N_775,N_1139);
nand U3614 (N_3614,N_2796,N_1919);
nand U3615 (N_3615,N_458,N_2963);
and U3616 (N_3616,N_160,N_2051);
xnor U3617 (N_3617,N_1640,N_1991);
nand U3618 (N_3618,N_1455,N_1557);
nor U3619 (N_3619,N_680,N_3117);
or U3620 (N_3620,N_2687,N_623);
and U3621 (N_3621,N_243,N_3112);
or U3622 (N_3622,N_2612,N_82);
nor U3623 (N_3623,N_795,N_2969);
xnor U3624 (N_3624,N_77,N_317);
nor U3625 (N_3625,N_2357,N_1168);
and U3626 (N_3626,N_2557,N_155);
nor U3627 (N_3627,N_1262,N_498);
xor U3628 (N_3628,N_2173,N_817);
xor U3629 (N_3629,N_2099,N_283);
or U3630 (N_3630,N_1261,N_2350);
or U3631 (N_3631,N_2966,N_1794);
nand U3632 (N_3632,N_556,N_1898);
nor U3633 (N_3633,N_2085,N_1520);
xor U3634 (N_3634,N_2667,N_1360);
or U3635 (N_3635,N_315,N_1517);
nor U3636 (N_3636,N_2870,N_380);
and U3637 (N_3637,N_1634,N_2892);
and U3638 (N_3638,N_2813,N_2474);
or U3639 (N_3639,N_2954,N_1196);
nor U3640 (N_3640,N_410,N_549);
or U3641 (N_3641,N_1452,N_2654);
xnor U3642 (N_3642,N_237,N_2365);
and U3643 (N_3643,N_442,N_2067);
nor U3644 (N_3644,N_1312,N_2999);
nand U3645 (N_3645,N_3009,N_2100);
nand U3646 (N_3646,N_2862,N_2240);
nor U3647 (N_3647,N_2490,N_1291);
nor U3648 (N_3648,N_1151,N_1270);
or U3649 (N_3649,N_585,N_1132);
and U3650 (N_3650,N_180,N_906);
and U3651 (N_3651,N_2901,N_1651);
and U3652 (N_3652,N_766,N_1985);
nor U3653 (N_3653,N_1609,N_1171);
xor U3654 (N_3654,N_2105,N_19);
xnor U3655 (N_3655,N_24,N_2851);
nand U3656 (N_3656,N_950,N_396);
or U3657 (N_3657,N_2021,N_2634);
xor U3658 (N_3658,N_2664,N_753);
or U3659 (N_3659,N_1915,N_2124);
or U3660 (N_3660,N_1038,N_1534);
nor U3661 (N_3661,N_787,N_1321);
or U3662 (N_3662,N_1983,N_1749);
nand U3663 (N_3663,N_2802,N_60);
nand U3664 (N_3664,N_479,N_1754);
xnor U3665 (N_3665,N_412,N_1121);
nand U3666 (N_3666,N_1989,N_2402);
and U3667 (N_3667,N_367,N_1986);
nand U3668 (N_3668,N_1461,N_2028);
nor U3669 (N_3669,N_1443,N_1441);
or U3670 (N_3670,N_2308,N_1141);
nand U3671 (N_3671,N_2009,N_1160);
nand U3672 (N_3672,N_1191,N_3020);
or U3673 (N_3673,N_2701,N_2503);
nor U3674 (N_3674,N_2265,N_389);
and U3675 (N_3675,N_2352,N_1111);
xnor U3676 (N_3676,N_907,N_1507);
nor U3677 (N_3677,N_69,N_1848);
or U3678 (N_3678,N_120,N_2544);
xnor U3679 (N_3679,N_2243,N_2304);
nor U3680 (N_3680,N_674,N_1511);
xor U3681 (N_3681,N_1095,N_1832);
nor U3682 (N_3682,N_2476,N_173);
xor U3683 (N_3683,N_692,N_608);
and U3684 (N_3684,N_1646,N_133);
xnor U3685 (N_3685,N_428,N_1223);
and U3686 (N_3686,N_1679,N_2434);
nor U3687 (N_3687,N_851,N_1040);
nor U3688 (N_3688,N_1819,N_1251);
and U3689 (N_3689,N_2920,N_2604);
or U3690 (N_3690,N_2015,N_1830);
nand U3691 (N_3691,N_885,N_2256);
and U3692 (N_3692,N_2050,N_2536);
nor U3693 (N_3693,N_1492,N_2012);
and U3694 (N_3694,N_488,N_806);
or U3695 (N_3695,N_2855,N_2677);
or U3696 (N_3696,N_1347,N_1565);
nor U3697 (N_3697,N_2049,N_1398);
xnor U3698 (N_3698,N_1988,N_1374);
or U3699 (N_3699,N_1478,N_1395);
nand U3700 (N_3700,N_1351,N_227);
or U3701 (N_3701,N_2293,N_1210);
or U3702 (N_3702,N_2930,N_1256);
or U3703 (N_3703,N_614,N_343);
nor U3704 (N_3704,N_1234,N_2889);
nand U3705 (N_3705,N_2717,N_1757);
nand U3706 (N_3706,N_2404,N_2202);
nand U3707 (N_3707,N_1778,N_384);
nand U3708 (N_3708,N_2961,N_340);
xnor U3709 (N_3709,N_1101,N_296);
nand U3710 (N_3710,N_302,N_2951);
and U3711 (N_3711,N_865,N_991);
xor U3712 (N_3712,N_1704,N_1536);
nor U3713 (N_3713,N_1594,N_1618);
and U3714 (N_3714,N_2158,N_1973);
nand U3715 (N_3715,N_2129,N_1524);
and U3716 (N_3716,N_1611,N_1570);
or U3717 (N_3717,N_2042,N_1338);
and U3718 (N_3718,N_1498,N_2583);
nor U3719 (N_3719,N_1354,N_1798);
nor U3720 (N_3720,N_2592,N_694);
or U3721 (N_3721,N_2520,N_1968);
nor U3722 (N_3722,N_2665,N_2884);
and U3723 (N_3723,N_455,N_1143);
nor U3724 (N_3724,N_2469,N_1893);
xor U3725 (N_3725,N_513,N_2326);
nor U3726 (N_3726,N_741,N_773);
xnor U3727 (N_3727,N_985,N_2989);
xor U3728 (N_3728,N_1479,N_955);
and U3729 (N_3729,N_473,N_540);
nor U3730 (N_3730,N_1339,N_999);
and U3731 (N_3731,N_824,N_244);
or U3732 (N_3732,N_2738,N_968);
nor U3733 (N_3733,N_2323,N_269);
nor U3734 (N_3734,N_116,N_2974);
or U3735 (N_3735,N_2367,N_586);
or U3736 (N_3736,N_530,N_2131);
xor U3737 (N_3737,N_2427,N_1057);
nor U3738 (N_3738,N_2360,N_864);
nand U3739 (N_3739,N_1964,N_1664);
or U3740 (N_3740,N_100,N_736);
nor U3741 (N_3741,N_2814,N_613);
nand U3742 (N_3742,N_552,N_667);
nand U3743 (N_3743,N_2465,N_1566);
nor U3744 (N_3744,N_2398,N_2082);
nand U3745 (N_3745,N_781,N_2056);
and U3746 (N_3746,N_3092,N_927);
and U3747 (N_3747,N_1796,N_3002);
nor U3748 (N_3748,N_1818,N_406);
and U3749 (N_3749,N_770,N_2335);
xor U3750 (N_3750,N_768,N_568);
xor U3751 (N_3751,N_1233,N_1916);
and U3752 (N_3752,N_2651,N_1269);
or U3753 (N_3753,N_2807,N_763);
nor U3754 (N_3754,N_2368,N_1777);
nor U3755 (N_3755,N_13,N_2488);
nand U3756 (N_3756,N_3015,N_2700);
nand U3757 (N_3757,N_1501,N_733);
xor U3758 (N_3758,N_453,N_1842);
nor U3759 (N_3759,N_647,N_905);
nor U3760 (N_3760,N_2471,N_1044);
and U3761 (N_3761,N_1280,N_2407);
nor U3762 (N_3762,N_2758,N_1004);
nand U3763 (N_3763,N_2895,N_3119);
nand U3764 (N_3764,N_889,N_1226);
or U3765 (N_3765,N_997,N_1841);
or U3766 (N_3766,N_1663,N_1772);
nand U3767 (N_3767,N_3035,N_1592);
or U3768 (N_3768,N_349,N_922);
or U3769 (N_3769,N_108,N_723);
and U3770 (N_3770,N_1034,N_843);
nor U3771 (N_3771,N_1042,N_810);
or U3772 (N_3772,N_1688,N_2587);
xor U3773 (N_3773,N_2157,N_1419);
or U3774 (N_3774,N_168,N_2198);
nor U3775 (N_3775,N_2689,N_179);
xnor U3776 (N_3776,N_1662,N_2683);
xor U3777 (N_3777,N_2955,N_1804);
nand U3778 (N_3778,N_422,N_414);
nand U3779 (N_3779,N_848,N_1091);
nand U3780 (N_3780,N_1789,N_3052);
xnor U3781 (N_3781,N_1204,N_704);
or U3782 (N_3782,N_1908,N_2885);
or U3783 (N_3783,N_1732,N_73);
nor U3784 (N_3784,N_445,N_31);
and U3785 (N_3785,N_1333,N_364);
or U3786 (N_3786,N_2176,N_2127);
nand U3787 (N_3787,N_532,N_3096);
nor U3788 (N_3788,N_2636,N_1363);
nor U3789 (N_3789,N_915,N_1349);
and U3790 (N_3790,N_2347,N_142);
nand U3791 (N_3791,N_2032,N_1341);
xnor U3792 (N_3792,N_187,N_1117);
nand U3793 (N_3793,N_631,N_385);
nor U3794 (N_3794,N_964,N_172);
or U3795 (N_3795,N_2315,N_2071);
or U3796 (N_3796,N_1922,N_2956);
nor U3797 (N_3797,N_3040,N_300);
xor U3798 (N_3798,N_1942,N_989);
or U3799 (N_3799,N_1182,N_3107);
nand U3800 (N_3800,N_1205,N_1058);
or U3801 (N_3801,N_1439,N_928);
or U3802 (N_3802,N_2370,N_2078);
or U3803 (N_3803,N_1153,N_152);
xnor U3804 (N_3804,N_1379,N_499);
or U3805 (N_3805,N_1462,N_725);
xnor U3806 (N_3806,N_415,N_1335);
nand U3807 (N_3807,N_3010,N_369);
or U3808 (N_3808,N_2123,N_2720);
xnor U3809 (N_3809,N_2593,N_3074);
or U3810 (N_3810,N_515,N_3097);
and U3811 (N_3811,N_690,N_1278);
xnor U3812 (N_3812,N_1537,N_373);
xor U3813 (N_3813,N_959,N_581);
nor U3814 (N_3814,N_2731,N_1304);
nand U3815 (N_3815,N_372,N_880);
xnor U3816 (N_3816,N_1800,N_209);
or U3817 (N_3817,N_275,N_696);
or U3818 (N_3818,N_1446,N_2175);
nor U3819 (N_3819,N_2497,N_682);
nand U3820 (N_3820,N_2562,N_2132);
xor U3821 (N_3821,N_2226,N_2020);
nor U3822 (N_3822,N_2199,N_1944);
nand U3823 (N_3823,N_1887,N_93);
or U3824 (N_3824,N_904,N_1860);
nor U3825 (N_3825,N_743,N_2502);
nor U3826 (N_3826,N_1561,N_2932);
nand U3827 (N_3827,N_1670,N_2838);
nand U3828 (N_3828,N_2399,N_2285);
xor U3829 (N_3829,N_2275,N_2169);
and U3830 (N_3830,N_2343,N_1905);
or U3831 (N_3831,N_162,N_1951);
or U3832 (N_3832,N_1539,N_1068);
and U3833 (N_3833,N_862,N_1816);
xor U3834 (N_3834,N_2046,N_1767);
and U3835 (N_3835,N_675,N_1906);
nand U3836 (N_3836,N_2600,N_2194);
nor U3837 (N_3837,N_1259,N_174);
or U3838 (N_3838,N_2101,N_2221);
or U3839 (N_3839,N_57,N_20);
and U3840 (N_3840,N_2447,N_995);
or U3841 (N_3841,N_1743,N_2528);
nor U3842 (N_3842,N_2400,N_1899);
and U3843 (N_3843,N_628,N_1923);
xor U3844 (N_3844,N_1931,N_2908);
xor U3845 (N_3845,N_2804,N_1383);
nand U3846 (N_3846,N_2207,N_2517);
and U3847 (N_3847,N_398,N_2096);
nand U3848 (N_3848,N_1009,N_1271);
or U3849 (N_3849,N_1845,N_681);
or U3850 (N_3850,N_1211,N_678);
and U3851 (N_3851,N_1856,N_3080);
and U3852 (N_3852,N_1579,N_2808);
and U3853 (N_3853,N_46,N_761);
nor U3854 (N_3854,N_1883,N_2584);
nand U3855 (N_3855,N_330,N_2541);
or U3856 (N_3856,N_2709,N_578);
xor U3857 (N_3857,N_2052,N_2369);
xnor U3858 (N_3858,N_1835,N_2510);
and U3859 (N_3859,N_1260,N_2388);
nand U3860 (N_3860,N_2183,N_1484);
nor U3861 (N_3861,N_2001,N_1150);
xor U3862 (N_3862,N_2481,N_1064);
and U3863 (N_3863,N_2877,N_559);
nor U3864 (N_3864,N_1502,N_1343);
and U3865 (N_3865,N_1821,N_1227);
xnor U3866 (N_3866,N_969,N_1970);
xor U3867 (N_3867,N_464,N_409);
and U3868 (N_3868,N_2495,N_566);
xor U3869 (N_3869,N_1834,N_651);
xnor U3870 (N_3870,N_752,N_2016);
xnor U3871 (N_3871,N_572,N_562);
xor U3872 (N_3872,N_161,N_310);
xnor U3873 (N_3873,N_510,N_2960);
or U3874 (N_3874,N_1564,N_2247);
nand U3875 (N_3875,N_1493,N_1011);
and U3876 (N_3876,N_1176,N_131);
or U3877 (N_3877,N_957,N_1766);
or U3878 (N_3878,N_247,N_2409);
or U3879 (N_3879,N_2330,N_2778);
xor U3880 (N_3880,N_9,N_360);
nor U3881 (N_3881,N_284,N_2245);
nor U3882 (N_3882,N_2756,N_328);
nand U3883 (N_3883,N_2292,N_2077);
nand U3884 (N_3884,N_1937,N_542);
or U3885 (N_3885,N_1629,N_977);
xor U3886 (N_3886,N_2212,N_1163);
xor U3887 (N_3887,N_3033,N_306);
xnor U3888 (N_3888,N_1061,N_2580);
or U3889 (N_3889,N_717,N_2290);
or U3890 (N_3890,N_1577,N_2609);
and U3891 (N_3891,N_1863,N_1666);
nor U3892 (N_3892,N_2,N_1473);
xor U3893 (N_3893,N_943,N_3065);
xnor U3894 (N_3894,N_1657,N_1963);
nand U3895 (N_3895,N_2715,N_1093);
nand U3896 (N_3896,N_2772,N_2331);
or U3897 (N_3897,N_1144,N_3028);
nand U3898 (N_3898,N_96,N_266);
nor U3899 (N_3899,N_2235,N_2287);
nor U3900 (N_3900,N_1807,N_882);
or U3901 (N_3901,N_2419,N_219);
nor U3902 (N_3902,N_2010,N_494);
or U3903 (N_3903,N_1913,N_1263);
and U3904 (N_3904,N_1569,N_151);
xor U3905 (N_3905,N_1910,N_553);
nor U3906 (N_3906,N_2215,N_1486);
nand U3907 (N_3907,N_85,N_1114);
nand U3908 (N_3908,N_1900,N_2926);
nand U3909 (N_3909,N_1126,N_2325);
or U3910 (N_3910,N_1806,N_2799);
nor U3911 (N_3911,N_261,N_2767);
or U3912 (N_3912,N_2234,N_2133);
or U3913 (N_3913,N_1340,N_2552);
nand U3914 (N_3914,N_278,N_21);
nor U3915 (N_3915,N_1680,N_2748);
xor U3916 (N_3916,N_2754,N_2155);
and U3917 (N_3917,N_641,N_1875);
nor U3918 (N_3918,N_1540,N_1958);
nand U3919 (N_3919,N_472,N_1356);
xnor U3920 (N_3920,N_492,N_2483);
or U3921 (N_3921,N_1023,N_1177);
or U3922 (N_3922,N_198,N_2937);
or U3923 (N_3923,N_2462,N_1828);
or U3924 (N_3924,N_2043,N_767);
and U3925 (N_3925,N_1311,N_80);
nor U3926 (N_3926,N_2378,N_260);
nand U3927 (N_3927,N_745,N_2405);
and U3928 (N_3928,N_2522,N_801);
and U3929 (N_3929,N_1902,N_993);
xnor U3930 (N_3930,N_973,N_95);
or U3931 (N_3931,N_1174,N_521);
or U3932 (N_3932,N_3023,N_2910);
nor U3933 (N_3933,N_1376,N_966);
or U3934 (N_3934,N_996,N_2523);
nor U3935 (N_3935,N_2678,N_2710);
nand U3936 (N_3936,N_1448,N_2422);
nor U3937 (N_3937,N_481,N_1820);
nand U3938 (N_3938,N_2039,N_1187);
nand U3939 (N_3939,N_1881,N_1288);
or U3940 (N_3940,N_1862,N_1616);
nor U3941 (N_3941,N_150,N_129);
nor U3942 (N_3942,N_1435,N_3064);
xor U3943 (N_3943,N_2064,N_2740);
or U3944 (N_3944,N_1596,N_1213);
or U3945 (N_3945,N_0,N_361);
nand U3946 (N_3946,N_2263,N_2011);
or U3947 (N_3947,N_979,N_2387);
nand U3948 (N_3948,N_1030,N_1731);
and U3949 (N_3949,N_124,N_1394);
xnor U3950 (N_3950,N_2670,N_2660);
xor U3951 (N_3951,N_1221,N_1192);
and U3952 (N_3952,N_2766,N_1081);
and U3953 (N_3953,N_2511,N_427);
xnor U3954 (N_3954,N_764,N_486);
nor U3955 (N_3955,N_2379,N_403);
or U3956 (N_3956,N_2055,N_1955);
xor U3957 (N_3957,N_1600,N_2831);
xor U3958 (N_3958,N_2770,N_789);
xor U3959 (N_3959,N_2965,N_1782);
or U3960 (N_3960,N_1274,N_1530);
nor U3961 (N_3961,N_2027,N_2817);
nand U3962 (N_3962,N_1890,N_35);
or U3963 (N_3963,N_976,N_1700);
nor U3964 (N_3964,N_1886,N_1045);
xnor U3965 (N_3965,N_702,N_1759);
or U3966 (N_3966,N_501,N_199);
nor U3967 (N_3967,N_716,N_1635);
and U3968 (N_3968,N_987,N_938);
and U3969 (N_3969,N_1748,N_2316);
nand U3970 (N_3970,N_2941,N_2206);
xor U3971 (N_3971,N_2140,N_2992);
nand U3972 (N_3972,N_2865,N_2159);
xor U3973 (N_3973,N_1122,N_1080);
or U3974 (N_3974,N_1070,N_2138);
or U3975 (N_3975,N_1946,N_2066);
or U3976 (N_3976,N_216,N_569);
nor U3977 (N_3977,N_2508,N_2575);
and U3978 (N_3978,N_693,N_1496);
nand U3979 (N_3979,N_2170,N_1310);
nand U3980 (N_3980,N_211,N_287);
nand U3981 (N_3981,N_1590,N_3027);
nor U3982 (N_3982,N_344,N_3075);
nor U3983 (N_3983,N_755,N_2923);
nand U3984 (N_3984,N_1175,N_3076);
nand U3985 (N_3985,N_1241,N_1325);
or U3986 (N_3986,N_2719,N_1699);
nor U3987 (N_3987,N_1202,N_582);
and U3988 (N_3988,N_1203,N_2161);
or U3989 (N_3989,N_2499,N_1185);
and U3990 (N_3990,N_2416,N_1673);
and U3991 (N_3991,N_1437,N_2338);
nand U3992 (N_3992,N_2436,N_1840);
xor U3993 (N_3993,N_1697,N_909);
and U3994 (N_3994,N_1444,N_2610);
xnor U3995 (N_3995,N_3016,N_1650);
xnor U3996 (N_3996,N_204,N_2733);
or U3997 (N_3997,N_1726,N_2008);
and U3998 (N_3998,N_52,N_470);
or U3999 (N_3999,N_650,N_2613);
xor U4000 (N_4000,N_547,N_571);
xnor U4001 (N_4001,N_1243,N_106);
xor U4002 (N_4002,N_1408,N_640);
xor U4003 (N_4003,N_331,N_661);
nand U4004 (N_4004,N_698,N_2504);
xnor U4005 (N_4005,N_811,N_203);
and U4006 (N_4006,N_371,N_2681);
xor U4007 (N_4007,N_2935,N_2938);
or U4008 (N_4008,N_2098,N_1328);
nand U4009 (N_4009,N_2532,N_495);
nor U4010 (N_4010,N_1971,N_982);
and U4011 (N_4011,N_505,N_250);
nor U4012 (N_4012,N_2125,N_550);
nand U4013 (N_4013,N_2022,N_2550);
nor U4014 (N_4014,N_2984,N_2907);
and U4015 (N_4015,N_934,N_3005);
nand U4016 (N_4016,N_25,N_584);
nor U4017 (N_4017,N_2833,N_929);
xor U4018 (N_4018,N_842,N_336);
or U4019 (N_4019,N_3116,N_2786);
or U4020 (N_4020,N_1432,N_185);
nand U4021 (N_4021,N_705,N_23);
and U4022 (N_4022,N_130,N_291);
xnor U4023 (N_4023,N_182,N_2752);
and U4024 (N_4024,N_2641,N_1581);
or U4025 (N_4025,N_1715,N_778);
xor U4026 (N_4026,N_56,N_323);
nor U4027 (N_4027,N_901,N_2200);
nor U4028 (N_4028,N_1786,N_493);
or U4029 (N_4029,N_892,N_2135);
xor U4030 (N_4030,N_64,N_952);
xor U4031 (N_4031,N_2911,N_1316);
and U4032 (N_4032,N_1686,N_567);
and U4033 (N_4033,N_111,N_2472);
xor U4034 (N_4034,N_2514,N_2535);
nor U4035 (N_4035,N_1781,N_1808);
and U4036 (N_4036,N_689,N_293);
or U4037 (N_4037,N_3066,N_670);
or U4038 (N_4038,N_1006,N_332);
and U4039 (N_4039,N_262,N_644);
xnor U4040 (N_4040,N_1133,N_713);
nor U4041 (N_4041,N_1740,N_1219);
nand U4042 (N_4042,N_2437,N_962);
xor U4043 (N_4043,N_536,N_2850);
or U4044 (N_4044,N_2224,N_3118);
and U4045 (N_4045,N_1885,N_1247);
nand U4046 (N_4046,N_846,N_1936);
and U4047 (N_4047,N_2894,N_2178);
nand U4048 (N_4048,N_1293,N_2904);
xor U4049 (N_4049,N_1652,N_193);
xnor U4050 (N_4050,N_762,N_3084);
xnor U4051 (N_4051,N_1621,N_1826);
xnor U4052 (N_4052,N_1532,N_1273);
xor U4053 (N_4053,N_491,N_2699);
nand U4054 (N_4054,N_2371,N_2424);
xnor U4055 (N_4055,N_738,N_899);
nor U4056 (N_4056,N_1140,N_780);
and U4057 (N_4057,N_2395,N_1268);
xnor U4058 (N_4058,N_2076,N_1457);
or U4059 (N_4059,N_954,N_2153);
xor U4060 (N_4060,N_26,N_2794);
xor U4061 (N_4061,N_829,N_2295);
xor U4062 (N_4062,N_1878,N_1161);
and U4063 (N_4063,N_2239,N_1813);
xnor U4064 (N_4064,N_245,N_2690);
nor U4065 (N_4065,N_1002,N_263);
nand U4066 (N_4066,N_2486,N_309);
or U4067 (N_4067,N_971,N_2924);
nor U4068 (N_4068,N_2615,N_28);
xnor U4069 (N_4069,N_2906,N_119);
or U4070 (N_4070,N_2211,N_33);
or U4071 (N_4071,N_1013,N_1966);
and U4072 (N_4072,N_1051,N_1188);
nor U4073 (N_4073,N_2917,N_2531);
nand U4074 (N_4074,N_637,N_1228);
xnor U4075 (N_4075,N_2684,N_722);
and U4076 (N_4076,N_657,N_2509);
xor U4077 (N_4077,N_875,N_2266);
nor U4078 (N_4078,N_2160,N_2915);
nor U4079 (N_4079,N_1967,N_1123);
or U4080 (N_4080,N_1505,N_1658);
xnor U4081 (N_4081,N_2812,N_895);
or U4082 (N_4082,N_2319,N_2017);
and U4083 (N_4083,N_2685,N_606);
or U4084 (N_4084,N_886,N_2418);
nand U4085 (N_4085,N_477,N_1982);
nor U4086 (N_4086,N_2674,N_1859);
xnor U4087 (N_4087,N_299,N_271);
xnor U4088 (N_4088,N_1981,N_1582);
nand U4089 (N_4089,N_1977,N_1568);
nor U4090 (N_4090,N_1714,N_1054);
nand U4091 (N_4091,N_305,N_1555);
xor U4092 (N_4092,N_2967,N_2697);
nor U4093 (N_4093,N_2236,N_2878);
nand U4094 (N_4094,N_1874,N_1012);
nor U4095 (N_4095,N_1385,N_1851);
xnor U4096 (N_4096,N_2463,N_1542);
nand U4097 (N_4097,N_89,N_230);
and U4098 (N_4098,N_2542,N_2327);
nor U4099 (N_4099,N_2364,N_2547);
nand U4100 (N_4100,N_2047,N_1506);
xor U4101 (N_4101,N_3045,N_1531);
nand U4102 (N_4102,N_1167,N_520);
or U4103 (N_4103,N_1113,N_1632);
or U4104 (N_4104,N_2771,N_254);
nor U4105 (N_4105,N_1802,N_117);
nor U4106 (N_4106,N_1738,N_1909);
and U4107 (N_4107,N_411,N_873);
and U4108 (N_4108,N_1125,N_2429);
nand U4109 (N_4109,N_2383,N_1157);
nor U4110 (N_4110,N_1366,N_2556);
nor U4111 (N_4111,N_1644,N_1768);
nor U4112 (N_4112,N_1578,N_2649);
nor U4113 (N_4113,N_1810,N_1021);
or U4114 (N_4114,N_2559,N_420);
nand U4115 (N_4115,N_1829,N_2512);
or U4116 (N_4116,N_1041,N_318);
nand U4117 (N_4117,N_2048,N_791);
or U4118 (N_4118,N_1846,N_1464);
xnor U4119 (N_4119,N_476,N_2166);
and U4120 (N_4120,N_39,N_2358);
nor U4121 (N_4121,N_2726,N_1674);
nand U4122 (N_4122,N_792,N_2184);
nor U4123 (N_4123,N_533,N_612);
nor U4124 (N_4124,N_2718,N_1159);
xnor U4125 (N_4125,N_2724,N_2203);
or U4126 (N_4126,N_2753,N_2059);
nand U4127 (N_4127,N_2986,N_2599);
or U4128 (N_4128,N_1378,N_1025);
xor U4129 (N_4129,N_1959,N_2276);
and U4130 (N_4130,N_632,N_1295);
and U4131 (N_4131,N_609,N_2361);
and U4132 (N_4132,N_1503,N_2784);
nor U4133 (N_4133,N_1162,N_1773);
or U4134 (N_4134,N_1292,N_164);
nand U4135 (N_4135,N_27,N_841);
nand U4136 (N_4136,N_1682,N_2083);
and U4137 (N_4137,N_816,N_2863);
nor U4138 (N_4138,N_132,N_1201);
nand U4139 (N_4139,N_684,N_2033);
xnor U4140 (N_4140,N_528,N_1342);
nor U4141 (N_4141,N_2672,N_2598);
and U4142 (N_4142,N_1668,N_2208);
nor U4143 (N_4143,N_1950,N_316);
nand U4144 (N_4144,N_718,N_621);
or U4145 (N_4145,N_1320,N_70);
or U4146 (N_4146,N_601,N_2790);
nor U4147 (N_4147,N_1266,N_504);
or U4148 (N_4148,N_1831,N_638);
nand U4149 (N_4149,N_1272,N_42);
xnor U4150 (N_4150,N_2007,N_804);
and U4151 (N_4151,N_1334,N_1711);
nor U4152 (N_4152,N_2351,N_2553);
nand U4153 (N_4153,N_273,N_3053);
or U4154 (N_4154,N_1580,N_776);
and U4155 (N_4155,N_102,N_1453);
nor U4156 (N_4156,N_2988,N_668);
xnor U4157 (N_4157,N_910,N_1350);
and U4158 (N_4158,N_355,N_471);
and U4159 (N_4159,N_3049,N_802);
or U4160 (N_4160,N_1056,N_2940);
or U4161 (N_4161,N_2971,N_1709);
xnor U4162 (N_4162,N_2570,N_1384);
and U4163 (N_4163,N_1997,N_790);
nand U4164 (N_4164,N_974,N_1858);
xnor U4165 (N_4165,N_235,N_2345);
nor U4166 (N_4166,N_1696,N_354);
and U4167 (N_4167,N_1643,N_2860);
and U4168 (N_4168,N_74,N_1267);
nand U4169 (N_4169,N_2445,N_2225);
nor U4170 (N_4170,N_2070,N_721);
or U4171 (N_4171,N_1765,N_588);
or U4172 (N_4172,N_311,N_893);
or U4173 (N_4173,N_2470,N_666);
nor U4174 (N_4174,N_1527,N_703);
nand U4175 (N_4175,N_2931,N_1145);
or U4176 (N_4176,N_1934,N_2180);
and U4177 (N_4177,N_1466,N_297);
or U4178 (N_4178,N_1294,N_672);
xor U4179 (N_4179,N_2561,N_564);
nor U4180 (N_4180,N_2949,N_2489);
nor U4181 (N_4181,N_1574,N_109);
nand U4182 (N_4182,N_857,N_730);
xnor U4183 (N_4183,N_2847,N_830);
or U4184 (N_4184,N_3018,N_362);
nand U4185 (N_4185,N_1037,N_2516);
and U4186 (N_4186,N_2560,N_2264);
xnor U4187 (N_4187,N_417,N_3061);
nor U4188 (N_4188,N_2595,N_429);
and U4189 (N_4189,N_2791,N_1638);
or U4190 (N_4190,N_1421,N_2355);
xor U4191 (N_4191,N_215,N_527);
nor U4192 (N_4192,N_660,N_1927);
nor U4193 (N_4193,N_147,N_1129);
nor U4194 (N_4194,N_2554,N_1074);
and U4195 (N_4195,N_1138,N_1752);
and U4196 (N_4196,N_1489,N_1487);
and U4197 (N_4197,N_1793,N_1827);
xnor U4198 (N_4198,N_1571,N_2579);
or U4199 (N_4199,N_2826,N_850);
xor U4200 (N_4200,N_2800,N_347);
or U4201 (N_4201,N_1867,N_2976);
and U4202 (N_4202,N_2617,N_1357);
nand U4203 (N_4203,N_1533,N_2565);
or U4204 (N_4204,N_387,N_2679);
or U4205 (N_4205,N_1560,N_812);
xnor U4206 (N_4206,N_1076,N_148);
and U4207 (N_4207,N_2277,N_2294);
xnor U4208 (N_4208,N_2250,N_6);
xnor U4209 (N_4209,N_2084,N_2089);
and U4210 (N_4210,N_2282,N_357);
xnor U4211 (N_4211,N_18,N_1488);
or U4212 (N_4212,N_956,N_2310);
nand U4213 (N_4213,N_1917,N_917);
xnor U4214 (N_4214,N_186,N_214);
and U4215 (N_4215,N_1301,N_729);
or U4216 (N_4216,N_894,N_838);
and U4217 (N_4217,N_2526,N_351);
and U4218 (N_4218,N_47,N_1463);
and U4219 (N_4219,N_937,N_2854);
nor U4220 (N_4220,N_1313,N_1010);
and U4221 (N_4221,N_732,N_2623);
nand U4222 (N_4222,N_708,N_827);
or U4223 (N_4223,N_1855,N_3111);
and U4224 (N_4224,N_1389,N_2281);
nor U4225 (N_4225,N_625,N_2990);
nor U4226 (N_4226,N_2318,N_482);
nand U4227 (N_4227,N_2030,N_1199);
or U4228 (N_4228,N_49,N_2466);
or U4229 (N_4229,N_1814,N_1425);
xor U4230 (N_4230,N_2525,N_103);
nor U4231 (N_4231,N_983,N_1914);
or U4232 (N_4232,N_759,N_1889);
nand U4233 (N_4233,N_462,N_1332);
xor U4234 (N_4234,N_847,N_1290);
and U4235 (N_4235,N_2274,N_2925);
or U4236 (N_4236,N_2815,N_137);
xor U4237 (N_4237,N_2410,N_2196);
and U4238 (N_4238,N_821,N_2188);
nor U4239 (N_4239,N_1617,N_1289);
nor U4240 (N_4240,N_1584,N_2094);
and U4241 (N_4241,N_2258,N_2858);
and U4242 (N_4242,N_312,N_1603);
nand U4243 (N_4243,N_683,N_1744);
xnor U4244 (N_4244,N_2611,N_757);
nand U4245 (N_4245,N_1554,N_822);
nor U4246 (N_4246,N_2069,N_652);
xnor U4247 (N_4247,N_3055,N_1238);
or U4248 (N_4248,N_935,N_115);
nor U4249 (N_4249,N_2479,N_248);
nor U4250 (N_4250,N_1990,N_634);
or U4251 (N_4251,N_3048,N_2148);
xor U4252 (N_4252,N_1954,N_159);
nand U4253 (N_4253,N_170,N_83);
nor U4254 (N_4254,N_2044,N_1737);
or U4255 (N_4255,N_3101,N_2167);
xor U4256 (N_4256,N_2823,N_2291);
or U4257 (N_4257,N_1282,N_1467);
or U4258 (N_4258,N_1750,N_2344);
or U4259 (N_4259,N_1615,N_2658);
nor U4260 (N_4260,N_1760,N_376);
xor U4261 (N_4261,N_407,N_1869);
and U4262 (N_4262,N_914,N_1513);
and U4263 (N_4263,N_1736,N_1108);
xnor U4264 (N_4264,N_2081,N_2606);
xnor U4265 (N_4265,N_677,N_272);
xnor U4266 (N_4266,N_2958,N_2666);
and U4267 (N_4267,N_1252,N_352);
xor U4268 (N_4268,N_2223,N_2566);
nor U4269 (N_4269,N_2411,N_1677);
or U4270 (N_4270,N_560,N_11);
or U4271 (N_4271,N_557,N_2372);
nor U4272 (N_4272,N_615,N_136);
nor U4273 (N_4273,N_2232,N_2406);
or U4274 (N_4274,N_1733,N_1279);
nor U4275 (N_4275,N_1170,N_2882);
or U4276 (N_4276,N_1326,N_1094);
or U4277 (N_4277,N_1331,N_2025);
or U4278 (N_4278,N_1258,N_2014);
nand U4279 (N_4279,N_2780,N_2970);
xnor U4280 (N_4280,N_720,N_257);
xor U4281 (N_4281,N_961,N_2774);
or U4282 (N_4282,N_3114,N_2622);
nor U4283 (N_4283,N_1996,N_879);
and U4284 (N_4284,N_2333,N_858);
and U4285 (N_4285,N_610,N_1932);
or U4286 (N_4286,N_2241,N_456);
xor U4287 (N_4287,N_1529,N_2305);
nor U4288 (N_4288,N_2491,N_1414);
and U4289 (N_4289,N_190,N_3026);
nand U4290 (N_4290,N_1551,N_368);
or U4291 (N_4291,N_1516,N_719);
xor U4292 (N_4292,N_947,N_1797);
or U4293 (N_4293,N_135,N_1062);
nand U4294 (N_4294,N_1764,N_3);
xor U4295 (N_4295,N_2311,N_2596);
xnor U4296 (N_4296,N_1218,N_1178);
xor U4297 (N_4297,N_1510,N_2810);
nand U4298 (N_4298,N_2630,N_1416);
nor U4299 (N_4299,N_101,N_574);
and U4300 (N_4300,N_709,N_1649);
xor U4301 (N_4301,N_1547,N_2864);
or U4302 (N_4302,N_1823,N_12);
nand U4303 (N_4303,N_1166,N_1172);
xnor U4304 (N_4304,N_2801,N_1984);
or U4305 (N_4305,N_2929,N_1433);
xor U4306 (N_4306,N_321,N_17);
nand U4307 (N_4307,N_2334,N_1755);
or U4308 (N_4308,N_3087,N_303);
nand U4309 (N_4309,N_2297,N_2819);
nor U4310 (N_4310,N_1368,N_1619);
xnor U4311 (N_4311,N_114,N_3077);
or U4312 (N_4312,N_1097,N_1358);
or U4313 (N_4313,N_2248,N_1253);
nor U4314 (N_4314,N_2068,N_3104);
nor U4315 (N_4315,N_55,N_1850);
and U4316 (N_4316,N_2273,N_1948);
nor U4317 (N_4317,N_1060,N_1083);
or U4318 (N_4318,N_2088,N_3013);
and U4319 (N_4319,N_967,N_3051);
nor U4320 (N_4320,N_2003,N_707);
nand U4321 (N_4321,N_2283,N_51);
or U4322 (N_4322,N_1546,N_859);
or U4323 (N_4323,N_839,N_548);
nand U4324 (N_4324,N_365,N_1303);
and U4325 (N_4325,N_2734,N_782);
and U4326 (N_4326,N_181,N_2393);
nor U4327 (N_4327,N_153,N_221);
nor U4328 (N_4328,N_1400,N_87);
or U4329 (N_4329,N_424,N_577);
or U4330 (N_4330,N_835,N_1788);
nand U4331 (N_4331,N_1298,N_591);
nand U4332 (N_4332,N_2723,N_576);
nand U4333 (N_4333,N_1610,N_2676);
or U4334 (N_4334,N_86,N_3094);
or U4335 (N_4335,N_1681,N_282);
xnor U4336 (N_4336,N_1302,N_1388);
or U4337 (N_4337,N_642,N_980);
xor U4338 (N_4338,N_771,N_2270);
nand U4339 (N_4339,N_118,N_143);
nor U4340 (N_4340,N_2341,N_242);
nand U4341 (N_4341,N_2569,N_175);
and U4342 (N_4342,N_3085,N_1538);
or U4343 (N_4343,N_158,N_1871);
nand U4344 (N_4344,N_2564,N_2104);
and U4345 (N_4345,N_394,N_2741);
nand U4346 (N_4346,N_285,N_747);
nor U4347 (N_4347,N_673,N_565);
xor U4348 (N_4348,N_1147,N_760);
or U4349 (N_4349,N_2507,N_439);
or U4350 (N_4350,N_2145,N_1998);
nor U4351 (N_4351,N_2827,N_2996);
or U4352 (N_4352,N_2698,N_140);
nand U4353 (N_4353,N_1065,N_1344);
or U4354 (N_4354,N_1672,N_509);
and U4355 (N_4355,N_382,N_2492);
nor U4356 (N_4356,N_1558,N_171);
nand U4357 (N_4357,N_1612,N_2313);
nor U4358 (N_4358,N_2905,N_3021);
xor U4359 (N_4359,N_16,N_3088);
nor U4360 (N_4360,N_3017,N_671);
nor U4361 (N_4361,N_1587,N_2568);
and U4362 (N_4362,N_122,N_2496);
and U4363 (N_4363,N_2430,N_1390);
xor U4364 (N_4364,N_2659,N_1116);
and U4365 (N_4365,N_2165,N_290);
xnor U4366 (N_4366,N_2062,N_2873);
nor U4367 (N_4367,N_1235,N_1112);
and U4368 (N_4368,N_2625,N_2809);
nand U4369 (N_4369,N_390,N_1103);
nand U4370 (N_4370,N_1361,N_1695);
or U4371 (N_4371,N_2380,N_1240);
nand U4372 (N_4372,N_1475,N_2114);
nor U4373 (N_4373,N_2783,N_487);
and U4374 (N_4374,N_2391,N_1173);
xor U4375 (N_4375,N_2189,N_593);
nand U4376 (N_4376,N_251,N_156);
nand U4377 (N_4377,N_617,N_2146);
and U4378 (N_4378,N_2446,N_998);
and U4379 (N_4379,N_1050,N_1401);
nor U4380 (N_4380,N_1879,N_1625);
nand U4381 (N_4381,N_497,N_931);
nand U4382 (N_4382,N_1545,N_75);
xor U4383 (N_4383,N_2607,N_1209);
and U4384 (N_4384,N_511,N_8);
xnor U4385 (N_4385,N_1490,N_2985);
xnor U4386 (N_4386,N_519,N_834);
nand U4387 (N_4387,N_2919,N_1518);
or U4388 (N_4388,N_575,N_1206);
and U4389 (N_4389,N_590,N_587);
nand U4390 (N_4390,N_1104,N_2629);
and U4391 (N_4391,N_3011,N_1962);
nand U4392 (N_4392,N_1008,N_363);
xnor U4393 (N_4393,N_353,N_1459);
or U4394 (N_4394,N_2382,N_1082);
xnor U4395 (N_4395,N_408,N_2900);
and U4396 (N_4396,N_2408,N_1654);
nand U4397 (N_4397,N_1120,N_2182);
nand U4398 (N_4398,N_1305,N_629);
and U4399 (N_4399,N_1943,N_1691);
nor U4400 (N_4400,N_2442,N_2142);
or U4401 (N_4401,N_1480,N_2219);
nand U4402 (N_4402,N_14,N_2922);
xor U4403 (N_4403,N_1156,N_1134);
nor U4404 (N_4404,N_2386,N_289);
nand U4405 (N_4405,N_523,N_2143);
nor U4406 (N_4406,N_2704,N_1665);
or U4407 (N_4407,N_1407,N_2638);
nor U4408 (N_4408,N_900,N_1865);
nor U4409 (N_4409,N_2428,N_1450);
or U4410 (N_4410,N_602,N_1053);
xnor U4411 (N_4411,N_1152,N_286);
and U4412 (N_4412,N_1928,N_544);
and U4413 (N_4413,N_1315,N_444);
or U4414 (N_4414,N_1701,N_1102);
nor U4415 (N_4415,N_157,N_443);
nand U4416 (N_4416,N_53,N_1604);
and U4417 (N_4417,N_1087,N_1193);
xor U4418 (N_4418,N_3036,N_2843);
or U4419 (N_4419,N_1096,N_3072);
or U4420 (N_4420,N_3025,N_1980);
nand U4421 (N_4421,N_184,N_1000);
nor U4422 (N_4422,N_3073,N_1442);
xor U4423 (N_4423,N_1220,N_994);
xor U4424 (N_4424,N_10,N_2242);
or U4425 (N_4425,N_3050,N_1690);
nor U4426 (N_4426,N_2846,N_78);
nand U4427 (N_4427,N_2377,N_1277);
nand U4428 (N_4428,N_2736,N_656);
xnor U4429 (N_4429,N_1181,N_3069);
xnor U4430 (N_4430,N_2711,N_877);
nor U4431 (N_4431,N_2309,N_2581);
nor U4432 (N_4432,N_751,N_2041);
nor U4433 (N_4433,N_944,N_1024);
or U4434 (N_4434,N_2501,N_2262);
xor U4435 (N_4435,N_1523,N_2213);
or U4436 (N_4436,N_2000,N_831);
and U4437 (N_4437,N_2519,N_2828);
or U4438 (N_4438,N_2118,N_779);
nor U4439 (N_4439,N_1231,N_992);
nand U4440 (N_4440,N_853,N_1960);
xor U4441 (N_4441,N_1809,N_1904);
nand U4442 (N_4442,N_2661,N_2018);
nand U4443 (N_4443,N_2943,N_2296);
nand U4444 (N_4444,N_2721,N_1995);
nand U4445 (N_4445,N_1556,N_2195);
nor U4446 (N_4446,N_607,N_249);
and U4447 (N_4447,N_138,N_395);
and U4448 (N_4448,N_438,N_1687);
or U4449 (N_4449,N_1713,N_2284);
and U4450 (N_4450,N_358,N_2805);
nor U4451 (N_4451,N_1474,N_1189);
xor U4452 (N_4452,N_1549,N_44);
xor U4453 (N_4453,N_2179,N_1003);
and U4454 (N_4454,N_2307,N_2994);
or U4455 (N_4455,N_622,N_912);
nor U4456 (N_4456,N_965,N_1217);
and U4457 (N_4457,N_59,N_2868);
xor U4458 (N_4458,N_3054,N_849);
xnor U4459 (N_4459,N_2029,N_2259);
nand U4460 (N_4460,N_580,N_2551);
nor U4461 (N_4461,N_1071,N_2872);
xnor U4462 (N_4462,N_669,N_2079);
nor U4463 (N_4463,N_1482,N_2928);
nand U4464 (N_4464,N_2346,N_2448);
nor U4465 (N_4465,N_1605,N_1575);
xor U4466 (N_4466,N_1894,N_1422);
and U4467 (N_4467,N_1559,N_281);
and U4468 (N_4468,N_2384,N_1833);
nand U4469 (N_4469,N_322,N_2883);
nor U4470 (N_4470,N_777,N_3056);
and U4471 (N_4471,N_1285,N_466);
or U4472 (N_4472,N_884,N_2959);
nand U4473 (N_4473,N_1415,N_2975);
xnor U4474 (N_4474,N_3062,N_986);
and U4475 (N_4475,N_939,N_823);
nand U4476 (N_4476,N_579,N_2279);
and U4477 (N_4477,N_2444,N_2150);
or U4478 (N_4478,N_1035,N_2054);
nor U4479 (N_4479,N_2139,N_61);
or U4480 (N_4480,N_1257,N_2154);
xnor U4481 (N_4481,N_1562,N_2876);
nand U4482 (N_4482,N_252,N_1925);
and U4483 (N_4483,N_1725,N_1364);
xor U4484 (N_4484,N_659,N_701);
xnor U4485 (N_4485,N_48,N_2563);
and U4486 (N_4486,N_860,N_1164);
nand U4487 (N_4487,N_324,N_2981);
xnor U4488 (N_4488,N_2742,N_2134);
and U4489 (N_4489,N_1622,N_1812);
nand U4490 (N_4490,N_2859,N_2785);
or U4491 (N_4491,N_154,N_1406);
xnor U4492 (N_4492,N_920,N_946);
and U4493 (N_4493,N_1597,N_1762);
or U4494 (N_4494,N_2633,N_2515);
and U4495 (N_4495,N_2394,N_819);
and U4496 (N_4496,N_246,N_1471);
nand U4497 (N_4497,N_2555,N_2775);
nand U4498 (N_4498,N_1776,N_1525);
nor U4499 (N_4499,N_951,N_459);
and U4500 (N_4500,N_2811,N_166);
or U4501 (N_4501,N_558,N_379);
nor U4502 (N_4502,N_292,N_1745);
and U4503 (N_4503,N_40,N_288);
nor U4504 (N_4504,N_1895,N_304);
nand U4505 (N_4505,N_478,N_3038);
nand U4506 (N_4506,N_1353,N_1595);
nor U4507 (N_4507,N_2755,N_2108);
nand U4508 (N_4508,N_1063,N_2119);
or U4509 (N_4509,N_3090,N_645);
and U4510 (N_4510,N_2197,N_2968);
nor U4511 (N_4511,N_1337,N_2914);
or U4512 (N_4512,N_871,N_1500);
xor U4513 (N_4513,N_1593,N_1741);
xor U4514 (N_4514,N_2627,N_923);
or U4515 (N_4515,N_2107,N_746);
or U4516 (N_4516,N_1468,N_1438);
and U4517 (N_4517,N_234,N_852);
nand U4518 (N_4518,N_434,N_2793);
or U4519 (N_4519,N_636,N_489);
or U4520 (N_4520,N_2349,N_2231);
nand U4521 (N_4521,N_2745,N_1703);
nor U4522 (N_4522,N_855,N_1655);
and U4523 (N_4523,N_1413,N_1365);
nand U4524 (N_4524,N_123,N_1330);
and U4525 (N_4525,N_3115,N_1694);
xor U4526 (N_4526,N_1387,N_1300);
xnor U4527 (N_4527,N_63,N_71);
nor U4528 (N_4528,N_2449,N_627);
nor U4529 (N_4529,N_1169,N_2317);
nand U4530 (N_4530,N_1712,N_3109);
xor U4531 (N_4531,N_1107,N_2543);
xnor U4532 (N_4532,N_2845,N_2712);
or U4533 (N_4533,N_2034,N_226);
nor U4534 (N_4534,N_840,N_2977);
nor U4535 (N_4535,N_1935,N_765);
nor U4536 (N_4536,N_2141,N_2714);
xnor U4537 (N_4537,N_402,N_258);
nor U4538 (N_4538,N_196,N_29);
nor U4539 (N_4539,N_447,N_3003);
or U4540 (N_4540,N_217,N_524);
and U4541 (N_4541,N_1631,N_1069);
or U4542 (N_4542,N_1573,N_128);
nor U4543 (N_4543,N_2228,N_1084);
nand U4544 (N_4544,N_218,N_1974);
nand U4545 (N_4545,N_2558,N_2475);
xor U4546 (N_4546,N_832,N_1245);
xor U4547 (N_4547,N_758,N_1803);
nor U4548 (N_4548,N_2005,N_348);
and U4549 (N_4549,N_2337,N_526);
nand U4550 (N_4550,N_534,N_960);
or U4551 (N_4551,N_2621,N_2354);
nor U4552 (N_4552,N_2252,N_1785);
nor U4553 (N_4553,N_431,N_921);
and U4554 (N_4554,N_81,N_1212);
nor U4555 (N_4555,N_737,N_2616);
xnor U4556 (N_4556,N_1606,N_2980);
nand U4557 (N_4557,N_220,N_1624);
xor U4558 (N_4558,N_2849,N_1763);
nand U4559 (N_4559,N_2539,N_496);
and U4560 (N_4560,N_595,N_1770);
xor U4561 (N_4561,N_2973,N_201);
nand U4562 (N_4562,N_2480,N_2342);
nor U4563 (N_4563,N_2867,N_2747);
or U4564 (N_4564,N_2891,N_2530);
nor U4565 (N_4565,N_2478,N_1608);
and U4566 (N_4566,N_930,N_772);
nand U4567 (N_4567,N_2061,N_1165);
xnor U4568 (N_4568,N_1190,N_2574);
nand U4569 (N_4569,N_97,N_1423);
nor U4570 (N_4570,N_239,N_1742);
and U4571 (N_4571,N_1645,N_2656);
xnor U4572 (N_4572,N_769,N_2903);
or U4573 (N_4573,N_1620,N_1896);
or U4574 (N_4574,N_169,N_2759);
or U4575 (N_4575,N_2257,N_1348);
nand U4576 (N_4576,N_2798,N_2688);
or U4577 (N_4577,N_1817,N_2332);
nor U4578 (N_4578,N_2572,N_1118);
nor U4579 (N_4579,N_2421,N_2415);
and U4580 (N_4580,N_1127,N_1048);
or U4581 (N_4581,N_1022,N_2879);
nor U4582 (N_4582,N_2037,N_2957);
nor U4583 (N_4583,N_2237,N_2111);
or U4584 (N_4584,N_121,N_2998);
and U4585 (N_4585,N_1576,N_1242);
xor U4586 (N_4586,N_2934,N_1872);
nor U4587 (N_4587,N_1992,N_2693);
or U4588 (N_4588,N_327,N_110);
nand U4589 (N_4589,N_679,N_2898);
xor U4590 (N_4590,N_1180,N_3102);
and U4591 (N_4591,N_726,N_1771);
or U4592 (N_4592,N_2893,N_805);
nand U4593 (N_4593,N_2825,N_881);
xnor U4594 (N_4594,N_1519,N_2762);
nor U4595 (N_4595,N_1007,N_2053);
and U4596 (N_4596,N_2848,N_2601);
nand U4597 (N_4597,N_2619,N_1659);
or U4598 (N_4598,N_1377,N_1386);
xor U4599 (N_4599,N_2498,N_240);
nand U4600 (N_4600,N_2663,N_1032);
and U4601 (N_4601,N_2286,N_1494);
nand U4602 (N_4602,N_815,N_663);
or U4603 (N_4603,N_1275,N_2777);
or U4604 (N_4604,N_878,N_2571);
xor U4605 (N_4605,N_2590,N_1015);
or U4606 (N_4606,N_2861,N_2881);
nand U4607 (N_4607,N_1705,N_113);
xor U4608 (N_4608,N_274,N_2152);
xor U4609 (N_4609,N_2443,N_1678);
nand U4610 (N_4610,N_3029,N_555);
xor U4611 (N_4611,N_1052,N_1882);
and U4612 (N_4612,N_2694,N_1314);
nor U4613 (N_4613,N_2432,N_2115);
nor U4614 (N_4614,N_1001,N_2413);
nand U4615 (N_4615,N_144,N_1716);
nand U4616 (N_4616,N_630,N_2874);
nand U4617 (N_4617,N_1373,N_1370);
and U4618 (N_4618,N_1930,N_3083);
xnor U4619 (N_4619,N_1633,N_1953);
nor U4620 (N_4620,N_366,N_2450);
nor U4621 (N_4621,N_433,N_326);
nand U4622 (N_4622,N_3071,N_535);
and U4623 (N_4623,N_1972,N_541);
and U4624 (N_4624,N_814,N_112);
or U4625 (N_4625,N_2795,N_512);
or U4626 (N_4626,N_1552,N_388);
or U4627 (N_4627,N_1639,N_783);
nand U4628 (N_4628,N_88,N_475);
or U4629 (N_4629,N_1420,N_1588);
or U4630 (N_4630,N_1844,N_1843);
nand U4631 (N_4631,N_2374,N_2439);
nand U4632 (N_4632,N_1130,N_270);
and U4633 (N_4633,N_2320,N_2635);
xnor U4634 (N_4634,N_1470,N_2065);
and U4635 (N_4635,N_514,N_2102);
nor U4636 (N_4636,N_2381,N_500);
and U4637 (N_4637,N_654,N_333);
nand U4638 (N_4638,N_981,N_2857);
and U4639 (N_4639,N_664,N_1460);
nor U4640 (N_4640,N_192,N_2093);
nor U4641 (N_4641,N_2707,N_30);
nor U4642 (N_4642,N_2686,N_2177);
or U4643 (N_4643,N_1046,N_2691);
nand U4644 (N_4644,N_1728,N_3067);
xor U4645 (N_4645,N_319,N_485);
nand U4646 (N_4646,N_1589,N_2933);
nand U4647 (N_4647,N_2441,N_2389);
nand U4648 (N_4648,N_1508,N_1751);
and U4649 (N_4649,N_3024,N_538);
nor U4650 (N_4650,N_2500,N_1306);
xnor U4651 (N_4651,N_1229,N_867);
nand U4652 (N_4652,N_1868,N_1861);
nand U4653 (N_4653,N_749,N_256);
nor U4654 (N_4654,N_314,N_793);
nand U4655 (N_4655,N_2024,N_2626);
nand U4656 (N_4656,N_2375,N_1901);
xor U4657 (N_4657,N_794,N_307);
or U4658 (N_4658,N_432,N_399);
nor U4659 (N_4659,N_2675,N_2708);
xor U4660 (N_4660,N_2484,N_3004);
nand U4661 (N_4661,N_1155,N_1897);
and U4662 (N_4662,N_1636,N_2451);
and U4663 (N_4663,N_3098,N_313);
and U4664 (N_4664,N_98,N_1735);
xor U4665 (N_4665,N_1497,N_1078);
nor U4666 (N_4666,N_2272,N_731);
nor U4667 (N_4667,N_916,N_797);
and U4668 (N_4668,N_1920,N_1929);
and U4669 (N_4669,N_1969,N_2217);
or U4670 (N_4670,N_189,N_1239);
and U4671 (N_4671,N_3063,N_2163);
and U4672 (N_4672,N_2269,N_826);
xnor U4673 (N_4673,N_2233,N_1734);
xnor U4674 (N_4674,N_734,N_2856);
xor U4675 (N_4675,N_2116,N_2109);
xnor U4676 (N_4676,N_570,N_41);
nor U4677 (N_4677,N_1372,N_1184);
xor U4678 (N_4678,N_1028,N_1200);
nor U4679 (N_4679,N_1381,N_66);
nor U4680 (N_4680,N_1601,N_1014);
nand U4681 (N_4681,N_1049,N_1195);
or U4682 (N_4682,N_1993,N_3030);
nand U4683 (N_4683,N_335,N_1729);
or U4684 (N_4684,N_177,N_2455);
xnor U4685 (N_4685,N_940,N_2214);
nand U4686 (N_4686,N_1098,N_3121);
and U4687 (N_4687,N_205,N_1529);
and U4688 (N_4688,N_3124,N_1023);
nor U4689 (N_4689,N_1167,N_394);
nor U4690 (N_4690,N_932,N_750);
nand U4691 (N_4691,N_1251,N_2118);
or U4692 (N_4692,N_2563,N_2711);
or U4693 (N_4693,N_3033,N_1765);
nand U4694 (N_4694,N_1531,N_226);
nand U4695 (N_4695,N_1859,N_1327);
xnor U4696 (N_4696,N_2514,N_2134);
xnor U4697 (N_4697,N_1995,N_2154);
xor U4698 (N_4698,N_1227,N_1717);
or U4699 (N_4699,N_1941,N_1327);
or U4700 (N_4700,N_547,N_883);
nor U4701 (N_4701,N_153,N_2652);
xnor U4702 (N_4702,N_1849,N_2833);
or U4703 (N_4703,N_2822,N_55);
xnor U4704 (N_4704,N_548,N_226);
nor U4705 (N_4705,N_1562,N_2272);
xnor U4706 (N_4706,N_1144,N_754);
xor U4707 (N_4707,N_2957,N_869);
and U4708 (N_4708,N_1847,N_1247);
and U4709 (N_4709,N_1816,N_2644);
or U4710 (N_4710,N_843,N_2385);
nor U4711 (N_4711,N_2970,N_1645);
xor U4712 (N_4712,N_694,N_2845);
and U4713 (N_4713,N_2836,N_1416);
and U4714 (N_4714,N_2543,N_1816);
and U4715 (N_4715,N_2217,N_2009);
nand U4716 (N_4716,N_1013,N_2511);
nand U4717 (N_4717,N_1400,N_1026);
or U4718 (N_4718,N_11,N_2674);
nand U4719 (N_4719,N_1790,N_2306);
nand U4720 (N_4720,N_1338,N_276);
nand U4721 (N_4721,N_448,N_645);
or U4722 (N_4722,N_2197,N_582);
nand U4723 (N_4723,N_167,N_2286);
and U4724 (N_4724,N_2176,N_1306);
xor U4725 (N_4725,N_2150,N_2043);
and U4726 (N_4726,N_590,N_2880);
xnor U4727 (N_4727,N_2294,N_124);
nand U4728 (N_4728,N_894,N_2339);
xnor U4729 (N_4729,N_1496,N_2325);
nor U4730 (N_4730,N_685,N_2530);
xnor U4731 (N_4731,N_1416,N_604);
nor U4732 (N_4732,N_1450,N_202);
xor U4733 (N_4733,N_481,N_115);
or U4734 (N_4734,N_1350,N_2383);
nor U4735 (N_4735,N_2294,N_599);
nand U4736 (N_4736,N_2222,N_1304);
and U4737 (N_4737,N_2796,N_912);
nor U4738 (N_4738,N_1717,N_227);
or U4739 (N_4739,N_2747,N_20);
nor U4740 (N_4740,N_917,N_585);
nand U4741 (N_4741,N_1008,N_105);
nor U4742 (N_4742,N_6,N_2116);
and U4743 (N_4743,N_2599,N_1041);
nand U4744 (N_4744,N_721,N_678);
nand U4745 (N_4745,N_1185,N_2051);
and U4746 (N_4746,N_367,N_96);
xor U4747 (N_4747,N_678,N_538);
or U4748 (N_4748,N_2069,N_613);
nand U4749 (N_4749,N_282,N_1218);
nor U4750 (N_4750,N_1060,N_1993);
nand U4751 (N_4751,N_738,N_2783);
and U4752 (N_4752,N_2567,N_2741);
nor U4753 (N_4753,N_2181,N_689);
nand U4754 (N_4754,N_1686,N_408);
xor U4755 (N_4755,N_2531,N_1735);
and U4756 (N_4756,N_1715,N_1406);
nor U4757 (N_4757,N_432,N_2053);
and U4758 (N_4758,N_1837,N_2406);
or U4759 (N_4759,N_1928,N_1401);
nand U4760 (N_4760,N_457,N_384);
xor U4761 (N_4761,N_1227,N_1298);
or U4762 (N_4762,N_917,N_1415);
or U4763 (N_4763,N_2189,N_790);
or U4764 (N_4764,N_329,N_2453);
xor U4765 (N_4765,N_618,N_1768);
or U4766 (N_4766,N_1432,N_1768);
nor U4767 (N_4767,N_1563,N_1570);
or U4768 (N_4768,N_1678,N_444);
nand U4769 (N_4769,N_454,N_1179);
and U4770 (N_4770,N_2,N_1317);
xnor U4771 (N_4771,N_533,N_2919);
or U4772 (N_4772,N_1055,N_1715);
xor U4773 (N_4773,N_955,N_1312);
and U4774 (N_4774,N_499,N_391);
xnor U4775 (N_4775,N_1527,N_3002);
xnor U4776 (N_4776,N_1909,N_1387);
and U4777 (N_4777,N_845,N_2509);
and U4778 (N_4778,N_784,N_1094);
and U4779 (N_4779,N_420,N_2539);
xor U4780 (N_4780,N_1743,N_2977);
xor U4781 (N_4781,N_2271,N_1074);
and U4782 (N_4782,N_1163,N_1636);
nor U4783 (N_4783,N_913,N_2500);
or U4784 (N_4784,N_192,N_68);
nand U4785 (N_4785,N_2152,N_737);
and U4786 (N_4786,N_1417,N_2014);
xnor U4787 (N_4787,N_213,N_2709);
and U4788 (N_4788,N_2984,N_1034);
xnor U4789 (N_4789,N_1360,N_2662);
or U4790 (N_4790,N_1343,N_1699);
and U4791 (N_4791,N_2969,N_2973);
xor U4792 (N_4792,N_2318,N_1974);
xor U4793 (N_4793,N_1570,N_1218);
and U4794 (N_4794,N_296,N_399);
or U4795 (N_4795,N_753,N_381);
and U4796 (N_4796,N_893,N_2773);
and U4797 (N_4797,N_370,N_599);
nand U4798 (N_4798,N_642,N_2739);
nand U4799 (N_4799,N_466,N_1097);
and U4800 (N_4800,N_2678,N_1254);
xnor U4801 (N_4801,N_2869,N_3061);
or U4802 (N_4802,N_1057,N_793);
nand U4803 (N_4803,N_1832,N_1011);
or U4804 (N_4804,N_1799,N_198);
and U4805 (N_4805,N_2918,N_700);
or U4806 (N_4806,N_2115,N_103);
or U4807 (N_4807,N_635,N_761);
nor U4808 (N_4808,N_1732,N_2563);
xnor U4809 (N_4809,N_413,N_1173);
xor U4810 (N_4810,N_2074,N_2764);
xnor U4811 (N_4811,N_629,N_1384);
nand U4812 (N_4812,N_138,N_733);
nand U4813 (N_4813,N_1063,N_2775);
xor U4814 (N_4814,N_1618,N_28);
nand U4815 (N_4815,N_2101,N_167);
and U4816 (N_4816,N_2553,N_3030);
xor U4817 (N_4817,N_2049,N_1720);
nand U4818 (N_4818,N_478,N_66);
nand U4819 (N_4819,N_884,N_363);
or U4820 (N_4820,N_2859,N_1156);
xnor U4821 (N_4821,N_711,N_1603);
nand U4822 (N_4822,N_2730,N_3087);
and U4823 (N_4823,N_1974,N_2196);
xnor U4824 (N_4824,N_1150,N_1903);
nand U4825 (N_4825,N_1765,N_2714);
nor U4826 (N_4826,N_1015,N_1090);
nor U4827 (N_4827,N_2303,N_1806);
and U4828 (N_4828,N_2414,N_729);
or U4829 (N_4829,N_2200,N_1901);
xnor U4830 (N_4830,N_567,N_530);
xnor U4831 (N_4831,N_874,N_2870);
nor U4832 (N_4832,N_2821,N_2848);
nand U4833 (N_4833,N_3111,N_599);
nor U4834 (N_4834,N_3001,N_1557);
nand U4835 (N_4835,N_2036,N_2573);
or U4836 (N_4836,N_1402,N_501);
nand U4837 (N_4837,N_1595,N_356);
nor U4838 (N_4838,N_556,N_2128);
and U4839 (N_4839,N_1840,N_672);
and U4840 (N_4840,N_2377,N_771);
or U4841 (N_4841,N_1955,N_244);
or U4842 (N_4842,N_1922,N_2029);
nand U4843 (N_4843,N_1582,N_2398);
or U4844 (N_4844,N_222,N_162);
or U4845 (N_4845,N_1560,N_599);
or U4846 (N_4846,N_2170,N_1960);
nand U4847 (N_4847,N_644,N_2332);
nand U4848 (N_4848,N_1413,N_194);
xnor U4849 (N_4849,N_1585,N_2397);
xnor U4850 (N_4850,N_2700,N_1134);
nor U4851 (N_4851,N_1837,N_482);
nand U4852 (N_4852,N_3123,N_2070);
nand U4853 (N_4853,N_1936,N_2382);
and U4854 (N_4854,N_433,N_1199);
or U4855 (N_4855,N_1355,N_2954);
xnor U4856 (N_4856,N_860,N_2215);
nand U4857 (N_4857,N_1547,N_1619);
xor U4858 (N_4858,N_889,N_2823);
nand U4859 (N_4859,N_2625,N_2004);
nand U4860 (N_4860,N_532,N_1077);
xor U4861 (N_4861,N_2241,N_1820);
nand U4862 (N_4862,N_853,N_2775);
or U4863 (N_4863,N_2237,N_804);
xor U4864 (N_4864,N_1282,N_902);
and U4865 (N_4865,N_1079,N_1060);
xor U4866 (N_4866,N_613,N_15);
nand U4867 (N_4867,N_1453,N_2017);
xor U4868 (N_4868,N_380,N_1827);
or U4869 (N_4869,N_589,N_592);
nor U4870 (N_4870,N_2987,N_1957);
nor U4871 (N_4871,N_681,N_352);
and U4872 (N_4872,N_3031,N_313);
nor U4873 (N_4873,N_2199,N_313);
xnor U4874 (N_4874,N_3077,N_449);
or U4875 (N_4875,N_2747,N_506);
and U4876 (N_4876,N_1490,N_2325);
xor U4877 (N_4877,N_1313,N_805);
xor U4878 (N_4878,N_1652,N_2037);
nand U4879 (N_4879,N_859,N_2068);
nor U4880 (N_4880,N_2007,N_1436);
and U4881 (N_4881,N_2074,N_1542);
nor U4882 (N_4882,N_2652,N_638);
nand U4883 (N_4883,N_1069,N_2820);
nand U4884 (N_4884,N_358,N_1660);
or U4885 (N_4885,N_207,N_532);
and U4886 (N_4886,N_1379,N_2371);
nand U4887 (N_4887,N_2238,N_2739);
nor U4888 (N_4888,N_1846,N_405);
nor U4889 (N_4889,N_662,N_959);
xnor U4890 (N_4890,N_1316,N_474);
nor U4891 (N_4891,N_664,N_2073);
nand U4892 (N_4892,N_162,N_59);
and U4893 (N_4893,N_2477,N_2745);
or U4894 (N_4894,N_113,N_932);
or U4895 (N_4895,N_2900,N_610);
xnor U4896 (N_4896,N_2864,N_1816);
nor U4897 (N_4897,N_2150,N_696);
nor U4898 (N_4898,N_1336,N_1219);
nand U4899 (N_4899,N_2248,N_234);
xnor U4900 (N_4900,N_1770,N_748);
nor U4901 (N_4901,N_2,N_2479);
nand U4902 (N_4902,N_2150,N_2962);
xnor U4903 (N_4903,N_2750,N_374);
xor U4904 (N_4904,N_1895,N_1845);
and U4905 (N_4905,N_2403,N_1761);
nand U4906 (N_4906,N_842,N_2560);
xnor U4907 (N_4907,N_1475,N_2681);
nand U4908 (N_4908,N_1471,N_740);
nand U4909 (N_4909,N_1009,N_691);
nand U4910 (N_4910,N_2328,N_1993);
nor U4911 (N_4911,N_2708,N_2484);
and U4912 (N_4912,N_2502,N_1641);
nand U4913 (N_4913,N_570,N_831);
nor U4914 (N_4914,N_2835,N_1687);
nor U4915 (N_4915,N_242,N_501);
nor U4916 (N_4916,N_1631,N_432);
xnor U4917 (N_4917,N_1390,N_2199);
nand U4918 (N_4918,N_736,N_1461);
xor U4919 (N_4919,N_1241,N_2106);
and U4920 (N_4920,N_2486,N_855);
and U4921 (N_4921,N_2438,N_1567);
nand U4922 (N_4922,N_2889,N_1807);
nor U4923 (N_4923,N_1259,N_318);
and U4924 (N_4924,N_1562,N_2831);
or U4925 (N_4925,N_948,N_1750);
nand U4926 (N_4926,N_840,N_972);
or U4927 (N_4927,N_2045,N_1215);
or U4928 (N_4928,N_2957,N_2021);
xnor U4929 (N_4929,N_2436,N_384);
nand U4930 (N_4930,N_1168,N_2252);
nor U4931 (N_4931,N_1837,N_1327);
nor U4932 (N_4932,N_2308,N_37);
or U4933 (N_4933,N_2840,N_2599);
xnor U4934 (N_4934,N_995,N_2174);
and U4935 (N_4935,N_2326,N_3030);
or U4936 (N_4936,N_2801,N_1632);
and U4937 (N_4937,N_2282,N_1041);
nand U4938 (N_4938,N_1668,N_2633);
or U4939 (N_4939,N_1788,N_179);
nor U4940 (N_4940,N_376,N_1007);
xnor U4941 (N_4941,N_8,N_1345);
and U4942 (N_4942,N_879,N_43);
xnor U4943 (N_4943,N_1197,N_2989);
nand U4944 (N_4944,N_2785,N_2367);
or U4945 (N_4945,N_2488,N_1434);
or U4946 (N_4946,N_925,N_2496);
nor U4947 (N_4947,N_910,N_2016);
and U4948 (N_4948,N_1960,N_2126);
nand U4949 (N_4949,N_1348,N_2523);
and U4950 (N_4950,N_1878,N_2825);
or U4951 (N_4951,N_522,N_15);
and U4952 (N_4952,N_223,N_2136);
or U4953 (N_4953,N_1184,N_3052);
nand U4954 (N_4954,N_2556,N_3047);
xnor U4955 (N_4955,N_101,N_1552);
or U4956 (N_4956,N_1627,N_1759);
nor U4957 (N_4957,N_3065,N_2945);
or U4958 (N_4958,N_990,N_634);
nor U4959 (N_4959,N_504,N_1501);
and U4960 (N_4960,N_576,N_3068);
or U4961 (N_4961,N_3064,N_119);
and U4962 (N_4962,N_2966,N_1824);
nand U4963 (N_4963,N_399,N_2466);
nor U4964 (N_4964,N_493,N_1749);
or U4965 (N_4965,N_1807,N_2020);
or U4966 (N_4966,N_1027,N_1143);
nand U4967 (N_4967,N_389,N_984);
or U4968 (N_4968,N_1135,N_2122);
and U4969 (N_4969,N_1248,N_1221);
or U4970 (N_4970,N_2924,N_1203);
nand U4971 (N_4971,N_2215,N_225);
nand U4972 (N_4972,N_1443,N_1553);
nand U4973 (N_4973,N_2318,N_2894);
nand U4974 (N_4974,N_410,N_2647);
nand U4975 (N_4975,N_2763,N_2308);
nor U4976 (N_4976,N_2003,N_652);
or U4977 (N_4977,N_1846,N_1314);
nand U4978 (N_4978,N_304,N_625);
and U4979 (N_4979,N_3050,N_1537);
xor U4980 (N_4980,N_275,N_363);
and U4981 (N_4981,N_1292,N_293);
nor U4982 (N_4982,N_3025,N_1348);
or U4983 (N_4983,N_2481,N_286);
nor U4984 (N_4984,N_2827,N_448);
xor U4985 (N_4985,N_2378,N_3118);
nor U4986 (N_4986,N_1837,N_1238);
nor U4987 (N_4987,N_2474,N_2945);
nand U4988 (N_4988,N_1805,N_447);
and U4989 (N_4989,N_2829,N_277);
xor U4990 (N_4990,N_626,N_2175);
nor U4991 (N_4991,N_1266,N_2901);
and U4992 (N_4992,N_1650,N_2058);
xor U4993 (N_4993,N_1863,N_3044);
and U4994 (N_4994,N_1318,N_527);
xor U4995 (N_4995,N_1070,N_2224);
nor U4996 (N_4996,N_2663,N_1729);
nand U4997 (N_4997,N_2712,N_315);
and U4998 (N_4998,N_2738,N_1228);
xor U4999 (N_4999,N_1838,N_1347);
nor U5000 (N_5000,N_218,N_2319);
xnor U5001 (N_5001,N_1281,N_1560);
and U5002 (N_5002,N_1502,N_558);
or U5003 (N_5003,N_2080,N_949);
nor U5004 (N_5004,N_1240,N_2459);
nor U5005 (N_5005,N_201,N_1519);
or U5006 (N_5006,N_0,N_1633);
nand U5007 (N_5007,N_2210,N_2770);
or U5008 (N_5008,N_3100,N_1569);
and U5009 (N_5009,N_1179,N_1622);
nand U5010 (N_5010,N_1802,N_277);
xnor U5011 (N_5011,N_1556,N_298);
nand U5012 (N_5012,N_1372,N_1861);
nand U5013 (N_5013,N_747,N_958);
or U5014 (N_5014,N_1204,N_178);
and U5015 (N_5015,N_1969,N_1376);
nand U5016 (N_5016,N_1428,N_3023);
and U5017 (N_5017,N_35,N_2109);
nor U5018 (N_5018,N_2203,N_765);
or U5019 (N_5019,N_373,N_2490);
or U5020 (N_5020,N_1774,N_1232);
or U5021 (N_5021,N_3091,N_1988);
or U5022 (N_5022,N_1070,N_2290);
nand U5023 (N_5023,N_1684,N_2847);
xnor U5024 (N_5024,N_2549,N_2938);
or U5025 (N_5025,N_1812,N_566);
nand U5026 (N_5026,N_19,N_1898);
nand U5027 (N_5027,N_1017,N_1792);
xor U5028 (N_5028,N_1462,N_2101);
nand U5029 (N_5029,N_1951,N_1720);
or U5030 (N_5030,N_1575,N_1369);
nand U5031 (N_5031,N_171,N_97);
xor U5032 (N_5032,N_509,N_1398);
nand U5033 (N_5033,N_2059,N_644);
xnor U5034 (N_5034,N_1010,N_207);
nor U5035 (N_5035,N_2124,N_635);
and U5036 (N_5036,N_1668,N_816);
nor U5037 (N_5037,N_2869,N_128);
nor U5038 (N_5038,N_697,N_1556);
nor U5039 (N_5039,N_1149,N_2701);
or U5040 (N_5040,N_2728,N_326);
nor U5041 (N_5041,N_798,N_2096);
or U5042 (N_5042,N_571,N_1068);
xnor U5043 (N_5043,N_113,N_2581);
or U5044 (N_5044,N_2467,N_25);
and U5045 (N_5045,N_917,N_844);
or U5046 (N_5046,N_1950,N_2481);
and U5047 (N_5047,N_2678,N_3058);
nand U5048 (N_5048,N_882,N_1037);
and U5049 (N_5049,N_1420,N_75);
nand U5050 (N_5050,N_666,N_1259);
xnor U5051 (N_5051,N_1525,N_2351);
or U5052 (N_5052,N_1050,N_1149);
nor U5053 (N_5053,N_2039,N_1015);
xnor U5054 (N_5054,N_2369,N_413);
or U5055 (N_5055,N_457,N_2059);
xnor U5056 (N_5056,N_54,N_1701);
and U5057 (N_5057,N_2359,N_895);
nor U5058 (N_5058,N_2158,N_1132);
nor U5059 (N_5059,N_2264,N_404);
nor U5060 (N_5060,N_576,N_747);
or U5061 (N_5061,N_446,N_1068);
nand U5062 (N_5062,N_411,N_498);
or U5063 (N_5063,N_1848,N_531);
nand U5064 (N_5064,N_371,N_2916);
nor U5065 (N_5065,N_773,N_1109);
nand U5066 (N_5066,N_1665,N_2926);
xnor U5067 (N_5067,N_931,N_1186);
or U5068 (N_5068,N_2489,N_493);
xnor U5069 (N_5069,N_2072,N_624);
xnor U5070 (N_5070,N_2673,N_20);
nor U5071 (N_5071,N_2097,N_2824);
nor U5072 (N_5072,N_1504,N_1513);
nor U5073 (N_5073,N_37,N_1032);
and U5074 (N_5074,N_2207,N_1621);
nand U5075 (N_5075,N_1827,N_661);
or U5076 (N_5076,N_2861,N_1808);
or U5077 (N_5077,N_1828,N_850);
and U5078 (N_5078,N_2727,N_2389);
nor U5079 (N_5079,N_414,N_272);
and U5080 (N_5080,N_1756,N_727);
nor U5081 (N_5081,N_3099,N_2969);
nand U5082 (N_5082,N_727,N_1077);
and U5083 (N_5083,N_1659,N_1817);
or U5084 (N_5084,N_369,N_208);
nor U5085 (N_5085,N_449,N_1882);
or U5086 (N_5086,N_806,N_1678);
and U5087 (N_5087,N_125,N_501);
and U5088 (N_5088,N_2146,N_2397);
nand U5089 (N_5089,N_349,N_2106);
xor U5090 (N_5090,N_2516,N_1480);
xor U5091 (N_5091,N_1428,N_670);
and U5092 (N_5092,N_976,N_2513);
xnor U5093 (N_5093,N_425,N_1088);
nor U5094 (N_5094,N_2785,N_1236);
nand U5095 (N_5095,N_303,N_1732);
and U5096 (N_5096,N_919,N_1626);
xor U5097 (N_5097,N_2933,N_386);
and U5098 (N_5098,N_1765,N_2722);
and U5099 (N_5099,N_2277,N_919);
and U5100 (N_5100,N_357,N_753);
and U5101 (N_5101,N_2720,N_2074);
nand U5102 (N_5102,N_173,N_1666);
nand U5103 (N_5103,N_2111,N_1436);
xnor U5104 (N_5104,N_2137,N_2209);
nand U5105 (N_5105,N_499,N_2514);
xnor U5106 (N_5106,N_51,N_1637);
nor U5107 (N_5107,N_603,N_2870);
nand U5108 (N_5108,N_527,N_2835);
nand U5109 (N_5109,N_794,N_2536);
nor U5110 (N_5110,N_883,N_1359);
or U5111 (N_5111,N_2813,N_3105);
or U5112 (N_5112,N_721,N_2816);
xnor U5113 (N_5113,N_239,N_1282);
xor U5114 (N_5114,N_1426,N_936);
or U5115 (N_5115,N_1722,N_261);
nand U5116 (N_5116,N_2468,N_1735);
nand U5117 (N_5117,N_127,N_1038);
or U5118 (N_5118,N_915,N_361);
xor U5119 (N_5119,N_63,N_1891);
nor U5120 (N_5120,N_2116,N_2002);
nor U5121 (N_5121,N_16,N_2910);
xor U5122 (N_5122,N_2635,N_3025);
xnor U5123 (N_5123,N_2838,N_1610);
xnor U5124 (N_5124,N_2261,N_2156);
xor U5125 (N_5125,N_1273,N_2884);
and U5126 (N_5126,N_106,N_1907);
nor U5127 (N_5127,N_983,N_1925);
nor U5128 (N_5128,N_1836,N_782);
nor U5129 (N_5129,N_3114,N_868);
nor U5130 (N_5130,N_1038,N_1222);
nor U5131 (N_5131,N_1412,N_1091);
nor U5132 (N_5132,N_1958,N_1063);
and U5133 (N_5133,N_965,N_335);
and U5134 (N_5134,N_1089,N_1210);
nand U5135 (N_5135,N_1410,N_215);
and U5136 (N_5136,N_1897,N_1359);
xor U5137 (N_5137,N_852,N_1357);
and U5138 (N_5138,N_2134,N_2653);
nand U5139 (N_5139,N_1280,N_2811);
xor U5140 (N_5140,N_773,N_841);
or U5141 (N_5141,N_2445,N_1263);
or U5142 (N_5142,N_1281,N_2492);
nor U5143 (N_5143,N_2021,N_623);
nor U5144 (N_5144,N_2816,N_1244);
nor U5145 (N_5145,N_2514,N_1435);
or U5146 (N_5146,N_481,N_1926);
and U5147 (N_5147,N_2343,N_2905);
and U5148 (N_5148,N_1082,N_1176);
xnor U5149 (N_5149,N_2272,N_1515);
and U5150 (N_5150,N_2086,N_255);
or U5151 (N_5151,N_2042,N_2435);
nor U5152 (N_5152,N_2823,N_2473);
nand U5153 (N_5153,N_1116,N_2065);
nor U5154 (N_5154,N_2758,N_823);
and U5155 (N_5155,N_2311,N_2787);
and U5156 (N_5156,N_2089,N_1649);
nor U5157 (N_5157,N_2600,N_2551);
nor U5158 (N_5158,N_648,N_2209);
and U5159 (N_5159,N_469,N_1919);
nor U5160 (N_5160,N_2560,N_1246);
xor U5161 (N_5161,N_2868,N_1497);
xor U5162 (N_5162,N_930,N_2595);
or U5163 (N_5163,N_410,N_1931);
nor U5164 (N_5164,N_2031,N_1086);
nand U5165 (N_5165,N_545,N_968);
nor U5166 (N_5166,N_97,N_438);
xor U5167 (N_5167,N_1807,N_2097);
xor U5168 (N_5168,N_826,N_1518);
or U5169 (N_5169,N_2912,N_2462);
or U5170 (N_5170,N_2527,N_622);
or U5171 (N_5171,N_2843,N_66);
or U5172 (N_5172,N_687,N_359);
or U5173 (N_5173,N_2803,N_1513);
or U5174 (N_5174,N_525,N_157);
nand U5175 (N_5175,N_1404,N_1968);
xnor U5176 (N_5176,N_1476,N_569);
and U5177 (N_5177,N_1306,N_2874);
nand U5178 (N_5178,N_3044,N_472);
and U5179 (N_5179,N_1613,N_431);
xor U5180 (N_5180,N_2194,N_1816);
and U5181 (N_5181,N_2869,N_1215);
nand U5182 (N_5182,N_1510,N_2539);
or U5183 (N_5183,N_2817,N_1749);
nor U5184 (N_5184,N_1854,N_2514);
or U5185 (N_5185,N_2821,N_1267);
and U5186 (N_5186,N_1571,N_868);
xnor U5187 (N_5187,N_2483,N_292);
or U5188 (N_5188,N_1782,N_3019);
or U5189 (N_5189,N_2528,N_1461);
nand U5190 (N_5190,N_966,N_714);
and U5191 (N_5191,N_1934,N_1865);
xnor U5192 (N_5192,N_199,N_2193);
xor U5193 (N_5193,N_1563,N_2398);
and U5194 (N_5194,N_986,N_563);
nand U5195 (N_5195,N_1537,N_1457);
and U5196 (N_5196,N_1892,N_3008);
nand U5197 (N_5197,N_2083,N_1305);
nor U5198 (N_5198,N_2503,N_2643);
or U5199 (N_5199,N_2454,N_815);
xnor U5200 (N_5200,N_82,N_1697);
xnor U5201 (N_5201,N_739,N_1793);
and U5202 (N_5202,N_347,N_2693);
nand U5203 (N_5203,N_247,N_1983);
or U5204 (N_5204,N_14,N_2707);
and U5205 (N_5205,N_513,N_1605);
or U5206 (N_5206,N_2664,N_1069);
xnor U5207 (N_5207,N_729,N_738);
xor U5208 (N_5208,N_927,N_1535);
nand U5209 (N_5209,N_956,N_391);
xor U5210 (N_5210,N_2716,N_1591);
nand U5211 (N_5211,N_2346,N_2128);
xor U5212 (N_5212,N_1101,N_1985);
and U5213 (N_5213,N_2225,N_1299);
xnor U5214 (N_5214,N_1114,N_2980);
and U5215 (N_5215,N_79,N_18);
or U5216 (N_5216,N_1396,N_1083);
xor U5217 (N_5217,N_3069,N_2614);
xor U5218 (N_5218,N_1775,N_2592);
xnor U5219 (N_5219,N_996,N_321);
nor U5220 (N_5220,N_917,N_1489);
and U5221 (N_5221,N_3118,N_1854);
and U5222 (N_5222,N_422,N_1217);
xor U5223 (N_5223,N_852,N_1793);
or U5224 (N_5224,N_1807,N_2114);
nand U5225 (N_5225,N_2489,N_1245);
and U5226 (N_5226,N_2756,N_1560);
and U5227 (N_5227,N_1909,N_1535);
and U5228 (N_5228,N_1466,N_1833);
or U5229 (N_5229,N_2204,N_111);
nor U5230 (N_5230,N_1402,N_288);
xor U5231 (N_5231,N_337,N_3051);
or U5232 (N_5232,N_1611,N_2063);
and U5233 (N_5233,N_30,N_1525);
xnor U5234 (N_5234,N_1699,N_1235);
nand U5235 (N_5235,N_1601,N_1718);
xor U5236 (N_5236,N_24,N_56);
or U5237 (N_5237,N_2564,N_829);
or U5238 (N_5238,N_1813,N_2570);
or U5239 (N_5239,N_767,N_2725);
or U5240 (N_5240,N_1334,N_286);
or U5241 (N_5241,N_515,N_2133);
and U5242 (N_5242,N_362,N_1975);
nor U5243 (N_5243,N_2838,N_1882);
xor U5244 (N_5244,N_981,N_2572);
xnor U5245 (N_5245,N_110,N_1387);
nor U5246 (N_5246,N_1854,N_2202);
nor U5247 (N_5247,N_1808,N_671);
nor U5248 (N_5248,N_1655,N_916);
nor U5249 (N_5249,N_2181,N_799);
nand U5250 (N_5250,N_12,N_2586);
nor U5251 (N_5251,N_3096,N_381);
and U5252 (N_5252,N_2299,N_1314);
nand U5253 (N_5253,N_196,N_2502);
or U5254 (N_5254,N_2820,N_290);
nand U5255 (N_5255,N_266,N_1612);
nor U5256 (N_5256,N_1395,N_932);
and U5257 (N_5257,N_1759,N_2096);
nand U5258 (N_5258,N_2240,N_2493);
xnor U5259 (N_5259,N_1512,N_2235);
nand U5260 (N_5260,N_501,N_2047);
nor U5261 (N_5261,N_1138,N_2008);
xnor U5262 (N_5262,N_963,N_875);
nand U5263 (N_5263,N_1447,N_726);
nand U5264 (N_5264,N_1942,N_2796);
and U5265 (N_5265,N_2,N_6);
nor U5266 (N_5266,N_2747,N_189);
xnor U5267 (N_5267,N_2598,N_1852);
or U5268 (N_5268,N_3115,N_184);
xor U5269 (N_5269,N_1321,N_2421);
or U5270 (N_5270,N_839,N_2723);
and U5271 (N_5271,N_677,N_1775);
nand U5272 (N_5272,N_837,N_1031);
xnor U5273 (N_5273,N_1979,N_2834);
nand U5274 (N_5274,N_2664,N_2848);
or U5275 (N_5275,N_84,N_2345);
nand U5276 (N_5276,N_33,N_204);
or U5277 (N_5277,N_2084,N_1348);
and U5278 (N_5278,N_1845,N_1764);
nor U5279 (N_5279,N_1291,N_2302);
nand U5280 (N_5280,N_983,N_827);
and U5281 (N_5281,N_1510,N_1310);
and U5282 (N_5282,N_717,N_883);
nor U5283 (N_5283,N_2679,N_1905);
and U5284 (N_5284,N_2491,N_1605);
nand U5285 (N_5285,N_3111,N_3112);
xor U5286 (N_5286,N_3123,N_1432);
or U5287 (N_5287,N_1534,N_453);
xor U5288 (N_5288,N_2723,N_375);
or U5289 (N_5289,N_1049,N_2179);
nor U5290 (N_5290,N_2035,N_1636);
nor U5291 (N_5291,N_691,N_1374);
nand U5292 (N_5292,N_776,N_2949);
or U5293 (N_5293,N_1743,N_1258);
nor U5294 (N_5294,N_2853,N_2849);
xnor U5295 (N_5295,N_2888,N_2817);
nor U5296 (N_5296,N_3035,N_990);
or U5297 (N_5297,N_1722,N_384);
and U5298 (N_5298,N_2606,N_2383);
and U5299 (N_5299,N_1537,N_226);
nor U5300 (N_5300,N_695,N_277);
or U5301 (N_5301,N_916,N_741);
xnor U5302 (N_5302,N_2872,N_1237);
and U5303 (N_5303,N_2886,N_1169);
nand U5304 (N_5304,N_196,N_3078);
xor U5305 (N_5305,N_3084,N_3088);
nor U5306 (N_5306,N_1762,N_1943);
nand U5307 (N_5307,N_261,N_2257);
and U5308 (N_5308,N_1653,N_1257);
xor U5309 (N_5309,N_592,N_1114);
xor U5310 (N_5310,N_91,N_1344);
nor U5311 (N_5311,N_108,N_465);
nor U5312 (N_5312,N_1959,N_2724);
nand U5313 (N_5313,N_2374,N_39);
xor U5314 (N_5314,N_2400,N_114);
nor U5315 (N_5315,N_132,N_1377);
and U5316 (N_5316,N_1739,N_419);
and U5317 (N_5317,N_496,N_176);
or U5318 (N_5318,N_3060,N_874);
and U5319 (N_5319,N_977,N_2877);
and U5320 (N_5320,N_1188,N_1333);
and U5321 (N_5321,N_2582,N_1726);
xor U5322 (N_5322,N_425,N_861);
or U5323 (N_5323,N_1146,N_1060);
nor U5324 (N_5324,N_2739,N_1700);
nor U5325 (N_5325,N_133,N_376);
nor U5326 (N_5326,N_1982,N_612);
or U5327 (N_5327,N_1,N_431);
xnor U5328 (N_5328,N_451,N_2214);
xor U5329 (N_5329,N_2949,N_810);
nand U5330 (N_5330,N_1314,N_344);
and U5331 (N_5331,N_1062,N_2028);
nor U5332 (N_5332,N_2320,N_115);
nor U5333 (N_5333,N_1434,N_796);
xor U5334 (N_5334,N_2986,N_1510);
or U5335 (N_5335,N_1338,N_2669);
or U5336 (N_5336,N_291,N_2224);
nor U5337 (N_5337,N_1536,N_2999);
or U5338 (N_5338,N_1074,N_1050);
xnor U5339 (N_5339,N_1064,N_2666);
nand U5340 (N_5340,N_1283,N_1039);
or U5341 (N_5341,N_2245,N_1452);
nor U5342 (N_5342,N_268,N_256);
and U5343 (N_5343,N_2278,N_948);
or U5344 (N_5344,N_682,N_1279);
nor U5345 (N_5345,N_156,N_2137);
xnor U5346 (N_5346,N_2839,N_263);
or U5347 (N_5347,N_2114,N_3040);
xnor U5348 (N_5348,N_1688,N_1693);
xnor U5349 (N_5349,N_2423,N_2282);
nor U5350 (N_5350,N_2326,N_2697);
xor U5351 (N_5351,N_1507,N_1027);
and U5352 (N_5352,N_1037,N_653);
nor U5353 (N_5353,N_2205,N_1704);
or U5354 (N_5354,N_914,N_1105);
nor U5355 (N_5355,N_2738,N_1004);
nor U5356 (N_5356,N_1533,N_1686);
nand U5357 (N_5357,N_165,N_2314);
or U5358 (N_5358,N_1408,N_2367);
nand U5359 (N_5359,N_1878,N_875);
nor U5360 (N_5360,N_2905,N_1978);
nor U5361 (N_5361,N_2526,N_2607);
nor U5362 (N_5362,N_1914,N_808);
xnor U5363 (N_5363,N_3107,N_1659);
nand U5364 (N_5364,N_1476,N_1202);
nand U5365 (N_5365,N_2682,N_1162);
xnor U5366 (N_5366,N_2514,N_2557);
nor U5367 (N_5367,N_22,N_927);
nor U5368 (N_5368,N_222,N_1468);
nor U5369 (N_5369,N_1074,N_16);
xnor U5370 (N_5370,N_731,N_2372);
xor U5371 (N_5371,N_20,N_2270);
and U5372 (N_5372,N_59,N_2984);
and U5373 (N_5373,N_44,N_855);
nand U5374 (N_5374,N_2194,N_2564);
nor U5375 (N_5375,N_5,N_2551);
and U5376 (N_5376,N_2942,N_1103);
xor U5377 (N_5377,N_917,N_152);
xor U5378 (N_5378,N_1580,N_314);
nand U5379 (N_5379,N_2230,N_935);
or U5380 (N_5380,N_260,N_2922);
nand U5381 (N_5381,N_1982,N_1433);
or U5382 (N_5382,N_1983,N_1311);
nand U5383 (N_5383,N_2436,N_2951);
and U5384 (N_5384,N_2606,N_724);
and U5385 (N_5385,N_2553,N_806);
nand U5386 (N_5386,N_2039,N_2976);
or U5387 (N_5387,N_1830,N_2234);
nand U5388 (N_5388,N_20,N_1486);
and U5389 (N_5389,N_1758,N_2429);
or U5390 (N_5390,N_140,N_1093);
nor U5391 (N_5391,N_2742,N_1725);
xor U5392 (N_5392,N_2432,N_804);
or U5393 (N_5393,N_1112,N_862);
nand U5394 (N_5394,N_1078,N_436);
nand U5395 (N_5395,N_1662,N_2254);
or U5396 (N_5396,N_3013,N_483);
or U5397 (N_5397,N_837,N_1949);
and U5398 (N_5398,N_2347,N_845);
and U5399 (N_5399,N_2688,N_1288);
nand U5400 (N_5400,N_2118,N_668);
nand U5401 (N_5401,N_1646,N_615);
nand U5402 (N_5402,N_1887,N_395);
nor U5403 (N_5403,N_2953,N_227);
or U5404 (N_5404,N_705,N_2484);
nand U5405 (N_5405,N_95,N_185);
and U5406 (N_5406,N_2725,N_2945);
nand U5407 (N_5407,N_1918,N_2273);
nor U5408 (N_5408,N_2534,N_1476);
nand U5409 (N_5409,N_2775,N_534);
and U5410 (N_5410,N_945,N_2345);
nand U5411 (N_5411,N_79,N_1858);
xnor U5412 (N_5412,N_50,N_2176);
and U5413 (N_5413,N_195,N_714);
nand U5414 (N_5414,N_1015,N_520);
or U5415 (N_5415,N_987,N_2545);
or U5416 (N_5416,N_1404,N_16);
and U5417 (N_5417,N_2312,N_163);
and U5418 (N_5418,N_1132,N_1241);
nor U5419 (N_5419,N_2584,N_1124);
and U5420 (N_5420,N_1221,N_2855);
xnor U5421 (N_5421,N_1369,N_1762);
nor U5422 (N_5422,N_407,N_2541);
nor U5423 (N_5423,N_2216,N_1862);
or U5424 (N_5424,N_2173,N_480);
xor U5425 (N_5425,N_2603,N_2414);
nor U5426 (N_5426,N_668,N_1890);
or U5427 (N_5427,N_2170,N_1736);
or U5428 (N_5428,N_2479,N_611);
or U5429 (N_5429,N_440,N_2549);
nand U5430 (N_5430,N_2201,N_3107);
or U5431 (N_5431,N_2282,N_32);
xor U5432 (N_5432,N_2237,N_3017);
and U5433 (N_5433,N_265,N_794);
and U5434 (N_5434,N_2900,N_1259);
xor U5435 (N_5435,N_1919,N_1344);
or U5436 (N_5436,N_2243,N_1166);
or U5437 (N_5437,N_2719,N_2833);
nor U5438 (N_5438,N_2754,N_932);
nand U5439 (N_5439,N_2521,N_2903);
or U5440 (N_5440,N_1282,N_2305);
or U5441 (N_5441,N_1302,N_2373);
nor U5442 (N_5442,N_546,N_2654);
nor U5443 (N_5443,N_2551,N_832);
nor U5444 (N_5444,N_267,N_771);
nand U5445 (N_5445,N_1016,N_1301);
and U5446 (N_5446,N_2348,N_638);
nand U5447 (N_5447,N_2268,N_3063);
and U5448 (N_5448,N_1745,N_1483);
or U5449 (N_5449,N_417,N_607);
nor U5450 (N_5450,N_194,N_2382);
and U5451 (N_5451,N_699,N_1159);
or U5452 (N_5452,N_1243,N_346);
nor U5453 (N_5453,N_2771,N_2606);
nand U5454 (N_5454,N_2126,N_1796);
nor U5455 (N_5455,N_1063,N_1014);
nand U5456 (N_5456,N_2193,N_869);
nor U5457 (N_5457,N_801,N_2615);
xnor U5458 (N_5458,N_1015,N_3038);
nor U5459 (N_5459,N_2931,N_1183);
and U5460 (N_5460,N_2435,N_2132);
xor U5461 (N_5461,N_1650,N_1615);
xor U5462 (N_5462,N_2869,N_784);
and U5463 (N_5463,N_2554,N_2792);
xor U5464 (N_5464,N_606,N_973);
or U5465 (N_5465,N_360,N_981);
and U5466 (N_5466,N_994,N_1418);
nor U5467 (N_5467,N_1067,N_1307);
and U5468 (N_5468,N_1791,N_249);
and U5469 (N_5469,N_508,N_2966);
or U5470 (N_5470,N_2056,N_249);
nand U5471 (N_5471,N_1040,N_2609);
or U5472 (N_5472,N_1305,N_2145);
nor U5473 (N_5473,N_1244,N_2862);
xnor U5474 (N_5474,N_2818,N_714);
or U5475 (N_5475,N_2051,N_1482);
nor U5476 (N_5476,N_2077,N_453);
nor U5477 (N_5477,N_3103,N_1111);
nor U5478 (N_5478,N_1488,N_1805);
nor U5479 (N_5479,N_2012,N_29);
or U5480 (N_5480,N_1669,N_2476);
or U5481 (N_5481,N_173,N_494);
nor U5482 (N_5482,N_2097,N_2745);
and U5483 (N_5483,N_2600,N_824);
and U5484 (N_5484,N_2279,N_94);
or U5485 (N_5485,N_2663,N_2270);
and U5486 (N_5486,N_2024,N_2979);
or U5487 (N_5487,N_2023,N_1683);
and U5488 (N_5488,N_54,N_760);
and U5489 (N_5489,N_1482,N_2835);
nand U5490 (N_5490,N_1852,N_2455);
or U5491 (N_5491,N_1451,N_2525);
nor U5492 (N_5492,N_1515,N_470);
xor U5493 (N_5493,N_2173,N_119);
and U5494 (N_5494,N_2623,N_2873);
and U5495 (N_5495,N_1397,N_2946);
and U5496 (N_5496,N_3063,N_153);
nand U5497 (N_5497,N_2593,N_1081);
xnor U5498 (N_5498,N_474,N_1005);
or U5499 (N_5499,N_1362,N_1612);
xnor U5500 (N_5500,N_495,N_1730);
or U5501 (N_5501,N_2671,N_2173);
and U5502 (N_5502,N_136,N_1746);
and U5503 (N_5503,N_1526,N_2987);
and U5504 (N_5504,N_1143,N_3015);
and U5505 (N_5505,N_2234,N_1036);
xnor U5506 (N_5506,N_2182,N_827);
xor U5507 (N_5507,N_1019,N_2788);
or U5508 (N_5508,N_1517,N_2751);
or U5509 (N_5509,N_2290,N_2194);
nand U5510 (N_5510,N_30,N_1818);
xnor U5511 (N_5511,N_995,N_899);
xnor U5512 (N_5512,N_963,N_288);
or U5513 (N_5513,N_1209,N_2269);
nor U5514 (N_5514,N_2001,N_1723);
or U5515 (N_5515,N_2616,N_1503);
or U5516 (N_5516,N_568,N_1975);
nand U5517 (N_5517,N_2473,N_1815);
xor U5518 (N_5518,N_750,N_2668);
and U5519 (N_5519,N_2851,N_912);
or U5520 (N_5520,N_643,N_1600);
nor U5521 (N_5521,N_290,N_2629);
or U5522 (N_5522,N_437,N_934);
and U5523 (N_5523,N_2108,N_1389);
or U5524 (N_5524,N_7,N_1671);
and U5525 (N_5525,N_957,N_2020);
nand U5526 (N_5526,N_97,N_1890);
and U5527 (N_5527,N_5,N_2921);
xor U5528 (N_5528,N_2072,N_1893);
and U5529 (N_5529,N_2220,N_1235);
xnor U5530 (N_5530,N_340,N_2138);
or U5531 (N_5531,N_1246,N_1976);
xor U5532 (N_5532,N_2288,N_733);
and U5533 (N_5533,N_1879,N_3004);
xnor U5534 (N_5534,N_1614,N_542);
nand U5535 (N_5535,N_2555,N_402);
xnor U5536 (N_5536,N_2743,N_113);
xnor U5537 (N_5537,N_929,N_2150);
or U5538 (N_5538,N_430,N_268);
nor U5539 (N_5539,N_1979,N_1859);
or U5540 (N_5540,N_2689,N_648);
or U5541 (N_5541,N_1243,N_1918);
or U5542 (N_5542,N_727,N_2063);
nor U5543 (N_5543,N_1516,N_2197);
or U5544 (N_5544,N_3076,N_684);
xnor U5545 (N_5545,N_1726,N_2631);
and U5546 (N_5546,N_3100,N_2265);
nor U5547 (N_5547,N_260,N_1580);
nand U5548 (N_5548,N_746,N_91);
xnor U5549 (N_5549,N_2341,N_1611);
nor U5550 (N_5550,N_1417,N_1448);
and U5551 (N_5551,N_1541,N_1778);
nand U5552 (N_5552,N_3085,N_2875);
xnor U5553 (N_5553,N_2261,N_1082);
and U5554 (N_5554,N_1513,N_2660);
nor U5555 (N_5555,N_69,N_181);
xnor U5556 (N_5556,N_954,N_2419);
xor U5557 (N_5557,N_1585,N_1189);
nor U5558 (N_5558,N_1714,N_2922);
nand U5559 (N_5559,N_2418,N_947);
nand U5560 (N_5560,N_3066,N_3061);
nor U5561 (N_5561,N_2396,N_1533);
and U5562 (N_5562,N_200,N_2833);
nor U5563 (N_5563,N_2144,N_2983);
or U5564 (N_5564,N_789,N_2451);
xnor U5565 (N_5565,N_280,N_1437);
and U5566 (N_5566,N_2687,N_515);
xor U5567 (N_5567,N_728,N_2916);
xor U5568 (N_5568,N_1478,N_1577);
nor U5569 (N_5569,N_2150,N_2615);
nor U5570 (N_5570,N_414,N_1547);
and U5571 (N_5571,N_3097,N_880);
nand U5572 (N_5572,N_308,N_877);
nand U5573 (N_5573,N_2763,N_2854);
nand U5574 (N_5574,N_2087,N_2312);
nand U5575 (N_5575,N_484,N_2101);
xnor U5576 (N_5576,N_666,N_842);
nand U5577 (N_5577,N_1909,N_2294);
xnor U5578 (N_5578,N_435,N_2382);
xnor U5579 (N_5579,N_2883,N_2147);
nor U5580 (N_5580,N_1945,N_2725);
and U5581 (N_5581,N_12,N_966);
nor U5582 (N_5582,N_442,N_1277);
or U5583 (N_5583,N_2244,N_1437);
and U5584 (N_5584,N_2784,N_2078);
nor U5585 (N_5585,N_346,N_760);
or U5586 (N_5586,N_1917,N_503);
and U5587 (N_5587,N_2093,N_615);
xor U5588 (N_5588,N_1440,N_2782);
nand U5589 (N_5589,N_2953,N_1284);
xnor U5590 (N_5590,N_1012,N_846);
and U5591 (N_5591,N_1690,N_2751);
nor U5592 (N_5592,N_1324,N_482);
or U5593 (N_5593,N_2908,N_961);
nor U5594 (N_5594,N_285,N_84);
or U5595 (N_5595,N_2854,N_825);
nand U5596 (N_5596,N_2777,N_1746);
xor U5597 (N_5597,N_668,N_782);
and U5598 (N_5598,N_181,N_2249);
nor U5599 (N_5599,N_2418,N_2513);
and U5600 (N_5600,N_657,N_75);
nand U5601 (N_5601,N_754,N_637);
nor U5602 (N_5602,N_544,N_662);
nor U5603 (N_5603,N_1193,N_282);
nand U5604 (N_5604,N_2381,N_880);
nand U5605 (N_5605,N_2568,N_1847);
or U5606 (N_5606,N_27,N_1446);
nor U5607 (N_5607,N_2919,N_2050);
or U5608 (N_5608,N_1655,N_1600);
or U5609 (N_5609,N_2664,N_40);
or U5610 (N_5610,N_1636,N_2165);
nor U5611 (N_5611,N_2715,N_600);
or U5612 (N_5612,N_2599,N_1098);
nand U5613 (N_5613,N_878,N_1487);
nor U5614 (N_5614,N_1820,N_1285);
nor U5615 (N_5615,N_1014,N_2020);
nor U5616 (N_5616,N_2166,N_1288);
and U5617 (N_5617,N_2651,N_2184);
or U5618 (N_5618,N_2936,N_601);
nor U5619 (N_5619,N_445,N_2229);
and U5620 (N_5620,N_341,N_2470);
or U5621 (N_5621,N_205,N_2672);
nand U5622 (N_5622,N_695,N_1693);
and U5623 (N_5623,N_1847,N_1422);
or U5624 (N_5624,N_899,N_1225);
nand U5625 (N_5625,N_762,N_1913);
nor U5626 (N_5626,N_382,N_162);
or U5627 (N_5627,N_1316,N_445);
nand U5628 (N_5628,N_3047,N_1071);
nor U5629 (N_5629,N_2960,N_1237);
or U5630 (N_5630,N_3080,N_446);
or U5631 (N_5631,N_276,N_1651);
nand U5632 (N_5632,N_210,N_1407);
and U5633 (N_5633,N_1770,N_359);
nor U5634 (N_5634,N_937,N_2746);
xor U5635 (N_5635,N_1714,N_648);
nor U5636 (N_5636,N_1420,N_1540);
or U5637 (N_5637,N_151,N_1996);
nand U5638 (N_5638,N_580,N_2878);
nor U5639 (N_5639,N_599,N_618);
nor U5640 (N_5640,N_2617,N_694);
nor U5641 (N_5641,N_927,N_1819);
nor U5642 (N_5642,N_1665,N_1521);
nor U5643 (N_5643,N_2211,N_2582);
xor U5644 (N_5644,N_2023,N_1323);
nand U5645 (N_5645,N_145,N_1264);
and U5646 (N_5646,N_570,N_2117);
and U5647 (N_5647,N_733,N_575);
nor U5648 (N_5648,N_2854,N_2276);
nor U5649 (N_5649,N_844,N_1123);
nor U5650 (N_5650,N_1506,N_543);
and U5651 (N_5651,N_1672,N_2319);
and U5652 (N_5652,N_806,N_2523);
nand U5653 (N_5653,N_96,N_2924);
xnor U5654 (N_5654,N_1284,N_386);
nand U5655 (N_5655,N_818,N_3077);
or U5656 (N_5656,N_2685,N_136);
nand U5657 (N_5657,N_1117,N_650);
nand U5658 (N_5658,N_842,N_1341);
nor U5659 (N_5659,N_465,N_682);
xnor U5660 (N_5660,N_287,N_141);
and U5661 (N_5661,N_2618,N_1059);
or U5662 (N_5662,N_753,N_789);
nor U5663 (N_5663,N_2248,N_1455);
nor U5664 (N_5664,N_1618,N_2537);
and U5665 (N_5665,N_580,N_865);
or U5666 (N_5666,N_2735,N_1302);
nor U5667 (N_5667,N_1332,N_1799);
xnor U5668 (N_5668,N_1338,N_991);
or U5669 (N_5669,N_1346,N_521);
and U5670 (N_5670,N_2899,N_446);
and U5671 (N_5671,N_3085,N_2076);
nand U5672 (N_5672,N_2953,N_2281);
nand U5673 (N_5673,N_1595,N_2175);
xor U5674 (N_5674,N_3040,N_2822);
xnor U5675 (N_5675,N_5,N_2648);
nor U5676 (N_5676,N_401,N_792);
nand U5677 (N_5677,N_420,N_540);
or U5678 (N_5678,N_994,N_535);
and U5679 (N_5679,N_3042,N_428);
or U5680 (N_5680,N_2564,N_625);
nand U5681 (N_5681,N_2231,N_2107);
xnor U5682 (N_5682,N_2425,N_2632);
nand U5683 (N_5683,N_3,N_2031);
nor U5684 (N_5684,N_1274,N_639);
nor U5685 (N_5685,N_2199,N_544);
xor U5686 (N_5686,N_504,N_2292);
or U5687 (N_5687,N_791,N_457);
and U5688 (N_5688,N_1664,N_1637);
or U5689 (N_5689,N_3123,N_2006);
xor U5690 (N_5690,N_559,N_1816);
nor U5691 (N_5691,N_631,N_397);
xor U5692 (N_5692,N_621,N_2022);
xnor U5693 (N_5693,N_1862,N_2787);
nand U5694 (N_5694,N_1903,N_1179);
and U5695 (N_5695,N_2725,N_3038);
or U5696 (N_5696,N_2125,N_973);
nor U5697 (N_5697,N_1370,N_168);
and U5698 (N_5698,N_2560,N_185);
xor U5699 (N_5699,N_1679,N_396);
xor U5700 (N_5700,N_1193,N_3004);
nor U5701 (N_5701,N_1950,N_2298);
or U5702 (N_5702,N_1542,N_603);
nor U5703 (N_5703,N_1273,N_2714);
nor U5704 (N_5704,N_1702,N_2458);
nand U5705 (N_5705,N_1019,N_1463);
or U5706 (N_5706,N_729,N_1122);
xnor U5707 (N_5707,N_2948,N_1919);
xor U5708 (N_5708,N_2246,N_1529);
xnor U5709 (N_5709,N_1202,N_2566);
nor U5710 (N_5710,N_414,N_1343);
or U5711 (N_5711,N_542,N_2166);
or U5712 (N_5712,N_1645,N_72);
xnor U5713 (N_5713,N_1524,N_2684);
nand U5714 (N_5714,N_2871,N_45);
or U5715 (N_5715,N_2274,N_305);
nor U5716 (N_5716,N_1527,N_2535);
and U5717 (N_5717,N_1679,N_2709);
or U5718 (N_5718,N_2166,N_1916);
or U5719 (N_5719,N_2689,N_494);
nand U5720 (N_5720,N_1095,N_844);
xor U5721 (N_5721,N_1585,N_2092);
nor U5722 (N_5722,N_1180,N_1568);
xor U5723 (N_5723,N_1210,N_2830);
nor U5724 (N_5724,N_1521,N_3095);
xnor U5725 (N_5725,N_2982,N_2793);
xnor U5726 (N_5726,N_2139,N_2201);
and U5727 (N_5727,N_7,N_1377);
and U5728 (N_5728,N_2747,N_1850);
xor U5729 (N_5729,N_2523,N_1468);
and U5730 (N_5730,N_278,N_2688);
nand U5731 (N_5731,N_264,N_607);
or U5732 (N_5732,N_418,N_314);
nand U5733 (N_5733,N_3000,N_2375);
nand U5734 (N_5734,N_2444,N_2757);
xnor U5735 (N_5735,N_1710,N_205);
xor U5736 (N_5736,N_477,N_2657);
nand U5737 (N_5737,N_1224,N_522);
nor U5738 (N_5738,N_2501,N_2781);
nor U5739 (N_5739,N_1010,N_1148);
xnor U5740 (N_5740,N_942,N_1049);
or U5741 (N_5741,N_3047,N_457);
nand U5742 (N_5742,N_2875,N_2545);
or U5743 (N_5743,N_812,N_1368);
and U5744 (N_5744,N_2872,N_715);
and U5745 (N_5745,N_1871,N_2612);
and U5746 (N_5746,N_2850,N_359);
and U5747 (N_5747,N_926,N_1268);
or U5748 (N_5748,N_863,N_2574);
xnor U5749 (N_5749,N_3114,N_2296);
xor U5750 (N_5750,N_2766,N_186);
and U5751 (N_5751,N_1220,N_1992);
xor U5752 (N_5752,N_1470,N_358);
nor U5753 (N_5753,N_544,N_1);
nand U5754 (N_5754,N_1206,N_556);
or U5755 (N_5755,N_2093,N_901);
and U5756 (N_5756,N_2008,N_3106);
or U5757 (N_5757,N_547,N_16);
nor U5758 (N_5758,N_2916,N_720);
nor U5759 (N_5759,N_1171,N_982);
or U5760 (N_5760,N_2137,N_587);
nor U5761 (N_5761,N_3024,N_2015);
or U5762 (N_5762,N_1664,N_988);
xnor U5763 (N_5763,N_375,N_1827);
nor U5764 (N_5764,N_835,N_2639);
and U5765 (N_5765,N_1978,N_1929);
xnor U5766 (N_5766,N_2041,N_2637);
xor U5767 (N_5767,N_2473,N_1126);
and U5768 (N_5768,N_2310,N_2464);
and U5769 (N_5769,N_1321,N_1884);
and U5770 (N_5770,N_654,N_1884);
and U5771 (N_5771,N_2422,N_1119);
and U5772 (N_5772,N_331,N_1750);
nand U5773 (N_5773,N_660,N_2383);
or U5774 (N_5774,N_572,N_20);
nor U5775 (N_5775,N_2057,N_1255);
and U5776 (N_5776,N_1956,N_3090);
or U5777 (N_5777,N_878,N_2103);
nand U5778 (N_5778,N_102,N_1983);
nand U5779 (N_5779,N_1465,N_1297);
or U5780 (N_5780,N_474,N_1792);
xnor U5781 (N_5781,N_1876,N_972);
nand U5782 (N_5782,N_2116,N_1460);
nor U5783 (N_5783,N_1520,N_693);
xnor U5784 (N_5784,N_2143,N_1909);
nand U5785 (N_5785,N_2450,N_1224);
or U5786 (N_5786,N_3041,N_514);
nand U5787 (N_5787,N_2392,N_2048);
xnor U5788 (N_5788,N_2787,N_2099);
or U5789 (N_5789,N_975,N_1453);
xor U5790 (N_5790,N_114,N_1182);
nor U5791 (N_5791,N_520,N_1310);
nor U5792 (N_5792,N_1281,N_315);
xor U5793 (N_5793,N_2652,N_2032);
and U5794 (N_5794,N_1774,N_2848);
xor U5795 (N_5795,N_2407,N_2936);
nand U5796 (N_5796,N_763,N_907);
xor U5797 (N_5797,N_1737,N_1772);
and U5798 (N_5798,N_53,N_2768);
or U5799 (N_5799,N_1820,N_1764);
and U5800 (N_5800,N_2029,N_570);
nand U5801 (N_5801,N_268,N_2017);
xnor U5802 (N_5802,N_699,N_1820);
nand U5803 (N_5803,N_2679,N_1164);
xor U5804 (N_5804,N_1317,N_2345);
nor U5805 (N_5805,N_2309,N_67);
and U5806 (N_5806,N_456,N_2640);
and U5807 (N_5807,N_1149,N_1706);
nand U5808 (N_5808,N_1517,N_1379);
and U5809 (N_5809,N_1537,N_3096);
xor U5810 (N_5810,N_59,N_1837);
nand U5811 (N_5811,N_2219,N_1267);
nand U5812 (N_5812,N_2741,N_2109);
nand U5813 (N_5813,N_2757,N_2875);
and U5814 (N_5814,N_705,N_834);
xor U5815 (N_5815,N_952,N_133);
nand U5816 (N_5816,N_2628,N_756);
xor U5817 (N_5817,N_2457,N_3077);
xnor U5818 (N_5818,N_2157,N_1186);
or U5819 (N_5819,N_314,N_971);
and U5820 (N_5820,N_2124,N_2139);
nand U5821 (N_5821,N_1819,N_353);
xnor U5822 (N_5822,N_216,N_762);
nand U5823 (N_5823,N_982,N_2787);
xor U5824 (N_5824,N_1559,N_3021);
nor U5825 (N_5825,N_2691,N_105);
nor U5826 (N_5826,N_1672,N_2268);
nor U5827 (N_5827,N_933,N_2489);
xnor U5828 (N_5828,N_527,N_699);
and U5829 (N_5829,N_2653,N_2422);
or U5830 (N_5830,N_162,N_346);
xnor U5831 (N_5831,N_595,N_46);
or U5832 (N_5832,N_2075,N_860);
or U5833 (N_5833,N_267,N_970);
nor U5834 (N_5834,N_2677,N_1778);
and U5835 (N_5835,N_3100,N_1287);
nand U5836 (N_5836,N_2018,N_569);
nand U5837 (N_5837,N_3111,N_1004);
xor U5838 (N_5838,N_2532,N_2697);
xnor U5839 (N_5839,N_391,N_2008);
xnor U5840 (N_5840,N_525,N_1016);
nor U5841 (N_5841,N_1042,N_1215);
xnor U5842 (N_5842,N_1321,N_963);
or U5843 (N_5843,N_860,N_677);
nor U5844 (N_5844,N_852,N_778);
or U5845 (N_5845,N_807,N_228);
or U5846 (N_5846,N_2486,N_3013);
nor U5847 (N_5847,N_1237,N_1152);
or U5848 (N_5848,N_201,N_1789);
and U5849 (N_5849,N_2470,N_2101);
nand U5850 (N_5850,N_545,N_2184);
and U5851 (N_5851,N_1611,N_842);
or U5852 (N_5852,N_392,N_1552);
or U5853 (N_5853,N_68,N_1962);
xnor U5854 (N_5854,N_2724,N_246);
nand U5855 (N_5855,N_2736,N_2315);
nand U5856 (N_5856,N_791,N_645);
and U5857 (N_5857,N_2709,N_799);
and U5858 (N_5858,N_2615,N_3120);
nand U5859 (N_5859,N_684,N_201);
xnor U5860 (N_5860,N_2295,N_1355);
and U5861 (N_5861,N_221,N_1081);
nor U5862 (N_5862,N_328,N_1557);
nand U5863 (N_5863,N_2679,N_1399);
xnor U5864 (N_5864,N_807,N_2779);
or U5865 (N_5865,N_2729,N_385);
nor U5866 (N_5866,N_422,N_1383);
xnor U5867 (N_5867,N_619,N_2643);
nor U5868 (N_5868,N_1002,N_2113);
nor U5869 (N_5869,N_3014,N_346);
and U5870 (N_5870,N_512,N_441);
xnor U5871 (N_5871,N_459,N_2368);
and U5872 (N_5872,N_621,N_942);
or U5873 (N_5873,N_807,N_1841);
nand U5874 (N_5874,N_2727,N_2853);
nor U5875 (N_5875,N_1977,N_2921);
or U5876 (N_5876,N_2191,N_890);
and U5877 (N_5877,N_1827,N_2056);
nor U5878 (N_5878,N_2134,N_1873);
or U5879 (N_5879,N_2080,N_1743);
nor U5880 (N_5880,N_3047,N_2340);
or U5881 (N_5881,N_1961,N_1590);
nand U5882 (N_5882,N_2822,N_2532);
nand U5883 (N_5883,N_383,N_2278);
xnor U5884 (N_5884,N_335,N_518);
and U5885 (N_5885,N_913,N_3112);
nand U5886 (N_5886,N_801,N_536);
nor U5887 (N_5887,N_159,N_2412);
nor U5888 (N_5888,N_2129,N_2617);
nand U5889 (N_5889,N_482,N_2344);
or U5890 (N_5890,N_2023,N_2605);
xor U5891 (N_5891,N_247,N_2925);
nor U5892 (N_5892,N_2838,N_1910);
xnor U5893 (N_5893,N_287,N_1571);
and U5894 (N_5894,N_1049,N_1769);
nand U5895 (N_5895,N_2169,N_2298);
xnor U5896 (N_5896,N_802,N_257);
and U5897 (N_5897,N_1324,N_1599);
nand U5898 (N_5898,N_2162,N_1923);
and U5899 (N_5899,N_979,N_773);
nand U5900 (N_5900,N_2635,N_2277);
and U5901 (N_5901,N_2689,N_1671);
nor U5902 (N_5902,N_2633,N_457);
nand U5903 (N_5903,N_3098,N_2895);
nand U5904 (N_5904,N_297,N_2562);
and U5905 (N_5905,N_2169,N_2526);
xor U5906 (N_5906,N_1313,N_2832);
xnor U5907 (N_5907,N_105,N_1163);
nand U5908 (N_5908,N_1685,N_1516);
and U5909 (N_5909,N_1790,N_248);
nor U5910 (N_5910,N_3005,N_2012);
or U5911 (N_5911,N_1638,N_510);
and U5912 (N_5912,N_1495,N_1839);
nor U5913 (N_5913,N_2641,N_1279);
and U5914 (N_5914,N_1901,N_2978);
or U5915 (N_5915,N_2337,N_1454);
or U5916 (N_5916,N_2293,N_2863);
xnor U5917 (N_5917,N_2290,N_1620);
nand U5918 (N_5918,N_216,N_2627);
nand U5919 (N_5919,N_2729,N_2554);
or U5920 (N_5920,N_663,N_189);
and U5921 (N_5921,N_74,N_364);
or U5922 (N_5922,N_1820,N_709);
nand U5923 (N_5923,N_3012,N_2918);
and U5924 (N_5924,N_1749,N_756);
nand U5925 (N_5925,N_1215,N_2873);
nand U5926 (N_5926,N_1420,N_945);
nor U5927 (N_5927,N_540,N_2966);
nand U5928 (N_5928,N_379,N_821);
nand U5929 (N_5929,N_1000,N_1888);
nand U5930 (N_5930,N_226,N_1564);
nand U5931 (N_5931,N_1021,N_1154);
xor U5932 (N_5932,N_554,N_1035);
and U5933 (N_5933,N_2294,N_148);
and U5934 (N_5934,N_2530,N_2336);
or U5935 (N_5935,N_1231,N_1312);
nor U5936 (N_5936,N_2163,N_2144);
xor U5937 (N_5937,N_1158,N_299);
nor U5938 (N_5938,N_2353,N_1349);
or U5939 (N_5939,N_1593,N_965);
or U5940 (N_5940,N_1402,N_2725);
or U5941 (N_5941,N_450,N_2546);
nor U5942 (N_5942,N_1284,N_2756);
and U5943 (N_5943,N_2590,N_207);
xor U5944 (N_5944,N_2417,N_161);
nand U5945 (N_5945,N_2745,N_1536);
or U5946 (N_5946,N_1698,N_1547);
nor U5947 (N_5947,N_2730,N_1150);
and U5948 (N_5948,N_1620,N_1104);
and U5949 (N_5949,N_1226,N_421);
nand U5950 (N_5950,N_2154,N_271);
and U5951 (N_5951,N_2618,N_2180);
nor U5952 (N_5952,N_366,N_1677);
xor U5953 (N_5953,N_816,N_1188);
nor U5954 (N_5954,N_1321,N_323);
xnor U5955 (N_5955,N_2399,N_2953);
or U5956 (N_5956,N_2411,N_1100);
or U5957 (N_5957,N_2337,N_2278);
nand U5958 (N_5958,N_2900,N_691);
nor U5959 (N_5959,N_2174,N_1645);
and U5960 (N_5960,N_2675,N_846);
nor U5961 (N_5961,N_1821,N_3102);
nand U5962 (N_5962,N_1027,N_2145);
or U5963 (N_5963,N_483,N_2450);
nor U5964 (N_5964,N_2284,N_1482);
nand U5965 (N_5965,N_2877,N_1815);
nor U5966 (N_5966,N_2673,N_1527);
xor U5967 (N_5967,N_1346,N_2444);
and U5968 (N_5968,N_1634,N_278);
nand U5969 (N_5969,N_1261,N_2130);
xnor U5970 (N_5970,N_1313,N_2269);
and U5971 (N_5971,N_1301,N_2275);
and U5972 (N_5972,N_203,N_1769);
and U5973 (N_5973,N_2411,N_1040);
or U5974 (N_5974,N_2409,N_1680);
xnor U5975 (N_5975,N_2375,N_3111);
xnor U5976 (N_5976,N_575,N_2066);
xnor U5977 (N_5977,N_288,N_2955);
nor U5978 (N_5978,N_360,N_1095);
xor U5979 (N_5979,N_743,N_2528);
nor U5980 (N_5980,N_5,N_542);
xor U5981 (N_5981,N_1738,N_2184);
nand U5982 (N_5982,N_1055,N_2115);
xor U5983 (N_5983,N_1765,N_677);
xnor U5984 (N_5984,N_1777,N_320);
and U5985 (N_5985,N_703,N_2704);
nor U5986 (N_5986,N_777,N_41);
nand U5987 (N_5987,N_2504,N_1312);
and U5988 (N_5988,N_762,N_2856);
nor U5989 (N_5989,N_1689,N_2043);
xnor U5990 (N_5990,N_826,N_403);
or U5991 (N_5991,N_690,N_2483);
or U5992 (N_5992,N_916,N_1151);
xnor U5993 (N_5993,N_1194,N_942);
or U5994 (N_5994,N_1907,N_2673);
xnor U5995 (N_5995,N_246,N_2101);
or U5996 (N_5996,N_2707,N_1780);
and U5997 (N_5997,N_688,N_2097);
or U5998 (N_5998,N_3054,N_185);
xor U5999 (N_5999,N_1663,N_1005);
nand U6000 (N_6000,N_24,N_2954);
xnor U6001 (N_6001,N_1333,N_139);
or U6002 (N_6002,N_1149,N_646);
nand U6003 (N_6003,N_2337,N_2141);
nor U6004 (N_6004,N_1265,N_2379);
and U6005 (N_6005,N_1950,N_1449);
nand U6006 (N_6006,N_2296,N_2396);
nor U6007 (N_6007,N_453,N_2918);
and U6008 (N_6008,N_2143,N_2845);
xnor U6009 (N_6009,N_1498,N_1671);
xor U6010 (N_6010,N_680,N_1316);
or U6011 (N_6011,N_2087,N_1174);
xnor U6012 (N_6012,N_2843,N_911);
xnor U6013 (N_6013,N_1275,N_2298);
xnor U6014 (N_6014,N_2508,N_1810);
xor U6015 (N_6015,N_1236,N_978);
and U6016 (N_6016,N_761,N_1183);
nand U6017 (N_6017,N_1313,N_2699);
or U6018 (N_6018,N_116,N_2422);
and U6019 (N_6019,N_1676,N_2389);
nand U6020 (N_6020,N_1233,N_2377);
xnor U6021 (N_6021,N_1370,N_2213);
nand U6022 (N_6022,N_1975,N_428);
and U6023 (N_6023,N_929,N_969);
nor U6024 (N_6024,N_1808,N_1999);
nor U6025 (N_6025,N_2582,N_1);
nor U6026 (N_6026,N_959,N_1389);
or U6027 (N_6027,N_665,N_2831);
xnor U6028 (N_6028,N_2307,N_1243);
or U6029 (N_6029,N_2936,N_1036);
nor U6030 (N_6030,N_722,N_1502);
xnor U6031 (N_6031,N_2641,N_2695);
and U6032 (N_6032,N_366,N_2246);
nand U6033 (N_6033,N_1235,N_1742);
or U6034 (N_6034,N_122,N_2920);
nor U6035 (N_6035,N_2642,N_2884);
and U6036 (N_6036,N_1914,N_1044);
xnor U6037 (N_6037,N_1969,N_166);
and U6038 (N_6038,N_2978,N_2507);
nand U6039 (N_6039,N_707,N_1072);
and U6040 (N_6040,N_2438,N_496);
nand U6041 (N_6041,N_1586,N_452);
xnor U6042 (N_6042,N_92,N_1923);
nor U6043 (N_6043,N_500,N_245);
nor U6044 (N_6044,N_2396,N_836);
and U6045 (N_6045,N_1758,N_1786);
and U6046 (N_6046,N_528,N_2951);
xor U6047 (N_6047,N_1844,N_2569);
and U6048 (N_6048,N_388,N_1061);
and U6049 (N_6049,N_618,N_2478);
xor U6050 (N_6050,N_1948,N_189);
and U6051 (N_6051,N_2074,N_1730);
and U6052 (N_6052,N_1096,N_2028);
xor U6053 (N_6053,N_1348,N_1775);
or U6054 (N_6054,N_3103,N_2470);
nor U6055 (N_6055,N_1846,N_2690);
xor U6056 (N_6056,N_2688,N_634);
nand U6057 (N_6057,N_1367,N_1709);
xnor U6058 (N_6058,N_614,N_1592);
nor U6059 (N_6059,N_1031,N_1386);
xnor U6060 (N_6060,N_1302,N_1231);
and U6061 (N_6061,N_250,N_48);
nor U6062 (N_6062,N_1865,N_2546);
nor U6063 (N_6063,N_1835,N_1563);
and U6064 (N_6064,N_2456,N_546);
nand U6065 (N_6065,N_3038,N_3114);
nor U6066 (N_6066,N_2707,N_2837);
or U6067 (N_6067,N_861,N_3084);
nand U6068 (N_6068,N_39,N_370);
xnor U6069 (N_6069,N_829,N_1368);
nand U6070 (N_6070,N_1500,N_2042);
nand U6071 (N_6071,N_586,N_1385);
and U6072 (N_6072,N_1859,N_2881);
nand U6073 (N_6073,N_478,N_2717);
nor U6074 (N_6074,N_3074,N_2236);
xnor U6075 (N_6075,N_1450,N_2621);
or U6076 (N_6076,N_1564,N_1125);
nor U6077 (N_6077,N_229,N_3003);
xor U6078 (N_6078,N_538,N_2466);
and U6079 (N_6079,N_1144,N_801);
or U6080 (N_6080,N_553,N_779);
and U6081 (N_6081,N_449,N_1636);
and U6082 (N_6082,N_2082,N_1405);
and U6083 (N_6083,N_2844,N_2098);
or U6084 (N_6084,N_2501,N_1756);
nor U6085 (N_6085,N_2138,N_723);
nand U6086 (N_6086,N_7,N_341);
and U6087 (N_6087,N_1799,N_2152);
nor U6088 (N_6088,N_2850,N_2841);
nor U6089 (N_6089,N_626,N_2453);
xor U6090 (N_6090,N_1430,N_223);
nand U6091 (N_6091,N_2617,N_2532);
xor U6092 (N_6092,N_1811,N_2519);
xor U6093 (N_6093,N_2699,N_2991);
or U6094 (N_6094,N_1588,N_649);
xor U6095 (N_6095,N_2371,N_1158);
nor U6096 (N_6096,N_782,N_3003);
xor U6097 (N_6097,N_25,N_2992);
nor U6098 (N_6098,N_815,N_384);
or U6099 (N_6099,N_395,N_2540);
or U6100 (N_6100,N_949,N_2347);
xnor U6101 (N_6101,N_1907,N_1012);
xor U6102 (N_6102,N_2742,N_156);
or U6103 (N_6103,N_939,N_3116);
or U6104 (N_6104,N_330,N_2438);
nand U6105 (N_6105,N_2818,N_2278);
xnor U6106 (N_6106,N_499,N_2533);
nand U6107 (N_6107,N_480,N_2240);
nor U6108 (N_6108,N_156,N_1517);
and U6109 (N_6109,N_1269,N_2101);
nor U6110 (N_6110,N_1439,N_1473);
or U6111 (N_6111,N_1493,N_2583);
nand U6112 (N_6112,N_1169,N_1046);
or U6113 (N_6113,N_1282,N_1042);
nor U6114 (N_6114,N_2841,N_1910);
xnor U6115 (N_6115,N_557,N_2757);
xor U6116 (N_6116,N_955,N_300);
nand U6117 (N_6117,N_1512,N_2906);
nor U6118 (N_6118,N_1001,N_375);
and U6119 (N_6119,N_618,N_2652);
nand U6120 (N_6120,N_53,N_721);
and U6121 (N_6121,N_1491,N_2531);
and U6122 (N_6122,N_79,N_546);
and U6123 (N_6123,N_2757,N_2788);
and U6124 (N_6124,N_2812,N_642);
nand U6125 (N_6125,N_295,N_1602);
nand U6126 (N_6126,N_309,N_3055);
or U6127 (N_6127,N_893,N_1671);
xnor U6128 (N_6128,N_217,N_1250);
nand U6129 (N_6129,N_1209,N_138);
xnor U6130 (N_6130,N_582,N_2005);
nor U6131 (N_6131,N_2431,N_2401);
or U6132 (N_6132,N_1428,N_1929);
and U6133 (N_6133,N_335,N_1593);
xor U6134 (N_6134,N_514,N_2086);
nor U6135 (N_6135,N_1657,N_2205);
and U6136 (N_6136,N_1345,N_2863);
nand U6137 (N_6137,N_2764,N_341);
nor U6138 (N_6138,N_71,N_538);
nor U6139 (N_6139,N_538,N_3001);
and U6140 (N_6140,N_1264,N_2023);
xor U6141 (N_6141,N_58,N_1807);
nand U6142 (N_6142,N_1554,N_2369);
nor U6143 (N_6143,N_1393,N_218);
nand U6144 (N_6144,N_1779,N_2114);
nand U6145 (N_6145,N_1336,N_625);
xnor U6146 (N_6146,N_2272,N_2986);
or U6147 (N_6147,N_125,N_1988);
and U6148 (N_6148,N_2676,N_1708);
and U6149 (N_6149,N_1704,N_1093);
and U6150 (N_6150,N_2263,N_1179);
nand U6151 (N_6151,N_677,N_2345);
xnor U6152 (N_6152,N_2774,N_149);
or U6153 (N_6153,N_336,N_1495);
xor U6154 (N_6154,N_335,N_205);
nand U6155 (N_6155,N_2891,N_1105);
or U6156 (N_6156,N_420,N_360);
or U6157 (N_6157,N_1098,N_3000);
xnor U6158 (N_6158,N_568,N_418);
or U6159 (N_6159,N_3038,N_180);
or U6160 (N_6160,N_2386,N_2713);
or U6161 (N_6161,N_1306,N_2146);
xnor U6162 (N_6162,N_586,N_2082);
or U6163 (N_6163,N_835,N_2873);
nand U6164 (N_6164,N_2749,N_1718);
and U6165 (N_6165,N_1589,N_849);
or U6166 (N_6166,N_2095,N_797);
nand U6167 (N_6167,N_2949,N_964);
nand U6168 (N_6168,N_2025,N_3100);
or U6169 (N_6169,N_2388,N_1407);
and U6170 (N_6170,N_1948,N_1464);
or U6171 (N_6171,N_994,N_1300);
and U6172 (N_6172,N_1490,N_1629);
nand U6173 (N_6173,N_2965,N_1571);
or U6174 (N_6174,N_1786,N_1351);
or U6175 (N_6175,N_1870,N_2749);
xnor U6176 (N_6176,N_63,N_1377);
or U6177 (N_6177,N_3052,N_1277);
and U6178 (N_6178,N_1084,N_306);
and U6179 (N_6179,N_934,N_2050);
or U6180 (N_6180,N_82,N_1587);
or U6181 (N_6181,N_255,N_1471);
xor U6182 (N_6182,N_779,N_2672);
nor U6183 (N_6183,N_1425,N_2642);
and U6184 (N_6184,N_2368,N_1290);
and U6185 (N_6185,N_897,N_681);
and U6186 (N_6186,N_2040,N_2140);
nand U6187 (N_6187,N_1904,N_452);
or U6188 (N_6188,N_42,N_2590);
nor U6189 (N_6189,N_2438,N_509);
and U6190 (N_6190,N_2520,N_1561);
and U6191 (N_6191,N_1982,N_1774);
nand U6192 (N_6192,N_1549,N_547);
and U6193 (N_6193,N_2497,N_681);
and U6194 (N_6194,N_2216,N_2551);
nor U6195 (N_6195,N_932,N_2617);
xor U6196 (N_6196,N_565,N_1864);
or U6197 (N_6197,N_2197,N_2359);
nor U6198 (N_6198,N_708,N_2856);
or U6199 (N_6199,N_1339,N_1073);
and U6200 (N_6200,N_1810,N_764);
and U6201 (N_6201,N_223,N_1423);
xnor U6202 (N_6202,N_3001,N_2971);
and U6203 (N_6203,N_1160,N_1726);
or U6204 (N_6204,N_2062,N_2292);
xnor U6205 (N_6205,N_2134,N_1186);
and U6206 (N_6206,N_2005,N_2842);
or U6207 (N_6207,N_1334,N_1743);
or U6208 (N_6208,N_1344,N_1038);
nand U6209 (N_6209,N_2642,N_1520);
xnor U6210 (N_6210,N_2317,N_2117);
nand U6211 (N_6211,N_368,N_665);
xor U6212 (N_6212,N_1674,N_955);
and U6213 (N_6213,N_2045,N_586);
nand U6214 (N_6214,N_1058,N_2621);
nand U6215 (N_6215,N_1337,N_3103);
and U6216 (N_6216,N_771,N_2321);
nand U6217 (N_6217,N_2208,N_2639);
nand U6218 (N_6218,N_1061,N_1842);
or U6219 (N_6219,N_440,N_132);
and U6220 (N_6220,N_484,N_2529);
xnor U6221 (N_6221,N_1236,N_1345);
nor U6222 (N_6222,N_1279,N_2618);
and U6223 (N_6223,N_152,N_1297);
and U6224 (N_6224,N_93,N_2865);
or U6225 (N_6225,N_872,N_992);
nand U6226 (N_6226,N_2809,N_2438);
and U6227 (N_6227,N_3030,N_677);
and U6228 (N_6228,N_1564,N_1049);
nand U6229 (N_6229,N_1387,N_1506);
and U6230 (N_6230,N_765,N_2861);
xor U6231 (N_6231,N_2747,N_2928);
nand U6232 (N_6232,N_1912,N_1195);
or U6233 (N_6233,N_2118,N_2287);
nand U6234 (N_6234,N_291,N_1159);
nor U6235 (N_6235,N_2143,N_2438);
and U6236 (N_6236,N_2661,N_890);
and U6237 (N_6237,N_143,N_2052);
xnor U6238 (N_6238,N_2492,N_2558);
and U6239 (N_6239,N_1118,N_2803);
nor U6240 (N_6240,N_2232,N_1246);
nor U6241 (N_6241,N_2330,N_1663);
or U6242 (N_6242,N_406,N_2416);
xnor U6243 (N_6243,N_2294,N_2856);
or U6244 (N_6244,N_1917,N_1160);
xnor U6245 (N_6245,N_1117,N_240);
or U6246 (N_6246,N_1250,N_1184);
xor U6247 (N_6247,N_1872,N_1943);
nor U6248 (N_6248,N_1938,N_169);
xor U6249 (N_6249,N_1664,N_1416);
nand U6250 (N_6250,N_3225,N_5980);
xor U6251 (N_6251,N_5993,N_5229);
nand U6252 (N_6252,N_3252,N_4473);
xnor U6253 (N_6253,N_4149,N_5770);
nand U6254 (N_6254,N_4675,N_5083);
nand U6255 (N_6255,N_3787,N_4871);
nand U6256 (N_6256,N_3561,N_4210);
nor U6257 (N_6257,N_3291,N_4360);
xnor U6258 (N_6258,N_4606,N_4730);
nand U6259 (N_6259,N_4094,N_4263);
nand U6260 (N_6260,N_3155,N_3442);
nand U6261 (N_6261,N_3952,N_4726);
or U6262 (N_6262,N_5403,N_4826);
nand U6263 (N_6263,N_4903,N_5413);
xnor U6264 (N_6264,N_4850,N_5658);
or U6265 (N_6265,N_3441,N_4275);
or U6266 (N_6266,N_6242,N_3609);
nand U6267 (N_6267,N_3314,N_4193);
nand U6268 (N_6268,N_3847,N_4357);
nor U6269 (N_6269,N_3264,N_4534);
or U6270 (N_6270,N_3914,N_5533);
or U6271 (N_6271,N_4757,N_5020);
or U6272 (N_6272,N_6158,N_4745);
nand U6273 (N_6273,N_4580,N_3910);
nor U6274 (N_6274,N_4371,N_5631);
or U6275 (N_6275,N_3200,N_4135);
xor U6276 (N_6276,N_3340,N_4869);
or U6277 (N_6277,N_5847,N_5066);
or U6278 (N_6278,N_5057,N_4996);
or U6279 (N_6279,N_6123,N_3204);
or U6280 (N_6280,N_4816,N_5481);
nor U6281 (N_6281,N_5349,N_4089);
or U6282 (N_6282,N_3182,N_6124);
nand U6283 (N_6283,N_4046,N_3529);
nand U6284 (N_6284,N_3604,N_5836);
or U6285 (N_6285,N_4634,N_4526);
nor U6286 (N_6286,N_3355,N_5292);
nand U6287 (N_6287,N_3147,N_5956);
xnor U6288 (N_6288,N_5394,N_6006);
xor U6289 (N_6289,N_6215,N_4594);
or U6290 (N_6290,N_4158,N_3421);
nand U6291 (N_6291,N_5855,N_5860);
or U6292 (N_6292,N_3364,N_5428);
nand U6293 (N_6293,N_3532,N_5414);
xnor U6294 (N_6294,N_5615,N_4027);
nand U6295 (N_6295,N_5086,N_3704);
xnor U6296 (N_6296,N_3190,N_5602);
nor U6297 (N_6297,N_5798,N_6004);
or U6298 (N_6298,N_5728,N_5887);
nand U6299 (N_6299,N_5402,N_3885);
nor U6300 (N_6300,N_3514,N_5144);
nor U6301 (N_6301,N_3668,N_5041);
and U6302 (N_6302,N_6220,N_5473);
and U6303 (N_6303,N_4909,N_4207);
nor U6304 (N_6304,N_5715,N_5900);
and U6305 (N_6305,N_6191,N_6164);
xnor U6306 (N_6306,N_4270,N_5737);
xnor U6307 (N_6307,N_4426,N_4103);
nand U6308 (N_6308,N_5157,N_5080);
nand U6309 (N_6309,N_5725,N_5444);
nand U6310 (N_6310,N_3217,N_3156);
nand U6311 (N_6311,N_3235,N_3886);
nand U6312 (N_6312,N_4657,N_4545);
nand U6313 (N_6313,N_5425,N_4699);
nor U6314 (N_6314,N_5613,N_5101);
nor U6315 (N_6315,N_5815,N_3231);
xnor U6316 (N_6316,N_4968,N_5743);
nand U6317 (N_6317,N_4319,N_5334);
nor U6318 (N_6318,N_4626,N_4057);
or U6319 (N_6319,N_4857,N_5659);
xor U6320 (N_6320,N_5825,N_3570);
and U6321 (N_6321,N_5657,N_4000);
nand U6322 (N_6322,N_3288,N_4405);
nor U6323 (N_6323,N_3989,N_3325);
nand U6324 (N_6324,N_3889,N_4115);
or U6325 (N_6325,N_5597,N_3500);
xor U6326 (N_6326,N_5548,N_3971);
and U6327 (N_6327,N_3319,N_4830);
nor U6328 (N_6328,N_5068,N_4333);
nand U6329 (N_6329,N_5799,N_5854);
or U6330 (N_6330,N_3766,N_3716);
nand U6331 (N_6331,N_3146,N_4544);
and U6332 (N_6332,N_4959,N_4465);
and U6333 (N_6333,N_5316,N_5146);
or U6334 (N_6334,N_5783,N_3328);
and U6335 (N_6335,N_4125,N_5485);
or U6336 (N_6336,N_4181,N_3650);
and U6337 (N_6337,N_5055,N_5243);
nand U6338 (N_6338,N_3483,N_5928);
nand U6339 (N_6339,N_3390,N_5518);
nor U6340 (N_6340,N_3911,N_3370);
or U6341 (N_6341,N_4225,N_3965);
nand U6342 (N_6342,N_3755,N_5383);
xor U6343 (N_6343,N_5257,N_4315);
nand U6344 (N_6344,N_5315,N_4852);
xor U6345 (N_6345,N_4940,N_4063);
and U6346 (N_6346,N_5116,N_4929);
xor U6347 (N_6347,N_3937,N_5733);
nor U6348 (N_6348,N_3138,N_4619);
nor U6349 (N_6349,N_4512,N_3440);
xor U6350 (N_6350,N_4382,N_3861);
or U6351 (N_6351,N_4993,N_5184);
nand U6352 (N_6352,N_3750,N_5430);
or U6353 (N_6353,N_3131,N_4229);
xor U6354 (N_6354,N_5270,N_3552);
or U6355 (N_6355,N_5271,N_3140);
or U6356 (N_6356,N_4530,N_4420);
or U6357 (N_6357,N_6175,N_4511);
nand U6358 (N_6358,N_5935,N_5756);
xnor U6359 (N_6359,N_4867,N_3218);
nor U6360 (N_6360,N_5189,N_4192);
nor U6361 (N_6361,N_5014,N_3259);
and U6362 (N_6362,N_6105,N_4246);
and U6363 (N_6363,N_4520,N_4516);
xor U6364 (N_6364,N_5067,N_3457);
nor U6365 (N_6365,N_5567,N_3664);
nand U6366 (N_6366,N_3625,N_4114);
nand U6367 (N_6367,N_4180,N_5065);
xnor U6368 (N_6368,N_5917,N_3667);
xnor U6369 (N_6369,N_5023,N_4839);
nand U6370 (N_6370,N_3834,N_5312);
or U6371 (N_6371,N_4444,N_5405);
nor U6372 (N_6372,N_4665,N_5497);
nand U6373 (N_6373,N_4820,N_5683);
or U6374 (N_6374,N_5447,N_4759);
xor U6375 (N_6375,N_4340,N_4196);
nor U6376 (N_6376,N_5303,N_4054);
nor U6377 (N_6377,N_5981,N_4779);
xnor U6378 (N_6378,N_3600,N_3841);
and U6379 (N_6379,N_4503,N_5151);
and U6380 (N_6380,N_3269,N_4195);
or U6381 (N_6381,N_3895,N_5311);
and U6382 (N_6382,N_3159,N_5620);
nor U6383 (N_6383,N_5344,N_3944);
and U6384 (N_6384,N_3286,N_5307);
and U6385 (N_6385,N_5685,N_5393);
xnor U6386 (N_6386,N_3682,N_3712);
nor U6387 (N_6387,N_5276,N_5761);
xor U6388 (N_6388,N_4936,N_3824);
or U6389 (N_6389,N_6082,N_4208);
xor U6390 (N_6390,N_5095,N_3747);
or U6391 (N_6391,N_4835,N_6161);
or U6392 (N_6392,N_3166,N_6093);
nand U6393 (N_6393,N_5472,N_4944);
or U6394 (N_6394,N_4965,N_3521);
and U6395 (N_6395,N_4716,N_4097);
nor U6396 (N_6396,N_5341,N_5650);
and U6397 (N_6397,N_3365,N_4219);
or U6398 (N_6398,N_5318,N_5532);
nor U6399 (N_6399,N_5289,N_5200);
xor U6400 (N_6400,N_4796,N_4399);
nand U6401 (N_6401,N_5872,N_5864);
and U6402 (N_6402,N_6075,N_3622);
and U6403 (N_6403,N_4264,N_5470);
xor U6404 (N_6404,N_3158,N_6016);
or U6405 (N_6405,N_4581,N_5585);
and U6406 (N_6406,N_3543,N_4577);
nor U6407 (N_6407,N_5668,N_4892);
xnor U6408 (N_6408,N_5118,N_3335);
nand U6409 (N_6409,N_5111,N_3617);
nand U6410 (N_6410,N_5009,N_4470);
or U6411 (N_6411,N_5480,N_3383);
xnor U6412 (N_6412,N_5734,N_5962);
nor U6413 (N_6413,N_3338,N_3608);
nand U6414 (N_6414,N_3707,N_5422);
xnor U6415 (N_6415,N_4744,N_5568);
xnor U6416 (N_6416,N_4065,N_4044);
or U6417 (N_6417,N_5489,N_4107);
nor U6418 (N_6418,N_4793,N_3374);
nand U6419 (N_6419,N_5600,N_3950);
and U6420 (N_6420,N_3362,N_3285);
nand U6421 (N_6421,N_5840,N_5436);
or U6422 (N_6422,N_3470,N_5103);
xor U6423 (N_6423,N_3638,N_5338);
xor U6424 (N_6424,N_4147,N_4937);
nand U6425 (N_6425,N_4754,N_5792);
xnor U6426 (N_6426,N_5274,N_5077);
or U6427 (N_6427,N_5508,N_5373);
and U6428 (N_6428,N_3693,N_4079);
xnor U6429 (N_6429,N_5535,N_5932);
xor U6430 (N_6430,N_5695,N_4277);
and U6431 (N_6431,N_5794,N_4553);
and U6432 (N_6432,N_5611,N_4926);
and U6433 (N_6433,N_4185,N_3385);
and U6434 (N_6434,N_5220,N_3813);
nand U6435 (N_6435,N_5176,N_5560);
or U6436 (N_6436,N_3498,N_4755);
nor U6437 (N_6437,N_3246,N_5022);
xnor U6438 (N_6438,N_4143,N_5700);
nor U6439 (N_6439,N_5329,N_4130);
nor U6440 (N_6440,N_6249,N_4279);
nand U6441 (N_6441,N_3560,N_4831);
nand U6442 (N_6442,N_4026,N_5681);
nor U6443 (N_6443,N_3864,N_4868);
nor U6444 (N_6444,N_6230,N_3884);
nor U6445 (N_6445,N_3628,N_4499);
nand U6446 (N_6446,N_5314,N_3292);
xor U6447 (N_6447,N_4407,N_4038);
nor U6448 (N_6448,N_3661,N_3271);
or U6449 (N_6449,N_5421,N_4408);
nand U6450 (N_6450,N_4659,N_4631);
and U6451 (N_6451,N_5596,N_3343);
nand U6452 (N_6452,N_4289,N_4660);
xor U6453 (N_6453,N_4756,N_5072);
xor U6454 (N_6454,N_6098,N_4463);
and U6455 (N_6455,N_4557,N_3918);
xor U6456 (N_6456,N_5539,N_3256);
and U6457 (N_6457,N_3783,N_5846);
nor U6458 (N_6458,N_5160,N_3781);
or U6459 (N_6459,N_5452,N_3236);
or U6460 (N_6460,N_5853,N_4596);
nand U6461 (N_6461,N_4623,N_5000);
nor U6462 (N_6462,N_5496,N_4785);
nand U6463 (N_6463,N_6059,N_3657);
or U6464 (N_6464,N_4108,N_5198);
nand U6465 (N_6465,N_4654,N_4256);
nor U6466 (N_6466,N_4422,N_5283);
xnor U6467 (N_6467,N_3729,N_3800);
or U6468 (N_6468,N_5167,N_5504);
xor U6469 (N_6469,N_5136,N_5375);
nor U6470 (N_6470,N_3565,N_3631);
nor U6471 (N_6471,N_4911,N_3582);
xor U6472 (N_6472,N_5340,N_6079);
or U6473 (N_6473,N_5032,N_5863);
nor U6474 (N_6474,N_3674,N_4259);
or U6475 (N_6475,N_4994,N_5925);
nand U6476 (N_6476,N_3391,N_3211);
xnor U6477 (N_6477,N_4050,N_4647);
nor U6478 (N_6478,N_6217,N_3192);
or U6479 (N_6479,N_3923,N_5260);
or U6480 (N_6480,N_5849,N_4638);
and U6481 (N_6481,N_5680,N_3724);
nand U6482 (N_6482,N_3473,N_5224);
and U6483 (N_6483,N_4471,N_4587);
nand U6484 (N_6484,N_3389,N_5453);
nor U6485 (N_6485,N_3411,N_5384);
or U6486 (N_6486,N_3445,N_4437);
and U6487 (N_6487,N_6214,N_3678);
nor U6488 (N_6488,N_5839,N_3614);
xor U6489 (N_6489,N_5360,N_5529);
and U6490 (N_6490,N_4295,N_4019);
and U6491 (N_6491,N_5305,N_5679);
or U6492 (N_6492,N_3405,N_4070);
xnor U6493 (N_6493,N_4554,N_4592);
xnor U6494 (N_6494,N_5476,N_4881);
xnor U6495 (N_6495,N_4972,N_4401);
nor U6496 (N_6496,N_6003,N_4244);
or U6497 (N_6497,N_4338,N_3170);
and U6498 (N_6498,N_3694,N_5026);
nor U6499 (N_6499,N_5324,N_4651);
nand U6500 (N_6500,N_6235,N_4339);
nand U6501 (N_6501,N_4069,N_5007);
nor U6502 (N_6502,N_4048,N_4737);
nor U6503 (N_6503,N_3949,N_6176);
and U6504 (N_6504,N_3127,N_4572);
xnor U6505 (N_6505,N_3804,N_5088);
nor U6506 (N_6506,N_3417,N_3202);
or U6507 (N_6507,N_6032,N_4591);
nor U6508 (N_6508,N_5630,N_5003);
and U6509 (N_6509,N_5502,N_3948);
nor U6510 (N_6510,N_3714,N_5286);
xor U6511 (N_6511,N_4569,N_3376);
and U6512 (N_6512,N_4578,N_6209);
nand U6513 (N_6513,N_4375,N_3629);
or U6514 (N_6514,N_5751,N_4062);
or U6515 (N_6515,N_5150,N_4679);
nand U6516 (N_6516,N_4469,N_5793);
xnor U6517 (N_6517,N_5262,N_5058);
nand U6518 (N_6518,N_3195,N_5653);
or U6519 (N_6519,N_3666,N_3808);
and U6520 (N_6520,N_4736,N_4693);
or U6521 (N_6521,N_4100,N_5181);
and U6522 (N_6522,N_3934,N_4507);
or U6523 (N_6523,N_5752,N_4589);
or U6524 (N_6524,N_5342,N_5309);
xnor U6525 (N_6525,N_3416,N_5845);
and U6526 (N_6526,N_3935,N_3515);
nor U6527 (N_6527,N_3562,N_3840);
and U6528 (N_6528,N_5127,N_6166);
nand U6529 (N_6529,N_4684,N_5703);
xnor U6530 (N_6530,N_4678,N_3566);
nor U6531 (N_6531,N_5805,N_3247);
and U6532 (N_6532,N_3660,N_5382);
xor U6533 (N_6533,N_5008,N_6101);
nand U6534 (N_6534,N_4200,N_3371);
xnor U6535 (N_6535,N_3904,N_3744);
and U6536 (N_6536,N_3439,N_5738);
and U6537 (N_6537,N_6226,N_3216);
or U6538 (N_6538,N_5905,N_4269);
nand U6539 (N_6539,N_6007,N_3702);
xnor U6540 (N_6540,N_5976,N_5191);
nand U6541 (N_6541,N_4637,N_6049);
nor U6542 (N_6542,N_3901,N_4935);
nor U6543 (N_6543,N_4919,N_3596);
nor U6544 (N_6544,N_5478,N_6145);
and U6545 (N_6545,N_4011,N_5520);
and U6546 (N_6546,N_5100,N_4024);
nand U6547 (N_6547,N_5048,N_4813);
nand U6548 (N_6548,N_3649,N_4539);
nand U6549 (N_6549,N_5284,N_4013);
nor U6550 (N_6550,N_5246,N_3654);
and U6551 (N_6551,N_4977,N_5339);
nand U6552 (N_6552,N_5780,N_5785);
and U6553 (N_6553,N_4117,N_5161);
or U6554 (N_6554,N_3799,N_3829);
or U6555 (N_6555,N_3485,N_3815);
or U6556 (N_6556,N_4917,N_5687);
or U6557 (N_6557,N_5711,N_5830);
and U6558 (N_6558,N_5484,N_4250);
or U6559 (N_6559,N_5878,N_4952);
and U6560 (N_6560,N_5186,N_3890);
nand U6561 (N_6561,N_3221,N_3577);
or U6562 (N_6562,N_4894,N_3451);
nand U6563 (N_6563,N_5590,N_4560);
xor U6564 (N_6564,N_3916,N_3822);
xor U6565 (N_6565,N_5219,N_5570);
nor U6566 (N_6566,N_5736,N_5786);
or U6567 (N_6567,N_5574,N_4309);
nand U6568 (N_6568,N_5215,N_4316);
nor U6569 (N_6569,N_6122,N_3873);
nor U6570 (N_6570,N_4843,N_3461);
nor U6571 (N_6571,N_3306,N_4663);
or U6572 (N_6572,N_3507,N_4688);
and U6573 (N_6573,N_4177,N_3867);
or U6574 (N_6574,N_3802,N_4846);
nor U6575 (N_6575,N_4624,N_5493);
or U6576 (N_6576,N_4153,N_4221);
nand U6577 (N_6577,N_5085,N_4049);
xor U6578 (N_6578,N_5275,N_5675);
or U6579 (N_6579,N_3234,N_4725);
and U6580 (N_6580,N_6018,N_3224);
nand U6581 (N_6581,N_5094,N_3506);
and U6582 (N_6582,N_4750,N_5998);
and U6583 (N_6583,N_5619,N_4567);
xor U6584 (N_6584,N_4808,N_5919);
or U6585 (N_6585,N_5718,N_4617);
or U6586 (N_6586,N_4670,N_4129);
nor U6587 (N_6587,N_4092,N_5945);
nand U6588 (N_6588,N_6083,N_4768);
nand U6589 (N_6589,N_5236,N_3871);
or U6590 (N_6590,N_4376,N_6223);
and U6591 (N_6591,N_4938,N_5731);
or U6592 (N_6592,N_3275,N_3710);
nor U6593 (N_6593,N_3511,N_4696);
nand U6594 (N_6594,N_4278,N_4329);
xor U6595 (N_6595,N_3266,N_4872);
nand U6596 (N_6596,N_3863,N_3375);
and U6597 (N_6597,N_6182,N_5944);
nor U6598 (N_6598,N_5479,N_3761);
and U6599 (N_6599,N_5359,N_5081);
xor U6600 (N_6600,N_4014,N_5129);
nor U6601 (N_6601,N_3180,N_5233);
nor U6602 (N_6602,N_3851,N_3825);
nand U6603 (N_6603,N_5208,N_5823);
xnor U6604 (N_6604,N_4713,N_4916);
nor U6605 (N_6605,N_4017,N_4967);
or U6606 (N_6606,N_3186,N_5278);
or U6607 (N_6607,N_5363,N_3776);
and U6608 (N_6608,N_3819,N_5955);
xnor U6609 (N_6609,N_3426,N_5506);
and U6610 (N_6610,N_5295,N_5656);
nand U6611 (N_6611,N_3606,N_5551);
xor U6612 (N_6612,N_5987,N_3768);
or U6613 (N_6613,N_6078,N_3648);
and U6614 (N_6614,N_4962,N_5367);
or U6615 (N_6615,N_6057,N_4220);
nand U6616 (N_6616,N_3139,N_5758);
nand U6617 (N_6617,N_5040,N_3663);
and U6618 (N_6618,N_3933,N_6070);
nand U6619 (N_6619,N_3765,N_5512);
nor U6620 (N_6620,N_3395,N_5120);
or U6621 (N_6621,N_3419,N_6150);
or U6622 (N_6622,N_3143,N_4337);
nor U6623 (N_6623,N_3311,N_3175);
nor U6624 (N_6624,N_3479,N_3164);
nand U6625 (N_6625,N_4483,N_4154);
and U6626 (N_6626,N_6021,N_4268);
and U6627 (N_6627,N_4897,N_4694);
nor U6628 (N_6628,N_4397,N_4173);
or U6629 (N_6629,N_5616,N_5643);
and U6630 (N_6630,N_5810,N_6110);
nand U6631 (N_6631,N_5104,N_4242);
or U6632 (N_6632,N_3359,N_4645);
nand U6633 (N_6633,N_5417,N_4136);
or U6634 (N_6634,N_6171,N_4294);
and U6635 (N_6635,N_4975,N_4595);
and U6636 (N_6636,N_3482,N_5709);
nor U6637 (N_6637,N_3459,N_4356);
and U6638 (N_6638,N_3887,N_3240);
nor U6639 (N_6639,N_5673,N_4383);
or U6640 (N_6640,N_5237,N_4308);
nor U6641 (N_6641,N_4817,N_4934);
nor U6642 (N_6642,N_5961,N_6151);
xor U6643 (N_6643,N_5556,N_3623);
nor U6644 (N_6644,N_3262,N_3484);
or U6645 (N_6645,N_4252,N_5951);
nand U6646 (N_6646,N_5689,N_3875);
nand U6647 (N_6647,N_5677,N_6241);
nand U6648 (N_6648,N_5832,N_4171);
and U6649 (N_6649,N_5017,N_5881);
and U6650 (N_6650,N_4441,N_5742);
nor U6651 (N_6651,N_4528,N_4406);
nor U6652 (N_6652,N_6060,N_3537);
and U6653 (N_6653,N_3436,N_3734);
nand U6654 (N_6654,N_5694,N_4486);
xor U6655 (N_6655,N_6100,N_4942);
nand U6656 (N_6656,N_5592,N_3399);
nor U6657 (N_6657,N_4671,N_5477);
and U6658 (N_6658,N_4690,N_3513);
nor U6659 (N_6659,N_3132,N_4535);
or U6660 (N_6660,N_5087,N_4387);
and U6661 (N_6661,N_4933,N_4317);
xnor U6662 (N_6662,N_5239,N_4332);
and U6663 (N_6663,N_3545,N_5922);
nand U6664 (N_6664,N_4343,N_5448);
nand U6665 (N_6665,N_3605,N_6170);
and U6666 (N_6666,N_3835,N_3151);
xor U6667 (N_6667,N_4468,N_4614);
or U6668 (N_6668,N_5416,N_3981);
nand U6669 (N_6669,N_5148,N_3926);
and U6670 (N_6670,N_4652,N_4385);
nand U6671 (N_6671,N_3534,N_4763);
nor U6672 (N_6672,N_6014,N_3850);
and U6673 (N_6673,N_4947,N_5222);
and U6674 (N_6674,N_3633,N_4840);
or U6675 (N_6675,N_4838,N_6087);
xor U6676 (N_6676,N_5440,N_6224);
nand U6677 (N_6677,N_5261,N_5851);
nor U6678 (N_6678,N_5230,N_3962);
or U6679 (N_6679,N_5979,N_6108);
nand U6680 (N_6680,N_5966,N_4081);
xnor U6681 (N_6681,N_5424,N_5531);
nor U6682 (N_6682,N_5105,N_5593);
and U6683 (N_6683,N_4982,N_4853);
xnor U6684 (N_6684,N_5024,N_3512);
nor U6685 (N_6685,N_3564,N_4106);
and U6686 (N_6686,N_3177,N_3982);
and U6687 (N_6687,N_5183,N_4178);
nand U6688 (N_6688,N_3632,N_5391);
xnor U6689 (N_6689,N_4293,N_3250);
nand U6690 (N_6690,N_5435,N_4218);
or U6691 (N_6691,N_5135,N_6157);
or U6692 (N_6692,N_5175,N_4893);
nor U6693 (N_6693,N_6073,N_3683);
or U6694 (N_6694,N_5698,N_5826);
nor U6695 (N_6695,N_5256,N_4474);
xnor U6696 (N_6696,N_4719,N_3305);
xor U6697 (N_6697,N_3637,N_5491);
and U6698 (N_6698,N_5691,N_6206);
or U6699 (N_6699,N_5902,N_5566);
and U6700 (N_6700,N_4334,N_3807);
or U6701 (N_6701,N_5062,N_5089);
and U6702 (N_6702,N_5906,N_6113);
xnor U6703 (N_6703,N_4832,N_5235);
and U6704 (N_6704,N_5883,N_5443);
or U6705 (N_6705,N_4734,N_6077);
nor U6706 (N_6706,N_4758,N_5714);
nor U6707 (N_6707,N_4562,N_3237);
nor U6708 (N_6708,N_3642,N_3220);
xor U6709 (N_6709,N_4425,N_4302);
xnor U6710 (N_6710,N_5720,N_5595);
nor U6711 (N_6711,N_3309,N_4604);
nor U6712 (N_6712,N_4751,N_5045);
nor U6713 (N_6713,N_4762,N_3762);
and U6714 (N_6714,N_4986,N_5407);
or U6715 (N_6715,N_4224,N_5494);
nor U6716 (N_6716,N_4039,N_5005);
xnor U6717 (N_6717,N_5251,N_3238);
or U6718 (N_6718,N_6198,N_3946);
and U6719 (N_6719,N_6172,N_3505);
nand U6720 (N_6720,N_6134,N_5459);
or U6721 (N_6721,N_5787,N_4951);
and U6722 (N_6722,N_5128,N_4007);
nor U6723 (N_6723,N_3640,N_3554);
or U6724 (N_6724,N_5126,N_3282);
nor U6725 (N_6725,N_4403,N_5130);
nand U6726 (N_6726,N_4601,N_3931);
xor U6727 (N_6727,N_5581,N_3881);
xnor U6728 (N_6728,N_3820,N_4016);
and U6729 (N_6729,N_3544,N_3454);
xnor U6730 (N_6730,N_6063,N_4849);
nand U6731 (N_6731,N_3626,N_5404);
nor U6732 (N_6732,N_6222,N_4320);
xor U6733 (N_6733,N_3351,N_4056);
xnor U6734 (N_6734,N_3809,N_4240);
xnor U6735 (N_6735,N_3277,N_3509);
nand U6736 (N_6736,N_6019,N_3902);
or U6737 (N_6737,N_6038,N_5368);
or U6738 (N_6738,N_3730,N_3478);
nand U6739 (N_6739,N_4747,N_4568);
or U6740 (N_6740,N_4508,N_4228);
and U6741 (N_6741,N_6035,N_5874);
nor U6742 (N_6742,N_3685,N_5612);
nand U6743 (N_6743,N_5795,N_3866);
xnor U6744 (N_6744,N_4841,N_5730);
nor U6745 (N_6745,N_3736,N_4430);
or U6746 (N_6746,N_4829,N_3341);
nand U6747 (N_6747,N_4448,N_4648);
or U6748 (N_6748,N_5877,N_5173);
and U6749 (N_6749,N_4365,N_3302);
and U6750 (N_6750,N_3510,N_4733);
xnor U6751 (N_6751,N_4212,N_4948);
and U6752 (N_6752,N_3208,N_4008);
nor U6753 (N_6753,N_4144,N_5899);
and U6754 (N_6754,N_5467,N_5753);
nor U6755 (N_6755,N_3369,N_6104);
and U6756 (N_6756,N_4174,N_3185);
or U6757 (N_6757,N_4707,N_5959);
and U6758 (N_6758,N_4131,N_5051);
nand U6759 (N_6759,N_3578,N_5999);
or U6760 (N_6760,N_5755,N_6202);
nor U6761 (N_6761,N_4067,N_5446);
xnor U6762 (N_6762,N_3174,N_5766);
and U6763 (N_6763,N_5121,N_4552);
or U6764 (N_6764,N_5776,N_6076);
nand U6765 (N_6765,N_3711,N_5850);
xnor U6766 (N_6766,N_6225,N_3969);
and U6767 (N_6767,N_4666,N_5573);
and U6768 (N_6768,N_4431,N_4137);
and U6769 (N_6769,N_4190,N_5242);
and U6770 (N_6770,N_4890,N_4211);
or U6771 (N_6771,N_4889,N_4668);
or U6772 (N_6772,N_4245,N_4021);
and U6773 (N_6773,N_5226,N_3812);
nor U6774 (N_6774,N_4418,N_3651);
or U6775 (N_6775,N_4451,N_6189);
nor U6776 (N_6776,N_4482,N_4402);
and U6777 (N_6777,N_4253,N_4002);
nand U6778 (N_6778,N_4656,N_5921);
nor U6779 (N_6779,N_5995,N_5699);
nor U6780 (N_6780,N_3517,N_3267);
and U6781 (N_6781,N_5117,N_5210);
or U6782 (N_6782,N_4206,N_4029);
nor U6783 (N_6783,N_6030,N_5973);
nand U6784 (N_6784,N_4574,N_5948);
or U6785 (N_6785,N_4718,N_6186);
nand U6786 (N_6786,N_4731,N_3464);
nor U6787 (N_6787,N_3244,N_5557);
nand U6788 (N_6788,N_4706,N_3976);
nor U6789 (N_6789,N_6195,N_4795);
and U6790 (N_6790,N_4477,N_5666);
or U6791 (N_6791,N_6129,N_4930);
and U6792 (N_6792,N_3187,N_4970);
nor U6793 (N_6793,N_6071,N_4939);
xor U6794 (N_6794,N_5796,N_3785);
and U6795 (N_6795,N_3641,N_5267);
or U6796 (N_6796,N_5124,N_3358);
nor U6797 (N_6797,N_5294,N_5598);
nand U6798 (N_6798,N_5941,N_5992);
nor U6799 (N_6799,N_4858,N_4961);
nand U6800 (N_6800,N_3646,N_5379);
nor U6801 (N_6801,N_3897,N_4182);
nor U6802 (N_6802,N_4685,N_4146);
nand U6803 (N_6803,N_4640,N_4901);
nor U6804 (N_6804,N_3432,N_5054);
xnor U6805 (N_6805,N_3833,N_3771);
and U6806 (N_6806,N_5063,N_4618);
nor U6807 (N_6807,N_4837,N_6103);
nand U6808 (N_6808,N_4603,N_3627);
or U6809 (N_6809,N_5500,N_5503);
xnor U6810 (N_6810,N_3831,N_5621);
or U6811 (N_6811,N_5577,N_4561);
xor U6812 (N_6812,N_4155,N_6152);
nor U6813 (N_6813,N_6155,N_6136);
or U6814 (N_6814,N_4262,N_6067);
nand U6815 (N_6815,N_6009,N_5434);
nand U6816 (N_6816,N_5091,N_5248);
xor U6817 (N_6817,N_3700,N_3437);
or U6818 (N_6818,N_5199,N_3842);
nand U6819 (N_6819,N_4184,N_5608);
nor U6820 (N_6820,N_5119,N_3675);
nand U6821 (N_6821,N_6207,N_4582);
or U6822 (N_6822,N_4045,N_4822);
nand U6823 (N_6823,N_3444,N_4746);
and U6824 (N_6824,N_5893,N_4336);
nand U6825 (N_6825,N_4998,N_5019);
or U6826 (N_6826,N_3449,N_3313);
or U6827 (N_6827,N_4394,N_4502);
nor U6828 (N_6828,N_5114,N_3924);
or U6829 (N_6829,N_3272,N_5693);
and U6830 (N_6830,N_3373,N_5523);
xor U6831 (N_6831,N_5591,N_3210);
nand U6832 (N_6832,N_3443,N_4845);
nor U6833 (N_6833,N_3689,N_3205);
xnor U6834 (N_6834,N_4384,N_5204);
nand U6835 (N_6835,N_5164,N_5519);
nor U6836 (N_6836,N_4099,N_5212);
and U6837 (N_6837,N_4980,N_3130);
or U6838 (N_6838,N_4722,N_4369);
and U6839 (N_6839,N_5377,N_3792);
nand U6840 (N_6840,N_4598,N_4605);
nand U6841 (N_6841,N_5745,N_4812);
xor U6842 (N_6842,N_3687,N_3838);
nand U6843 (N_6843,N_6232,N_3930);
nand U6844 (N_6844,N_5398,N_3307);
xor U6845 (N_6845,N_5876,N_4362);
xnor U6846 (N_6846,N_5464,N_4898);
or U6847 (N_6847,N_3721,N_4161);
nand U6848 (N_6848,N_5410,N_3476);
xnor U6849 (N_6849,N_5300,N_4292);
and U6850 (N_6850,N_3853,N_5814);
and U6851 (N_6851,N_4197,N_3731);
and U6852 (N_6852,N_4851,N_5115);
or U6853 (N_6853,N_5588,N_3435);
nor U6854 (N_6854,N_4819,N_5958);
nand U6855 (N_6855,N_3818,N_5923);
nand U6856 (N_6856,N_3496,N_3129);
and U6857 (N_6857,N_3882,N_3811);
nor U6858 (N_6858,N_4272,N_3584);
or U6859 (N_6859,N_4531,N_5056);
nand U6860 (N_6860,N_4030,N_3161);
xor U6861 (N_6861,N_6081,N_4653);
xor U6862 (N_6862,N_6041,N_3284);
xnor U6863 (N_6863,N_4781,N_5188);
nor U6864 (N_6864,N_4814,N_5559);
nand U6865 (N_6865,N_6000,N_5837);
and U6866 (N_6866,N_6120,N_6169);
xor U6867 (N_6867,N_3701,N_4818);
xnor U6868 (N_6868,N_3896,N_3985);
xor U6869 (N_6869,N_5607,N_4226);
nand U6870 (N_6870,N_4321,N_4882);
and U6871 (N_6871,N_4023,N_4836);
or U6872 (N_6872,N_6156,N_3839);
or U6873 (N_6873,N_5006,N_3852);
xor U6874 (N_6874,N_4954,N_3980);
nor U6875 (N_6875,N_3579,N_5174);
nand U6876 (N_6876,N_5717,N_4366);
nand U6877 (N_6877,N_6137,N_3974);
xor U6878 (N_6878,N_5449,N_5674);
and U6879 (N_6879,N_4035,N_3858);
or U6880 (N_6880,N_3688,N_4740);
nor U6881 (N_6881,N_5073,N_5280);
nor U6882 (N_6882,N_3927,N_5165);
or U6883 (N_6883,N_3898,N_5336);
nand U6884 (N_6884,N_5511,N_4140);
xor U6885 (N_6885,N_4995,N_5301);
or U6886 (N_6886,N_4299,N_5554);
nand U6887 (N_6887,N_5252,N_3332);
nand U6888 (N_6888,N_5254,N_5565);
or U6889 (N_6889,N_4563,N_3337);
nand U6890 (N_6890,N_3717,N_3795);
or U6891 (N_6891,N_3719,N_4711);
and U6892 (N_6892,N_4495,N_4692);
and U6893 (N_6893,N_4285,N_3758);
nand U6894 (N_6894,N_5552,N_4466);
nand U6895 (N_6895,N_5916,N_6002);
xor U6896 (N_6896,N_3438,N_4170);
nand U6897 (N_6897,N_3740,N_3676);
nand U6898 (N_6898,N_4481,N_4551);
or U6899 (N_6899,N_6142,N_6047);
or U6900 (N_6900,N_4419,N_6011);
nor U6901 (N_6901,N_3176,N_5910);
nand U6902 (N_6902,N_5697,N_4484);
or U6903 (N_6903,N_3764,N_4411);
nand U6904 (N_6904,N_5669,N_3477);
and U6905 (N_6905,N_4698,N_3352);
or U6906 (N_6906,N_5033,N_3967);
xor U6907 (N_6907,N_5895,N_4318);
and U6908 (N_6908,N_3726,N_4931);
and U6909 (N_6909,N_5950,N_3287);
or U6910 (N_6910,N_3535,N_3988);
nand U6911 (N_6911,N_4649,N_5092);
nand U6912 (N_6912,N_3699,N_3594);
xnor U6913 (N_6913,N_5990,N_5991);
xor U6914 (N_6914,N_4602,N_4296);
and U6915 (N_6915,N_5667,N_5972);
nand U6916 (N_6916,N_4548,N_5381);
xor U6917 (N_6917,N_3708,N_4241);
nor U6918 (N_6918,N_4990,N_5660);
xor U6919 (N_6919,N_5043,N_3751);
nand U6920 (N_6920,N_5937,N_3905);
xor U6921 (N_6921,N_4844,N_3480);
or U6922 (N_6922,N_4672,N_3893);
or U6923 (N_6923,N_3697,N_6162);
and U6924 (N_6924,N_5171,N_5155);
xnor U6925 (N_6925,N_3778,N_4257);
nand U6926 (N_6926,N_5486,N_4204);
or U6927 (N_6927,N_5744,N_4187);
nand U6928 (N_6928,N_5903,N_4667);
nand U6929 (N_6929,N_5706,N_4636);
nand U6930 (N_6930,N_4714,N_5152);
xnor U6931 (N_6931,N_6227,N_5399);
nand U6932 (N_6932,N_4913,N_4842);
xor U6933 (N_6933,N_4632,N_4689);
nand U6934 (N_6934,N_3384,N_4920);
nand U6935 (N_6935,N_5918,N_5202);
nor U6936 (N_6936,N_3748,N_4460);
xor U6937 (N_6937,N_3681,N_4729);
nand U6938 (N_6938,N_5870,N_5978);
xor U6939 (N_6939,N_5536,N_5661);
and U6940 (N_6940,N_3289,N_6183);
or U6941 (N_6941,N_3763,N_5265);
nand U6942 (N_6942,N_4395,N_4720);
nor U6943 (N_6943,N_5060,N_5885);
nor U6944 (N_6944,N_4509,N_5337);
nand U6945 (N_6945,N_3951,N_3420);
xnor U6946 (N_6946,N_4216,N_5888);
or U6947 (N_6947,N_4827,N_5866);
and U6948 (N_6948,N_3280,N_5763);
and U6949 (N_6949,N_4449,N_6187);
or U6950 (N_6950,N_4721,N_5460);
or U6951 (N_6951,N_3686,N_3531);
xor U6952 (N_6952,N_4232,N_3703);
nor U6953 (N_6953,N_6005,N_5070);
xnor U6954 (N_6954,N_3869,N_6116);
nand U6955 (N_6955,N_6036,N_5018);
nand U6956 (N_6956,N_5401,N_3524);
xnor U6957 (N_6957,N_3466,N_4875);
nor U6958 (N_6958,N_5325,N_4612);
xor U6959 (N_6959,N_4527,N_5084);
nor U6960 (N_6960,N_4464,N_5211);
nor U6961 (N_6961,N_5039,N_4393);
and U6962 (N_6962,N_4176,N_3945);
nor U6963 (N_6963,N_3888,N_4148);
nor U6964 (N_6964,N_3742,N_5564);
nor U6965 (N_6965,N_5187,N_4536);
xor U6966 (N_6966,N_4367,N_5047);
or U6967 (N_6967,N_3141,N_5159);
or U6968 (N_6968,N_5926,N_3261);
nor U6969 (N_6969,N_3372,N_3919);
xnor U6970 (N_6970,N_5369,N_4786);
xor U6971 (N_6971,N_3490,N_6160);
and U6972 (N_6972,N_3644,N_5561);
and U6973 (N_6973,N_3458,N_4453);
or U6974 (N_6974,N_3601,N_4347);
or U6975 (N_6975,N_5521,N_4074);
or U6976 (N_6976,N_4203,N_3907);
nor U6977 (N_6977,N_6148,N_4330);
or U6978 (N_6978,N_6221,N_5201);
nor U6979 (N_6979,N_6178,N_4194);
nand U6980 (N_6980,N_4791,N_3705);
nor U6981 (N_6981,N_5828,N_5896);
or U6982 (N_6982,N_4121,N_4811);
xor U6983 (N_6983,N_3572,N_5385);
nand U6984 (N_6984,N_5050,N_3488);
nand U6985 (N_6985,N_5587,N_4001);
xnor U6986 (N_6986,N_5423,N_4724);
or U6987 (N_6987,N_5784,N_4620);
nand U6988 (N_6988,N_4416,N_4078);
xnor U6989 (N_6989,N_3403,N_4611);
nor U6990 (N_6990,N_3413,N_3157);
and U6991 (N_6991,N_3669,N_3961);
and U6992 (N_6992,N_3388,N_6084);
nor U6993 (N_6993,N_4879,N_5195);
and U6994 (N_6994,N_3856,N_3854);
nor U6995 (N_6995,N_4607,N_3784);
and U6996 (N_6996,N_3214,N_4124);
and U6997 (N_6997,N_3806,N_5203);
nor U6998 (N_6998,N_3541,N_5791);
nand U6999 (N_6999,N_5663,N_3733);
and U7000 (N_7000,N_3163,N_4036);
xnor U7001 (N_7001,N_4072,N_3251);
xor U7002 (N_7002,N_3308,N_4379);
xor U7003 (N_7003,N_4139,N_6210);
and U7004 (N_7004,N_5488,N_4515);
nand U7005 (N_7005,N_5406,N_5331);
or U7006 (N_7006,N_4798,N_5907);
nand U7007 (N_7007,N_3230,N_3909);
nor U7008 (N_7008,N_5190,N_4848);
or U7009 (N_7009,N_4300,N_5821);
xor U7010 (N_7010,N_4609,N_6159);
nor U7011 (N_7011,N_5617,N_5357);
or U7012 (N_7012,N_6168,N_4127);
or U7013 (N_7013,N_4742,N_5579);
nand U7014 (N_7014,N_3181,N_3749);
nand U7015 (N_7015,N_4088,N_3573);
nor U7016 (N_7016,N_4325,N_3722);
xor U7017 (N_7017,N_4311,N_3990);
or U7018 (N_7018,N_5372,N_4958);
xnor U7019 (N_7019,N_3983,N_4400);
and U7020 (N_7020,N_3558,N_6010);
nor U7021 (N_7021,N_3677,N_3786);
nor U7022 (N_7022,N_3547,N_4803);
nor U7023 (N_7023,N_6143,N_4927);
and U7024 (N_7024,N_5690,N_4433);
xor U7025 (N_7025,N_5671,N_4924);
nand U7026 (N_7026,N_4303,N_4538);
xor U7027 (N_7027,N_4492,N_3964);
and U7028 (N_7028,N_4828,N_5739);
xnor U7029 (N_7029,N_4753,N_5240);
nand U7030 (N_7030,N_4058,N_5727);
and U7031 (N_7031,N_6147,N_5293);
and U7032 (N_7032,N_5974,N_4997);
nor U7033 (N_7033,N_3448,N_4168);
nand U7034 (N_7034,N_3922,N_6243);
nor U7035 (N_7035,N_5516,N_5015);
and U7036 (N_7036,N_5765,N_5412);
xor U7037 (N_7037,N_3878,N_5064);
nand U7038 (N_7038,N_5390,N_3398);
and U7039 (N_7039,N_5614,N_3533);
nor U7040 (N_7040,N_4905,N_4209);
and U7041 (N_7041,N_5358,N_5652);
xnor U7042 (N_7042,N_3659,N_5938);
or U7043 (N_7043,N_3900,N_3692);
nand U7044 (N_7044,N_5010,N_5802);
nand U7045 (N_7045,N_3320,N_4255);
and U7046 (N_7046,N_4372,N_4172);
xnor U7047 (N_7047,N_6043,N_3862);
nand U7048 (N_7048,N_5985,N_4227);
or U7049 (N_7049,N_5306,N_6128);
or U7050 (N_7050,N_5740,N_5323);
nand U7051 (N_7051,N_5769,N_3446);
nor U7052 (N_7052,N_5433,N_3273);
xor U7053 (N_7053,N_4966,N_4584);
and U7054 (N_7054,N_5356,N_3920);
or U7055 (N_7055,N_3720,N_4133);
xnor U7056 (N_7056,N_5954,N_3408);
xnor U7057 (N_7057,N_6188,N_6048);
and U7058 (N_7058,N_4943,N_5253);
xnor U7059 (N_7059,N_3868,N_4529);
nand U7060 (N_7060,N_5983,N_5163);
or U7061 (N_7061,N_3455,N_3406);
nand U7062 (N_7062,N_3986,N_5196);
and U7063 (N_7063,N_5797,N_6244);
and U7064 (N_7064,N_4031,N_5166);
xnor U7065 (N_7065,N_5712,N_4415);
xnor U7066 (N_7066,N_6131,N_5857);
and U7067 (N_7067,N_4434,N_5268);
or U7068 (N_7068,N_3300,N_3415);
nand U7069 (N_7069,N_6132,N_3212);
xnor U7070 (N_7070,N_3645,N_4462);
xor U7071 (N_7071,N_5911,N_3404);
or U7072 (N_7072,N_3142,N_4251);
nor U7073 (N_7073,N_4664,N_5288);
nand U7074 (N_7074,N_4805,N_4518);
or U7075 (N_7075,N_5192,N_3450);
xor U7076 (N_7076,N_3805,N_4579);
or U7077 (N_7077,N_5636,N_3723);
or U7078 (N_7078,N_3789,N_3345);
and U7079 (N_7079,N_3489,N_4313);
xnor U7080 (N_7080,N_5353,N_4532);
xnor U7081 (N_7081,N_5078,N_3329);
and U7082 (N_7082,N_4412,N_5626);
and U7083 (N_7083,N_4476,N_4585);
xor U7084 (N_7084,N_4728,N_4307);
and U7085 (N_7085,N_3226,N_5330);
xnor U7086 (N_7086,N_5411,N_5361);
and U7087 (N_7087,N_6192,N_4351);
xor U7088 (N_7088,N_6072,N_5934);
or U7089 (N_7089,N_5772,N_5678);
or U7090 (N_7090,N_5483,N_3586);
nand U7091 (N_7091,N_3497,N_6177);
nand U7092 (N_7092,N_4712,N_5931);
and U7093 (N_7093,N_4424,N_3526);
or U7094 (N_7094,N_5313,N_3612);
or U7095 (N_7095,N_3936,N_5844);
and U7096 (N_7096,N_6008,N_6119);
nand U7097 (N_7097,N_5492,N_4613);
xor U7098 (N_7098,N_5259,N_3752);
nor U7099 (N_7099,N_4784,N_4646);
xnor U7100 (N_7100,N_5782,N_4373);
nand U7101 (N_7101,N_4417,N_6139);
or U7102 (N_7102,N_3670,N_5380);
or U7103 (N_7103,N_5156,N_6085);
and U7104 (N_7104,N_5609,N_4600);
nor U7105 (N_7105,N_5455,N_3519);
or U7106 (N_7106,N_4655,N_5969);
nand U7107 (N_7107,N_5264,N_4110);
nand U7108 (N_7108,N_4436,N_5310);
nor U7109 (N_7109,N_4885,N_4126);
nand U7110 (N_7110,N_5471,N_6111);
nor U7111 (N_7111,N_3152,N_6031);
nor U7112 (N_7112,N_4374,N_3598);
and U7113 (N_7113,N_6236,N_5131);
or U7114 (N_7114,N_3263,N_4327);
xor U7115 (N_7115,N_3360,N_5320);
or U7116 (N_7116,N_4974,N_4151);
nor U7117 (N_7117,N_3150,N_5811);
nor U7118 (N_7118,N_4950,N_5638);
nand U7119 (N_7119,N_5546,N_5635);
or U7120 (N_7120,N_4273,N_5030);
xnor U7121 (N_7121,N_4566,N_5122);
nand U7122 (N_7122,N_4314,N_4877);
and U7123 (N_7123,N_4141,N_5771);
or U7124 (N_7124,N_3381,N_3463);
or U7125 (N_7125,N_4547,N_4428);
nand U7126 (N_7126,N_3298,N_5831);
or U7127 (N_7127,N_5370,N_4949);
or U7128 (N_7128,N_6020,N_4546);
nand U7129 (N_7129,N_3652,N_5507);
xnor U7130 (N_7130,N_4205,N_5490);
or U7131 (N_7131,N_4150,N_6228);
nor U7132 (N_7132,N_3382,N_3844);
xnor U7133 (N_7133,N_3199,N_4423);
xor U7134 (N_7134,N_4517,N_3879);
nor U7135 (N_7135,N_4398,N_3334);
nand U7136 (N_7136,N_4335,N_3603);
or U7137 (N_7137,N_4522,N_5960);
xnor U7138 (N_7138,N_4138,N_4459);
xnor U7139 (N_7139,N_5505,N_5474);
and U7140 (N_7140,N_5153,N_4723);
nand U7141 (N_7141,N_3709,N_4500);
nor U7142 (N_7142,N_4261,N_4608);
or U7143 (N_7143,N_5942,N_5862);
nand U7144 (N_7144,N_3274,N_3732);
and U7145 (N_7145,N_5589,N_4310);
and U7146 (N_7146,N_3770,N_3304);
and U7147 (N_7147,N_3422,N_3301);
and U7148 (N_7148,N_3991,N_5431);
and U7149 (N_7149,N_3571,N_5705);
xor U7150 (N_7150,N_4378,N_3330);
xnor U7151 (N_7151,N_4167,N_6054);
nor U7152 (N_7152,N_3607,N_6027);
nand U7153 (N_7153,N_4790,N_4291);
nand U7154 (N_7154,N_3323,N_5646);
xnor U7155 (N_7155,N_3243,N_3975);
nor U7156 (N_7156,N_5541,N_5082);
and U7157 (N_7157,N_4865,N_4777);
and U7158 (N_7158,N_4708,N_5037);
nor U7159 (N_7159,N_5255,N_3213);
nor U7160 (N_7160,N_3239,N_3567);
xnor U7161 (N_7161,N_5046,N_5266);
and U7162 (N_7162,N_5967,N_3525);
nand U7163 (N_7163,N_4955,N_3754);
xor U7164 (N_7164,N_5290,N_4988);
nand U7165 (N_7165,N_5527,N_3401);
and U7166 (N_7166,N_5818,N_4941);
or U7167 (N_7167,N_4162,N_4891);
xnor U7168 (N_7168,N_5618,N_4095);
xor U7169 (N_7169,N_4134,N_3992);
or U7170 (N_7170,N_6037,N_3520);
nand U7171 (N_7171,N_5984,N_5170);
or U7172 (N_7172,N_3662,N_4377);
nand U7173 (N_7173,N_5285,N_6052);
nand U7174 (N_7174,N_3363,N_5145);
and U7175 (N_7175,N_4231,N_5781);
nor U7176 (N_7176,N_6013,N_4680);
xor U7177 (N_7177,N_4908,N_4105);
and U7178 (N_7178,N_4860,N_4748);
xor U7179 (N_7179,N_5696,N_3465);
and U7180 (N_7180,N_3928,N_4284);
nor U7181 (N_7181,N_5898,N_4804);
or U7182 (N_7182,N_6140,N_3634);
nor U7183 (N_7183,N_4346,N_4249);
and U7184 (N_7184,N_4286,N_5584);
nand U7185 (N_7185,N_3791,N_5466);
xor U7186 (N_7186,N_5540,N_4077);
and U7187 (N_7187,N_4080,N_3283);
nor U7188 (N_7188,N_5915,N_6180);
or U7189 (N_7189,N_6201,N_5890);
or U7190 (N_7190,N_4673,N_3523);
nor U7191 (N_7191,N_3679,N_4643);
and U7192 (N_7192,N_3940,N_3219);
nand U7193 (N_7193,N_4348,N_4328);
or U7194 (N_7194,N_4570,N_5816);
xnor U7195 (N_7195,N_4989,N_4918);
nand U7196 (N_7196,N_4489,N_3877);
xor U7197 (N_7197,N_6066,N_5319);
and U7198 (N_7198,N_4661,N_5789);
nor U7199 (N_7199,N_3312,N_4564);
nor U7200 (N_7200,N_3917,N_3874);
xnor U7201 (N_7201,N_5482,N_4104);
nand U7202 (N_7202,N_5125,N_4455);
or U7203 (N_7203,N_6154,N_5858);
xnor U7204 (N_7204,N_3528,N_5197);
or U7205 (N_7205,N_4490,N_3493);
xor U7206 (N_7206,N_4976,N_3491);
or U7207 (N_7207,N_3647,N_4345);
nor U7208 (N_7208,N_3743,N_4438);
nand U7209 (N_7209,N_5004,N_3128);
or U7210 (N_7210,N_5366,N_4076);
nand U7211 (N_7211,N_5889,N_5522);
nand U7212 (N_7212,N_5247,N_5949);
or U7213 (N_7213,N_5625,N_5028);
and U7214 (N_7214,N_3899,N_5879);
and U7215 (N_7215,N_6023,N_3794);
xnor U7216 (N_7216,N_3207,N_4283);
and U7217 (N_7217,N_4404,N_6212);
and U7218 (N_7218,N_6229,N_5975);
nor U7219 (N_7219,N_5069,N_3836);
or U7220 (N_7220,N_3378,N_4979);
and U7221 (N_7221,N_3303,N_6029);
nand U7222 (N_7222,N_5813,N_5576);
xor U7223 (N_7223,N_3698,N_3745);
and U7224 (N_7224,N_4388,N_3979);
xnor U7225 (N_7225,N_4349,N_4214);
or U7226 (N_7226,N_3184,N_3728);
or U7227 (N_7227,N_5465,N_3494);
nor U7228 (N_7228,N_3790,N_4041);
nand U7229 (N_7229,N_4112,N_5515);
xnor U7230 (N_7230,N_3258,N_4003);
nor U7231 (N_7231,N_3684,N_6231);
nand U7232 (N_7232,N_4597,N_3209);
or U7233 (N_7233,N_3848,N_3706);
or U7234 (N_7234,N_3602,N_5741);
or U7235 (N_7235,N_5297,N_3613);
nand U7236 (N_7236,N_3796,N_5684);
or U7237 (N_7237,N_3892,N_5649);
nand U7238 (N_7238,N_5670,N_6034);
nand U7239 (N_7239,N_3630,N_5133);
or U7240 (N_7240,N_4364,N_3295);
or U7241 (N_7241,N_5346,N_5134);
and U7242 (N_7242,N_5750,N_4969);
or U7243 (N_7243,N_4776,N_3366);
or U7244 (N_7244,N_3581,N_5812);
nor U7245 (N_7245,N_4715,N_4238);
xnor U7246 (N_7246,N_5132,N_4700);
or U7247 (N_7247,N_4410,N_5904);
nand U7248 (N_7248,N_3133,N_4432);
xor U7249 (N_7249,N_4789,N_4635);
xor U7250 (N_7250,N_4739,N_3165);
nand U7251 (N_7251,N_5871,N_6117);
or U7252 (N_7252,N_5437,N_3620);
nor U7253 (N_7253,N_4217,N_3316);
nor U7254 (N_7254,N_4494,N_3135);
xnor U7255 (N_7255,N_6194,N_5225);
nor U7256 (N_7256,N_5308,N_3793);
nand U7257 (N_7257,N_6141,N_5462);
nor U7258 (N_7258,N_5400,N_3656);
and U7259 (N_7259,N_4165,N_5158);
xor U7260 (N_7260,N_4324,N_5141);
nor U7261 (N_7261,N_3843,N_5637);
nor U7262 (N_7262,N_5534,N_3592);
or U7263 (N_7263,N_5525,N_4358);
xor U7264 (N_7264,N_5605,N_3148);
and U7265 (N_7265,N_5610,N_3580);
and U7266 (N_7266,N_5775,N_5732);
xnor U7267 (N_7267,N_4442,N_3741);
and U7268 (N_7268,N_4355,N_5767);
xor U7269 (N_7269,N_5807,N_3144);
xor U7270 (N_7270,N_4301,N_6204);
nor U7271 (N_7271,N_5777,N_3953);
or U7272 (N_7272,N_6239,N_4156);
or U7273 (N_7273,N_4787,N_3189);
nor U7274 (N_7274,N_3680,N_4501);
nor U7275 (N_7275,N_4625,N_5553);
or U7276 (N_7276,N_5322,N_3746);
and U7277 (N_7277,N_6135,N_5647);
and U7278 (N_7278,N_4928,N_5364);
nand U7279 (N_7279,N_5345,N_4824);
nor U7280 (N_7280,N_4119,N_4306);
nor U7281 (N_7281,N_3803,N_5013);
and U7282 (N_7282,N_4899,N_3349);
and U7283 (N_7283,N_4887,N_5764);
xnor U7284 (N_7284,N_6091,N_4735);
nor U7285 (N_7285,N_4902,N_4222);
nor U7286 (N_7286,N_6247,N_4354);
xor U7287 (N_7287,N_5509,N_3255);
and U7288 (N_7288,N_5321,N_4274);
or U7289 (N_7289,N_3447,N_3775);
nand U7290 (N_7290,N_5272,N_6112);
nand U7291 (N_7291,N_5547,N_3407);
nand U7292 (N_7292,N_5279,N_4287);
xnor U7293 (N_7293,N_5747,N_4878);
xor U7294 (N_7294,N_5450,N_4704);
or U7295 (N_7295,N_4610,N_4599);
xor U7296 (N_7296,N_4098,N_4485);
and U7297 (N_7297,N_5542,N_5628);
nor U7298 (N_7298,N_3474,N_3801);
or U7299 (N_7299,N_4142,N_4505);
nor U7300 (N_7300,N_5790,N_3178);
xor U7301 (N_7301,N_3522,N_5843);
nor U7302 (N_7302,N_3658,N_3938);
xnor U7303 (N_7303,N_3757,N_4331);
and U7304 (N_7304,N_3756,N_4621);
nand U7305 (N_7305,N_4863,N_5644);
or U7306 (N_7306,N_5052,N_4874);
and U7307 (N_7307,N_5415,N_6064);
nor U7308 (N_7308,N_5442,N_4519);
or U7309 (N_7309,N_5957,N_3427);
and U7310 (N_7310,N_3551,N_4297);
xnor U7311 (N_7311,N_5147,N_3941);
xor U7312 (N_7312,N_5571,N_4963);
or U7313 (N_7313,N_5149,N_5820);
and U7314 (N_7314,N_5031,N_4549);
or U7315 (N_7315,N_5475,N_4896);
nand U7316 (N_7316,N_4802,N_5920);
nand U7317 (N_7317,N_4052,N_6133);
and U7318 (N_7318,N_4487,N_4288);
nor U7319 (N_7319,N_3431,N_3915);
nor U7320 (N_7320,N_5397,N_4859);
xnor U7321 (N_7321,N_5108,N_3859);
xor U7322 (N_7322,N_4370,N_3615);
nand U7323 (N_7323,N_3984,N_6102);
xor U7324 (N_7324,N_5989,N_6001);
and U7325 (N_7325,N_5106,N_5172);
xnor U7326 (N_7326,N_4101,N_4981);
and U7327 (N_7327,N_5099,N_4235);
and U7328 (N_7328,N_5362,N_4461);
xor U7329 (N_7329,N_4550,N_5389);
nand U7330 (N_7330,N_3471,N_4510);
xor U7331 (N_7331,N_5376,N_5193);
and U7332 (N_7332,N_5946,N_5749);
nor U7333 (N_7333,N_4380,N_5138);
or U7334 (N_7334,N_5833,N_6179);
and U7335 (N_7335,N_5185,N_6080);
nand U7336 (N_7336,N_5606,N_6046);
nor U7337 (N_7337,N_4102,N_3814);
nor U7338 (N_7338,N_3715,N_5169);
or U7339 (N_7339,N_3995,N_5408);
or U7340 (N_7340,N_4179,N_3206);
nor U7341 (N_7341,N_5291,N_3162);
and U7342 (N_7342,N_4234,N_3423);
or U7343 (N_7343,N_6033,N_3997);
nor U7344 (N_7344,N_4213,N_4973);
nor U7345 (N_7345,N_3501,N_6238);
and U7346 (N_7346,N_3963,N_5774);
nand U7347 (N_7347,N_5298,N_3908);
xor U7348 (N_7348,N_3837,N_4305);
and U7349 (N_7349,N_5514,N_3883);
xnor U7350 (N_7350,N_5206,N_4391);
xor U7351 (N_7351,N_4323,N_4281);
and U7352 (N_7352,N_5545,N_5528);
xor U7353 (N_7353,N_3585,N_3241);
or U7354 (N_7354,N_3357,N_4783);
nor U7355 (N_7355,N_3616,N_3499);
nor U7356 (N_7356,N_4576,N_4475);
and U7357 (N_7357,N_4764,N_3870);
and U7358 (N_7358,N_4732,N_4421);
nand U7359 (N_7359,N_5648,N_6099);
nor U7360 (N_7360,N_3549,N_4066);
nor U7361 (N_7361,N_6090,N_4188);
or U7362 (N_7362,N_4683,N_5469);
xor U7363 (N_7363,N_6245,N_4254);
xnor U7364 (N_7364,N_5838,N_5963);
and U7365 (N_7365,N_4012,N_6024);
nor U7366 (N_7366,N_5829,N_5662);
nand U7367 (N_7367,N_4923,N_6203);
nor U7368 (N_7368,N_5042,N_4794);
or U7369 (N_7369,N_3960,N_5386);
nand U7370 (N_7370,N_4160,N_3179);
and U7371 (N_7371,N_3321,N_5258);
or U7372 (N_7372,N_6109,N_5392);
nor U7373 (N_7373,N_3538,N_5808);
xnor U7374 (N_7374,N_3987,N_4342);
xor U7375 (N_7375,N_3590,N_5599);
nand U7376 (N_7376,N_4043,N_5027);
xnor U7377 (N_7377,N_3845,N_4265);
or U7378 (N_7378,N_4856,N_3278);
xnor U7379 (N_7379,N_6055,N_5988);
nand U7380 (N_7380,N_5665,N_4590);
xor U7381 (N_7381,N_5374,N_4034);
nor U7382 (N_7382,N_3188,N_3530);
nor U7383 (N_7383,N_3925,N_3618);
nand U7384 (N_7384,N_4042,N_5757);
nor U7385 (N_7385,N_4677,N_6086);
nor U7386 (N_7386,N_3559,N_4953);
or U7387 (N_7387,N_3760,N_5651);
nand U7388 (N_7388,N_4248,N_4760);
nor U7389 (N_7389,N_3414,N_5550);
xnor U7390 (N_7390,N_6149,N_3487);
xnor U7391 (N_7391,N_5335,N_5035);
nand U7392 (N_7392,N_4266,N_4687);
nor U7393 (N_7393,N_6126,N_4641);
xnor U7394 (N_7394,N_4571,N_5686);
nor U7395 (N_7395,N_3735,N_6028);
nor U7396 (N_7396,N_6015,N_6053);
nor U7397 (N_7397,N_4615,N_3168);
nand U7398 (N_7398,N_5578,N_5327);
and U7399 (N_7399,N_4189,N_3773);
nand U7400 (N_7400,N_5760,N_4005);
or U7401 (N_7401,N_5641,N_5273);
nor U7402 (N_7402,N_5943,N_5947);
nor U7403 (N_7403,N_5634,N_4533);
or U7404 (N_7404,N_5632,N_4166);
nand U7405 (N_7405,N_5001,N_4392);
xor U7406 (N_7406,N_4086,N_6062);
xor U7407 (N_7407,N_5371,N_4964);
xnor U7408 (N_7408,N_4068,N_3589);
or U7409 (N_7409,N_4120,N_4191);
xnor U7410 (N_7410,N_3553,N_3460);
nor U7411 (N_7411,N_4386,N_4506);
and U7412 (N_7412,N_5365,N_3453);
or U7413 (N_7413,N_5012,N_3690);
or U7414 (N_7414,N_3380,N_3593);
or U7415 (N_7415,N_5387,N_5759);
and U7416 (N_7416,N_5707,N_4873);
nand U7417 (N_7417,N_5704,N_6074);
or U7418 (N_7418,N_5891,N_4093);
or U7419 (N_7419,N_4341,N_4223);
nand U7420 (N_7420,N_5326,N_5965);
xnor U7421 (N_7421,N_5708,N_5594);
or U7422 (N_7422,N_4907,N_4888);
and U7423 (N_7423,N_6121,N_3145);
xnor U7424 (N_7424,N_4493,N_3550);
or U7425 (N_7425,N_3193,N_4326);
nor U7426 (N_7426,N_5468,N_5445);
nor U7427 (N_7427,N_4087,N_5487);
or U7428 (N_7428,N_3137,N_3412);
xnor U7429 (N_7429,N_3429,N_4409);
nand U7430 (N_7430,N_3518,N_3410);
nand U7431 (N_7431,N_3223,N_4801);
nor U7432 (N_7432,N_3996,N_4025);
xor U7433 (N_7433,N_5213,N_6012);
nand U7434 (N_7434,N_5562,N_5097);
xor U7435 (N_7435,N_4691,N_3611);
xnor U7436 (N_7436,N_3233,N_3418);
xnor U7437 (N_7437,N_3228,N_3939);
or U7438 (N_7438,N_3673,N_3621);
nor U7439 (N_7439,N_3527,N_5822);
nand U7440 (N_7440,N_4866,N_6095);
xor U7441 (N_7441,N_5729,N_5457);
nand U7442 (N_7442,N_5655,N_5762);
or U7443 (N_7443,N_5396,N_4091);
xor U7444 (N_7444,N_6017,N_4312);
xnor U7445 (N_7445,N_3171,N_3978);
nand U7446 (N_7446,N_3279,N_5865);
and U7447 (N_7447,N_4004,N_5848);
or U7448 (N_7448,N_3942,N_3957);
nor U7449 (N_7449,N_5061,N_4985);
nand U7450 (N_7450,N_4513,N_4984);
nor U7451 (N_7451,N_4109,N_5701);
nor U7452 (N_7452,N_3356,N_4010);
nor U7453 (N_7453,N_4033,N_6107);
nor U7454 (N_7454,N_3828,N_5842);
and U7455 (N_7455,N_3977,N_4669);
nand U7456 (N_7456,N_5180,N_3956);
or U7457 (N_7457,N_4132,N_6246);
nor U7458 (N_7458,N_4414,N_4910);
nand U7459 (N_7459,N_3568,N_5735);
or U7460 (N_7460,N_6025,N_6174);
nand U7461 (N_7461,N_6190,N_5263);
and U7462 (N_7462,N_5601,N_5439);
xnor U7463 (N_7463,N_5924,N_4703);
or U7464 (N_7464,N_6056,N_4864);
nor U7465 (N_7465,N_6199,N_4773);
xnor U7466 (N_7466,N_3229,N_4389);
xnor U7467 (N_7467,N_5107,N_3932);
nor U7468 (N_7468,N_4630,N_3392);
xnor U7469 (N_7469,N_5719,N_4202);
nor U7470 (N_7470,N_4983,N_6118);
xnor U7471 (N_7471,N_3597,N_3575);
nor U7472 (N_7472,N_4815,N_4524);
or U7473 (N_7473,N_4239,N_3947);
nand U7474 (N_7474,N_3467,N_5722);
nand U7475 (N_7475,N_3548,N_4116);
xnor U7476 (N_7476,N_4847,N_4472);
or U7477 (N_7477,N_5930,N_4390);
or U7478 (N_7478,N_6184,N_5530);
nand U7479 (N_7479,N_4083,N_3906);
nand U7480 (N_7480,N_6061,N_4788);
and U7481 (N_7481,N_4053,N_3318);
nand U7482 (N_7482,N_4123,N_5544);
nand U7483 (N_7483,N_5501,N_3830);
nor U7484 (N_7484,N_4697,N_3772);
and U7485 (N_7485,N_4061,N_5801);
xor U7486 (N_7486,N_5140,N_5016);
or U7487 (N_7487,N_3959,N_3368);
nand U7488 (N_7488,N_5296,N_3402);
or U7489 (N_7489,N_3574,N_4020);
nor U7490 (N_7490,N_5079,N_4201);
nand U7491 (N_7491,N_3610,N_5090);
or U7492 (N_7492,N_4932,N_4573);
xnor U7493 (N_7493,N_5074,N_3160);
xor U7494 (N_7494,N_4771,N_4575);
and U7495 (N_7495,N_3994,N_4260);
nand U7496 (N_7496,N_5970,N_5513);
and U7497 (N_7497,N_5179,N_5304);
nand U7498 (N_7498,N_4946,N_3780);
nor U7499 (N_7499,N_5723,N_4922);
nor U7500 (N_7500,N_4681,N_5021);
xor U7501 (N_7501,N_5277,N_5726);
or U7502 (N_7502,N_3153,N_3587);
xor U7503 (N_7503,N_3149,N_5154);
xor U7504 (N_7504,N_5558,N_3782);
or U7505 (N_7505,N_4113,N_5672);
nor U7506 (N_7506,N_5645,N_5526);
xnor U7507 (N_7507,N_5986,N_4458);
nand U7508 (N_7508,N_4247,N_3253);
xnor U7509 (N_7509,N_5964,N_5178);
and U7510 (N_7510,N_5517,N_4267);
and U7511 (N_7511,N_4028,N_4298);
nor U7512 (N_7512,N_3810,N_5419);
nor U7513 (N_7513,N_5835,N_4622);
nor U7514 (N_7514,N_3386,N_5044);
nor U7515 (N_7515,N_4778,N_4290);
nor U7516 (N_7516,N_4543,N_4823);
or U7517 (N_7517,N_5269,N_4686);
and U7518 (N_7518,N_3336,N_5788);
or U7519 (N_7519,N_4541,N_5458);
nand U7520 (N_7520,N_3196,N_5702);
nand U7521 (N_7521,N_3943,N_3452);
and U7522 (N_7522,N_3475,N_3342);
nor U7523 (N_7523,N_4639,N_4230);
nand U7524 (N_7524,N_5463,N_5333);
xor U7525 (N_7525,N_5038,N_4705);
nand U7526 (N_7526,N_3821,N_5429);
and U7527 (N_7527,N_3817,N_3400);
xnor U7528 (N_7528,N_4457,N_5827);
and U7529 (N_7529,N_5328,N_5555);
or U7530 (N_7530,N_6130,N_3317);
nand U7531 (N_7531,N_3348,N_6115);
nor U7532 (N_7532,N_5249,N_4912);
nor U7533 (N_7533,N_3583,N_3563);
xor U7534 (N_7534,N_5137,N_5778);
or U7535 (N_7535,N_5886,N_4304);
nor U7536 (N_7536,N_3966,N_3331);
and U7537 (N_7537,N_3860,N_3929);
xnor U7538 (N_7538,N_3958,N_3198);
nand U7539 (N_7539,N_3556,N_5228);
and U7540 (N_7540,N_3242,N_5768);
nor U7541 (N_7541,N_6237,N_3347);
or U7542 (N_7542,N_5388,N_6197);
xor U7543 (N_7543,N_5461,N_5287);
nand U7544 (N_7544,N_4440,N_5299);
or U7545 (N_7545,N_3713,N_5441);
xor U7546 (N_7546,N_5688,N_4770);
and U7547 (N_7547,N_4709,N_3767);
or U7548 (N_7548,N_4987,N_4454);
nor U7549 (N_7549,N_4479,N_4456);
or U7550 (N_7550,N_5250,N_3788);
nand U7551 (N_7551,N_3265,N_3326);
and U7552 (N_7552,N_5897,N_4854);
and U7553 (N_7553,N_5112,N_3434);
and U7554 (N_7554,N_4175,N_3999);
or U7555 (N_7555,N_4157,N_5537);
and U7556 (N_7556,N_4413,N_5912);
and U7557 (N_7557,N_3276,N_6040);
nand U7558 (N_7558,N_3393,N_5817);
or U7559 (N_7559,N_5034,N_3595);
xnor U7560 (N_7560,N_4883,N_4738);
nor U7561 (N_7561,N_5623,N_3154);
xor U7562 (N_7562,N_4629,N_5892);
nor U7563 (N_7563,N_6205,N_4445);
nor U7564 (N_7564,N_3425,N_3769);
or U7565 (N_7565,N_4055,N_4521);
or U7566 (N_7566,N_4833,N_5395);
nor U7567 (N_7567,N_6216,N_4583);
and U7568 (N_7568,N_6248,N_4085);
and U7569 (N_7569,N_3718,N_4825);
nand U7570 (N_7570,N_5350,N_4352);
or U7571 (N_7571,N_4593,N_4775);
xor U7572 (N_7572,N_5968,N_4233);
and U7573 (N_7573,N_3481,N_4525);
nand U7574 (N_7574,N_5682,N_6213);
nor U7575 (N_7575,N_5347,N_4855);
xnor U7576 (N_7576,N_6218,N_5011);
and U7577 (N_7577,N_4145,N_4090);
nand U7578 (N_7578,N_3855,N_4957);
nor U7579 (N_7579,N_5244,N_6193);
or U7580 (N_7580,N_3469,N_3346);
and U7581 (N_7581,N_3691,N_3655);
or U7582 (N_7582,N_4556,N_5873);
nand U7583 (N_7583,N_3639,N_5676);
nand U7584 (N_7584,N_5096,N_5909);
xor U7585 (N_7585,N_6088,N_3245);
nand U7586 (N_7586,N_4496,N_5710);
or U7587 (N_7587,N_4199,N_3913);
or U7588 (N_7588,N_4682,N_4588);
or U7589 (N_7589,N_4164,N_5971);
and U7590 (N_7590,N_4051,N_6167);
xor U7591 (N_7591,N_5868,N_5162);
nor U7592 (N_7592,N_5994,N_4642);
and U7593 (N_7593,N_5803,N_3665);
nand U7594 (N_7594,N_5563,N_4710);
or U7595 (N_7595,N_5076,N_4766);
nand U7596 (N_7596,N_4555,N_4780);
or U7597 (N_7597,N_4558,N_5102);
nand U7598 (N_7598,N_3502,N_4198);
xnor U7599 (N_7599,N_4396,N_3468);
nand U7600 (N_7600,N_4047,N_3993);
nor U7601 (N_7601,N_5029,N_5852);
or U7602 (N_7602,N_3268,N_5317);
or U7603 (N_7603,N_5809,N_4633);
and U7604 (N_7604,N_3894,N_4806);
and U7605 (N_7605,N_4032,N_6173);
nand U7606 (N_7606,N_5880,N_4271);
or U7607 (N_7607,N_4956,N_5583);
nor U7608 (N_7608,N_5627,N_6181);
and U7609 (N_7609,N_3968,N_5859);
or U7610 (N_7610,N_4540,N_6125);
or U7611 (N_7611,N_5834,N_5586);
or U7612 (N_7612,N_3322,N_4807);
and U7613 (N_7613,N_3636,N_5427);
or U7614 (N_7614,N_5582,N_5779);
nor U7615 (N_7615,N_5953,N_3424);
nand U7616 (N_7616,N_6146,N_4800);
or U7617 (N_7617,N_5575,N_5754);
nand U7618 (N_7618,N_3849,N_4040);
or U7619 (N_7619,N_5059,N_5231);
and U7620 (N_7620,N_4792,N_4163);
nand U7621 (N_7621,N_4183,N_5332);
nand U7622 (N_7622,N_5214,N_6094);
nand U7623 (N_7623,N_3396,N_6165);
and U7624 (N_7624,N_5221,N_5624);
nor U7625 (N_7625,N_4018,N_3387);
or U7626 (N_7626,N_6044,N_4467);
or U7627 (N_7627,N_5952,N_3557);
nor U7628 (N_7628,N_3260,N_4236);
or U7629 (N_7629,N_5352,N_3327);
nand U7630 (N_7630,N_5901,N_4446);
nor U7631 (N_7631,N_4435,N_5438);
nor U7632 (N_7632,N_3296,N_3576);
nand U7633 (N_7633,N_4978,N_4662);
nand U7634 (N_7634,N_6208,N_5913);
xnor U7635 (N_7635,N_4443,N_5245);
nand U7636 (N_7636,N_3294,N_4862);
nand U7637 (N_7637,N_4084,N_5216);
nand U7638 (N_7638,N_3759,N_5420);
nor U7639 (N_7639,N_4429,N_6138);
or U7640 (N_7640,N_4999,N_4559);
and U7641 (N_7641,N_3495,N_4650);
nand U7642 (N_7642,N_5773,N_4169);
nand U7643 (N_7643,N_5861,N_4900);
xnor U7644 (N_7644,N_3591,N_4497);
and U7645 (N_7645,N_3281,N_5234);
nand U7646 (N_7646,N_5075,N_5495);
xnor U7647 (N_7647,N_3134,N_4616);
xor U7648 (N_7648,N_3293,N_3299);
nand U7649 (N_7649,N_5841,N_4925);
xor U7650 (N_7650,N_5348,N_3394);
nor U7651 (N_7651,N_3173,N_4075);
and U7652 (N_7652,N_3672,N_5177);
xor U7653 (N_7653,N_4243,N_4960);
xnor U7654 (N_7654,N_4628,N_3880);
nand U7655 (N_7655,N_3857,N_5168);
xnor U7656 (N_7656,N_4701,N_5908);
xnor U7657 (N_7657,N_3569,N_3492);
or U7658 (N_7658,N_5824,N_4799);
or U7659 (N_7659,N_3876,N_4749);
or U7660 (N_7660,N_4353,N_3191);
nor U7661 (N_7661,N_3169,N_4674);
or U7662 (N_7662,N_4870,N_5205);
and U7663 (N_7663,N_6211,N_5543);
nor U7664 (N_7664,N_5281,N_5025);
nor U7665 (N_7665,N_3826,N_5640);
and U7666 (N_7666,N_3955,N_3891);
xnor U7667 (N_7667,N_4884,N_5927);
and U7668 (N_7668,N_3344,N_4752);
nor U7669 (N_7669,N_5354,N_4809);
nor U7670 (N_7670,N_3409,N_4782);
nor U7671 (N_7671,N_3290,N_4904);
nand U7672 (N_7672,N_3430,N_3727);
or U7673 (N_7673,N_4258,N_3739);
or U7674 (N_7674,N_3970,N_5110);
and U7675 (N_7675,N_3354,N_4914);
nand U7676 (N_7676,N_4368,N_4498);
xor U7677 (N_7677,N_5432,N_4658);
nor U7678 (N_7678,N_6127,N_6196);
xor U7679 (N_7679,N_3248,N_5139);
or U7680 (N_7680,N_3194,N_4797);
xor U7681 (N_7681,N_4060,N_4186);
or U7682 (N_7682,N_3921,N_5227);
xor U7683 (N_7683,N_5232,N_5238);
or U7684 (N_7684,N_4322,N_4991);
xnor U7685 (N_7685,N_3197,N_3539);
and U7686 (N_7686,N_4876,N_3954);
nor U7687 (N_7687,N_4504,N_5142);
or U7688 (N_7688,N_3695,N_4915);
nor U7689 (N_7689,N_3973,N_5982);
nand U7690 (N_7690,N_5207,N_3397);
nand U7691 (N_7691,N_5894,N_4514);
or U7692 (N_7692,N_6114,N_5977);
nor U7693 (N_7693,N_4774,N_5499);
xnor U7694 (N_7694,N_6045,N_4359);
xor U7695 (N_7695,N_3433,N_4717);
and U7696 (N_7696,N_4767,N_5933);
or U7697 (N_7697,N_3777,N_5875);
nand U7698 (N_7698,N_3125,N_5806);
xnor U7699 (N_7699,N_4073,N_4009);
nor U7700 (N_7700,N_4128,N_3797);
xnor U7701 (N_7701,N_5182,N_5642);
or U7702 (N_7702,N_6089,N_3738);
xnor U7703 (N_7703,N_6240,N_3508);
xor U7704 (N_7704,N_5748,N_3428);
nand U7705 (N_7705,N_5716,N_4280);
nor U7706 (N_7706,N_4523,N_5936);
xor U7707 (N_7707,N_5939,N_4361);
nor U7708 (N_7708,N_5113,N_3297);
and U7709 (N_7709,N_5002,N_5569);
xnor U7710 (N_7710,N_4761,N_4447);
and U7711 (N_7711,N_4282,N_5223);
or U7712 (N_7712,N_3798,N_4743);
nor U7713 (N_7713,N_3136,N_4015);
and U7714 (N_7714,N_3599,N_3201);
or U7715 (N_7715,N_4152,N_3536);
nand U7716 (N_7716,N_3203,N_5538);
or U7717 (N_7717,N_5633,N_5036);
or U7718 (N_7718,N_6022,N_4880);
or U7719 (N_7719,N_6097,N_4676);
nand U7720 (N_7720,N_4765,N_3361);
or U7721 (N_7721,N_5524,N_5217);
or U7722 (N_7722,N_3753,N_3696);
nand U7723 (N_7723,N_4537,N_5549);
xnor U7724 (N_7724,N_3270,N_5724);
xnor U7725 (N_7725,N_3315,N_4059);
xnor U7726 (N_7726,N_3486,N_3555);
or U7727 (N_7727,N_5418,N_6219);
and U7728 (N_7728,N_3635,N_3816);
and U7729 (N_7729,N_5218,N_6234);
or U7730 (N_7730,N_5604,N_3588);
or U7731 (N_7731,N_3516,N_3172);
xor U7732 (N_7732,N_6144,N_4491);
or U7733 (N_7733,N_3903,N_4344);
nand U7734 (N_7734,N_5884,N_5882);
nor U7735 (N_7735,N_5804,N_4037);
nand U7736 (N_7736,N_5093,N_4006);
nor U7737 (N_7737,N_5664,N_3624);
and U7738 (N_7738,N_4542,N_3462);
and U7739 (N_7739,N_3254,N_3379);
xor U7740 (N_7740,N_6096,N_3367);
or U7741 (N_7741,N_4741,N_3872);
xnor U7742 (N_7742,N_4834,N_3671);
xor U7743 (N_7743,N_5869,N_4096);
xor U7744 (N_7744,N_4478,N_3324);
or U7745 (N_7745,N_5098,N_3333);
nand U7746 (N_7746,N_3546,N_3504);
nand U7747 (N_7747,N_4350,N_3542);
nor U7748 (N_7748,N_5143,N_4215);
nand U7749 (N_7749,N_5451,N_4810);
nand U7750 (N_7750,N_6153,N_3998);
and U7751 (N_7751,N_3827,N_5929);
and U7752 (N_7752,N_5194,N_4159);
nor U7753 (N_7753,N_6233,N_4439);
and U7754 (N_7754,N_5071,N_4071);
or U7755 (N_7755,N_5572,N_4821);
and U7756 (N_7756,N_5622,N_3737);
and U7757 (N_7757,N_3972,N_3472);
or U7758 (N_7758,N_4122,N_4118);
nand U7759 (N_7759,N_4565,N_4695);
and U7760 (N_7760,N_3249,N_3619);
and U7761 (N_7761,N_3865,N_3353);
nand U7762 (N_7762,N_3823,N_3540);
or U7763 (N_7763,N_3643,N_4480);
xnor U7764 (N_7764,N_5049,N_3456);
or U7765 (N_7765,N_5109,N_6058);
nand U7766 (N_7766,N_4276,N_3503);
and U7767 (N_7767,N_5996,N_4971);
nand U7768 (N_7768,N_5426,N_4064);
or U7769 (N_7769,N_3779,N_4772);
and U7770 (N_7770,N_4427,N_3257);
or U7771 (N_7771,N_4906,N_5454);
xor U7772 (N_7772,N_4644,N_5282);
and U7773 (N_7773,N_3222,N_3846);
or U7774 (N_7774,N_5914,N_3377);
xnor U7775 (N_7775,N_4363,N_4237);
xnor U7776 (N_7776,N_5378,N_5302);
nand U7777 (N_7777,N_5819,N_3774);
nor U7778 (N_7778,N_5997,N_6050);
and U7779 (N_7779,N_4452,N_5510);
or U7780 (N_7780,N_5721,N_4586);
and U7781 (N_7781,N_4702,N_3832);
and U7782 (N_7782,N_4861,N_4921);
nand U7783 (N_7783,N_5603,N_4727);
or U7784 (N_7784,N_4111,N_3232);
and U7785 (N_7785,N_6026,N_4488);
xor U7786 (N_7786,N_6039,N_6185);
or U7787 (N_7787,N_5856,N_3725);
and U7788 (N_7788,N_6068,N_3167);
nor U7789 (N_7789,N_4627,N_6200);
nand U7790 (N_7790,N_3310,N_4450);
nand U7791 (N_7791,N_3912,N_5713);
nand U7792 (N_7792,N_4381,N_5456);
nand U7793 (N_7793,N_5343,N_3350);
nor U7794 (N_7794,N_5209,N_3339);
nor U7795 (N_7795,N_5053,N_5580);
or U7796 (N_7796,N_4769,N_5498);
and U7797 (N_7797,N_4082,N_6065);
nor U7798 (N_7798,N_5940,N_5409);
xor U7799 (N_7799,N_3126,N_4886);
nor U7800 (N_7800,N_5692,N_3227);
and U7801 (N_7801,N_4022,N_6092);
nand U7802 (N_7802,N_4945,N_5746);
xnor U7803 (N_7803,N_4992,N_5123);
and U7804 (N_7804,N_6163,N_3653);
and U7805 (N_7805,N_5629,N_5800);
nor U7806 (N_7806,N_5867,N_6106);
and U7807 (N_7807,N_5639,N_6051);
nand U7808 (N_7808,N_5654,N_5241);
xor U7809 (N_7809,N_5355,N_4895);
or U7810 (N_7810,N_5351,N_6069);
xnor U7811 (N_7811,N_3183,N_3215);
nor U7812 (N_7812,N_6042,N_5941);
or U7813 (N_7813,N_4948,N_4202);
xor U7814 (N_7814,N_4765,N_4371);
or U7815 (N_7815,N_5623,N_4492);
xor U7816 (N_7816,N_5526,N_6006);
nor U7817 (N_7817,N_4357,N_6024);
nor U7818 (N_7818,N_3612,N_4337);
nor U7819 (N_7819,N_5294,N_4547);
or U7820 (N_7820,N_4923,N_4829);
nand U7821 (N_7821,N_4102,N_3173);
nand U7822 (N_7822,N_4587,N_4809);
and U7823 (N_7823,N_4518,N_6096);
nor U7824 (N_7824,N_4832,N_5431);
or U7825 (N_7825,N_4062,N_6097);
nand U7826 (N_7826,N_3924,N_5507);
nand U7827 (N_7827,N_5712,N_3956);
or U7828 (N_7828,N_4284,N_6145);
nor U7829 (N_7829,N_4165,N_5890);
and U7830 (N_7830,N_4729,N_3700);
nor U7831 (N_7831,N_3194,N_3274);
nand U7832 (N_7832,N_5979,N_5465);
and U7833 (N_7833,N_5863,N_4921);
nor U7834 (N_7834,N_4529,N_4162);
nor U7835 (N_7835,N_5417,N_4303);
xnor U7836 (N_7836,N_4922,N_4005);
nand U7837 (N_7837,N_3815,N_4169);
and U7838 (N_7838,N_3877,N_3303);
nor U7839 (N_7839,N_3632,N_5029);
and U7840 (N_7840,N_4931,N_6165);
nand U7841 (N_7841,N_4237,N_5956);
or U7842 (N_7842,N_6123,N_6162);
or U7843 (N_7843,N_3454,N_5665);
xnor U7844 (N_7844,N_5512,N_5345);
nor U7845 (N_7845,N_5228,N_5998);
or U7846 (N_7846,N_5614,N_5714);
xor U7847 (N_7847,N_3190,N_3781);
xnor U7848 (N_7848,N_3362,N_3395);
nor U7849 (N_7849,N_4759,N_5765);
nand U7850 (N_7850,N_4954,N_6118);
or U7851 (N_7851,N_5665,N_5712);
and U7852 (N_7852,N_3900,N_5315);
nand U7853 (N_7853,N_5588,N_5704);
and U7854 (N_7854,N_3331,N_5766);
nand U7855 (N_7855,N_3891,N_5285);
xnor U7856 (N_7856,N_5425,N_4369);
nor U7857 (N_7857,N_4934,N_6010);
and U7858 (N_7858,N_6134,N_4630);
and U7859 (N_7859,N_5411,N_5699);
nor U7860 (N_7860,N_5836,N_3323);
nor U7861 (N_7861,N_3327,N_4237);
and U7862 (N_7862,N_6078,N_5685);
and U7863 (N_7863,N_4349,N_3612);
and U7864 (N_7864,N_4024,N_4964);
xor U7865 (N_7865,N_3728,N_5442);
xnor U7866 (N_7866,N_5637,N_3899);
nor U7867 (N_7867,N_3236,N_3861);
nor U7868 (N_7868,N_4903,N_4614);
xnor U7869 (N_7869,N_4646,N_4685);
nand U7870 (N_7870,N_3524,N_4995);
or U7871 (N_7871,N_4016,N_5919);
xor U7872 (N_7872,N_5633,N_5419);
or U7873 (N_7873,N_5470,N_3367);
nand U7874 (N_7874,N_4356,N_3199);
or U7875 (N_7875,N_5488,N_5867);
nand U7876 (N_7876,N_5265,N_4419);
or U7877 (N_7877,N_3655,N_5904);
xor U7878 (N_7878,N_4784,N_5837);
nor U7879 (N_7879,N_4594,N_3282);
or U7880 (N_7880,N_3555,N_5704);
or U7881 (N_7881,N_4085,N_3828);
nor U7882 (N_7882,N_5457,N_4820);
nor U7883 (N_7883,N_4843,N_3990);
nand U7884 (N_7884,N_5289,N_5642);
xnor U7885 (N_7885,N_5770,N_5163);
nor U7886 (N_7886,N_5386,N_3801);
xor U7887 (N_7887,N_3836,N_3468);
and U7888 (N_7888,N_4558,N_5032);
nor U7889 (N_7889,N_3511,N_3675);
or U7890 (N_7890,N_5169,N_6241);
nor U7891 (N_7891,N_4757,N_3944);
nor U7892 (N_7892,N_5943,N_5717);
nand U7893 (N_7893,N_4379,N_3526);
or U7894 (N_7894,N_5055,N_3326);
nand U7895 (N_7895,N_5249,N_4265);
xnor U7896 (N_7896,N_5926,N_4753);
xnor U7897 (N_7897,N_6060,N_5951);
or U7898 (N_7898,N_5700,N_3547);
nand U7899 (N_7899,N_6205,N_3792);
and U7900 (N_7900,N_5668,N_3669);
nor U7901 (N_7901,N_5218,N_5983);
nand U7902 (N_7902,N_4515,N_3952);
and U7903 (N_7903,N_4881,N_4281);
xnor U7904 (N_7904,N_4619,N_4559);
nand U7905 (N_7905,N_3209,N_3412);
nand U7906 (N_7906,N_4566,N_6225);
nand U7907 (N_7907,N_5687,N_3610);
or U7908 (N_7908,N_3341,N_4821);
xor U7909 (N_7909,N_5164,N_5675);
nand U7910 (N_7910,N_4508,N_6191);
nor U7911 (N_7911,N_5682,N_4889);
or U7912 (N_7912,N_4744,N_5329);
and U7913 (N_7913,N_3212,N_6073);
nor U7914 (N_7914,N_3234,N_6154);
or U7915 (N_7915,N_4911,N_4165);
xnor U7916 (N_7916,N_3960,N_4170);
nor U7917 (N_7917,N_3999,N_4661);
nor U7918 (N_7918,N_4899,N_5042);
xor U7919 (N_7919,N_4856,N_4426);
nor U7920 (N_7920,N_5827,N_5417);
xor U7921 (N_7921,N_3248,N_4360);
or U7922 (N_7922,N_3659,N_4815);
and U7923 (N_7923,N_3931,N_3531);
xor U7924 (N_7924,N_4343,N_3955);
nor U7925 (N_7925,N_4792,N_3252);
or U7926 (N_7926,N_5679,N_4373);
and U7927 (N_7927,N_4202,N_5578);
xnor U7928 (N_7928,N_4084,N_4796);
nor U7929 (N_7929,N_5688,N_4021);
nand U7930 (N_7930,N_6110,N_3212);
xor U7931 (N_7931,N_4988,N_4776);
nor U7932 (N_7932,N_5220,N_3254);
nor U7933 (N_7933,N_3932,N_5284);
nand U7934 (N_7934,N_3361,N_4659);
nand U7935 (N_7935,N_5769,N_5991);
nand U7936 (N_7936,N_4408,N_5759);
nor U7937 (N_7937,N_6120,N_4440);
nor U7938 (N_7938,N_4094,N_4096);
nor U7939 (N_7939,N_5321,N_3402);
nor U7940 (N_7940,N_4532,N_4708);
nand U7941 (N_7941,N_5947,N_3911);
nor U7942 (N_7942,N_5850,N_3527);
nand U7943 (N_7943,N_3513,N_3147);
xnor U7944 (N_7944,N_5993,N_4738);
nand U7945 (N_7945,N_6113,N_4811);
xor U7946 (N_7946,N_4969,N_5844);
xnor U7947 (N_7947,N_5065,N_4610);
and U7948 (N_7948,N_3157,N_4800);
nand U7949 (N_7949,N_4768,N_3803);
and U7950 (N_7950,N_5654,N_5952);
nor U7951 (N_7951,N_3258,N_4157);
and U7952 (N_7952,N_4646,N_3370);
and U7953 (N_7953,N_4195,N_4303);
xnor U7954 (N_7954,N_3391,N_6139);
and U7955 (N_7955,N_5003,N_3924);
and U7956 (N_7956,N_4177,N_5776);
nor U7957 (N_7957,N_4856,N_5143);
nand U7958 (N_7958,N_5034,N_4863);
xor U7959 (N_7959,N_5441,N_4136);
nor U7960 (N_7960,N_3494,N_4269);
or U7961 (N_7961,N_5769,N_5122);
or U7962 (N_7962,N_3632,N_5441);
nand U7963 (N_7963,N_6032,N_5769);
xor U7964 (N_7964,N_4668,N_5785);
nand U7965 (N_7965,N_4414,N_5300);
or U7966 (N_7966,N_4329,N_3948);
nand U7967 (N_7967,N_3286,N_4927);
and U7968 (N_7968,N_5991,N_3835);
nor U7969 (N_7969,N_4036,N_3946);
or U7970 (N_7970,N_5862,N_3533);
xnor U7971 (N_7971,N_5084,N_4438);
and U7972 (N_7972,N_4432,N_4826);
xnor U7973 (N_7973,N_3235,N_3579);
nor U7974 (N_7974,N_5981,N_4289);
nor U7975 (N_7975,N_3791,N_5379);
nor U7976 (N_7976,N_5934,N_3163);
nand U7977 (N_7977,N_3920,N_4383);
nand U7978 (N_7978,N_3716,N_4753);
and U7979 (N_7979,N_5720,N_5001);
or U7980 (N_7980,N_3316,N_3369);
nand U7981 (N_7981,N_3420,N_4242);
and U7982 (N_7982,N_3666,N_4654);
nor U7983 (N_7983,N_6058,N_4929);
xor U7984 (N_7984,N_3691,N_4483);
and U7985 (N_7985,N_5488,N_4135);
nor U7986 (N_7986,N_5032,N_5925);
xnor U7987 (N_7987,N_5163,N_4794);
nand U7988 (N_7988,N_4657,N_4960);
nor U7989 (N_7989,N_3396,N_4497);
nand U7990 (N_7990,N_3563,N_5318);
nor U7991 (N_7991,N_6081,N_4265);
xor U7992 (N_7992,N_6059,N_4957);
nand U7993 (N_7993,N_5214,N_4082);
xnor U7994 (N_7994,N_5509,N_6175);
or U7995 (N_7995,N_3367,N_5002);
xnor U7996 (N_7996,N_5458,N_5030);
and U7997 (N_7997,N_6221,N_5524);
xnor U7998 (N_7998,N_4420,N_5560);
nor U7999 (N_7999,N_4596,N_4801);
nor U8000 (N_8000,N_3347,N_4634);
or U8001 (N_8001,N_5756,N_5316);
nor U8002 (N_8002,N_5513,N_3707);
or U8003 (N_8003,N_4447,N_6164);
and U8004 (N_8004,N_5345,N_5149);
and U8005 (N_8005,N_3639,N_3759);
xnor U8006 (N_8006,N_4372,N_5548);
or U8007 (N_8007,N_3765,N_3645);
and U8008 (N_8008,N_4476,N_3527);
xor U8009 (N_8009,N_3964,N_3394);
and U8010 (N_8010,N_5823,N_4985);
nand U8011 (N_8011,N_5618,N_6185);
xnor U8012 (N_8012,N_4444,N_5596);
xnor U8013 (N_8013,N_4097,N_3893);
nor U8014 (N_8014,N_6109,N_3315);
nor U8015 (N_8015,N_3223,N_4065);
and U8016 (N_8016,N_5712,N_3691);
nand U8017 (N_8017,N_5540,N_3685);
nor U8018 (N_8018,N_6187,N_3529);
xnor U8019 (N_8019,N_5499,N_4094);
xor U8020 (N_8020,N_6223,N_4507);
and U8021 (N_8021,N_3290,N_6098);
nor U8022 (N_8022,N_3151,N_3292);
and U8023 (N_8023,N_5078,N_4101);
and U8024 (N_8024,N_5278,N_3844);
and U8025 (N_8025,N_3856,N_4471);
and U8026 (N_8026,N_4811,N_3271);
xor U8027 (N_8027,N_4052,N_3241);
and U8028 (N_8028,N_4003,N_5088);
and U8029 (N_8029,N_4549,N_5476);
nor U8030 (N_8030,N_5135,N_5641);
nand U8031 (N_8031,N_5187,N_5262);
or U8032 (N_8032,N_5166,N_6169);
nand U8033 (N_8033,N_4374,N_3943);
and U8034 (N_8034,N_6238,N_6038);
xnor U8035 (N_8035,N_4355,N_6246);
and U8036 (N_8036,N_4035,N_5470);
nor U8037 (N_8037,N_4045,N_5582);
or U8038 (N_8038,N_3883,N_4560);
or U8039 (N_8039,N_5026,N_3390);
nand U8040 (N_8040,N_5359,N_5592);
nand U8041 (N_8041,N_3812,N_5803);
or U8042 (N_8042,N_5059,N_6218);
or U8043 (N_8043,N_3138,N_6120);
or U8044 (N_8044,N_4277,N_5031);
and U8045 (N_8045,N_5833,N_4321);
or U8046 (N_8046,N_5397,N_3134);
and U8047 (N_8047,N_5556,N_6139);
or U8048 (N_8048,N_4927,N_6096);
nand U8049 (N_8049,N_3920,N_6102);
and U8050 (N_8050,N_4176,N_4787);
xnor U8051 (N_8051,N_3720,N_6121);
and U8052 (N_8052,N_3306,N_5016);
and U8053 (N_8053,N_6073,N_5886);
and U8054 (N_8054,N_4361,N_5244);
nor U8055 (N_8055,N_4907,N_3674);
or U8056 (N_8056,N_6108,N_4906);
and U8057 (N_8057,N_4491,N_3396);
nand U8058 (N_8058,N_3407,N_4271);
and U8059 (N_8059,N_3619,N_5412);
and U8060 (N_8060,N_4685,N_6144);
or U8061 (N_8061,N_4479,N_4077);
nand U8062 (N_8062,N_3707,N_3443);
xor U8063 (N_8063,N_4773,N_3585);
xor U8064 (N_8064,N_3889,N_5248);
xor U8065 (N_8065,N_5446,N_6031);
or U8066 (N_8066,N_5620,N_4814);
nor U8067 (N_8067,N_3245,N_3721);
nand U8068 (N_8068,N_5221,N_5674);
or U8069 (N_8069,N_3838,N_5263);
nand U8070 (N_8070,N_5546,N_4162);
nor U8071 (N_8071,N_4134,N_5817);
or U8072 (N_8072,N_3946,N_4755);
xor U8073 (N_8073,N_5689,N_3837);
xnor U8074 (N_8074,N_5630,N_3608);
or U8075 (N_8075,N_5961,N_5518);
and U8076 (N_8076,N_4067,N_6198);
xnor U8077 (N_8077,N_5190,N_5387);
nand U8078 (N_8078,N_3579,N_4352);
nand U8079 (N_8079,N_3147,N_6044);
nor U8080 (N_8080,N_5293,N_5163);
xnor U8081 (N_8081,N_4896,N_5080);
and U8082 (N_8082,N_4443,N_3963);
xnor U8083 (N_8083,N_5044,N_3793);
nand U8084 (N_8084,N_4734,N_6074);
xor U8085 (N_8085,N_4040,N_5133);
or U8086 (N_8086,N_5785,N_4596);
or U8087 (N_8087,N_3718,N_4399);
nand U8088 (N_8088,N_5531,N_3299);
xnor U8089 (N_8089,N_5917,N_5808);
or U8090 (N_8090,N_5490,N_3909);
nand U8091 (N_8091,N_4493,N_3789);
xor U8092 (N_8092,N_6134,N_5958);
or U8093 (N_8093,N_6183,N_5074);
or U8094 (N_8094,N_3626,N_5021);
xnor U8095 (N_8095,N_4897,N_5424);
nor U8096 (N_8096,N_5998,N_3570);
nand U8097 (N_8097,N_5484,N_5137);
and U8098 (N_8098,N_4885,N_5384);
nand U8099 (N_8099,N_3279,N_5481);
nor U8100 (N_8100,N_3652,N_4582);
nor U8101 (N_8101,N_6007,N_6190);
and U8102 (N_8102,N_5529,N_5768);
nand U8103 (N_8103,N_6050,N_6232);
or U8104 (N_8104,N_4068,N_5943);
and U8105 (N_8105,N_5827,N_6051);
nand U8106 (N_8106,N_3904,N_4714);
and U8107 (N_8107,N_5916,N_3640);
and U8108 (N_8108,N_5540,N_3886);
nor U8109 (N_8109,N_3630,N_5053);
or U8110 (N_8110,N_5912,N_5669);
or U8111 (N_8111,N_4665,N_5074);
xor U8112 (N_8112,N_4380,N_4475);
nor U8113 (N_8113,N_5985,N_5458);
or U8114 (N_8114,N_3393,N_5074);
xnor U8115 (N_8115,N_3776,N_4099);
or U8116 (N_8116,N_4410,N_3164);
nand U8117 (N_8117,N_5478,N_5926);
nor U8118 (N_8118,N_3837,N_4221);
xnor U8119 (N_8119,N_6191,N_4061);
nor U8120 (N_8120,N_4030,N_5852);
nand U8121 (N_8121,N_3890,N_3634);
nor U8122 (N_8122,N_3739,N_3528);
or U8123 (N_8123,N_4655,N_4486);
nor U8124 (N_8124,N_4618,N_3598);
nor U8125 (N_8125,N_4555,N_3990);
and U8126 (N_8126,N_3948,N_4299);
xnor U8127 (N_8127,N_3658,N_5384);
xnor U8128 (N_8128,N_4658,N_4709);
nor U8129 (N_8129,N_5061,N_4901);
xor U8130 (N_8130,N_5466,N_4702);
and U8131 (N_8131,N_3426,N_5708);
nand U8132 (N_8132,N_5660,N_3991);
nor U8133 (N_8133,N_3628,N_5871);
xor U8134 (N_8134,N_5369,N_5891);
nor U8135 (N_8135,N_6158,N_4128);
or U8136 (N_8136,N_4872,N_5236);
xnor U8137 (N_8137,N_5178,N_4305);
or U8138 (N_8138,N_5445,N_5893);
or U8139 (N_8139,N_3755,N_4029);
and U8140 (N_8140,N_5229,N_3471);
nand U8141 (N_8141,N_5145,N_3296);
nand U8142 (N_8142,N_4663,N_3610);
nor U8143 (N_8143,N_4651,N_4600);
and U8144 (N_8144,N_3526,N_5205);
or U8145 (N_8145,N_6245,N_3632);
or U8146 (N_8146,N_5758,N_4674);
nor U8147 (N_8147,N_3863,N_5292);
nand U8148 (N_8148,N_6211,N_4475);
nand U8149 (N_8149,N_5669,N_4267);
and U8150 (N_8150,N_3205,N_5290);
nand U8151 (N_8151,N_3596,N_3627);
and U8152 (N_8152,N_6230,N_5894);
or U8153 (N_8153,N_4682,N_3770);
or U8154 (N_8154,N_4231,N_4072);
or U8155 (N_8155,N_6154,N_4935);
nand U8156 (N_8156,N_4003,N_3846);
or U8157 (N_8157,N_5398,N_6026);
xnor U8158 (N_8158,N_3588,N_5700);
xnor U8159 (N_8159,N_3873,N_4585);
nor U8160 (N_8160,N_4297,N_6103);
xnor U8161 (N_8161,N_6024,N_4531);
xnor U8162 (N_8162,N_4751,N_4753);
nor U8163 (N_8163,N_4090,N_6121);
and U8164 (N_8164,N_4241,N_3262);
nand U8165 (N_8165,N_5540,N_3513);
nand U8166 (N_8166,N_4642,N_6183);
and U8167 (N_8167,N_4926,N_3632);
or U8168 (N_8168,N_4129,N_4882);
xor U8169 (N_8169,N_5800,N_5252);
nor U8170 (N_8170,N_4529,N_5493);
or U8171 (N_8171,N_5995,N_6111);
nor U8172 (N_8172,N_5231,N_5841);
or U8173 (N_8173,N_3396,N_5611);
xnor U8174 (N_8174,N_4851,N_4321);
xor U8175 (N_8175,N_3693,N_5535);
nor U8176 (N_8176,N_4644,N_4303);
nor U8177 (N_8177,N_3451,N_4648);
nor U8178 (N_8178,N_3580,N_5267);
xnor U8179 (N_8179,N_5571,N_4751);
nor U8180 (N_8180,N_3537,N_5624);
and U8181 (N_8181,N_4401,N_4089);
xnor U8182 (N_8182,N_3854,N_3240);
or U8183 (N_8183,N_3541,N_4099);
nand U8184 (N_8184,N_4249,N_4630);
xnor U8185 (N_8185,N_5287,N_4374);
nor U8186 (N_8186,N_6179,N_4659);
and U8187 (N_8187,N_4350,N_3976);
nand U8188 (N_8188,N_4387,N_3968);
xor U8189 (N_8189,N_4854,N_4959);
xor U8190 (N_8190,N_4542,N_3437);
xnor U8191 (N_8191,N_5518,N_6071);
xnor U8192 (N_8192,N_4509,N_5791);
nand U8193 (N_8193,N_3147,N_4212);
and U8194 (N_8194,N_6162,N_4453);
or U8195 (N_8195,N_3369,N_5681);
nand U8196 (N_8196,N_3860,N_4087);
nand U8197 (N_8197,N_4514,N_3504);
and U8198 (N_8198,N_4063,N_4207);
or U8199 (N_8199,N_5044,N_4076);
xnor U8200 (N_8200,N_4048,N_5179);
or U8201 (N_8201,N_3659,N_5785);
nor U8202 (N_8202,N_5463,N_3230);
xnor U8203 (N_8203,N_5882,N_3435);
nor U8204 (N_8204,N_3977,N_4038);
or U8205 (N_8205,N_4785,N_4068);
or U8206 (N_8206,N_5260,N_4442);
xnor U8207 (N_8207,N_3367,N_3798);
nor U8208 (N_8208,N_4754,N_3405);
nor U8209 (N_8209,N_3485,N_4150);
and U8210 (N_8210,N_4995,N_5283);
nor U8211 (N_8211,N_6113,N_6084);
nor U8212 (N_8212,N_5899,N_5556);
or U8213 (N_8213,N_3734,N_5628);
or U8214 (N_8214,N_3721,N_5722);
nor U8215 (N_8215,N_3584,N_5267);
or U8216 (N_8216,N_3691,N_3278);
nand U8217 (N_8217,N_3812,N_3624);
xor U8218 (N_8218,N_4045,N_5291);
nor U8219 (N_8219,N_5523,N_4283);
nor U8220 (N_8220,N_5123,N_5379);
and U8221 (N_8221,N_3898,N_3478);
nor U8222 (N_8222,N_5498,N_4684);
or U8223 (N_8223,N_5909,N_3906);
nand U8224 (N_8224,N_4637,N_4289);
and U8225 (N_8225,N_5831,N_4145);
or U8226 (N_8226,N_5963,N_3738);
or U8227 (N_8227,N_3476,N_5030);
nand U8228 (N_8228,N_3769,N_5024);
or U8229 (N_8229,N_4784,N_6176);
nor U8230 (N_8230,N_3892,N_4125);
and U8231 (N_8231,N_4375,N_4312);
nor U8232 (N_8232,N_4161,N_3367);
nand U8233 (N_8233,N_3836,N_3849);
xor U8234 (N_8234,N_3686,N_5207);
xor U8235 (N_8235,N_5572,N_4652);
or U8236 (N_8236,N_5903,N_5941);
xor U8237 (N_8237,N_4133,N_4822);
xor U8238 (N_8238,N_4352,N_4672);
or U8239 (N_8239,N_3765,N_5200);
xor U8240 (N_8240,N_5032,N_5677);
nand U8241 (N_8241,N_3136,N_5743);
and U8242 (N_8242,N_5096,N_4176);
nand U8243 (N_8243,N_6118,N_3396);
or U8244 (N_8244,N_4362,N_5670);
nor U8245 (N_8245,N_4566,N_4616);
and U8246 (N_8246,N_4502,N_5934);
nor U8247 (N_8247,N_5037,N_5011);
or U8248 (N_8248,N_4525,N_5528);
nor U8249 (N_8249,N_5761,N_4579);
nor U8250 (N_8250,N_4558,N_6106);
and U8251 (N_8251,N_5865,N_4665);
xnor U8252 (N_8252,N_6186,N_4253);
and U8253 (N_8253,N_5469,N_6205);
or U8254 (N_8254,N_3810,N_5405);
nand U8255 (N_8255,N_4620,N_4870);
xnor U8256 (N_8256,N_5607,N_5007);
and U8257 (N_8257,N_4878,N_3445);
and U8258 (N_8258,N_4304,N_5391);
and U8259 (N_8259,N_3717,N_5061);
nand U8260 (N_8260,N_4223,N_4202);
nand U8261 (N_8261,N_5063,N_4322);
xor U8262 (N_8262,N_5659,N_4659);
nor U8263 (N_8263,N_4045,N_3879);
or U8264 (N_8264,N_4108,N_6140);
nand U8265 (N_8265,N_3303,N_5099);
or U8266 (N_8266,N_5601,N_4116);
nand U8267 (N_8267,N_3652,N_5504);
and U8268 (N_8268,N_5604,N_3178);
and U8269 (N_8269,N_4834,N_5513);
or U8270 (N_8270,N_5237,N_3505);
or U8271 (N_8271,N_3934,N_4733);
xor U8272 (N_8272,N_4331,N_4937);
nor U8273 (N_8273,N_3682,N_4738);
nand U8274 (N_8274,N_5702,N_5143);
or U8275 (N_8275,N_4482,N_4737);
xor U8276 (N_8276,N_5523,N_3199);
and U8277 (N_8277,N_5427,N_5309);
and U8278 (N_8278,N_3680,N_5471);
and U8279 (N_8279,N_6100,N_4125);
and U8280 (N_8280,N_5446,N_3783);
nand U8281 (N_8281,N_5923,N_5085);
nor U8282 (N_8282,N_3433,N_3753);
xor U8283 (N_8283,N_5738,N_3702);
and U8284 (N_8284,N_4351,N_4020);
nor U8285 (N_8285,N_3199,N_3487);
and U8286 (N_8286,N_5582,N_4133);
nand U8287 (N_8287,N_5204,N_6017);
xor U8288 (N_8288,N_3276,N_6130);
xor U8289 (N_8289,N_3887,N_4202);
and U8290 (N_8290,N_3475,N_4827);
xnor U8291 (N_8291,N_3786,N_3274);
and U8292 (N_8292,N_4809,N_4683);
and U8293 (N_8293,N_3727,N_5149);
nand U8294 (N_8294,N_4357,N_5434);
or U8295 (N_8295,N_3572,N_3217);
nor U8296 (N_8296,N_3268,N_5216);
nor U8297 (N_8297,N_4938,N_3349);
nor U8298 (N_8298,N_5773,N_5112);
xnor U8299 (N_8299,N_6146,N_3427);
and U8300 (N_8300,N_3864,N_5124);
nand U8301 (N_8301,N_4428,N_3906);
xor U8302 (N_8302,N_4094,N_5136);
nor U8303 (N_8303,N_6178,N_4453);
or U8304 (N_8304,N_4064,N_4198);
nor U8305 (N_8305,N_4756,N_4155);
nor U8306 (N_8306,N_4801,N_3615);
nand U8307 (N_8307,N_5381,N_3249);
nor U8308 (N_8308,N_4320,N_4007);
and U8309 (N_8309,N_3800,N_5656);
nand U8310 (N_8310,N_5818,N_3266);
nor U8311 (N_8311,N_4325,N_3443);
xnor U8312 (N_8312,N_3514,N_5065);
nand U8313 (N_8313,N_6032,N_5767);
and U8314 (N_8314,N_4424,N_6133);
xnor U8315 (N_8315,N_3308,N_3160);
and U8316 (N_8316,N_4940,N_5839);
xnor U8317 (N_8317,N_5711,N_5692);
nand U8318 (N_8318,N_5897,N_5605);
nand U8319 (N_8319,N_4954,N_5146);
nor U8320 (N_8320,N_4152,N_4879);
xor U8321 (N_8321,N_4965,N_3796);
nand U8322 (N_8322,N_3780,N_6142);
nand U8323 (N_8323,N_5900,N_3384);
nor U8324 (N_8324,N_4799,N_4853);
or U8325 (N_8325,N_6111,N_5111);
nand U8326 (N_8326,N_4193,N_4273);
nor U8327 (N_8327,N_3504,N_4209);
xor U8328 (N_8328,N_5825,N_5944);
nand U8329 (N_8329,N_3607,N_4492);
nand U8330 (N_8330,N_5282,N_3607);
and U8331 (N_8331,N_6246,N_5849);
xor U8332 (N_8332,N_5919,N_5560);
xnor U8333 (N_8333,N_3743,N_4621);
nand U8334 (N_8334,N_5970,N_5468);
xnor U8335 (N_8335,N_3453,N_3180);
or U8336 (N_8336,N_4504,N_4457);
and U8337 (N_8337,N_3134,N_5054);
or U8338 (N_8338,N_4296,N_4643);
nor U8339 (N_8339,N_4091,N_4002);
nor U8340 (N_8340,N_4655,N_3689);
xor U8341 (N_8341,N_5928,N_5729);
and U8342 (N_8342,N_5395,N_3913);
xor U8343 (N_8343,N_4203,N_4323);
and U8344 (N_8344,N_5565,N_5324);
nor U8345 (N_8345,N_3401,N_4069);
xnor U8346 (N_8346,N_5015,N_4951);
xnor U8347 (N_8347,N_4432,N_4767);
xor U8348 (N_8348,N_3699,N_4414);
nand U8349 (N_8349,N_5078,N_3292);
nor U8350 (N_8350,N_6003,N_4268);
and U8351 (N_8351,N_3216,N_3401);
nor U8352 (N_8352,N_6103,N_3340);
or U8353 (N_8353,N_5443,N_4299);
xnor U8354 (N_8354,N_5613,N_3802);
nor U8355 (N_8355,N_3566,N_5081);
xnor U8356 (N_8356,N_5003,N_5132);
or U8357 (N_8357,N_6228,N_5848);
nor U8358 (N_8358,N_4068,N_4783);
nor U8359 (N_8359,N_4081,N_3556);
xor U8360 (N_8360,N_5621,N_5332);
nor U8361 (N_8361,N_4471,N_5885);
nand U8362 (N_8362,N_3967,N_5678);
xor U8363 (N_8363,N_4968,N_4362);
nor U8364 (N_8364,N_3183,N_6194);
nand U8365 (N_8365,N_5372,N_4216);
nor U8366 (N_8366,N_3836,N_5691);
and U8367 (N_8367,N_4667,N_4712);
xnor U8368 (N_8368,N_4045,N_5458);
nand U8369 (N_8369,N_3488,N_3922);
nand U8370 (N_8370,N_5786,N_5591);
nor U8371 (N_8371,N_3137,N_3589);
or U8372 (N_8372,N_5986,N_5574);
xnor U8373 (N_8373,N_5418,N_4001);
and U8374 (N_8374,N_5165,N_5440);
nand U8375 (N_8375,N_4620,N_5103);
xnor U8376 (N_8376,N_5747,N_4533);
nor U8377 (N_8377,N_3379,N_5538);
nor U8378 (N_8378,N_5481,N_4910);
nor U8379 (N_8379,N_3607,N_3224);
xnor U8380 (N_8380,N_5777,N_3770);
or U8381 (N_8381,N_4042,N_4473);
nor U8382 (N_8382,N_4475,N_5503);
nand U8383 (N_8383,N_6046,N_3408);
nor U8384 (N_8384,N_5802,N_3879);
nor U8385 (N_8385,N_4898,N_5007);
xnor U8386 (N_8386,N_3555,N_6223);
xor U8387 (N_8387,N_5535,N_5667);
xor U8388 (N_8388,N_3853,N_4561);
nor U8389 (N_8389,N_5301,N_5954);
or U8390 (N_8390,N_5979,N_4777);
nor U8391 (N_8391,N_3155,N_3726);
nor U8392 (N_8392,N_4646,N_3664);
xor U8393 (N_8393,N_4389,N_3967);
and U8394 (N_8394,N_3132,N_4411);
or U8395 (N_8395,N_5369,N_5446);
nor U8396 (N_8396,N_4068,N_3799);
and U8397 (N_8397,N_3526,N_5576);
nor U8398 (N_8398,N_5600,N_5258);
nand U8399 (N_8399,N_5181,N_5470);
nor U8400 (N_8400,N_4140,N_3353);
and U8401 (N_8401,N_5557,N_6008);
or U8402 (N_8402,N_4828,N_4476);
or U8403 (N_8403,N_5398,N_5656);
or U8404 (N_8404,N_4711,N_4691);
nand U8405 (N_8405,N_3602,N_3944);
xnor U8406 (N_8406,N_5784,N_5037);
and U8407 (N_8407,N_6037,N_3648);
xnor U8408 (N_8408,N_5294,N_3715);
nand U8409 (N_8409,N_3728,N_4867);
and U8410 (N_8410,N_4674,N_3868);
and U8411 (N_8411,N_4190,N_5715);
nor U8412 (N_8412,N_5343,N_4443);
nor U8413 (N_8413,N_5949,N_4528);
or U8414 (N_8414,N_5189,N_5468);
xnor U8415 (N_8415,N_4737,N_5770);
nor U8416 (N_8416,N_4310,N_4163);
or U8417 (N_8417,N_3981,N_4344);
and U8418 (N_8418,N_4989,N_3702);
nor U8419 (N_8419,N_3567,N_5480);
or U8420 (N_8420,N_6112,N_5286);
xor U8421 (N_8421,N_6223,N_5444);
xnor U8422 (N_8422,N_5437,N_3669);
or U8423 (N_8423,N_5175,N_3125);
nand U8424 (N_8424,N_5576,N_3918);
nand U8425 (N_8425,N_5139,N_4007);
or U8426 (N_8426,N_4750,N_4470);
or U8427 (N_8427,N_4060,N_3983);
nor U8428 (N_8428,N_4572,N_4674);
or U8429 (N_8429,N_3578,N_5258);
nor U8430 (N_8430,N_4010,N_3645);
and U8431 (N_8431,N_5834,N_3716);
xnor U8432 (N_8432,N_5492,N_4746);
xor U8433 (N_8433,N_5749,N_4888);
nor U8434 (N_8434,N_5203,N_5674);
nand U8435 (N_8435,N_5732,N_3135);
nand U8436 (N_8436,N_4757,N_5424);
nor U8437 (N_8437,N_5620,N_3188);
nand U8438 (N_8438,N_3380,N_3459);
or U8439 (N_8439,N_4190,N_3591);
or U8440 (N_8440,N_5733,N_3863);
nor U8441 (N_8441,N_4967,N_5594);
nor U8442 (N_8442,N_3300,N_4141);
nand U8443 (N_8443,N_4644,N_3702);
or U8444 (N_8444,N_3304,N_5086);
nor U8445 (N_8445,N_3986,N_3740);
or U8446 (N_8446,N_4871,N_5598);
and U8447 (N_8447,N_5430,N_3527);
nand U8448 (N_8448,N_3598,N_3600);
nand U8449 (N_8449,N_5115,N_6024);
nand U8450 (N_8450,N_6208,N_3427);
xnor U8451 (N_8451,N_4661,N_4651);
nand U8452 (N_8452,N_4800,N_5258);
or U8453 (N_8453,N_5121,N_4734);
nor U8454 (N_8454,N_4231,N_5480);
or U8455 (N_8455,N_3235,N_4762);
and U8456 (N_8456,N_4290,N_5749);
or U8457 (N_8457,N_5190,N_4415);
and U8458 (N_8458,N_5777,N_5357);
xnor U8459 (N_8459,N_5083,N_5014);
or U8460 (N_8460,N_5131,N_5096);
xnor U8461 (N_8461,N_5453,N_3229);
or U8462 (N_8462,N_5560,N_3662);
xor U8463 (N_8463,N_3627,N_5278);
xnor U8464 (N_8464,N_5451,N_4224);
nor U8465 (N_8465,N_5905,N_4325);
and U8466 (N_8466,N_5583,N_3763);
or U8467 (N_8467,N_6055,N_3622);
nand U8468 (N_8468,N_5743,N_5231);
or U8469 (N_8469,N_4793,N_4728);
xor U8470 (N_8470,N_3625,N_3593);
nor U8471 (N_8471,N_3733,N_4676);
or U8472 (N_8472,N_5205,N_5980);
and U8473 (N_8473,N_5179,N_3611);
nand U8474 (N_8474,N_3370,N_4079);
and U8475 (N_8475,N_4178,N_6083);
nor U8476 (N_8476,N_5304,N_4819);
nor U8477 (N_8477,N_3529,N_6121);
nand U8478 (N_8478,N_4820,N_4718);
nand U8479 (N_8479,N_4515,N_4251);
or U8480 (N_8480,N_3260,N_4385);
nand U8481 (N_8481,N_3700,N_5465);
or U8482 (N_8482,N_4143,N_4946);
nor U8483 (N_8483,N_3321,N_3203);
xnor U8484 (N_8484,N_3939,N_4893);
nand U8485 (N_8485,N_4039,N_5167);
and U8486 (N_8486,N_3355,N_4359);
xor U8487 (N_8487,N_4205,N_3677);
nor U8488 (N_8488,N_4239,N_3219);
or U8489 (N_8489,N_4287,N_5478);
nor U8490 (N_8490,N_5241,N_4645);
or U8491 (N_8491,N_4034,N_5794);
or U8492 (N_8492,N_3393,N_4163);
and U8493 (N_8493,N_3215,N_6174);
or U8494 (N_8494,N_4247,N_4951);
nor U8495 (N_8495,N_5034,N_3766);
and U8496 (N_8496,N_5688,N_4248);
nor U8497 (N_8497,N_4571,N_4906);
xor U8498 (N_8498,N_4482,N_4211);
and U8499 (N_8499,N_4657,N_4168);
nand U8500 (N_8500,N_3905,N_3645);
or U8501 (N_8501,N_4990,N_5643);
xor U8502 (N_8502,N_4201,N_3214);
or U8503 (N_8503,N_5404,N_4952);
nor U8504 (N_8504,N_4058,N_4789);
and U8505 (N_8505,N_3139,N_5134);
xnor U8506 (N_8506,N_4658,N_4366);
nand U8507 (N_8507,N_4451,N_5242);
nand U8508 (N_8508,N_4417,N_4494);
or U8509 (N_8509,N_3854,N_5153);
nor U8510 (N_8510,N_3976,N_5813);
nor U8511 (N_8511,N_4371,N_4093);
nand U8512 (N_8512,N_5986,N_3887);
nand U8513 (N_8513,N_5395,N_6172);
nor U8514 (N_8514,N_4702,N_5690);
nand U8515 (N_8515,N_5638,N_4426);
nand U8516 (N_8516,N_5786,N_5247);
and U8517 (N_8517,N_5040,N_3790);
nor U8518 (N_8518,N_5524,N_5038);
nand U8519 (N_8519,N_5317,N_5660);
xnor U8520 (N_8520,N_5715,N_5068);
xor U8521 (N_8521,N_5142,N_5918);
and U8522 (N_8522,N_3245,N_4666);
and U8523 (N_8523,N_6059,N_5859);
nor U8524 (N_8524,N_5421,N_3667);
xnor U8525 (N_8525,N_3429,N_6170);
and U8526 (N_8526,N_5657,N_3513);
nand U8527 (N_8527,N_4796,N_3949);
xor U8528 (N_8528,N_3401,N_5932);
nand U8529 (N_8529,N_4727,N_4773);
and U8530 (N_8530,N_3615,N_3491);
or U8531 (N_8531,N_6100,N_4108);
and U8532 (N_8532,N_4768,N_4573);
and U8533 (N_8533,N_5729,N_5809);
nor U8534 (N_8534,N_3926,N_4253);
xnor U8535 (N_8535,N_5923,N_5115);
and U8536 (N_8536,N_6171,N_5709);
nor U8537 (N_8537,N_3296,N_5031);
nand U8538 (N_8538,N_5471,N_5117);
nor U8539 (N_8539,N_5739,N_3665);
or U8540 (N_8540,N_4439,N_5519);
and U8541 (N_8541,N_5059,N_3730);
xor U8542 (N_8542,N_3964,N_5159);
xnor U8543 (N_8543,N_4538,N_3501);
or U8544 (N_8544,N_4937,N_6245);
xor U8545 (N_8545,N_5125,N_5158);
and U8546 (N_8546,N_5348,N_4016);
xnor U8547 (N_8547,N_3143,N_3469);
or U8548 (N_8548,N_3175,N_5233);
xor U8549 (N_8549,N_4313,N_4429);
nor U8550 (N_8550,N_5519,N_6181);
or U8551 (N_8551,N_5253,N_6220);
xnor U8552 (N_8552,N_4597,N_4809);
xnor U8553 (N_8553,N_3201,N_3654);
xor U8554 (N_8554,N_5988,N_5592);
or U8555 (N_8555,N_5139,N_3425);
xor U8556 (N_8556,N_3676,N_4684);
nor U8557 (N_8557,N_3184,N_6245);
and U8558 (N_8558,N_6029,N_4304);
nor U8559 (N_8559,N_6183,N_5492);
nor U8560 (N_8560,N_3329,N_3343);
nand U8561 (N_8561,N_3277,N_4131);
nor U8562 (N_8562,N_4570,N_5629);
nand U8563 (N_8563,N_5635,N_5394);
and U8564 (N_8564,N_5526,N_4849);
and U8565 (N_8565,N_5392,N_6210);
or U8566 (N_8566,N_4728,N_4253);
xor U8567 (N_8567,N_3554,N_5415);
xor U8568 (N_8568,N_3308,N_4067);
or U8569 (N_8569,N_6176,N_5559);
nand U8570 (N_8570,N_4587,N_4963);
and U8571 (N_8571,N_4666,N_3291);
and U8572 (N_8572,N_5872,N_3295);
nor U8573 (N_8573,N_5025,N_4518);
or U8574 (N_8574,N_3776,N_5387);
and U8575 (N_8575,N_3660,N_5684);
nor U8576 (N_8576,N_3507,N_5936);
or U8577 (N_8577,N_3197,N_5036);
nand U8578 (N_8578,N_4117,N_4391);
xor U8579 (N_8579,N_3165,N_5136);
and U8580 (N_8580,N_3896,N_6083);
nor U8581 (N_8581,N_5022,N_3425);
xor U8582 (N_8582,N_6078,N_4096);
nor U8583 (N_8583,N_5958,N_4884);
nand U8584 (N_8584,N_3135,N_5663);
and U8585 (N_8585,N_3681,N_4452);
nand U8586 (N_8586,N_5750,N_5121);
xnor U8587 (N_8587,N_4151,N_5423);
or U8588 (N_8588,N_6216,N_4588);
nor U8589 (N_8589,N_5957,N_3375);
xor U8590 (N_8590,N_3782,N_4335);
or U8591 (N_8591,N_3229,N_4078);
or U8592 (N_8592,N_4558,N_5226);
xnor U8593 (N_8593,N_3320,N_3862);
nor U8594 (N_8594,N_5895,N_5692);
or U8595 (N_8595,N_5415,N_4538);
xnor U8596 (N_8596,N_5703,N_4509);
and U8597 (N_8597,N_4037,N_5908);
nand U8598 (N_8598,N_4083,N_4506);
nand U8599 (N_8599,N_5165,N_4648);
nand U8600 (N_8600,N_4372,N_6001);
and U8601 (N_8601,N_4834,N_6230);
and U8602 (N_8602,N_4070,N_6094);
nand U8603 (N_8603,N_4570,N_5059);
and U8604 (N_8604,N_3815,N_4813);
nand U8605 (N_8605,N_5985,N_4575);
nor U8606 (N_8606,N_6081,N_5953);
and U8607 (N_8607,N_3924,N_3230);
and U8608 (N_8608,N_4976,N_4759);
nor U8609 (N_8609,N_3459,N_5608);
nand U8610 (N_8610,N_4506,N_4627);
xnor U8611 (N_8611,N_4164,N_5474);
and U8612 (N_8612,N_4421,N_5203);
and U8613 (N_8613,N_5078,N_4618);
or U8614 (N_8614,N_5374,N_3167);
nand U8615 (N_8615,N_4702,N_3173);
nand U8616 (N_8616,N_3691,N_5521);
nand U8617 (N_8617,N_4846,N_5834);
xnor U8618 (N_8618,N_4871,N_3625);
nor U8619 (N_8619,N_3753,N_6091);
xnor U8620 (N_8620,N_5853,N_3621);
or U8621 (N_8621,N_4975,N_5886);
xor U8622 (N_8622,N_4294,N_4064);
or U8623 (N_8623,N_4030,N_3227);
nand U8624 (N_8624,N_4711,N_6196);
nor U8625 (N_8625,N_5040,N_5786);
or U8626 (N_8626,N_6082,N_4020);
and U8627 (N_8627,N_4154,N_6106);
nor U8628 (N_8628,N_4065,N_3800);
xnor U8629 (N_8629,N_3979,N_4760);
nand U8630 (N_8630,N_6163,N_4116);
or U8631 (N_8631,N_3317,N_4925);
nand U8632 (N_8632,N_3678,N_5397);
xnor U8633 (N_8633,N_3495,N_4361);
and U8634 (N_8634,N_4343,N_5438);
and U8635 (N_8635,N_4303,N_4131);
nor U8636 (N_8636,N_3632,N_3975);
and U8637 (N_8637,N_4734,N_6094);
and U8638 (N_8638,N_3597,N_3838);
nand U8639 (N_8639,N_3446,N_5604);
xnor U8640 (N_8640,N_6012,N_5858);
or U8641 (N_8641,N_3711,N_6153);
xnor U8642 (N_8642,N_4559,N_5082);
xnor U8643 (N_8643,N_5886,N_4052);
or U8644 (N_8644,N_5549,N_4877);
or U8645 (N_8645,N_3855,N_5824);
or U8646 (N_8646,N_5332,N_5859);
and U8647 (N_8647,N_4354,N_3303);
and U8648 (N_8648,N_4155,N_4731);
nor U8649 (N_8649,N_4231,N_4094);
xnor U8650 (N_8650,N_3428,N_3759);
and U8651 (N_8651,N_4825,N_6243);
or U8652 (N_8652,N_5773,N_3251);
nor U8653 (N_8653,N_5450,N_3676);
nor U8654 (N_8654,N_5619,N_4796);
or U8655 (N_8655,N_3725,N_5949);
nand U8656 (N_8656,N_5853,N_3495);
and U8657 (N_8657,N_3356,N_5504);
or U8658 (N_8658,N_4669,N_4841);
nor U8659 (N_8659,N_5498,N_4174);
nor U8660 (N_8660,N_5266,N_3724);
nor U8661 (N_8661,N_5466,N_4954);
xor U8662 (N_8662,N_4342,N_3172);
xor U8663 (N_8663,N_5660,N_4258);
or U8664 (N_8664,N_5385,N_5912);
nor U8665 (N_8665,N_3577,N_5017);
and U8666 (N_8666,N_3565,N_5460);
and U8667 (N_8667,N_4425,N_3641);
or U8668 (N_8668,N_3333,N_3518);
nor U8669 (N_8669,N_5576,N_6112);
nor U8670 (N_8670,N_5590,N_6111);
and U8671 (N_8671,N_4622,N_5268);
nand U8672 (N_8672,N_3283,N_5736);
nand U8673 (N_8673,N_4543,N_5472);
and U8674 (N_8674,N_4393,N_6020);
xnor U8675 (N_8675,N_5585,N_5318);
xor U8676 (N_8676,N_5589,N_5637);
nor U8677 (N_8677,N_4048,N_3398);
nor U8678 (N_8678,N_5875,N_4257);
nand U8679 (N_8679,N_4366,N_4200);
or U8680 (N_8680,N_5027,N_3548);
xnor U8681 (N_8681,N_3457,N_5966);
and U8682 (N_8682,N_3837,N_3411);
nor U8683 (N_8683,N_5908,N_6233);
xor U8684 (N_8684,N_3734,N_5809);
or U8685 (N_8685,N_4403,N_4593);
nand U8686 (N_8686,N_5936,N_4481);
nand U8687 (N_8687,N_5604,N_4508);
nor U8688 (N_8688,N_4944,N_4378);
or U8689 (N_8689,N_3186,N_5808);
or U8690 (N_8690,N_3558,N_3593);
nor U8691 (N_8691,N_6038,N_4885);
xnor U8692 (N_8692,N_4697,N_4535);
or U8693 (N_8693,N_3143,N_3657);
nand U8694 (N_8694,N_4311,N_4799);
xor U8695 (N_8695,N_3920,N_4609);
nand U8696 (N_8696,N_5860,N_3711);
nor U8697 (N_8697,N_4064,N_4997);
xor U8698 (N_8698,N_3665,N_4373);
or U8699 (N_8699,N_4264,N_3156);
or U8700 (N_8700,N_4893,N_4549);
xnor U8701 (N_8701,N_4634,N_4378);
nor U8702 (N_8702,N_4883,N_4585);
nor U8703 (N_8703,N_4994,N_3783);
xor U8704 (N_8704,N_3220,N_4340);
or U8705 (N_8705,N_3175,N_5064);
and U8706 (N_8706,N_5190,N_3270);
or U8707 (N_8707,N_3204,N_6195);
nand U8708 (N_8708,N_5267,N_4421);
or U8709 (N_8709,N_4668,N_4744);
nand U8710 (N_8710,N_5555,N_3824);
xor U8711 (N_8711,N_4451,N_4911);
or U8712 (N_8712,N_3585,N_4532);
and U8713 (N_8713,N_6008,N_3153);
nor U8714 (N_8714,N_4440,N_3508);
nand U8715 (N_8715,N_6053,N_4885);
nor U8716 (N_8716,N_5556,N_5834);
nand U8717 (N_8717,N_4164,N_3790);
and U8718 (N_8718,N_4187,N_5835);
xor U8719 (N_8719,N_3871,N_3154);
or U8720 (N_8720,N_4667,N_5561);
nand U8721 (N_8721,N_5970,N_5844);
or U8722 (N_8722,N_4038,N_4074);
and U8723 (N_8723,N_5139,N_6242);
and U8724 (N_8724,N_4549,N_4586);
xor U8725 (N_8725,N_5997,N_3994);
or U8726 (N_8726,N_4429,N_3401);
and U8727 (N_8727,N_4195,N_3722);
or U8728 (N_8728,N_3465,N_4849);
xnor U8729 (N_8729,N_5623,N_5337);
nand U8730 (N_8730,N_5554,N_3979);
and U8731 (N_8731,N_3372,N_4082);
or U8732 (N_8732,N_3902,N_4200);
and U8733 (N_8733,N_5943,N_3546);
or U8734 (N_8734,N_3354,N_3422);
or U8735 (N_8735,N_3226,N_3130);
nand U8736 (N_8736,N_4020,N_4015);
and U8737 (N_8737,N_6241,N_5464);
xor U8738 (N_8738,N_4557,N_3465);
and U8739 (N_8739,N_4525,N_6021);
and U8740 (N_8740,N_5617,N_5968);
nor U8741 (N_8741,N_5117,N_3862);
nor U8742 (N_8742,N_3513,N_5677);
nand U8743 (N_8743,N_3772,N_3665);
nand U8744 (N_8744,N_4533,N_5609);
or U8745 (N_8745,N_3244,N_5671);
xor U8746 (N_8746,N_3226,N_3910);
nand U8747 (N_8747,N_4026,N_4265);
nor U8748 (N_8748,N_4924,N_5658);
or U8749 (N_8749,N_3305,N_3663);
xor U8750 (N_8750,N_4481,N_6247);
and U8751 (N_8751,N_4567,N_4534);
and U8752 (N_8752,N_4329,N_4807);
nor U8753 (N_8753,N_5151,N_6192);
nand U8754 (N_8754,N_5435,N_5414);
or U8755 (N_8755,N_4410,N_3222);
xnor U8756 (N_8756,N_6065,N_3535);
or U8757 (N_8757,N_3759,N_6039);
and U8758 (N_8758,N_5946,N_6133);
and U8759 (N_8759,N_3718,N_6228);
and U8760 (N_8760,N_3586,N_4485);
nor U8761 (N_8761,N_3739,N_3296);
xor U8762 (N_8762,N_3656,N_3126);
nand U8763 (N_8763,N_5260,N_6150);
and U8764 (N_8764,N_6102,N_3907);
and U8765 (N_8765,N_3586,N_3901);
or U8766 (N_8766,N_3301,N_3606);
and U8767 (N_8767,N_5008,N_5134);
nor U8768 (N_8768,N_5799,N_4285);
nor U8769 (N_8769,N_4371,N_3754);
and U8770 (N_8770,N_5281,N_5105);
and U8771 (N_8771,N_3274,N_4488);
or U8772 (N_8772,N_6064,N_4390);
or U8773 (N_8773,N_4322,N_5736);
nand U8774 (N_8774,N_5651,N_5232);
xnor U8775 (N_8775,N_3600,N_3270);
xor U8776 (N_8776,N_4949,N_5292);
xor U8777 (N_8777,N_5821,N_5652);
nor U8778 (N_8778,N_4271,N_3966);
nand U8779 (N_8779,N_3259,N_3960);
and U8780 (N_8780,N_4978,N_5391);
and U8781 (N_8781,N_5754,N_5573);
nor U8782 (N_8782,N_4243,N_4752);
nand U8783 (N_8783,N_4880,N_5524);
and U8784 (N_8784,N_4446,N_5167);
and U8785 (N_8785,N_3839,N_4531);
or U8786 (N_8786,N_3952,N_3460);
xor U8787 (N_8787,N_4778,N_4164);
and U8788 (N_8788,N_4751,N_6196);
nand U8789 (N_8789,N_3413,N_5704);
and U8790 (N_8790,N_4654,N_5309);
or U8791 (N_8791,N_5510,N_5418);
nand U8792 (N_8792,N_3257,N_3403);
nor U8793 (N_8793,N_3588,N_4981);
nor U8794 (N_8794,N_3722,N_4705);
or U8795 (N_8795,N_4799,N_5222);
nor U8796 (N_8796,N_5385,N_4360);
and U8797 (N_8797,N_3790,N_4239);
nor U8798 (N_8798,N_3724,N_5155);
and U8799 (N_8799,N_5930,N_5875);
xor U8800 (N_8800,N_6207,N_4198);
xor U8801 (N_8801,N_4613,N_5412);
nand U8802 (N_8802,N_5690,N_5391);
xor U8803 (N_8803,N_3495,N_5676);
or U8804 (N_8804,N_3586,N_5368);
nor U8805 (N_8805,N_3412,N_3341);
and U8806 (N_8806,N_5947,N_5494);
nand U8807 (N_8807,N_5176,N_3815);
and U8808 (N_8808,N_4198,N_4230);
nand U8809 (N_8809,N_3158,N_4254);
xor U8810 (N_8810,N_4732,N_4978);
or U8811 (N_8811,N_5056,N_4813);
and U8812 (N_8812,N_3463,N_4646);
or U8813 (N_8813,N_5061,N_4339);
nand U8814 (N_8814,N_3807,N_3909);
and U8815 (N_8815,N_3223,N_5814);
xor U8816 (N_8816,N_3724,N_4207);
or U8817 (N_8817,N_5561,N_6082);
xor U8818 (N_8818,N_3479,N_5723);
nand U8819 (N_8819,N_5206,N_3919);
nand U8820 (N_8820,N_3153,N_4420);
xor U8821 (N_8821,N_5804,N_5642);
xor U8822 (N_8822,N_4950,N_3173);
or U8823 (N_8823,N_4277,N_3853);
xor U8824 (N_8824,N_4996,N_3554);
nor U8825 (N_8825,N_4295,N_4344);
nor U8826 (N_8826,N_4636,N_5249);
xnor U8827 (N_8827,N_5154,N_6246);
xnor U8828 (N_8828,N_5203,N_5164);
and U8829 (N_8829,N_5811,N_4515);
nand U8830 (N_8830,N_5129,N_5544);
and U8831 (N_8831,N_6132,N_3598);
nand U8832 (N_8832,N_5461,N_4390);
or U8833 (N_8833,N_4049,N_4951);
nand U8834 (N_8834,N_4574,N_5620);
nor U8835 (N_8835,N_3909,N_3509);
and U8836 (N_8836,N_4358,N_6228);
nor U8837 (N_8837,N_4690,N_5558);
nor U8838 (N_8838,N_5131,N_5209);
and U8839 (N_8839,N_4484,N_4231);
xor U8840 (N_8840,N_3414,N_5012);
and U8841 (N_8841,N_3817,N_4998);
or U8842 (N_8842,N_5489,N_4661);
nor U8843 (N_8843,N_5198,N_5807);
and U8844 (N_8844,N_5391,N_5483);
or U8845 (N_8845,N_6011,N_3755);
nand U8846 (N_8846,N_6245,N_5922);
nor U8847 (N_8847,N_4842,N_5939);
xor U8848 (N_8848,N_3837,N_4589);
and U8849 (N_8849,N_4624,N_4753);
xnor U8850 (N_8850,N_5312,N_3881);
nand U8851 (N_8851,N_6028,N_3551);
nor U8852 (N_8852,N_4122,N_5967);
or U8853 (N_8853,N_3773,N_3253);
or U8854 (N_8854,N_5883,N_4018);
or U8855 (N_8855,N_5494,N_5362);
and U8856 (N_8856,N_4514,N_3910);
and U8857 (N_8857,N_3166,N_3797);
or U8858 (N_8858,N_4098,N_4594);
and U8859 (N_8859,N_5420,N_3611);
nor U8860 (N_8860,N_4898,N_5019);
or U8861 (N_8861,N_6024,N_3198);
and U8862 (N_8862,N_6108,N_5387);
and U8863 (N_8863,N_3323,N_4113);
nand U8864 (N_8864,N_5142,N_3438);
xor U8865 (N_8865,N_5838,N_5030);
and U8866 (N_8866,N_3662,N_3845);
xnor U8867 (N_8867,N_4339,N_5645);
xor U8868 (N_8868,N_4654,N_3680);
and U8869 (N_8869,N_5325,N_5549);
nor U8870 (N_8870,N_5113,N_5267);
nand U8871 (N_8871,N_5666,N_5723);
xor U8872 (N_8872,N_5509,N_5943);
nand U8873 (N_8873,N_5973,N_3946);
xnor U8874 (N_8874,N_5302,N_5148);
or U8875 (N_8875,N_5537,N_5847);
nor U8876 (N_8876,N_3753,N_5982);
or U8877 (N_8877,N_5633,N_4913);
nand U8878 (N_8878,N_4866,N_3773);
or U8879 (N_8879,N_5043,N_4157);
nor U8880 (N_8880,N_6230,N_4915);
nor U8881 (N_8881,N_4812,N_4902);
xnor U8882 (N_8882,N_5490,N_4477);
and U8883 (N_8883,N_4739,N_4049);
xor U8884 (N_8884,N_5305,N_3587);
xor U8885 (N_8885,N_5769,N_5446);
nor U8886 (N_8886,N_3565,N_6224);
nor U8887 (N_8887,N_4098,N_6005);
nor U8888 (N_8888,N_4098,N_4179);
or U8889 (N_8889,N_3608,N_4314);
xnor U8890 (N_8890,N_5323,N_3590);
nand U8891 (N_8891,N_3858,N_5011);
xnor U8892 (N_8892,N_4483,N_3869);
nor U8893 (N_8893,N_4580,N_5197);
or U8894 (N_8894,N_4102,N_3960);
xnor U8895 (N_8895,N_6211,N_4169);
and U8896 (N_8896,N_3767,N_3787);
and U8897 (N_8897,N_3949,N_5443);
nand U8898 (N_8898,N_3771,N_3334);
or U8899 (N_8899,N_5440,N_5389);
xnor U8900 (N_8900,N_5742,N_5482);
and U8901 (N_8901,N_5530,N_5488);
xor U8902 (N_8902,N_3244,N_5718);
and U8903 (N_8903,N_4693,N_5406);
or U8904 (N_8904,N_3888,N_4624);
or U8905 (N_8905,N_5718,N_5219);
or U8906 (N_8906,N_4294,N_4184);
xnor U8907 (N_8907,N_3536,N_4307);
xnor U8908 (N_8908,N_5890,N_4571);
nor U8909 (N_8909,N_5641,N_3705);
nor U8910 (N_8910,N_6218,N_4797);
nor U8911 (N_8911,N_5181,N_5635);
nand U8912 (N_8912,N_3275,N_5442);
nor U8913 (N_8913,N_5913,N_5370);
nor U8914 (N_8914,N_4911,N_5770);
and U8915 (N_8915,N_3634,N_6214);
or U8916 (N_8916,N_3431,N_5725);
and U8917 (N_8917,N_3243,N_6119);
or U8918 (N_8918,N_5995,N_4671);
xor U8919 (N_8919,N_5418,N_3990);
and U8920 (N_8920,N_5732,N_3707);
xor U8921 (N_8921,N_3172,N_3635);
nor U8922 (N_8922,N_3372,N_3276);
xor U8923 (N_8923,N_4175,N_4086);
or U8924 (N_8924,N_3887,N_6120);
nor U8925 (N_8925,N_3156,N_5299);
xnor U8926 (N_8926,N_5986,N_4303);
or U8927 (N_8927,N_4521,N_6170);
and U8928 (N_8928,N_3888,N_3326);
nand U8929 (N_8929,N_4468,N_5494);
nor U8930 (N_8930,N_4687,N_4042);
and U8931 (N_8931,N_5083,N_4067);
xor U8932 (N_8932,N_5348,N_4106);
xnor U8933 (N_8933,N_5719,N_5127);
nand U8934 (N_8934,N_5153,N_6134);
nor U8935 (N_8935,N_3354,N_5493);
and U8936 (N_8936,N_3693,N_5591);
or U8937 (N_8937,N_5640,N_4699);
nor U8938 (N_8938,N_4229,N_3450);
nor U8939 (N_8939,N_4298,N_3225);
or U8940 (N_8940,N_5374,N_4568);
nor U8941 (N_8941,N_3908,N_5531);
nand U8942 (N_8942,N_4575,N_5308);
xnor U8943 (N_8943,N_3877,N_3322);
nor U8944 (N_8944,N_3656,N_6016);
and U8945 (N_8945,N_3376,N_6239);
and U8946 (N_8946,N_3645,N_4288);
or U8947 (N_8947,N_4887,N_4990);
nor U8948 (N_8948,N_5313,N_3576);
and U8949 (N_8949,N_3664,N_3267);
or U8950 (N_8950,N_3885,N_6111);
nor U8951 (N_8951,N_5754,N_3507);
or U8952 (N_8952,N_5570,N_5472);
and U8953 (N_8953,N_6092,N_5709);
nand U8954 (N_8954,N_3745,N_5060);
xnor U8955 (N_8955,N_4275,N_4442);
and U8956 (N_8956,N_5115,N_5898);
and U8957 (N_8957,N_5413,N_5273);
and U8958 (N_8958,N_4577,N_4405);
nand U8959 (N_8959,N_6225,N_5974);
xor U8960 (N_8960,N_4497,N_4644);
or U8961 (N_8961,N_3576,N_3612);
and U8962 (N_8962,N_4829,N_5063);
nand U8963 (N_8963,N_5383,N_6158);
and U8964 (N_8964,N_5548,N_5905);
xnor U8965 (N_8965,N_5365,N_3433);
or U8966 (N_8966,N_4777,N_5564);
xor U8967 (N_8967,N_4406,N_5980);
and U8968 (N_8968,N_3383,N_5274);
or U8969 (N_8969,N_5139,N_4110);
nand U8970 (N_8970,N_5801,N_5230);
nand U8971 (N_8971,N_4367,N_5585);
xnor U8972 (N_8972,N_4692,N_3561);
or U8973 (N_8973,N_4823,N_5617);
and U8974 (N_8974,N_4371,N_3904);
nor U8975 (N_8975,N_3240,N_4941);
nor U8976 (N_8976,N_5297,N_3635);
or U8977 (N_8977,N_3720,N_4388);
or U8978 (N_8978,N_4812,N_5988);
nor U8979 (N_8979,N_4507,N_5551);
nor U8980 (N_8980,N_5481,N_6166);
and U8981 (N_8981,N_3662,N_5469);
nand U8982 (N_8982,N_5558,N_6060);
or U8983 (N_8983,N_5292,N_5119);
xor U8984 (N_8984,N_5473,N_4495);
and U8985 (N_8985,N_4455,N_4238);
xnor U8986 (N_8986,N_4418,N_3219);
xor U8987 (N_8987,N_3983,N_4008);
xor U8988 (N_8988,N_5499,N_3959);
and U8989 (N_8989,N_4055,N_4965);
nand U8990 (N_8990,N_3722,N_4060);
nor U8991 (N_8991,N_3131,N_5827);
nand U8992 (N_8992,N_3687,N_5202);
and U8993 (N_8993,N_4019,N_4220);
or U8994 (N_8994,N_6064,N_3322);
and U8995 (N_8995,N_5670,N_4350);
and U8996 (N_8996,N_3229,N_5702);
xnor U8997 (N_8997,N_4332,N_3222);
and U8998 (N_8998,N_3293,N_3909);
and U8999 (N_8999,N_5879,N_4819);
and U9000 (N_9000,N_4888,N_4909);
xnor U9001 (N_9001,N_5481,N_4833);
nand U9002 (N_9002,N_3313,N_3286);
xnor U9003 (N_9003,N_4649,N_4040);
xor U9004 (N_9004,N_6245,N_4240);
and U9005 (N_9005,N_5089,N_3308);
xor U9006 (N_9006,N_5148,N_4291);
and U9007 (N_9007,N_4445,N_4208);
xnor U9008 (N_9008,N_4756,N_6128);
xor U9009 (N_9009,N_3218,N_4892);
nor U9010 (N_9010,N_5412,N_4535);
xnor U9011 (N_9011,N_5472,N_5840);
xnor U9012 (N_9012,N_3747,N_6045);
nand U9013 (N_9013,N_4052,N_4580);
and U9014 (N_9014,N_3549,N_4681);
and U9015 (N_9015,N_5796,N_5027);
xor U9016 (N_9016,N_6150,N_3246);
xor U9017 (N_9017,N_3718,N_3826);
nor U9018 (N_9018,N_5360,N_3368);
nand U9019 (N_9019,N_5679,N_5742);
or U9020 (N_9020,N_4394,N_5565);
and U9021 (N_9021,N_3196,N_5802);
nor U9022 (N_9022,N_5711,N_5723);
xnor U9023 (N_9023,N_3389,N_5999);
nand U9024 (N_9024,N_4758,N_3487);
nand U9025 (N_9025,N_3468,N_3998);
xnor U9026 (N_9026,N_4160,N_4490);
nor U9027 (N_9027,N_5649,N_3694);
xnor U9028 (N_9028,N_3637,N_4252);
nor U9029 (N_9029,N_4909,N_6156);
nor U9030 (N_9030,N_5173,N_4761);
xor U9031 (N_9031,N_5091,N_3566);
nand U9032 (N_9032,N_6015,N_5650);
nand U9033 (N_9033,N_4189,N_4705);
xor U9034 (N_9034,N_5257,N_4833);
or U9035 (N_9035,N_6229,N_5086);
xor U9036 (N_9036,N_3264,N_5327);
and U9037 (N_9037,N_6053,N_5895);
nand U9038 (N_9038,N_3161,N_6032);
nand U9039 (N_9039,N_5801,N_4654);
and U9040 (N_9040,N_6133,N_5516);
and U9041 (N_9041,N_6011,N_3585);
nand U9042 (N_9042,N_5978,N_6022);
or U9043 (N_9043,N_3709,N_3290);
or U9044 (N_9044,N_5225,N_4582);
nor U9045 (N_9045,N_4842,N_4452);
nor U9046 (N_9046,N_5395,N_5599);
and U9047 (N_9047,N_5838,N_4885);
or U9048 (N_9048,N_5171,N_5438);
nand U9049 (N_9049,N_4631,N_4909);
or U9050 (N_9050,N_6193,N_6140);
nor U9051 (N_9051,N_4371,N_4151);
or U9052 (N_9052,N_3493,N_4661);
xor U9053 (N_9053,N_3222,N_4556);
or U9054 (N_9054,N_5963,N_3584);
xnor U9055 (N_9055,N_5007,N_3386);
nand U9056 (N_9056,N_3717,N_5190);
nor U9057 (N_9057,N_3357,N_4485);
and U9058 (N_9058,N_4896,N_5524);
nand U9059 (N_9059,N_3434,N_5911);
and U9060 (N_9060,N_3968,N_4901);
or U9061 (N_9061,N_3914,N_4875);
and U9062 (N_9062,N_4852,N_5078);
or U9063 (N_9063,N_3902,N_5501);
nand U9064 (N_9064,N_5146,N_5025);
xor U9065 (N_9065,N_6149,N_3773);
and U9066 (N_9066,N_4581,N_4216);
nor U9067 (N_9067,N_5980,N_5985);
nor U9068 (N_9068,N_3148,N_3179);
or U9069 (N_9069,N_5017,N_4623);
and U9070 (N_9070,N_3269,N_4821);
and U9071 (N_9071,N_4038,N_3251);
xor U9072 (N_9072,N_6073,N_3840);
nor U9073 (N_9073,N_6223,N_3940);
nand U9074 (N_9074,N_5202,N_3130);
nor U9075 (N_9075,N_3666,N_4829);
or U9076 (N_9076,N_4942,N_4035);
or U9077 (N_9077,N_4937,N_4899);
nand U9078 (N_9078,N_4360,N_3990);
or U9079 (N_9079,N_5254,N_5649);
and U9080 (N_9080,N_6150,N_5789);
or U9081 (N_9081,N_6111,N_5616);
nor U9082 (N_9082,N_5485,N_5922);
or U9083 (N_9083,N_3767,N_5290);
nor U9084 (N_9084,N_5289,N_4238);
nor U9085 (N_9085,N_6232,N_3812);
or U9086 (N_9086,N_3255,N_5539);
nand U9087 (N_9087,N_5087,N_4225);
and U9088 (N_9088,N_4778,N_3401);
nand U9089 (N_9089,N_4468,N_4622);
or U9090 (N_9090,N_4616,N_5446);
nand U9091 (N_9091,N_6244,N_3568);
and U9092 (N_9092,N_4487,N_5134);
xnor U9093 (N_9093,N_4310,N_6247);
and U9094 (N_9094,N_4543,N_5828);
xor U9095 (N_9095,N_4032,N_5024);
xor U9096 (N_9096,N_4512,N_3285);
or U9097 (N_9097,N_4027,N_3270);
xnor U9098 (N_9098,N_5458,N_4566);
nor U9099 (N_9099,N_3744,N_5997);
nor U9100 (N_9100,N_5273,N_3724);
nor U9101 (N_9101,N_4436,N_3811);
xnor U9102 (N_9102,N_4496,N_5753);
and U9103 (N_9103,N_5473,N_5998);
nand U9104 (N_9104,N_6043,N_4902);
and U9105 (N_9105,N_4353,N_4765);
nor U9106 (N_9106,N_4869,N_3279);
or U9107 (N_9107,N_5454,N_5550);
or U9108 (N_9108,N_5031,N_5972);
nand U9109 (N_9109,N_3978,N_3709);
nand U9110 (N_9110,N_5536,N_5395);
or U9111 (N_9111,N_5827,N_5502);
nand U9112 (N_9112,N_5862,N_3962);
and U9113 (N_9113,N_3481,N_5297);
and U9114 (N_9114,N_5055,N_3796);
xor U9115 (N_9115,N_3759,N_5319);
xor U9116 (N_9116,N_5518,N_4805);
or U9117 (N_9117,N_4326,N_4904);
nor U9118 (N_9118,N_5846,N_5783);
xnor U9119 (N_9119,N_5111,N_5948);
nor U9120 (N_9120,N_3302,N_5299);
nand U9121 (N_9121,N_4377,N_5525);
nor U9122 (N_9122,N_5728,N_5404);
xnor U9123 (N_9123,N_6005,N_3677);
and U9124 (N_9124,N_5375,N_3341);
xnor U9125 (N_9125,N_4164,N_4536);
or U9126 (N_9126,N_5712,N_5130);
and U9127 (N_9127,N_4880,N_3738);
nand U9128 (N_9128,N_5668,N_4108);
nor U9129 (N_9129,N_4341,N_5915);
nand U9130 (N_9130,N_4070,N_5432);
and U9131 (N_9131,N_3729,N_3832);
nor U9132 (N_9132,N_4700,N_4173);
or U9133 (N_9133,N_5175,N_5007);
or U9134 (N_9134,N_3825,N_3183);
nor U9135 (N_9135,N_6057,N_3345);
and U9136 (N_9136,N_5641,N_4018);
xnor U9137 (N_9137,N_4016,N_5229);
nor U9138 (N_9138,N_5624,N_4277);
nand U9139 (N_9139,N_3767,N_6163);
and U9140 (N_9140,N_5309,N_5164);
xor U9141 (N_9141,N_5251,N_6177);
nand U9142 (N_9142,N_4907,N_5734);
and U9143 (N_9143,N_3440,N_6188);
xor U9144 (N_9144,N_3755,N_6178);
nand U9145 (N_9145,N_4708,N_3916);
nor U9146 (N_9146,N_3662,N_3492);
or U9147 (N_9147,N_5118,N_5945);
nand U9148 (N_9148,N_6152,N_5913);
nor U9149 (N_9149,N_6209,N_4183);
xnor U9150 (N_9150,N_3609,N_6229);
or U9151 (N_9151,N_5278,N_4435);
nor U9152 (N_9152,N_3463,N_3275);
nand U9153 (N_9153,N_4613,N_6173);
xnor U9154 (N_9154,N_4931,N_5603);
or U9155 (N_9155,N_5251,N_3573);
nor U9156 (N_9156,N_3211,N_4264);
or U9157 (N_9157,N_5873,N_4924);
nand U9158 (N_9158,N_3891,N_3899);
xnor U9159 (N_9159,N_3863,N_4529);
xor U9160 (N_9160,N_3939,N_4105);
and U9161 (N_9161,N_4778,N_4348);
and U9162 (N_9162,N_5725,N_3804);
and U9163 (N_9163,N_5682,N_5647);
and U9164 (N_9164,N_5262,N_4189);
nor U9165 (N_9165,N_4914,N_5416);
nand U9166 (N_9166,N_3414,N_3509);
and U9167 (N_9167,N_6053,N_3826);
and U9168 (N_9168,N_3468,N_5673);
and U9169 (N_9169,N_3805,N_5283);
or U9170 (N_9170,N_3628,N_6207);
nor U9171 (N_9171,N_3413,N_3212);
or U9172 (N_9172,N_4368,N_5678);
nor U9173 (N_9173,N_3804,N_4482);
xor U9174 (N_9174,N_4992,N_4597);
xor U9175 (N_9175,N_5498,N_5818);
nor U9176 (N_9176,N_5211,N_4667);
or U9177 (N_9177,N_3376,N_4838);
and U9178 (N_9178,N_3809,N_5116);
or U9179 (N_9179,N_5730,N_5100);
xnor U9180 (N_9180,N_3242,N_4054);
nand U9181 (N_9181,N_5969,N_5646);
xor U9182 (N_9182,N_6159,N_4891);
nand U9183 (N_9183,N_4915,N_4816);
and U9184 (N_9184,N_3790,N_6053);
or U9185 (N_9185,N_4859,N_5393);
or U9186 (N_9186,N_4093,N_4334);
xor U9187 (N_9187,N_4194,N_4592);
or U9188 (N_9188,N_5738,N_5290);
and U9189 (N_9189,N_3931,N_3650);
xnor U9190 (N_9190,N_6198,N_3483);
or U9191 (N_9191,N_4437,N_4978);
xnor U9192 (N_9192,N_5702,N_3320);
nand U9193 (N_9193,N_4975,N_4213);
nand U9194 (N_9194,N_3986,N_3163);
nand U9195 (N_9195,N_4138,N_5609);
xor U9196 (N_9196,N_3264,N_3517);
nor U9197 (N_9197,N_3542,N_5434);
nand U9198 (N_9198,N_5354,N_5705);
or U9199 (N_9199,N_5676,N_5760);
nor U9200 (N_9200,N_4365,N_4563);
or U9201 (N_9201,N_5308,N_3985);
nand U9202 (N_9202,N_6009,N_5722);
and U9203 (N_9203,N_5061,N_4721);
or U9204 (N_9204,N_3723,N_4145);
xor U9205 (N_9205,N_5890,N_4604);
nor U9206 (N_9206,N_3754,N_5668);
or U9207 (N_9207,N_6216,N_4529);
or U9208 (N_9208,N_4117,N_6086);
xnor U9209 (N_9209,N_5055,N_3294);
nor U9210 (N_9210,N_5717,N_4017);
and U9211 (N_9211,N_5823,N_3823);
nand U9212 (N_9212,N_3249,N_5520);
xnor U9213 (N_9213,N_5729,N_3366);
xnor U9214 (N_9214,N_5837,N_3974);
or U9215 (N_9215,N_3646,N_3993);
nand U9216 (N_9216,N_5862,N_5074);
nor U9217 (N_9217,N_5560,N_5428);
nor U9218 (N_9218,N_5002,N_4376);
nand U9219 (N_9219,N_4953,N_4739);
nand U9220 (N_9220,N_4986,N_5669);
or U9221 (N_9221,N_4687,N_3977);
xor U9222 (N_9222,N_4333,N_4790);
and U9223 (N_9223,N_3988,N_4024);
xor U9224 (N_9224,N_4034,N_4127);
nand U9225 (N_9225,N_5123,N_5182);
nand U9226 (N_9226,N_5830,N_3644);
nor U9227 (N_9227,N_5576,N_4603);
or U9228 (N_9228,N_5181,N_5157);
and U9229 (N_9229,N_5317,N_3998);
and U9230 (N_9230,N_4906,N_5092);
and U9231 (N_9231,N_3923,N_5739);
nor U9232 (N_9232,N_5222,N_4300);
or U9233 (N_9233,N_3745,N_5581);
nand U9234 (N_9234,N_5220,N_5249);
or U9235 (N_9235,N_4075,N_4284);
or U9236 (N_9236,N_5626,N_5414);
or U9237 (N_9237,N_4487,N_4446);
nand U9238 (N_9238,N_5131,N_4729);
or U9239 (N_9239,N_3146,N_5923);
nand U9240 (N_9240,N_4349,N_5619);
and U9241 (N_9241,N_4072,N_5923);
nand U9242 (N_9242,N_5822,N_3953);
or U9243 (N_9243,N_3353,N_3834);
and U9244 (N_9244,N_4986,N_5963);
or U9245 (N_9245,N_3956,N_5357);
or U9246 (N_9246,N_4014,N_5760);
nand U9247 (N_9247,N_3479,N_6050);
xnor U9248 (N_9248,N_3836,N_3156);
or U9249 (N_9249,N_3623,N_3527);
and U9250 (N_9250,N_3645,N_5908);
xor U9251 (N_9251,N_4690,N_4890);
nor U9252 (N_9252,N_3297,N_6188);
or U9253 (N_9253,N_6243,N_4634);
and U9254 (N_9254,N_4764,N_5809);
nor U9255 (N_9255,N_5162,N_4874);
nand U9256 (N_9256,N_4129,N_3516);
or U9257 (N_9257,N_3990,N_3888);
nor U9258 (N_9258,N_6103,N_5783);
and U9259 (N_9259,N_5595,N_4401);
nand U9260 (N_9260,N_6194,N_5131);
nand U9261 (N_9261,N_4848,N_3128);
nor U9262 (N_9262,N_4607,N_3375);
and U9263 (N_9263,N_5614,N_4635);
xor U9264 (N_9264,N_4312,N_4231);
xor U9265 (N_9265,N_6248,N_4601);
nand U9266 (N_9266,N_4009,N_5253);
or U9267 (N_9267,N_6103,N_5242);
nor U9268 (N_9268,N_4665,N_5564);
nand U9269 (N_9269,N_4750,N_5617);
xor U9270 (N_9270,N_5373,N_6038);
nor U9271 (N_9271,N_5521,N_5298);
nand U9272 (N_9272,N_3256,N_4787);
or U9273 (N_9273,N_4689,N_6230);
nand U9274 (N_9274,N_3851,N_4188);
or U9275 (N_9275,N_4875,N_5130);
nand U9276 (N_9276,N_5845,N_3853);
nor U9277 (N_9277,N_4761,N_3958);
nand U9278 (N_9278,N_5766,N_5015);
nor U9279 (N_9279,N_3711,N_3230);
nand U9280 (N_9280,N_4005,N_3181);
xnor U9281 (N_9281,N_4357,N_4153);
nor U9282 (N_9282,N_5637,N_3949);
nor U9283 (N_9283,N_4915,N_5343);
nor U9284 (N_9284,N_3500,N_4943);
and U9285 (N_9285,N_3696,N_4490);
and U9286 (N_9286,N_3542,N_5889);
or U9287 (N_9287,N_5577,N_3481);
nor U9288 (N_9288,N_5120,N_3734);
nor U9289 (N_9289,N_3551,N_4175);
nor U9290 (N_9290,N_4938,N_4751);
nor U9291 (N_9291,N_5474,N_6054);
nor U9292 (N_9292,N_4137,N_3721);
nor U9293 (N_9293,N_3686,N_3249);
nand U9294 (N_9294,N_3498,N_3591);
nand U9295 (N_9295,N_5023,N_4325);
nand U9296 (N_9296,N_5697,N_5816);
nor U9297 (N_9297,N_6019,N_3594);
or U9298 (N_9298,N_6137,N_3140);
nor U9299 (N_9299,N_5209,N_3410);
nand U9300 (N_9300,N_3656,N_3977);
and U9301 (N_9301,N_3835,N_4576);
nor U9302 (N_9302,N_4437,N_5268);
nor U9303 (N_9303,N_5316,N_3811);
or U9304 (N_9304,N_3627,N_3552);
nor U9305 (N_9305,N_3772,N_4932);
nor U9306 (N_9306,N_5792,N_5583);
and U9307 (N_9307,N_5001,N_5821);
nor U9308 (N_9308,N_5377,N_5984);
xnor U9309 (N_9309,N_4609,N_4856);
xnor U9310 (N_9310,N_6168,N_3890);
and U9311 (N_9311,N_5316,N_3964);
and U9312 (N_9312,N_3188,N_4482);
and U9313 (N_9313,N_3289,N_4422);
or U9314 (N_9314,N_5482,N_4072);
nor U9315 (N_9315,N_6076,N_5130);
xnor U9316 (N_9316,N_6084,N_5503);
or U9317 (N_9317,N_3439,N_4156);
nand U9318 (N_9318,N_4152,N_5457);
xor U9319 (N_9319,N_3731,N_3558);
xor U9320 (N_9320,N_4353,N_3399);
nor U9321 (N_9321,N_3589,N_5830);
nand U9322 (N_9322,N_3609,N_5383);
and U9323 (N_9323,N_5264,N_3444);
xor U9324 (N_9324,N_5990,N_4603);
xor U9325 (N_9325,N_3317,N_5995);
nor U9326 (N_9326,N_5972,N_4810);
nor U9327 (N_9327,N_4089,N_5761);
or U9328 (N_9328,N_3512,N_4054);
nor U9329 (N_9329,N_4299,N_3205);
nand U9330 (N_9330,N_5250,N_3137);
nor U9331 (N_9331,N_4106,N_3925);
nand U9332 (N_9332,N_5368,N_5487);
or U9333 (N_9333,N_3270,N_5799);
xnor U9334 (N_9334,N_5177,N_3950);
xor U9335 (N_9335,N_5706,N_5929);
and U9336 (N_9336,N_5665,N_4662);
xnor U9337 (N_9337,N_3567,N_5545);
nor U9338 (N_9338,N_3590,N_3449);
or U9339 (N_9339,N_4849,N_5715);
xor U9340 (N_9340,N_4855,N_4405);
nand U9341 (N_9341,N_4750,N_3842);
nand U9342 (N_9342,N_3580,N_3314);
xor U9343 (N_9343,N_4606,N_5687);
or U9344 (N_9344,N_3546,N_4784);
xor U9345 (N_9345,N_3268,N_3274);
nand U9346 (N_9346,N_4079,N_3240);
nor U9347 (N_9347,N_3903,N_4499);
nand U9348 (N_9348,N_5509,N_3174);
xnor U9349 (N_9349,N_4946,N_5322);
xnor U9350 (N_9350,N_4809,N_5855);
and U9351 (N_9351,N_5960,N_4283);
nor U9352 (N_9352,N_4454,N_6105);
or U9353 (N_9353,N_5918,N_3575);
nor U9354 (N_9354,N_3180,N_4503);
and U9355 (N_9355,N_5657,N_5400);
nor U9356 (N_9356,N_4283,N_5164);
nand U9357 (N_9357,N_3487,N_5964);
and U9358 (N_9358,N_5966,N_3198);
nand U9359 (N_9359,N_5543,N_4788);
nor U9360 (N_9360,N_5228,N_5427);
xor U9361 (N_9361,N_4140,N_4955);
or U9362 (N_9362,N_3128,N_4101);
nor U9363 (N_9363,N_3197,N_4980);
and U9364 (N_9364,N_3619,N_3964);
and U9365 (N_9365,N_5474,N_5103);
xnor U9366 (N_9366,N_4322,N_3650);
xnor U9367 (N_9367,N_5567,N_4389);
nor U9368 (N_9368,N_4950,N_3800);
nand U9369 (N_9369,N_5836,N_4849);
nor U9370 (N_9370,N_3319,N_5853);
or U9371 (N_9371,N_5922,N_5929);
xnor U9372 (N_9372,N_4911,N_4297);
or U9373 (N_9373,N_4634,N_5020);
nand U9374 (N_9374,N_6159,N_5800);
and U9375 (N_9375,N_8466,N_7481);
and U9376 (N_9376,N_7572,N_6388);
nand U9377 (N_9377,N_9255,N_7409);
xnor U9378 (N_9378,N_6433,N_7161);
nor U9379 (N_9379,N_8038,N_9160);
nand U9380 (N_9380,N_6581,N_7862);
and U9381 (N_9381,N_7410,N_6450);
and U9382 (N_9382,N_7855,N_8076);
and U9383 (N_9383,N_8932,N_8473);
or U9384 (N_9384,N_6992,N_7851);
nand U9385 (N_9385,N_7835,N_6756);
or U9386 (N_9386,N_6725,N_7643);
nor U9387 (N_9387,N_8111,N_7813);
and U9388 (N_9388,N_7511,N_8701);
nand U9389 (N_9389,N_7273,N_9225);
nor U9390 (N_9390,N_7727,N_8313);
or U9391 (N_9391,N_6825,N_6389);
nor U9392 (N_9392,N_8833,N_7622);
nand U9393 (N_9393,N_6885,N_8642);
nand U9394 (N_9394,N_6552,N_7430);
nor U9395 (N_9395,N_7571,N_8788);
or U9396 (N_9396,N_6928,N_7558);
xnor U9397 (N_9397,N_7889,N_7756);
xor U9398 (N_9398,N_7929,N_7610);
and U9399 (N_9399,N_6630,N_8534);
xnor U9400 (N_9400,N_7499,N_8538);
nand U9401 (N_9401,N_7767,N_7704);
or U9402 (N_9402,N_9054,N_8875);
nand U9403 (N_9403,N_6976,N_8964);
nor U9404 (N_9404,N_9170,N_8748);
nand U9405 (N_9405,N_8605,N_6390);
or U9406 (N_9406,N_7554,N_7212);
xnor U9407 (N_9407,N_6577,N_6599);
or U9408 (N_9408,N_8384,N_6662);
xor U9409 (N_9409,N_6872,N_8753);
and U9410 (N_9410,N_8958,N_7260);
and U9411 (N_9411,N_8310,N_8557);
nor U9412 (N_9412,N_8755,N_8287);
xor U9413 (N_9413,N_6923,N_7111);
xnor U9414 (N_9414,N_7600,N_9175);
xor U9415 (N_9415,N_8357,N_7897);
nand U9416 (N_9416,N_7004,N_7760);
and U9417 (N_9417,N_6322,N_8798);
or U9418 (N_9418,N_6408,N_7715);
and U9419 (N_9419,N_8147,N_9156);
or U9420 (N_9420,N_6684,N_7561);
nor U9421 (N_9421,N_7313,N_7706);
and U9422 (N_9422,N_8648,N_8714);
and U9423 (N_9423,N_7799,N_7315);
xnor U9424 (N_9424,N_8823,N_7596);
or U9425 (N_9425,N_7143,N_6698);
nand U9426 (N_9426,N_9226,N_8962);
or U9427 (N_9427,N_9277,N_9005);
xor U9428 (N_9428,N_8026,N_8304);
nor U9429 (N_9429,N_7175,N_8156);
and U9430 (N_9430,N_9245,N_7408);
and U9431 (N_9431,N_7562,N_9114);
nand U9432 (N_9432,N_8807,N_8834);
or U9433 (N_9433,N_8355,N_6357);
xnor U9434 (N_9434,N_6472,N_7689);
and U9435 (N_9435,N_6501,N_7682);
xnor U9436 (N_9436,N_9167,N_7364);
nand U9437 (N_9437,N_8426,N_6980);
and U9438 (N_9438,N_8924,N_7263);
nand U9439 (N_9439,N_7310,N_7136);
and U9440 (N_9440,N_6373,N_8035);
nor U9441 (N_9441,N_7493,N_7538);
nor U9442 (N_9442,N_8526,N_7265);
and U9443 (N_9443,N_8133,N_6283);
nor U9444 (N_9444,N_6724,N_7083);
xnor U9445 (N_9445,N_8090,N_7747);
and U9446 (N_9446,N_8439,N_6528);
nand U9447 (N_9447,N_7342,N_9107);
or U9448 (N_9448,N_7729,N_7589);
nor U9449 (N_9449,N_8941,N_6848);
xnor U9450 (N_9450,N_7033,N_6302);
nand U9451 (N_9451,N_7158,N_6739);
and U9452 (N_9452,N_7658,N_7061);
xnor U9453 (N_9453,N_8786,N_8578);
xnor U9454 (N_9454,N_8951,N_7761);
nor U9455 (N_9455,N_7051,N_7288);
nor U9456 (N_9456,N_7241,N_6371);
nand U9457 (N_9457,N_7619,N_8105);
xnor U9458 (N_9458,N_6958,N_8849);
and U9459 (N_9459,N_6913,N_6447);
nor U9460 (N_9460,N_7476,N_6732);
xor U9461 (N_9461,N_6515,N_6588);
nand U9462 (N_9462,N_7529,N_7047);
nor U9463 (N_9463,N_7854,N_6748);
nand U9464 (N_9464,N_7565,N_6328);
nand U9465 (N_9465,N_8937,N_7043);
xor U9466 (N_9466,N_6961,N_8194);
or U9467 (N_9467,N_6579,N_8570);
and U9468 (N_9468,N_8174,N_6644);
nand U9469 (N_9469,N_6652,N_9230);
nor U9470 (N_9470,N_9066,N_8416);
or U9471 (N_9471,N_7036,N_8083);
nand U9472 (N_9472,N_8303,N_6726);
or U9473 (N_9473,N_8375,N_6353);
xnor U9474 (N_9474,N_7464,N_8424);
nand U9475 (N_9475,N_8281,N_9016);
xor U9476 (N_9476,N_7293,N_7868);
or U9477 (N_9477,N_7954,N_6944);
or U9478 (N_9478,N_8922,N_8977);
and U9479 (N_9479,N_9145,N_7216);
nand U9480 (N_9480,N_9110,N_6657);
and U9481 (N_9481,N_7318,N_6808);
or U9482 (N_9482,N_7392,N_7469);
nor U9483 (N_9483,N_9261,N_6769);
or U9484 (N_9484,N_8978,N_8627);
xor U9485 (N_9485,N_8617,N_7080);
or U9486 (N_9486,N_7181,N_6763);
and U9487 (N_9487,N_8521,N_8167);
nand U9488 (N_9488,N_6266,N_7594);
and U9489 (N_9489,N_8134,N_6558);
or U9490 (N_9490,N_7259,N_8609);
and U9491 (N_9491,N_6999,N_8612);
xnor U9492 (N_9492,N_8270,N_6770);
nand U9493 (N_9493,N_6379,N_8395);
or U9494 (N_9494,N_6533,N_7305);
and U9495 (N_9495,N_8241,N_9007);
xnor U9496 (N_9496,N_6274,N_8649);
nor U9497 (N_9497,N_7074,N_6643);
xnor U9498 (N_9498,N_7001,N_7830);
and U9499 (N_9499,N_6585,N_8278);
and U9500 (N_9500,N_6674,N_7450);
and U9501 (N_9501,N_6950,N_8884);
or U9502 (N_9502,N_7840,N_7962);
xnor U9503 (N_9503,N_9142,N_7133);
nand U9504 (N_9504,N_6440,N_8293);
nand U9505 (N_9505,N_7362,N_7483);
and U9506 (N_9506,N_8269,N_8496);
nor U9507 (N_9507,N_7875,N_6667);
nand U9508 (N_9508,N_6418,N_7953);
xnor U9509 (N_9509,N_6295,N_6859);
and U9510 (N_9510,N_8647,N_6776);
or U9511 (N_9511,N_8120,N_6300);
or U9512 (N_9512,N_8117,N_8498);
or U9513 (N_9513,N_6460,N_9311);
or U9514 (N_9514,N_8663,N_9303);
or U9515 (N_9515,N_7322,N_7921);
xnor U9516 (N_9516,N_7327,N_8660);
or U9517 (N_9517,N_6653,N_9089);
nand U9518 (N_9518,N_9320,N_8816);
and U9519 (N_9519,N_7946,N_7349);
nor U9520 (N_9520,N_9258,N_7809);
or U9521 (N_9521,N_8773,N_7130);
nand U9522 (N_9522,N_7871,N_6613);
and U9523 (N_9523,N_6890,N_8979);
nand U9524 (N_9524,N_7970,N_7787);
nand U9525 (N_9525,N_8193,N_6995);
nor U9526 (N_9526,N_6733,N_6744);
nor U9527 (N_9527,N_7780,N_6939);
and U9528 (N_9528,N_7247,N_7724);
or U9529 (N_9529,N_6555,N_8427);
and U9530 (N_9530,N_6735,N_7888);
nor U9531 (N_9531,N_6781,N_7695);
nor U9532 (N_9532,N_9214,N_7505);
nand U9533 (N_9533,N_8210,N_7959);
nand U9534 (N_9534,N_7354,N_8691);
xnor U9535 (N_9535,N_7307,N_8731);
xnor U9536 (N_9536,N_6773,N_8852);
and U9537 (N_9537,N_7431,N_7226);
and U9538 (N_9538,N_7118,N_7574);
and U9539 (N_9539,N_8409,N_7188);
or U9540 (N_9540,N_8213,N_9361);
or U9541 (N_9541,N_6278,N_9048);
nor U9542 (N_9542,N_6696,N_8228);
and U9543 (N_9543,N_8668,N_6719);
and U9544 (N_9544,N_6737,N_8780);
nor U9545 (N_9545,N_9331,N_9201);
nand U9546 (N_9546,N_9003,N_7943);
or U9547 (N_9547,N_8616,N_7530);
xor U9548 (N_9548,N_7473,N_6441);
nor U9549 (N_9549,N_7991,N_7150);
or U9550 (N_9550,N_6453,N_7420);
or U9551 (N_9551,N_7580,N_9124);
nand U9552 (N_9552,N_7053,N_6953);
xor U9553 (N_9553,N_6801,N_7416);
and U9554 (N_9554,N_7687,N_8596);
nor U9555 (N_9555,N_8464,N_8611);
or U9556 (N_9556,N_8018,N_6749);
xnor U9557 (N_9557,N_7942,N_7478);
nand U9558 (N_9558,N_9266,N_7979);
xor U9559 (N_9559,N_8713,N_8592);
and U9560 (N_9560,N_9295,N_7365);
nand U9561 (N_9561,N_8170,N_7350);
or U9562 (N_9562,N_7725,N_6396);
nand U9563 (N_9563,N_8399,N_8672);
nand U9564 (N_9564,N_8494,N_8207);
or U9565 (N_9565,N_8577,N_6766);
or U9566 (N_9566,N_8805,N_8726);
nor U9567 (N_9567,N_6843,N_8141);
nor U9568 (N_9568,N_8721,N_8106);
xnor U9569 (N_9569,N_6655,N_7534);
and U9570 (N_9570,N_8022,N_6506);
xor U9571 (N_9571,N_8190,N_8636);
xnor U9572 (N_9572,N_9158,N_8275);
xnor U9573 (N_9573,N_7272,N_6339);
nor U9574 (N_9574,N_8012,N_7746);
and U9575 (N_9575,N_9302,N_8926);
or U9576 (N_9576,N_8728,N_7249);
xnor U9577 (N_9577,N_9132,N_9011);
xnor U9578 (N_9578,N_7264,N_6865);
or U9579 (N_9579,N_8499,N_6443);
nor U9580 (N_9580,N_7474,N_7820);
and U9581 (N_9581,N_9351,N_8305);
xnor U9582 (N_9582,N_7944,N_7831);
or U9583 (N_9583,N_6356,N_9210);
nand U9584 (N_9584,N_8420,N_6341);
or U9585 (N_9585,N_8793,N_7964);
nor U9586 (N_9586,N_8178,N_7200);
nand U9587 (N_9587,N_6629,N_8583);
nor U9588 (N_9588,N_6586,N_6967);
nand U9589 (N_9589,N_7583,N_9056);
nor U9590 (N_9590,N_7577,N_7328);
xor U9591 (N_9591,N_9161,N_9026);
and U9592 (N_9592,N_8478,N_8162);
or U9593 (N_9593,N_8573,N_6805);
or U9594 (N_9594,N_6260,N_6779);
and U9595 (N_9595,N_6642,N_8891);
nor U9596 (N_9596,N_8812,N_9122);
and U9597 (N_9597,N_7590,N_7193);
nor U9598 (N_9598,N_9013,N_6512);
and U9599 (N_9599,N_7904,N_6659);
or U9600 (N_9600,N_7123,N_6831);
nand U9601 (N_9601,N_8486,N_8931);
nor U9602 (N_9602,N_8048,N_6718);
xnor U9603 (N_9603,N_6888,N_6432);
xnor U9604 (N_9604,N_8936,N_7177);
or U9605 (N_9605,N_9061,N_9123);
nor U9606 (N_9606,N_6271,N_7935);
nand U9607 (N_9607,N_8692,N_8010);
xnor U9608 (N_9608,N_9355,N_8382);
and U9609 (N_9609,N_7939,N_6827);
or U9610 (N_9610,N_7765,N_7543);
nand U9611 (N_9611,N_6452,N_8121);
or U9612 (N_9612,N_6618,N_8238);
or U9613 (N_9613,N_6332,N_8738);
nand U9614 (N_9614,N_7106,N_6741);
nor U9615 (N_9615,N_8890,N_8835);
xnor U9616 (N_9616,N_8242,N_7743);
nand U9617 (N_9617,N_6985,N_8846);
nor U9618 (N_9618,N_8719,N_7256);
nand U9619 (N_9619,N_7826,N_7646);
or U9620 (N_9620,N_6331,N_6790);
nand U9621 (N_9621,N_8710,N_7545);
nor U9622 (N_9622,N_6968,N_7320);
nor U9623 (N_9623,N_8227,N_6706);
and U9624 (N_9624,N_8320,N_6437);
and U9625 (N_9625,N_6660,N_8002);
xor U9626 (N_9626,N_8272,N_7022);
or U9627 (N_9627,N_7209,N_6812);
nor U9628 (N_9628,N_8109,N_8024);
xor U9629 (N_9629,N_8969,N_7205);
xnor U9630 (N_9630,N_7269,N_7628);
xor U9631 (N_9631,N_7852,N_8075);
nand U9632 (N_9632,N_6394,N_8838);
nand U9633 (N_9633,N_8665,N_6424);
xnor U9634 (N_9634,N_6678,N_8667);
nor U9635 (N_9635,N_9165,N_8944);
or U9636 (N_9636,N_6477,N_7699);
nor U9637 (N_9637,N_6947,N_7599);
nor U9638 (N_9638,N_6656,N_8327);
xnor U9639 (N_9639,N_8172,N_7220);
and U9640 (N_9640,N_8907,N_7718);
nand U9641 (N_9641,N_8234,N_6858);
nor U9642 (N_9642,N_9280,N_8436);
and U9643 (N_9643,N_7708,N_6596);
and U9644 (N_9644,N_8548,N_9119);
nor U9645 (N_9645,N_7721,N_6896);
xnor U9646 (N_9646,N_8959,N_7870);
nand U9647 (N_9647,N_7611,N_6454);
xor U9648 (N_9648,N_7109,N_9330);
or U9649 (N_9649,N_9128,N_8481);
or U9650 (N_9650,N_7500,N_8935);
nand U9651 (N_9651,N_8462,N_8998);
nor U9652 (N_9652,N_8380,N_7941);
and U9653 (N_9653,N_8894,N_7267);
nand U9654 (N_9654,N_8232,N_7988);
nor U9655 (N_9655,N_6583,N_6905);
nand U9656 (N_9656,N_6612,N_8608);
nand U9657 (N_9657,N_8550,N_8973);
nor U9658 (N_9658,N_7463,N_6608);
and U9659 (N_9659,N_8068,N_8604);
nand U9660 (N_9660,N_6638,N_8370);
nor U9661 (N_9661,N_7506,N_6291);
nor U9662 (N_9662,N_7148,N_7861);
nor U9663 (N_9663,N_7012,N_7686);
nor U9664 (N_9664,N_6764,N_6720);
or U9665 (N_9665,N_8869,N_9273);
or U9666 (N_9666,N_8376,N_7225);
or U9667 (N_9667,N_8470,N_6935);
xnor U9668 (N_9668,N_7117,N_6987);
nor U9669 (N_9669,N_8872,N_6270);
or U9670 (N_9670,N_7383,N_6716);
and U9671 (N_9671,N_7395,N_6826);
xnor U9672 (N_9672,N_8552,N_8334);
nor U9673 (N_9673,N_7849,N_7020);
xnor U9674 (N_9674,N_8743,N_7556);
xnor U9675 (N_9675,N_8744,N_6646);
nand U9676 (N_9676,N_6308,N_8960);
nand U9677 (N_9677,N_7903,N_8994);
and U9678 (N_9678,N_7211,N_8880);
or U9679 (N_9679,N_6839,N_6411);
and U9680 (N_9680,N_6800,N_8980);
or U9681 (N_9681,N_6884,N_7893);
nor U9682 (N_9682,N_8523,N_7741);
xor U9683 (N_9683,N_7905,N_9004);
nand U9684 (N_9684,N_9234,N_9324);
xor U9685 (N_9685,N_9130,N_7048);
nand U9686 (N_9686,N_7125,N_8878);
or U9687 (N_9687,N_7279,N_7966);
or U9688 (N_9688,N_7795,N_8483);
xnor U9689 (N_9689,N_7424,N_9106);
and U9690 (N_9690,N_7544,N_8367);
and U9691 (N_9691,N_8346,N_7494);
and U9692 (N_9692,N_7974,N_9012);
or U9693 (N_9693,N_9162,N_6478);
nor U9694 (N_9694,N_9293,N_8408);
nor U9695 (N_9695,N_8332,N_6574);
xor U9696 (N_9696,N_9323,N_7208);
nand U9697 (N_9697,N_6435,N_8383);
xor U9698 (N_9698,N_6866,N_6530);
or U9699 (N_9699,N_6787,N_8992);
and U9700 (N_9700,N_6677,N_7955);
nor U9701 (N_9701,N_9365,N_8019);
nor U9702 (N_9702,N_8271,N_8673);
xor U9703 (N_9703,N_7027,N_6610);
and U9704 (N_9704,N_8267,N_8542);
nand U9705 (N_9705,N_9038,N_6407);
or U9706 (N_9706,N_7050,N_6863);
or U9707 (N_9707,N_7798,N_7013);
or U9708 (N_9708,N_9035,N_6795);
and U9709 (N_9709,N_6650,N_8853);
and U9710 (N_9710,N_6742,N_9077);
xnor U9711 (N_9711,N_8511,N_7999);
or U9712 (N_9712,N_6484,N_7294);
or U9713 (N_9713,N_6523,N_8110);
nand U9714 (N_9714,N_8794,N_7372);
xnor U9715 (N_9715,N_7178,N_9197);
nor U9716 (N_9716,N_8779,N_8211);
nand U9717 (N_9717,N_8457,N_8956);
nand U9718 (N_9718,N_7857,N_6768);
and U9719 (N_9719,N_6938,N_7489);
or U9720 (N_9720,N_8413,N_7901);
nor U9721 (N_9721,N_7238,N_6820);
nand U9722 (N_9722,N_6286,N_6346);
xnor U9723 (N_9723,N_7195,N_7201);
and U9724 (N_9724,N_8707,N_8968);
nor U9725 (N_9725,N_8686,N_7387);
or U9726 (N_9726,N_6310,N_8594);
or U9727 (N_9727,N_8173,N_8288);
or U9728 (N_9728,N_9072,N_6933);
xor U9729 (N_9729,N_7927,N_8326);
and U9730 (N_9730,N_6648,N_6458);
nor U9731 (N_9731,N_8345,N_8634);
nand U9732 (N_9732,N_6397,N_8154);
nand U9733 (N_9733,N_9209,N_7366);
xnor U9734 (N_9734,N_7186,N_6974);
xnor U9735 (N_9735,N_9206,N_9271);
xnor U9736 (N_9736,N_8056,N_6774);
and U9737 (N_9737,N_9236,N_7821);
nand U9738 (N_9738,N_8306,N_7122);
nor U9739 (N_9739,N_7551,N_9363);
nand U9740 (N_9740,N_9166,N_6651);
nand U9741 (N_9741,N_7906,N_7958);
and U9742 (N_9742,N_6500,N_6714);
and U9743 (N_9743,N_8803,N_8114);
nor U9744 (N_9744,N_6319,N_6609);
nor U9745 (N_9745,N_7784,N_6936);
or U9746 (N_9746,N_8323,N_8644);
nor U9747 (N_9747,N_8214,N_7184);
or U9748 (N_9748,N_8829,N_7251);
xnor U9749 (N_9749,N_6513,N_7341);
nand U9750 (N_9750,N_7025,N_8429);
xor U9751 (N_9751,N_6707,N_6889);
nand U9752 (N_9752,N_9334,N_6793);
nand U9753 (N_9753,N_9086,N_7427);
nor U9754 (N_9754,N_9100,N_6280);
nor U9755 (N_9755,N_6922,N_6367);
xnor U9756 (N_9756,N_8450,N_9317);
xnor U9757 (N_9757,N_8325,N_6311);
and U9758 (N_9758,N_8438,N_7847);
or U9759 (N_9759,N_8599,N_7128);
xnor U9760 (N_9760,N_7413,N_8045);
and U9761 (N_9761,N_6264,N_7710);
xnor U9762 (N_9762,N_6654,N_8089);
nor U9763 (N_9763,N_6519,N_7429);
or U9764 (N_9764,N_7948,N_9136);
xnor U9765 (N_9765,N_6544,N_6900);
or U9766 (N_9766,N_8940,N_8443);
xnor U9767 (N_9767,N_7446,N_7626);
nor U9768 (N_9768,N_7656,N_9050);
and U9769 (N_9769,N_6853,N_6497);
nor U9770 (N_9770,N_6546,N_7353);
nand U9771 (N_9771,N_8171,N_9370);
and U9772 (N_9772,N_7018,N_7252);
and U9773 (N_9773,N_9058,N_7522);
and U9774 (N_9774,N_8250,N_7603);
or U9775 (N_9775,N_8082,N_6814);
and U9776 (N_9776,N_8365,N_8913);
nor U9777 (N_9777,N_8736,N_7700);
and U9778 (N_9778,N_8784,N_8991);
nor U9779 (N_9779,N_8097,N_7286);
or U9780 (N_9780,N_6430,N_6597);
nand U9781 (N_9781,N_8311,N_8842);
nor U9782 (N_9782,N_9008,N_7652);
xnor U9783 (N_9783,N_7271,N_9265);
and U9784 (N_9784,N_6451,N_6897);
nor U9785 (N_9785,N_8757,N_8993);
nor U9786 (N_9786,N_7262,N_7093);
nand U9787 (N_9787,N_9143,N_7638);
xnor U9788 (N_9788,N_7236,N_7709);
xnor U9789 (N_9789,N_9071,N_6697);
and U9790 (N_9790,N_7221,N_6312);
nor U9791 (N_9791,N_9290,N_8440);
nor U9792 (N_9792,N_7641,N_7455);
nand U9793 (N_9793,N_6504,N_6626);
or U9794 (N_9794,N_9139,N_8296);
nor U9795 (N_9795,N_8001,N_7865);
xnor U9796 (N_9796,N_6767,N_6337);
and U9797 (N_9797,N_8766,N_8863);
xnor U9798 (N_9798,N_7996,N_8204);
xnor U9799 (N_9799,N_7065,N_9297);
and U9800 (N_9800,N_8387,N_8813);
and U9801 (N_9801,N_8815,N_6804);
xor U9802 (N_9802,N_8340,N_6746);
nor U9803 (N_9803,N_6604,N_7488);
xnor U9804 (N_9804,N_7266,N_6797);
xnor U9805 (N_9805,N_8220,N_8143);
xnor U9806 (N_9806,N_9272,N_7369);
or U9807 (N_9807,N_7711,N_8830);
and U9808 (N_9808,N_7087,N_8546);
and U9809 (N_9809,N_8430,N_9037);
nand U9810 (N_9810,N_9354,N_6669);
and U9811 (N_9811,N_8484,N_8014);
nor U9812 (N_9812,N_7067,N_6536);
and U9813 (N_9813,N_6565,N_6493);
nand U9814 (N_9814,N_6329,N_8292);
nor U9815 (N_9815,N_6284,N_6316);
nor U9816 (N_9816,N_8411,N_8831);
nand U9817 (N_9817,N_8914,N_8059);
xor U9818 (N_9818,N_6541,N_9034);
nor U9819 (N_9819,N_7470,N_7194);
xor U9820 (N_9820,N_8047,N_6632);
and U9821 (N_9821,N_8290,N_7564);
nor U9822 (N_9822,N_8585,N_6867);
nand U9823 (N_9823,N_8150,N_7425);
nand U9824 (N_9824,N_6907,N_9246);
nor U9825 (N_9825,N_8297,N_7245);
nor U9826 (N_9826,N_6279,N_6874);
and U9827 (N_9827,N_6870,N_7152);
nand U9828 (N_9828,N_6862,N_7933);
nor U9829 (N_9829,N_7578,N_7972);
or U9830 (N_9830,N_7400,N_8225);
or U9831 (N_9831,N_8509,N_7762);
nor U9832 (N_9832,N_7153,N_6305);
nand U9833 (N_9833,N_6971,N_8144);
or U9834 (N_9834,N_9239,N_8683);
xor U9835 (N_9835,N_7503,N_7566);
nor U9836 (N_9836,N_6979,N_7716);
and U9837 (N_9837,N_8801,N_9294);
nor U9838 (N_9838,N_8650,N_8360);
nand U9839 (N_9839,N_7797,N_6347);
xnor U9840 (N_9840,N_8525,N_6702);
nand U9841 (N_9841,N_8754,N_7398);
nor U9842 (N_9842,N_6465,N_8641);
xor U9843 (N_9843,N_7466,N_8752);
or U9844 (N_9844,N_7171,N_7844);
nor U9845 (N_9845,N_7298,N_6837);
and U9846 (N_9846,N_6649,N_6860);
nand U9847 (N_9847,N_7872,N_9319);
nand U9848 (N_9848,N_8976,N_6956);
xnor U9849 (N_9849,N_8329,N_7287);
nand U9850 (N_9850,N_6772,N_7777);
nor U9851 (N_9851,N_7361,N_8189);
nand U9852 (N_9852,N_7537,N_7640);
or U9853 (N_9853,N_6832,N_8566);
nor U9854 (N_9854,N_8851,N_8338);
and U9855 (N_9855,N_8747,N_9141);
nor U9856 (N_9856,N_6469,N_6780);
xnor U9857 (N_9857,N_7358,N_7121);
and U9858 (N_9858,N_8989,N_7015);
and U9859 (N_9859,N_7850,N_6645);
xnor U9860 (N_9860,N_6934,N_6338);
xor U9861 (N_9861,N_7671,N_6798);
nand U9862 (N_9862,N_6965,N_7802);
nand U9863 (N_9863,N_8301,N_8028);
or U9864 (N_9864,N_7460,N_7176);
nand U9865 (N_9865,N_8398,N_9018);
nor U9866 (N_9866,N_9149,N_7441);
or U9867 (N_9867,N_9275,N_7138);
or U9868 (N_9868,N_7547,N_6809);
nor U9869 (N_9869,N_7911,N_6351);
nand U9870 (N_9870,N_6691,N_9259);
or U9871 (N_9871,N_7764,N_8129);
or U9872 (N_9872,N_7145,N_6851);
xnor U9873 (N_9873,N_7846,N_9282);
xor U9874 (N_9874,N_7807,N_8351);
or U9875 (N_9875,N_8910,N_7011);
xor U9876 (N_9876,N_7951,N_8385);
xnor U9877 (N_9877,N_8274,N_9325);
xnor U9878 (N_9878,N_6481,N_8079);
or U9879 (N_9879,N_7768,N_7172);
xnor U9880 (N_9880,N_8164,N_7402);
nor U9881 (N_9881,N_8388,N_8434);
xor U9882 (N_9882,N_7334,N_7099);
nand U9883 (N_9883,N_8735,N_6761);
nor U9884 (N_9884,N_7546,N_8060);
and U9885 (N_9885,N_6842,N_8854);
xor U9886 (N_9886,N_6514,N_8553);
xor U9887 (N_9887,N_7060,N_7678);
xnor U9888 (N_9888,N_6562,N_8781);
nand U9889 (N_9889,N_7019,N_9291);
nor U9890 (N_9890,N_7078,N_8905);
nand U9891 (N_9891,N_7005,N_8750);
and U9892 (N_9892,N_8053,N_8988);
or U9893 (N_9893,N_6273,N_7276);
or U9894 (N_9894,N_9321,N_8695);
and U9895 (N_9895,N_9344,N_8597);
nor U9896 (N_9896,N_7137,N_6973);
or U9897 (N_9897,N_7705,N_9039);
or U9898 (N_9898,N_9276,N_9336);
nand U9899 (N_9899,N_8459,N_8229);
nand U9900 (N_9900,N_8545,N_7443);
or U9901 (N_9901,N_9359,N_9188);
nor U9902 (N_9902,N_8544,N_9080);
nand U9903 (N_9903,N_6502,N_9240);
xnor U9904 (N_9904,N_8814,N_8148);
or U9905 (N_9905,N_8446,N_8391);
and U9906 (N_9906,N_6395,N_7520);
nor U9907 (N_9907,N_6419,N_8651);
xnor U9908 (N_9908,N_9346,N_9349);
xor U9909 (N_9909,N_6695,N_8072);
nand U9910 (N_9910,N_9084,N_9308);
xnor U9911 (N_9911,N_8767,N_7308);
and U9912 (N_9912,N_7884,N_6627);
or U9913 (N_9913,N_7591,N_6412);
xnor U9914 (N_9914,N_8503,N_8613);
and U9915 (N_9915,N_8113,N_7203);
nor U9916 (N_9916,N_9264,N_7920);
nor U9917 (N_9917,N_7909,N_6560);
or U9918 (N_9918,N_6892,N_6532);
xor U9919 (N_9919,N_8586,N_8036);
nor U9920 (N_9920,N_8778,N_7000);
nand U9921 (N_9921,N_7931,N_7141);
xnor U9922 (N_9922,N_6671,N_6693);
xor U9923 (N_9923,N_7164,N_6635);
nor U9924 (N_9924,N_6925,N_7378);
and U9925 (N_9925,N_6547,N_8253);
or U9926 (N_9926,N_6380,N_6573);
nor U9927 (N_9927,N_6548,N_8285);
and U9928 (N_9928,N_8918,N_8423);
nor U9929 (N_9929,N_9137,N_6817);
and U9930 (N_9930,N_6333,N_9027);
or U9931 (N_9931,N_6792,N_6349);
nor U9932 (N_9932,N_7039,N_7976);
or U9933 (N_9933,N_7753,N_6878);
xor U9934 (N_9934,N_7144,N_8809);
xnor U9935 (N_9935,N_7472,N_8390);
nor U9936 (N_9936,N_6489,N_8751);
or U9937 (N_9937,N_8684,N_7598);
xor U9938 (N_9938,N_9163,N_7684);
and U9939 (N_9939,N_6806,N_6261);
and U9940 (N_9940,N_6325,N_6615);
xor U9941 (N_9941,N_8811,N_6920);
or U9942 (N_9942,N_8142,N_6762);
or U9943 (N_9943,N_6736,N_6456);
nand U9944 (N_9944,N_7841,N_8929);
nor U9945 (N_9945,N_8705,N_6914);
nand U9946 (N_9946,N_8888,N_8762);
nand U9947 (N_9947,N_7187,N_7803);
nor U9948 (N_9948,N_7607,N_6263);
nand U9949 (N_9949,N_8856,N_7299);
and U9950 (N_9950,N_6811,N_7407);
or U9951 (N_9951,N_7436,N_6771);
xnor U9952 (N_9952,N_8307,N_8074);
and U9953 (N_9953,N_8237,N_7277);
nand U9954 (N_9954,N_8092,N_9284);
nor U9955 (N_9955,N_8062,N_6551);
or U9956 (N_9956,N_8700,N_8043);
nand U9957 (N_9957,N_6363,N_8575);
and U9958 (N_9958,N_7376,N_9314);
nor U9959 (N_9959,N_6898,N_6365);
nand U9960 (N_9960,N_8246,N_6520);
nand U9961 (N_9961,N_8046,N_7668);
nand U9962 (N_9962,N_8987,N_8800);
and U9963 (N_9963,N_8268,N_7679);
and U9964 (N_9964,N_8972,N_8912);
or U9965 (N_9965,N_8655,N_8373);
xnor U9966 (N_9966,N_9287,N_7016);
nor U9967 (N_9967,N_8887,N_7575);
nor U9968 (N_9968,N_6258,N_7819);
nor U9969 (N_9969,N_7627,N_9151);
nand U9970 (N_9970,N_7088,N_8364);
and U9971 (N_9971,N_8254,N_6666);
nor U9972 (N_9972,N_8539,N_7796);
and U9973 (N_9973,N_8362,N_9229);
and U9974 (N_9974,N_8741,N_8352);
and U9975 (N_9975,N_6723,N_7623);
nand U9976 (N_9976,N_7902,N_8160);
xor U9977 (N_9977,N_8244,N_6592);
nor U9978 (N_9978,N_6522,N_6783);
nand U9979 (N_9979,N_8058,N_7794);
or U9980 (N_9980,N_7981,N_7032);
or U9981 (N_9981,N_7776,N_8151);
and U9982 (N_9982,N_9207,N_8069);
xor U9983 (N_9983,N_8050,N_7126);
and U9984 (N_9984,N_9063,N_7539);
or U9985 (N_9985,N_7214,N_8040);
or U9986 (N_9986,N_7295,N_8675);
or U9987 (N_9987,N_6975,N_8717);
or U9988 (N_9988,N_9099,N_8795);
and U9989 (N_9989,N_6688,N_8354);
or U9990 (N_9990,N_8432,N_7278);
or U9991 (N_9991,N_7763,N_6590);
or U9992 (N_9992,N_9373,N_7754);
nor U9993 (N_9993,N_6759,N_7932);
nand U9994 (N_9994,N_7261,N_8495);
xor U9995 (N_9995,N_8950,N_8505);
nand U9996 (N_9996,N_8681,N_8774);
nor U9997 (N_9997,N_6703,N_6705);
and U9998 (N_9998,N_8864,N_7593);
xor U9999 (N_9999,N_7616,N_9098);
and U10000 (N_10000,N_7887,N_7869);
and U10001 (N_10001,N_6387,N_7268);
nor U10002 (N_10002,N_7120,N_6256);
or U10003 (N_10003,N_9335,N_7462);
xor U10004 (N_10004,N_6285,N_8230);
or U10005 (N_10005,N_7510,N_6297);
nand U10006 (N_10006,N_7926,N_8671);
or U10007 (N_10007,N_6740,N_7077);
nor U10008 (N_10008,N_8485,N_6882);
and U10009 (N_10009,N_9248,N_6384);
or U10010 (N_10010,N_8103,N_7774);
and U10011 (N_10011,N_8152,N_9023);
and U10012 (N_10012,N_6620,N_8080);
nor U10013 (N_10013,N_7239,N_8897);
xnor U10014 (N_10014,N_6446,N_7496);
or U10015 (N_10015,N_8468,N_7617);
xor U10016 (N_10016,N_7934,N_8460);
and U10017 (N_10017,N_8218,N_7227);
nor U10018 (N_10018,N_8957,N_8188);
nand U10019 (N_10019,N_6462,N_7097);
nand U10020 (N_10020,N_8433,N_6845);
or U10021 (N_10021,N_8369,N_8614);
nand U10022 (N_10022,N_9368,N_7731);
and U10023 (N_10023,N_6569,N_6830);
and U10024 (N_10024,N_8379,N_7977);
nand U10025 (N_10025,N_8697,N_9357);
nor U10026 (N_10026,N_7222,N_7606);
xor U10027 (N_10027,N_7531,N_8745);
and U10028 (N_10028,N_8456,N_7612);
nor U10029 (N_10029,N_6600,N_8996);
xor U10030 (N_10030,N_6564,N_7614);
or U10031 (N_10031,N_8406,N_9010);
nor U10032 (N_10032,N_6468,N_7480);
xnor U10033 (N_10033,N_6471,N_8017);
nor U10034 (N_10034,N_8571,N_6883);
and U10035 (N_10035,N_8904,N_8115);
or U10036 (N_10036,N_7597,N_9064);
nor U10037 (N_10037,N_8175,N_9182);
nand U10038 (N_10038,N_7667,N_7235);
nand U10039 (N_10039,N_8501,N_7169);
nor U10040 (N_10040,N_6841,N_6734);
xnor U10041 (N_10041,N_8704,N_8298);
or U10042 (N_10042,N_8768,N_7134);
nor U10043 (N_10043,N_7848,N_8725);
nand U10044 (N_10044,N_6383,N_6524);
nand U10045 (N_10045,N_8759,N_8953);
nand U10046 (N_10046,N_7084,N_7915);
xnor U10047 (N_10047,N_8836,N_9032);
nor U10048 (N_10048,N_8547,N_6699);
nand U10049 (N_10049,N_7475,N_7028);
nor U10050 (N_10050,N_8020,N_7389);
and U10051 (N_10051,N_7952,N_9269);
nand U10052 (N_10052,N_9065,N_6582);
and U10053 (N_10053,N_7453,N_6701);
and U10054 (N_10054,N_9339,N_8698);
and U10055 (N_10055,N_8455,N_7625);
and U10056 (N_10056,N_7244,N_6949);
nand U10057 (N_10057,N_8942,N_8209);
nor U10058 (N_10058,N_6919,N_8258);
and U10059 (N_10059,N_8259,N_6946);
nand U10060 (N_10060,N_6943,N_9129);
and U10061 (N_10061,N_6578,N_7749);
xor U10062 (N_10062,N_9152,N_7008);
nor U10063 (N_10063,N_6683,N_7370);
or U10064 (N_10064,N_8344,N_6293);
nor U10065 (N_10065,N_8790,N_7738);
nand U10066 (N_10066,N_8569,N_9176);
xnor U10067 (N_10067,N_6903,N_8057);
nor U10068 (N_10068,N_6658,N_8528);
nand U10069 (N_10069,N_8772,N_6752);
and U10070 (N_10070,N_7839,N_7649);
xnor U10071 (N_10071,N_8331,N_7916);
nand U10072 (N_10072,N_6880,N_7127);
nor U10073 (N_10073,N_6345,N_8312);
nand U10074 (N_10074,N_7923,N_7192);
xnor U10075 (N_10075,N_9237,N_6368);
or U10076 (N_10076,N_7390,N_8223);
or U10077 (N_10077,N_6628,N_9150);
xor U10078 (N_10078,N_7698,N_6253);
or U10079 (N_10079,N_9185,N_8064);
nor U10080 (N_10080,N_7371,N_7246);
and U10081 (N_10081,N_8104,N_6499);
or U10082 (N_10082,N_8938,N_7391);
or U10083 (N_10083,N_9347,N_8990);
nand U10084 (N_10084,N_8986,N_6480);
or U10085 (N_10085,N_9345,N_8480);
nor U10086 (N_10086,N_8482,N_8065);
and U10087 (N_10087,N_7393,N_7166);
or U10088 (N_10088,N_7585,N_7913);
nor U10089 (N_10089,N_8911,N_6984);
nor U10090 (N_10090,N_8169,N_8011);
and U10091 (N_10091,N_6313,N_7517);
or U10092 (N_10092,N_8670,N_9060);
nand U10093 (N_10093,N_8314,N_9301);
and U10094 (N_10094,N_8696,N_6315);
nor U10095 (N_10095,N_7584,N_7680);
xor U10096 (N_10096,N_8674,N_9251);
xnor U10097 (N_10097,N_6436,N_9256);
and U10098 (N_10098,N_8758,N_6614);
and U10099 (N_10099,N_8176,N_8260);
and U10100 (N_10100,N_6838,N_7345);
nor U10101 (N_10101,N_7535,N_9074);
nor U10102 (N_10102,N_6802,N_8182);
nand U10103 (N_10103,N_8620,N_8465);
xor U10104 (N_10104,N_8186,N_8600);
and U10105 (N_10105,N_6381,N_6603);
or U10106 (N_10106,N_8625,N_7073);
or U10107 (N_10107,N_6624,N_6794);
xnor U10108 (N_10108,N_7647,N_8283);
nand U10109 (N_10109,N_8381,N_7810);
xor U10110 (N_10110,N_7891,N_8677);
or U10111 (N_10111,N_6299,N_6791);
nor U10112 (N_10112,N_7132,N_7989);
nor U10113 (N_10113,N_8412,N_7692);
xnor U10114 (N_10114,N_6358,N_8341);
nand U10115 (N_10115,N_8372,N_8163);
or U10116 (N_10116,N_8203,N_6400);
and U10117 (N_10117,N_6428,N_7281);
or U10118 (N_10118,N_7312,N_7631);
xor U10119 (N_10119,N_7081,N_6952);
nor U10120 (N_10120,N_7017,N_7757);
and U10121 (N_10121,N_9329,N_6901);
xnor U10122 (N_10122,N_8560,N_9059);
and U10123 (N_10123,N_8348,N_8619);
xnor U10124 (N_10124,N_6282,N_6978);
nand U10125 (N_10125,N_8949,N_6483);
xor U10126 (N_10126,N_7723,N_6382);
or U10127 (N_10127,N_6572,N_7336);
and U10128 (N_10128,N_6929,N_6554);
or U10129 (N_10129,N_9093,N_7961);
nor U10130 (N_10130,N_7789,N_6306);
or U10131 (N_10131,N_7563,N_6969);
or U10132 (N_10132,N_8633,N_7576);
or U10133 (N_10133,N_7971,N_8125);
or U10134 (N_10134,N_7090,N_7995);
xor U10135 (N_10135,N_8184,N_6605);
xor U10136 (N_10136,N_6529,N_7773);
xor U10137 (N_10137,N_7879,N_8073);
nor U10138 (N_10138,N_7076,N_6267);
nor U10139 (N_10139,N_6709,N_6941);
xnor U10140 (N_10140,N_8208,N_8850);
and U10141 (N_10141,N_6301,N_7912);
or U10142 (N_10142,N_8945,N_7595);
xnor U10143 (N_10143,N_8453,N_6593);
nand U10144 (N_10144,N_6977,N_8107);
and U10145 (N_10145,N_7502,N_9183);
nand U10146 (N_10146,N_7987,N_8787);
xnor U10147 (N_10147,N_7242,N_8166);
nor U10148 (N_10148,N_7359,N_6661);
nand U10149 (N_10149,N_7592,N_9333);
and U10150 (N_10150,N_7282,N_6405);
xnor U10151 (N_10151,N_9148,N_9195);
and U10152 (N_10152,N_8810,N_6747);
xor U10153 (N_10153,N_9313,N_6507);
nor U10154 (N_10154,N_9356,N_6327);
or U10155 (N_10155,N_8961,N_6728);
xor U10156 (N_10156,N_8537,N_7101);
nor U10157 (N_10157,N_8130,N_7291);
and U10158 (N_10158,N_7386,N_9147);
and U10159 (N_10159,N_6587,N_8027);
and U10160 (N_10160,N_6835,N_8822);
nor U10161 (N_10161,N_7189,N_6344);
and U10162 (N_10162,N_7054,N_8967);
and U10163 (N_10163,N_7940,N_7772);
xnor U10164 (N_10164,N_9157,N_7292);
or U10165 (N_10165,N_6818,N_9021);
nor U10166 (N_10166,N_9189,N_7665);
and U10167 (N_10167,N_6262,N_8646);
and U10168 (N_10168,N_8722,N_8866);
nand U10169 (N_10169,N_6542,N_9171);
xnor U10170 (N_10170,N_7818,N_8393);
nand U10171 (N_10171,N_8817,N_6485);
and U10172 (N_10172,N_7650,N_8541);
and U10173 (N_10173,N_7630,N_7975);
xnor U10174 (N_10174,N_6932,N_7174);
nor U10175 (N_10175,N_6970,N_8656);
or U10176 (N_10176,N_8324,N_7002);
or U10177 (N_10177,N_7644,N_9360);
or U10178 (N_10178,N_6250,N_7311);
or U10179 (N_10179,N_8231,N_8855);
xnor U10180 (N_10180,N_6757,N_6288);
nand U10181 (N_10181,N_9036,N_8602);
xnor U10182 (N_10182,N_8158,N_7458);
nor U10183 (N_10183,N_8279,N_7512);
or U10184 (N_10184,N_7938,N_7918);
nand U10185 (N_10185,N_7142,N_8044);
and U10186 (N_10186,N_9307,N_7170);
or U10187 (N_10187,N_9285,N_9057);
or U10188 (N_10188,N_8715,N_8955);
nand U10189 (N_10189,N_6591,N_8248);
and U10190 (N_10190,N_6745,N_7038);
nor U10191 (N_10191,N_8428,N_8149);
nand U10192 (N_10192,N_8720,N_7274);
xnor U10193 (N_10193,N_7823,N_9177);
nand U10194 (N_10194,N_6692,N_6496);
xnor U10195 (N_10195,N_9337,N_9198);
xor U10196 (N_10196,N_7707,N_6416);
nor U10197 (N_10197,N_7089,N_6378);
or U10198 (N_10198,N_6553,N_6664);
nor U10199 (N_10199,N_8333,N_8302);
nand U10200 (N_10200,N_7258,N_7124);
or U10201 (N_10201,N_7223,N_8740);
xnor U10202 (N_10202,N_8123,N_6955);
or U10203 (N_10203,N_8661,N_8576);
and U10204 (N_10204,N_8591,N_7908);
nand U10205 (N_10205,N_6887,N_7604);
nor U10206 (N_10206,N_8226,N_8118);
xor U10207 (N_10207,N_7309,N_8461);
nand U10208 (N_10208,N_8895,N_7886);
and U10209 (N_10209,N_6687,N_8678);
nand U10210 (N_10210,N_6807,N_8524);
or U10211 (N_10211,N_7876,N_8206);
nand U10212 (N_10212,N_8008,N_7373);
xnor U10213 (N_10213,N_8874,N_6633);
xor U10214 (N_10214,N_8479,N_6292);
nand U10215 (N_10215,N_7058,N_7993);
or U10216 (N_10216,N_7816,N_8716);
nor U10217 (N_10217,N_8487,N_8943);
nor U10218 (N_10218,N_8792,N_8245);
and U10219 (N_10219,N_6959,N_7885);
xnor U10220 (N_10220,N_8532,N_6821);
and U10221 (N_10221,N_8948,N_7963);
nor U10222 (N_10222,N_8514,N_8447);
nand U10223 (N_10223,N_8316,N_7352);
or U10224 (N_10224,N_8007,N_8066);
nor U10225 (N_10225,N_6490,N_9053);
xnor U10226 (N_10226,N_8294,N_6930);
and U10227 (N_10227,N_7655,N_6417);
xor U10228 (N_10228,N_6871,N_8598);
and U10229 (N_10229,N_6881,N_8081);
nand U10230 (N_10230,N_6571,N_8084);
xnor U10231 (N_10231,N_9126,N_8138);
or U10232 (N_10232,N_8356,N_9168);
or U10233 (N_10233,N_9049,N_9017);
nand U10234 (N_10234,N_8041,N_8517);
xnor U10235 (N_10235,N_9155,N_7750);
or U10236 (N_10236,N_8321,N_9283);
xnor U10237 (N_10237,N_8643,N_7477);
or U10238 (N_10238,N_8233,N_6785);
or U10239 (N_10239,N_8236,N_7421);
and U10240 (N_10240,N_9305,N_6799);
or U10241 (N_10241,N_7899,N_6550);
or U10242 (N_10242,N_7479,N_7457);
xnor U10243 (N_10243,N_8630,N_7237);
nand U10244 (N_10244,N_7632,N_6694);
nand U10245 (N_10245,N_9116,N_8126);
nor U10246 (N_10246,N_6894,N_7119);
nor U10247 (N_10247,N_9205,N_7368);
nor U10248 (N_10248,N_8770,N_8431);
nand U10249 (N_10249,N_7284,N_6423);
and U10250 (N_10250,N_8727,N_6364);
and U10251 (N_10251,N_8319,N_7316);
and U10252 (N_10252,N_8518,N_6991);
nor U10253 (N_10253,N_6738,N_9372);
xor U10254 (N_10254,N_6486,N_7253);
nand U10255 (N_10255,N_8927,N_8624);
xor U10256 (N_10256,N_7945,N_7335);
nor U10257 (N_10257,N_9088,N_7605);
xor U10258 (N_10258,N_8445,N_6931);
and U10259 (N_10259,N_8889,N_7791);
nand U10260 (N_10260,N_7557,N_7465);
xnor U10261 (N_10261,N_6340,N_9220);
xor U10262 (N_10262,N_7434,N_6639);
xnor U10263 (N_10263,N_8098,N_8402);
and U10264 (N_10264,N_7485,N_8615);
and U10265 (N_10265,N_7401,N_6951);
and U10266 (N_10266,N_7231,N_9184);
nor U10267 (N_10267,N_8540,N_6868);
and U10268 (N_10268,N_8694,N_9338);
xor U10269 (N_10269,N_6700,N_6294);
and U10270 (N_10270,N_9103,N_7863);
or U10271 (N_10271,N_8712,N_8146);
nor U10272 (N_10272,N_6689,N_8658);
and U10273 (N_10273,N_8567,N_8796);
xnor U10274 (N_10274,N_9082,N_9090);
xnor U10275 (N_10275,N_7555,N_7197);
or U10276 (N_10276,N_7527,N_9299);
or U10277 (N_10277,N_7898,N_6473);
xor U10278 (N_10278,N_8582,N_8414);
and U10279 (N_10279,N_7859,N_9238);
or U10280 (N_10280,N_7442,N_7779);
nor U10281 (N_10281,N_8049,N_7808);
and U10282 (N_10282,N_6475,N_8645);
or U10283 (N_10283,N_9241,N_9193);
or U10284 (N_10284,N_6623,N_7042);
nand U10285 (N_10285,N_7154,N_9223);
or U10286 (N_10286,N_7255,N_6290);
and U10287 (N_10287,N_8595,N_8791);
nand U10288 (N_10288,N_7202,N_7586);
nand U10289 (N_10289,N_8215,N_7568);
xor U10290 (N_10290,N_6272,N_8777);
nor U10291 (N_10291,N_8840,N_7396);
xor U10292 (N_10292,N_8472,N_7049);
nand U10293 (N_10293,N_8657,N_8276);
xnor U10294 (N_10294,N_9045,N_9131);
nand U10295 (N_10295,N_7232,N_9041);
xnor U10296 (N_10296,N_6990,N_6850);
xnor U10297 (N_10297,N_8930,N_8200);
or U10298 (N_10298,N_8892,N_6813);
nand U10299 (N_10299,N_7570,N_6445);
nor U10300 (N_10300,N_7363,N_8623);
nor U10301 (N_10301,N_9069,N_7635);
and U10302 (N_10302,N_7147,N_6466);
xor U10303 (N_10303,N_7986,N_6682);
nand U10304 (N_10304,N_7415,N_7086);
xnor U10305 (N_10305,N_7982,N_7340);
or U10306 (N_10306,N_8475,N_7003);
nor U10307 (N_10307,N_6576,N_8039);
or U10308 (N_10308,N_7459,N_6556);
xnor U10309 (N_10309,N_7666,N_9120);
or U10310 (N_10310,N_8886,N_7217);
nand U10311 (N_10311,N_7445,N_7348);
nand U10312 (N_10312,N_6410,N_9014);
and U10313 (N_10313,N_8335,N_8785);
nand U10314 (N_10314,N_8782,N_7759);
nor U10315 (N_10315,N_8639,N_8183);
xor U10316 (N_10316,N_8746,N_8555);
and U10317 (N_10317,N_6372,N_8797);
or U10318 (N_10318,N_6402,N_8180);
or U10319 (N_10319,N_7524,N_8689);
and U10320 (N_10320,N_7621,N_7021);
and U10321 (N_10321,N_8100,N_8580);
nand U10322 (N_10322,N_7082,N_7775);
nand U10323 (N_10323,N_9218,N_7495);
nand U10324 (N_10324,N_7157,N_8037);
and U10325 (N_10325,N_6753,N_8579);
nor U10326 (N_10326,N_6879,N_6998);
xnor U10327 (N_10327,N_8112,N_8477);
and U10328 (N_10328,N_8366,N_7079);
nand U10329 (N_10329,N_6425,N_8139);
nor U10330 (N_10330,N_7691,N_6393);
nor U10331 (N_10331,N_8593,N_8898);
nand U10332 (N_10332,N_7726,N_7740);
nand U10333 (N_10333,N_6455,N_8308);
nand U10334 (N_10334,N_6602,N_6966);
and U10335 (N_10335,N_9044,N_6915);
and U10336 (N_10336,N_8531,N_8709);
nand U10337 (N_10337,N_6672,N_9070);
and U10338 (N_10338,N_7379,N_7324);
xnor U10339 (N_10339,N_9328,N_7168);
or U10340 (N_10340,N_6434,N_9366);
or U10341 (N_10341,N_7696,N_6580);
and U10342 (N_10342,N_6686,N_7732);
nand U10343 (N_10343,N_8919,N_8504);
and U10344 (N_10344,N_8131,N_8448);
and U10345 (N_10345,N_6824,N_7484);
nor U10346 (N_10346,N_6815,N_9092);
nand U10347 (N_10347,N_6374,N_7233);
nand U10348 (N_10348,N_6721,N_7967);
or U10349 (N_10349,N_9113,N_9025);
or U10350 (N_10350,N_7559,N_8622);
nand U10351 (N_10351,N_6369,N_9187);
nand U10352 (N_10352,N_9212,N_7733);
nand U10353 (N_10353,N_9350,N_6426);
nand U10354 (N_10354,N_8841,N_7542);
or U10355 (N_10355,N_6775,N_9304);
or U10356 (N_10356,N_8820,N_9192);
xnor U10357 (N_10357,N_8034,N_7672);
or U10358 (N_10358,N_6685,N_8621);
xnor U10359 (N_10359,N_6414,N_6563);
and U10360 (N_10360,N_9115,N_8828);
and U10361 (N_10361,N_9075,N_8915);
xnor U10362 (N_10362,N_7146,N_7100);
nand U10363 (N_10363,N_7947,N_8419);
nor U10364 (N_10364,N_6334,N_7550);
and U10365 (N_10365,N_9211,N_9179);
and U10366 (N_10366,N_7497,N_8359);
and U10367 (N_10367,N_7736,N_9068);
nand U10368 (N_10368,N_7856,N_8925);
nor U10369 (N_10369,N_6375,N_7653);
nor U10370 (N_10370,N_7114,N_8739);
nor U10371 (N_10371,N_7104,N_8966);
nor U10372 (N_10372,N_7636,N_8410);
nand U10373 (N_10373,N_8085,N_8859);
and U10374 (N_10374,N_8249,N_8264);
xor U10375 (N_10375,N_8177,N_7014);
nand U10376 (N_10376,N_9232,N_8153);
nor U10377 (N_10377,N_8711,N_6442);
or U10378 (N_10378,N_6534,N_7618);
xnor U10379 (N_10379,N_7968,N_6303);
nand U10380 (N_10380,N_7302,N_6415);
or U10381 (N_10381,N_6575,N_6503);
xor U10382 (N_10382,N_8771,N_8063);
nor U10383 (N_10383,N_9108,N_7419);
and U10384 (N_10384,N_8629,N_6819);
and U10385 (N_10385,N_8733,N_7159);
nand U10386 (N_10386,N_7602,N_7023);
nor U10387 (N_10387,N_7864,N_6668);
and U10388 (N_10388,N_7526,N_9006);
and U10389 (N_10389,N_8626,N_8243);
nand U10390 (N_10390,N_7301,N_6616);
and U10391 (N_10391,N_9094,N_7064);
and U10392 (N_10392,N_6844,N_8003);
and U10393 (N_10393,N_7115,N_8516);
nor U10394 (N_10394,N_9352,N_8289);
nor U10395 (N_10395,N_8240,N_6861);
nor U10396 (N_10396,N_7639,N_7405);
nand U10397 (N_10397,N_7355,N_7874);
and U10398 (N_10398,N_7112,N_7536);
and U10399 (N_10399,N_7582,N_7827);
xor U10400 (N_10400,N_8108,N_6598);
or U10401 (N_10401,N_7098,N_7105);
xnor U10402 (N_10402,N_8664,N_7683);
nor U10403 (N_10403,N_7160,N_8703);
or U10404 (N_10404,N_8783,N_9312);
or U10405 (N_10405,N_8676,N_8806);
nor U10406 (N_10406,N_6852,N_6361);
and U10407 (N_10407,N_6463,N_6945);
and U10408 (N_10408,N_9278,N_8702);
xor U10409 (N_10409,N_8737,N_6665);
and U10410 (N_10410,N_9029,N_9228);
and U10411 (N_10411,N_9316,N_9217);
and U10412 (N_10412,N_6509,N_7950);
and U10413 (N_10413,N_6948,N_7800);
xnor U10414 (N_10414,N_8554,N_8688);
and U10415 (N_10415,N_6317,N_8205);
and U10416 (N_10416,N_8016,N_8165);
nor U10417 (N_10417,N_7056,N_8273);
xor U10418 (N_10418,N_6362,N_8263);
and U10419 (N_10419,N_8051,N_8500);
and U10420 (N_10420,N_8096,N_7337);
or U10421 (N_10421,N_9020,N_6778);
nor U10422 (N_10422,N_7673,N_8843);
nand U10423 (N_10423,N_8295,N_8871);
nor U10424 (N_10424,N_7085,N_7403);
nand U10425 (N_10425,N_8212,N_6309);
and U10426 (N_10426,N_8520,N_8159);
nor U10427 (N_10427,N_7347,N_9046);
nand U10428 (N_10428,N_7553,N_8507);
nand U10429 (N_10429,N_9140,N_6712);
xnor U10430 (N_10430,N_8493,N_6916);
and U10431 (N_10431,N_7717,N_9254);
xor U10432 (N_10432,N_8137,N_6715);
or U10433 (N_10433,N_6754,N_7285);
or U10434 (N_10434,N_8561,N_7071);
nand U10435 (N_10435,N_8563,N_8086);
or U10436 (N_10436,N_7045,N_6398);
nor U10437 (N_10437,N_7448,N_8116);
nor U10438 (N_10438,N_6422,N_9085);
and U10439 (N_10439,N_9127,N_7010);
nand U10440 (N_10440,N_6823,N_6996);
and U10441 (N_10441,N_8848,N_8847);
xnor U10442 (N_10442,N_6803,N_6467);
and U10443 (N_10443,N_6488,N_7880);
xnor U10444 (N_10444,N_7009,N_7471);
nor U10445 (N_10445,N_8908,N_7411);
or U10446 (N_10446,N_7331,N_9118);
and U10447 (N_10447,N_9343,N_8132);
nor U10448 (N_10448,N_9173,N_7735);
nand U10449 (N_10449,N_7615,N_7770);
xor U10450 (N_10450,N_6972,N_8185);
and U10451 (N_10451,N_7608,N_6377);
and U10452 (N_10452,N_7467,N_8901);
or U10453 (N_10453,N_7645,N_7351);
or U10454 (N_10454,N_9281,N_8091);
nor U10455 (N_10455,N_7319,N_8685);
nand U10456 (N_10456,N_7581,N_8565);
or U10457 (N_10457,N_8251,N_7343);
or U10458 (N_10458,N_8508,N_8971);
and U10459 (N_10459,N_8804,N_6918);
or U10460 (N_10460,N_7894,N_8386);
nand U10461 (N_10461,N_6676,N_6487);
xor U10462 (N_10462,N_6265,N_6413);
xor U10463 (N_10463,N_9322,N_8403);
xor U10464 (N_10464,N_8562,N_7969);
or U10465 (N_10465,N_8881,N_7075);
or U10466 (N_10466,N_8374,N_8997);
xor U10467 (N_10467,N_9215,N_8708);
nor U10468 (N_10468,N_7432,N_8764);
or U10469 (N_10469,N_7722,N_8054);
nor U10470 (N_10470,N_7397,N_7270);
nand U10471 (N_10471,N_8896,N_8729);
nand U10472 (N_10472,N_6619,N_6625);
and U10473 (N_10473,N_6954,N_8277);
nand U10474 (N_10474,N_8394,N_7601);
nand U10475 (N_10475,N_7997,N_8909);
xnor U10476 (N_10476,N_7676,N_8946);
and U10477 (N_10477,N_8015,N_9208);
and U10478 (N_10478,N_7783,N_8491);
and U10479 (N_10479,N_9031,N_7533);
or U10480 (N_10480,N_8730,N_8603);
xnor U10481 (N_10481,N_7752,N_6476);
xnor U10482 (N_10482,N_7374,N_8145);
nor U10483 (N_10483,N_8315,N_7451);
nor U10484 (N_10484,N_7228,N_9083);
and U10485 (N_10485,N_9102,N_8476);
nand U10486 (N_10486,N_9153,N_8857);
nor U10487 (N_10487,N_6622,N_8799);
nand U10488 (N_10488,N_6330,N_8216);
nand U10489 (N_10489,N_8071,N_7642);
nand U10490 (N_10490,N_8680,N_7290);
xnor U10491 (N_10491,N_6343,N_9371);
xnor U10492 (N_10492,N_7423,N_7521);
nor U10493 (N_10493,N_9270,N_9117);
or U10494 (N_10494,N_6690,N_7675);
xnor U10495 (N_10495,N_7007,N_7240);
or U10496 (N_10496,N_8099,N_6385);
nand U10497 (N_10497,N_9009,N_6491);
or U10498 (N_10498,N_7070,N_8763);
xnor U10499 (N_10499,N_7323,N_7659);
and U10500 (N_10500,N_6640,N_9091);
and U10501 (N_10501,N_9112,N_7303);
nor U10502 (N_10502,N_7030,N_7110);
nand U10503 (N_10503,N_6538,N_8975);
or U10504 (N_10504,N_9144,N_7304);
xnor U10505 (N_10505,N_8584,N_8122);
nor U10506 (N_10506,N_6621,N_9000);
nor U10507 (N_10507,N_6251,N_6854);
xnor U10508 (N_10508,N_9200,N_6336);
nor U10509 (N_10509,N_8637,N_8094);
or U10510 (N_10510,N_6869,N_7433);
and U10511 (N_10511,N_7702,N_9213);
and U10512 (N_10512,N_9289,N_6924);
nor U10513 (N_10513,N_9178,N_9095);
nand U10514 (N_10514,N_7380,N_8928);
xor U10515 (N_10515,N_7669,N_6997);
nor U10516 (N_10516,N_9268,N_9174);
nand U10517 (N_10517,N_8732,N_6508);
nand U10518 (N_10518,N_7041,N_7243);
and U10519 (N_10519,N_7739,N_6893);
xor U10520 (N_10520,N_7326,N_7297);
or U10521 (N_10521,N_7296,N_8581);
nand U10522 (N_10522,N_8235,N_8157);
or U10523 (N_10523,N_8101,N_7382);
nor U10524 (N_10524,N_8070,N_7806);
or U10525 (N_10525,N_7519,N_8181);
nand U10526 (N_10526,N_8342,N_9318);
and U10527 (N_10527,N_6431,N_7507);
or U10528 (N_10528,N_8415,N_8031);
and U10529 (N_10529,N_9047,N_8749);
or U10530 (N_10530,N_8140,N_9076);
xor U10531 (N_10531,N_8052,N_6760);
or U10532 (N_10532,N_9288,N_6981);
xnor U10533 (N_10533,N_6963,N_7454);
nor U10534 (N_10534,N_6782,N_7873);
nand U10535 (N_10535,N_7892,N_8825);
nor U10536 (N_10536,N_8417,N_9315);
and U10537 (N_10537,N_7883,N_8471);
nand U10538 (N_10538,N_9253,N_8161);
nand U10539 (N_10539,N_9043,N_8510);
nand U10540 (N_10540,N_8920,N_6595);
or U10541 (N_10541,N_8601,N_9096);
nor U10542 (N_10542,N_7824,N_8756);
and U10543 (N_10543,N_8564,N_7766);
xnor U10544 (N_10544,N_8030,N_7629);
nand U10545 (N_10545,N_7140,N_7490);
and U10546 (N_10546,N_9222,N_7514);
nand U10547 (N_10547,N_9310,N_7024);
nor U10548 (N_10548,N_7280,N_6296);
or U10549 (N_10549,N_9204,N_8845);
or U10550 (N_10550,N_7674,N_6926);
xnor U10551 (N_10551,N_6704,N_9097);
or U10552 (N_10552,N_8378,N_8033);
or U10553 (N_10553,N_7207,N_7230);
and U10554 (N_10554,N_7654,N_7509);
or U10555 (N_10555,N_7412,N_8549);
or U10556 (N_10556,N_7198,N_7254);
nor U10557 (N_10557,N_8266,N_6906);
nor U10558 (N_10558,N_7624,N_6539);
nand U10559 (N_10559,N_8882,N_8970);
nor U10560 (N_10560,N_8568,N_7701);
nor U10561 (N_10561,N_6348,N_6765);
or U10562 (N_10562,N_8087,N_7406);
xnor U10563 (N_10563,N_9191,N_8934);
xor U10564 (N_10564,N_8983,N_7540);
or U10565 (N_10565,N_7965,N_6634);
nor U10566 (N_10566,N_7173,N_7785);
xnor U10567 (N_10567,N_6743,N_6281);
xor U10568 (N_10568,N_9374,N_6335);
nor U10569 (N_10569,N_8488,N_9133);
and U10570 (N_10570,N_6891,N_8300);
and U10571 (N_10571,N_6568,N_8802);
and U10572 (N_10572,N_6429,N_7185);
nor U10573 (N_10573,N_7843,N_8127);
or U10574 (N_10574,N_7330,N_6810);
nand U10575 (N_10575,N_8318,N_8265);
nor U10576 (N_10576,N_7435,N_8765);
or U10577 (N_10577,N_6521,N_9296);
xor U10578 (N_10578,N_8873,N_7439);
or U10579 (N_10579,N_6675,N_8155);
or U10580 (N_10580,N_6989,N_8963);
xnor U10581 (N_10581,N_6607,N_8463);
xnor U10582 (N_10582,N_7289,N_7179);
nand U10583 (N_10583,N_9247,N_7664);
or U10584 (N_10584,N_6498,N_8965);
and U10585 (N_10585,N_6670,N_6492);
nor U10586 (N_10586,N_8789,N_8061);
or U10587 (N_10587,N_6537,N_6320);
nand U10588 (N_10588,N_8021,N_7573);
or U10589 (N_10589,N_7719,N_7107);
xor U10590 (N_10590,N_8095,N_6899);
or U10591 (N_10591,N_8025,N_6404);
xnor U10592 (N_10592,N_6921,N_7440);
nand U10593 (N_10593,N_6902,N_8995);
nor U10594 (N_10594,N_6982,N_9015);
and U10595 (N_10595,N_6518,N_9367);
nor U10596 (N_10596,N_7219,N_6927);
and U10597 (N_10597,N_7812,N_6940);
or U10598 (N_10598,N_9358,N_6495);
xnor U10599 (N_10599,N_8377,N_8221);
xnor U10600 (N_10600,N_7960,N_7525);
or U10601 (N_10601,N_7697,N_7984);
and U10602 (N_10602,N_7275,N_6601);
nor U10603 (N_10603,N_8309,N_7651);
xor U10604 (N_10604,N_9342,N_7191);
nor U10605 (N_10605,N_9051,N_9109);
or U10606 (N_10606,N_9249,N_8631);
nand U10607 (N_10607,N_7837,N_7482);
nor U10608 (N_10608,N_8196,N_9001);
xor U10609 (N_10609,N_7360,N_6505);
or U10610 (N_10610,N_6856,N_6904);
and U10611 (N_10611,N_7377,N_8906);
and U10612 (N_10612,N_6257,N_6983);
or U10613 (N_10613,N_8239,N_8529);
or U10614 (N_10614,N_6324,N_8055);
nor U10615 (N_10615,N_7755,N_6370);
or U10616 (N_10616,N_6304,N_8201);
nand U10617 (N_10617,N_6663,N_6545);
nor U10618 (N_10618,N_6912,N_6321);
xnor U10619 (N_10619,N_6482,N_6777);
or U10620 (N_10620,N_7980,N_7877);
and U10621 (N_10621,N_7103,N_7062);
nor U10622 (N_10622,N_8659,N_7867);
nand U10623 (N_10623,N_8776,N_6708);
nor U10624 (N_10624,N_8005,N_7620);
nor U10625 (N_10625,N_9219,N_6474);
nor U10626 (N_10626,N_6606,N_7516);
or U10627 (N_10627,N_7300,N_8407);
nand U10628 (N_10628,N_7057,N_7092);
xor U10629 (N_10629,N_8742,N_8009);
xnor U10630 (N_10630,N_7314,N_6540);
xor U10631 (N_10631,N_7367,N_7491);
xor U10632 (N_10632,N_7059,N_6710);
or U10633 (N_10633,N_8734,N_7815);
nor U10634 (N_10634,N_9154,N_6449);
xnor U10635 (N_10635,N_7151,N_6788);
nand U10636 (N_10636,N_6409,N_7066);
xnor U10637 (N_10637,N_7588,N_7437);
and U10638 (N_10638,N_7998,N_8826);
nand U10639 (N_10639,N_8396,N_9309);
xor U10640 (N_10640,N_6750,N_8077);
xor U10641 (N_10641,N_8808,N_7156);
xnor U10642 (N_10642,N_8128,N_8985);
nor U10643 (N_10643,N_7648,N_8442);
and U10644 (N_10644,N_8336,N_7713);
or U10645 (N_10645,N_7786,N_9242);
nand U10646 (N_10646,N_6298,N_7438);
nor U10647 (N_10647,N_8982,N_9028);
nand U10648 (N_10648,N_8392,N_6549);
xor U10649 (N_10649,N_6751,N_7498);
nor U10650 (N_10650,N_9121,N_6895);
and U10651 (N_10651,N_8923,N_8761);
xor U10652 (N_10652,N_8662,N_9221);
nor U10653 (N_10653,N_9022,N_8224);
nor U10654 (N_10654,N_7026,N_6855);
nand U10655 (N_10655,N_8202,N_6836);
nor U10656 (N_10656,N_8947,N_8723);
nand U10657 (N_10657,N_7329,N_8824);
xor U10658 (N_10658,N_7907,N_8361);
and U10659 (N_10659,N_7685,N_7139);
and U10660 (N_10660,N_7663,N_7046);
nor U10661 (N_10661,N_8358,N_9300);
xor U10662 (N_10662,N_9055,N_7422);
or U10663 (N_10663,N_6570,N_7737);
nor U10664 (N_10664,N_7992,N_9172);
xnor U10665 (N_10665,N_7957,N_6849);
and U10666 (N_10666,N_7882,N_8337);
xor U10667 (N_10667,N_6420,N_7190);
xnor U10668 (N_10668,N_6876,N_7418);
and U10669 (N_10669,N_6647,N_9164);
or U10670 (N_10670,N_6531,N_8654);
or U10671 (N_10671,N_8179,N_7501);
nand U10672 (N_10672,N_7196,N_7782);
xnor U10673 (N_10673,N_6834,N_9052);
or U10674 (N_10674,N_7634,N_8917);
xnor U10675 (N_10675,N_8515,N_7858);
nand U10676 (N_10676,N_8900,N_7734);
nor U10677 (N_10677,N_8262,N_8640);
or U10678 (N_10678,N_8635,N_6857);
xnor U10679 (N_10679,N_8883,N_9369);
and U10680 (N_10680,N_7781,N_7155);
nand U10681 (N_10681,N_8397,N_6276);
nor U10682 (N_10682,N_8876,N_7919);
nor U10683 (N_10683,N_7549,N_7881);
nand U10684 (N_10684,N_8291,N_7325);
or U10685 (N_10685,N_9203,N_7518);
nor U10686 (N_10686,N_7224,N_7792);
xnor U10687 (N_10687,N_7375,N_7063);
nand U10688 (N_10688,N_6406,N_9101);
or U10689 (N_10689,N_9181,N_7346);
or U10690 (N_10690,N_9216,N_9292);
xnor U10691 (N_10691,N_8441,N_8590);
and U10692 (N_10692,N_7560,N_6459);
or U10693 (N_10693,N_6864,N_7790);
xnor U10694 (N_10694,N_8317,N_9105);
and U10695 (N_10695,N_7213,N_8607);
or U10696 (N_10696,N_8832,N_6589);
nand U10697 (N_10697,N_7548,N_9180);
or U10698 (N_10698,N_6828,N_7532);
xor U10699 (N_10699,N_9326,N_8422);
xor U10700 (N_10700,N_7113,N_8954);
xnor U10701 (N_10701,N_8522,N_8819);
nor U10702 (N_10702,N_8042,N_8933);
and U10703 (N_10703,N_6617,N_7102);
nand U10704 (N_10704,N_8974,N_8299);
or U10705 (N_10705,N_7094,N_6908);
or U10706 (N_10706,N_6846,N_7637);
and U10707 (N_10707,N_8821,N_7399);
or U10708 (N_10708,N_8088,N_6822);
and U10709 (N_10709,N_7165,N_6847);
nor U10710 (N_10710,N_6318,N_9353);
xor U10711 (N_10711,N_6840,N_9073);
nand U10712 (N_10712,N_8222,N_7930);
or U10713 (N_10713,N_7758,N_7229);
nand U10714 (N_10714,N_7199,N_7332);
and U10715 (N_10715,N_8458,N_7552);
or U10716 (N_10716,N_8330,N_7356);
nand U10717 (N_10717,N_6386,N_7788);
and U10718 (N_10718,N_9340,N_9079);
xor U10719 (N_10719,N_6427,N_8023);
xor U10720 (N_10720,N_7385,N_6910);
nand U10721 (N_10721,N_7860,N_7523);
nor U10722 (N_10722,N_8006,N_7936);
and U10723 (N_10723,N_7044,N_7513);
nand U10724 (N_10724,N_7569,N_7822);
nor U10725 (N_10725,N_7183,N_6399);
xor U10726 (N_10726,N_8004,N_7452);
nor U10727 (N_10727,N_7135,N_8861);
or U10728 (N_10728,N_8404,N_9257);
and U10729 (N_10729,N_9081,N_7688);
nand U10730 (N_10730,N_6510,N_9135);
and U10731 (N_10731,N_7694,N_8451);
and U10732 (N_10732,N_8588,N_9202);
xnor U10733 (N_10733,N_7508,N_7690);
nor U10734 (N_10734,N_7129,N_9279);
xnor U10735 (N_10735,N_7866,N_7579);
nand U10736 (N_10736,N_8862,N_8119);
and U10737 (N_10737,N_7949,N_6566);
nor U10738 (N_10738,N_8589,N_9267);
nor U10739 (N_10739,N_8952,N_8610);
or U10740 (N_10740,N_6993,N_9040);
or U10741 (N_10741,N_6439,N_8879);
xor U10742 (N_10742,N_7983,N_6833);
nand U10743 (N_10743,N_7381,N_9262);
nand U10744 (N_10744,N_7834,N_7703);
xor U10745 (N_10745,N_8421,N_6526);
or U10746 (N_10746,N_6917,N_9252);
or U10747 (N_10747,N_7662,N_6567);
xnor U10748 (N_10748,N_9125,N_7922);
xnor U10749 (N_10749,N_7730,N_7712);
and U10750 (N_10750,N_8687,N_9332);
nand U10751 (N_10751,N_7006,N_8191);
nor U10752 (N_10752,N_7180,N_6255);
and U10753 (N_10753,N_7567,N_7167);
xnor U10754 (N_10754,N_7937,N_8353);
or U10755 (N_10755,N_8192,N_8533);
nand U10756 (N_10756,N_7910,N_7681);
nor U10757 (N_10757,N_6681,N_7778);
and U10758 (N_10758,N_9134,N_6494);
or U10759 (N_10759,N_7333,N_8837);
or U10760 (N_10760,N_7978,N_6730);
nand U10761 (N_10761,N_8425,N_8198);
or U10762 (N_10762,N_7990,N_7069);
xnor U10763 (N_10763,N_6516,N_9260);
or U10764 (N_10764,N_8168,N_8587);
nor U10765 (N_10765,N_7814,N_8877);
xnor U10766 (N_10766,N_8512,N_6342);
xor U10767 (N_10767,N_7149,N_9186);
and U10768 (N_10768,N_8371,N_7162);
nor U10769 (N_10769,N_7052,N_8916);
xnor U10770 (N_10770,N_8492,N_6829);
nor U10771 (N_10771,N_7587,N_7805);
and U10772 (N_10772,N_9199,N_7613);
nor U10773 (N_10773,N_7744,N_7492);
nand U10774 (N_10774,N_8000,N_6911);
nand U10775 (N_10775,N_7900,N_7388);
xnor U10776 (N_10776,N_6557,N_7609);
nor U10777 (N_10777,N_6525,N_6731);
and U10778 (N_10778,N_6886,N_6877);
xnor U10779 (N_10779,N_9111,N_7836);
or U10780 (N_10780,N_6360,N_8284);
nor U10781 (N_10781,N_8347,N_8256);
or U10782 (N_10782,N_7528,N_7394);
xor U10783 (N_10783,N_8693,N_9024);
or U10784 (N_10784,N_8899,N_9286);
or U10785 (N_10785,N_7745,N_7461);
xor U10786 (N_10786,N_9233,N_7693);
xnor U10787 (N_10787,N_7091,N_7040);
nand U10788 (N_10788,N_6594,N_6784);
and U10789 (N_10789,N_8217,N_7769);
or U10790 (N_10790,N_8444,N_8102);
nor U10791 (N_10791,N_7925,N_7257);
nand U10792 (N_10792,N_9244,N_8556);
nand U10793 (N_10793,N_7890,N_8769);
or U10794 (N_10794,N_7108,N_7486);
nor U10795 (N_10795,N_8405,N_6727);
or U10796 (N_10796,N_7384,N_9190);
nand U10797 (N_10797,N_6636,N_7924);
nand U10798 (N_10798,N_6354,N_6444);
nor U10799 (N_10799,N_6269,N_7771);
nand U10800 (N_10800,N_7035,N_9159);
nand U10801 (N_10801,N_6464,N_6680);
nand U10802 (N_10802,N_8282,N_7804);
nor U10803 (N_10803,N_7321,N_9196);
xor U10804 (N_10804,N_9243,N_7456);
and U10805 (N_10805,N_8490,N_8860);
xnor U10806 (N_10806,N_8280,N_8286);
or U10807 (N_10807,N_8343,N_6631);
xnor U10808 (N_10808,N_7832,N_9306);
or U10809 (N_10809,N_6816,N_7414);
nor U10810 (N_10810,N_8984,N_8867);
nand U10811 (N_10811,N_8474,N_6559);
nand U10812 (N_10812,N_7801,N_7633);
xnor U10813 (N_10813,N_7055,N_6511);
xnor U10814 (N_10814,N_9030,N_8261);
or U10815 (N_10815,N_9298,N_7215);
xnor U10816 (N_10816,N_7914,N_7720);
and U10817 (N_10817,N_6611,N_6796);
nor U10818 (N_10818,N_6391,N_6584);
or U10819 (N_10819,N_8706,N_7468);
nand U10820 (N_10820,N_6307,N_7838);
xor U10821 (N_10821,N_6535,N_8902);
nor U10822 (N_10822,N_7853,N_7250);
xor U10823 (N_10823,N_9042,N_7728);
nor U10824 (N_10824,N_7449,N_7447);
xnor U10825 (N_10825,N_6789,N_7096);
and U10826 (N_10826,N_6641,N_7131);
xor U10827 (N_10827,N_8322,N_6461);
xnor U10828 (N_10828,N_6942,N_6457);
and U10829 (N_10829,N_8536,N_8497);
or U10830 (N_10830,N_8255,N_6957);
or U10831 (N_10831,N_8032,N_6717);
or U10832 (N_10832,N_8467,N_8981);
xor U10833 (N_10833,N_8718,N_8328);
nor U10834 (N_10834,N_9146,N_7417);
nand U10835 (N_10835,N_6259,N_7842);
xor U10836 (N_10836,N_8724,N_8574);
and U10837 (N_10837,N_7751,N_6517);
xnor U10838 (N_10838,N_7742,N_8999);
xor U10839 (N_10839,N_9194,N_7817);
xnor U10840 (N_10840,N_8435,N_7833);
nand U10841 (N_10841,N_6448,N_6350);
nor U10842 (N_10842,N_8543,N_7985);
nor U10843 (N_10843,N_8252,N_8513);
or U10844 (N_10844,N_8187,N_8489);
nand U10845 (N_10845,N_8454,N_6561);
nand U10846 (N_10846,N_7670,N_6287);
or U10847 (N_10847,N_8679,N_6470);
nor U10848 (N_10848,N_8067,N_6711);
nand U10849 (N_10849,N_7068,N_8350);
xor U10850 (N_10850,N_7515,N_7029);
nand U10851 (N_10851,N_8530,N_7928);
nor U10852 (N_10852,N_9364,N_8078);
or U10853 (N_10853,N_8136,N_6479);
xor U10854 (N_10854,N_7218,N_8652);
and U10855 (N_10855,N_9348,N_8682);
nor U10856 (N_10856,N_6755,N_9341);
and U10857 (N_10857,N_7956,N_8699);
and U10858 (N_10858,N_8551,N_8572);
and U10859 (N_10859,N_8519,N_7204);
xor U10860 (N_10860,N_7896,N_6994);
nor U10861 (N_10861,N_6421,N_6964);
and U10862 (N_10862,N_9263,N_8865);
and U10863 (N_10863,N_9227,N_8618);
and U10864 (N_10864,N_8452,N_8093);
and U10865 (N_10865,N_6986,N_6355);
and U10866 (N_10866,N_7072,N_6875);
or U10867 (N_10867,N_6326,N_8135);
nor U10868 (N_10868,N_7660,N_6527);
nor U10869 (N_10869,N_8195,N_7895);
or U10870 (N_10870,N_7878,N_9250);
and U10871 (N_10871,N_7357,N_6401);
nand U10872 (N_10872,N_8893,N_9169);
or U10873 (N_10873,N_8638,N_7917);
or U10874 (N_10874,N_8535,N_8257);
or U10875 (N_10875,N_6637,N_7428);
nor U10876 (N_10876,N_8349,N_9104);
or U10877 (N_10877,N_8368,N_8527);
xor U10878 (N_10878,N_7748,N_8632);
and U10879 (N_10879,N_8199,N_8903);
nand U10880 (N_10880,N_8666,N_8013);
xor U10881 (N_10881,N_7037,N_6252);
nor U10882 (N_10882,N_6722,N_7234);
xor U10883 (N_10883,N_6254,N_7829);
and U10884 (N_10884,N_7994,N_6909);
nor U10885 (N_10885,N_9067,N_9362);
or U10886 (N_10886,N_8818,N_6543);
nand U10887 (N_10887,N_7811,N_7677);
xor U10888 (N_10888,N_8827,N_6438);
or U10889 (N_10889,N_9062,N_8858);
and U10890 (N_10890,N_8197,N_6962);
nand U10891 (N_10891,N_6275,N_8029);
or U10892 (N_10892,N_8559,N_8939);
or U10893 (N_10893,N_8437,N_7317);
xor U10894 (N_10894,N_7248,N_7504);
nand U10895 (N_10895,N_8839,N_6786);
or U10896 (N_10896,N_9327,N_8247);
or U10897 (N_10897,N_8844,N_8400);
nand U10898 (N_10898,N_7210,N_7095);
xnor U10899 (N_10899,N_6352,N_7206);
and U10900 (N_10900,N_7845,N_6392);
nor U10901 (N_10901,N_6729,N_8219);
nand U10902 (N_10902,N_9274,N_6713);
nor U10903 (N_10903,N_8669,N_9078);
and U10904 (N_10904,N_7661,N_9019);
nor U10905 (N_10905,N_6277,N_8690);
xnor U10906 (N_10906,N_7426,N_7339);
or U10907 (N_10907,N_6873,N_8418);
and U10908 (N_10908,N_8653,N_7825);
and U10909 (N_10909,N_6323,N_7541);
or U10910 (N_10910,N_6403,N_6289);
nor U10911 (N_10911,N_6937,N_8389);
xor U10912 (N_10912,N_6314,N_8628);
xnor U10913 (N_10913,N_7034,N_9235);
or U10914 (N_10914,N_6679,N_7657);
nand U10915 (N_10915,N_6960,N_6359);
nand U10916 (N_10916,N_9002,N_8921);
and U10917 (N_10917,N_7487,N_8870);
nor U10918 (N_10918,N_8469,N_7182);
nor U10919 (N_10919,N_6376,N_8339);
xor U10920 (N_10920,N_8606,N_7344);
nand U10921 (N_10921,N_8124,N_7793);
xnor U10922 (N_10922,N_7714,N_6988);
and U10923 (N_10923,N_8502,N_7973);
nor U10924 (N_10924,N_6758,N_6366);
or U10925 (N_10925,N_8401,N_9231);
and U10926 (N_10926,N_7283,N_9138);
nand U10927 (N_10927,N_6268,N_9087);
nand U10928 (N_10928,N_7306,N_8775);
nand U10929 (N_10929,N_9033,N_7828);
nor U10930 (N_10930,N_8868,N_8558);
or U10931 (N_10931,N_7116,N_7031);
and U10932 (N_10932,N_6673,N_7444);
and U10933 (N_10933,N_8363,N_8885);
and U10934 (N_10934,N_9224,N_7163);
xnor U10935 (N_10935,N_8506,N_8449);
and U10936 (N_10936,N_8760,N_7404);
nand U10937 (N_10937,N_7338,N_7353);
and U10938 (N_10938,N_7356,N_8084);
and U10939 (N_10939,N_8422,N_7334);
and U10940 (N_10940,N_7494,N_7977);
or U10941 (N_10941,N_6611,N_9291);
and U10942 (N_10942,N_8980,N_9227);
or U10943 (N_10943,N_6535,N_7820);
and U10944 (N_10944,N_6438,N_7110);
nor U10945 (N_10945,N_8450,N_8338);
nand U10946 (N_10946,N_6801,N_7312);
nand U10947 (N_10947,N_8069,N_7272);
nor U10948 (N_10948,N_7759,N_6251);
or U10949 (N_10949,N_9160,N_7878);
and U10950 (N_10950,N_7345,N_6913);
nand U10951 (N_10951,N_7108,N_6452);
or U10952 (N_10952,N_8622,N_7599);
nor U10953 (N_10953,N_9357,N_8863);
nand U10954 (N_10954,N_9356,N_8475);
xor U10955 (N_10955,N_7576,N_8384);
xor U10956 (N_10956,N_6874,N_9145);
or U10957 (N_10957,N_9183,N_8194);
nor U10958 (N_10958,N_8178,N_6884);
nand U10959 (N_10959,N_7382,N_6565);
nor U10960 (N_10960,N_8919,N_8501);
xor U10961 (N_10961,N_6436,N_8549);
and U10962 (N_10962,N_6659,N_7158);
nand U10963 (N_10963,N_6300,N_6773);
or U10964 (N_10964,N_6855,N_8313);
xor U10965 (N_10965,N_6717,N_8432);
nand U10966 (N_10966,N_7805,N_6799);
xor U10967 (N_10967,N_6604,N_7478);
xnor U10968 (N_10968,N_8509,N_8566);
and U10969 (N_10969,N_7289,N_6798);
xor U10970 (N_10970,N_7051,N_9206);
and U10971 (N_10971,N_8602,N_7437);
xnor U10972 (N_10972,N_7311,N_6380);
nor U10973 (N_10973,N_9039,N_9280);
and U10974 (N_10974,N_6768,N_6614);
nand U10975 (N_10975,N_7777,N_7262);
or U10976 (N_10976,N_7874,N_8882);
nor U10977 (N_10977,N_9137,N_8091);
nand U10978 (N_10978,N_7431,N_7502);
xnor U10979 (N_10979,N_7846,N_7590);
and U10980 (N_10980,N_8340,N_6699);
xor U10981 (N_10981,N_7755,N_7821);
nand U10982 (N_10982,N_6993,N_7736);
nor U10983 (N_10983,N_7619,N_6398);
nor U10984 (N_10984,N_7736,N_7188);
xor U10985 (N_10985,N_8377,N_6776);
xor U10986 (N_10986,N_7371,N_7514);
nor U10987 (N_10987,N_8604,N_6880);
xnor U10988 (N_10988,N_8633,N_8063);
xor U10989 (N_10989,N_6295,N_7613);
and U10990 (N_10990,N_8173,N_6373);
or U10991 (N_10991,N_8127,N_7396);
xor U10992 (N_10992,N_6526,N_7406);
nand U10993 (N_10993,N_7061,N_8801);
nor U10994 (N_10994,N_6878,N_8285);
and U10995 (N_10995,N_7462,N_6760);
or U10996 (N_10996,N_6829,N_7388);
xnor U10997 (N_10997,N_8617,N_7397);
or U10998 (N_10998,N_7154,N_8258);
and U10999 (N_10999,N_6714,N_9150);
and U11000 (N_11000,N_6620,N_9277);
xor U11001 (N_11001,N_7049,N_8856);
and U11002 (N_11002,N_7741,N_7652);
nand U11003 (N_11003,N_7112,N_8735);
and U11004 (N_11004,N_6286,N_7648);
nand U11005 (N_11005,N_7709,N_7542);
nand U11006 (N_11006,N_7487,N_6548);
nand U11007 (N_11007,N_8762,N_7961);
nand U11008 (N_11008,N_8625,N_6379);
or U11009 (N_11009,N_8135,N_9116);
xnor U11010 (N_11010,N_8315,N_6735);
nand U11011 (N_11011,N_9287,N_6560);
xnor U11012 (N_11012,N_8633,N_7292);
and U11013 (N_11013,N_7503,N_6322);
nor U11014 (N_11014,N_7682,N_7294);
or U11015 (N_11015,N_7725,N_6307);
nand U11016 (N_11016,N_9316,N_7564);
nand U11017 (N_11017,N_6862,N_7871);
or U11018 (N_11018,N_8146,N_6782);
and U11019 (N_11019,N_7002,N_7833);
and U11020 (N_11020,N_6913,N_8900);
and U11021 (N_11021,N_8670,N_7439);
nor U11022 (N_11022,N_8272,N_9272);
nor U11023 (N_11023,N_7725,N_8745);
xnor U11024 (N_11024,N_6284,N_6860);
or U11025 (N_11025,N_8871,N_8572);
or U11026 (N_11026,N_7492,N_7919);
nor U11027 (N_11027,N_7489,N_7100);
and U11028 (N_11028,N_8599,N_7744);
nor U11029 (N_11029,N_6417,N_9271);
xnor U11030 (N_11030,N_8932,N_7579);
nor U11031 (N_11031,N_8208,N_6251);
nor U11032 (N_11032,N_6608,N_8281);
and U11033 (N_11033,N_8438,N_7840);
nor U11034 (N_11034,N_6727,N_6260);
nand U11035 (N_11035,N_6401,N_6957);
nor U11036 (N_11036,N_8800,N_6909);
or U11037 (N_11037,N_7966,N_6863);
or U11038 (N_11038,N_6894,N_6912);
or U11039 (N_11039,N_9088,N_6597);
xnor U11040 (N_11040,N_8713,N_7290);
xnor U11041 (N_11041,N_8853,N_9248);
and U11042 (N_11042,N_7123,N_6367);
or U11043 (N_11043,N_7281,N_8473);
nor U11044 (N_11044,N_7380,N_9273);
and U11045 (N_11045,N_7418,N_6287);
and U11046 (N_11046,N_7216,N_7456);
xor U11047 (N_11047,N_8913,N_7989);
nor U11048 (N_11048,N_8242,N_8241);
nor U11049 (N_11049,N_7388,N_9228);
and U11050 (N_11050,N_9152,N_9295);
nor U11051 (N_11051,N_6382,N_8798);
xnor U11052 (N_11052,N_6783,N_8447);
and U11053 (N_11053,N_6649,N_7814);
and U11054 (N_11054,N_8439,N_8810);
or U11055 (N_11055,N_7297,N_7121);
nor U11056 (N_11056,N_7429,N_6523);
nor U11057 (N_11057,N_8780,N_6887);
nor U11058 (N_11058,N_9338,N_8955);
or U11059 (N_11059,N_6751,N_8909);
or U11060 (N_11060,N_8020,N_6455);
and U11061 (N_11061,N_8894,N_8321);
or U11062 (N_11062,N_9096,N_6709);
nand U11063 (N_11063,N_7055,N_8197);
nand U11064 (N_11064,N_6368,N_6276);
or U11065 (N_11065,N_8484,N_6752);
xnor U11066 (N_11066,N_7048,N_7588);
nand U11067 (N_11067,N_7659,N_6256);
or U11068 (N_11068,N_7348,N_8734);
nand U11069 (N_11069,N_6965,N_9324);
nand U11070 (N_11070,N_7935,N_8379);
xor U11071 (N_11071,N_6913,N_7181);
nor U11072 (N_11072,N_9367,N_7567);
or U11073 (N_11073,N_8437,N_8898);
xor U11074 (N_11074,N_6896,N_7406);
nand U11075 (N_11075,N_8153,N_6982);
and U11076 (N_11076,N_6417,N_7137);
xnor U11077 (N_11077,N_8982,N_9185);
or U11078 (N_11078,N_8129,N_7553);
nand U11079 (N_11079,N_7189,N_7273);
and U11080 (N_11080,N_6948,N_6566);
nand U11081 (N_11081,N_7866,N_9044);
xnor U11082 (N_11082,N_8979,N_9113);
or U11083 (N_11083,N_8943,N_9024);
xnor U11084 (N_11084,N_7695,N_7018);
nor U11085 (N_11085,N_7364,N_8817);
or U11086 (N_11086,N_8875,N_7756);
or U11087 (N_11087,N_7601,N_7588);
nand U11088 (N_11088,N_7979,N_7324);
nand U11089 (N_11089,N_8021,N_6342);
nor U11090 (N_11090,N_7259,N_9178);
and U11091 (N_11091,N_8130,N_8232);
nand U11092 (N_11092,N_6595,N_7923);
nand U11093 (N_11093,N_9248,N_6998);
nor U11094 (N_11094,N_6327,N_6838);
and U11095 (N_11095,N_7910,N_6347);
nand U11096 (N_11096,N_9146,N_8173);
xor U11097 (N_11097,N_8197,N_7758);
xor U11098 (N_11098,N_7800,N_7767);
or U11099 (N_11099,N_9185,N_7746);
nand U11100 (N_11100,N_6354,N_8692);
nand U11101 (N_11101,N_6464,N_6459);
nor U11102 (N_11102,N_7581,N_6915);
and U11103 (N_11103,N_9340,N_8919);
nor U11104 (N_11104,N_6392,N_8889);
and U11105 (N_11105,N_8229,N_9268);
xor U11106 (N_11106,N_6629,N_7519);
nor U11107 (N_11107,N_9168,N_7533);
nand U11108 (N_11108,N_8998,N_6905);
nand U11109 (N_11109,N_8441,N_7478);
nand U11110 (N_11110,N_7094,N_8173);
xnor U11111 (N_11111,N_6621,N_9026);
and U11112 (N_11112,N_7788,N_6890);
nand U11113 (N_11113,N_6275,N_8746);
or U11114 (N_11114,N_7880,N_6526);
nor U11115 (N_11115,N_9100,N_7180);
or U11116 (N_11116,N_7239,N_9288);
nor U11117 (N_11117,N_6727,N_7718);
xnor U11118 (N_11118,N_9024,N_6362);
and U11119 (N_11119,N_8788,N_7889);
nor U11120 (N_11120,N_6894,N_8635);
nor U11121 (N_11121,N_6402,N_8010);
nand U11122 (N_11122,N_7555,N_6865);
nor U11123 (N_11123,N_6303,N_6674);
nand U11124 (N_11124,N_8906,N_7320);
nor U11125 (N_11125,N_8662,N_7401);
nor U11126 (N_11126,N_8675,N_9169);
or U11127 (N_11127,N_6471,N_7111);
xnor U11128 (N_11128,N_8392,N_6550);
nand U11129 (N_11129,N_9043,N_8768);
and U11130 (N_11130,N_8664,N_7475);
nor U11131 (N_11131,N_7771,N_8944);
nor U11132 (N_11132,N_8554,N_6355);
nor U11133 (N_11133,N_7449,N_6630);
xnor U11134 (N_11134,N_7288,N_7332);
or U11135 (N_11135,N_9091,N_7590);
or U11136 (N_11136,N_7557,N_7488);
nor U11137 (N_11137,N_8699,N_7877);
nor U11138 (N_11138,N_8356,N_7135);
or U11139 (N_11139,N_8386,N_6995);
and U11140 (N_11140,N_7396,N_7400);
or U11141 (N_11141,N_7593,N_9262);
and U11142 (N_11142,N_6953,N_7461);
xor U11143 (N_11143,N_6996,N_6818);
and U11144 (N_11144,N_7866,N_9048);
xor U11145 (N_11145,N_7123,N_7260);
nand U11146 (N_11146,N_6957,N_7076);
nand U11147 (N_11147,N_8480,N_8963);
nand U11148 (N_11148,N_6527,N_7249);
nor U11149 (N_11149,N_8387,N_9200);
and U11150 (N_11150,N_8937,N_6291);
nand U11151 (N_11151,N_6639,N_7368);
or U11152 (N_11152,N_6488,N_7468);
or U11153 (N_11153,N_7126,N_8433);
and U11154 (N_11154,N_7234,N_7443);
nand U11155 (N_11155,N_9268,N_6578);
nand U11156 (N_11156,N_7147,N_7284);
nor U11157 (N_11157,N_7855,N_7182);
and U11158 (N_11158,N_8132,N_7797);
nand U11159 (N_11159,N_8067,N_7473);
nand U11160 (N_11160,N_8710,N_6380);
and U11161 (N_11161,N_7761,N_7735);
xor U11162 (N_11162,N_7845,N_7524);
nand U11163 (N_11163,N_7935,N_7255);
or U11164 (N_11164,N_6861,N_8097);
and U11165 (N_11165,N_8565,N_8779);
nand U11166 (N_11166,N_8514,N_8416);
or U11167 (N_11167,N_9333,N_7934);
nand U11168 (N_11168,N_9172,N_6561);
nand U11169 (N_11169,N_6728,N_8716);
or U11170 (N_11170,N_6898,N_7178);
nor U11171 (N_11171,N_7029,N_6805);
nand U11172 (N_11172,N_8038,N_8367);
and U11173 (N_11173,N_8277,N_7679);
xor U11174 (N_11174,N_9210,N_6347);
and U11175 (N_11175,N_8363,N_8058);
and U11176 (N_11176,N_9191,N_7801);
nor U11177 (N_11177,N_7290,N_7054);
nor U11178 (N_11178,N_8088,N_6675);
and U11179 (N_11179,N_6996,N_6565);
or U11180 (N_11180,N_7381,N_7341);
nand U11181 (N_11181,N_8387,N_6397);
or U11182 (N_11182,N_8121,N_8829);
or U11183 (N_11183,N_7926,N_7210);
xor U11184 (N_11184,N_6500,N_6286);
nor U11185 (N_11185,N_9010,N_6981);
nor U11186 (N_11186,N_7757,N_8117);
xnor U11187 (N_11187,N_9335,N_8072);
nand U11188 (N_11188,N_9069,N_6740);
or U11189 (N_11189,N_6767,N_6701);
xor U11190 (N_11190,N_6577,N_7023);
nor U11191 (N_11191,N_7808,N_6488);
nor U11192 (N_11192,N_7043,N_6642);
or U11193 (N_11193,N_8362,N_7411);
nand U11194 (N_11194,N_7096,N_7536);
nor U11195 (N_11195,N_7360,N_7975);
xor U11196 (N_11196,N_8872,N_7022);
xor U11197 (N_11197,N_6467,N_7738);
nand U11198 (N_11198,N_7580,N_8691);
nand U11199 (N_11199,N_8358,N_8052);
and U11200 (N_11200,N_7427,N_6380);
nand U11201 (N_11201,N_6811,N_7894);
nand U11202 (N_11202,N_8097,N_8168);
or U11203 (N_11203,N_9153,N_8876);
nor U11204 (N_11204,N_8412,N_7880);
and U11205 (N_11205,N_6898,N_7228);
or U11206 (N_11206,N_7525,N_7710);
or U11207 (N_11207,N_7579,N_8743);
and U11208 (N_11208,N_6510,N_6309);
nand U11209 (N_11209,N_6638,N_7090);
xnor U11210 (N_11210,N_6447,N_7636);
nor U11211 (N_11211,N_6798,N_6347);
and U11212 (N_11212,N_9104,N_7716);
nand U11213 (N_11213,N_8711,N_7272);
xnor U11214 (N_11214,N_7974,N_8787);
or U11215 (N_11215,N_9184,N_9039);
and U11216 (N_11216,N_7490,N_8042);
xnor U11217 (N_11217,N_7878,N_7775);
xor U11218 (N_11218,N_8030,N_7464);
nor U11219 (N_11219,N_6664,N_7772);
xor U11220 (N_11220,N_7495,N_8413);
nand U11221 (N_11221,N_7262,N_6740);
nand U11222 (N_11222,N_8636,N_7109);
or U11223 (N_11223,N_7267,N_6311);
nand U11224 (N_11224,N_8083,N_7802);
or U11225 (N_11225,N_9060,N_6502);
nand U11226 (N_11226,N_7210,N_6614);
and U11227 (N_11227,N_6597,N_8547);
and U11228 (N_11228,N_6771,N_7826);
or U11229 (N_11229,N_7206,N_7796);
nand U11230 (N_11230,N_7690,N_7357);
nand U11231 (N_11231,N_6545,N_7132);
nor U11232 (N_11232,N_7632,N_6509);
nand U11233 (N_11233,N_7150,N_8405);
and U11234 (N_11234,N_8413,N_7105);
and U11235 (N_11235,N_9292,N_8737);
nor U11236 (N_11236,N_9160,N_7933);
xnor U11237 (N_11237,N_6572,N_6396);
xnor U11238 (N_11238,N_8270,N_7897);
or U11239 (N_11239,N_9179,N_7531);
and U11240 (N_11240,N_9228,N_7898);
xor U11241 (N_11241,N_8748,N_7841);
and U11242 (N_11242,N_7797,N_6990);
or U11243 (N_11243,N_7691,N_6868);
nor U11244 (N_11244,N_7818,N_7861);
nand U11245 (N_11245,N_7834,N_7220);
xnor U11246 (N_11246,N_8649,N_6949);
and U11247 (N_11247,N_6672,N_7089);
or U11248 (N_11248,N_8120,N_6668);
and U11249 (N_11249,N_8556,N_7228);
xnor U11250 (N_11250,N_8545,N_8034);
and U11251 (N_11251,N_8690,N_7150);
or U11252 (N_11252,N_6347,N_8527);
nor U11253 (N_11253,N_7162,N_8895);
nand U11254 (N_11254,N_6885,N_8149);
xnor U11255 (N_11255,N_9015,N_9005);
xor U11256 (N_11256,N_6891,N_9252);
or U11257 (N_11257,N_7825,N_6271);
xnor U11258 (N_11258,N_6308,N_6275);
and U11259 (N_11259,N_8084,N_9035);
nand U11260 (N_11260,N_8376,N_8254);
nor U11261 (N_11261,N_7847,N_8665);
nand U11262 (N_11262,N_8166,N_8832);
xor U11263 (N_11263,N_8243,N_7683);
nand U11264 (N_11264,N_8542,N_7819);
nor U11265 (N_11265,N_7121,N_7853);
nor U11266 (N_11266,N_9246,N_8974);
xor U11267 (N_11267,N_9019,N_7231);
nand U11268 (N_11268,N_8274,N_9199);
xor U11269 (N_11269,N_7297,N_8344);
or U11270 (N_11270,N_6480,N_6511);
xor U11271 (N_11271,N_9272,N_6326);
xnor U11272 (N_11272,N_7272,N_8898);
xnor U11273 (N_11273,N_7145,N_7634);
and U11274 (N_11274,N_7097,N_7089);
xor U11275 (N_11275,N_8463,N_7271);
or U11276 (N_11276,N_7291,N_7711);
and U11277 (N_11277,N_8152,N_7196);
or U11278 (N_11278,N_6922,N_6740);
nor U11279 (N_11279,N_6486,N_7107);
and U11280 (N_11280,N_6518,N_9252);
and U11281 (N_11281,N_8605,N_8260);
and U11282 (N_11282,N_9225,N_9319);
xor U11283 (N_11283,N_7186,N_7649);
xnor U11284 (N_11284,N_7129,N_7255);
and U11285 (N_11285,N_7683,N_7194);
or U11286 (N_11286,N_7189,N_7179);
and U11287 (N_11287,N_6761,N_7637);
nor U11288 (N_11288,N_7578,N_8726);
xor U11289 (N_11289,N_6535,N_6992);
nand U11290 (N_11290,N_6351,N_6804);
xnor U11291 (N_11291,N_8658,N_8265);
xor U11292 (N_11292,N_6289,N_8340);
and U11293 (N_11293,N_7960,N_9034);
nor U11294 (N_11294,N_7137,N_9237);
nand U11295 (N_11295,N_8351,N_8706);
and U11296 (N_11296,N_9290,N_6798);
xor U11297 (N_11297,N_6471,N_7049);
and U11298 (N_11298,N_8546,N_7302);
or U11299 (N_11299,N_8745,N_8584);
nor U11300 (N_11300,N_7083,N_6618);
xnor U11301 (N_11301,N_7786,N_7712);
or U11302 (N_11302,N_6757,N_9244);
or U11303 (N_11303,N_7324,N_7507);
or U11304 (N_11304,N_6575,N_8780);
or U11305 (N_11305,N_8758,N_9327);
and U11306 (N_11306,N_7741,N_7277);
or U11307 (N_11307,N_6551,N_8784);
and U11308 (N_11308,N_8532,N_7249);
and U11309 (N_11309,N_7928,N_7762);
nand U11310 (N_11310,N_7171,N_8411);
or U11311 (N_11311,N_8319,N_8452);
and U11312 (N_11312,N_6524,N_7985);
or U11313 (N_11313,N_8259,N_6357);
or U11314 (N_11314,N_9354,N_8975);
and U11315 (N_11315,N_7052,N_6704);
and U11316 (N_11316,N_9261,N_8555);
nand U11317 (N_11317,N_7862,N_7390);
or U11318 (N_11318,N_8160,N_8167);
and U11319 (N_11319,N_8636,N_8797);
xnor U11320 (N_11320,N_6331,N_7862);
xnor U11321 (N_11321,N_6730,N_7926);
nor U11322 (N_11322,N_9327,N_6832);
and U11323 (N_11323,N_7265,N_8796);
xor U11324 (N_11324,N_7143,N_8035);
or U11325 (N_11325,N_8565,N_8569);
and U11326 (N_11326,N_8192,N_8535);
nor U11327 (N_11327,N_6287,N_8315);
or U11328 (N_11328,N_8295,N_8677);
nand U11329 (N_11329,N_8338,N_7923);
nand U11330 (N_11330,N_9144,N_6778);
nor U11331 (N_11331,N_9312,N_6320);
xnor U11332 (N_11332,N_7880,N_9028);
and U11333 (N_11333,N_8231,N_7799);
nand U11334 (N_11334,N_7846,N_8666);
nand U11335 (N_11335,N_7304,N_7357);
nor U11336 (N_11336,N_9102,N_7310);
nand U11337 (N_11337,N_7277,N_9150);
nand U11338 (N_11338,N_7445,N_8097);
xor U11339 (N_11339,N_9037,N_6580);
xor U11340 (N_11340,N_6754,N_6251);
or U11341 (N_11341,N_9056,N_7444);
nor U11342 (N_11342,N_7430,N_8269);
xnor U11343 (N_11343,N_9300,N_8649);
xnor U11344 (N_11344,N_7361,N_7498);
nor U11345 (N_11345,N_8726,N_8788);
xnor U11346 (N_11346,N_8971,N_6579);
and U11347 (N_11347,N_6421,N_9085);
and U11348 (N_11348,N_8243,N_9288);
and U11349 (N_11349,N_9128,N_7012);
nand U11350 (N_11350,N_8495,N_7162);
xor U11351 (N_11351,N_6823,N_7721);
xnor U11352 (N_11352,N_7168,N_6897);
and U11353 (N_11353,N_7058,N_7423);
nor U11354 (N_11354,N_6430,N_7559);
xor U11355 (N_11355,N_6784,N_6843);
nor U11356 (N_11356,N_7215,N_8430);
nand U11357 (N_11357,N_7266,N_7930);
nand U11358 (N_11358,N_8648,N_8805);
or U11359 (N_11359,N_7189,N_6526);
or U11360 (N_11360,N_7912,N_7561);
xnor U11361 (N_11361,N_7774,N_7848);
nor U11362 (N_11362,N_6498,N_7086);
xnor U11363 (N_11363,N_7230,N_7188);
and U11364 (N_11364,N_9363,N_7356);
nand U11365 (N_11365,N_9134,N_7625);
nand U11366 (N_11366,N_8126,N_8196);
and U11367 (N_11367,N_8561,N_7530);
nor U11368 (N_11368,N_9278,N_7989);
nand U11369 (N_11369,N_6658,N_7925);
xnor U11370 (N_11370,N_9249,N_7039);
nor U11371 (N_11371,N_7227,N_6444);
nand U11372 (N_11372,N_9145,N_9027);
nand U11373 (N_11373,N_8368,N_6924);
and U11374 (N_11374,N_7039,N_7074);
or U11375 (N_11375,N_8733,N_7730);
or U11376 (N_11376,N_8798,N_7900);
xnor U11377 (N_11377,N_6949,N_6675);
or U11378 (N_11378,N_6983,N_6433);
nor U11379 (N_11379,N_6687,N_9281);
and U11380 (N_11380,N_8766,N_8045);
or U11381 (N_11381,N_8346,N_9180);
and U11382 (N_11382,N_6483,N_9066);
xor U11383 (N_11383,N_7086,N_7972);
nand U11384 (N_11384,N_8066,N_7167);
and U11385 (N_11385,N_7172,N_8991);
nor U11386 (N_11386,N_9324,N_6924);
xnor U11387 (N_11387,N_6897,N_7111);
nand U11388 (N_11388,N_6702,N_6625);
and U11389 (N_11389,N_8027,N_7428);
or U11390 (N_11390,N_8919,N_8750);
nor U11391 (N_11391,N_6267,N_7738);
or U11392 (N_11392,N_7429,N_6809);
xor U11393 (N_11393,N_7745,N_6495);
and U11394 (N_11394,N_7675,N_7742);
or U11395 (N_11395,N_7392,N_6307);
and U11396 (N_11396,N_8860,N_6403);
nand U11397 (N_11397,N_7380,N_7868);
and U11398 (N_11398,N_6573,N_7255);
xnor U11399 (N_11399,N_8387,N_9014);
nand U11400 (N_11400,N_8026,N_7979);
and U11401 (N_11401,N_7202,N_6728);
and U11402 (N_11402,N_8927,N_8627);
xor U11403 (N_11403,N_8923,N_9001);
xnor U11404 (N_11404,N_6813,N_9290);
nand U11405 (N_11405,N_8701,N_9036);
nor U11406 (N_11406,N_7650,N_6450);
and U11407 (N_11407,N_8902,N_6781);
or U11408 (N_11408,N_8835,N_8924);
xnor U11409 (N_11409,N_8021,N_6679);
xnor U11410 (N_11410,N_7184,N_6584);
or U11411 (N_11411,N_8110,N_8158);
nor U11412 (N_11412,N_8798,N_6886);
or U11413 (N_11413,N_7823,N_7472);
nor U11414 (N_11414,N_8741,N_6391);
nand U11415 (N_11415,N_9132,N_7391);
and U11416 (N_11416,N_7702,N_6923);
xor U11417 (N_11417,N_8742,N_8165);
nand U11418 (N_11418,N_9171,N_6781);
or U11419 (N_11419,N_7449,N_7474);
nand U11420 (N_11420,N_9192,N_8266);
or U11421 (N_11421,N_7032,N_8235);
nor U11422 (N_11422,N_6614,N_6382);
nor U11423 (N_11423,N_9055,N_7712);
nor U11424 (N_11424,N_8724,N_6820);
xnor U11425 (N_11425,N_8496,N_6767);
xor U11426 (N_11426,N_8582,N_6584);
and U11427 (N_11427,N_7259,N_8498);
nand U11428 (N_11428,N_6699,N_8125);
nand U11429 (N_11429,N_7895,N_8558);
xor U11430 (N_11430,N_7800,N_8588);
and U11431 (N_11431,N_8224,N_9070);
and U11432 (N_11432,N_7717,N_9105);
xnor U11433 (N_11433,N_8199,N_7329);
and U11434 (N_11434,N_8182,N_6251);
and U11435 (N_11435,N_8481,N_6574);
or U11436 (N_11436,N_8092,N_8569);
and U11437 (N_11437,N_6572,N_8740);
nand U11438 (N_11438,N_6991,N_6738);
and U11439 (N_11439,N_6813,N_6280);
xor U11440 (N_11440,N_6929,N_7686);
nor U11441 (N_11441,N_7902,N_7138);
nor U11442 (N_11442,N_8733,N_9155);
and U11443 (N_11443,N_7232,N_7878);
or U11444 (N_11444,N_7805,N_7594);
xor U11445 (N_11445,N_6331,N_7804);
nor U11446 (N_11446,N_8376,N_8157);
nor U11447 (N_11447,N_9353,N_8062);
xor U11448 (N_11448,N_8002,N_9141);
xnor U11449 (N_11449,N_7542,N_9342);
or U11450 (N_11450,N_7128,N_6634);
and U11451 (N_11451,N_7098,N_6655);
nand U11452 (N_11452,N_7597,N_7744);
xnor U11453 (N_11453,N_8841,N_7995);
xnor U11454 (N_11454,N_7435,N_8511);
nor U11455 (N_11455,N_8744,N_6744);
nand U11456 (N_11456,N_8063,N_7512);
nand U11457 (N_11457,N_8789,N_8329);
xnor U11458 (N_11458,N_9185,N_7198);
xnor U11459 (N_11459,N_7263,N_6722);
and U11460 (N_11460,N_8282,N_8390);
xnor U11461 (N_11461,N_6390,N_7675);
nand U11462 (N_11462,N_6843,N_9012);
or U11463 (N_11463,N_9173,N_8999);
nor U11464 (N_11464,N_7853,N_8400);
xor U11465 (N_11465,N_7267,N_7049);
or U11466 (N_11466,N_7150,N_7400);
xor U11467 (N_11467,N_7294,N_6606);
or U11468 (N_11468,N_7394,N_7682);
nand U11469 (N_11469,N_9204,N_9196);
xnor U11470 (N_11470,N_9373,N_8315);
xor U11471 (N_11471,N_8978,N_7835);
nand U11472 (N_11472,N_6690,N_9292);
or U11473 (N_11473,N_7342,N_7065);
or U11474 (N_11474,N_8108,N_6739);
xor U11475 (N_11475,N_7978,N_7730);
or U11476 (N_11476,N_6561,N_6324);
xor U11477 (N_11477,N_8281,N_8630);
nor U11478 (N_11478,N_9110,N_7566);
or U11479 (N_11479,N_8953,N_7186);
or U11480 (N_11480,N_9285,N_8265);
and U11481 (N_11481,N_7231,N_9241);
xnor U11482 (N_11482,N_9295,N_7520);
and U11483 (N_11483,N_6640,N_8200);
nand U11484 (N_11484,N_9147,N_8387);
xor U11485 (N_11485,N_8303,N_7817);
or U11486 (N_11486,N_6706,N_7759);
nand U11487 (N_11487,N_8020,N_6802);
and U11488 (N_11488,N_8573,N_6902);
or U11489 (N_11489,N_7067,N_8989);
nand U11490 (N_11490,N_7220,N_9131);
and U11491 (N_11491,N_9274,N_9314);
and U11492 (N_11492,N_6312,N_6920);
and U11493 (N_11493,N_7169,N_8215);
nor U11494 (N_11494,N_8477,N_8264);
or U11495 (N_11495,N_8915,N_8496);
and U11496 (N_11496,N_7942,N_7955);
or U11497 (N_11497,N_6421,N_8006);
or U11498 (N_11498,N_6561,N_6982);
nor U11499 (N_11499,N_8977,N_7919);
xnor U11500 (N_11500,N_7595,N_6634);
xnor U11501 (N_11501,N_7573,N_7468);
nand U11502 (N_11502,N_6657,N_8694);
xnor U11503 (N_11503,N_8912,N_8173);
nand U11504 (N_11504,N_6315,N_8025);
and U11505 (N_11505,N_6712,N_7750);
xnor U11506 (N_11506,N_8483,N_7904);
and U11507 (N_11507,N_8559,N_7356);
xnor U11508 (N_11508,N_7851,N_7596);
nor U11509 (N_11509,N_8206,N_8023);
or U11510 (N_11510,N_9181,N_7449);
or U11511 (N_11511,N_8086,N_8758);
or U11512 (N_11512,N_6822,N_7259);
or U11513 (N_11513,N_8104,N_9195);
and U11514 (N_11514,N_6315,N_7492);
and U11515 (N_11515,N_7912,N_7145);
and U11516 (N_11516,N_9048,N_7415);
xnor U11517 (N_11517,N_7392,N_6323);
or U11518 (N_11518,N_7482,N_7598);
nor U11519 (N_11519,N_6263,N_6524);
nand U11520 (N_11520,N_8809,N_7202);
and U11521 (N_11521,N_6838,N_9308);
and U11522 (N_11522,N_8286,N_8527);
or U11523 (N_11523,N_8654,N_6540);
and U11524 (N_11524,N_8992,N_6933);
or U11525 (N_11525,N_7460,N_8653);
or U11526 (N_11526,N_7469,N_6973);
nand U11527 (N_11527,N_9001,N_7727);
nor U11528 (N_11528,N_6906,N_6633);
and U11529 (N_11529,N_8211,N_8771);
nor U11530 (N_11530,N_7639,N_6719);
and U11531 (N_11531,N_7218,N_8886);
or U11532 (N_11532,N_6630,N_8505);
xnor U11533 (N_11533,N_6833,N_9013);
xnor U11534 (N_11534,N_8795,N_6954);
and U11535 (N_11535,N_7224,N_6895);
nand U11536 (N_11536,N_7925,N_8068);
xor U11537 (N_11537,N_8896,N_7194);
nor U11538 (N_11538,N_8773,N_6711);
and U11539 (N_11539,N_7326,N_6516);
nand U11540 (N_11540,N_7202,N_8948);
or U11541 (N_11541,N_7155,N_8218);
or U11542 (N_11542,N_8889,N_6559);
or U11543 (N_11543,N_8837,N_8050);
nand U11544 (N_11544,N_8661,N_8848);
or U11545 (N_11545,N_8380,N_6515);
nand U11546 (N_11546,N_7151,N_9349);
and U11547 (N_11547,N_6358,N_6450);
or U11548 (N_11548,N_7067,N_9128);
nor U11549 (N_11549,N_8392,N_8408);
xor U11550 (N_11550,N_8459,N_6412);
nand U11551 (N_11551,N_7182,N_8667);
or U11552 (N_11552,N_7342,N_7565);
and U11553 (N_11553,N_7746,N_8605);
or U11554 (N_11554,N_8292,N_6716);
xor U11555 (N_11555,N_7634,N_8695);
xnor U11556 (N_11556,N_6982,N_6411);
nor U11557 (N_11557,N_6572,N_6375);
or U11558 (N_11558,N_6585,N_7567);
xnor U11559 (N_11559,N_8495,N_7388);
nand U11560 (N_11560,N_8081,N_7466);
nand U11561 (N_11561,N_6415,N_8514);
xnor U11562 (N_11562,N_7475,N_8920);
nor U11563 (N_11563,N_7646,N_6741);
or U11564 (N_11564,N_7043,N_6682);
nand U11565 (N_11565,N_7522,N_7926);
nand U11566 (N_11566,N_6827,N_7278);
and U11567 (N_11567,N_7818,N_7875);
nand U11568 (N_11568,N_7150,N_8894);
and U11569 (N_11569,N_8797,N_9190);
or U11570 (N_11570,N_8498,N_7972);
nor U11571 (N_11571,N_8069,N_8507);
nor U11572 (N_11572,N_8054,N_7263);
and U11573 (N_11573,N_8385,N_8451);
xor U11574 (N_11574,N_8599,N_6900);
or U11575 (N_11575,N_7602,N_8205);
nand U11576 (N_11576,N_7611,N_7207);
nand U11577 (N_11577,N_6823,N_8473);
nor U11578 (N_11578,N_7021,N_7494);
nor U11579 (N_11579,N_8976,N_6409);
and U11580 (N_11580,N_6310,N_6588);
and U11581 (N_11581,N_6985,N_8354);
or U11582 (N_11582,N_7155,N_8425);
or U11583 (N_11583,N_7155,N_8696);
and U11584 (N_11584,N_9136,N_7662);
nor U11585 (N_11585,N_6328,N_7790);
nor U11586 (N_11586,N_9073,N_8190);
nand U11587 (N_11587,N_8829,N_9326);
and U11588 (N_11588,N_7062,N_7041);
nor U11589 (N_11589,N_7812,N_8390);
or U11590 (N_11590,N_8246,N_6850);
or U11591 (N_11591,N_7832,N_6513);
nand U11592 (N_11592,N_8098,N_8914);
nand U11593 (N_11593,N_7551,N_7165);
nand U11594 (N_11594,N_7906,N_7780);
xnor U11595 (N_11595,N_8095,N_7935);
or U11596 (N_11596,N_6837,N_7503);
nand U11597 (N_11597,N_8472,N_7360);
nor U11598 (N_11598,N_8483,N_8610);
nor U11599 (N_11599,N_8994,N_8423);
and U11600 (N_11600,N_7554,N_8913);
nor U11601 (N_11601,N_6655,N_9093);
or U11602 (N_11602,N_7541,N_9270);
nor U11603 (N_11603,N_9055,N_9242);
nor U11604 (N_11604,N_7171,N_8624);
and U11605 (N_11605,N_9148,N_8542);
nor U11606 (N_11606,N_8542,N_7449);
nor U11607 (N_11607,N_7724,N_7208);
or U11608 (N_11608,N_9303,N_6948);
or U11609 (N_11609,N_7470,N_6387);
and U11610 (N_11610,N_8402,N_6616);
or U11611 (N_11611,N_6967,N_7909);
nor U11612 (N_11612,N_7399,N_9186);
and U11613 (N_11613,N_8205,N_9070);
nor U11614 (N_11614,N_6587,N_7937);
nor U11615 (N_11615,N_8645,N_7690);
or U11616 (N_11616,N_6746,N_8263);
and U11617 (N_11617,N_8761,N_7612);
xor U11618 (N_11618,N_6590,N_7304);
and U11619 (N_11619,N_8810,N_8828);
nor U11620 (N_11620,N_8405,N_8069);
or U11621 (N_11621,N_8475,N_8933);
and U11622 (N_11622,N_6695,N_6880);
nand U11623 (N_11623,N_8669,N_7412);
nor U11624 (N_11624,N_8946,N_8061);
nand U11625 (N_11625,N_6743,N_9180);
or U11626 (N_11626,N_6790,N_9285);
xor U11627 (N_11627,N_6422,N_7374);
xor U11628 (N_11628,N_9152,N_6658);
nand U11629 (N_11629,N_7113,N_7719);
nor U11630 (N_11630,N_8349,N_8645);
nor U11631 (N_11631,N_6467,N_8669);
and U11632 (N_11632,N_8346,N_6363);
xnor U11633 (N_11633,N_8023,N_9305);
xnor U11634 (N_11634,N_8680,N_8030);
nor U11635 (N_11635,N_9329,N_7189);
nor U11636 (N_11636,N_7827,N_9151);
xnor U11637 (N_11637,N_6936,N_6644);
nand U11638 (N_11638,N_8117,N_9191);
xor U11639 (N_11639,N_7765,N_8995);
or U11640 (N_11640,N_8774,N_7796);
nand U11641 (N_11641,N_8791,N_7982);
and U11642 (N_11642,N_6698,N_8968);
xnor U11643 (N_11643,N_9066,N_7547);
nor U11644 (N_11644,N_6545,N_8527);
nand U11645 (N_11645,N_8892,N_6464);
nor U11646 (N_11646,N_8003,N_7385);
and U11647 (N_11647,N_6579,N_7681);
xor U11648 (N_11648,N_7521,N_7539);
or U11649 (N_11649,N_8241,N_6650);
nand U11650 (N_11650,N_7497,N_7872);
or U11651 (N_11651,N_8230,N_8092);
xor U11652 (N_11652,N_6622,N_8382);
and U11653 (N_11653,N_7928,N_8684);
and U11654 (N_11654,N_8061,N_7101);
nor U11655 (N_11655,N_9051,N_7228);
xnor U11656 (N_11656,N_6775,N_7117);
nand U11657 (N_11657,N_8608,N_7099);
nor U11658 (N_11658,N_6321,N_8460);
nand U11659 (N_11659,N_6932,N_8145);
nor U11660 (N_11660,N_7077,N_8145);
nor U11661 (N_11661,N_7120,N_9287);
and U11662 (N_11662,N_7098,N_6454);
or U11663 (N_11663,N_8172,N_7170);
nor U11664 (N_11664,N_6402,N_8890);
and U11665 (N_11665,N_9334,N_8551);
or U11666 (N_11666,N_8349,N_8890);
xor U11667 (N_11667,N_7788,N_6809);
nor U11668 (N_11668,N_8146,N_8228);
nand U11669 (N_11669,N_8393,N_8632);
or U11670 (N_11670,N_6921,N_8251);
or U11671 (N_11671,N_9202,N_7898);
xnor U11672 (N_11672,N_8933,N_7077);
xor U11673 (N_11673,N_6809,N_6717);
xnor U11674 (N_11674,N_9062,N_6852);
or U11675 (N_11675,N_8302,N_8750);
or U11676 (N_11676,N_8672,N_8628);
nor U11677 (N_11677,N_8887,N_8847);
nor U11678 (N_11678,N_8540,N_9108);
and U11679 (N_11679,N_6261,N_8975);
nor U11680 (N_11680,N_9136,N_8970);
xnor U11681 (N_11681,N_7415,N_8429);
and U11682 (N_11682,N_6809,N_8449);
and U11683 (N_11683,N_9050,N_6760);
xor U11684 (N_11684,N_7853,N_8799);
nand U11685 (N_11685,N_8530,N_8537);
xnor U11686 (N_11686,N_7179,N_8148);
nor U11687 (N_11687,N_6811,N_6876);
or U11688 (N_11688,N_8062,N_8420);
xnor U11689 (N_11689,N_8589,N_8424);
or U11690 (N_11690,N_7250,N_9373);
nand U11691 (N_11691,N_9355,N_8459);
nand U11692 (N_11692,N_7643,N_7053);
and U11693 (N_11693,N_6887,N_8852);
or U11694 (N_11694,N_7921,N_6927);
xnor U11695 (N_11695,N_7966,N_7804);
nand U11696 (N_11696,N_7377,N_8612);
xnor U11697 (N_11697,N_6533,N_6647);
and U11698 (N_11698,N_8501,N_8492);
or U11699 (N_11699,N_6786,N_7164);
xor U11700 (N_11700,N_8598,N_8031);
and U11701 (N_11701,N_7096,N_9245);
nand U11702 (N_11702,N_7461,N_7466);
or U11703 (N_11703,N_8525,N_7870);
xnor U11704 (N_11704,N_9039,N_6377);
nor U11705 (N_11705,N_6882,N_8084);
and U11706 (N_11706,N_6338,N_8793);
and U11707 (N_11707,N_9280,N_7735);
nand U11708 (N_11708,N_7650,N_7925);
nor U11709 (N_11709,N_9123,N_6638);
and U11710 (N_11710,N_7995,N_6945);
xor U11711 (N_11711,N_8059,N_7049);
and U11712 (N_11712,N_8497,N_7268);
or U11713 (N_11713,N_8678,N_8646);
xnor U11714 (N_11714,N_6889,N_8746);
nor U11715 (N_11715,N_9052,N_6670);
nor U11716 (N_11716,N_7636,N_6819);
nand U11717 (N_11717,N_7079,N_8562);
nand U11718 (N_11718,N_8146,N_6900);
nand U11719 (N_11719,N_6939,N_9271);
nor U11720 (N_11720,N_8796,N_7911);
or U11721 (N_11721,N_9156,N_7033);
and U11722 (N_11722,N_8030,N_6857);
nor U11723 (N_11723,N_9239,N_7132);
xnor U11724 (N_11724,N_7684,N_8874);
xnor U11725 (N_11725,N_6488,N_7677);
or U11726 (N_11726,N_8848,N_7880);
nand U11727 (N_11727,N_7863,N_7029);
and U11728 (N_11728,N_6456,N_9073);
nor U11729 (N_11729,N_9107,N_6600);
nor U11730 (N_11730,N_9098,N_9043);
nor U11731 (N_11731,N_8248,N_6766);
nand U11732 (N_11732,N_6987,N_8723);
and U11733 (N_11733,N_8052,N_8246);
or U11734 (N_11734,N_9001,N_8250);
and U11735 (N_11735,N_8601,N_7090);
nor U11736 (N_11736,N_7679,N_7491);
xor U11737 (N_11737,N_6390,N_6488);
nor U11738 (N_11738,N_6827,N_7806);
or U11739 (N_11739,N_7080,N_9241);
nand U11740 (N_11740,N_7803,N_6701);
nor U11741 (N_11741,N_8802,N_7111);
nor U11742 (N_11742,N_7380,N_9199);
xnor U11743 (N_11743,N_6401,N_7796);
nand U11744 (N_11744,N_7596,N_7593);
or U11745 (N_11745,N_8797,N_7770);
xor U11746 (N_11746,N_9143,N_7834);
and U11747 (N_11747,N_7306,N_8885);
nand U11748 (N_11748,N_8147,N_8780);
and U11749 (N_11749,N_6347,N_8485);
xor U11750 (N_11750,N_8388,N_6802);
and U11751 (N_11751,N_6817,N_8805);
nand U11752 (N_11752,N_7408,N_9083);
nor U11753 (N_11753,N_7883,N_6416);
and U11754 (N_11754,N_8181,N_7997);
xnor U11755 (N_11755,N_6828,N_6318);
nand U11756 (N_11756,N_9167,N_7837);
nand U11757 (N_11757,N_7515,N_7796);
xnor U11758 (N_11758,N_7311,N_8350);
nand U11759 (N_11759,N_8792,N_7653);
or U11760 (N_11760,N_6641,N_6879);
xnor U11761 (N_11761,N_8071,N_9155);
nor U11762 (N_11762,N_6875,N_6902);
or U11763 (N_11763,N_9098,N_7325);
and U11764 (N_11764,N_6798,N_6364);
and U11765 (N_11765,N_8403,N_9324);
or U11766 (N_11766,N_7806,N_8887);
and U11767 (N_11767,N_8842,N_7684);
nand U11768 (N_11768,N_8199,N_7338);
nor U11769 (N_11769,N_9129,N_8564);
xor U11770 (N_11770,N_6290,N_7846);
and U11771 (N_11771,N_9159,N_9062);
xnor U11772 (N_11772,N_7104,N_7944);
nor U11773 (N_11773,N_7658,N_7716);
nor U11774 (N_11774,N_8759,N_8377);
nor U11775 (N_11775,N_9152,N_6880);
nor U11776 (N_11776,N_9054,N_8687);
nand U11777 (N_11777,N_7714,N_6583);
xnor U11778 (N_11778,N_8862,N_7166);
nand U11779 (N_11779,N_7712,N_7500);
nand U11780 (N_11780,N_6712,N_9285);
xor U11781 (N_11781,N_8407,N_6657);
and U11782 (N_11782,N_9147,N_8955);
xor U11783 (N_11783,N_9258,N_7390);
and U11784 (N_11784,N_7018,N_7506);
nand U11785 (N_11785,N_6834,N_6302);
nor U11786 (N_11786,N_8816,N_7487);
and U11787 (N_11787,N_7633,N_6830);
nand U11788 (N_11788,N_6719,N_8122);
xnor U11789 (N_11789,N_7946,N_9311);
nor U11790 (N_11790,N_7307,N_8044);
nand U11791 (N_11791,N_6309,N_6492);
xor U11792 (N_11792,N_8433,N_7206);
xnor U11793 (N_11793,N_8365,N_7343);
xnor U11794 (N_11794,N_9342,N_6409);
or U11795 (N_11795,N_8746,N_6307);
and U11796 (N_11796,N_9161,N_8962);
nor U11797 (N_11797,N_8760,N_8746);
or U11798 (N_11798,N_9017,N_6406);
or U11799 (N_11799,N_7936,N_7403);
nand U11800 (N_11800,N_6327,N_7252);
xor U11801 (N_11801,N_8084,N_8208);
or U11802 (N_11802,N_7205,N_9293);
or U11803 (N_11803,N_7520,N_7360);
nand U11804 (N_11804,N_7930,N_6605);
xnor U11805 (N_11805,N_7950,N_7859);
nand U11806 (N_11806,N_9367,N_9052);
xor U11807 (N_11807,N_6527,N_7608);
and U11808 (N_11808,N_7783,N_6912);
or U11809 (N_11809,N_7314,N_8662);
and U11810 (N_11810,N_7742,N_6751);
xnor U11811 (N_11811,N_6622,N_8338);
or U11812 (N_11812,N_8240,N_6899);
nand U11813 (N_11813,N_8579,N_8077);
xor U11814 (N_11814,N_8281,N_7916);
xnor U11815 (N_11815,N_6751,N_6668);
xor U11816 (N_11816,N_6759,N_8476);
nand U11817 (N_11817,N_9020,N_8925);
nand U11818 (N_11818,N_8639,N_7960);
nor U11819 (N_11819,N_7628,N_6680);
and U11820 (N_11820,N_6706,N_9073);
xnor U11821 (N_11821,N_6321,N_6677);
or U11822 (N_11822,N_7787,N_9232);
nor U11823 (N_11823,N_8287,N_7627);
or U11824 (N_11824,N_9203,N_9239);
and U11825 (N_11825,N_7049,N_6744);
nand U11826 (N_11826,N_6817,N_6881);
nand U11827 (N_11827,N_8322,N_8088);
and U11828 (N_11828,N_7719,N_7196);
xnor U11829 (N_11829,N_9104,N_7446);
and U11830 (N_11830,N_8643,N_8263);
nand U11831 (N_11831,N_6609,N_7125);
nand U11832 (N_11832,N_9216,N_7693);
nand U11833 (N_11833,N_6664,N_9119);
xor U11834 (N_11834,N_8728,N_7729);
nand U11835 (N_11835,N_7033,N_6848);
or U11836 (N_11836,N_6366,N_6846);
xnor U11837 (N_11837,N_7593,N_7701);
or U11838 (N_11838,N_6609,N_6883);
xnor U11839 (N_11839,N_8540,N_9182);
nand U11840 (N_11840,N_9274,N_8454);
nor U11841 (N_11841,N_9071,N_6961);
and U11842 (N_11842,N_9301,N_8194);
and U11843 (N_11843,N_7002,N_7655);
xnor U11844 (N_11844,N_6863,N_7524);
nand U11845 (N_11845,N_8518,N_7012);
and U11846 (N_11846,N_6967,N_8491);
nor U11847 (N_11847,N_6916,N_8477);
and U11848 (N_11848,N_8147,N_8747);
nand U11849 (N_11849,N_6287,N_7406);
nor U11850 (N_11850,N_7257,N_8856);
nor U11851 (N_11851,N_7676,N_7030);
nor U11852 (N_11852,N_8460,N_6539);
nand U11853 (N_11853,N_7890,N_7058);
or U11854 (N_11854,N_8915,N_8824);
xnor U11855 (N_11855,N_7125,N_6450);
xnor U11856 (N_11856,N_7587,N_6362);
or U11857 (N_11857,N_6486,N_8147);
nor U11858 (N_11858,N_8536,N_8730);
or U11859 (N_11859,N_6953,N_7684);
or U11860 (N_11860,N_6901,N_8113);
and U11861 (N_11861,N_8212,N_7134);
nand U11862 (N_11862,N_9080,N_8241);
and U11863 (N_11863,N_8918,N_8217);
or U11864 (N_11864,N_9023,N_7121);
xor U11865 (N_11865,N_7987,N_6830);
xor U11866 (N_11866,N_6871,N_6594);
or U11867 (N_11867,N_6525,N_7441);
nand U11868 (N_11868,N_8119,N_6916);
nand U11869 (N_11869,N_7607,N_6698);
nand U11870 (N_11870,N_8392,N_7332);
and U11871 (N_11871,N_8670,N_8028);
or U11872 (N_11872,N_8370,N_8700);
and U11873 (N_11873,N_8906,N_6973);
or U11874 (N_11874,N_8246,N_6340);
nor U11875 (N_11875,N_8636,N_8606);
nor U11876 (N_11876,N_9330,N_8281);
nand U11877 (N_11877,N_6621,N_7315);
xor U11878 (N_11878,N_6642,N_9358);
or U11879 (N_11879,N_6434,N_6893);
nor U11880 (N_11880,N_6595,N_6969);
and U11881 (N_11881,N_7434,N_7884);
nand U11882 (N_11882,N_9229,N_7373);
nor U11883 (N_11883,N_8938,N_9013);
xnor U11884 (N_11884,N_7703,N_8097);
and U11885 (N_11885,N_9057,N_6390);
and U11886 (N_11886,N_6332,N_7142);
nand U11887 (N_11887,N_7250,N_7129);
nand U11888 (N_11888,N_7723,N_8536);
or U11889 (N_11889,N_9028,N_6690);
nand U11890 (N_11890,N_8372,N_7143);
nor U11891 (N_11891,N_9026,N_8230);
xnor U11892 (N_11892,N_8332,N_8777);
nand U11893 (N_11893,N_8824,N_7253);
or U11894 (N_11894,N_6412,N_8023);
and U11895 (N_11895,N_7314,N_8816);
nor U11896 (N_11896,N_6346,N_8251);
xor U11897 (N_11897,N_7489,N_7536);
and U11898 (N_11898,N_6570,N_7125);
xor U11899 (N_11899,N_7783,N_9225);
or U11900 (N_11900,N_9142,N_7656);
or U11901 (N_11901,N_8922,N_7232);
nand U11902 (N_11902,N_6475,N_6859);
xor U11903 (N_11903,N_8377,N_7437);
nor U11904 (N_11904,N_7012,N_9096);
and U11905 (N_11905,N_8893,N_6846);
and U11906 (N_11906,N_8201,N_8835);
nor U11907 (N_11907,N_6587,N_7210);
nand U11908 (N_11908,N_8752,N_6939);
and U11909 (N_11909,N_9203,N_8665);
and U11910 (N_11910,N_7785,N_8713);
and U11911 (N_11911,N_7963,N_9363);
nor U11912 (N_11912,N_8220,N_8687);
xnor U11913 (N_11913,N_8032,N_7586);
and U11914 (N_11914,N_6798,N_7762);
nor U11915 (N_11915,N_8661,N_6342);
xor U11916 (N_11916,N_7129,N_6773);
nand U11917 (N_11917,N_6377,N_7308);
and U11918 (N_11918,N_8883,N_8670);
and U11919 (N_11919,N_7075,N_8433);
and U11920 (N_11920,N_6736,N_8355);
nor U11921 (N_11921,N_6251,N_6877);
xnor U11922 (N_11922,N_6377,N_7526);
nor U11923 (N_11923,N_7539,N_7340);
or U11924 (N_11924,N_8060,N_8317);
nor U11925 (N_11925,N_8556,N_7489);
and U11926 (N_11926,N_8939,N_7207);
or U11927 (N_11927,N_7540,N_8595);
nand U11928 (N_11928,N_8798,N_9367);
and U11929 (N_11929,N_7891,N_6276);
xor U11930 (N_11930,N_8867,N_8740);
nor U11931 (N_11931,N_6795,N_8157);
or U11932 (N_11932,N_6965,N_8618);
and U11933 (N_11933,N_9278,N_9256);
or U11934 (N_11934,N_7283,N_8022);
nand U11935 (N_11935,N_6860,N_9007);
and U11936 (N_11936,N_8271,N_6825);
nor U11937 (N_11937,N_9073,N_8886);
or U11938 (N_11938,N_7975,N_7991);
and U11939 (N_11939,N_7114,N_8199);
nor U11940 (N_11940,N_8080,N_7984);
or U11941 (N_11941,N_7688,N_6694);
xnor U11942 (N_11942,N_8432,N_6822);
xor U11943 (N_11943,N_7866,N_7164);
nand U11944 (N_11944,N_9126,N_8749);
and U11945 (N_11945,N_6596,N_8583);
nand U11946 (N_11946,N_6735,N_8108);
or U11947 (N_11947,N_8422,N_7646);
and U11948 (N_11948,N_8188,N_6597);
and U11949 (N_11949,N_8441,N_6816);
nor U11950 (N_11950,N_7229,N_6694);
nand U11951 (N_11951,N_9122,N_6664);
nand U11952 (N_11952,N_7982,N_8326);
xor U11953 (N_11953,N_8483,N_6938);
xor U11954 (N_11954,N_6396,N_6517);
nand U11955 (N_11955,N_7391,N_7471);
nand U11956 (N_11956,N_7894,N_7133);
or U11957 (N_11957,N_7228,N_7215);
nor U11958 (N_11958,N_8611,N_7008);
xnor U11959 (N_11959,N_6612,N_6665);
or U11960 (N_11960,N_7536,N_6970);
nor U11961 (N_11961,N_6451,N_7423);
or U11962 (N_11962,N_8004,N_7483);
and U11963 (N_11963,N_7584,N_8785);
nor U11964 (N_11964,N_6797,N_7556);
nand U11965 (N_11965,N_9252,N_9067);
nand U11966 (N_11966,N_6516,N_8176);
and U11967 (N_11967,N_8118,N_7728);
nor U11968 (N_11968,N_8956,N_8382);
and U11969 (N_11969,N_8974,N_6368);
xnor U11970 (N_11970,N_7241,N_8333);
or U11971 (N_11971,N_7104,N_6768);
and U11972 (N_11972,N_8845,N_6679);
and U11973 (N_11973,N_7749,N_7540);
or U11974 (N_11974,N_6334,N_9011);
xor U11975 (N_11975,N_9306,N_8915);
nor U11976 (N_11976,N_8229,N_9157);
nand U11977 (N_11977,N_7946,N_6423);
and U11978 (N_11978,N_7990,N_8023);
xor U11979 (N_11979,N_7701,N_7683);
xor U11980 (N_11980,N_8227,N_9157);
nand U11981 (N_11981,N_8700,N_7646);
nor U11982 (N_11982,N_7199,N_8521);
and U11983 (N_11983,N_8598,N_7207);
or U11984 (N_11984,N_9044,N_8805);
nand U11985 (N_11985,N_6292,N_7676);
or U11986 (N_11986,N_7352,N_6876);
nand U11987 (N_11987,N_8913,N_8977);
or U11988 (N_11988,N_8603,N_7041);
or U11989 (N_11989,N_8678,N_8312);
xor U11990 (N_11990,N_7234,N_8932);
nand U11991 (N_11991,N_8718,N_6588);
nand U11992 (N_11992,N_8047,N_9266);
nor U11993 (N_11993,N_8737,N_9263);
xnor U11994 (N_11994,N_7638,N_8764);
nor U11995 (N_11995,N_8483,N_9002);
xnor U11996 (N_11996,N_7118,N_7695);
nand U11997 (N_11997,N_8869,N_7243);
or U11998 (N_11998,N_7665,N_8762);
or U11999 (N_11999,N_9085,N_7525);
or U12000 (N_12000,N_6272,N_7022);
nand U12001 (N_12001,N_7054,N_8056);
and U12002 (N_12002,N_7438,N_7999);
nand U12003 (N_12003,N_7536,N_9084);
xor U12004 (N_12004,N_7491,N_9119);
nor U12005 (N_12005,N_8505,N_7853);
and U12006 (N_12006,N_6556,N_7130);
and U12007 (N_12007,N_8147,N_7266);
nor U12008 (N_12008,N_6288,N_9159);
nand U12009 (N_12009,N_7796,N_8583);
nor U12010 (N_12010,N_7569,N_8866);
nor U12011 (N_12011,N_8756,N_7673);
nor U12012 (N_12012,N_9120,N_8575);
or U12013 (N_12013,N_8013,N_6971);
or U12014 (N_12014,N_8376,N_7884);
xor U12015 (N_12015,N_6887,N_8349);
and U12016 (N_12016,N_6426,N_7688);
and U12017 (N_12017,N_7065,N_9293);
or U12018 (N_12018,N_6607,N_6949);
and U12019 (N_12019,N_7336,N_9163);
nor U12020 (N_12020,N_8590,N_7029);
or U12021 (N_12021,N_6716,N_7851);
nand U12022 (N_12022,N_8888,N_8825);
nand U12023 (N_12023,N_6638,N_7699);
and U12024 (N_12024,N_6400,N_9222);
and U12025 (N_12025,N_9084,N_7535);
xnor U12026 (N_12026,N_8778,N_8837);
xor U12027 (N_12027,N_7653,N_6764);
xnor U12028 (N_12028,N_7137,N_8401);
xnor U12029 (N_12029,N_7745,N_8373);
and U12030 (N_12030,N_7351,N_7687);
xnor U12031 (N_12031,N_7342,N_6729);
or U12032 (N_12032,N_7938,N_7146);
nor U12033 (N_12033,N_8910,N_7095);
xnor U12034 (N_12034,N_9169,N_8532);
nor U12035 (N_12035,N_6520,N_8986);
xor U12036 (N_12036,N_9337,N_9115);
nand U12037 (N_12037,N_8000,N_7208);
xor U12038 (N_12038,N_7005,N_7452);
xor U12039 (N_12039,N_7261,N_8843);
nand U12040 (N_12040,N_6568,N_6769);
and U12041 (N_12041,N_7931,N_8592);
and U12042 (N_12042,N_8462,N_8393);
nor U12043 (N_12043,N_8452,N_6462);
nor U12044 (N_12044,N_6390,N_7085);
or U12045 (N_12045,N_6383,N_7800);
xor U12046 (N_12046,N_9151,N_6690);
nand U12047 (N_12047,N_7958,N_7748);
and U12048 (N_12048,N_6798,N_8019);
and U12049 (N_12049,N_6653,N_6268);
or U12050 (N_12050,N_8431,N_8297);
and U12051 (N_12051,N_8897,N_6326);
and U12052 (N_12052,N_6585,N_8380);
and U12053 (N_12053,N_8674,N_8707);
xor U12054 (N_12054,N_8657,N_8458);
nor U12055 (N_12055,N_7952,N_9206);
nand U12056 (N_12056,N_8841,N_9262);
or U12057 (N_12057,N_6677,N_8680);
or U12058 (N_12058,N_6772,N_8524);
and U12059 (N_12059,N_6358,N_7000);
nor U12060 (N_12060,N_8294,N_8420);
and U12061 (N_12061,N_7416,N_7028);
or U12062 (N_12062,N_6773,N_8349);
xor U12063 (N_12063,N_6991,N_7995);
nand U12064 (N_12064,N_6257,N_7741);
xor U12065 (N_12065,N_8299,N_7789);
and U12066 (N_12066,N_9222,N_9181);
nor U12067 (N_12067,N_7770,N_8890);
and U12068 (N_12068,N_6533,N_6965);
and U12069 (N_12069,N_8270,N_7346);
xnor U12070 (N_12070,N_8767,N_6415);
and U12071 (N_12071,N_8708,N_6521);
nand U12072 (N_12072,N_9202,N_9022);
nor U12073 (N_12073,N_7522,N_8334);
nand U12074 (N_12074,N_7201,N_9209);
nor U12075 (N_12075,N_9224,N_7317);
or U12076 (N_12076,N_7986,N_8121);
xnor U12077 (N_12077,N_7238,N_8902);
nand U12078 (N_12078,N_7070,N_6977);
nor U12079 (N_12079,N_7338,N_8914);
nor U12080 (N_12080,N_6320,N_7374);
and U12081 (N_12081,N_9268,N_7626);
or U12082 (N_12082,N_7077,N_6538);
nand U12083 (N_12083,N_7128,N_8489);
nand U12084 (N_12084,N_6345,N_8556);
or U12085 (N_12085,N_7159,N_7141);
nor U12086 (N_12086,N_7384,N_7285);
nand U12087 (N_12087,N_8508,N_6482);
or U12088 (N_12088,N_6766,N_7184);
xor U12089 (N_12089,N_8247,N_8221);
xor U12090 (N_12090,N_7962,N_7326);
or U12091 (N_12091,N_6532,N_6265);
xnor U12092 (N_12092,N_8295,N_8135);
nor U12093 (N_12093,N_7395,N_7225);
nand U12094 (N_12094,N_8041,N_9299);
nor U12095 (N_12095,N_8692,N_7888);
and U12096 (N_12096,N_6985,N_8099);
nand U12097 (N_12097,N_9068,N_7142);
nand U12098 (N_12098,N_7663,N_6748);
nor U12099 (N_12099,N_6921,N_9010);
nor U12100 (N_12100,N_7784,N_7710);
nand U12101 (N_12101,N_8857,N_8479);
and U12102 (N_12102,N_8177,N_9054);
and U12103 (N_12103,N_8918,N_8928);
or U12104 (N_12104,N_7512,N_6496);
and U12105 (N_12105,N_7507,N_7854);
xor U12106 (N_12106,N_8748,N_8825);
and U12107 (N_12107,N_6298,N_7811);
nand U12108 (N_12108,N_7393,N_8829);
nand U12109 (N_12109,N_6656,N_7688);
xnor U12110 (N_12110,N_8337,N_8165);
nand U12111 (N_12111,N_9350,N_6257);
nand U12112 (N_12112,N_7559,N_8688);
xor U12113 (N_12113,N_7182,N_7464);
and U12114 (N_12114,N_8182,N_7157);
nor U12115 (N_12115,N_9364,N_8056);
or U12116 (N_12116,N_6404,N_8188);
nor U12117 (N_12117,N_7230,N_6707);
nor U12118 (N_12118,N_8345,N_6454);
nor U12119 (N_12119,N_6887,N_9262);
or U12120 (N_12120,N_8185,N_8233);
xor U12121 (N_12121,N_8183,N_7471);
nand U12122 (N_12122,N_8560,N_8844);
and U12123 (N_12123,N_8967,N_7518);
or U12124 (N_12124,N_6550,N_7503);
nand U12125 (N_12125,N_7494,N_7381);
and U12126 (N_12126,N_6415,N_8540);
xor U12127 (N_12127,N_7436,N_7636);
nand U12128 (N_12128,N_8301,N_8518);
xnor U12129 (N_12129,N_6898,N_6823);
or U12130 (N_12130,N_7936,N_8418);
nand U12131 (N_12131,N_9336,N_7891);
nand U12132 (N_12132,N_7357,N_9373);
nand U12133 (N_12133,N_7032,N_7591);
or U12134 (N_12134,N_7701,N_6757);
or U12135 (N_12135,N_8273,N_9245);
or U12136 (N_12136,N_7862,N_9009);
nor U12137 (N_12137,N_7673,N_7296);
nand U12138 (N_12138,N_7714,N_8371);
or U12139 (N_12139,N_9082,N_7242);
or U12140 (N_12140,N_6910,N_8140);
nand U12141 (N_12141,N_8842,N_8821);
xnor U12142 (N_12142,N_7145,N_9031);
nand U12143 (N_12143,N_7093,N_7128);
xnor U12144 (N_12144,N_7647,N_8240);
xnor U12145 (N_12145,N_7797,N_9045);
nor U12146 (N_12146,N_8336,N_8844);
or U12147 (N_12147,N_6263,N_7481);
nor U12148 (N_12148,N_7682,N_8457);
and U12149 (N_12149,N_9079,N_7163);
nand U12150 (N_12150,N_9287,N_7676);
nor U12151 (N_12151,N_7829,N_7114);
and U12152 (N_12152,N_8168,N_7012);
nand U12153 (N_12153,N_8398,N_8123);
or U12154 (N_12154,N_8605,N_7734);
or U12155 (N_12155,N_9281,N_6774);
nor U12156 (N_12156,N_6527,N_9007);
and U12157 (N_12157,N_9294,N_7397);
xnor U12158 (N_12158,N_9211,N_7727);
and U12159 (N_12159,N_6814,N_6381);
xnor U12160 (N_12160,N_8460,N_9020);
or U12161 (N_12161,N_6918,N_8569);
nand U12162 (N_12162,N_6849,N_7293);
or U12163 (N_12163,N_7160,N_8089);
nor U12164 (N_12164,N_7747,N_6900);
nand U12165 (N_12165,N_9313,N_9182);
and U12166 (N_12166,N_6955,N_8826);
or U12167 (N_12167,N_8876,N_8899);
or U12168 (N_12168,N_7381,N_7640);
or U12169 (N_12169,N_7035,N_8495);
nand U12170 (N_12170,N_9262,N_8046);
or U12171 (N_12171,N_6720,N_8296);
nor U12172 (N_12172,N_6559,N_7479);
xnor U12173 (N_12173,N_8850,N_7316);
or U12174 (N_12174,N_7687,N_7207);
and U12175 (N_12175,N_6908,N_7632);
xor U12176 (N_12176,N_9015,N_9107);
or U12177 (N_12177,N_7902,N_8660);
nand U12178 (N_12178,N_7823,N_9107);
nor U12179 (N_12179,N_8091,N_9112);
nand U12180 (N_12180,N_7888,N_8751);
nor U12181 (N_12181,N_7248,N_8219);
and U12182 (N_12182,N_6681,N_8765);
xnor U12183 (N_12183,N_7569,N_9057);
nor U12184 (N_12184,N_7299,N_7423);
nand U12185 (N_12185,N_7661,N_6988);
nor U12186 (N_12186,N_8503,N_7195);
nor U12187 (N_12187,N_8801,N_8954);
nor U12188 (N_12188,N_7685,N_8013);
nand U12189 (N_12189,N_7322,N_7103);
nor U12190 (N_12190,N_7115,N_8057);
nor U12191 (N_12191,N_8170,N_8405);
nor U12192 (N_12192,N_8775,N_8576);
xnor U12193 (N_12193,N_7136,N_8722);
or U12194 (N_12194,N_7774,N_7863);
nand U12195 (N_12195,N_6452,N_9040);
or U12196 (N_12196,N_9324,N_7343);
and U12197 (N_12197,N_8339,N_7122);
and U12198 (N_12198,N_8789,N_6847);
and U12199 (N_12199,N_8618,N_6789);
nor U12200 (N_12200,N_6493,N_6330);
nand U12201 (N_12201,N_7234,N_6559);
nor U12202 (N_12202,N_8815,N_8393);
xnor U12203 (N_12203,N_6766,N_7580);
nor U12204 (N_12204,N_7012,N_6978);
or U12205 (N_12205,N_8787,N_7090);
and U12206 (N_12206,N_6935,N_8948);
xor U12207 (N_12207,N_8081,N_7528);
nand U12208 (N_12208,N_8858,N_7017);
nand U12209 (N_12209,N_7400,N_8669);
nor U12210 (N_12210,N_8682,N_6820);
or U12211 (N_12211,N_7737,N_7288);
nor U12212 (N_12212,N_7509,N_9327);
and U12213 (N_12213,N_9227,N_6820);
and U12214 (N_12214,N_6754,N_7201);
or U12215 (N_12215,N_8153,N_6657);
and U12216 (N_12216,N_7958,N_8823);
nor U12217 (N_12217,N_6611,N_8147);
or U12218 (N_12218,N_7414,N_6486);
and U12219 (N_12219,N_8222,N_9069);
nand U12220 (N_12220,N_6969,N_7374);
or U12221 (N_12221,N_9339,N_8540);
nor U12222 (N_12222,N_6601,N_8924);
or U12223 (N_12223,N_7623,N_6517);
nor U12224 (N_12224,N_7488,N_8458);
or U12225 (N_12225,N_8592,N_6510);
and U12226 (N_12226,N_7983,N_7046);
and U12227 (N_12227,N_7759,N_8515);
and U12228 (N_12228,N_7725,N_9128);
nor U12229 (N_12229,N_8526,N_8586);
xnor U12230 (N_12230,N_7743,N_6657);
nor U12231 (N_12231,N_7705,N_6581);
nand U12232 (N_12232,N_8575,N_7258);
or U12233 (N_12233,N_6695,N_8697);
nor U12234 (N_12234,N_8900,N_8785);
nand U12235 (N_12235,N_7277,N_6833);
or U12236 (N_12236,N_7200,N_7128);
and U12237 (N_12237,N_8554,N_6899);
and U12238 (N_12238,N_6714,N_6390);
or U12239 (N_12239,N_7945,N_9277);
xnor U12240 (N_12240,N_9186,N_8592);
nand U12241 (N_12241,N_8165,N_8566);
xnor U12242 (N_12242,N_7454,N_8932);
nor U12243 (N_12243,N_6356,N_7037);
nor U12244 (N_12244,N_7998,N_8249);
nor U12245 (N_12245,N_8377,N_7379);
xnor U12246 (N_12246,N_7930,N_9267);
nor U12247 (N_12247,N_8209,N_8466);
nand U12248 (N_12248,N_8966,N_8494);
xnor U12249 (N_12249,N_6448,N_8600);
or U12250 (N_12250,N_7987,N_7700);
nand U12251 (N_12251,N_7924,N_7825);
and U12252 (N_12252,N_7162,N_9016);
and U12253 (N_12253,N_7391,N_9218);
and U12254 (N_12254,N_8308,N_8317);
nor U12255 (N_12255,N_7892,N_8839);
and U12256 (N_12256,N_7607,N_7634);
nand U12257 (N_12257,N_9162,N_7509);
nor U12258 (N_12258,N_8368,N_7306);
nor U12259 (N_12259,N_9190,N_9229);
or U12260 (N_12260,N_8026,N_9042);
xor U12261 (N_12261,N_8619,N_7748);
nor U12262 (N_12262,N_9092,N_9113);
and U12263 (N_12263,N_9291,N_9023);
nor U12264 (N_12264,N_9193,N_6451);
xor U12265 (N_12265,N_8178,N_6889);
and U12266 (N_12266,N_8020,N_8022);
nor U12267 (N_12267,N_8766,N_7086);
and U12268 (N_12268,N_7526,N_6792);
and U12269 (N_12269,N_7745,N_7721);
or U12270 (N_12270,N_9365,N_8483);
xnor U12271 (N_12271,N_6905,N_8151);
xnor U12272 (N_12272,N_8331,N_8457);
and U12273 (N_12273,N_6565,N_9099);
nor U12274 (N_12274,N_7651,N_7303);
nor U12275 (N_12275,N_6430,N_7698);
and U12276 (N_12276,N_8156,N_9014);
and U12277 (N_12277,N_8595,N_6812);
and U12278 (N_12278,N_7838,N_6899);
xnor U12279 (N_12279,N_9155,N_9019);
nor U12280 (N_12280,N_7124,N_8979);
nand U12281 (N_12281,N_6642,N_6279);
and U12282 (N_12282,N_7743,N_8685);
and U12283 (N_12283,N_7669,N_8098);
xnor U12284 (N_12284,N_7138,N_6335);
and U12285 (N_12285,N_7450,N_8884);
nand U12286 (N_12286,N_7851,N_7527);
or U12287 (N_12287,N_8939,N_6808);
and U12288 (N_12288,N_6763,N_7681);
or U12289 (N_12289,N_7636,N_7150);
nand U12290 (N_12290,N_6404,N_6686);
nor U12291 (N_12291,N_8771,N_6913);
and U12292 (N_12292,N_8091,N_6419);
nand U12293 (N_12293,N_6586,N_8751);
nor U12294 (N_12294,N_8191,N_8951);
or U12295 (N_12295,N_6421,N_9144);
and U12296 (N_12296,N_6505,N_8823);
nor U12297 (N_12297,N_8808,N_8476);
or U12298 (N_12298,N_7844,N_9200);
nor U12299 (N_12299,N_6588,N_6697);
or U12300 (N_12300,N_7411,N_8798);
and U12301 (N_12301,N_6897,N_9246);
nand U12302 (N_12302,N_8860,N_6335);
or U12303 (N_12303,N_9262,N_6789);
nor U12304 (N_12304,N_6943,N_9246);
nor U12305 (N_12305,N_6365,N_7240);
nor U12306 (N_12306,N_7892,N_8347);
nor U12307 (N_12307,N_6712,N_8340);
or U12308 (N_12308,N_6305,N_6633);
nand U12309 (N_12309,N_8745,N_8288);
or U12310 (N_12310,N_9139,N_7494);
nor U12311 (N_12311,N_8581,N_7423);
nor U12312 (N_12312,N_8376,N_6814);
or U12313 (N_12313,N_8070,N_7078);
or U12314 (N_12314,N_6778,N_7863);
xor U12315 (N_12315,N_7249,N_7809);
nor U12316 (N_12316,N_6743,N_6882);
and U12317 (N_12317,N_7270,N_7039);
or U12318 (N_12318,N_7451,N_9289);
nand U12319 (N_12319,N_7128,N_6973);
or U12320 (N_12320,N_7796,N_7718);
or U12321 (N_12321,N_7812,N_7779);
nand U12322 (N_12322,N_7243,N_8225);
and U12323 (N_12323,N_9047,N_8430);
nand U12324 (N_12324,N_8518,N_7511);
nand U12325 (N_12325,N_7943,N_7602);
or U12326 (N_12326,N_6267,N_9042);
nand U12327 (N_12327,N_8890,N_7241);
or U12328 (N_12328,N_8216,N_9197);
and U12329 (N_12329,N_6890,N_8624);
xnor U12330 (N_12330,N_6796,N_7145);
or U12331 (N_12331,N_8529,N_6540);
xnor U12332 (N_12332,N_8832,N_8524);
or U12333 (N_12333,N_8337,N_7775);
and U12334 (N_12334,N_7648,N_7720);
and U12335 (N_12335,N_7844,N_6858);
or U12336 (N_12336,N_6605,N_7093);
or U12337 (N_12337,N_6832,N_9274);
xor U12338 (N_12338,N_7508,N_8622);
nor U12339 (N_12339,N_8870,N_6927);
xnor U12340 (N_12340,N_6263,N_9284);
xnor U12341 (N_12341,N_6997,N_7836);
or U12342 (N_12342,N_6956,N_7039);
xor U12343 (N_12343,N_8262,N_8748);
xnor U12344 (N_12344,N_8873,N_7948);
and U12345 (N_12345,N_6979,N_7786);
and U12346 (N_12346,N_8946,N_8539);
nand U12347 (N_12347,N_7266,N_6284);
nor U12348 (N_12348,N_8732,N_8453);
and U12349 (N_12349,N_7366,N_8032);
xnor U12350 (N_12350,N_6921,N_6538);
or U12351 (N_12351,N_8760,N_9044);
xnor U12352 (N_12352,N_8354,N_7601);
nor U12353 (N_12353,N_7292,N_8409);
nor U12354 (N_12354,N_6336,N_6787);
and U12355 (N_12355,N_7712,N_7072);
xor U12356 (N_12356,N_6799,N_9030);
and U12357 (N_12357,N_7792,N_6723);
nor U12358 (N_12358,N_7097,N_8977);
or U12359 (N_12359,N_7028,N_6574);
or U12360 (N_12360,N_7963,N_8492);
or U12361 (N_12361,N_6482,N_8697);
or U12362 (N_12362,N_6267,N_7017);
nor U12363 (N_12363,N_8812,N_8889);
and U12364 (N_12364,N_8159,N_7706);
xnor U12365 (N_12365,N_8979,N_9222);
xor U12366 (N_12366,N_8229,N_7608);
and U12367 (N_12367,N_7163,N_8372);
nor U12368 (N_12368,N_8107,N_6889);
and U12369 (N_12369,N_8277,N_7715);
nor U12370 (N_12370,N_7150,N_7118);
and U12371 (N_12371,N_8831,N_8845);
and U12372 (N_12372,N_6425,N_9123);
xor U12373 (N_12373,N_9039,N_7173);
and U12374 (N_12374,N_6377,N_7181);
nor U12375 (N_12375,N_7168,N_6294);
nor U12376 (N_12376,N_7016,N_6888);
or U12377 (N_12377,N_7751,N_8918);
and U12378 (N_12378,N_9250,N_7458);
or U12379 (N_12379,N_6849,N_7255);
or U12380 (N_12380,N_8634,N_7927);
or U12381 (N_12381,N_6870,N_9127);
nor U12382 (N_12382,N_6335,N_7023);
or U12383 (N_12383,N_8395,N_6689);
nand U12384 (N_12384,N_7546,N_8887);
xnor U12385 (N_12385,N_8128,N_6296);
nand U12386 (N_12386,N_8720,N_7375);
and U12387 (N_12387,N_7602,N_7321);
nand U12388 (N_12388,N_8625,N_9273);
and U12389 (N_12389,N_6265,N_8969);
and U12390 (N_12390,N_8193,N_7831);
or U12391 (N_12391,N_7299,N_7160);
or U12392 (N_12392,N_9177,N_6500);
or U12393 (N_12393,N_8355,N_7085);
or U12394 (N_12394,N_8882,N_9296);
and U12395 (N_12395,N_6690,N_6843);
or U12396 (N_12396,N_6692,N_6760);
or U12397 (N_12397,N_9310,N_8816);
or U12398 (N_12398,N_6412,N_7615);
and U12399 (N_12399,N_6360,N_7063);
or U12400 (N_12400,N_6869,N_7130);
xor U12401 (N_12401,N_7806,N_6405);
nor U12402 (N_12402,N_8856,N_6947);
nand U12403 (N_12403,N_7595,N_6880);
nor U12404 (N_12404,N_9316,N_7415);
or U12405 (N_12405,N_9286,N_7539);
or U12406 (N_12406,N_7964,N_6306);
nor U12407 (N_12407,N_6313,N_7515);
xor U12408 (N_12408,N_7727,N_7903);
xnor U12409 (N_12409,N_9325,N_7130);
nor U12410 (N_12410,N_7592,N_7879);
or U12411 (N_12411,N_7186,N_6544);
nand U12412 (N_12412,N_9090,N_6751);
xor U12413 (N_12413,N_6405,N_8133);
or U12414 (N_12414,N_6747,N_9070);
xor U12415 (N_12415,N_8136,N_8677);
xor U12416 (N_12416,N_6252,N_8742);
or U12417 (N_12417,N_9036,N_8693);
xnor U12418 (N_12418,N_9067,N_7340);
nand U12419 (N_12419,N_8891,N_7666);
nand U12420 (N_12420,N_8343,N_8550);
nor U12421 (N_12421,N_7374,N_8544);
nand U12422 (N_12422,N_7352,N_7563);
nor U12423 (N_12423,N_7618,N_8339);
nor U12424 (N_12424,N_9173,N_7666);
nor U12425 (N_12425,N_8531,N_8980);
or U12426 (N_12426,N_7203,N_7566);
and U12427 (N_12427,N_7862,N_9315);
or U12428 (N_12428,N_9356,N_7329);
and U12429 (N_12429,N_7823,N_7005);
or U12430 (N_12430,N_7237,N_7216);
nor U12431 (N_12431,N_7316,N_8045);
or U12432 (N_12432,N_6793,N_7144);
xnor U12433 (N_12433,N_9370,N_7188);
or U12434 (N_12434,N_6785,N_8553);
nand U12435 (N_12435,N_9367,N_7418);
or U12436 (N_12436,N_8418,N_6747);
nand U12437 (N_12437,N_9000,N_9149);
nand U12438 (N_12438,N_6586,N_9123);
and U12439 (N_12439,N_6935,N_9208);
or U12440 (N_12440,N_6951,N_8639);
and U12441 (N_12441,N_6579,N_6853);
xnor U12442 (N_12442,N_8879,N_8120);
xor U12443 (N_12443,N_6800,N_8412);
nand U12444 (N_12444,N_6424,N_8348);
xnor U12445 (N_12445,N_9340,N_8854);
and U12446 (N_12446,N_7414,N_8909);
or U12447 (N_12447,N_8043,N_8387);
or U12448 (N_12448,N_7326,N_9027);
or U12449 (N_12449,N_7650,N_7881);
or U12450 (N_12450,N_7442,N_6367);
nand U12451 (N_12451,N_7714,N_6301);
or U12452 (N_12452,N_7559,N_9240);
xnor U12453 (N_12453,N_6810,N_7745);
or U12454 (N_12454,N_6564,N_9215);
nor U12455 (N_12455,N_6855,N_7835);
and U12456 (N_12456,N_9142,N_6571);
nor U12457 (N_12457,N_7266,N_7093);
nand U12458 (N_12458,N_8059,N_6713);
or U12459 (N_12459,N_8950,N_8281);
and U12460 (N_12460,N_6957,N_9283);
nor U12461 (N_12461,N_7208,N_8308);
xor U12462 (N_12462,N_8537,N_6657);
xor U12463 (N_12463,N_8596,N_7575);
nand U12464 (N_12464,N_7807,N_7276);
nand U12465 (N_12465,N_7868,N_9081);
xnor U12466 (N_12466,N_7085,N_7245);
nor U12467 (N_12467,N_7309,N_8285);
nand U12468 (N_12468,N_8273,N_8806);
nand U12469 (N_12469,N_6373,N_6786);
or U12470 (N_12470,N_9165,N_6887);
or U12471 (N_12471,N_8342,N_6767);
nand U12472 (N_12472,N_7970,N_8729);
and U12473 (N_12473,N_7088,N_8110);
nor U12474 (N_12474,N_8696,N_6594);
or U12475 (N_12475,N_7504,N_6407);
nand U12476 (N_12476,N_8509,N_7326);
and U12477 (N_12477,N_9146,N_8790);
and U12478 (N_12478,N_7659,N_9352);
xor U12479 (N_12479,N_7997,N_6284);
and U12480 (N_12480,N_7426,N_7814);
nand U12481 (N_12481,N_7812,N_8589);
or U12482 (N_12482,N_7619,N_7922);
and U12483 (N_12483,N_6464,N_7319);
or U12484 (N_12484,N_8204,N_9119);
or U12485 (N_12485,N_6864,N_7252);
nor U12486 (N_12486,N_7596,N_6746);
or U12487 (N_12487,N_6824,N_8589);
xor U12488 (N_12488,N_7267,N_8840);
or U12489 (N_12489,N_8519,N_8197);
or U12490 (N_12490,N_6918,N_7566);
nor U12491 (N_12491,N_7164,N_9224);
and U12492 (N_12492,N_9065,N_9117);
nand U12493 (N_12493,N_9346,N_7358);
or U12494 (N_12494,N_8375,N_9278);
nand U12495 (N_12495,N_7530,N_8531);
or U12496 (N_12496,N_8948,N_8298);
and U12497 (N_12497,N_6952,N_7797);
and U12498 (N_12498,N_6705,N_8053);
xor U12499 (N_12499,N_9374,N_9147);
xor U12500 (N_12500,N_11557,N_9451);
xnor U12501 (N_12501,N_9658,N_10433);
nand U12502 (N_12502,N_10027,N_12425);
nand U12503 (N_12503,N_11328,N_12201);
nand U12504 (N_12504,N_10933,N_11718);
or U12505 (N_12505,N_11969,N_9797);
and U12506 (N_12506,N_11354,N_9722);
or U12507 (N_12507,N_10637,N_11780);
nand U12508 (N_12508,N_11228,N_11192);
or U12509 (N_12509,N_12051,N_11060);
nor U12510 (N_12510,N_9701,N_12370);
nand U12511 (N_12511,N_9907,N_10522);
xnor U12512 (N_12512,N_12423,N_11137);
and U12513 (N_12513,N_9683,N_11753);
nor U12514 (N_12514,N_10159,N_10183);
and U12515 (N_12515,N_10271,N_9444);
nor U12516 (N_12516,N_11380,N_12159);
xor U12517 (N_12517,N_10026,N_11761);
xnor U12518 (N_12518,N_12315,N_12093);
nor U12519 (N_12519,N_10405,N_10654);
nand U12520 (N_12520,N_11588,N_10961);
xor U12521 (N_12521,N_10584,N_10655);
or U12522 (N_12522,N_12234,N_10249);
xor U12523 (N_12523,N_11393,N_11420);
nor U12524 (N_12524,N_10479,N_11158);
or U12525 (N_12525,N_12071,N_9473);
and U12526 (N_12526,N_12145,N_11376);
nand U12527 (N_12527,N_10947,N_12161);
and U12528 (N_12528,N_11801,N_9665);
and U12529 (N_12529,N_12366,N_9791);
xnor U12530 (N_12530,N_11502,N_10029);
and U12531 (N_12531,N_12121,N_11472);
xor U12532 (N_12532,N_11889,N_9422);
or U12533 (N_12533,N_9922,N_11930);
nand U12534 (N_12534,N_9673,N_10207);
nor U12535 (N_12535,N_11675,N_10838);
or U12536 (N_12536,N_10975,N_11994);
or U12537 (N_12537,N_10043,N_10987);
nand U12538 (N_12538,N_10340,N_11288);
or U12539 (N_12539,N_11130,N_9738);
and U12540 (N_12540,N_10321,N_10318);
nand U12541 (N_12541,N_9868,N_12453);
or U12542 (N_12542,N_11534,N_10101);
nor U12543 (N_12543,N_10598,N_11359);
nand U12544 (N_12544,N_10325,N_10824);
and U12545 (N_12545,N_11307,N_9419);
nor U12546 (N_12546,N_9742,N_11519);
nand U12547 (N_12547,N_10127,N_10739);
or U12548 (N_12548,N_11574,N_11148);
xor U12549 (N_12549,N_11119,N_10526);
or U12550 (N_12550,N_11898,N_10005);
nor U12551 (N_12551,N_11135,N_9775);
or U12552 (N_12552,N_9932,N_12382);
and U12553 (N_12553,N_10107,N_10345);
nor U12554 (N_12554,N_10648,N_11261);
and U12555 (N_12555,N_12003,N_9729);
and U12556 (N_12556,N_11145,N_10721);
nand U12557 (N_12557,N_9719,N_11394);
nor U12558 (N_12558,N_10888,N_11657);
or U12559 (N_12559,N_11474,N_11373);
nand U12560 (N_12560,N_11643,N_11642);
nor U12561 (N_12561,N_12231,N_9455);
nor U12562 (N_12562,N_11701,N_10876);
or U12563 (N_12563,N_11841,N_9593);
and U12564 (N_12564,N_10121,N_10951);
xnor U12565 (N_12565,N_10532,N_11835);
nor U12566 (N_12566,N_12123,N_11853);
or U12567 (N_12567,N_12205,N_12210);
nor U12568 (N_12568,N_11647,N_10822);
nand U12569 (N_12569,N_9434,N_11721);
xnor U12570 (N_12570,N_11606,N_11322);
nand U12571 (N_12571,N_11506,N_9467);
or U12572 (N_12572,N_11034,N_10173);
nor U12573 (N_12573,N_12172,N_10455);
nor U12574 (N_12574,N_11608,N_12066);
xnor U12575 (N_12575,N_11447,N_11515);
nor U12576 (N_12576,N_10725,N_9957);
xor U12577 (N_12577,N_12289,N_9675);
or U12578 (N_12578,N_11844,N_9380);
and U12579 (N_12579,N_11090,N_10084);
xnor U12580 (N_12580,N_9395,N_11958);
or U12581 (N_12581,N_10176,N_10150);
nor U12582 (N_12582,N_9551,N_9713);
nand U12583 (N_12583,N_10421,N_10042);
xor U12584 (N_12584,N_9602,N_12449);
xor U12585 (N_12585,N_10643,N_11976);
or U12586 (N_12586,N_9777,N_11790);
xnor U12587 (N_12587,N_11103,N_10069);
nor U12588 (N_12588,N_9959,N_9962);
or U12589 (N_12589,N_11662,N_12222);
nand U12590 (N_12590,N_12469,N_12369);
nor U12591 (N_12591,N_12153,N_11399);
xnor U12592 (N_12592,N_12428,N_9747);
xor U12593 (N_12593,N_9681,N_11243);
xnor U12594 (N_12594,N_11395,N_11882);
or U12595 (N_12595,N_9820,N_11986);
xnor U12596 (N_12596,N_9877,N_11385);
and U12597 (N_12597,N_9656,N_11754);
and U12598 (N_12598,N_11859,N_12088);
or U12599 (N_12599,N_9408,N_9532);
xnor U12600 (N_12600,N_11398,N_11477);
nor U12601 (N_12601,N_11631,N_10125);
xor U12602 (N_12602,N_12048,N_10324);
nor U12603 (N_12603,N_10904,N_10449);
nand U12604 (N_12604,N_9426,N_10428);
xor U12605 (N_12605,N_9859,N_10308);
and U12606 (N_12606,N_12143,N_11171);
nor U12607 (N_12607,N_10067,N_11644);
xor U12608 (N_12608,N_10098,N_10148);
nand U12609 (N_12609,N_11838,N_11150);
nand U12610 (N_12610,N_10305,N_10141);
nand U12611 (N_12611,N_11939,N_11457);
or U12612 (N_12612,N_12266,N_9813);
and U12613 (N_12613,N_10264,N_12459);
and U12614 (N_12614,N_10041,N_9428);
nor U12615 (N_12615,N_9411,N_12399);
or U12616 (N_12616,N_12012,N_11475);
or U12617 (N_12617,N_11727,N_11639);
or U12618 (N_12618,N_9518,N_10400);
nor U12619 (N_12619,N_10561,N_11665);
and U12620 (N_12620,N_10260,N_10379);
nor U12621 (N_12621,N_9595,N_9889);
nor U12622 (N_12622,N_11524,N_12202);
nand U12623 (N_12623,N_9802,N_11873);
xor U12624 (N_12624,N_10863,N_12258);
nor U12625 (N_12625,N_12444,N_11944);
or U12626 (N_12626,N_9840,N_10074);
nor U12627 (N_12627,N_11156,N_12291);
nor U12628 (N_12628,N_11962,N_11972);
nand U12629 (N_12629,N_11071,N_12166);
nor U12630 (N_12630,N_11595,N_10454);
and U12631 (N_12631,N_12194,N_10918);
nand U12632 (N_12632,N_10233,N_11735);
or U12633 (N_12633,N_11527,N_9377);
nor U12634 (N_12634,N_12069,N_10446);
and U12635 (N_12635,N_11566,N_11061);
and U12636 (N_12636,N_10247,N_10699);
nand U12637 (N_12637,N_12294,N_12211);
and U12638 (N_12638,N_11811,N_9482);
nand U12639 (N_12639,N_11428,N_10900);
xor U12640 (N_12640,N_11031,N_12424);
or U12641 (N_12641,N_10778,N_9884);
and U12642 (N_12642,N_9787,N_9383);
and U12643 (N_12643,N_10160,N_9764);
nor U12644 (N_12644,N_10157,N_12059);
or U12645 (N_12645,N_10527,N_11212);
and U12646 (N_12646,N_10988,N_11531);
and U12647 (N_12647,N_10774,N_11717);
xnor U12648 (N_12648,N_10460,N_10520);
and U12649 (N_12649,N_9420,N_11567);
or U12650 (N_12650,N_10311,N_11802);
nor U12651 (N_12651,N_10779,N_11175);
xnor U12652 (N_12652,N_9967,N_11169);
nand U12653 (N_12653,N_9397,N_11798);
and U12654 (N_12654,N_10465,N_9730);
or U12655 (N_12655,N_9899,N_10187);
nor U12656 (N_12656,N_11523,N_11950);
nor U12657 (N_12657,N_10389,N_11051);
and U12658 (N_12658,N_10880,N_11846);
nand U12659 (N_12659,N_11746,N_11612);
or U12660 (N_12660,N_11493,N_10109);
or U12661 (N_12661,N_9429,N_11568);
and U12662 (N_12662,N_10943,N_11951);
xor U12663 (N_12663,N_11147,N_11864);
nor U12664 (N_12664,N_11234,N_9400);
nor U12665 (N_12665,N_9872,N_12152);
or U12666 (N_12666,N_11592,N_10765);
nor U12667 (N_12667,N_11286,N_9390);
nor U12668 (N_12668,N_10875,N_11940);
nor U12669 (N_12669,N_12317,N_12324);
nor U12670 (N_12670,N_11538,N_11869);
and U12671 (N_12671,N_9971,N_10147);
xnor U12672 (N_12672,N_9632,N_11489);
and U12673 (N_12673,N_9575,N_12075);
xor U12674 (N_12674,N_10035,N_10444);
xnor U12675 (N_12675,N_10129,N_12497);
xnor U12676 (N_12676,N_10222,N_10163);
xnor U12677 (N_12677,N_12192,N_10510);
nor U12678 (N_12678,N_9990,N_11292);
xnor U12679 (N_12679,N_10840,N_10979);
or U12680 (N_12680,N_9666,N_9534);
nor U12681 (N_12681,N_11163,N_9445);
nand U12682 (N_12682,N_12214,N_9671);
and U12683 (N_12683,N_10429,N_11315);
nand U12684 (N_12684,N_9672,N_9389);
nor U12685 (N_12685,N_10601,N_10694);
or U12686 (N_12686,N_11582,N_9960);
xnor U12687 (N_12687,N_10877,N_11351);
xor U12688 (N_12688,N_10945,N_11526);
nor U12689 (N_12689,N_12267,N_9762);
xor U12690 (N_12690,N_11299,N_11706);
nor U12691 (N_12691,N_11319,N_10870);
xor U12692 (N_12692,N_10331,N_10797);
nor U12693 (N_12693,N_10011,N_10813);
or U12694 (N_12694,N_9414,N_11876);
xnor U12695 (N_12695,N_10178,N_9677);
or U12696 (N_12696,N_11661,N_10133);
xnor U12697 (N_12697,N_11993,N_12353);
and U12698 (N_12698,N_11303,N_9424);
xor U12699 (N_12699,N_11056,N_9489);
or U12700 (N_12700,N_10594,N_11863);
or U12701 (N_12701,N_12436,N_11610);
xor U12702 (N_12702,N_10664,N_11217);
and U12703 (N_12703,N_9988,N_11903);
and U12704 (N_12704,N_9682,N_11808);
or U12705 (N_12705,N_10610,N_9376);
nand U12706 (N_12706,N_9963,N_12415);
nand U12707 (N_12707,N_11695,N_10899);
and U12708 (N_12708,N_12154,N_11855);
nand U12709 (N_12709,N_10806,N_10451);
nor U12710 (N_12710,N_10060,N_10291);
xnor U12711 (N_12711,N_9514,N_10737);
or U12712 (N_12712,N_10882,N_9494);
or U12713 (N_12713,N_10450,N_9793);
nand U12714 (N_12714,N_10910,N_9509);
and U12715 (N_12715,N_11082,N_10593);
xor U12716 (N_12716,N_9752,N_12349);
nand U12717 (N_12717,N_10589,N_11280);
and U12718 (N_12718,N_11205,N_11178);
or U12719 (N_12719,N_10905,N_10086);
xnor U12720 (N_12720,N_11374,N_12004);
and U12721 (N_12721,N_11905,N_11714);
xor U12722 (N_12722,N_11188,N_11249);
xor U12723 (N_12723,N_10030,N_10501);
nor U12724 (N_12724,N_11666,N_10403);
xor U12725 (N_12725,N_11312,N_10186);
xnor U12726 (N_12726,N_11929,N_11828);
nand U12727 (N_12727,N_9823,N_10008);
or U12728 (N_12728,N_11805,N_10518);
nor U12729 (N_12729,N_10269,N_10749);
or U12730 (N_12730,N_12014,N_10235);
nand U12731 (N_12731,N_11854,N_11659);
nor U12732 (N_12732,N_11029,N_10211);
nor U12733 (N_12733,N_9893,N_11155);
nand U12734 (N_12734,N_10033,N_11111);
nor U12735 (N_12735,N_10563,N_11674);
nor U12736 (N_12736,N_10327,N_11356);
or U12737 (N_12737,N_11776,N_11244);
and U12738 (N_12738,N_11933,N_10371);
nor U12739 (N_12739,N_10179,N_9880);
and U12740 (N_12740,N_10976,N_10969);
xnor U12741 (N_12741,N_9497,N_12218);
nand U12742 (N_12742,N_9921,N_12239);
or U12743 (N_12743,N_10798,N_12318);
or U12744 (N_12744,N_10748,N_10761);
or U12745 (N_12745,N_9405,N_9997);
nand U12746 (N_12746,N_11881,N_12476);
and U12747 (N_12747,N_10731,N_11470);
and U12748 (N_12748,N_11480,N_10754);
and U12749 (N_12749,N_12306,N_12160);
nand U12750 (N_12750,N_11340,N_10085);
nor U12751 (N_12751,N_10294,N_12302);
nand U12752 (N_12752,N_9594,N_10673);
nor U12753 (N_12753,N_11942,N_11529);
nand U12754 (N_12754,N_10075,N_10917);
nor U12755 (N_12755,N_10714,N_11732);
nand U12756 (N_12756,N_11166,N_12000);
or U12757 (N_12757,N_9382,N_12191);
and U12758 (N_12758,N_10695,N_12383);
nand U12759 (N_12759,N_11817,N_10712);
xor U12760 (N_12760,N_12460,N_11908);
and U12761 (N_12761,N_9588,N_10683);
or U12762 (N_12762,N_11093,N_10836);
nor U12763 (N_12763,N_10177,N_10016);
xnor U12764 (N_12764,N_12033,N_11274);
and U12765 (N_12765,N_11453,N_11609);
xor U12766 (N_12766,N_12485,N_10356);
nand U12767 (N_12767,N_10240,N_11125);
and U12768 (N_12768,N_9978,N_10262);
xnor U12769 (N_12769,N_9638,N_10878);
nor U12770 (N_12770,N_10804,N_10873);
and U12771 (N_12771,N_11065,N_11837);
xor U12772 (N_12772,N_9911,N_10815);
or U12773 (N_12773,N_10989,N_9816);
nor U12774 (N_12774,N_9973,N_9413);
nor U12775 (N_12775,N_10794,N_10441);
nand U12776 (N_12776,N_10558,N_11787);
nand U12777 (N_12777,N_12017,N_11232);
xor U12778 (N_12778,N_9982,N_12112);
nor U12779 (N_12779,N_11785,N_10828);
or U12780 (N_12780,N_11597,N_12401);
and U12781 (N_12781,N_9892,N_10885);
and U12782 (N_12782,N_11922,N_12396);
nor U12783 (N_12783,N_9447,N_10009);
or U12784 (N_12784,N_11865,N_12120);
and U12785 (N_12785,N_10632,N_9789);
xor U12786 (N_12786,N_9800,N_10184);
nand U12787 (N_12787,N_9460,N_12386);
nor U12788 (N_12788,N_10082,N_12471);
xor U12789 (N_12789,N_9449,N_9410);
and U12790 (N_12790,N_10088,N_9394);
xor U12791 (N_12791,N_9576,N_10785);
or U12792 (N_12792,N_11806,N_11707);
nand U12793 (N_12793,N_11036,N_11300);
xor U12794 (N_12794,N_12050,N_9586);
nand U12795 (N_12795,N_11210,N_10825);
xor U12796 (N_12796,N_11513,N_12101);
nand U12797 (N_12797,N_10508,N_10155);
xor U12798 (N_12798,N_10397,N_12344);
xor U12799 (N_12799,N_10528,N_9517);
or U12800 (N_12800,N_11043,N_11616);
and U12801 (N_12801,N_9941,N_12233);
or U12802 (N_12802,N_10134,N_10923);
or U12803 (N_12803,N_10046,N_9601);
xor U12804 (N_12804,N_11948,N_9568);
nand U12805 (N_12805,N_10162,N_11273);
or U12806 (N_12806,N_9996,N_10021);
or U12807 (N_12807,N_10152,N_9678);
nor U12808 (N_12808,N_11278,N_10808);
xor U12809 (N_12809,N_10199,N_11943);
nand U12810 (N_12810,N_11581,N_10320);
xor U12811 (N_12811,N_10409,N_10942);
nor U12812 (N_12812,N_10470,N_11416);
or U12813 (N_12813,N_10469,N_9505);
nor U12814 (N_12814,N_11058,N_11895);
xnor U12815 (N_12815,N_10434,N_9476);
nand U12816 (N_12816,N_10997,N_12010);
nand U12817 (N_12817,N_11450,N_9898);
nand U12818 (N_12818,N_10747,N_9403);
or U12819 (N_12819,N_9749,N_10866);
xor U12820 (N_12820,N_10368,N_10227);
or U12821 (N_12821,N_12013,N_9379);
nor U12822 (N_12822,N_12058,N_9852);
nor U12823 (N_12823,N_10919,N_10415);
nand U12824 (N_12824,N_11471,N_10827);
or U12825 (N_12825,N_10795,N_11751);
nor U12826 (N_12826,N_12379,N_11104);
and U12827 (N_12827,N_10841,N_11343);
xor U12828 (N_12828,N_12316,N_10472);
or U12829 (N_12829,N_11432,N_11214);
or U12830 (N_12830,N_12490,N_9731);
nor U12831 (N_12831,N_10427,N_10750);
or U12832 (N_12832,N_9544,N_10932);
or U12833 (N_12833,N_11935,N_11454);
xnor U12834 (N_12834,N_9808,N_10079);
or U12835 (N_12835,N_12107,N_10002);
nor U12836 (N_12836,N_11815,N_9825);
nand U12837 (N_12837,N_11803,N_10474);
and U12838 (N_12838,N_11964,N_12464);
nor U12839 (N_12839,N_10057,N_11240);
and U12840 (N_12840,N_10114,N_12078);
and U12841 (N_12841,N_10251,N_9788);
xor U12842 (N_12842,N_10566,N_12165);
nor U12843 (N_12843,N_9831,N_12252);
and U12844 (N_12844,N_10711,N_9409);
or U12845 (N_12845,N_9766,N_11073);
and U12846 (N_12846,N_10590,N_10944);
nand U12847 (N_12847,N_11615,N_11460);
and U12848 (N_12848,N_10414,N_9860);
nand U12849 (N_12849,N_9768,N_11341);
and U12850 (N_12850,N_12284,N_11005);
nor U12851 (N_12851,N_11885,N_9589);
nor U12852 (N_12852,N_11342,N_12297);
nand U12853 (N_12853,N_9432,N_12200);
nand U12854 (N_12854,N_12131,N_10662);
and U12855 (N_12855,N_10359,N_10225);
nand U12856 (N_12856,N_10642,N_11733);
nor U12857 (N_12857,N_12164,N_10545);
nor U12858 (N_12858,N_9975,N_9667);
and U12859 (N_12859,N_12024,N_11741);
or U12860 (N_12860,N_11847,N_11025);
nand U12861 (N_12861,N_11211,N_9779);
and U12862 (N_12862,N_10336,N_9483);
or U12863 (N_12863,N_11900,N_10334);
and U12864 (N_12864,N_10534,N_9533);
and U12865 (N_12865,N_12269,N_10145);
or U12866 (N_12866,N_12206,N_11369);
nand U12867 (N_12867,N_12385,N_12285);
nand U12868 (N_12868,N_9524,N_11064);
nand U12869 (N_12869,N_10916,N_10554);
and U12870 (N_12870,N_10758,N_10034);
xnor U12871 (N_12871,N_10887,N_9803);
and U12872 (N_12872,N_10071,N_9661);
xor U12873 (N_12873,N_11168,N_10971);
or U12874 (N_12874,N_12335,N_12094);
nor U12875 (N_12875,N_11542,N_11172);
xor U12876 (N_12876,N_11936,N_11443);
or U12877 (N_12877,N_11079,N_11251);
nand U12878 (N_12878,N_10775,N_11893);
xor U12879 (N_12879,N_12413,N_11194);
xnor U12880 (N_12880,N_10599,N_11760);
nand U12881 (N_12881,N_9508,N_9538);
nand U12882 (N_12882,N_10647,N_9986);
and U12883 (N_12883,N_10623,N_9690);
xor U12884 (N_12884,N_10883,N_11723);
xnor U12885 (N_12885,N_12357,N_11584);
nor U12886 (N_12886,N_10037,N_12044);
and U12887 (N_12887,N_10591,N_12328);
nand U12888 (N_12888,N_11038,N_12188);
nand U12889 (N_12889,N_12421,N_11242);
nor U12890 (N_12890,N_10439,N_9744);
nor U12891 (N_12891,N_12080,N_10467);
nor U12892 (N_12892,N_11934,N_12377);
nand U12893 (N_12893,N_12227,N_10653);
xnor U12894 (N_12894,N_11009,N_12352);
or U12895 (N_12895,N_9415,N_11982);
xnor U12896 (N_12896,N_11830,N_10241);
xnor U12897 (N_12897,N_9983,N_11209);
nor U12898 (N_12898,N_10459,N_9727);
or U12899 (N_12899,N_9485,N_11338);
xor U12900 (N_12900,N_10745,N_12027);
nand U12901 (N_12901,N_9829,N_11276);
nand U12902 (N_12902,N_9585,N_10966);
nor U12903 (N_12903,N_11270,N_11579);
or U12904 (N_12904,N_10784,N_11311);
nor U12905 (N_12905,N_10646,N_11991);
and U12906 (N_12906,N_9861,N_10906);
or U12907 (N_12907,N_9778,N_11762);
and U12908 (N_12908,N_9670,N_11998);
and U12909 (N_12909,N_12097,N_12009);
nor U12910 (N_12910,N_11027,N_10164);
xor U12911 (N_12911,N_10938,N_12198);
nor U12912 (N_12912,N_12090,N_11530);
nor U12913 (N_12913,N_11362,N_11495);
xnor U12914 (N_12914,N_12245,N_12354);
nor U12915 (N_12915,N_11266,N_12282);
and U12916 (N_12916,N_10214,N_11304);
and U12917 (N_12917,N_11007,N_10728);
xnor U12918 (N_12918,N_10629,N_12230);
xnor U12919 (N_12919,N_9391,N_10014);
and U12920 (N_12920,N_12358,N_10398);
nand U12921 (N_12921,N_10756,N_11795);
and U12922 (N_12922,N_12103,N_12204);
xnor U12923 (N_12923,N_10028,N_11884);
and U12924 (N_12924,N_11827,N_12495);
nor U12925 (N_12925,N_10649,N_11669);
nand U12926 (N_12926,N_10752,N_10705);
or U12927 (N_12927,N_12074,N_10174);
xnor U12928 (N_12928,N_12420,N_10540);
or U12929 (N_12929,N_9611,N_10377);
or U12930 (N_12930,N_9901,N_11649);
xnor U12931 (N_12931,N_11078,N_11451);
xor U12932 (N_12932,N_12255,N_10874);
and U12933 (N_12933,N_11752,N_11314);
and U12934 (N_12934,N_10032,N_12193);
nand U12935 (N_12935,N_10793,N_9561);
or U12936 (N_12936,N_11983,N_9549);
or U12937 (N_12937,N_10865,N_11224);
or U12938 (N_12938,N_11851,N_11326);
nor U12939 (N_12939,N_12465,N_10358);
nand U12940 (N_12940,N_10862,N_9753);
or U12941 (N_12941,N_9881,N_11965);
nor U12942 (N_12942,N_9446,N_9631);
nor U12943 (N_12943,N_11804,N_12063);
nand U12944 (N_12944,N_11238,N_11652);
and U12945 (N_12945,N_9545,N_12376);
nor U12946 (N_12946,N_9459,N_10972);
nor U12947 (N_12947,N_10161,N_12177);
or U12948 (N_12948,N_10483,N_10312);
or U12949 (N_12949,N_12134,N_10210);
xor U12950 (N_12950,N_10478,N_11562);
nor U12951 (N_12951,N_10425,N_11325);
or U12952 (N_12952,N_11907,N_10402);
or U12953 (N_12953,N_10696,N_11852);
nand U12954 (N_12954,N_9522,N_10684);
xor U12955 (N_12955,N_9637,N_11365);
xor U12956 (N_12956,N_11834,N_10665);
nand U12957 (N_12957,N_11917,N_9520);
nand U12958 (N_12958,N_9378,N_10044);
nor U12959 (N_12959,N_9702,N_11586);
nor U12960 (N_12960,N_10530,N_11687);
nand U12961 (N_12961,N_11115,N_11849);
and U12962 (N_12962,N_12248,N_10805);
and U12963 (N_12963,N_12380,N_11767);
nor U12964 (N_12964,N_11203,N_12489);
and U12965 (N_12965,N_11412,N_11862);
or U12966 (N_12966,N_11970,N_12187);
and U12967 (N_12967,N_12463,N_11857);
nand U12968 (N_12968,N_11053,N_10137);
and U12969 (N_12969,N_10963,N_9906);
or U12970 (N_12970,N_11831,N_10858);
xnor U12971 (N_12971,N_9743,N_11525);
nor U12972 (N_12972,N_10180,N_10000);
nor U12973 (N_12973,N_10719,N_10381);
or U12974 (N_12974,N_10635,N_10690);
or U12975 (N_12975,N_10167,N_12155);
xor U12976 (N_12976,N_10280,N_9974);
xnor U12977 (N_12977,N_10013,N_11461);
and U12978 (N_12978,N_12456,N_11910);
xor U12979 (N_12979,N_9993,N_12437);
xnor U12980 (N_12980,N_10065,N_10579);
and U12981 (N_12981,N_10316,N_12190);
or U12982 (N_12982,N_9919,N_11010);
or U12983 (N_12983,N_10897,N_11729);
and U12984 (N_12984,N_12035,N_10996);
nand U12985 (N_12985,N_11880,N_10886);
nor U12986 (N_12986,N_10053,N_9760);
nand U12987 (N_12987,N_10702,N_10245);
or U12988 (N_12988,N_9598,N_10261);
and U12989 (N_12989,N_10031,N_10730);
or U12990 (N_12990,N_10505,N_9407);
nand U12991 (N_12991,N_10826,N_11814);
xor U12992 (N_12992,N_12089,N_12462);
nor U12993 (N_12993,N_10577,N_11357);
or U12994 (N_12994,N_11747,N_10516);
nand U12995 (N_12995,N_10023,N_11308);
nor U12996 (N_12996,N_10675,N_11622);
or U12997 (N_12997,N_9624,N_11139);
and U12998 (N_12998,N_11793,N_11438);
and U12999 (N_12999,N_9412,N_11677);
nor U13000 (N_13000,N_12298,N_11505);
xnor U13001 (N_13001,N_9750,N_10871);
nor U13002 (N_13002,N_9582,N_11572);
nor U13003 (N_13003,N_10354,N_10236);
nand U13004 (N_13004,N_10218,N_12110);
xor U13005 (N_13005,N_10220,N_10195);
or U13006 (N_13006,N_9955,N_12077);
nand U13007 (N_13007,N_10482,N_11902);
or U13008 (N_13008,N_12483,N_12029);
and U13009 (N_13009,N_10821,N_12183);
and U13010 (N_13010,N_10608,N_12323);
and U13011 (N_13011,N_11054,N_12367);
nand U13012 (N_13012,N_10831,N_11411);
and U13013 (N_13013,N_11423,N_12273);
nand U13014 (N_13014,N_9552,N_10792);
and U13015 (N_13015,N_10276,N_12124);
xnor U13016 (N_13016,N_10597,N_9388);
or U13017 (N_13017,N_11818,N_11636);
and U13018 (N_13018,N_12220,N_9625);
nand U13019 (N_13019,N_11310,N_9854);
xnor U13020 (N_13020,N_10560,N_9929);
or U13021 (N_13021,N_11237,N_11730);
nor U13022 (N_13022,N_12179,N_10985);
and U13023 (N_13023,N_10927,N_11092);
and U13024 (N_13024,N_10352,N_11225);
xnor U13025 (N_13025,N_10746,N_12361);
or U13026 (N_13026,N_12387,N_12397);
or U13027 (N_13027,N_11952,N_10376);
nand U13028 (N_13028,N_12237,N_10385);
or U13029 (N_13029,N_9610,N_10845);
nand U13030 (N_13030,N_11548,N_11309);
nand U13031 (N_13031,N_10369,N_10787);
nand U13032 (N_13032,N_12036,N_11946);
or U13033 (N_13033,N_11372,N_12168);
nand U13034 (N_13034,N_12244,N_10040);
and U13035 (N_13035,N_10329,N_10612);
xnor U13036 (N_13036,N_10128,N_9464);
nor U13037 (N_13037,N_10620,N_11966);
xnor U13038 (N_13038,N_9865,N_11095);
xor U13039 (N_13039,N_10197,N_11685);
nand U13040 (N_13040,N_11207,N_10781);
nand U13041 (N_13041,N_9879,N_11504);
nand U13042 (N_13042,N_9599,N_10275);
xor U13043 (N_13043,N_11182,N_9528);
nor U13044 (N_13044,N_10438,N_9936);
xnor U13045 (N_13045,N_11528,N_10586);
xor U13046 (N_13046,N_11658,N_9645);
and U13047 (N_13047,N_9946,N_10567);
or U13048 (N_13048,N_11545,N_9418);
nand U13049 (N_13049,N_10243,N_10087);
and U13050 (N_13050,N_9692,N_11129);
or U13051 (N_13051,N_11216,N_11126);
nand U13052 (N_13052,N_11921,N_9836);
and U13053 (N_13053,N_9845,N_10674);
xor U13054 (N_13054,N_11187,N_9939);
or U13055 (N_13055,N_12163,N_10296);
or U13056 (N_13056,N_11206,N_11105);
nor U13057 (N_13057,N_11167,N_9550);
nand U13058 (N_13058,N_10140,N_10307);
and U13059 (N_13059,N_11444,N_11117);
nand U13060 (N_13060,N_10801,N_10983);
or U13061 (N_13061,N_10656,N_10998);
or U13062 (N_13062,N_11439,N_11204);
nor U13063 (N_13063,N_12406,N_12310);
nor U13064 (N_13064,N_10372,N_12186);
nand U13065 (N_13065,N_9496,N_12280);
nor U13066 (N_13066,N_10266,N_9393);
nand U13067 (N_13067,N_12492,N_10511);
xor U13068 (N_13068,N_11345,N_9989);
xor U13069 (N_13069,N_9774,N_11483);
or U13070 (N_13070,N_11514,N_9700);
xnor U13071 (N_13071,N_10463,N_11522);
and U13072 (N_13072,N_10273,N_12113);
and U13073 (N_13073,N_11046,N_11868);
nor U13074 (N_13074,N_12207,N_11563);
or U13075 (N_13075,N_10844,N_11389);
nor U13076 (N_13076,N_9853,N_10889);
nor U13077 (N_13077,N_11152,N_9384);
xnor U13078 (N_13078,N_11954,N_10293);
or U13079 (N_13079,N_10734,N_10182);
nor U13080 (N_13080,N_10595,N_10634);
xnor U13081 (N_13081,N_9927,N_10386);
or U13082 (N_13082,N_10476,N_10529);
and U13083 (N_13083,N_12411,N_9699);
xnor U13084 (N_13084,N_12130,N_9819);
nand U13085 (N_13085,N_9785,N_12251);
xor U13086 (N_13086,N_10553,N_9540);
nand U13087 (N_13087,N_9519,N_11773);
or U13088 (N_13088,N_10362,N_10717);
and U13089 (N_13089,N_10094,N_12060);
nand U13090 (N_13090,N_9695,N_10753);
xor U13091 (N_13091,N_9563,N_10854);
nor U13092 (N_13092,N_10936,N_9725);
and U13093 (N_13093,N_10626,N_11364);
or U13094 (N_13094,N_10303,N_11112);
or U13095 (N_13095,N_9995,N_11603);
nor U13096 (N_13096,N_11223,N_11465);
xnor U13097 (N_13097,N_9472,N_11267);
or U13098 (N_13098,N_11856,N_12491);
and U13099 (N_13099,N_10348,N_11672);
nor U13100 (N_13100,N_10257,N_11809);
or U13101 (N_13101,N_10903,N_9562);
nand U13102 (N_13102,N_12219,N_11241);
xor U13103 (N_13103,N_12281,N_11977);
nand U13104 (N_13104,N_9976,N_10494);
nand U13105 (N_13105,N_10281,N_11252);
or U13106 (N_13106,N_11626,N_12182);
nand U13107 (N_13107,N_9900,N_10120);
nor U13108 (N_13108,N_12484,N_10440);
nand U13109 (N_13109,N_10070,N_12095);
nand U13110 (N_13110,N_10770,N_10592);
or U13111 (N_13111,N_9716,N_11875);
and U13112 (N_13112,N_9537,N_9940);
xnor U13113 (N_13113,N_12470,N_11375);
nand U13114 (N_13114,N_11591,N_9674);
and U13115 (N_13115,N_10641,N_11564);
nor U13116 (N_13116,N_9498,N_12146);
or U13117 (N_13117,N_9873,N_10565);
nor U13118 (N_13118,N_11140,N_9581);
or U13119 (N_13119,N_9633,N_11201);
nand U13120 (N_13120,N_10893,N_12487);
nand U13121 (N_13121,N_12005,N_9641);
nor U13122 (N_13122,N_12435,N_10958);
nand U13123 (N_13123,N_10475,N_12482);
and U13124 (N_13124,N_11402,N_11068);
and U13125 (N_13125,N_12348,N_11768);
nor U13126 (N_13126,N_10990,N_10272);
and U13127 (N_13127,N_9984,N_12300);
nand U13128 (N_13128,N_11198,N_12041);
nand U13129 (N_13129,N_11190,N_10751);
or U13130 (N_13130,N_12392,N_11925);
nor U13131 (N_13131,N_9790,N_10017);
or U13132 (N_13132,N_12311,N_12457);
or U13133 (N_13133,N_11549,N_10811);
xnor U13134 (N_13134,N_10122,N_9830);
nor U13135 (N_13135,N_12304,N_11697);
nand U13136 (N_13136,N_11667,N_11149);
nand U13137 (N_13137,N_11026,N_10682);
xnor U13138 (N_13138,N_10624,N_10668);
nor U13139 (N_13139,N_11947,N_10412);
and U13140 (N_13140,N_10299,N_10502);
nand U13141 (N_13141,N_10513,N_12046);
xnor U13142 (N_13142,N_11887,N_12065);
and U13143 (N_13143,N_11937,N_11245);
nor U13144 (N_13144,N_11195,N_11306);
nor U13145 (N_13145,N_10355,N_11346);
and U13146 (N_13146,N_9944,N_11017);
xor U13147 (N_13147,N_10322,N_9634);
and U13148 (N_13148,N_11452,N_9798);
xor U13149 (N_13149,N_11544,N_12345);
or U13150 (N_13150,N_10361,N_10279);
nand U13151 (N_13151,N_11928,N_10112);
and U13152 (N_13152,N_11473,N_11066);
nand U13153 (N_13153,N_10956,N_10410);
or U13154 (N_13154,N_12330,N_9639);
nor U13155 (N_13155,N_10572,N_9630);
xnor U13156 (N_13156,N_12320,N_10708);
or U13157 (N_13157,N_9908,N_12342);
xnor U13158 (N_13158,N_9516,N_10791);
xnor U13159 (N_13159,N_10404,N_12295);
nor U13160 (N_13160,N_12301,N_12151);
nor U13161 (N_13161,N_10928,N_9607);
or U13162 (N_13162,N_9525,N_10300);
nand U13163 (N_13163,N_10773,N_9721);
xor U13164 (N_13164,N_12478,N_11400);
xnor U13165 (N_13165,N_12212,N_10146);
or U13166 (N_13166,N_11222,N_10817);
xor U13167 (N_13167,N_11750,N_9711);
nor U13168 (N_13168,N_9772,N_12129);
or U13169 (N_13169,N_9741,N_10660);
and U13170 (N_13170,N_10135,N_10934);
and U13171 (N_13171,N_10676,N_12254);
or U13172 (N_13172,N_10149,N_10993);
nand U13173 (N_13173,N_10481,N_11271);
nor U13174 (N_13174,N_11180,N_12283);
nor U13175 (N_13175,N_12241,N_10852);
nand U13176 (N_13176,N_11604,N_9622);
nand U13177 (N_13177,N_11551,N_9841);
nand U13178 (N_13178,N_11709,N_9462);
nand U13179 (N_13179,N_9783,N_9604);
and U13180 (N_13180,N_11629,N_11388);
xor U13181 (N_13181,N_10607,N_11327);
or U13182 (N_13182,N_10864,N_11558);
nand U13183 (N_13183,N_9923,N_11063);
or U13184 (N_13184,N_10962,N_9425);
nand U13185 (N_13185,N_12253,N_10603);
xor U13186 (N_13186,N_12426,N_11492);
or U13187 (N_13187,N_10050,N_11100);
and U13188 (N_13188,N_12189,N_9915);
nor U13189 (N_13189,N_10205,N_11289);
nand U13190 (N_13190,N_10548,N_9686);
and U13191 (N_13191,N_9886,N_11042);
and U13192 (N_13192,N_10206,N_12100);
nand U13193 (N_13193,N_12322,N_11599);
and U13194 (N_13194,N_12412,N_11409);
or U13195 (N_13195,N_10736,N_12475);
and U13196 (N_13196,N_10471,N_10426);
or U13197 (N_13197,N_9621,N_11874);
xor U13198 (N_13198,N_10803,N_12360);
and U13199 (N_13199,N_10869,N_11789);
xnor U13200 (N_13200,N_10103,N_12148);
and U13201 (N_13201,N_11269,N_12197);
nand U13202 (N_13202,N_11971,N_12170);
or U13203 (N_13203,N_9998,N_10047);
or U13204 (N_13204,N_10480,N_10301);
nand U13205 (N_13205,N_11737,N_11879);
and U13206 (N_13206,N_9487,N_10740);
nand U13207 (N_13207,N_10506,N_10931);
and U13208 (N_13208,N_12087,N_9737);
and U13209 (N_13209,N_10922,N_11174);
nand U13210 (N_13210,N_10600,N_9401);
xnor U13211 (N_13211,N_11715,N_11430);
xor U13212 (N_13212,N_9736,N_10396);
nor U13213 (N_13213,N_10867,N_11832);
and U13214 (N_13214,N_12020,N_9867);
and U13215 (N_13215,N_10571,N_10650);
and U13216 (N_13216,N_11350,N_9510);
and U13217 (N_13217,N_11690,N_10898);
xnor U13218 (N_13218,N_9697,N_10216);
nand U13219 (N_13219,N_10406,N_10418);
and U13220 (N_13220,N_10709,N_11556);
or U13221 (N_13221,N_10399,N_11445);
xor U13222 (N_13222,N_10517,N_9970);
nand U13223 (N_13223,N_11153,N_11487);
or U13224 (N_13224,N_11580,N_11277);
xor U13225 (N_13225,N_10574,N_11783);
nor U13226 (N_13226,N_12417,N_11170);
and U13227 (N_13227,N_9456,N_12499);
and U13228 (N_13228,N_9440,N_10680);
or U13229 (N_13229,N_12422,N_11177);
or U13230 (N_13230,N_12257,N_10692);
nand U13231 (N_13231,N_10491,N_10772);
xor U13232 (N_13232,N_12429,N_10485);
and U13233 (N_13233,N_12018,N_11926);
nor U13234 (N_13234,N_10810,N_11419);
and U13235 (N_13235,N_9530,N_11488);
nor U13236 (N_13236,N_10252,N_10503);
and U13237 (N_13237,N_11333,N_12346);
and U13238 (N_13238,N_11185,N_11349);
nor U13239 (N_13239,N_10964,N_12022);
nor U13240 (N_13240,N_11116,N_11541);
and U13241 (N_13241,N_12040,N_11000);
nor U13242 (N_13242,N_11469,N_9535);
nor U13243 (N_13243,N_12038,N_10628);
or U13244 (N_13244,N_10297,N_12128);
and U13245 (N_13245,N_11537,N_9404);
or U13246 (N_13246,N_12313,N_11191);
nor U13247 (N_13247,N_11997,N_9557);
xnor U13248 (N_13248,N_9958,N_11507);
nand U13249 (N_13249,N_10384,N_11097);
xor U13250 (N_13250,N_11587,N_11573);
nand U13251 (N_13251,N_10126,N_10658);
nor U13252 (N_13252,N_10196,N_10263);
nand U13253 (N_13253,N_11039,N_10583);
and U13254 (N_13254,N_11259,N_11128);
nand U13255 (N_13255,N_10045,N_11655);
nand U13256 (N_13256,N_11749,N_10436);
or U13257 (N_13257,N_12032,N_12158);
xor U13258 (N_13258,N_10657,N_11840);
nand U13259 (N_13259,N_11956,N_11463);
xor U13260 (N_13260,N_9930,N_11360);
nand U13261 (N_13261,N_11246,N_11692);
xor U13262 (N_13262,N_10742,N_11458);
or U13263 (N_13263,N_9430,N_9956);
nand U13264 (N_13264,N_9385,N_11532);
and U13265 (N_13265,N_9463,N_12199);
or U13266 (N_13266,N_11745,N_11996);
nor U13267 (N_13267,N_12427,N_9846);
and U13268 (N_13268,N_10202,N_11102);
xnor U13269 (N_13269,N_10104,N_12016);
nand U13270 (N_13270,N_10244,N_9584);
nor U13271 (N_13271,N_9981,N_10292);
xnor U13272 (N_13272,N_10115,N_11317);
nand U13273 (N_13273,N_10732,N_10401);
xnor U13274 (N_13274,N_10490,N_10010);
nor U13275 (N_13275,N_11536,N_10298);
xnor U13276 (N_13276,N_11637,N_10796);
xnor U13277 (N_13277,N_12068,N_11999);
xnor U13278 (N_13278,N_10788,N_10059);
or U13279 (N_13279,N_10507,N_9580);
or U13280 (N_13280,N_10191,N_10328);
nand U13281 (N_13281,N_11381,N_10556);
and U13282 (N_13282,N_10849,N_10515);
xor U13283 (N_13283,N_9416,N_12454);
xor U13284 (N_13284,N_9653,N_9554);
or U13285 (N_13285,N_10550,N_12374);
xor U13286 (N_13286,N_11990,N_9583);
and U13287 (N_13287,N_10535,N_10170);
and U13288 (N_13288,N_11331,N_10847);
xnor U13289 (N_13289,N_11786,N_9458);
and U13290 (N_13290,N_9817,N_9838);
nor U13291 (N_13291,N_12262,N_11539);
nand U13292 (N_13292,N_11268,N_10239);
or U13293 (N_13293,N_10652,N_11797);
xor U13294 (N_13294,N_12173,N_11016);
or U13295 (N_13295,N_11485,N_9696);
or U13296 (N_13296,N_9869,N_11136);
and U13297 (N_13297,N_11218,N_11272);
and U13298 (N_13298,N_9876,N_9539);
or U13299 (N_13299,N_11923,N_10733);
nor U13300 (N_13300,N_11006,N_11540);
xnor U13301 (N_13301,N_10681,N_12321);
xor U13302 (N_13302,N_11253,N_10939);
nor U13303 (N_13303,N_10912,N_10514);
nand U13304 (N_13304,N_12432,N_10973);
or U13305 (N_13305,N_11316,N_10189);
nand U13306 (N_13306,N_9757,N_9488);
and U13307 (N_13307,N_11968,N_9399);
nor U13308 (N_13308,N_12115,N_9669);
xnor U13309 (N_13309,N_12045,N_10171);
nand U13310 (N_13310,N_11466,N_11108);
or U13311 (N_13311,N_12261,N_11467);
and U13312 (N_13312,N_10913,N_12175);
or U13313 (N_13313,N_10738,N_9654);
xor U13314 (N_13314,N_12384,N_12102);
and U13315 (N_13315,N_11263,N_10422);
and U13316 (N_13316,N_11708,N_9531);
nand U13317 (N_13317,N_11656,N_9606);
xor U13318 (N_13318,N_10270,N_11256);
xor U13319 (N_13319,N_9954,N_11848);
nand U13320 (N_13320,N_11638,N_11686);
or U13321 (N_13321,N_11221,N_9897);
nor U13322 (N_13322,N_9724,N_10609);
or U13323 (N_13323,N_11062,N_9465);
and U13324 (N_13324,N_9943,N_10432);
and U13325 (N_13325,N_10596,N_11646);
xnor U13326 (N_13326,N_9574,N_10413);
nand U13327 (N_13327,N_11008,N_11756);
or U13328 (N_13328,N_12167,N_10335);
nand U13329 (N_13329,N_11434,N_9600);
nor U13330 (N_13330,N_11778,N_11219);
xnor U13331 (N_13331,N_11861,N_10915);
nand U13332 (N_13332,N_10259,N_9945);
and U13333 (N_13333,N_12156,N_12147);
nand U13334 (N_13334,N_9635,N_11867);
or U13335 (N_13335,N_9423,N_12049);
or U13336 (N_13336,N_12171,N_10366);
nand U13337 (N_13337,N_9457,N_9439);
xor U13338 (N_13338,N_10022,N_11759);
or U13339 (N_13339,N_10073,N_11377);
nor U13340 (N_13340,N_10981,N_9735);
or U13341 (N_13341,N_12086,N_11144);
xor U13342 (N_13342,N_10814,N_11711);
and U13343 (N_13343,N_9821,N_10557);
xor U13344 (N_13344,N_9902,N_9417);
nand U13345 (N_13345,N_10616,N_10812);
xor U13346 (N_13346,N_9629,N_11403);
nand U13347 (N_13347,N_10056,N_11264);
and U13348 (N_13348,N_9612,N_12351);
nor U13349 (N_13349,N_11501,N_11305);
and U13350 (N_13350,N_11236,N_10131);
and U13351 (N_13351,N_11700,N_10068);
and U13352 (N_13352,N_10537,N_9529);
or U13353 (N_13353,N_10666,N_11023);
and U13354 (N_13354,N_11771,N_11127);
xor U13355 (N_13355,N_11076,N_9618);
and U13356 (N_13356,N_11109,N_12308);
xnor U13357 (N_13357,N_9651,N_9636);
nand U13358 (N_13358,N_11499,N_11293);
and U13359 (N_13359,N_10622,N_9985);
and U13360 (N_13360,N_12181,N_10445);
or U13361 (N_13361,N_12256,N_12117);
xor U13362 (N_13362,N_11691,N_11618);
or U13363 (N_13363,N_9680,N_11987);
and U13364 (N_13364,N_10286,N_10066);
nand U13365 (N_13365,N_11871,N_9453);
nand U13366 (N_13366,N_10832,N_9375);
nor U13367 (N_13367,N_10707,N_11114);
xor U13368 (N_13368,N_12091,N_9691);
and U13369 (N_13369,N_11543,N_11694);
and U13370 (N_13370,N_10111,N_11918);
nor U13371 (N_13371,N_10466,N_10724);
nor U13372 (N_13372,N_9748,N_11414);
nor U13373 (N_13373,N_11213,N_12356);
nand U13374 (N_13374,N_11892,N_10544);
nor U13375 (N_13375,N_11476,N_10081);
and U13376 (N_13376,N_11909,N_12368);
nor U13377 (N_13377,N_11019,N_11621);
xor U13378 (N_13378,N_10238,N_10881);
nor U13379 (N_13379,N_12085,N_11378);
xor U13380 (N_13380,N_12126,N_9402);
nand U13381 (N_13381,N_10343,N_11091);
or U13382 (N_13382,N_12111,N_11408);
nand U13383 (N_13383,N_10663,N_12332);
or U13384 (N_13384,N_12098,N_10255);
xnor U13385 (N_13385,N_9579,N_11820);
nor U13386 (N_13386,N_12398,N_9438);
nand U13387 (N_13387,N_9796,N_10855);
nor U13388 (N_13388,N_12271,N_11617);
nor U13389 (N_13389,N_12458,N_11748);
or U13390 (N_13390,N_11069,N_10274);
or U13391 (N_13391,N_10083,N_11202);
nand U13392 (N_13392,N_10391,N_9461);
or U13393 (N_13393,N_11980,N_12246);
nand U13394 (N_13394,N_10217,N_10349);
and U13395 (N_13395,N_10346,N_11554);
xnor U13396 (N_13396,N_10701,N_11594);
nor U13397 (N_13397,N_11226,N_11577);
and U13398 (N_13398,N_11992,N_12125);
or U13399 (N_13399,N_10012,N_10347);
nand U13400 (N_13400,N_10192,N_10940);
or U13401 (N_13401,N_11689,N_11494);
nor U13402 (N_13402,N_11725,N_12419);
or U13403 (N_13403,N_11353,N_10948);
xor U13404 (N_13404,N_9979,N_11757);
nor U13405 (N_13405,N_11571,N_9776);
nor U13406 (N_13406,N_11456,N_9558);
xor U13407 (N_13407,N_10763,N_12133);
xor U13408 (N_13408,N_12178,N_9891);
and U13409 (N_13409,N_11435,N_10223);
nand U13410 (N_13410,N_10201,N_10489);
nand U13411 (N_13411,N_11679,N_9746);
nand U13412 (N_13412,N_11047,N_11387);
nor U13413 (N_13413,N_12343,N_12132);
and U13414 (N_13414,N_11678,N_11478);
and U13415 (N_13415,N_9427,N_9626);
xor U13416 (N_13416,N_11176,N_11057);
and U13417 (N_13417,N_11482,N_11810);
nor U13418 (N_13418,N_11052,N_9857);
xor U13419 (N_13419,N_11858,N_10175);
or U13420 (N_13420,N_10937,N_11738);
xnor U13421 (N_13421,N_12109,N_10373);
xor U13422 (N_13422,N_11576,N_9499);
and U13423 (N_13423,N_10365,N_10130);
and U13424 (N_13424,N_11683,N_11960);
nor U13425 (N_13425,N_10390,N_12440);
and U13426 (N_13426,N_11720,N_10670);
or U13427 (N_13427,N_11067,N_9977);
and U13428 (N_13428,N_11426,N_11569);
nor U13429 (N_13429,N_10879,N_10986);
nand U13430 (N_13430,N_10703,N_11089);
and U13431 (N_13431,N_10789,N_12226);
nor U13432 (N_13432,N_9848,N_10106);
xnor U13433 (N_13433,N_11985,N_10551);
and U13434 (N_13434,N_11070,N_10357);
nand U13435 (N_13435,N_10630,N_10645);
nor U13436 (N_13436,N_11836,N_10430);
or U13437 (N_13437,N_11624,N_12275);
xor U13438 (N_13438,N_9784,N_9536);
xor U13439 (N_13439,N_10437,N_11535);
nor U13440 (N_13440,N_11151,N_12092);
or U13441 (N_13441,N_9780,N_9920);
xnor U13442 (N_13442,N_10991,N_9526);
xnor U13443 (N_13443,N_10078,N_12430);
or U13444 (N_13444,N_11348,N_12378);
and U13445 (N_13445,N_10926,N_11654);
xnor U13446 (N_13446,N_10213,N_10039);
xnor U13447 (N_13447,N_9501,N_11845);
nand U13448 (N_13448,N_11941,N_10492);
nor U13449 (N_13449,N_12268,N_12334);
xnor U13450 (N_13450,N_10423,N_12061);
nand U13451 (N_13451,N_11164,N_12096);
or U13452 (N_13452,N_11648,N_10890);
or U13453 (N_13453,N_10839,N_10338);
nor U13454 (N_13454,N_11590,N_10688);
or U13455 (N_13455,N_9511,N_11796);
nand U13456 (N_13456,N_12249,N_11370);
nand U13457 (N_13457,N_11184,N_11974);
or U13458 (N_13458,N_10387,N_9883);
xor U13459 (N_13459,N_12467,N_12002);
and U13460 (N_13460,N_9450,N_12481);
and U13461 (N_13461,N_10559,N_9909);
nor U13462 (N_13462,N_11651,N_11630);
nor U13463 (N_13463,N_9755,N_10549);
or U13464 (N_13464,N_12438,N_11973);
or U13465 (N_13465,N_11860,N_10290);
nor U13466 (N_13466,N_11812,N_10001);
nor U13467 (N_13467,N_12391,N_12405);
or U13468 (N_13468,N_11634,N_10061);
xnor U13469 (N_13469,N_10230,N_9726);
xnor U13470 (N_13470,N_10907,N_12118);
or U13471 (N_13471,N_11410,N_12287);
and U13472 (N_13472,N_9548,N_11320);
nand U13473 (N_13473,N_10759,N_10113);
xnor U13474 (N_13474,N_9966,N_9560);
nand U13475 (N_13475,N_11142,N_11696);
and U13476 (N_13476,N_10621,N_9870);
or U13477 (N_13477,N_10052,N_9822);
and U13478 (N_13478,N_11989,N_10168);
nor U13479 (N_13479,N_9442,N_12371);
or U13480 (N_13480,N_12277,N_10456);
or U13481 (N_13481,N_12407,N_10999);
nor U13482 (N_13482,N_9834,N_12488);
nor U13483 (N_13483,N_11765,N_10064);
xnor U13484 (N_13484,N_11891,N_12047);
or U13485 (N_13485,N_9613,N_9863);
nor U13486 (N_13486,N_10486,N_10720);
xor U13487 (N_13487,N_10570,N_10509);
or U13488 (N_13488,N_10097,N_11775);
xnor U13489 (N_13489,N_12104,N_12479);
xnor U13490 (N_13490,N_11872,N_12494);
xnor U13491 (N_13491,N_11883,N_11988);
nand U13492 (N_13492,N_12259,N_10718);
nor U13493 (N_13493,N_11739,N_10896);
nand U13494 (N_13494,N_11429,N_10585);
nand U13495 (N_13495,N_11358,N_11468);
xnor U13496 (N_13496,N_9566,N_11197);
nand U13497 (N_13497,N_10287,N_9504);
or U13498 (N_13498,N_11938,N_9662);
nor U13499 (N_13499,N_12213,N_11298);
and U13500 (N_13500,N_9874,N_9882);
xnor U13501 (N_13501,N_11391,N_9502);
or U13502 (N_13502,N_10250,N_11313);
nor U13503 (N_13503,N_11520,N_12247);
xnor U13504 (N_13504,N_10581,N_11799);
and U13505 (N_13505,N_11995,N_11596);
or U13506 (N_13506,N_9812,N_11110);
or U13507 (N_13507,N_12099,N_11084);
and U13508 (N_13508,N_9421,N_9657);
or U13509 (N_13509,N_12064,N_11614);
nor U13510 (N_13510,N_12229,N_11763);
or U13511 (N_13511,N_10857,N_12442);
xnor U13512 (N_13512,N_10221,N_9503);
or U13513 (N_13513,N_9433,N_12340);
nand U13514 (N_13514,N_10284,N_10268);
or U13515 (N_13515,N_9740,N_10519);
and U13516 (N_13516,N_9578,N_11724);
nor U13517 (N_13517,N_9685,N_9596);
nor U13518 (N_13518,N_10659,N_12037);
xnor U13519 (N_13519,N_9643,N_9824);
xnor U13520 (N_13520,N_12403,N_9720);
xnor U13521 (N_13521,N_11287,N_10209);
xor U13522 (N_13522,N_9706,N_9795);
nor U13523 (N_13523,N_11096,N_11415);
nor U13524 (N_13524,N_9466,N_12264);
xor U13525 (N_13525,N_11332,N_11123);
xnor U13526 (N_13526,N_10957,N_10253);
or U13527 (N_13527,N_11022,N_9818);
or U13528 (N_13528,N_10807,N_11508);
and U13529 (N_13529,N_11668,N_12238);
or U13530 (N_13530,N_10891,N_9871);
and U13531 (N_13531,N_11282,N_11455);
or U13532 (N_13532,N_9987,N_12319);
xnor U13533 (N_13533,N_11436,N_11361);
nor U13534 (N_13534,N_11919,N_10378);
or U13535 (N_13535,N_10920,N_10842);
xnor U13536 (N_13536,N_9436,N_11726);
nand U13537 (N_13537,N_11030,N_12232);
and U13538 (N_13538,N_11173,N_11878);
or U13539 (N_13539,N_9773,N_9759);
and U13540 (N_13540,N_11772,N_10229);
xnor U13541 (N_13541,N_11645,N_11301);
xor U13542 (N_13542,N_9512,N_12472);
nand U13543 (N_13543,N_9928,N_9847);
nand U13544 (N_13544,N_11911,N_10970);
nand U13545 (N_13545,N_9479,N_10697);
and U13546 (N_13546,N_11247,N_10484);
and U13547 (N_13547,N_10142,N_9468);
nor U13548 (N_13548,N_11914,N_10782);
xnor U13549 (N_13549,N_9965,N_11321);
and U13550 (N_13550,N_10153,N_11734);
nand U13551 (N_13551,N_9693,N_10219);
nor U13552 (N_13552,N_10498,N_9470);
or U13553 (N_13553,N_11040,N_12083);
nor U13554 (N_13554,N_11640,N_9953);
nand U13555 (N_13555,N_10295,N_11088);
and U13556 (N_13556,N_9381,N_10523);
and U13557 (N_13557,N_12431,N_12337);
and U13558 (N_13558,N_11758,N_11405);
and U13559 (N_13559,N_11257,N_9555);
nand U13560 (N_13560,N_11813,N_9917);
nor U13561 (N_13561,N_11955,N_12031);
nor U13562 (N_13562,N_12402,N_11037);
nand U13563 (N_13563,N_10092,N_10138);
and U13564 (N_13564,N_11777,N_12314);
and U13565 (N_13565,N_10777,N_10370);
xor U13566 (N_13566,N_11021,N_9827);
nand U13567 (N_13567,N_9912,N_11183);
nor U13568 (N_13568,N_10868,N_10619);
or U13569 (N_13569,N_10447,N_12081);
xor U13570 (N_13570,N_10859,N_12265);
xor U13571 (N_13571,N_12184,N_11620);
and U13572 (N_13572,N_10512,N_11406);
xor U13573 (N_13573,N_10226,N_10339);
or U13574 (N_13574,N_12030,N_9615);
and U13575 (N_13575,N_10242,N_10302);
xor U13576 (N_13576,N_12127,N_12486);
or U13577 (N_13577,N_10769,N_11628);
nor U13578 (N_13578,N_10124,N_10363);
xor U13579 (N_13579,N_10995,N_11819);
xnor U13580 (N_13580,N_10723,N_10468);
or U13581 (N_13581,N_9849,N_9952);
or U13582 (N_13582,N_9937,N_9490);
nor U13583 (N_13583,N_10602,N_10564);
or U13584 (N_13584,N_12034,N_12326);
and U13585 (N_13585,N_11553,N_10541);
and U13586 (N_13586,N_11979,N_12067);
and U13587 (N_13587,N_11106,N_11693);
nor U13588 (N_13588,N_11920,N_9758);
nand U13589 (N_13589,N_10333,N_9664);
or U13590 (N_13590,N_11281,N_12468);
and U13591 (N_13591,N_12404,N_11583);
nor U13592 (N_13592,N_10743,N_12079);
nand U13593 (N_13593,N_11113,N_12290);
or U13594 (N_13594,N_11497,N_9999);
xor U13595 (N_13595,N_12054,N_11912);
nand U13596 (N_13596,N_10569,N_10790);
nand U13597 (N_13597,N_9448,N_11570);
nor U13598 (N_13598,N_9443,N_9523);
nand U13599 (N_13599,N_9926,N_10353);
nand U13600 (N_13600,N_11418,N_11699);
and U13601 (N_13601,N_12144,N_9815);
and U13602 (N_13602,N_12209,N_11728);
xor U13603 (N_13603,N_10419,N_11018);
or U13604 (N_13604,N_9617,N_10497);
nor U13605 (N_13605,N_10613,N_10538);
xor U13606 (N_13606,N_10700,N_11698);
xor U13607 (N_13607,N_11713,N_11500);
xnor U13608 (N_13608,N_10234,N_11984);
xor U13609 (N_13609,N_9842,N_9826);
xor U13610 (N_13610,N_11764,N_10786);
xor U13611 (N_13611,N_11766,N_12325);
or U13612 (N_13612,N_11719,N_9642);
xor U13613 (N_13613,N_11512,N_11660);
nand U13614 (N_13614,N_11821,N_11099);
or U13615 (N_13615,N_12162,N_10984);
or U13616 (N_13616,N_10158,N_12336);
and U13617 (N_13617,N_9890,N_10588);
and U13618 (N_13618,N_11141,N_11050);
and U13619 (N_13619,N_9679,N_10062);
nor U13620 (N_13620,N_10605,N_10691);
and U13621 (N_13621,N_9663,N_11602);
nand U13622 (N_13622,N_9792,N_12434);
or U13623 (N_13623,N_9708,N_11550);
xor U13624 (N_13624,N_9714,N_9968);
xor U13625 (N_13625,N_10580,N_10698);
or U13626 (N_13626,N_10224,N_10715);
nor U13627 (N_13627,N_12333,N_11424);
and U13628 (N_13628,N_11371,N_11625);
xor U13629 (N_13629,N_11742,N_11296);
and U13630 (N_13630,N_11366,N_9406);
nand U13631 (N_13631,N_12260,N_9931);
nor U13632 (N_13632,N_11850,N_12023);
nor U13633 (N_13633,N_10317,N_10314);
and U13634 (N_13634,N_12480,N_11924);
and U13635 (N_13635,N_10685,N_9771);
xnor U13636 (N_13636,N_11680,N_12474);
xnor U13637 (N_13637,N_10058,N_10661);
or U13638 (N_13638,N_11565,N_9947);
and U13639 (N_13639,N_10604,N_10582);
nand U13640 (N_13640,N_11839,N_9572);
xnor U13641 (N_13641,N_9969,N_10935);
or U13642 (N_13642,N_11044,N_12221);
or U13643 (N_13643,N_11906,N_11963);
nor U13644 (N_13644,N_11159,N_9650);
nor U13645 (N_13645,N_9386,N_10819);
xor U13646 (N_13646,N_10843,N_11337);
nand U13647 (N_13647,N_12466,N_12236);
nand U13648 (N_13648,N_9441,N_12225);
xnor U13649 (N_13649,N_11193,N_11355);
or U13650 (N_13650,N_10077,N_12414);
nand U13651 (N_13651,N_9913,N_11981);
xnor U13652 (N_13652,N_12122,N_11352);
nor U13653 (N_13653,N_10408,N_11279);
xnor U13654 (N_13654,N_11448,N_10687);
and U13655 (N_13655,N_10473,N_11442);
nor U13656 (N_13656,N_10994,N_11559);
xnor U13657 (N_13657,N_11449,N_10967);
and U13658 (N_13658,N_11386,N_12142);
nor U13659 (N_13659,N_12082,N_12393);
nor U13660 (N_13660,N_10977,N_10323);
xnor U13661 (N_13661,N_12135,N_11712);
or U13662 (N_13662,N_10208,N_10722);
nor U13663 (N_13663,N_10848,N_9668);
nand U13664 (N_13664,N_11404,N_9649);
nor U13665 (N_13665,N_9398,N_9605);
or U13666 (N_13666,N_12455,N_10693);
xor U13667 (N_13667,N_10054,N_9799);
nand U13668 (N_13668,N_10729,N_12243);
or U13669 (N_13669,N_11235,N_11015);
xnor U13670 (N_13670,N_11318,N_9527);
or U13671 (N_13671,N_10799,N_10651);
or U13672 (N_13672,N_11041,N_9547);
nand U13673 (N_13673,N_11120,N_11231);
xnor U13674 (N_13674,N_9801,N_10099);
nor U13675 (N_13675,N_11392,N_11899);
nand U13676 (N_13676,N_12307,N_10360);
and U13677 (N_13677,N_10818,N_11284);
or U13678 (N_13678,N_10193,N_10829);
and U13679 (N_13679,N_10640,N_10533);
or U13680 (N_13680,N_9951,N_9933);
and U13681 (N_13681,N_11215,N_9553);
xor U13682 (N_13682,N_12157,N_9567);
or U13683 (N_13683,N_11425,N_10677);
or U13684 (N_13684,N_11897,N_9935);
xor U13685 (N_13685,N_10380,N_11012);
or U13686 (N_13686,N_10248,N_11302);
and U13687 (N_13687,N_9895,N_10285);
xor U13688 (N_13688,N_10304,N_9910);
nand U13689 (N_13689,N_9660,N_11446);
and U13690 (N_13690,N_9991,N_11510);
or U13691 (N_13691,N_10536,N_10982);
nor U13692 (N_13692,N_10820,N_9875);
or U13693 (N_13693,N_9994,N_9495);
or U13694 (N_13694,N_10771,N_9597);
or U13695 (N_13695,N_9894,N_9619);
nand U13696 (N_13696,N_10020,N_11101);
nor U13697 (N_13697,N_11949,N_11186);
and U13698 (N_13698,N_12176,N_11323);
or U13699 (N_13699,N_9676,N_11496);
nor U13700 (N_13700,N_12108,N_10388);
xor U13701 (N_13701,N_9878,N_12006);
or U13702 (N_13702,N_11262,N_10644);
nor U13703 (N_13703,N_11791,N_10096);
xnor U13704 (N_13704,N_10955,N_11324);
and U13705 (N_13705,N_10278,N_11521);
or U13706 (N_13706,N_11518,N_9474);
and U13707 (N_13707,N_9652,N_10488);
nor U13708 (N_13708,N_11098,N_9709);
or U13709 (N_13709,N_11254,N_10851);
or U13710 (N_13710,N_10136,N_12042);
or U13711 (N_13711,N_9571,N_11189);
nand U13712 (N_13712,N_9980,N_10946);
or U13713 (N_13713,N_9832,N_11877);
or U13714 (N_13714,N_10741,N_11833);
nand U13715 (N_13715,N_12439,N_11157);
or U13716 (N_13716,N_12076,N_10636);
and U13717 (N_13717,N_11927,N_12138);
nand U13718 (N_13718,N_11916,N_9698);
nand U13719 (N_13719,N_12008,N_11462);
and U13720 (N_13720,N_12451,N_11605);
nand U13721 (N_13721,N_12305,N_12053);
nor U13722 (N_13722,N_11179,N_9896);
and U13723 (N_13723,N_12279,N_11143);
xnor U13724 (N_13724,N_11230,N_10198);
and U13725 (N_13725,N_9396,N_12139);
nand U13726 (N_13726,N_10457,N_11208);
or U13727 (N_13727,N_11131,N_12196);
xor U13728 (N_13728,N_11866,N_11382);
and U13729 (N_13729,N_12359,N_10762);
xnor U13730 (N_13730,N_9703,N_10573);
and U13731 (N_13731,N_10495,N_12373);
xor U13732 (N_13732,N_11894,N_9794);
or U13733 (N_13733,N_10908,N_11077);
and U13734 (N_13734,N_11650,N_11975);
or U13735 (N_13735,N_10587,N_10706);
nand U13736 (N_13736,N_12224,N_10265);
nor U13737 (N_13737,N_10063,N_10188);
nand U13738 (N_13738,N_10710,N_11258);
xor U13739 (N_13739,N_11481,N_9992);
or U13740 (N_13740,N_9704,N_11087);
xnor U13741 (N_13741,N_11959,N_10036);
or U13742 (N_13742,N_11517,N_11843);
or U13743 (N_13743,N_12493,N_11146);
and U13744 (N_13744,N_10091,N_10894);
and U13745 (N_13745,N_11578,N_11407);
nand U13746 (N_13746,N_9763,N_10667);
and U13747 (N_13747,N_11132,N_11045);
and U13748 (N_13748,N_12250,N_11229);
or U13749 (N_13749,N_12195,N_10143);
xnor U13750 (N_13750,N_9603,N_9934);
nor U13751 (N_13751,N_12350,N_12240);
and U13752 (N_13752,N_10015,N_12409);
and U13753 (N_13753,N_11676,N_11842);
xor U13754 (N_13754,N_12084,N_12150);
nand U13755 (N_13755,N_10453,N_12395);
nor U13756 (N_13756,N_10568,N_10169);
nor U13757 (N_13757,N_11781,N_11227);
nand U13758 (N_13758,N_11823,N_10959);
or U13759 (N_13759,N_11437,N_10464);
nand U13760 (N_13760,N_12274,N_10735);
and U13761 (N_13761,N_10055,N_11807);
or U13762 (N_13762,N_11623,N_11283);
nor U13763 (N_13763,N_9616,N_10704);
xor U13764 (N_13764,N_11329,N_10631);
or U13765 (N_13765,N_12242,N_9644);
nand U13766 (N_13766,N_9972,N_11239);
xor U13767 (N_13767,N_10960,N_10768);
nor U13768 (N_13768,N_11653,N_10833);
nand U13769 (N_13769,N_11703,N_11953);
xnor U13770 (N_13770,N_11427,N_11784);
or U13771 (N_13771,N_11363,N_10611);
or U13772 (N_13772,N_11800,N_12410);
and U13773 (N_13773,N_11704,N_12339);
and U13774 (N_13774,N_10417,N_10552);
or U13775 (N_13775,N_9828,N_9437);
nor U13776 (N_13776,N_9850,N_12347);
and U13777 (N_13777,N_10392,N_12007);
or U13778 (N_13778,N_9542,N_10856);
xor U13779 (N_13779,N_9964,N_12039);
nor U13780 (N_13780,N_10895,N_10783);
nand U13781 (N_13781,N_12445,N_12390);
nor U13782 (N_13782,N_11396,N_11285);
nand U13783 (N_13783,N_10679,N_11511);
nor U13784 (N_13784,N_11888,N_9905);
xor U13785 (N_13785,N_11417,N_10606);
and U13786 (N_13786,N_11161,N_9843);
nand U13787 (N_13787,N_10830,N_9805);
nand U13788 (N_13788,N_9684,N_11681);
or U13789 (N_13789,N_11632,N_10172);
nor U13790 (N_13790,N_10978,N_10246);
and U13791 (N_13791,N_9565,N_10929);
nand U13792 (N_13792,N_10578,N_10539);
xnor U13793 (N_13793,N_9855,N_11957);
or U13794 (N_13794,N_9705,N_11633);
nor U13795 (N_13795,N_12331,N_9573);
nor U13796 (N_13796,N_11886,N_10424);
or U13797 (N_13797,N_10151,N_11397);
xor U13798 (N_13798,N_12448,N_12174);
or U13799 (N_13799,N_9887,N_12364);
xor U13800 (N_13800,N_12052,N_10452);
xor U13801 (N_13801,N_9587,N_11533);
or U13802 (N_13802,N_10499,N_9454);
nor U13803 (N_13803,N_9570,N_10123);
and U13804 (N_13804,N_10341,N_10326);
nor U13805 (N_13805,N_12303,N_12394);
nand U13806 (N_13806,N_12312,N_9715);
nor U13807 (N_13807,N_10614,N_9837);
nor U13808 (N_13808,N_12381,N_11074);
or U13809 (N_13809,N_10525,N_10576);
and U13810 (N_13810,N_11049,N_10393);
xnor U13811 (N_13811,N_11740,N_10231);
and U13812 (N_13812,N_10760,N_12408);
or U13813 (N_13813,N_10531,N_9862);
nor U13814 (N_13814,N_9948,N_10215);
xor U13815 (N_13815,N_10019,N_11561);
nand U13816 (N_13816,N_11250,N_10767);
nor U13817 (N_13817,N_10200,N_10949);
nor U13818 (N_13818,N_11961,N_11744);
nor U13819 (N_13819,N_10090,N_9856);
xor U13820 (N_13820,N_11165,N_10232);
nor U13821 (N_13821,N_9814,N_11611);
nand U13822 (N_13822,N_12447,N_9506);
and U13823 (N_13823,N_11367,N_11220);
and U13824 (N_13824,N_11032,N_9623);
xnor U13825 (N_13825,N_9687,N_11673);
nor U13826 (N_13826,N_11755,N_12375);
xor U13827 (N_13827,N_9835,N_10165);
xor U13828 (N_13828,N_11048,N_11085);
nand U13829 (N_13829,N_10185,N_11641);
nor U13830 (N_13830,N_9559,N_10283);
nor U13831 (N_13831,N_10689,N_11383);
and U13832 (N_13832,N_10816,N_10892);
and U13833 (N_13833,N_10351,N_10669);
nor U13834 (N_13834,N_10884,N_10546);
or U13835 (N_13835,N_11011,N_10374);
nor U13836 (N_13836,N_10780,N_11931);
and U13837 (N_13837,N_10116,N_9728);
nor U13838 (N_13838,N_10846,N_12278);
nand U13839 (N_13839,N_11122,N_10965);
and U13840 (N_13840,N_10407,N_12015);
nand U13841 (N_13841,N_11255,N_10367);
and U13842 (N_13842,N_10992,N_12011);
nor U13843 (N_13843,N_12363,N_9806);
xor U13844 (N_13844,N_11769,N_9781);
xnor U13845 (N_13845,N_11547,N_9717);
or U13846 (N_13846,N_12217,N_11670);
nand U13847 (N_13847,N_10095,N_9961);
or U13848 (N_13848,N_11825,N_12215);
or U13849 (N_13849,N_11682,N_12057);
and U13850 (N_13850,N_10003,N_11248);
and U13851 (N_13851,N_11422,N_9712);
or U13852 (N_13852,N_10448,N_11896);
and U13853 (N_13853,N_9608,N_11330);
or U13854 (N_13854,N_11134,N_9938);
or U13855 (N_13855,N_11552,N_11575);
and U13856 (N_13856,N_9452,N_10672);
and U13857 (N_13857,N_10493,N_12043);
nand U13858 (N_13858,N_10435,N_10487);
xnor U13859 (N_13859,N_12169,N_10909);
nor U13860 (N_13860,N_11589,N_10726);
nor U13861 (N_13861,N_9648,N_11431);
or U13862 (N_13862,N_12263,N_11199);
xor U13863 (N_13863,N_9556,N_10477);
xor U13864 (N_13864,N_11297,N_9770);
nor U13865 (N_13865,N_10267,N_10132);
and U13866 (N_13866,N_9950,N_10633);
xor U13867 (N_13867,N_11684,N_11978);
xnor U13868 (N_13868,N_11035,N_10835);
or U13869 (N_13869,N_10051,N_9844);
nand U13870 (N_13870,N_9767,N_11870);
and U13871 (N_13871,N_9809,N_12136);
nand U13872 (N_13872,N_11368,N_11033);
nand U13873 (N_13873,N_11627,N_11479);
xnor U13874 (N_13874,N_10382,N_12025);
nor U13875 (N_13875,N_11743,N_10181);
nor U13876 (N_13876,N_9486,N_12019);
and U13877 (N_13877,N_11421,N_10615);
or U13878 (N_13878,N_10007,N_10344);
xnor U13879 (N_13879,N_11181,N_12140);
xnor U13880 (N_13880,N_9761,N_11601);
nand U13881 (N_13881,N_9569,N_10194);
nor U13882 (N_13882,N_9591,N_9916);
and U13883 (N_13883,N_11915,N_10776);
and U13884 (N_13884,N_9754,N_11344);
xor U13885 (N_13885,N_11788,N_10953);
xnor U13886 (N_13886,N_11440,N_10800);
xnor U13887 (N_13887,N_11486,N_10914);
xnor U13888 (N_13888,N_11716,N_12372);
xnor U13889 (N_13889,N_11585,N_12028);
or U13890 (N_13890,N_10500,N_9493);
nor U13891 (N_13891,N_10853,N_10411);
xnor U13892 (N_13892,N_10671,N_9718);
or U13893 (N_13893,N_9387,N_10954);
and U13894 (N_13894,N_10713,N_11081);
and U13895 (N_13895,N_12362,N_11822);
nor U13896 (N_13896,N_11413,N_12276);
or U13897 (N_13897,N_11384,N_10618);
or U13898 (N_13898,N_11401,N_10921);
nand U13899 (N_13899,N_11598,N_10837);
nand U13900 (N_13900,N_12452,N_9484);
or U13901 (N_13901,N_10901,N_12450);
nand U13902 (N_13902,N_12389,N_12293);
and U13903 (N_13903,N_11335,N_9851);
nor U13904 (N_13904,N_11671,N_10093);
nand U13905 (N_13905,N_10049,N_10625);
and U13906 (N_13906,N_9769,N_9491);
nand U13907 (N_13907,N_10004,N_12001);
xor U13908 (N_13908,N_9431,N_9521);
nand U13909 (N_13909,N_10076,N_10755);
nand U13910 (N_13910,N_9515,N_10350);
or U13911 (N_13911,N_10156,N_9756);
nand U13912 (N_13912,N_11196,N_11291);
or U13913 (N_13913,N_10313,N_12114);
xor U13914 (N_13914,N_11433,N_10850);
xor U13915 (N_13915,N_9655,N_10757);
xor U13916 (N_13916,N_11555,N_9478);
and U13917 (N_13917,N_9627,N_11503);
nand U13918 (N_13918,N_10309,N_10204);
and U13919 (N_13919,N_12185,N_12073);
nor U13920 (N_13920,N_11546,N_9707);
nand U13921 (N_13921,N_9733,N_10911);
or U13922 (N_13922,N_11059,N_12496);
or U13923 (N_13923,N_11498,N_11731);
xor U13924 (N_13924,N_10823,N_11967);
nor U13925 (N_13925,N_10203,N_10395);
and U13926 (N_13926,N_11705,N_12026);
nand U13927 (N_13927,N_10834,N_11770);
nor U13928 (N_13928,N_12388,N_9745);
nor U13929 (N_13929,N_9541,N_10442);
xor U13930 (N_13930,N_11162,N_9833);
nand U13931 (N_13931,N_9513,N_10108);
and U13932 (N_13932,N_9592,N_11133);
or U13933 (N_13933,N_10802,N_9885);
and U13934 (N_13934,N_9925,N_12180);
nand U13935 (N_13935,N_11020,N_9590);
xnor U13936 (N_13936,N_11774,N_10038);
nor U13937 (N_13937,N_12021,N_11124);
or U13938 (N_13938,N_10383,N_10319);
nor U13939 (N_13939,N_9689,N_10686);
nand U13940 (N_13940,N_11233,N_10555);
and U13941 (N_13941,N_12270,N_11710);
xnor U13942 (N_13942,N_10727,N_10766);
nand U13943 (N_13943,N_9804,N_11600);
nor U13944 (N_13944,N_10950,N_9392);
nand U13945 (N_13945,N_12235,N_10764);
nand U13946 (N_13946,N_12056,N_10306);
and U13947 (N_13947,N_10364,N_12137);
nand U13948 (N_13948,N_11702,N_11664);
xnor U13949 (N_13949,N_12216,N_11295);
nor U13950 (N_13950,N_9628,N_9469);
xnor U13951 (N_13951,N_10289,N_11490);
nor U13952 (N_13952,N_12292,N_10375);
xnor U13953 (N_13953,N_11816,N_10118);
or U13954 (N_13954,N_11779,N_10744);
xnor U13955 (N_13955,N_10342,N_12341);
or U13956 (N_13956,N_10443,N_10100);
or U13957 (N_13957,N_11260,N_10105);
nand U13958 (N_13958,N_11824,N_10119);
and U13959 (N_13959,N_10941,N_11794);
nor U13960 (N_13960,N_11826,N_12208);
and U13961 (N_13961,N_12296,N_11901);
or U13962 (N_13962,N_12062,N_12473);
and U13963 (N_13963,N_11121,N_12441);
nor U13964 (N_13964,N_9640,N_10006);
nor U13965 (N_13965,N_10902,N_12477);
or U13966 (N_13966,N_9903,N_12055);
nand U13967 (N_13967,N_10924,N_10288);
and U13968 (N_13968,N_11347,N_10639);
xnor U13969 (N_13969,N_10102,N_11792);
or U13970 (N_13970,N_11688,N_9688);
or U13971 (N_13971,N_9477,N_12072);
nand U13972 (N_13972,N_9659,N_10139);
nand U13973 (N_13973,N_10617,N_10974);
nor U13974 (N_13974,N_12355,N_9492);
or U13975 (N_13975,N_11154,N_12329);
and U13976 (N_13976,N_11004,N_10080);
xor U13977 (N_13977,N_9858,N_10416);
nand U13978 (N_13978,N_12149,N_11275);
nor U13979 (N_13979,N_9694,N_11945);
nand U13980 (N_13980,N_12228,N_11028);
xor U13981 (N_13981,N_10018,N_10089);
or U13982 (N_13982,N_11138,N_10521);
nand U13983 (N_13983,N_11334,N_9914);
xor U13984 (N_13984,N_9646,N_9480);
and U13985 (N_13985,N_11118,N_10461);
or U13986 (N_13986,N_11560,N_9949);
and U13987 (N_13987,N_10254,N_10332);
xnor U13988 (N_13988,N_12141,N_11890);
and U13989 (N_13989,N_9904,N_11441);
and U13990 (N_13990,N_10872,N_10980);
or U13991 (N_13991,N_10638,N_12461);
nor U13992 (N_13992,N_12327,N_11619);
nand U13993 (N_13993,N_11593,N_11913);
and U13994 (N_13994,N_10925,N_11491);
and U13995 (N_13995,N_12223,N_11003);
xor U13996 (N_13996,N_9786,N_11072);
and U13997 (N_13997,N_10277,N_10524);
nor U13998 (N_13998,N_11002,N_10258);
nor U13999 (N_13999,N_11829,N_11613);
xor U14000 (N_14000,N_11055,N_11516);
or U14001 (N_14001,N_9564,N_10110);
xor U14002 (N_14002,N_9481,N_10575);
nand U14003 (N_14003,N_12070,N_10462);
or U14004 (N_14004,N_9614,N_10627);
and U14005 (N_14005,N_9888,N_9918);
and U14006 (N_14006,N_9723,N_12443);
xor U14007 (N_14007,N_9866,N_11390);
xnor U14008 (N_14008,N_9471,N_9810);
nand U14009 (N_14009,N_11459,N_10496);
and U14010 (N_14010,N_12446,N_9751);
and U14011 (N_14011,N_11722,N_9475);
nor U14012 (N_14012,N_9807,N_12365);
nor U14013 (N_14013,N_10048,N_10212);
nor U14014 (N_14014,N_9765,N_11339);
xnor U14015 (N_14015,N_12433,N_10543);
xor U14016 (N_14016,N_11607,N_10237);
or U14017 (N_14017,N_12299,N_9710);
nor U14018 (N_14018,N_9811,N_9620);
nand U14019 (N_14019,N_11464,N_11484);
nand U14020 (N_14020,N_10310,N_9739);
xor U14021 (N_14021,N_12106,N_10024);
or U14022 (N_14022,N_9500,N_12309);
and U14023 (N_14023,N_12418,N_9647);
xor U14024 (N_14024,N_9924,N_10072);
xor U14025 (N_14025,N_9435,N_9864);
xnor U14026 (N_14026,N_10716,N_11024);
nor U14027 (N_14027,N_11014,N_10678);
and U14028 (N_14028,N_10860,N_12286);
and U14029 (N_14029,N_10394,N_11290);
nor U14030 (N_14030,N_10542,N_9782);
nand U14031 (N_14031,N_10190,N_9507);
and U14032 (N_14032,N_11075,N_9546);
xnor U14033 (N_14033,N_10315,N_10952);
and U14034 (N_14034,N_9732,N_10025);
and U14035 (N_14035,N_10154,N_11265);
nor U14036 (N_14036,N_10431,N_9609);
or U14037 (N_14037,N_11736,N_12338);
nand U14038 (N_14038,N_11663,N_9839);
xor U14039 (N_14039,N_10458,N_10117);
nor U14040 (N_14040,N_10968,N_12272);
nand U14041 (N_14041,N_10337,N_10228);
and U14042 (N_14042,N_10562,N_12498);
nor U14043 (N_14043,N_12105,N_12203);
nand U14044 (N_14044,N_11379,N_9543);
xnor U14045 (N_14045,N_10930,N_10282);
or U14046 (N_14046,N_12288,N_9734);
and U14047 (N_14047,N_11904,N_10504);
xnor U14048 (N_14048,N_10861,N_10809);
xnor U14049 (N_14049,N_10256,N_11200);
nor U14050 (N_14050,N_12119,N_12116);
nand U14051 (N_14051,N_9942,N_11160);
or U14052 (N_14052,N_10166,N_10144);
nor U14053 (N_14053,N_11001,N_11294);
nor U14054 (N_14054,N_9577,N_11086);
or U14055 (N_14055,N_11509,N_11013);
xor U14056 (N_14056,N_12416,N_10420);
and U14057 (N_14057,N_11080,N_11782);
and U14058 (N_14058,N_12400,N_11336);
xnor U14059 (N_14059,N_10330,N_10547);
nand U14060 (N_14060,N_11094,N_11107);
nor U14061 (N_14061,N_11932,N_11635);
or U14062 (N_14062,N_11083,N_11344);
and U14063 (N_14063,N_11875,N_10983);
nor U14064 (N_14064,N_10756,N_10008);
nor U14065 (N_14065,N_10324,N_9380);
xor U14066 (N_14066,N_11685,N_12400);
nand U14067 (N_14067,N_9991,N_11470);
nor U14068 (N_14068,N_10424,N_9631);
xnor U14069 (N_14069,N_9486,N_10711);
nand U14070 (N_14070,N_11716,N_10098);
or U14071 (N_14071,N_12188,N_11358);
xnor U14072 (N_14072,N_9965,N_10304);
nor U14073 (N_14073,N_12196,N_12189);
nor U14074 (N_14074,N_11874,N_10859);
nand U14075 (N_14075,N_11482,N_12497);
xor U14076 (N_14076,N_10141,N_12268);
or U14077 (N_14077,N_10013,N_11584);
xor U14078 (N_14078,N_10417,N_10997);
nor U14079 (N_14079,N_10210,N_11771);
and U14080 (N_14080,N_10758,N_10451);
xnor U14081 (N_14081,N_10894,N_10691);
nand U14082 (N_14082,N_9511,N_11490);
nand U14083 (N_14083,N_10664,N_11600);
nor U14084 (N_14084,N_10093,N_10012);
nand U14085 (N_14085,N_10795,N_10925);
xnor U14086 (N_14086,N_10435,N_11145);
xor U14087 (N_14087,N_9443,N_11048);
and U14088 (N_14088,N_12463,N_11047);
or U14089 (N_14089,N_12252,N_10340);
nor U14090 (N_14090,N_10925,N_10706);
and U14091 (N_14091,N_10741,N_10253);
or U14092 (N_14092,N_11707,N_11804);
nor U14093 (N_14093,N_11100,N_11318);
nor U14094 (N_14094,N_12338,N_10262);
nor U14095 (N_14095,N_10092,N_10660);
nor U14096 (N_14096,N_11804,N_11284);
and U14097 (N_14097,N_10147,N_10273);
and U14098 (N_14098,N_9567,N_11982);
nor U14099 (N_14099,N_9830,N_12407);
xnor U14100 (N_14100,N_11553,N_11749);
and U14101 (N_14101,N_9762,N_11756);
xor U14102 (N_14102,N_12290,N_11896);
or U14103 (N_14103,N_11526,N_11572);
xnor U14104 (N_14104,N_11894,N_10021);
and U14105 (N_14105,N_11275,N_11442);
nor U14106 (N_14106,N_10444,N_10916);
and U14107 (N_14107,N_11534,N_11688);
and U14108 (N_14108,N_9407,N_10843);
or U14109 (N_14109,N_12251,N_10384);
nor U14110 (N_14110,N_11555,N_11335);
xor U14111 (N_14111,N_11878,N_10331);
and U14112 (N_14112,N_10423,N_10904);
xor U14113 (N_14113,N_9393,N_10069);
xnor U14114 (N_14114,N_11501,N_9635);
and U14115 (N_14115,N_11500,N_11820);
nand U14116 (N_14116,N_10463,N_10779);
nor U14117 (N_14117,N_11889,N_11618);
nor U14118 (N_14118,N_11293,N_11603);
xnor U14119 (N_14119,N_11357,N_11040);
nand U14120 (N_14120,N_11148,N_10213);
xnor U14121 (N_14121,N_9644,N_9453);
or U14122 (N_14122,N_10933,N_10738);
xor U14123 (N_14123,N_10364,N_10268);
and U14124 (N_14124,N_11078,N_11322);
xor U14125 (N_14125,N_9539,N_12329);
nand U14126 (N_14126,N_10353,N_11624);
nor U14127 (N_14127,N_9396,N_9410);
or U14128 (N_14128,N_11091,N_10101);
xor U14129 (N_14129,N_12228,N_9797);
xnor U14130 (N_14130,N_12076,N_10279);
or U14131 (N_14131,N_10825,N_9827);
nand U14132 (N_14132,N_9859,N_10165);
and U14133 (N_14133,N_10809,N_11168);
xnor U14134 (N_14134,N_10458,N_10906);
nand U14135 (N_14135,N_10818,N_10507);
nand U14136 (N_14136,N_9819,N_10536);
or U14137 (N_14137,N_9966,N_11466);
and U14138 (N_14138,N_11999,N_10679);
xor U14139 (N_14139,N_9811,N_9896);
and U14140 (N_14140,N_11412,N_10361);
and U14141 (N_14141,N_9726,N_10026);
or U14142 (N_14142,N_9764,N_11893);
nand U14143 (N_14143,N_11665,N_11348);
nor U14144 (N_14144,N_10719,N_9395);
xor U14145 (N_14145,N_11130,N_12420);
nor U14146 (N_14146,N_11347,N_12048);
or U14147 (N_14147,N_10431,N_11537);
and U14148 (N_14148,N_10015,N_10330);
or U14149 (N_14149,N_9597,N_10278);
or U14150 (N_14150,N_12268,N_11111);
xnor U14151 (N_14151,N_11246,N_11741);
or U14152 (N_14152,N_10366,N_11749);
xor U14153 (N_14153,N_11286,N_11901);
or U14154 (N_14154,N_11330,N_11839);
xor U14155 (N_14155,N_10433,N_10988);
nor U14156 (N_14156,N_9977,N_9591);
nand U14157 (N_14157,N_10012,N_10563);
nor U14158 (N_14158,N_11589,N_10012);
and U14159 (N_14159,N_10186,N_10086);
nand U14160 (N_14160,N_10071,N_10394);
nand U14161 (N_14161,N_11932,N_10505);
nand U14162 (N_14162,N_9490,N_9465);
nor U14163 (N_14163,N_12274,N_12432);
xor U14164 (N_14164,N_12107,N_12368);
xor U14165 (N_14165,N_9761,N_11077);
and U14166 (N_14166,N_11329,N_10766);
or U14167 (N_14167,N_11678,N_9397);
nand U14168 (N_14168,N_10199,N_12180);
nand U14169 (N_14169,N_12412,N_11872);
xnor U14170 (N_14170,N_10814,N_11454);
nor U14171 (N_14171,N_10558,N_10302);
nor U14172 (N_14172,N_9491,N_10371);
xnor U14173 (N_14173,N_12474,N_11406);
and U14174 (N_14174,N_11566,N_11214);
xnor U14175 (N_14175,N_11280,N_12093);
nand U14176 (N_14176,N_11122,N_11328);
and U14177 (N_14177,N_11175,N_10872);
and U14178 (N_14178,N_10062,N_12016);
or U14179 (N_14179,N_9375,N_10124);
nor U14180 (N_14180,N_9931,N_11891);
or U14181 (N_14181,N_10777,N_10562);
xnor U14182 (N_14182,N_10653,N_10907);
nand U14183 (N_14183,N_11285,N_11461);
nand U14184 (N_14184,N_12010,N_11655);
nor U14185 (N_14185,N_10564,N_12365);
nor U14186 (N_14186,N_10806,N_9749);
nand U14187 (N_14187,N_11913,N_11928);
and U14188 (N_14188,N_10592,N_11129);
xor U14189 (N_14189,N_10857,N_11102);
nand U14190 (N_14190,N_12481,N_10775);
and U14191 (N_14191,N_10242,N_12137);
nor U14192 (N_14192,N_10996,N_10533);
xor U14193 (N_14193,N_9396,N_11512);
nor U14194 (N_14194,N_9987,N_10226);
or U14195 (N_14195,N_12292,N_10273);
and U14196 (N_14196,N_11942,N_10924);
xnor U14197 (N_14197,N_11863,N_11222);
nor U14198 (N_14198,N_12266,N_11066);
or U14199 (N_14199,N_11549,N_10270);
or U14200 (N_14200,N_11461,N_10317);
or U14201 (N_14201,N_9538,N_10693);
or U14202 (N_14202,N_10152,N_9720);
xnor U14203 (N_14203,N_9848,N_9985);
nor U14204 (N_14204,N_9514,N_12403);
and U14205 (N_14205,N_11767,N_10883);
or U14206 (N_14206,N_10115,N_9799);
or U14207 (N_14207,N_9426,N_10491);
nand U14208 (N_14208,N_11810,N_10918);
nand U14209 (N_14209,N_9673,N_12022);
nand U14210 (N_14210,N_12217,N_11710);
and U14211 (N_14211,N_11060,N_9544);
nand U14212 (N_14212,N_11703,N_10691);
nand U14213 (N_14213,N_9963,N_9432);
nor U14214 (N_14214,N_12350,N_10058);
nor U14215 (N_14215,N_12243,N_10963);
nor U14216 (N_14216,N_10437,N_9628);
xnor U14217 (N_14217,N_10996,N_10723);
or U14218 (N_14218,N_10738,N_10789);
or U14219 (N_14219,N_10012,N_10442);
or U14220 (N_14220,N_9992,N_11454);
xnor U14221 (N_14221,N_9766,N_12257);
or U14222 (N_14222,N_9862,N_10004);
nand U14223 (N_14223,N_10563,N_10627);
nand U14224 (N_14224,N_10322,N_11274);
or U14225 (N_14225,N_11809,N_10930);
and U14226 (N_14226,N_11541,N_9617);
or U14227 (N_14227,N_10315,N_10116);
and U14228 (N_14228,N_9606,N_10356);
nor U14229 (N_14229,N_10115,N_9716);
nor U14230 (N_14230,N_12217,N_11904);
nand U14231 (N_14231,N_11450,N_10910);
nand U14232 (N_14232,N_11615,N_11741);
xor U14233 (N_14233,N_12154,N_11075);
nor U14234 (N_14234,N_9721,N_11829);
nor U14235 (N_14235,N_11103,N_10463);
or U14236 (N_14236,N_12000,N_11244);
or U14237 (N_14237,N_11047,N_11136);
and U14238 (N_14238,N_11014,N_11521);
and U14239 (N_14239,N_11062,N_10774);
or U14240 (N_14240,N_10332,N_11849);
xnor U14241 (N_14241,N_11298,N_11032);
nor U14242 (N_14242,N_9639,N_10862);
xor U14243 (N_14243,N_11514,N_11415);
nor U14244 (N_14244,N_11431,N_11474);
xor U14245 (N_14245,N_12266,N_9827);
or U14246 (N_14246,N_12085,N_11433);
and U14247 (N_14247,N_11359,N_10538);
and U14248 (N_14248,N_11302,N_10189);
xnor U14249 (N_14249,N_10052,N_12129);
nand U14250 (N_14250,N_11586,N_12317);
nor U14251 (N_14251,N_10327,N_11766);
nand U14252 (N_14252,N_12106,N_10849);
nand U14253 (N_14253,N_12092,N_10654);
or U14254 (N_14254,N_11593,N_12335);
and U14255 (N_14255,N_10877,N_11218);
and U14256 (N_14256,N_12220,N_10013);
nand U14257 (N_14257,N_11764,N_9594);
and U14258 (N_14258,N_11534,N_11454);
xor U14259 (N_14259,N_12347,N_11675);
and U14260 (N_14260,N_12034,N_10569);
nand U14261 (N_14261,N_12104,N_12043);
xnor U14262 (N_14262,N_11960,N_9418);
or U14263 (N_14263,N_9590,N_10395);
nor U14264 (N_14264,N_10357,N_10127);
and U14265 (N_14265,N_11223,N_11136);
nor U14266 (N_14266,N_11442,N_9510);
nor U14267 (N_14267,N_10994,N_9601);
nand U14268 (N_14268,N_11863,N_10804);
and U14269 (N_14269,N_10371,N_12202);
or U14270 (N_14270,N_11283,N_11624);
or U14271 (N_14271,N_10694,N_12311);
and U14272 (N_14272,N_10630,N_11779);
nor U14273 (N_14273,N_10256,N_12135);
nand U14274 (N_14274,N_11734,N_11912);
or U14275 (N_14275,N_11553,N_11492);
and U14276 (N_14276,N_11312,N_11772);
or U14277 (N_14277,N_10404,N_10022);
nor U14278 (N_14278,N_9551,N_11315);
nor U14279 (N_14279,N_12197,N_9489);
nor U14280 (N_14280,N_12114,N_11973);
xor U14281 (N_14281,N_10092,N_11601);
and U14282 (N_14282,N_10768,N_11941);
and U14283 (N_14283,N_11050,N_9659);
or U14284 (N_14284,N_11872,N_11618);
nor U14285 (N_14285,N_10694,N_10234);
xnor U14286 (N_14286,N_10408,N_11259);
or U14287 (N_14287,N_11484,N_10541);
or U14288 (N_14288,N_10309,N_9643);
nand U14289 (N_14289,N_10322,N_10834);
nand U14290 (N_14290,N_11988,N_10238);
or U14291 (N_14291,N_11107,N_10327);
xor U14292 (N_14292,N_9897,N_10960);
xnor U14293 (N_14293,N_10475,N_11283);
or U14294 (N_14294,N_10659,N_11125);
or U14295 (N_14295,N_11503,N_9991);
xor U14296 (N_14296,N_12360,N_9890);
or U14297 (N_14297,N_10995,N_11092);
or U14298 (N_14298,N_11600,N_10275);
xor U14299 (N_14299,N_10762,N_11114);
or U14300 (N_14300,N_10827,N_11509);
xor U14301 (N_14301,N_9528,N_11185);
nor U14302 (N_14302,N_10652,N_10032);
xor U14303 (N_14303,N_10836,N_9893);
and U14304 (N_14304,N_9385,N_12081);
or U14305 (N_14305,N_10215,N_9849);
or U14306 (N_14306,N_11208,N_10649);
nor U14307 (N_14307,N_11092,N_10827);
and U14308 (N_14308,N_11102,N_9434);
nor U14309 (N_14309,N_9907,N_10512);
xor U14310 (N_14310,N_10739,N_11678);
and U14311 (N_14311,N_11166,N_9457);
and U14312 (N_14312,N_12265,N_9666);
nand U14313 (N_14313,N_10770,N_11103);
and U14314 (N_14314,N_9997,N_9863);
and U14315 (N_14315,N_11210,N_9816);
nor U14316 (N_14316,N_12221,N_9622);
xor U14317 (N_14317,N_11438,N_9909);
nand U14318 (N_14318,N_9649,N_12116);
and U14319 (N_14319,N_11935,N_9668);
and U14320 (N_14320,N_10363,N_10270);
nand U14321 (N_14321,N_9852,N_12059);
nor U14322 (N_14322,N_11792,N_9766);
or U14323 (N_14323,N_11405,N_10178);
xnor U14324 (N_14324,N_11488,N_10212);
nand U14325 (N_14325,N_12299,N_9570);
xor U14326 (N_14326,N_9649,N_11149);
or U14327 (N_14327,N_11215,N_11863);
and U14328 (N_14328,N_10133,N_11196);
and U14329 (N_14329,N_10226,N_11536);
nor U14330 (N_14330,N_12161,N_11205);
nand U14331 (N_14331,N_10195,N_11750);
or U14332 (N_14332,N_9773,N_12388);
and U14333 (N_14333,N_10335,N_11183);
xor U14334 (N_14334,N_11333,N_11228);
nand U14335 (N_14335,N_9651,N_11710);
nand U14336 (N_14336,N_11092,N_11305);
or U14337 (N_14337,N_11933,N_9393);
nor U14338 (N_14338,N_12398,N_9737);
nand U14339 (N_14339,N_11947,N_10357);
and U14340 (N_14340,N_11549,N_10149);
nand U14341 (N_14341,N_11073,N_11667);
and U14342 (N_14342,N_12440,N_10304);
or U14343 (N_14343,N_10737,N_11485);
nand U14344 (N_14344,N_11078,N_9961);
nand U14345 (N_14345,N_10908,N_11272);
nand U14346 (N_14346,N_10172,N_9674);
xor U14347 (N_14347,N_10556,N_10903);
nor U14348 (N_14348,N_9828,N_11737);
xnor U14349 (N_14349,N_12105,N_11276);
and U14350 (N_14350,N_9487,N_11237);
or U14351 (N_14351,N_11493,N_10458);
xor U14352 (N_14352,N_10807,N_9853);
nand U14353 (N_14353,N_9829,N_10827);
and U14354 (N_14354,N_10908,N_10281);
or U14355 (N_14355,N_10889,N_11064);
and U14356 (N_14356,N_11552,N_9611);
nor U14357 (N_14357,N_11139,N_10672);
nand U14358 (N_14358,N_10288,N_10227);
nor U14359 (N_14359,N_10508,N_10120);
nand U14360 (N_14360,N_12097,N_10627);
or U14361 (N_14361,N_9924,N_12117);
or U14362 (N_14362,N_10330,N_11377);
or U14363 (N_14363,N_11141,N_10930);
and U14364 (N_14364,N_11910,N_11762);
xor U14365 (N_14365,N_12269,N_11130);
nor U14366 (N_14366,N_11058,N_11847);
or U14367 (N_14367,N_9998,N_11811);
xor U14368 (N_14368,N_9901,N_11371);
nand U14369 (N_14369,N_10239,N_9793);
xor U14370 (N_14370,N_11331,N_10930);
xor U14371 (N_14371,N_11327,N_10387);
xor U14372 (N_14372,N_9930,N_12314);
and U14373 (N_14373,N_12372,N_10875);
and U14374 (N_14374,N_10985,N_11170);
nor U14375 (N_14375,N_12366,N_11803);
xor U14376 (N_14376,N_10519,N_12305);
nand U14377 (N_14377,N_11242,N_11367);
or U14378 (N_14378,N_9468,N_10575);
and U14379 (N_14379,N_11113,N_9689);
xor U14380 (N_14380,N_11712,N_11881);
nand U14381 (N_14381,N_11939,N_9428);
nor U14382 (N_14382,N_10934,N_10138);
nand U14383 (N_14383,N_11303,N_9924);
nor U14384 (N_14384,N_12112,N_11676);
xor U14385 (N_14385,N_11574,N_9556);
and U14386 (N_14386,N_10361,N_12171);
xor U14387 (N_14387,N_9685,N_12011);
nor U14388 (N_14388,N_11479,N_11454);
xnor U14389 (N_14389,N_11477,N_10534);
nand U14390 (N_14390,N_10076,N_12085);
nand U14391 (N_14391,N_11042,N_10056);
nand U14392 (N_14392,N_9585,N_11696);
or U14393 (N_14393,N_12346,N_11372);
nand U14394 (N_14394,N_9779,N_9560);
or U14395 (N_14395,N_10400,N_10150);
and U14396 (N_14396,N_12207,N_11756);
xor U14397 (N_14397,N_11991,N_12401);
nor U14398 (N_14398,N_10322,N_10667);
nor U14399 (N_14399,N_10947,N_11125);
and U14400 (N_14400,N_10699,N_10187);
and U14401 (N_14401,N_11781,N_10750);
xnor U14402 (N_14402,N_11102,N_9968);
xnor U14403 (N_14403,N_10082,N_11976);
and U14404 (N_14404,N_9746,N_11781);
nand U14405 (N_14405,N_11430,N_10011);
nand U14406 (N_14406,N_11496,N_12031);
and U14407 (N_14407,N_10941,N_12241);
xor U14408 (N_14408,N_10686,N_11152);
xor U14409 (N_14409,N_9753,N_11870);
nand U14410 (N_14410,N_11386,N_12406);
xnor U14411 (N_14411,N_11431,N_11632);
xor U14412 (N_14412,N_12178,N_10959);
and U14413 (N_14413,N_10794,N_10440);
and U14414 (N_14414,N_12401,N_11238);
or U14415 (N_14415,N_10268,N_10702);
nand U14416 (N_14416,N_11648,N_10361);
nor U14417 (N_14417,N_9677,N_10451);
nand U14418 (N_14418,N_11602,N_11087);
nor U14419 (N_14419,N_11324,N_12210);
nor U14420 (N_14420,N_10540,N_10870);
or U14421 (N_14421,N_10126,N_11669);
and U14422 (N_14422,N_10682,N_12361);
nor U14423 (N_14423,N_10750,N_11235);
nand U14424 (N_14424,N_9737,N_11893);
nand U14425 (N_14425,N_12146,N_11972);
or U14426 (N_14426,N_12288,N_9577);
nor U14427 (N_14427,N_10322,N_12032);
nor U14428 (N_14428,N_10683,N_12025);
nand U14429 (N_14429,N_11847,N_9743);
nand U14430 (N_14430,N_12370,N_9506);
nand U14431 (N_14431,N_11287,N_12064);
nor U14432 (N_14432,N_11410,N_10622);
nor U14433 (N_14433,N_12228,N_11840);
nor U14434 (N_14434,N_12283,N_11492);
nor U14435 (N_14435,N_9643,N_10641);
and U14436 (N_14436,N_10431,N_10422);
nand U14437 (N_14437,N_12336,N_10596);
xnor U14438 (N_14438,N_9675,N_10784);
nor U14439 (N_14439,N_10077,N_9532);
nor U14440 (N_14440,N_11068,N_9847);
nand U14441 (N_14441,N_10272,N_12047);
nor U14442 (N_14442,N_11928,N_9884);
and U14443 (N_14443,N_12437,N_9772);
or U14444 (N_14444,N_11354,N_9418);
xor U14445 (N_14445,N_11331,N_9984);
xor U14446 (N_14446,N_12319,N_11803);
or U14447 (N_14447,N_12400,N_9376);
nand U14448 (N_14448,N_12248,N_9722);
nand U14449 (N_14449,N_9723,N_10508);
nor U14450 (N_14450,N_10296,N_11594);
and U14451 (N_14451,N_10244,N_11272);
and U14452 (N_14452,N_11273,N_9605);
nand U14453 (N_14453,N_12047,N_10102);
and U14454 (N_14454,N_10480,N_10566);
nand U14455 (N_14455,N_9999,N_10478);
nor U14456 (N_14456,N_11012,N_12071);
nand U14457 (N_14457,N_12236,N_10997);
nor U14458 (N_14458,N_10568,N_9747);
nor U14459 (N_14459,N_12078,N_10436);
and U14460 (N_14460,N_11791,N_12179);
or U14461 (N_14461,N_11417,N_10458);
nand U14462 (N_14462,N_11899,N_9945);
xnor U14463 (N_14463,N_10399,N_10500);
or U14464 (N_14464,N_11123,N_11986);
and U14465 (N_14465,N_10767,N_12326);
and U14466 (N_14466,N_10069,N_9399);
xnor U14467 (N_14467,N_11389,N_10451);
nor U14468 (N_14468,N_9544,N_12158);
xnor U14469 (N_14469,N_9810,N_11393);
xor U14470 (N_14470,N_10360,N_12390);
or U14471 (N_14471,N_11544,N_10731);
nor U14472 (N_14472,N_9466,N_11537);
nor U14473 (N_14473,N_10717,N_9769);
xor U14474 (N_14474,N_11884,N_11224);
nand U14475 (N_14475,N_10075,N_9562);
nand U14476 (N_14476,N_9411,N_10955);
or U14477 (N_14477,N_12027,N_12459);
nand U14478 (N_14478,N_12318,N_11196);
nand U14479 (N_14479,N_11132,N_11447);
nor U14480 (N_14480,N_9971,N_12266);
nand U14481 (N_14481,N_10618,N_10522);
nor U14482 (N_14482,N_12132,N_12291);
xor U14483 (N_14483,N_11956,N_10524);
xor U14484 (N_14484,N_10601,N_10863);
or U14485 (N_14485,N_11363,N_10461);
xor U14486 (N_14486,N_11628,N_12100);
xor U14487 (N_14487,N_10822,N_10008);
nor U14488 (N_14488,N_9594,N_9512);
nor U14489 (N_14489,N_11420,N_11990);
and U14490 (N_14490,N_10019,N_11666);
nand U14491 (N_14491,N_10582,N_11735);
xor U14492 (N_14492,N_10701,N_11986);
xnor U14493 (N_14493,N_9927,N_12466);
nor U14494 (N_14494,N_10353,N_10940);
and U14495 (N_14495,N_11692,N_11140);
xnor U14496 (N_14496,N_9911,N_9418);
xnor U14497 (N_14497,N_9549,N_11174);
or U14498 (N_14498,N_10092,N_9727);
nor U14499 (N_14499,N_11055,N_12486);
and U14500 (N_14500,N_9984,N_12246);
nor U14501 (N_14501,N_9406,N_10181);
xor U14502 (N_14502,N_9753,N_10994);
xnor U14503 (N_14503,N_11502,N_10355);
nand U14504 (N_14504,N_12021,N_11468);
or U14505 (N_14505,N_12407,N_10107);
xnor U14506 (N_14506,N_12093,N_10472);
and U14507 (N_14507,N_11292,N_9904);
xor U14508 (N_14508,N_10793,N_9594);
xor U14509 (N_14509,N_10053,N_11924);
nand U14510 (N_14510,N_12149,N_10227);
xor U14511 (N_14511,N_9586,N_11873);
nand U14512 (N_14512,N_10137,N_12190);
nand U14513 (N_14513,N_9825,N_9721);
xor U14514 (N_14514,N_10806,N_12014);
nand U14515 (N_14515,N_11622,N_11836);
or U14516 (N_14516,N_10620,N_10093);
or U14517 (N_14517,N_12286,N_10580);
nor U14518 (N_14518,N_10417,N_11874);
or U14519 (N_14519,N_10538,N_11776);
xnor U14520 (N_14520,N_12248,N_9501);
or U14521 (N_14521,N_9999,N_11907);
or U14522 (N_14522,N_11952,N_11028);
nand U14523 (N_14523,N_12062,N_11112);
and U14524 (N_14524,N_10125,N_11804);
and U14525 (N_14525,N_11153,N_10874);
or U14526 (N_14526,N_12025,N_10770);
and U14527 (N_14527,N_12236,N_12287);
or U14528 (N_14528,N_9639,N_10490);
nor U14529 (N_14529,N_10594,N_11553);
nor U14530 (N_14530,N_10139,N_9547);
nand U14531 (N_14531,N_11892,N_9394);
nand U14532 (N_14532,N_12390,N_9860);
nand U14533 (N_14533,N_12170,N_9710);
and U14534 (N_14534,N_10331,N_12142);
xnor U14535 (N_14535,N_11839,N_10751);
or U14536 (N_14536,N_11549,N_10137);
nand U14537 (N_14537,N_10405,N_12102);
nor U14538 (N_14538,N_9536,N_11732);
nand U14539 (N_14539,N_11014,N_11998);
xnor U14540 (N_14540,N_11067,N_12041);
xnor U14541 (N_14541,N_12150,N_9615);
xnor U14542 (N_14542,N_11425,N_9512);
xor U14543 (N_14543,N_11575,N_9774);
nor U14544 (N_14544,N_10799,N_11919);
xnor U14545 (N_14545,N_11523,N_11426);
nor U14546 (N_14546,N_10198,N_10510);
nand U14547 (N_14547,N_12273,N_10214);
or U14548 (N_14548,N_10926,N_11705);
nor U14549 (N_14549,N_10639,N_10143);
nand U14550 (N_14550,N_12223,N_11043);
nor U14551 (N_14551,N_10306,N_11249);
nor U14552 (N_14552,N_11645,N_9687);
nor U14553 (N_14553,N_11380,N_12262);
nor U14554 (N_14554,N_11976,N_9931);
xor U14555 (N_14555,N_10566,N_10983);
nand U14556 (N_14556,N_9531,N_12263);
nor U14557 (N_14557,N_11722,N_11052);
nor U14558 (N_14558,N_10753,N_10268);
nor U14559 (N_14559,N_10622,N_11601);
or U14560 (N_14560,N_10651,N_10785);
or U14561 (N_14561,N_12113,N_11580);
nand U14562 (N_14562,N_10516,N_9973);
or U14563 (N_14563,N_12164,N_11949);
nor U14564 (N_14564,N_11308,N_11156);
or U14565 (N_14565,N_11538,N_11300);
xor U14566 (N_14566,N_10713,N_11009);
nor U14567 (N_14567,N_11300,N_9898);
xor U14568 (N_14568,N_11352,N_10126);
xor U14569 (N_14569,N_11418,N_12429);
nor U14570 (N_14570,N_9917,N_10667);
and U14571 (N_14571,N_12414,N_12266);
nand U14572 (N_14572,N_11981,N_10485);
nor U14573 (N_14573,N_10906,N_10030);
or U14574 (N_14574,N_11576,N_11384);
xnor U14575 (N_14575,N_9377,N_10859);
or U14576 (N_14576,N_9438,N_10875);
nor U14577 (N_14577,N_12378,N_11661);
and U14578 (N_14578,N_12160,N_11649);
nand U14579 (N_14579,N_9913,N_9978);
nand U14580 (N_14580,N_11743,N_9960);
and U14581 (N_14581,N_11140,N_12495);
nand U14582 (N_14582,N_12148,N_9866);
or U14583 (N_14583,N_9737,N_11759);
xnor U14584 (N_14584,N_12141,N_11161);
nor U14585 (N_14585,N_9409,N_9500);
or U14586 (N_14586,N_11167,N_12041);
or U14587 (N_14587,N_9994,N_12199);
xor U14588 (N_14588,N_12226,N_10701);
nor U14589 (N_14589,N_11151,N_11652);
xor U14590 (N_14590,N_11309,N_9848);
nand U14591 (N_14591,N_9494,N_11209);
xor U14592 (N_14592,N_11131,N_11880);
nor U14593 (N_14593,N_10014,N_10215);
or U14594 (N_14594,N_11307,N_11364);
xor U14595 (N_14595,N_11527,N_9952);
and U14596 (N_14596,N_9730,N_9636);
xnor U14597 (N_14597,N_11843,N_9504);
nand U14598 (N_14598,N_10998,N_10103);
xnor U14599 (N_14599,N_11808,N_11680);
xnor U14600 (N_14600,N_10177,N_10977);
nand U14601 (N_14601,N_10602,N_9757);
or U14602 (N_14602,N_11232,N_12117);
xor U14603 (N_14603,N_11701,N_10555);
and U14604 (N_14604,N_12318,N_9545);
or U14605 (N_14605,N_10435,N_9972);
and U14606 (N_14606,N_11975,N_12066);
xor U14607 (N_14607,N_11085,N_11569);
or U14608 (N_14608,N_12422,N_10334);
nor U14609 (N_14609,N_9818,N_11969);
nand U14610 (N_14610,N_10597,N_11612);
nor U14611 (N_14611,N_10011,N_11832);
and U14612 (N_14612,N_11353,N_10203);
nand U14613 (N_14613,N_10667,N_9662);
xnor U14614 (N_14614,N_12080,N_12229);
nand U14615 (N_14615,N_11207,N_11551);
xor U14616 (N_14616,N_10352,N_9460);
nand U14617 (N_14617,N_11659,N_11565);
and U14618 (N_14618,N_12273,N_10331);
and U14619 (N_14619,N_12279,N_11914);
and U14620 (N_14620,N_12195,N_11023);
xnor U14621 (N_14621,N_11448,N_11515);
or U14622 (N_14622,N_11059,N_11691);
nor U14623 (N_14623,N_12473,N_10175);
xor U14624 (N_14624,N_11504,N_9766);
nand U14625 (N_14625,N_10168,N_9664);
and U14626 (N_14626,N_11146,N_11632);
nand U14627 (N_14627,N_12164,N_11934);
nor U14628 (N_14628,N_10575,N_9390);
xor U14629 (N_14629,N_9988,N_9911);
xnor U14630 (N_14630,N_9892,N_10900);
xnor U14631 (N_14631,N_9992,N_9599);
and U14632 (N_14632,N_9502,N_10406);
or U14633 (N_14633,N_10696,N_10138);
and U14634 (N_14634,N_12462,N_10772);
and U14635 (N_14635,N_9795,N_10509);
nor U14636 (N_14636,N_10438,N_12341);
xnor U14637 (N_14637,N_11055,N_11899);
nand U14638 (N_14638,N_10910,N_11048);
or U14639 (N_14639,N_9745,N_10151);
xnor U14640 (N_14640,N_11733,N_10470);
xor U14641 (N_14641,N_12462,N_12333);
or U14642 (N_14642,N_10371,N_11972);
xnor U14643 (N_14643,N_9803,N_12346);
xnor U14644 (N_14644,N_11152,N_11562);
xnor U14645 (N_14645,N_9802,N_12253);
nor U14646 (N_14646,N_10795,N_12084);
and U14647 (N_14647,N_9967,N_11942);
xnor U14648 (N_14648,N_10975,N_10309);
nand U14649 (N_14649,N_9708,N_10467);
xor U14650 (N_14650,N_11971,N_10502);
and U14651 (N_14651,N_9862,N_11096);
or U14652 (N_14652,N_9822,N_12399);
nand U14653 (N_14653,N_11830,N_11647);
or U14654 (N_14654,N_10324,N_11139);
nor U14655 (N_14655,N_11409,N_10822);
nand U14656 (N_14656,N_12097,N_11943);
or U14657 (N_14657,N_9823,N_10308);
nand U14658 (N_14658,N_12303,N_9624);
nand U14659 (N_14659,N_10966,N_10470);
and U14660 (N_14660,N_9599,N_10722);
and U14661 (N_14661,N_9409,N_9568);
nand U14662 (N_14662,N_10864,N_10853);
or U14663 (N_14663,N_10948,N_11161);
nor U14664 (N_14664,N_12324,N_9458);
and U14665 (N_14665,N_12214,N_10323);
or U14666 (N_14666,N_9692,N_10349);
nor U14667 (N_14667,N_11970,N_10254);
or U14668 (N_14668,N_11454,N_11640);
xnor U14669 (N_14669,N_11970,N_12479);
xor U14670 (N_14670,N_10919,N_12341);
or U14671 (N_14671,N_10069,N_10603);
nor U14672 (N_14672,N_10156,N_10042);
and U14673 (N_14673,N_10027,N_10763);
and U14674 (N_14674,N_10738,N_10265);
or U14675 (N_14675,N_10515,N_12376);
and U14676 (N_14676,N_12129,N_11964);
and U14677 (N_14677,N_9790,N_12360);
nand U14678 (N_14678,N_12297,N_12075);
xor U14679 (N_14679,N_12120,N_10157);
nand U14680 (N_14680,N_10823,N_11846);
nor U14681 (N_14681,N_11411,N_11561);
or U14682 (N_14682,N_9505,N_9375);
nand U14683 (N_14683,N_11268,N_9503);
nand U14684 (N_14684,N_9787,N_11431);
xor U14685 (N_14685,N_10448,N_11784);
nand U14686 (N_14686,N_11584,N_10450);
nor U14687 (N_14687,N_12209,N_11157);
xnor U14688 (N_14688,N_9843,N_9599);
xor U14689 (N_14689,N_10848,N_12430);
or U14690 (N_14690,N_10629,N_12169);
nand U14691 (N_14691,N_11020,N_11209);
and U14692 (N_14692,N_11975,N_10340);
and U14693 (N_14693,N_9393,N_10473);
nand U14694 (N_14694,N_11403,N_10500);
or U14695 (N_14695,N_10721,N_11412);
nor U14696 (N_14696,N_10148,N_10855);
nor U14697 (N_14697,N_11329,N_9647);
nand U14698 (N_14698,N_11150,N_10387);
nor U14699 (N_14699,N_9493,N_9943);
and U14700 (N_14700,N_11728,N_9491);
xnor U14701 (N_14701,N_11721,N_12494);
nand U14702 (N_14702,N_11934,N_12009);
and U14703 (N_14703,N_9426,N_11253);
or U14704 (N_14704,N_12100,N_11995);
and U14705 (N_14705,N_11100,N_11409);
nor U14706 (N_14706,N_12269,N_10926);
xnor U14707 (N_14707,N_11825,N_11090);
or U14708 (N_14708,N_10947,N_10212);
xor U14709 (N_14709,N_9996,N_9641);
and U14710 (N_14710,N_9987,N_11198);
xor U14711 (N_14711,N_9645,N_10279);
xor U14712 (N_14712,N_11046,N_9597);
and U14713 (N_14713,N_11749,N_11212);
and U14714 (N_14714,N_12293,N_10103);
nand U14715 (N_14715,N_11560,N_11940);
and U14716 (N_14716,N_11196,N_12168);
nand U14717 (N_14717,N_9619,N_10933);
nor U14718 (N_14718,N_11052,N_9819);
and U14719 (N_14719,N_11949,N_12071);
xnor U14720 (N_14720,N_11793,N_11705);
nand U14721 (N_14721,N_12430,N_11899);
or U14722 (N_14722,N_11081,N_10853);
nand U14723 (N_14723,N_12172,N_11952);
xnor U14724 (N_14724,N_10280,N_9826);
or U14725 (N_14725,N_11883,N_12112);
and U14726 (N_14726,N_10790,N_11767);
and U14727 (N_14727,N_10157,N_9907);
xor U14728 (N_14728,N_10698,N_10192);
xnor U14729 (N_14729,N_10180,N_10322);
nor U14730 (N_14730,N_11454,N_10749);
nor U14731 (N_14731,N_9716,N_9952);
xor U14732 (N_14732,N_9401,N_11194);
xnor U14733 (N_14733,N_10664,N_10929);
and U14734 (N_14734,N_10047,N_12379);
nor U14735 (N_14735,N_10114,N_9730);
and U14736 (N_14736,N_9575,N_9713);
xor U14737 (N_14737,N_10331,N_10345);
nor U14738 (N_14738,N_11186,N_11131);
nand U14739 (N_14739,N_9549,N_11470);
nor U14740 (N_14740,N_11528,N_11817);
xor U14741 (N_14741,N_11862,N_10220);
nand U14742 (N_14742,N_9795,N_9538);
or U14743 (N_14743,N_11465,N_9694);
or U14744 (N_14744,N_10726,N_11223);
or U14745 (N_14745,N_11126,N_12083);
nand U14746 (N_14746,N_10717,N_10021);
or U14747 (N_14747,N_10235,N_10658);
nand U14748 (N_14748,N_11376,N_11730);
nor U14749 (N_14749,N_11063,N_10341);
nand U14750 (N_14750,N_11282,N_9785);
xor U14751 (N_14751,N_11014,N_12113);
or U14752 (N_14752,N_10801,N_10602);
or U14753 (N_14753,N_11577,N_12079);
or U14754 (N_14754,N_11822,N_9702);
xor U14755 (N_14755,N_12033,N_11349);
and U14756 (N_14756,N_10543,N_12352);
nand U14757 (N_14757,N_12063,N_10880);
xor U14758 (N_14758,N_11263,N_10645);
nor U14759 (N_14759,N_12260,N_9477);
xor U14760 (N_14760,N_11566,N_9384);
xnor U14761 (N_14761,N_10842,N_11046);
nor U14762 (N_14762,N_9745,N_12208);
nand U14763 (N_14763,N_11361,N_12126);
xnor U14764 (N_14764,N_10326,N_11941);
or U14765 (N_14765,N_11833,N_9696);
or U14766 (N_14766,N_10338,N_11585);
and U14767 (N_14767,N_9416,N_11466);
nor U14768 (N_14768,N_10998,N_12089);
nand U14769 (N_14769,N_11705,N_11637);
xnor U14770 (N_14770,N_10785,N_10212);
nor U14771 (N_14771,N_9445,N_10091);
nand U14772 (N_14772,N_9675,N_11578);
and U14773 (N_14773,N_11919,N_9462);
nand U14774 (N_14774,N_12039,N_12357);
nand U14775 (N_14775,N_10228,N_9654);
and U14776 (N_14776,N_11205,N_11816);
xor U14777 (N_14777,N_10708,N_9630);
and U14778 (N_14778,N_11201,N_11896);
nor U14779 (N_14779,N_10742,N_10562);
nor U14780 (N_14780,N_11819,N_10135);
or U14781 (N_14781,N_11692,N_9742);
or U14782 (N_14782,N_12289,N_9437);
nor U14783 (N_14783,N_11970,N_10683);
or U14784 (N_14784,N_11193,N_11232);
nor U14785 (N_14785,N_12249,N_11231);
nor U14786 (N_14786,N_10328,N_9605);
and U14787 (N_14787,N_10548,N_12125);
nor U14788 (N_14788,N_11649,N_11802);
xnor U14789 (N_14789,N_9678,N_9835);
xnor U14790 (N_14790,N_9863,N_11180);
nor U14791 (N_14791,N_12068,N_10876);
nand U14792 (N_14792,N_12006,N_9660);
nand U14793 (N_14793,N_10560,N_11888);
xor U14794 (N_14794,N_11688,N_9557);
nand U14795 (N_14795,N_11881,N_10578);
nor U14796 (N_14796,N_11414,N_10875);
and U14797 (N_14797,N_11349,N_12419);
nand U14798 (N_14798,N_10107,N_9395);
nand U14799 (N_14799,N_12294,N_11198);
nand U14800 (N_14800,N_11045,N_10813);
or U14801 (N_14801,N_12496,N_10272);
or U14802 (N_14802,N_10095,N_10792);
and U14803 (N_14803,N_9915,N_11458);
xnor U14804 (N_14804,N_12496,N_10880);
and U14805 (N_14805,N_11820,N_10122);
nor U14806 (N_14806,N_12346,N_10721);
and U14807 (N_14807,N_12374,N_11526);
nor U14808 (N_14808,N_11283,N_10780);
xor U14809 (N_14809,N_10400,N_10814);
nand U14810 (N_14810,N_12203,N_12062);
and U14811 (N_14811,N_11914,N_10864);
nor U14812 (N_14812,N_11496,N_9451);
xnor U14813 (N_14813,N_11230,N_10988);
or U14814 (N_14814,N_11882,N_11523);
nor U14815 (N_14815,N_10203,N_11630);
and U14816 (N_14816,N_12007,N_10711);
and U14817 (N_14817,N_12493,N_10445);
nor U14818 (N_14818,N_9813,N_10626);
or U14819 (N_14819,N_10349,N_10842);
nor U14820 (N_14820,N_11795,N_9591);
xor U14821 (N_14821,N_10613,N_10626);
or U14822 (N_14822,N_11376,N_9563);
and U14823 (N_14823,N_9721,N_11965);
nor U14824 (N_14824,N_11194,N_10174);
and U14825 (N_14825,N_11929,N_10218);
or U14826 (N_14826,N_9719,N_11878);
nand U14827 (N_14827,N_10115,N_12076);
nand U14828 (N_14828,N_9922,N_11597);
or U14829 (N_14829,N_10106,N_12246);
nor U14830 (N_14830,N_11445,N_9648);
nor U14831 (N_14831,N_11997,N_10833);
xnor U14832 (N_14832,N_10520,N_11958);
nor U14833 (N_14833,N_11725,N_11570);
or U14834 (N_14834,N_11104,N_9733);
nor U14835 (N_14835,N_11773,N_11107);
nand U14836 (N_14836,N_10277,N_10434);
and U14837 (N_14837,N_10572,N_10512);
nor U14838 (N_14838,N_10744,N_11439);
xor U14839 (N_14839,N_10852,N_12245);
or U14840 (N_14840,N_11243,N_12233);
nor U14841 (N_14841,N_12377,N_12168);
and U14842 (N_14842,N_9974,N_11824);
or U14843 (N_14843,N_11840,N_11105);
nor U14844 (N_14844,N_12084,N_12003);
nor U14845 (N_14845,N_10196,N_10636);
or U14846 (N_14846,N_9953,N_9675);
xor U14847 (N_14847,N_12111,N_10169);
xnor U14848 (N_14848,N_12275,N_11733);
or U14849 (N_14849,N_10022,N_10828);
nand U14850 (N_14850,N_12035,N_11188);
nand U14851 (N_14851,N_10236,N_9719);
xnor U14852 (N_14852,N_11249,N_11024);
and U14853 (N_14853,N_9865,N_12385);
xnor U14854 (N_14854,N_11320,N_12027);
or U14855 (N_14855,N_10822,N_12415);
xor U14856 (N_14856,N_11070,N_9559);
nor U14857 (N_14857,N_12237,N_11081);
nor U14858 (N_14858,N_9643,N_12377);
or U14859 (N_14859,N_9947,N_11520);
nand U14860 (N_14860,N_11896,N_9733);
and U14861 (N_14861,N_10794,N_9780);
nand U14862 (N_14862,N_10033,N_10346);
and U14863 (N_14863,N_11362,N_11197);
nor U14864 (N_14864,N_11154,N_12284);
nand U14865 (N_14865,N_11899,N_9934);
nand U14866 (N_14866,N_11471,N_10121);
nand U14867 (N_14867,N_10056,N_11527);
nand U14868 (N_14868,N_10652,N_9748);
or U14869 (N_14869,N_11092,N_10797);
and U14870 (N_14870,N_11634,N_11533);
nand U14871 (N_14871,N_11288,N_11617);
xnor U14872 (N_14872,N_10022,N_10463);
and U14873 (N_14873,N_11227,N_11054);
or U14874 (N_14874,N_11900,N_9904);
nand U14875 (N_14875,N_9380,N_9836);
xnor U14876 (N_14876,N_11594,N_12439);
nor U14877 (N_14877,N_11313,N_12430);
nor U14878 (N_14878,N_9385,N_12170);
or U14879 (N_14879,N_10097,N_12024);
nor U14880 (N_14880,N_11346,N_9625);
nor U14881 (N_14881,N_12170,N_10803);
nand U14882 (N_14882,N_9452,N_9882);
and U14883 (N_14883,N_9819,N_11331);
nor U14884 (N_14884,N_11070,N_11758);
nand U14885 (N_14885,N_10519,N_9510);
or U14886 (N_14886,N_11632,N_10030);
and U14887 (N_14887,N_11669,N_9894);
and U14888 (N_14888,N_11903,N_10018);
xnor U14889 (N_14889,N_10528,N_10728);
or U14890 (N_14890,N_11958,N_9463);
nand U14891 (N_14891,N_10966,N_12032);
and U14892 (N_14892,N_10497,N_9622);
or U14893 (N_14893,N_10981,N_10405);
nor U14894 (N_14894,N_10556,N_10565);
or U14895 (N_14895,N_12164,N_11701);
or U14896 (N_14896,N_9837,N_11960);
xor U14897 (N_14897,N_9934,N_9489);
and U14898 (N_14898,N_12290,N_11526);
or U14899 (N_14899,N_10383,N_10531);
and U14900 (N_14900,N_11614,N_11657);
or U14901 (N_14901,N_11978,N_12385);
nor U14902 (N_14902,N_11716,N_11958);
or U14903 (N_14903,N_10361,N_11083);
nor U14904 (N_14904,N_11690,N_12289);
or U14905 (N_14905,N_11471,N_10318);
or U14906 (N_14906,N_12296,N_9663);
or U14907 (N_14907,N_12365,N_9855);
nand U14908 (N_14908,N_9559,N_9421);
or U14909 (N_14909,N_10848,N_11773);
nor U14910 (N_14910,N_10888,N_11268);
or U14911 (N_14911,N_11498,N_12048);
xnor U14912 (N_14912,N_12018,N_12458);
or U14913 (N_14913,N_10473,N_11718);
nor U14914 (N_14914,N_9646,N_12005);
nor U14915 (N_14915,N_12196,N_10492);
and U14916 (N_14916,N_10356,N_12269);
nand U14917 (N_14917,N_11494,N_12342);
and U14918 (N_14918,N_12446,N_11007);
xnor U14919 (N_14919,N_9560,N_11204);
nor U14920 (N_14920,N_9517,N_9654);
and U14921 (N_14921,N_9744,N_11774);
xor U14922 (N_14922,N_9500,N_11105);
or U14923 (N_14923,N_11256,N_9981);
and U14924 (N_14924,N_9975,N_12481);
nand U14925 (N_14925,N_11032,N_12289);
nor U14926 (N_14926,N_11065,N_10114);
xor U14927 (N_14927,N_10339,N_9647);
or U14928 (N_14928,N_10184,N_9811);
and U14929 (N_14929,N_10661,N_9435);
or U14930 (N_14930,N_10645,N_9839);
nor U14931 (N_14931,N_10872,N_9562);
nand U14932 (N_14932,N_11095,N_11142);
xnor U14933 (N_14933,N_10882,N_10605);
xor U14934 (N_14934,N_9665,N_9780);
and U14935 (N_14935,N_11031,N_11226);
xor U14936 (N_14936,N_10233,N_9424);
xor U14937 (N_14937,N_12221,N_12148);
xor U14938 (N_14938,N_10796,N_9546);
or U14939 (N_14939,N_10860,N_12075);
nor U14940 (N_14940,N_12065,N_11795);
xor U14941 (N_14941,N_11634,N_10418);
or U14942 (N_14942,N_12394,N_11896);
nor U14943 (N_14943,N_11694,N_11601);
nand U14944 (N_14944,N_10645,N_11432);
or U14945 (N_14945,N_9833,N_10583);
and U14946 (N_14946,N_12363,N_10673);
nand U14947 (N_14947,N_10986,N_10505);
and U14948 (N_14948,N_10426,N_12011);
nor U14949 (N_14949,N_9425,N_9387);
xor U14950 (N_14950,N_10668,N_11641);
xor U14951 (N_14951,N_11571,N_10928);
and U14952 (N_14952,N_11236,N_9549);
or U14953 (N_14953,N_11863,N_11638);
xnor U14954 (N_14954,N_11315,N_9702);
or U14955 (N_14955,N_9519,N_9758);
or U14956 (N_14956,N_12060,N_11905);
nand U14957 (N_14957,N_9864,N_9456);
and U14958 (N_14958,N_12120,N_9668);
xnor U14959 (N_14959,N_10324,N_11101);
xnor U14960 (N_14960,N_11316,N_10123);
or U14961 (N_14961,N_11067,N_11878);
and U14962 (N_14962,N_11956,N_12289);
or U14963 (N_14963,N_10332,N_11416);
xor U14964 (N_14964,N_11306,N_10936);
and U14965 (N_14965,N_9412,N_9394);
or U14966 (N_14966,N_9776,N_10054);
or U14967 (N_14967,N_10488,N_12415);
or U14968 (N_14968,N_9625,N_11414);
and U14969 (N_14969,N_11927,N_11206);
and U14970 (N_14970,N_12106,N_11225);
xor U14971 (N_14971,N_9628,N_11088);
or U14972 (N_14972,N_9897,N_12079);
nor U14973 (N_14973,N_11764,N_11986);
and U14974 (N_14974,N_10222,N_9403);
nand U14975 (N_14975,N_9714,N_12184);
xor U14976 (N_14976,N_12326,N_10952);
xor U14977 (N_14977,N_10305,N_11284);
and U14978 (N_14978,N_11367,N_12255);
nand U14979 (N_14979,N_9478,N_10689);
xnor U14980 (N_14980,N_12396,N_11691);
nor U14981 (N_14981,N_11763,N_12296);
nor U14982 (N_14982,N_10768,N_11215);
nand U14983 (N_14983,N_9456,N_10950);
xor U14984 (N_14984,N_9916,N_11021);
nand U14985 (N_14985,N_11418,N_10023);
xnor U14986 (N_14986,N_12080,N_9685);
xor U14987 (N_14987,N_10121,N_10341);
or U14988 (N_14988,N_9938,N_11858);
nand U14989 (N_14989,N_10844,N_11508);
nor U14990 (N_14990,N_10022,N_9429);
nand U14991 (N_14991,N_11200,N_10535);
nor U14992 (N_14992,N_11329,N_10701);
nor U14993 (N_14993,N_9913,N_10509);
xnor U14994 (N_14994,N_10388,N_9492);
nand U14995 (N_14995,N_9593,N_10606);
nor U14996 (N_14996,N_12418,N_9414);
nand U14997 (N_14997,N_10562,N_10417);
and U14998 (N_14998,N_12185,N_9701);
nor U14999 (N_14999,N_10047,N_9936);
or U15000 (N_15000,N_10279,N_10984);
and U15001 (N_15001,N_9430,N_11488);
or U15002 (N_15002,N_10373,N_12237);
or U15003 (N_15003,N_9837,N_9378);
nor U15004 (N_15004,N_10186,N_10145);
and U15005 (N_15005,N_12126,N_11270);
xnor U15006 (N_15006,N_9924,N_10525);
nand U15007 (N_15007,N_10504,N_9691);
or U15008 (N_15008,N_10984,N_11468);
xor U15009 (N_15009,N_10586,N_10141);
or U15010 (N_15010,N_9939,N_9673);
xnor U15011 (N_15011,N_11378,N_10759);
nor U15012 (N_15012,N_12257,N_11835);
nand U15013 (N_15013,N_11671,N_12227);
nand U15014 (N_15014,N_9708,N_9668);
and U15015 (N_15015,N_11921,N_10535);
and U15016 (N_15016,N_11713,N_11868);
or U15017 (N_15017,N_12373,N_12118);
and U15018 (N_15018,N_11590,N_10025);
nand U15019 (N_15019,N_11402,N_10090);
and U15020 (N_15020,N_9376,N_12197);
nor U15021 (N_15021,N_12197,N_9548);
xor U15022 (N_15022,N_12037,N_10617);
or U15023 (N_15023,N_11621,N_9582);
nand U15024 (N_15024,N_9922,N_11535);
xor U15025 (N_15025,N_10730,N_11687);
and U15026 (N_15026,N_12062,N_12404);
and U15027 (N_15027,N_10805,N_10027);
or U15028 (N_15028,N_10459,N_11838);
or U15029 (N_15029,N_11332,N_10085);
nor U15030 (N_15030,N_11289,N_9584);
and U15031 (N_15031,N_9613,N_11260);
nor U15032 (N_15032,N_12314,N_11754);
or U15033 (N_15033,N_10738,N_12170);
nand U15034 (N_15034,N_10946,N_11965);
xnor U15035 (N_15035,N_9706,N_11511);
nand U15036 (N_15036,N_12284,N_10509);
or U15037 (N_15037,N_9497,N_11171);
xnor U15038 (N_15038,N_10605,N_10617);
and U15039 (N_15039,N_11735,N_10891);
nand U15040 (N_15040,N_9662,N_9992);
xnor U15041 (N_15041,N_10578,N_10003);
and U15042 (N_15042,N_12132,N_9818);
xor U15043 (N_15043,N_11834,N_10384);
xor U15044 (N_15044,N_9503,N_12266);
and U15045 (N_15045,N_9577,N_11500);
and U15046 (N_15046,N_10354,N_11205);
xnor U15047 (N_15047,N_10943,N_10376);
or U15048 (N_15048,N_10287,N_12366);
xor U15049 (N_15049,N_12141,N_11762);
or U15050 (N_15050,N_10598,N_11784);
xor U15051 (N_15051,N_10695,N_11198);
and U15052 (N_15052,N_10304,N_11940);
xnor U15053 (N_15053,N_12161,N_10865);
or U15054 (N_15054,N_12276,N_9703);
and U15055 (N_15055,N_11419,N_9880);
nor U15056 (N_15056,N_10717,N_11080);
or U15057 (N_15057,N_10425,N_9620);
and U15058 (N_15058,N_10806,N_11160);
xnor U15059 (N_15059,N_11856,N_10102);
and U15060 (N_15060,N_11410,N_10571);
and U15061 (N_15061,N_10636,N_10198);
xor U15062 (N_15062,N_11546,N_11596);
xnor U15063 (N_15063,N_11240,N_12235);
and U15064 (N_15064,N_11054,N_11153);
nor U15065 (N_15065,N_9682,N_11505);
nand U15066 (N_15066,N_10983,N_11406);
nor U15067 (N_15067,N_12134,N_12338);
nand U15068 (N_15068,N_12433,N_12139);
nor U15069 (N_15069,N_12426,N_12234);
nor U15070 (N_15070,N_11500,N_10770);
nand U15071 (N_15071,N_10464,N_10453);
xnor U15072 (N_15072,N_9467,N_12261);
xor U15073 (N_15073,N_10348,N_11032);
nand U15074 (N_15074,N_11892,N_12169);
nand U15075 (N_15075,N_12396,N_9978);
or U15076 (N_15076,N_10109,N_10345);
nand U15077 (N_15077,N_9919,N_10067);
or U15078 (N_15078,N_10233,N_11805);
xor U15079 (N_15079,N_11633,N_11274);
and U15080 (N_15080,N_12182,N_10452);
or U15081 (N_15081,N_10708,N_10690);
nor U15082 (N_15082,N_11746,N_10836);
or U15083 (N_15083,N_11538,N_11146);
nand U15084 (N_15084,N_12293,N_12137);
or U15085 (N_15085,N_9736,N_10451);
nand U15086 (N_15086,N_11012,N_12112);
nor U15087 (N_15087,N_12491,N_12173);
xnor U15088 (N_15088,N_9926,N_10539);
xor U15089 (N_15089,N_10509,N_11490);
or U15090 (N_15090,N_10183,N_10527);
nand U15091 (N_15091,N_10592,N_10641);
or U15092 (N_15092,N_9547,N_11818);
xnor U15093 (N_15093,N_11239,N_10868);
and U15094 (N_15094,N_11693,N_9719);
nand U15095 (N_15095,N_11832,N_9655);
and U15096 (N_15096,N_12460,N_11851);
and U15097 (N_15097,N_11672,N_12034);
nand U15098 (N_15098,N_9420,N_9414);
xor U15099 (N_15099,N_10965,N_9791);
xor U15100 (N_15100,N_12304,N_9568);
and U15101 (N_15101,N_10155,N_12496);
nand U15102 (N_15102,N_10063,N_10761);
and U15103 (N_15103,N_9721,N_10576);
and U15104 (N_15104,N_9423,N_10052);
or U15105 (N_15105,N_9784,N_10348);
or U15106 (N_15106,N_9894,N_10560);
and U15107 (N_15107,N_11091,N_11053);
xnor U15108 (N_15108,N_12274,N_12328);
or U15109 (N_15109,N_10065,N_12258);
or U15110 (N_15110,N_11356,N_11973);
xnor U15111 (N_15111,N_11651,N_11867);
or U15112 (N_15112,N_11088,N_11679);
nor U15113 (N_15113,N_9494,N_12064);
nand U15114 (N_15114,N_11901,N_10676);
nor U15115 (N_15115,N_10431,N_11879);
nand U15116 (N_15116,N_10739,N_10893);
nor U15117 (N_15117,N_9868,N_9468);
xor U15118 (N_15118,N_9896,N_11641);
nand U15119 (N_15119,N_11051,N_9619);
and U15120 (N_15120,N_9627,N_9552);
or U15121 (N_15121,N_11353,N_11961);
xnor U15122 (N_15122,N_11221,N_11628);
nor U15123 (N_15123,N_11703,N_10772);
and U15124 (N_15124,N_10441,N_10762);
nor U15125 (N_15125,N_9753,N_11761);
and U15126 (N_15126,N_11944,N_11063);
or U15127 (N_15127,N_9804,N_10707);
nor U15128 (N_15128,N_11847,N_11282);
and U15129 (N_15129,N_10248,N_10049);
nor U15130 (N_15130,N_10293,N_10539);
nand U15131 (N_15131,N_11436,N_9554);
nor U15132 (N_15132,N_10425,N_10446);
and U15133 (N_15133,N_11709,N_10292);
or U15134 (N_15134,N_10924,N_11591);
and U15135 (N_15135,N_10223,N_12261);
nor U15136 (N_15136,N_10821,N_12492);
and U15137 (N_15137,N_9772,N_10435);
nand U15138 (N_15138,N_10289,N_11721);
xnor U15139 (N_15139,N_10785,N_12370);
or U15140 (N_15140,N_12365,N_9411);
nor U15141 (N_15141,N_11886,N_10100);
and U15142 (N_15142,N_11252,N_10080);
or U15143 (N_15143,N_10498,N_9393);
xor U15144 (N_15144,N_11021,N_11198);
nand U15145 (N_15145,N_11168,N_9819);
and U15146 (N_15146,N_12314,N_9729);
nand U15147 (N_15147,N_11937,N_11405);
nor U15148 (N_15148,N_9419,N_11778);
nand U15149 (N_15149,N_10489,N_12391);
and U15150 (N_15150,N_11112,N_10758);
nor U15151 (N_15151,N_11516,N_11631);
and U15152 (N_15152,N_12258,N_12457);
nand U15153 (N_15153,N_11251,N_11295);
or U15154 (N_15154,N_11709,N_9475);
nor U15155 (N_15155,N_10684,N_10981);
nor U15156 (N_15156,N_10757,N_9779);
and U15157 (N_15157,N_9380,N_10082);
xor U15158 (N_15158,N_9459,N_9719);
nor U15159 (N_15159,N_11186,N_12370);
nor U15160 (N_15160,N_12118,N_11756);
and U15161 (N_15161,N_9816,N_11665);
xnor U15162 (N_15162,N_12358,N_10744);
nand U15163 (N_15163,N_11444,N_11514);
or U15164 (N_15164,N_11889,N_10203);
nor U15165 (N_15165,N_9675,N_10598);
or U15166 (N_15166,N_10337,N_11008);
nand U15167 (N_15167,N_9578,N_9875);
xnor U15168 (N_15168,N_9935,N_11039);
and U15169 (N_15169,N_10958,N_11954);
or U15170 (N_15170,N_12286,N_11113);
xor U15171 (N_15171,N_10387,N_12448);
and U15172 (N_15172,N_11649,N_11394);
nand U15173 (N_15173,N_12157,N_9710);
nand U15174 (N_15174,N_10879,N_11515);
nor U15175 (N_15175,N_11615,N_10837);
xnor U15176 (N_15176,N_10336,N_10352);
xor U15177 (N_15177,N_12267,N_10592);
nor U15178 (N_15178,N_10137,N_11568);
nand U15179 (N_15179,N_9463,N_12045);
and U15180 (N_15180,N_10749,N_10522);
nor U15181 (N_15181,N_12468,N_11029);
xor U15182 (N_15182,N_10190,N_10812);
nand U15183 (N_15183,N_12369,N_10389);
and U15184 (N_15184,N_9523,N_9381);
nor U15185 (N_15185,N_12051,N_10973);
xnor U15186 (N_15186,N_11912,N_9967);
xnor U15187 (N_15187,N_10093,N_11184);
and U15188 (N_15188,N_10024,N_12376);
nor U15189 (N_15189,N_10233,N_10886);
nor U15190 (N_15190,N_10024,N_10602);
nand U15191 (N_15191,N_12220,N_11150);
nand U15192 (N_15192,N_12492,N_10943);
xnor U15193 (N_15193,N_10100,N_11616);
and U15194 (N_15194,N_12398,N_10518);
xnor U15195 (N_15195,N_12375,N_10667);
nor U15196 (N_15196,N_11329,N_12463);
nand U15197 (N_15197,N_10663,N_10978);
nand U15198 (N_15198,N_9987,N_10184);
nand U15199 (N_15199,N_10899,N_11300);
nor U15200 (N_15200,N_11057,N_10153);
or U15201 (N_15201,N_10637,N_10556);
nand U15202 (N_15202,N_11394,N_12183);
nand U15203 (N_15203,N_9773,N_10296);
and U15204 (N_15204,N_10936,N_11287);
xor U15205 (N_15205,N_11661,N_11316);
nor U15206 (N_15206,N_12393,N_11937);
and U15207 (N_15207,N_11559,N_12117);
or U15208 (N_15208,N_10585,N_9816);
nor U15209 (N_15209,N_11878,N_10490);
nor U15210 (N_15210,N_11890,N_11377);
nor U15211 (N_15211,N_11780,N_11011);
xnor U15212 (N_15212,N_10473,N_12109);
nand U15213 (N_15213,N_10506,N_11110);
nand U15214 (N_15214,N_12373,N_11441);
nor U15215 (N_15215,N_12489,N_11426);
xnor U15216 (N_15216,N_9993,N_11562);
nand U15217 (N_15217,N_10417,N_10923);
or U15218 (N_15218,N_9693,N_12091);
and U15219 (N_15219,N_11475,N_11820);
xnor U15220 (N_15220,N_12389,N_11216);
or U15221 (N_15221,N_11104,N_9916);
nand U15222 (N_15222,N_11805,N_10999);
xor U15223 (N_15223,N_12403,N_11297);
and U15224 (N_15224,N_10017,N_10405);
nand U15225 (N_15225,N_11758,N_10809);
nand U15226 (N_15226,N_11266,N_10891);
and U15227 (N_15227,N_11034,N_11236);
xor U15228 (N_15228,N_12420,N_12091);
nand U15229 (N_15229,N_12249,N_10949);
nand U15230 (N_15230,N_9433,N_11196);
or U15231 (N_15231,N_11984,N_9955);
and U15232 (N_15232,N_10827,N_10329);
nor U15233 (N_15233,N_11443,N_11073);
nand U15234 (N_15234,N_9658,N_10171);
nand U15235 (N_15235,N_11418,N_11704);
nor U15236 (N_15236,N_11375,N_12321);
or U15237 (N_15237,N_12204,N_9483);
xnor U15238 (N_15238,N_12057,N_10234);
and U15239 (N_15239,N_9489,N_12373);
or U15240 (N_15240,N_12078,N_9933);
nor U15241 (N_15241,N_10421,N_10838);
nor U15242 (N_15242,N_9833,N_10705);
and U15243 (N_15243,N_11495,N_10605);
nand U15244 (N_15244,N_12456,N_9712);
and U15245 (N_15245,N_9721,N_9401);
or U15246 (N_15246,N_10686,N_11527);
nor U15247 (N_15247,N_10971,N_9597);
and U15248 (N_15248,N_11725,N_9773);
and U15249 (N_15249,N_10038,N_11226);
and U15250 (N_15250,N_9659,N_9688);
or U15251 (N_15251,N_10913,N_10205);
or U15252 (N_15252,N_11228,N_9706);
nor U15253 (N_15253,N_12183,N_11914);
or U15254 (N_15254,N_10736,N_11958);
nand U15255 (N_15255,N_10333,N_10873);
nor U15256 (N_15256,N_12394,N_10113);
or U15257 (N_15257,N_9759,N_11770);
and U15258 (N_15258,N_11631,N_11406);
or U15259 (N_15259,N_9829,N_10148);
xor U15260 (N_15260,N_11105,N_12107);
or U15261 (N_15261,N_11844,N_10654);
nor U15262 (N_15262,N_10645,N_10808);
and U15263 (N_15263,N_10678,N_12394);
and U15264 (N_15264,N_10055,N_9991);
nor U15265 (N_15265,N_12488,N_9830);
nand U15266 (N_15266,N_12126,N_11929);
and U15267 (N_15267,N_10616,N_10235);
or U15268 (N_15268,N_11075,N_10057);
and U15269 (N_15269,N_11168,N_10206);
or U15270 (N_15270,N_10237,N_9949);
or U15271 (N_15271,N_10792,N_10264);
or U15272 (N_15272,N_11662,N_11735);
and U15273 (N_15273,N_9477,N_9606);
or U15274 (N_15274,N_9811,N_9538);
xnor U15275 (N_15275,N_10830,N_9485);
and U15276 (N_15276,N_10082,N_11331);
nor U15277 (N_15277,N_11148,N_10345);
or U15278 (N_15278,N_11900,N_12238);
xnor U15279 (N_15279,N_12065,N_9609);
and U15280 (N_15280,N_11214,N_10763);
and U15281 (N_15281,N_10625,N_11335);
or U15282 (N_15282,N_11328,N_11010);
nor U15283 (N_15283,N_10237,N_11230);
xor U15284 (N_15284,N_10113,N_12226);
xnor U15285 (N_15285,N_12038,N_9853);
nor U15286 (N_15286,N_11424,N_11909);
and U15287 (N_15287,N_10964,N_9614);
or U15288 (N_15288,N_9887,N_10759);
and U15289 (N_15289,N_11845,N_10249);
and U15290 (N_15290,N_11020,N_9643);
or U15291 (N_15291,N_12215,N_11168);
or U15292 (N_15292,N_11828,N_10064);
or U15293 (N_15293,N_12000,N_11361);
nor U15294 (N_15294,N_11718,N_12337);
nor U15295 (N_15295,N_12435,N_10235);
and U15296 (N_15296,N_9866,N_11458);
or U15297 (N_15297,N_11049,N_12183);
or U15298 (N_15298,N_12127,N_9868);
xor U15299 (N_15299,N_12070,N_10660);
nand U15300 (N_15300,N_12399,N_11362);
and U15301 (N_15301,N_11181,N_10158);
nand U15302 (N_15302,N_9733,N_11302);
xor U15303 (N_15303,N_10522,N_10191);
nand U15304 (N_15304,N_9440,N_12018);
xnor U15305 (N_15305,N_11870,N_10918);
nand U15306 (N_15306,N_11758,N_10209);
or U15307 (N_15307,N_10454,N_9641);
and U15308 (N_15308,N_12423,N_9751);
nor U15309 (N_15309,N_9853,N_11220);
and U15310 (N_15310,N_11712,N_11905);
nand U15311 (N_15311,N_11670,N_11073);
xnor U15312 (N_15312,N_10590,N_11627);
or U15313 (N_15313,N_10995,N_11710);
nand U15314 (N_15314,N_10658,N_11156);
and U15315 (N_15315,N_11356,N_12275);
nand U15316 (N_15316,N_11427,N_9469);
nor U15317 (N_15317,N_10411,N_11372);
and U15318 (N_15318,N_11849,N_11343);
and U15319 (N_15319,N_10398,N_12330);
xor U15320 (N_15320,N_11111,N_11159);
xnor U15321 (N_15321,N_10050,N_10258);
nor U15322 (N_15322,N_12023,N_10721);
nor U15323 (N_15323,N_11141,N_11644);
or U15324 (N_15324,N_9926,N_9923);
xor U15325 (N_15325,N_11545,N_10052);
xnor U15326 (N_15326,N_11573,N_11958);
or U15327 (N_15327,N_10433,N_12463);
xnor U15328 (N_15328,N_11702,N_12288);
or U15329 (N_15329,N_12213,N_11602);
and U15330 (N_15330,N_11624,N_11864);
nor U15331 (N_15331,N_10205,N_11233);
or U15332 (N_15332,N_12252,N_11516);
xnor U15333 (N_15333,N_11945,N_11855);
and U15334 (N_15334,N_9610,N_12384);
nor U15335 (N_15335,N_11337,N_11705);
nor U15336 (N_15336,N_9499,N_9860);
xnor U15337 (N_15337,N_10760,N_10197);
and U15338 (N_15338,N_12145,N_11081);
xnor U15339 (N_15339,N_10753,N_11541);
xnor U15340 (N_15340,N_11969,N_11458);
xnor U15341 (N_15341,N_11647,N_9964);
nand U15342 (N_15342,N_9676,N_12099);
nor U15343 (N_15343,N_11095,N_11108);
nor U15344 (N_15344,N_10874,N_9517);
and U15345 (N_15345,N_11651,N_10949);
nor U15346 (N_15346,N_10909,N_11366);
or U15347 (N_15347,N_10717,N_9457);
nor U15348 (N_15348,N_11589,N_10203);
xor U15349 (N_15349,N_10744,N_10544);
or U15350 (N_15350,N_11476,N_10995);
or U15351 (N_15351,N_11474,N_10417);
or U15352 (N_15352,N_10108,N_10771);
and U15353 (N_15353,N_12347,N_11502);
xnor U15354 (N_15354,N_11427,N_10905);
nand U15355 (N_15355,N_12467,N_10858);
nand U15356 (N_15356,N_11756,N_10845);
and U15357 (N_15357,N_12469,N_11183);
or U15358 (N_15358,N_11939,N_10272);
xor U15359 (N_15359,N_10307,N_9538);
or U15360 (N_15360,N_9992,N_10028);
or U15361 (N_15361,N_9874,N_10810);
and U15362 (N_15362,N_11493,N_10600);
or U15363 (N_15363,N_11562,N_12321);
xnor U15364 (N_15364,N_10841,N_11047);
and U15365 (N_15365,N_11142,N_11821);
nor U15366 (N_15366,N_12323,N_11914);
nor U15367 (N_15367,N_11055,N_11946);
or U15368 (N_15368,N_12428,N_11616);
or U15369 (N_15369,N_12012,N_12440);
nand U15370 (N_15370,N_11778,N_12014);
nand U15371 (N_15371,N_10860,N_9501);
nand U15372 (N_15372,N_9845,N_12128);
or U15373 (N_15373,N_12219,N_10004);
nor U15374 (N_15374,N_9712,N_10615);
and U15375 (N_15375,N_9693,N_11980);
nor U15376 (N_15376,N_9681,N_11648);
or U15377 (N_15377,N_11972,N_12252);
or U15378 (N_15378,N_10601,N_9603);
nor U15379 (N_15379,N_9505,N_11147);
nand U15380 (N_15380,N_10783,N_12310);
nor U15381 (N_15381,N_10906,N_11911);
and U15382 (N_15382,N_11030,N_11867);
or U15383 (N_15383,N_12461,N_9928);
nand U15384 (N_15384,N_11228,N_9895);
and U15385 (N_15385,N_12425,N_10035);
nand U15386 (N_15386,N_12251,N_11524);
or U15387 (N_15387,N_11788,N_9601);
nand U15388 (N_15388,N_11587,N_12440);
nor U15389 (N_15389,N_11988,N_9757);
xnor U15390 (N_15390,N_11087,N_10484);
xor U15391 (N_15391,N_12249,N_9943);
or U15392 (N_15392,N_10433,N_11653);
nand U15393 (N_15393,N_11041,N_12371);
nor U15394 (N_15394,N_11777,N_12300);
or U15395 (N_15395,N_10461,N_11211);
and U15396 (N_15396,N_12058,N_10670);
xor U15397 (N_15397,N_12479,N_9935);
nor U15398 (N_15398,N_11721,N_11356);
and U15399 (N_15399,N_10658,N_11265);
xor U15400 (N_15400,N_12001,N_11260);
nand U15401 (N_15401,N_11431,N_9940);
and U15402 (N_15402,N_9378,N_12109);
nor U15403 (N_15403,N_9994,N_11112);
xnor U15404 (N_15404,N_9376,N_11255);
xnor U15405 (N_15405,N_10732,N_11177);
nand U15406 (N_15406,N_11419,N_10159);
and U15407 (N_15407,N_9966,N_12275);
nor U15408 (N_15408,N_9745,N_12262);
nor U15409 (N_15409,N_11806,N_10503);
or U15410 (N_15410,N_10747,N_9465);
nand U15411 (N_15411,N_10401,N_10037);
xnor U15412 (N_15412,N_9701,N_10391);
xnor U15413 (N_15413,N_11163,N_12240);
or U15414 (N_15414,N_10252,N_10613);
and U15415 (N_15415,N_11789,N_9419);
nor U15416 (N_15416,N_11194,N_12101);
and U15417 (N_15417,N_9998,N_10376);
and U15418 (N_15418,N_11482,N_9896);
xnor U15419 (N_15419,N_10182,N_11189);
xnor U15420 (N_15420,N_9822,N_9478);
or U15421 (N_15421,N_10357,N_9617);
xnor U15422 (N_15422,N_10683,N_11695);
nand U15423 (N_15423,N_10363,N_10661);
and U15424 (N_15424,N_11608,N_11503);
xnor U15425 (N_15425,N_11935,N_12096);
nand U15426 (N_15426,N_11498,N_11638);
and U15427 (N_15427,N_11785,N_10904);
nor U15428 (N_15428,N_10627,N_11342);
nor U15429 (N_15429,N_10898,N_10956);
or U15430 (N_15430,N_10860,N_12315);
xnor U15431 (N_15431,N_10204,N_12243);
nor U15432 (N_15432,N_9766,N_10512);
or U15433 (N_15433,N_10567,N_9519);
and U15434 (N_15434,N_11796,N_11577);
nor U15435 (N_15435,N_11418,N_9375);
nor U15436 (N_15436,N_11461,N_11930);
xnor U15437 (N_15437,N_10342,N_10801);
xor U15438 (N_15438,N_11478,N_9416);
nor U15439 (N_15439,N_11849,N_12153);
nor U15440 (N_15440,N_11365,N_12130);
nand U15441 (N_15441,N_11099,N_10572);
or U15442 (N_15442,N_11569,N_11268);
or U15443 (N_15443,N_10541,N_9495);
xnor U15444 (N_15444,N_12007,N_11392);
xnor U15445 (N_15445,N_9534,N_10222);
xnor U15446 (N_15446,N_9978,N_11666);
nor U15447 (N_15447,N_10964,N_10435);
and U15448 (N_15448,N_11629,N_12351);
nor U15449 (N_15449,N_12091,N_10687);
nor U15450 (N_15450,N_10749,N_11837);
or U15451 (N_15451,N_9943,N_10225);
nor U15452 (N_15452,N_10169,N_12296);
nor U15453 (N_15453,N_12168,N_9600);
nand U15454 (N_15454,N_10600,N_10422);
or U15455 (N_15455,N_12317,N_11943);
and U15456 (N_15456,N_10937,N_11963);
nor U15457 (N_15457,N_10878,N_10351);
xnor U15458 (N_15458,N_11975,N_9806);
nor U15459 (N_15459,N_10156,N_12223);
or U15460 (N_15460,N_9438,N_9708);
or U15461 (N_15461,N_11949,N_10981);
nand U15462 (N_15462,N_10402,N_9959);
or U15463 (N_15463,N_12241,N_10280);
nand U15464 (N_15464,N_11933,N_12378);
or U15465 (N_15465,N_10293,N_11047);
and U15466 (N_15466,N_10421,N_10728);
and U15467 (N_15467,N_9421,N_9390);
nor U15468 (N_15468,N_10281,N_10247);
nor U15469 (N_15469,N_10547,N_10767);
or U15470 (N_15470,N_10289,N_10279);
nand U15471 (N_15471,N_11772,N_9698);
nand U15472 (N_15472,N_12296,N_12146);
nor U15473 (N_15473,N_12447,N_10404);
nand U15474 (N_15474,N_11671,N_9995);
nor U15475 (N_15475,N_10425,N_11770);
or U15476 (N_15476,N_11421,N_11819);
or U15477 (N_15477,N_10176,N_12446);
nand U15478 (N_15478,N_10544,N_9562);
xnor U15479 (N_15479,N_11788,N_10928);
and U15480 (N_15480,N_12363,N_9610);
xnor U15481 (N_15481,N_10579,N_9804);
nor U15482 (N_15482,N_9650,N_9912);
and U15483 (N_15483,N_10118,N_10536);
xor U15484 (N_15484,N_12318,N_10357);
xor U15485 (N_15485,N_9992,N_10972);
or U15486 (N_15486,N_10456,N_11049);
xor U15487 (N_15487,N_12110,N_10526);
nor U15488 (N_15488,N_10299,N_9709);
nand U15489 (N_15489,N_10625,N_9632);
and U15490 (N_15490,N_12040,N_11712);
nor U15491 (N_15491,N_10499,N_12380);
nand U15492 (N_15492,N_10926,N_10232);
xnor U15493 (N_15493,N_11598,N_11977);
or U15494 (N_15494,N_9846,N_9927);
xnor U15495 (N_15495,N_12168,N_11766);
and U15496 (N_15496,N_9773,N_12155);
xor U15497 (N_15497,N_10721,N_9748);
or U15498 (N_15498,N_10523,N_9917);
or U15499 (N_15499,N_10184,N_11679);
xnor U15500 (N_15500,N_10627,N_11372);
and U15501 (N_15501,N_10847,N_10111);
nor U15502 (N_15502,N_10545,N_11204);
or U15503 (N_15503,N_11336,N_10307);
nand U15504 (N_15504,N_11771,N_10074);
xnor U15505 (N_15505,N_10466,N_9940);
or U15506 (N_15506,N_9822,N_12118);
nand U15507 (N_15507,N_12243,N_11575);
nand U15508 (N_15508,N_9992,N_12218);
or U15509 (N_15509,N_12392,N_11751);
or U15510 (N_15510,N_12034,N_11360);
nor U15511 (N_15511,N_9911,N_10545);
nand U15512 (N_15512,N_11025,N_10648);
nor U15513 (N_15513,N_10190,N_11779);
xnor U15514 (N_15514,N_10645,N_10011);
xnor U15515 (N_15515,N_10243,N_10587);
and U15516 (N_15516,N_10571,N_12023);
and U15517 (N_15517,N_11162,N_12236);
xor U15518 (N_15518,N_10640,N_11226);
or U15519 (N_15519,N_12241,N_11471);
and U15520 (N_15520,N_11193,N_10594);
nor U15521 (N_15521,N_9447,N_11578);
or U15522 (N_15522,N_10207,N_11631);
nand U15523 (N_15523,N_11602,N_11366);
and U15524 (N_15524,N_9959,N_10540);
xor U15525 (N_15525,N_11782,N_11930);
and U15526 (N_15526,N_10687,N_10038);
xnor U15527 (N_15527,N_9847,N_11320);
and U15528 (N_15528,N_10825,N_10379);
xnor U15529 (N_15529,N_11171,N_10962);
and U15530 (N_15530,N_12064,N_11351);
nand U15531 (N_15531,N_12140,N_11299);
nor U15532 (N_15532,N_9715,N_11187);
or U15533 (N_15533,N_11613,N_10734);
or U15534 (N_15534,N_11646,N_10903);
nand U15535 (N_15535,N_9561,N_11351);
nand U15536 (N_15536,N_11273,N_10490);
xor U15537 (N_15537,N_11202,N_11764);
or U15538 (N_15538,N_10214,N_10684);
nor U15539 (N_15539,N_10427,N_9986);
nand U15540 (N_15540,N_9672,N_10343);
nor U15541 (N_15541,N_10517,N_10463);
and U15542 (N_15542,N_10012,N_11671);
nand U15543 (N_15543,N_11373,N_9840);
nor U15544 (N_15544,N_12231,N_11495);
and U15545 (N_15545,N_11476,N_11463);
and U15546 (N_15546,N_11016,N_11005);
xor U15547 (N_15547,N_10671,N_11693);
or U15548 (N_15548,N_10982,N_11565);
nor U15549 (N_15549,N_12407,N_12194);
or U15550 (N_15550,N_10841,N_12194);
and U15551 (N_15551,N_9641,N_11997);
xnor U15552 (N_15552,N_9726,N_10808);
xnor U15553 (N_15553,N_11077,N_10112);
nor U15554 (N_15554,N_10349,N_12406);
nand U15555 (N_15555,N_12219,N_9716);
nand U15556 (N_15556,N_11138,N_10641);
nor U15557 (N_15557,N_9618,N_11015);
nand U15558 (N_15558,N_10961,N_11510);
or U15559 (N_15559,N_10002,N_11015);
and U15560 (N_15560,N_12075,N_11910);
nand U15561 (N_15561,N_12293,N_10104);
nor U15562 (N_15562,N_11185,N_12354);
nand U15563 (N_15563,N_12210,N_11334);
or U15564 (N_15564,N_11398,N_9390);
and U15565 (N_15565,N_11136,N_11080);
nand U15566 (N_15566,N_12019,N_10542);
nor U15567 (N_15567,N_11429,N_9526);
xor U15568 (N_15568,N_9631,N_10968);
xnor U15569 (N_15569,N_11347,N_10459);
nand U15570 (N_15570,N_9458,N_11114);
nand U15571 (N_15571,N_11471,N_11224);
and U15572 (N_15572,N_11617,N_10191);
and U15573 (N_15573,N_10446,N_11500);
and U15574 (N_15574,N_9888,N_11895);
or U15575 (N_15575,N_9665,N_10508);
or U15576 (N_15576,N_10125,N_9469);
or U15577 (N_15577,N_9602,N_9846);
nand U15578 (N_15578,N_11330,N_10373);
and U15579 (N_15579,N_11201,N_11933);
nor U15580 (N_15580,N_11175,N_9536);
or U15581 (N_15581,N_12126,N_11691);
and U15582 (N_15582,N_9857,N_9895);
nand U15583 (N_15583,N_11742,N_12098);
nand U15584 (N_15584,N_11476,N_11157);
nand U15585 (N_15585,N_11608,N_11378);
xnor U15586 (N_15586,N_9731,N_9601);
nor U15587 (N_15587,N_12285,N_11849);
nor U15588 (N_15588,N_11048,N_10567);
nor U15589 (N_15589,N_10489,N_10294);
nand U15590 (N_15590,N_10073,N_11770);
and U15591 (N_15591,N_9902,N_9832);
xor U15592 (N_15592,N_11884,N_9919);
or U15593 (N_15593,N_10199,N_11918);
nand U15594 (N_15594,N_11233,N_12028);
nor U15595 (N_15595,N_11308,N_10085);
xnor U15596 (N_15596,N_10145,N_11029);
nor U15597 (N_15597,N_12049,N_10384);
nand U15598 (N_15598,N_10730,N_10400);
nor U15599 (N_15599,N_9662,N_10267);
or U15600 (N_15600,N_10239,N_10589);
xor U15601 (N_15601,N_11227,N_11644);
nand U15602 (N_15602,N_10404,N_11194);
or U15603 (N_15603,N_12234,N_10459);
and U15604 (N_15604,N_10377,N_9892);
nand U15605 (N_15605,N_9765,N_11358);
nand U15606 (N_15606,N_9722,N_12303);
nand U15607 (N_15607,N_11405,N_9626);
nand U15608 (N_15608,N_10662,N_12336);
and U15609 (N_15609,N_12088,N_11779);
and U15610 (N_15610,N_10305,N_10168);
nand U15611 (N_15611,N_9602,N_10364);
xnor U15612 (N_15612,N_12099,N_12334);
and U15613 (N_15613,N_11030,N_9669);
nor U15614 (N_15614,N_11498,N_11476);
nand U15615 (N_15615,N_9581,N_10411);
or U15616 (N_15616,N_9460,N_11137);
and U15617 (N_15617,N_9581,N_10087);
and U15618 (N_15618,N_11444,N_9780);
xnor U15619 (N_15619,N_9520,N_9721);
nor U15620 (N_15620,N_10986,N_11355);
nor U15621 (N_15621,N_10092,N_10433);
nor U15622 (N_15622,N_12163,N_10919);
nand U15623 (N_15623,N_10478,N_12301);
nand U15624 (N_15624,N_9432,N_11993);
nor U15625 (N_15625,N_13240,N_15311);
nand U15626 (N_15626,N_14436,N_14340);
and U15627 (N_15627,N_14180,N_12768);
xnor U15628 (N_15628,N_12608,N_15039);
nand U15629 (N_15629,N_13294,N_14251);
nand U15630 (N_15630,N_14461,N_13287);
or U15631 (N_15631,N_13266,N_15451);
xnor U15632 (N_15632,N_13536,N_12852);
nand U15633 (N_15633,N_13637,N_15009);
and U15634 (N_15634,N_12509,N_13223);
nand U15635 (N_15635,N_14162,N_15493);
and U15636 (N_15636,N_13473,N_12804);
nor U15637 (N_15637,N_15334,N_13032);
nand U15638 (N_15638,N_12823,N_15436);
xor U15639 (N_15639,N_13366,N_12859);
and U15640 (N_15640,N_15526,N_13910);
or U15641 (N_15641,N_13087,N_12692);
or U15642 (N_15642,N_14151,N_14469);
or U15643 (N_15643,N_13876,N_14752);
xor U15644 (N_15644,N_12862,N_15123);
xnor U15645 (N_15645,N_13355,N_14944);
nor U15646 (N_15646,N_13357,N_14870);
or U15647 (N_15647,N_14607,N_13128);
or U15648 (N_15648,N_14428,N_14226);
nor U15649 (N_15649,N_15180,N_15139);
nor U15650 (N_15650,N_15549,N_15126);
and U15651 (N_15651,N_13220,N_14505);
nor U15652 (N_15652,N_14680,N_14143);
nand U15653 (N_15653,N_14099,N_12764);
and U15654 (N_15654,N_12558,N_12906);
and U15655 (N_15655,N_14523,N_15524);
and U15656 (N_15656,N_14253,N_13392);
nor U15657 (N_15657,N_14715,N_12958);
nor U15658 (N_15658,N_14077,N_15019);
nor U15659 (N_15659,N_12663,N_12886);
nor U15660 (N_15660,N_12996,N_14093);
nor U15661 (N_15661,N_12536,N_14332);
or U15662 (N_15662,N_13347,N_13216);
nor U15663 (N_15663,N_13629,N_13335);
or U15664 (N_15664,N_14274,N_14916);
nor U15665 (N_15665,N_13088,N_12552);
or U15666 (N_15666,N_12725,N_15392);
xor U15667 (N_15667,N_13172,N_13089);
nor U15668 (N_15668,N_15067,N_12907);
nand U15669 (N_15669,N_15597,N_13821);
nor U15670 (N_15670,N_14361,N_15568);
xor U15671 (N_15671,N_15514,N_13655);
xor U15672 (N_15672,N_13874,N_12734);
xnor U15673 (N_15673,N_14412,N_14603);
nand U15674 (N_15674,N_13479,N_12526);
and U15675 (N_15675,N_13160,N_14167);
and U15676 (N_15676,N_13635,N_12518);
xnor U15677 (N_15677,N_13367,N_13183);
nand U15678 (N_15678,N_13095,N_14137);
nor U15679 (N_15679,N_13455,N_13959);
nor U15680 (N_15680,N_13945,N_14216);
and U15681 (N_15681,N_14262,N_15248);
nand U15682 (N_15682,N_13498,N_15192);
and U15683 (N_15683,N_12601,N_12675);
xor U15684 (N_15684,N_15048,N_15441);
nor U15685 (N_15685,N_15577,N_13836);
xnor U15686 (N_15686,N_12635,N_15435);
xnor U15687 (N_15687,N_13072,N_15558);
nor U15688 (N_15688,N_14693,N_13570);
and U15689 (N_15689,N_13450,N_12869);
and U15690 (N_15690,N_12850,N_12715);
and U15691 (N_15691,N_14481,N_14401);
or U15692 (N_15692,N_15381,N_14853);
and U15693 (N_15693,N_14073,N_13299);
xnor U15694 (N_15694,N_13110,N_15464);
nor U15695 (N_15695,N_15165,N_12875);
nand U15696 (N_15696,N_12729,N_15282);
nand U15697 (N_15697,N_14341,N_15036);
nand U15698 (N_15698,N_13327,N_15460);
nand U15699 (N_15699,N_14559,N_14733);
nand U15700 (N_15700,N_15251,N_13061);
or U15701 (N_15701,N_14899,N_14169);
xnor U15702 (N_15702,N_15147,N_15382);
nor U15703 (N_15703,N_13151,N_13682);
xor U15704 (N_15704,N_13171,N_13077);
xnor U15705 (N_15705,N_14437,N_13238);
nand U15706 (N_15706,N_13757,N_15100);
nand U15707 (N_15707,N_13296,N_13428);
or U15708 (N_15708,N_13701,N_13002);
nor U15709 (N_15709,N_14528,N_15153);
nand U15710 (N_15710,N_14369,N_13215);
nand U15711 (N_15711,N_14185,N_15604);
nand U15712 (N_15712,N_12830,N_14996);
nand U15713 (N_15713,N_15053,N_15098);
nand U15714 (N_15714,N_14782,N_15058);
and U15715 (N_15715,N_15348,N_14628);
xor U15716 (N_15716,N_14466,N_14681);
and U15717 (N_15717,N_15047,N_14156);
xnor U15718 (N_15718,N_15115,N_14533);
xnor U15719 (N_15719,N_12720,N_14491);
nand U15720 (N_15720,N_12501,N_15567);
and U15721 (N_15721,N_14610,N_12980);
nor U15722 (N_15722,N_13565,N_13272);
nor U15723 (N_15723,N_15322,N_14872);
or U15724 (N_15724,N_14705,N_13532);
nor U15725 (N_15725,N_15371,N_13439);
and U15726 (N_15726,N_14506,N_15317);
nor U15727 (N_15727,N_12796,N_13583);
or U15728 (N_15728,N_13548,N_13678);
nand U15729 (N_15729,N_14336,N_15209);
xnor U15730 (N_15730,N_15160,N_15233);
nand U15731 (N_15731,N_13092,N_15150);
nand U15732 (N_15732,N_12941,N_14471);
or U15733 (N_15733,N_14653,N_15375);
nand U15734 (N_15734,N_13751,N_14558);
nor U15735 (N_15735,N_15571,N_13178);
or U15736 (N_15736,N_14738,N_15280);
nand U15737 (N_15737,N_12808,N_13680);
xnor U15738 (N_15738,N_13610,N_14214);
nor U15739 (N_15739,N_15134,N_13530);
nand U15740 (N_15740,N_14120,N_15120);
or U15741 (N_15741,N_14416,N_13199);
nand U15742 (N_15742,N_13600,N_12506);
nor U15743 (N_15743,N_13879,N_15104);
or U15744 (N_15744,N_14240,N_15481);
nand U15745 (N_15745,N_15175,N_14703);
xor U15746 (N_15746,N_13053,N_13919);
nor U15747 (N_15747,N_14021,N_14764);
xor U15748 (N_15748,N_12668,N_12638);
nor U15749 (N_15749,N_15356,N_13803);
and U15750 (N_15750,N_13903,N_12508);
nor U15751 (N_15751,N_13139,N_13405);
nor U15752 (N_15752,N_15228,N_14816);
and U15753 (N_15753,N_14885,N_14871);
nor U15754 (N_15754,N_12927,N_14513);
nand U15755 (N_15755,N_12545,N_13854);
nand U15756 (N_15756,N_13957,N_13711);
nor U15757 (N_15757,N_15310,N_14792);
xnor U15758 (N_15758,N_13982,N_13958);
or U15759 (N_15759,N_15543,N_13603);
nand U15760 (N_15760,N_13602,N_13323);
or U15761 (N_15761,N_14883,N_12737);
or U15762 (N_15762,N_14668,N_14258);
nor U15763 (N_15763,N_14699,N_13971);
nor U15764 (N_15764,N_15199,N_12695);
nor U15765 (N_15765,N_15091,N_15454);
nor U15766 (N_15766,N_12595,N_14904);
nand U15767 (N_15767,N_14122,N_14183);
or U15768 (N_15768,N_15601,N_15389);
xor U15769 (N_15769,N_13650,N_14585);
nand U15770 (N_15770,N_15620,N_12593);
xor U15771 (N_15771,N_14299,N_14330);
and U15772 (N_15772,N_13589,N_14464);
nor U15773 (N_15773,N_15584,N_13411);
nand U15774 (N_15774,N_14874,N_12763);
nor U15775 (N_15775,N_13358,N_12870);
nor U15776 (N_15776,N_13098,N_13121);
xor U15777 (N_15777,N_14431,N_14514);
and U15778 (N_15778,N_15480,N_13349);
xnor U15779 (N_15779,N_12904,N_14832);
nor U15780 (N_15780,N_14370,N_13809);
nor U15781 (N_15781,N_12562,N_14589);
or U15782 (N_15782,N_14114,N_15602);
and U15783 (N_15783,N_15502,N_14422);
nor U15784 (N_15784,N_13526,N_13912);
nand U15785 (N_15785,N_13624,N_13227);
or U15786 (N_15786,N_14754,N_13188);
and U15787 (N_15787,N_15574,N_13560);
xnor U15788 (N_15788,N_13625,N_15443);
nand U15789 (N_15789,N_14671,N_14468);
nand U15790 (N_15790,N_13567,N_13927);
and U15791 (N_15791,N_12930,N_14810);
or U15792 (N_15792,N_15598,N_12643);
nor U15793 (N_15793,N_15097,N_14696);
nor U15794 (N_15794,N_13279,N_14873);
nor U15795 (N_15795,N_12868,N_12682);
xnor U15796 (N_15796,N_13606,N_13553);
and U15797 (N_15797,N_14684,N_15548);
xor U15798 (N_15798,N_13662,N_13165);
nor U15799 (N_15799,N_15294,N_15390);
nor U15800 (N_15800,N_13307,N_14493);
and U15801 (N_15801,N_14002,N_15327);
xnor U15802 (N_15802,N_15466,N_12997);
nand U15803 (N_15803,N_13750,N_12833);
xor U15804 (N_15804,N_14269,N_14859);
xor U15805 (N_15805,N_14414,N_12987);
nand U15806 (N_15806,N_13503,N_13547);
xor U15807 (N_15807,N_13343,N_13642);
or U15808 (N_15808,N_14893,N_13324);
nand U15809 (N_15809,N_13396,N_15622);
and U15810 (N_15810,N_13772,N_15238);
xnor U15811 (N_15811,N_13737,N_13952);
xor U15812 (N_15812,N_14560,N_13947);
or U15813 (N_15813,N_13310,N_13442);
nand U15814 (N_15814,N_14868,N_14982);
and U15815 (N_15815,N_14088,N_15021);
nor U15816 (N_15816,N_15397,N_13715);
and U15817 (N_15817,N_13398,N_12664);
xor U15818 (N_15818,N_14391,N_13669);
nor U15819 (N_15819,N_13695,N_13724);
nand U15820 (N_15820,N_15137,N_13923);
nand U15821 (N_15821,N_14435,N_14081);
nor U15822 (N_15822,N_15266,N_13247);
nand U15823 (N_15823,N_13993,N_14990);
and U15824 (N_15824,N_14731,N_15218);
nor U15825 (N_15825,N_15336,N_13723);
nand U15826 (N_15826,N_12564,N_12936);
nand U15827 (N_15827,N_14001,N_13995);
and U15828 (N_15828,N_12848,N_12861);
nor U15829 (N_15829,N_13161,N_14107);
nand U15830 (N_15830,N_13471,N_13382);
or U15831 (N_15831,N_15186,N_13595);
nor U15832 (N_15832,N_13152,N_12991);
xor U15833 (N_15833,N_14935,N_13133);
and U15834 (N_15834,N_12644,N_14504);
nand U15835 (N_15835,N_14835,N_12798);
or U15836 (N_15836,N_14385,N_13623);
xor U15837 (N_15837,N_14182,N_13890);
or U15838 (N_15838,N_13675,N_12618);
or U15839 (N_15839,N_13146,N_14132);
nor U15840 (N_15840,N_14923,N_12757);
or U15841 (N_15841,N_13293,N_12983);
and U15842 (N_15842,N_14376,N_12673);
nand U15843 (N_15843,N_13696,N_13608);
nor U15844 (N_15844,N_15572,N_13925);
and U15845 (N_15845,N_13867,N_12606);
xnor U15846 (N_15846,N_13273,N_13064);
and U15847 (N_15847,N_12575,N_13672);
and U15848 (N_15848,N_13023,N_14521);
nor U15849 (N_15849,N_14882,N_15346);
nand U15850 (N_15850,N_15055,N_14255);
and U15851 (N_15851,N_13155,N_14264);
or U15852 (N_15852,N_13852,N_14356);
nor U15853 (N_15853,N_13420,N_14490);
or U15854 (N_15854,N_13755,N_13265);
nand U15855 (N_15855,N_13045,N_12752);
nor U15856 (N_15856,N_13915,N_14296);
xnor U15857 (N_15857,N_13877,N_13419);
nand U15858 (N_15858,N_12809,N_15338);
xor U15859 (N_15859,N_14069,N_15507);
nor U15860 (N_15860,N_13404,N_14321);
and U15861 (N_15861,N_12879,N_13738);
or U15862 (N_15862,N_15286,N_13244);
nor U15863 (N_15863,N_13260,N_15398);
or U15864 (N_15864,N_15035,N_15262);
or U15865 (N_15865,N_14282,N_14305);
or U15866 (N_15866,N_14193,N_14146);
xor U15867 (N_15867,N_14095,N_13488);
nor U15868 (N_15868,N_14273,N_15223);
xor U15869 (N_15869,N_14345,N_13054);
and U15870 (N_15870,N_14819,N_12747);
nor U15871 (N_15871,N_15118,N_14366);
and U15872 (N_15872,N_13459,N_15079);
or U15873 (N_15873,N_13861,N_13869);
xnor U15874 (N_15874,N_15086,N_13898);
xnor U15875 (N_15875,N_14420,N_13660);
nand U15876 (N_15876,N_14903,N_14569);
nor U15877 (N_15877,N_14492,N_14993);
nand U15878 (N_15878,N_13164,N_15345);
nand U15879 (N_15879,N_14475,N_12527);
xor U15880 (N_15880,N_14943,N_14244);
or U15881 (N_15881,N_14054,N_12831);
xor U15882 (N_15882,N_15203,N_15422);
and U15883 (N_15883,N_12903,N_15065);
xor U15884 (N_15884,N_13802,N_13326);
nor U15885 (N_15885,N_13081,N_14338);
or U15886 (N_15886,N_13305,N_13531);
nor U15887 (N_15887,N_12700,N_15561);
nand U15888 (N_15888,N_13856,N_13012);
nor U15889 (N_15889,N_14160,N_14259);
nand U15890 (N_15890,N_14925,N_12957);
nand U15891 (N_15891,N_13955,N_13557);
and U15892 (N_15892,N_13538,N_12874);
and U15893 (N_15893,N_12580,N_12774);
nor U15894 (N_15894,N_13581,N_12567);
nand U15895 (N_15895,N_13502,N_13946);
and U15896 (N_15896,N_14398,N_14236);
nor U15897 (N_15897,N_13934,N_13686);
nor U15898 (N_15898,N_14458,N_14836);
nor U15899 (N_15899,N_13786,N_14148);
xor U15900 (N_15900,N_13849,N_13517);
nor U15901 (N_15901,N_13494,N_15029);
xor U15902 (N_15902,N_13550,N_13831);
or U15903 (N_15903,N_13074,N_12802);
and U15904 (N_15904,N_12588,N_13933);
or U15905 (N_15905,N_13440,N_13897);
nor U15906 (N_15906,N_12662,N_13016);
xnor U15907 (N_15907,N_14248,N_14115);
xor U15908 (N_15908,N_12970,N_13566);
nor U15909 (N_15909,N_14322,N_15075);
or U15910 (N_15910,N_14119,N_15552);
nor U15911 (N_15911,N_14657,N_14427);
and U15912 (N_15912,N_13813,N_13791);
nand U15913 (N_15913,N_13492,N_12557);
nand U15914 (N_15914,N_13328,N_13424);
xnor U15915 (N_15915,N_14445,N_14987);
xnor U15916 (N_15916,N_13372,N_12748);
or U15917 (N_15917,N_12612,N_14415);
xor U15918 (N_15918,N_12728,N_12994);
xor U15919 (N_15919,N_13163,N_13951);
or U15920 (N_15920,N_15257,N_12919);
and U15921 (N_15921,N_12532,N_14622);
nand U15922 (N_15922,N_13969,N_13776);
nand U15923 (N_15923,N_13881,N_12780);
or U15924 (N_15924,N_13114,N_14199);
nor U15925 (N_15925,N_14512,N_15504);
xor U15926 (N_15926,N_13425,N_13830);
nand U15927 (N_15927,N_15313,N_14822);
nand U15928 (N_15928,N_12926,N_13014);
nor U15929 (N_15929,N_15285,N_15341);
nor U15930 (N_15930,N_15372,N_13515);
or U15931 (N_15931,N_14865,N_13697);
xnor U15932 (N_15932,N_14438,N_13872);
nand U15933 (N_15933,N_14914,N_12587);
nand U15934 (N_15934,N_12961,N_15073);
nand U15935 (N_15935,N_13040,N_14683);
or U15936 (N_15936,N_14735,N_13871);
nand U15937 (N_15937,N_14544,N_13137);
nand U15938 (N_15938,N_13362,N_13730);
or U15939 (N_15939,N_12585,N_13069);
and U15940 (N_15940,N_12594,N_12538);
xor U15941 (N_15941,N_14397,N_13798);
and U15942 (N_15942,N_12947,N_15049);
nor U15943 (N_15943,N_13278,N_13036);
or U15944 (N_15944,N_15162,N_14465);
nand U15945 (N_15945,N_14746,N_15467);
and U15946 (N_15946,N_14063,N_13640);
nand U15947 (N_15947,N_12990,N_15252);
or U15948 (N_15948,N_15246,N_14474);
nor U15949 (N_15949,N_15169,N_13679);
and U15950 (N_15950,N_13834,N_13099);
or U15951 (N_15951,N_13983,N_14106);
and U15952 (N_15952,N_13926,N_14888);
or U15953 (N_15953,N_13806,N_12547);
nor U15954 (N_15954,N_13722,N_13844);
or U15955 (N_15955,N_13559,N_14172);
nor U15956 (N_15956,N_12881,N_14830);
xnor U15957 (N_15957,N_13415,N_14526);
xor U15958 (N_15958,N_15066,N_14334);
nor U15959 (N_15959,N_13017,N_13258);
nand U15960 (N_15960,N_12882,N_13692);
nor U15961 (N_15961,N_14967,N_15156);
nand U15962 (N_15962,N_14019,N_15510);
nor U15963 (N_15963,N_15155,N_15061);
nand U15964 (N_15964,N_12989,N_14880);
or U15965 (N_15965,N_14869,N_12952);
nand U15966 (N_15966,N_15052,N_15581);
xor U15967 (N_15967,N_15438,N_14165);
and U15968 (N_15968,N_13618,N_12723);
nand U15969 (N_15969,N_14405,N_13713);
xnor U15970 (N_15970,N_13201,N_13304);
xor U15971 (N_15971,N_13921,N_15092);
xnor U15972 (N_15972,N_15088,N_14787);
nand U15973 (N_15973,N_14252,N_15391);
nand U15974 (N_15974,N_12837,N_15269);
nand U15975 (N_15975,N_15471,N_12620);
nand U15976 (N_15976,N_14745,N_13239);
xor U15977 (N_15977,N_15437,N_14234);
nor U15978 (N_15978,N_13233,N_13541);
and U15979 (N_15979,N_13820,N_14009);
nand U15980 (N_15980,N_14265,N_15378);
or U15981 (N_15981,N_12738,N_15108);
nand U15982 (N_15982,N_14110,N_14423);
nand U15983 (N_15983,N_15613,N_14737);
and U15984 (N_15984,N_15012,N_13794);
nand U15985 (N_15985,N_15332,N_12627);
nand U15986 (N_15986,N_13699,N_13251);
nand U15987 (N_15987,N_15562,N_14897);
nand U15988 (N_15988,N_14808,N_14333);
nand U15989 (N_15989,N_13298,N_14522);
or U15990 (N_15990,N_13200,N_14613);
or U15991 (N_15991,N_13018,N_13989);
and U15992 (N_15992,N_14968,N_13892);
nor U15993 (N_15993,N_15420,N_13249);
nor U15994 (N_15994,N_13038,N_13523);
and U15995 (N_15995,N_15585,N_15492);
xnor U15996 (N_15996,N_15363,N_14166);
and U15997 (N_15997,N_12818,N_15535);
or U15998 (N_15998,N_13136,N_14302);
and U15999 (N_15999,N_14038,N_12937);
nor U16000 (N_16000,N_12625,N_15407);
or U16001 (N_16001,N_15517,N_13612);
nand U16002 (N_16002,N_13173,N_14157);
and U16003 (N_16003,N_13719,N_13905);
nor U16004 (N_16004,N_14007,N_14128);
nand U16005 (N_16005,N_13482,N_12541);
and U16006 (N_16006,N_14697,N_15284);
nand U16007 (N_16007,N_13150,N_13329);
xnor U16008 (N_16008,N_13426,N_15131);
and U16009 (N_16009,N_13135,N_14767);
or U16010 (N_16010,N_14291,N_14140);
nor U16011 (N_16011,N_14074,N_15330);
xor U16012 (N_16012,N_13748,N_15198);
nand U16013 (N_16013,N_14994,N_12711);
and U16014 (N_16014,N_14663,N_13225);
or U16015 (N_16015,N_14288,N_12807);
or U16016 (N_16016,N_13552,N_14644);
and U16017 (N_16017,N_14202,N_15352);
nor U16018 (N_16018,N_14682,N_12697);
and U16019 (N_16019,N_13192,N_14948);
and U16020 (N_16020,N_13817,N_13862);
xnor U16021 (N_16021,N_15042,N_12836);
xor U16022 (N_16022,N_13256,N_13907);
nand U16023 (N_16023,N_12613,N_12916);
nor U16024 (N_16024,N_14089,N_15401);
xnor U16025 (N_16025,N_15416,N_14351);
xor U16026 (N_16026,N_13558,N_14201);
nor U16027 (N_16027,N_12579,N_13687);
and U16028 (N_16028,N_13102,N_13285);
or U16029 (N_16029,N_12560,N_13937);
or U16030 (N_16030,N_12946,N_15468);
nor U16031 (N_16031,N_13453,N_13149);
nand U16032 (N_16032,N_12857,N_15074);
and U16033 (N_16033,N_14582,N_15367);
or U16034 (N_16034,N_14542,N_13705);
or U16035 (N_16035,N_15290,N_12535);
nor U16036 (N_16036,N_12999,N_12901);
or U16037 (N_16037,N_15094,N_14494);
nand U16038 (N_16038,N_14472,N_15178);
and U16039 (N_16039,N_13850,N_12826);
nor U16040 (N_16040,N_14755,N_15498);
and U16041 (N_16041,N_15054,N_13648);
nand U16042 (N_16042,N_14649,N_15051);
nor U16043 (N_16043,N_13274,N_13100);
nand U16044 (N_16044,N_14821,N_13994);
and U16045 (N_16045,N_14145,N_15528);
nor U16046 (N_16046,N_14860,N_12993);
and U16047 (N_16047,N_12607,N_13563);
nor U16048 (N_16048,N_12691,N_13378);
or U16049 (N_16049,N_12722,N_14344);
nor U16050 (N_16050,N_13785,N_12650);
xnor U16051 (N_16051,N_14463,N_14775);
or U16052 (N_16052,N_15022,N_12679);
nand U16053 (N_16053,N_12979,N_12688);
xor U16054 (N_16054,N_13319,N_15083);
and U16055 (N_16055,N_12972,N_12888);
or U16056 (N_16056,N_15217,N_13351);
and U16057 (N_16057,N_14176,N_13234);
or U16058 (N_16058,N_13902,N_12977);
and U16059 (N_16059,N_14831,N_14802);
nand U16060 (N_16060,N_15606,N_12843);
or U16061 (N_16061,N_13505,N_15619);
nand U16062 (N_16062,N_14005,N_14700);
and U16063 (N_16063,N_15143,N_14555);
nor U16064 (N_16064,N_13497,N_14794);
nor U16065 (N_16065,N_15006,N_13716);
and U16066 (N_16066,N_13524,N_14660);
nor U16067 (N_16067,N_13665,N_14955);
or U16068 (N_16068,N_14643,N_13375);
xor U16069 (N_16069,N_14066,N_14780);
and U16070 (N_16070,N_14197,N_13747);
nand U16071 (N_16071,N_13438,N_13066);
and U16072 (N_16072,N_14355,N_12940);
and U16073 (N_16073,N_12656,N_13315);
or U16074 (N_16074,N_15179,N_14300);
nor U16075 (N_16075,N_14768,N_13511);
and U16076 (N_16076,N_15000,N_14619);
or U16077 (N_16077,N_13858,N_14317);
nand U16078 (N_16078,N_13141,N_14879);
xnor U16079 (N_16079,N_12933,N_14665);
nor U16080 (N_16080,N_15413,N_15130);
or U16081 (N_16081,N_12591,N_15167);
and U16082 (N_16082,N_12925,N_15521);
or U16083 (N_16083,N_14690,N_14055);
nand U16084 (N_16084,N_13142,N_12914);
or U16085 (N_16085,N_14950,N_13300);
or U16086 (N_16086,N_13996,N_14997);
or U16087 (N_16087,N_14803,N_13932);
xor U16088 (N_16088,N_13084,N_12712);
xnor U16089 (N_16089,N_12880,N_15462);
nor U16090 (N_16090,N_14309,N_12521);
xnor U16091 (N_16091,N_13887,N_15423);
nor U16092 (N_16092,N_14630,N_12670);
and U16093 (N_16093,N_12770,N_13714);
xor U16094 (N_16094,N_15089,N_14963);
and U16095 (N_16095,N_14383,N_13041);
and U16096 (N_16096,N_14926,N_14191);
xor U16097 (N_16097,N_13988,N_12948);
xor U16098 (N_16098,N_14206,N_13280);
or U16099 (N_16099,N_15387,N_13050);
and U16100 (N_16100,N_12701,N_15007);
xnor U16101 (N_16101,N_14985,N_13543);
and U16102 (N_16102,N_13709,N_12924);
xnor U16103 (N_16103,N_13773,N_15596);
or U16104 (N_16104,N_13119,N_13853);
and U16105 (N_16105,N_13394,N_14751);
nand U16106 (N_16106,N_15211,N_15184);
or U16107 (N_16107,N_15560,N_15109);
and U16108 (N_16108,N_14090,N_15511);
nand U16109 (N_16109,N_13076,N_14231);
nand U16110 (N_16110,N_15592,N_15541);
nor U16111 (N_16111,N_14912,N_12840);
or U16112 (N_16112,N_14406,N_12865);
nand U16113 (N_16113,N_15101,N_14006);
xnor U16114 (N_16114,N_13539,N_14432);
nor U16115 (N_16115,N_14900,N_15024);
nor U16116 (N_16116,N_15570,N_13732);
nor U16117 (N_16117,N_13734,N_13960);
nand U16118 (N_16118,N_14678,N_13241);
nand U16119 (N_16119,N_14281,N_13109);
nand U16120 (N_16120,N_12913,N_14581);
and U16121 (N_16121,N_15292,N_13638);
nor U16122 (N_16122,N_15177,N_13677);
and U16123 (N_16123,N_14478,N_13667);
xor U16124 (N_16124,N_14761,N_15062);
and U16125 (N_16125,N_13037,N_15273);
xor U16126 (N_16126,N_14278,N_15183);
nor U16127 (N_16127,N_14549,N_15050);
xnor U16128 (N_16128,N_15288,N_13055);
xor U16129 (N_16129,N_13520,N_12740);
and U16130 (N_16130,N_13782,N_13117);
xor U16131 (N_16131,N_13605,N_14824);
or U16132 (N_16132,N_14297,N_14220);
or U16133 (N_16133,N_15573,N_14026);
nand U16134 (N_16134,N_13377,N_15404);
xor U16135 (N_16135,N_13022,N_13138);
xnor U16136 (N_16136,N_14930,N_14348);
and U16137 (N_16137,N_15281,N_12794);
and U16138 (N_16138,N_13804,N_15253);
xnor U16139 (N_16139,N_12769,N_14488);
xnor U16140 (N_16140,N_12703,N_14600);
xor U16141 (N_16141,N_12824,N_15339);
and U16142 (N_16142,N_14655,N_13434);
nand U16143 (N_16143,N_14983,N_14823);
nand U16144 (N_16144,N_15197,N_13389);
nor U16145 (N_16145,N_14147,N_14689);
xnor U16146 (N_16146,N_13829,N_14225);
and U16147 (N_16147,N_14271,N_13093);
nand U16148 (N_16148,N_14187,N_15174);
nor U16149 (N_16149,N_12998,N_13718);
nand U16150 (N_16150,N_15244,N_14543);
and U16151 (N_16151,N_14820,N_14529);
nor U16152 (N_16152,N_13354,N_14459);
or U16153 (N_16153,N_14638,N_15265);
nor U16154 (N_16154,N_14723,N_13407);
nor U16155 (N_16155,N_14434,N_13592);
nor U16156 (N_16156,N_13104,N_12845);
xor U16157 (N_16157,N_13801,N_14130);
nor U16158 (N_16158,N_13421,N_14509);
xor U16159 (N_16159,N_15445,N_13079);
and U16160 (N_16160,N_15431,N_13401);
xnor U16161 (N_16161,N_13468,N_14329);
nand U16162 (N_16162,N_14541,N_13049);
and U16163 (N_16163,N_15354,N_14242);
nand U16164 (N_16164,N_14625,N_13027);
and U16165 (N_16165,N_14211,N_14959);
nand U16166 (N_16166,N_15475,N_12775);
nand U16167 (N_16167,N_15107,N_14457);
or U16168 (N_16168,N_15316,N_15011);
nand U16169 (N_16169,N_13938,N_13762);
nor U16170 (N_16170,N_14477,N_13930);
nand U16171 (N_16171,N_15110,N_12844);
and U16172 (N_16172,N_15342,N_14708);
nand U16173 (N_16173,N_13271,N_15547);
and U16174 (N_16174,N_14346,N_14629);
and U16175 (N_16175,N_13452,N_13057);
xor U16176 (N_16176,N_12639,N_13232);
or U16177 (N_16177,N_13519,N_14992);
and U16178 (N_16178,N_14765,N_12500);
and U16179 (N_16179,N_13540,N_13270);
nand U16180 (N_16180,N_13864,N_14012);
nor U16181 (N_16181,N_13478,N_14098);
and U16182 (N_16182,N_15105,N_13292);
or U16183 (N_16183,N_14070,N_13390);
nand U16184 (N_16184,N_14651,N_12867);
and U16185 (N_16185,N_12791,N_14064);
and U16186 (N_16186,N_15208,N_14917);
xnor U16187 (N_16187,N_14763,N_14396);
nand U16188 (N_16188,N_14343,N_14503);
xnor U16189 (N_16189,N_13613,N_15512);
nand U16190 (N_16190,N_14050,N_15323);
nand U16191 (N_16191,N_14372,N_15433);
xor U16192 (N_16192,N_15427,N_13622);
nor U16193 (N_16193,N_15506,N_13179);
nor U16194 (N_16194,N_14855,N_15497);
nor U16195 (N_16195,N_14190,N_13616);
xnor U16196 (N_16196,N_15081,N_12651);
or U16197 (N_16197,N_12754,N_15461);
or U16198 (N_16198,N_14818,N_14902);
xor U16199 (N_16199,N_13308,N_14325);
nor U16200 (N_16200,N_13676,N_13551);
nor U16201 (N_16201,N_13028,N_12767);
and U16202 (N_16202,N_14777,N_15538);
nand U16203 (N_16203,N_13659,N_13230);
nand U16204 (N_16204,N_14349,N_14142);
or U16205 (N_16205,N_14710,N_15268);
nand U16206 (N_16206,N_14519,N_13763);
nor U16207 (N_16207,N_13105,N_13948);
nand U16208 (N_16208,N_14108,N_15259);
or U16209 (N_16209,N_15523,N_14139);
and U16210 (N_16210,N_15491,N_14284);
nand U16211 (N_16211,N_15070,N_14238);
and U16212 (N_16212,N_13710,N_13620);
xnor U16213 (N_16213,N_14911,N_12687);
nor U16214 (N_16214,N_13198,N_15299);
nor U16215 (N_16215,N_13860,N_12623);
and U16216 (N_16216,N_13735,N_15271);
or U16217 (N_16217,N_14104,N_13997);
or U16218 (N_16218,N_13210,N_15037);
and U16219 (N_16219,N_13739,N_14901);
nor U16220 (N_16220,N_13427,N_15556);
or U16221 (N_16221,N_14170,N_14194);
nor U16222 (N_16222,N_14245,N_14377);
nand U16223 (N_16223,N_13097,N_15458);
xor U16224 (N_16224,N_14267,N_12741);
nand U16225 (N_16225,N_13129,N_13360);
nand U16226 (N_16226,N_13352,N_13704);
xor U16227 (N_16227,N_12749,N_15030);
and U16228 (N_16228,N_13922,N_15364);
or U16229 (N_16229,N_12745,N_14695);
or U16230 (N_16230,N_14327,N_14123);
nand U16231 (N_16231,N_14363,N_14260);
nand U16232 (N_16232,N_14518,N_15242);
nor U16233 (N_16233,N_13970,N_12995);
and U16234 (N_16234,N_14688,N_13597);
nor U16235 (N_16235,N_14056,N_14947);
xor U16236 (N_16236,N_13371,N_12519);
or U16237 (N_16237,N_13369,N_14953);
xnor U16238 (N_16238,N_15149,N_14706);
nand U16239 (N_16239,N_13339,N_12899);
xor U16240 (N_16240,N_12842,N_14045);
nor U16241 (N_16241,N_14717,N_13506);
and U16242 (N_16242,N_13917,N_14482);
nand U16243 (N_16243,N_15428,N_15525);
nand U16244 (N_16244,N_13978,N_14083);
nor U16245 (N_16245,N_14384,N_12694);
nand U16246 (N_16246,N_12801,N_13579);
nand U16247 (N_16247,N_15575,N_12953);
xor U16248 (N_16248,N_14924,N_14894);
or U16249 (N_16249,N_14168,N_12676);
and U16250 (N_16250,N_15148,N_12931);
xnor U16251 (N_16251,N_13387,N_12549);
and U16252 (N_16252,N_12971,N_14375);
or U16253 (N_16253,N_15550,N_12637);
and U16254 (N_16254,N_13961,N_14347);
and U16255 (N_16255,N_12726,N_13340);
and U16256 (N_16256,N_13731,N_15383);
xnor U16257 (N_16257,N_14850,N_15555);
and U16258 (N_16258,N_12928,N_12884);
or U16259 (N_16259,N_14105,N_15368);
nor U16260 (N_16260,N_15059,N_13187);
nor U16261 (N_16261,N_14446,N_13127);
xor U16262 (N_16262,N_15444,N_14112);
nand U16263 (N_16263,N_14283,N_12896);
nand U16264 (N_16264,N_14748,N_12583);
nand U16265 (N_16265,N_12599,N_12950);
or U16266 (N_16266,N_14379,N_14659);
and U16267 (N_16267,N_13703,N_13564);
and U16268 (N_16268,N_12816,N_15261);
nor U16269 (N_16269,N_13003,N_14381);
xor U16270 (N_16270,N_12810,N_12502);
xor U16271 (N_16271,N_13611,N_12572);
and U16272 (N_16272,N_13333,N_13418);
or U16273 (N_16273,N_13359,N_14539);
nor U16274 (N_16274,N_14936,N_15159);
nand U16275 (N_16275,N_13391,N_12640);
nand U16276 (N_16276,N_13626,N_12524);
nor U16277 (N_16277,N_12762,N_13493);
and U16278 (N_16278,N_13627,N_13968);
nor U16279 (N_16279,N_12598,N_15289);
or U16280 (N_16280,N_12709,N_14286);
nor U16281 (N_16281,N_13302,N_14774);
or U16282 (N_16282,N_14250,N_14228);
xor U16283 (N_16283,N_13826,N_15034);
xor U16284 (N_16284,N_14813,N_15539);
nand U16285 (N_16285,N_12847,N_14817);
xnor U16286 (N_16286,N_14421,N_13656);
or U16287 (N_16287,N_13122,N_14602);
nand U16288 (N_16288,N_15388,N_14141);
nor U16289 (N_16289,N_15344,N_14161);
and U16290 (N_16290,N_15005,N_12596);
nand U16291 (N_16291,N_13005,N_13010);
and U16292 (N_16292,N_12902,N_13047);
xor U16293 (N_16293,N_13528,N_13544);
and U16294 (N_16294,N_15172,N_13744);
xnor U16295 (N_16295,N_13966,N_13193);
nand U16296 (N_16296,N_14308,N_15473);
xnor U16297 (N_16297,N_14154,N_13781);
nor U16298 (N_16298,N_13819,N_14030);
or U16299 (N_16299,N_14337,N_14799);
or U16300 (N_16300,N_12864,N_15230);
and U16301 (N_16301,N_14862,N_13474);
nand U16302 (N_16302,N_13261,N_12956);
nand U16303 (N_16303,N_13364,N_15157);
xor U16304 (N_16304,N_13941,N_15519);
nand U16305 (N_16305,N_13694,N_14965);
nand U16306 (N_16306,N_14411,N_14980);
nand U16307 (N_16307,N_13733,N_12590);
and U16308 (N_16308,N_13313,N_14101);
nand U16309 (N_16309,N_12872,N_12716);
nor U16310 (N_16310,N_14712,N_12605);
xnor U16311 (N_16311,N_12539,N_13370);
nand U16312 (N_16312,N_15457,N_12659);
and U16313 (N_16313,N_12514,N_14280);
nor U16314 (N_16314,N_14789,N_13847);
nand U16315 (N_16315,N_12530,N_12788);
or U16316 (N_16316,N_15017,N_14806);
xnor U16317 (N_16317,N_15578,N_14623);
or U16318 (N_16318,N_13126,N_13195);
or U16319 (N_16319,N_13658,N_13030);
and U16320 (N_16320,N_14719,N_14642);
nand U16321 (N_16321,N_15056,N_13025);
nand U16322 (N_16322,N_14951,N_14887);
xnor U16323 (N_16323,N_13476,N_15494);
xnor U16324 (N_16324,N_12654,N_15196);
nor U16325 (N_16325,N_12755,N_12897);
nor U16326 (N_16326,N_12853,N_14766);
or U16327 (N_16327,N_15231,N_13522);
xnor U16328 (N_16328,N_14373,N_15362);
nor U16329 (N_16329,N_13664,N_15430);
nand U16330 (N_16330,N_14744,N_13033);
nor U16331 (N_16331,N_14937,N_15080);
nor U16332 (N_16332,N_13322,N_14540);
nand U16333 (N_16333,N_14232,N_14928);
nand U16334 (N_16334,N_14929,N_12717);
nor U16335 (N_16335,N_14749,N_14266);
nand U16336 (N_16336,N_14626,N_14109);
or U16337 (N_16337,N_14829,N_12976);
nor U16338 (N_16338,N_13228,N_14554);
nor U16339 (N_16339,N_14212,N_12512);
nand U16340 (N_16340,N_13451,N_13683);
nand U16341 (N_16341,N_14358,N_13397);
or U16342 (N_16342,N_12513,N_15483);
xor U16343 (N_16343,N_14072,N_15087);
and U16344 (N_16344,N_14915,N_12706);
and U16345 (N_16345,N_14004,N_14790);
xnor U16346 (N_16346,N_13094,N_14701);
or U16347 (N_16347,N_13756,N_13046);
nor U16348 (N_16348,N_15090,N_13467);
nand U16349 (N_16349,N_15113,N_13555);
nor U16350 (N_16350,N_14218,N_13771);
xnor U16351 (N_16351,N_12647,N_14016);
nor U16352 (N_16352,N_15045,N_14453);
nor U16353 (N_16353,N_13590,N_14740);
or U16354 (N_16354,N_14442,N_13191);
xor U16355 (N_16355,N_15260,N_14235);
xor U16356 (N_16356,N_13031,N_14440);
nand U16357 (N_16357,N_13768,N_13654);
nor U16358 (N_16358,N_14973,N_15095);
nand U16359 (N_16359,N_14840,N_15312);
xnor U16360 (N_16360,N_13931,N_15331);
xnor U16361 (N_16361,N_12878,N_15509);
nand U16362 (N_16362,N_13736,N_14189);
nand U16363 (N_16363,N_14035,N_13209);
or U16364 (N_16364,N_14339,N_15154);
or U16365 (N_16365,N_12672,N_15301);
xor U16366 (N_16366,N_15361,N_14949);
and U16367 (N_16367,N_13885,N_13706);
nor U16368 (N_16368,N_15533,N_15315);
xnor U16369 (N_16369,N_15554,N_13513);
or U16370 (N_16370,N_14648,N_15295);
and U16371 (N_16371,N_15232,N_14667);
and U16372 (N_16372,N_12719,N_15465);
nor U16373 (N_16373,N_15393,N_14076);
xor U16374 (N_16374,N_14174,N_13621);
or U16375 (N_16375,N_14595,N_13604);
nor U16376 (N_16376,N_13928,N_15025);
and U16377 (N_16377,N_14204,N_13486);
nand U16378 (N_16378,N_14094,N_13158);
nor U16379 (N_16379,N_15041,N_13365);
nor U16380 (N_16380,N_12806,N_14946);
and U16381 (N_16381,N_14078,N_15350);
and U16382 (N_16382,N_13015,N_14023);
nand U16383 (N_16383,N_14954,N_13236);
nor U16384 (N_16384,N_13725,N_13649);
nor U16385 (N_16385,N_12820,N_13111);
or U16386 (N_16386,N_12609,N_14295);
nor U16387 (N_16387,N_15116,N_14545);
nor U16388 (N_16388,N_14661,N_12516);
nor U16389 (N_16389,N_14676,N_14410);
xor U16390 (N_16390,N_13634,N_14298);
xor U16391 (N_16391,N_14756,N_14845);
or U16392 (N_16392,N_14223,N_13384);
or U16393 (N_16393,N_13878,N_14747);
nor U16394 (N_16394,N_14425,N_13901);
and U16395 (N_16395,N_14082,N_12893);
nor U16396 (N_16396,N_14633,N_14516);
or U16397 (N_16397,N_15496,N_13698);
xnor U16398 (N_16398,N_13875,N_14075);
nor U16399 (N_16399,N_15040,N_12838);
nor U16400 (N_16400,N_14910,N_12683);
nand U16401 (N_16401,N_12968,N_14807);
and U16402 (N_16402,N_15447,N_15237);
or U16403 (N_16403,N_12511,N_12510);
xor U16404 (N_16404,N_15530,N_12891);
nor U16405 (N_16405,N_13855,N_13759);
or U16406 (N_16406,N_13103,N_13507);
and U16407 (N_16407,N_13108,N_15202);
and U16408 (N_16408,N_14127,N_14979);
nand U16409 (N_16409,N_13742,N_15616);
and U16410 (N_16410,N_15594,N_14520);
or U16411 (N_16411,N_14939,N_12892);
or U16412 (N_16412,N_12667,N_13645);
xnor U16413 (N_16413,N_14586,N_14179);
nor U16414 (N_16414,N_14815,N_12645);
and U16415 (N_16415,N_14085,N_15003);
and U16416 (N_16416,N_13491,N_13500);
xor U16417 (N_16417,N_12610,N_15142);
nor U16418 (N_16418,N_13689,N_15250);
and U16419 (N_16419,N_14694,N_14732);
nor U16420 (N_16420,N_14538,N_13546);
nand U16421 (N_16421,N_12787,N_14590);
nand U16422 (N_16422,N_15185,N_14646);
and U16423 (N_16423,N_13609,N_12621);
xor U16424 (N_16424,N_15599,N_12905);
nand U16425 (N_16425,N_12975,N_13845);
or U16426 (N_16426,N_13311,N_15226);
or U16427 (N_16427,N_13644,N_15329);
and U16428 (N_16428,N_13430,N_12674);
nand U16429 (N_16429,N_13203,N_12805);
xor U16430 (N_16430,N_12566,N_14429);
or U16431 (N_16431,N_13229,N_13116);
or U16432 (N_16432,N_13029,N_13288);
or U16433 (N_16433,N_13818,N_13832);
xor U16434 (N_16434,N_13106,N_13758);
xor U16435 (N_16435,N_14186,N_14966);
and U16436 (N_16436,N_13571,N_15349);
or U16437 (N_16437,N_15279,N_15275);
nand U16438 (N_16438,N_13363,N_13414);
or U16439 (N_16439,N_15181,N_13044);
and U16440 (N_16440,N_15559,N_14713);
and U16441 (N_16441,N_15077,N_13402);
nand U16442 (N_16442,N_14029,N_13042);
nor U16443 (N_16443,N_14441,N_15424);
nand U16444 (N_16444,N_13218,N_14285);
xor U16445 (N_16445,N_15112,N_14584);
xor U16446 (N_16446,N_13935,N_12789);
nand U16447 (N_16447,N_14884,N_13805);
xnor U16448 (N_16448,N_15057,N_14508);
or U16449 (N_16449,N_15546,N_14467);
nand U16450 (N_16450,N_14084,N_13422);
or U16451 (N_16451,N_13019,N_14452);
and U16452 (N_16452,N_14460,N_12887);
nor U16453 (N_16453,N_13828,N_14640);
nor U16454 (N_16454,N_15145,N_13630);
xnor U16455 (N_16455,N_14233,N_12883);
nor U16456 (N_16456,N_12690,N_13460);
and U16457 (N_16457,N_12563,N_14673);
nor U16458 (N_16458,N_14444,N_14033);
xor U16459 (N_16459,N_14593,N_12555);
and U16460 (N_16460,N_13841,N_15453);
xor U16461 (N_16461,N_13035,N_15505);
or U16462 (N_16462,N_12786,N_13674);
or U16463 (N_16463,N_12822,N_14362);
and U16464 (N_16464,N_14858,N_14662);
xor U16465 (N_16465,N_13857,N_13096);
or U16466 (N_16466,N_14149,N_14757);
xor U16467 (N_16467,N_13998,N_13598);
nor U16468 (N_16468,N_13991,N_12939);
nand U16469 (N_16469,N_13518,N_13316);
nand U16470 (N_16470,N_14323,N_15161);
and U16471 (N_16471,N_14866,N_12900);
nor U16472 (N_16472,N_13226,N_12945);
nand U16473 (N_16473,N_12657,N_14413);
or U16474 (N_16474,N_13026,N_13769);
and U16475 (N_16475,N_14318,N_13639);
nand U16476 (N_16476,N_14814,N_15369);
and U16477 (N_16477,N_13577,N_14498);
or U16478 (N_16478,N_14352,N_15256);
nor U16479 (N_16479,N_14580,N_13578);
nand U16480 (N_16480,N_12665,N_14927);
nand U16481 (N_16481,N_13956,N_12921);
and U16482 (N_16482,N_15264,N_13462);
nand U16483 (N_16483,N_13641,N_14117);
nand U16484 (N_16484,N_15173,N_13586);
nand U16485 (N_16485,N_15229,N_12707);
nand U16486 (N_16486,N_14350,N_14677);
xor U16487 (N_16487,N_14795,N_13796);
or U16488 (N_16488,N_14587,N_14881);
or U16489 (N_16489,N_15277,N_13433);
nor U16490 (N_16490,N_12922,N_14922);
nand U16491 (N_16491,N_13174,N_15023);
xor U16492 (N_16492,N_12849,N_12985);
nor U16493 (N_16493,N_13264,N_15365);
xnor U16494 (N_16494,N_14892,N_13588);
nand U16495 (N_16495,N_13653,N_14188);
and U16496 (N_16496,N_14399,N_14312);
nand U16497 (N_16497,N_12832,N_13987);
nor U16498 (N_16498,N_12954,N_12698);
nor U16499 (N_16499,N_13214,N_13317);
xor U16500 (N_16500,N_13000,N_13726);
and U16501 (N_16501,N_14612,N_14360);
nand U16502 (N_16502,N_13062,N_12671);
and U16503 (N_16503,N_14387,N_14184);
nor U16504 (N_16504,N_14502,N_13469);
nor U16505 (N_16505,N_12646,N_12631);
xor U16506 (N_16506,N_15044,N_13545);
xnor U16507 (N_16507,N_13267,N_13204);
or U16508 (N_16508,N_14034,N_12730);
or U16509 (N_16509,N_13435,N_14268);
xor U16510 (N_16510,N_15318,N_13909);
xnor U16511 (N_16511,N_13443,N_12619);
nand U16512 (N_16512,N_14275,N_15501);
nor U16513 (N_16513,N_12705,N_13159);
and U16514 (N_16514,N_12911,N_14511);
nand U16515 (N_16515,N_13259,N_14027);
and U16516 (N_16516,N_14961,N_14058);
and U16517 (N_16517,N_14592,N_15258);
or U16518 (N_16518,N_12568,N_12507);
nor U16519 (N_16519,N_13380,N_12876);
nand U16520 (N_16520,N_15243,N_15333);
nand U16521 (N_16521,N_12617,N_13840);
and U16522 (N_16522,N_12988,N_15588);
nand U16523 (N_16523,N_13123,N_12721);
xor U16524 (N_16524,N_14249,N_13681);
and U16525 (N_16525,N_15611,N_15084);
xnor U16526 (N_16526,N_14786,N_12520);
nor U16527 (N_16527,N_14480,N_12525);
and U16528 (N_16528,N_15300,N_12858);
and U16529 (N_16529,N_13784,N_14772);
nor U16530 (N_16530,N_13269,N_14618);
nor U16531 (N_16531,N_13070,N_15276);
and U16532 (N_16532,N_14224,N_14551);
nor U16533 (N_16533,N_13441,N_13965);
or U16534 (N_16534,N_15583,N_14256);
and U16535 (N_16535,N_14293,N_14159);
nor U16536 (N_16536,N_15415,N_15534);
or U16537 (N_16537,N_15210,N_14886);
and U16538 (N_16538,N_12505,N_14065);
nor U16539 (N_16539,N_15163,N_13889);
nor U16540 (N_16540,N_15018,N_12540);
nand U16541 (N_16541,N_12577,N_13973);
nand U16542 (N_16542,N_12986,N_13208);
or U16543 (N_16543,N_12731,N_12951);
xnor U16544 (N_16544,N_15400,N_13481);
and U16545 (N_16545,N_13975,N_15063);
and U16546 (N_16546,N_14053,N_12632);
and U16547 (N_16547,N_14430,N_14741);
and U16548 (N_16548,N_14135,N_13985);
and U16549 (N_16549,N_13388,N_14730);
nand U16550 (N_16550,N_15412,N_15124);
xnor U16551 (N_16551,N_13529,N_14692);
and U16552 (N_16552,N_12649,N_14958);
nand U16553 (N_16553,N_13342,N_14207);
nor U16554 (N_16554,N_12856,N_15031);
or U16555 (N_16555,N_13963,N_12603);
nand U16556 (N_16556,N_12761,N_14931);
nor U16557 (N_16557,N_12917,N_13284);
nand U16558 (N_16558,N_14111,N_13615);
nand U16559 (N_16559,N_15495,N_13807);
nor U16560 (N_16560,N_15016,N_14454);
or U16561 (N_16561,N_15353,N_14557);
nand U16562 (N_16562,N_15297,N_14403);
xor U16563 (N_16563,N_12959,N_12574);
or U16564 (N_16564,N_14290,N_14530);
and U16565 (N_16565,N_13337,N_12984);
xor U16566 (N_16566,N_14448,N_15376);
nand U16567 (N_16567,N_13134,N_13297);
nor U16568 (N_16568,N_14641,N_12978);
nor U16569 (N_16569,N_14778,N_14604);
and U16570 (N_16570,N_12811,N_14670);
and U16571 (N_16571,N_14277,N_14704);
and U16572 (N_16572,N_13972,N_15489);
and U16573 (N_16573,N_14960,N_13838);
nand U16574 (N_16574,N_14501,N_14153);
xor U16575 (N_16575,N_13839,N_13177);
or U16576 (N_16576,N_12622,N_15610);
or U16577 (N_16577,N_13501,N_13291);
nand U16578 (N_16578,N_15122,N_15617);
xor U16579 (N_16579,N_12553,N_15121);
xor U16580 (N_16580,N_13211,N_13576);
and U16581 (N_16581,N_14289,N_13413);
and U16582 (N_16582,N_14941,N_13976);
nand U16583 (N_16583,N_13717,N_14152);
nor U16584 (N_16584,N_15219,N_12636);
or U16585 (N_16585,N_14686,N_14675);
and U16586 (N_16586,N_12846,N_14013);
and U16587 (N_16587,N_13341,N_14784);
and U16588 (N_16588,N_13569,N_13052);
nor U16589 (N_16589,N_13423,N_13670);
nand U16590 (N_16590,N_13690,N_13512);
nor U16591 (N_16591,N_15324,N_13437);
or U16592 (N_16592,N_15103,N_13812);
and U16593 (N_16593,N_14827,N_12960);
and U16594 (N_16594,N_13913,N_15099);
nor U16595 (N_16595,N_14116,N_14039);
or U16596 (N_16596,N_12890,N_15500);
and U16597 (N_16597,N_14068,N_14402);
or U16598 (N_16598,N_14567,N_12592);
xor U16599 (N_16599,N_14131,N_15221);
nor U16600 (N_16600,N_12611,N_13379);
or U16601 (N_16601,N_12776,N_15520);
and U16602 (N_16602,N_14531,N_14417);
and U16603 (N_16603,N_14890,N_12974);
nand U16604 (N_16604,N_12727,N_14597);
and U16605 (N_16605,N_14957,N_13495);
xnor U16606 (N_16606,N_13509,N_13400);
nor U16607 (N_16607,N_13145,N_13924);
and U16608 (N_16608,N_14096,N_12814);
xnor U16609 (N_16609,N_13685,N_13436);
xor U16610 (N_16610,N_14834,N_15136);
or U16611 (N_16611,N_13953,N_14311);
nand U16612 (N_16612,N_13814,N_13185);
nand U16613 (N_16613,N_14788,N_12578);
and U16614 (N_16614,N_12779,N_15014);
nand U16615 (N_16615,N_14952,N_13811);
nor U16616 (N_16616,N_15605,N_15490);
nand U16617 (N_16617,N_12828,N_13067);
or U16618 (N_16618,N_12732,N_15254);
nand U16619 (N_16619,N_14483,N_12550);
or U16620 (N_16620,N_14462,N_14018);
nor U16621 (N_16621,N_14577,N_12615);
and U16622 (N_16622,N_13950,N_15158);
nand U16623 (N_16623,N_15565,N_13219);
and U16624 (N_16624,N_12724,N_14192);
and U16625 (N_16625,N_12771,N_12969);
nand U16626 (N_16626,N_14315,N_12797);
and U16627 (N_16627,N_13180,N_15170);
nor U16628 (N_16628,N_13873,N_12582);
and U16629 (N_16629,N_15117,N_13535);
xor U16630 (N_16630,N_15522,N_13120);
nand U16631 (N_16631,N_14791,N_15564);
and U16632 (N_16632,N_15249,N_14227);
and U16633 (N_16633,N_15456,N_14877);
and U16634 (N_16634,N_13870,N_13345);
nand U16635 (N_16635,N_14669,N_14596);
xor U16636 (N_16636,N_14553,N_13661);
or U16637 (N_16637,N_13043,N_14736);
nor U16638 (N_16638,N_15478,N_13168);
nand U16639 (N_16639,N_15307,N_13224);
xnor U16640 (N_16640,N_15140,N_13466);
xnor U16641 (N_16641,N_14536,N_13749);
nor U16642 (N_16642,N_14895,N_15425);
nand U16643 (N_16643,N_14995,N_14368);
and U16644 (N_16644,N_12965,N_13908);
or U16645 (N_16645,N_12973,N_12573);
or U16646 (N_16646,N_15477,N_13842);
nand U16647 (N_16647,N_13880,N_13242);
nand U16648 (N_16648,N_14479,N_13263);
and U16649 (N_16649,N_12841,N_12777);
nor U16650 (N_16650,N_14221,N_14804);
nand U16651 (N_16651,N_15168,N_13585);
xnor U16652 (N_16652,N_14304,N_15623);
or U16653 (N_16653,N_13504,N_13461);
xor U16654 (N_16654,N_15093,N_13056);
nor U16655 (N_16655,N_15414,N_12616);
nor U16656 (N_16656,N_13004,N_14842);
nor U16657 (N_16657,N_15476,N_14687);
nand U16658 (N_16658,N_14097,N_14243);
xor U16659 (N_16659,N_13904,N_13986);
nand U16660 (N_16660,N_13939,N_13888);
and U16661 (N_16661,N_12943,N_15138);
or U16662 (N_16662,N_14485,N_14854);
nor U16663 (N_16663,N_14920,N_14599);
xor U16664 (N_16664,N_15164,N_13666);
nand U16665 (N_16665,N_12633,N_13729);
nand U16666 (N_16666,N_15406,N_15046);
xor U16667 (N_16667,N_13651,N_14010);
or U16668 (N_16668,N_13822,N_14210);
xnor U16669 (N_16669,N_14805,N_15191);
and U16670 (N_16670,N_13246,N_15026);
or U16671 (N_16671,N_14205,N_13900);
and U16672 (N_16672,N_14022,N_13194);
nor U16673 (N_16673,N_13942,N_12684);
nand U16674 (N_16674,N_13207,N_15278);
or U16675 (N_16675,N_15085,N_15358);
nand U16676 (N_16676,N_15518,N_13601);
or U16677 (N_16677,N_15078,N_12648);
or U16678 (N_16678,N_14499,N_12561);
or U16679 (N_16679,N_14138,N_14672);
and U16680 (N_16680,N_14976,N_14495);
or U16681 (N_16681,N_12944,N_15309);
or U16682 (N_16682,N_13107,N_15240);
or U16683 (N_16683,N_13795,N_12835);
or U16684 (N_16684,N_14407,N_13508);
nand U16685 (N_16685,N_14714,N_14940);
nor U16686 (N_16686,N_14057,N_13693);
or U16687 (N_16687,N_14898,N_14975);
and U16688 (N_16688,N_15503,N_12658);
nand U16689 (N_16689,N_14981,N_12753);
xor U16690 (N_16690,N_14825,N_15306);
xnor U16691 (N_16691,N_14515,N_14303);
nor U16692 (N_16692,N_14905,N_13799);
or U16693 (N_16693,N_15463,N_13895);
nand U16694 (N_16694,N_13475,N_12581);
nand U16695 (N_16695,N_13753,N_15337);
nand U16696 (N_16696,N_14734,N_15305);
and U16697 (N_16697,N_12799,N_15171);
xnor U16698 (N_16698,N_13221,N_13386);
and U16699 (N_16699,N_13657,N_13783);
nor U16700 (N_16700,N_15609,N_14844);
and U16701 (N_16701,N_12718,N_15589);
or U16702 (N_16702,N_13980,N_13338);
or U16703 (N_16703,N_14801,N_15426);
nand U16704 (N_16704,N_14847,N_13330);
nand U16705 (N_16705,N_14969,N_13824);
nor U16706 (N_16706,N_14588,N_13765);
nor U16707 (N_16707,N_14843,N_15326);
or U16708 (N_16708,N_13196,N_15220);
xnor U16709 (N_16709,N_13591,N_13395);
and U16710 (N_16710,N_14878,N_13465);
xor U16711 (N_16711,N_14650,N_15429);
xnor U16712 (N_16712,N_14913,N_13073);
and U16713 (N_16713,N_12785,N_12920);
nor U16714 (N_16714,N_14720,N_13788);
nand U16715 (N_16715,N_15267,N_15241);
or U16716 (N_16716,N_13295,N_13990);
and U16717 (N_16717,N_13521,N_13448);
nand U16718 (N_16718,N_13534,N_13584);
and U16719 (N_16719,N_13607,N_12812);
nor U16720 (N_16720,N_14071,N_14367);
nor U16721 (N_16721,N_14041,N_13489);
nor U16722 (N_16722,N_14800,N_15370);
or U16723 (N_16723,N_14525,N_13668);
nand U16724 (N_16724,N_14364,N_12655);
xor U16725 (N_16725,N_13125,N_13891);
or U16726 (N_16726,N_13684,N_14758);
or U16727 (N_16727,N_15321,N_13712);
or U16728 (N_16728,N_15325,N_14270);
nand U16729 (N_16729,N_12967,N_15319);
nor U16730 (N_16730,N_12910,N_14357);
nand U16731 (N_16731,N_14921,N_14770);
or U16732 (N_16732,N_14059,N_15129);
xor U16733 (N_16733,N_13184,N_12641);
or U16734 (N_16734,N_13549,N_14716);
and U16735 (N_16735,N_14769,N_14718);
or U16736 (N_16736,N_15566,N_14711);
nor U16737 (N_16737,N_12736,N_12871);
and U16738 (N_16738,N_13202,N_14828);
and U16739 (N_16739,N_14246,N_14217);
xnor U16740 (N_16740,N_14456,N_14918);
nor U16741 (N_16741,N_15128,N_12860);
or U16742 (N_16742,N_13992,N_15417);
xor U16743 (N_16743,N_13078,N_13837);
or U16744 (N_16744,N_13542,N_14907);
or U16745 (N_16745,N_14335,N_15421);
nor U16746 (N_16746,N_14359,N_13447);
xor U16747 (N_16747,N_15144,N_13024);
or U16748 (N_16748,N_12929,N_14978);
and U16749 (N_16749,N_14578,N_13764);
or U16750 (N_16750,N_15270,N_15607);
xor U16751 (N_16751,N_13312,N_14552);
and U16752 (N_16752,N_12576,N_12702);
nor U16753 (N_16753,N_13020,N_15472);
nand U16754 (N_16754,N_12714,N_13766);
nor U16755 (N_16755,N_15366,N_14753);
xor U16756 (N_16756,N_14393,N_12584);
or U16757 (N_16757,N_14124,N_14215);
or U16758 (N_16758,N_12634,N_15418);
nor U16759 (N_16759,N_14556,N_15536);
nor U16760 (N_16760,N_14032,N_14426);
and U16761 (N_16761,N_13409,N_13894);
and U16762 (N_16762,N_13131,N_15359);
nor U16763 (N_16763,N_12677,N_14991);
nor U16764 (N_16764,N_12546,N_14287);
xnor U16765 (N_16765,N_15215,N_15010);
xor U16766 (N_16766,N_15563,N_14759);
xnor U16767 (N_16767,N_14080,N_13429);
or U16768 (N_16768,N_12626,N_14408);
nand U16769 (N_16769,N_12854,N_14036);
or U16770 (N_16770,N_14229,N_13514);
and U16771 (N_16771,N_14709,N_14574);
nand U16772 (N_16772,N_15576,N_14319);
and U16773 (N_16773,N_15544,N_15302);
nand U16774 (N_16774,N_15455,N_15432);
nor U16775 (N_16775,N_12735,N_13222);
nand U16776 (N_16776,N_13572,N_15200);
xnor U16777 (N_16777,N_14571,N_14876);
nor U16778 (N_16778,N_13318,N_15614);
nor U16779 (N_16779,N_13205,N_14727);
nand U16780 (N_16780,N_14614,N_15206);
nand U16781 (N_16781,N_13245,N_13883);
and U16782 (N_16782,N_15214,N_14896);
nor U16783 (N_16783,N_15379,N_14606);
and U16784 (N_16784,N_13101,N_15001);
nor U16785 (N_16785,N_15590,N_14848);
or U16786 (N_16786,N_15133,N_14047);
and U16787 (N_16787,N_14793,N_14797);
xnor U16788 (N_16788,N_15499,N_14583);
nand U16789 (N_16789,N_14196,N_12600);
xnor U16790 (N_16790,N_13868,N_14307);
and U16791 (N_16791,N_13383,N_14473);
nor U16792 (N_16792,N_14424,N_14970);
nor U16793 (N_16793,N_14489,N_14566);
xor U16794 (N_16794,N_14400,N_15207);
nand U16795 (N_16795,N_13156,N_13974);
xor U16796 (N_16796,N_14177,N_13851);
nor U16797 (N_16797,N_14306,N_15004);
xor U16798 (N_16798,N_13086,N_13348);
nand U16799 (N_16799,N_15482,N_14118);
nor U16800 (N_16800,N_12571,N_15135);
nand U16801 (N_16801,N_13516,N_12589);
xor U16802 (N_16802,N_12533,N_14635);
xnor U16803 (N_16803,N_13827,N_15283);
xnor U16804 (N_16804,N_12704,N_13562);
or U16805 (N_16805,N_14158,N_12915);
and U16806 (N_16806,N_14020,N_15236);
nand U16807 (N_16807,N_14945,N_14439);
nor U16808 (N_16808,N_13252,N_14390);
or U16809 (N_16809,N_14043,N_15469);
or U16810 (N_16810,N_15532,N_13943);
nor U16811 (N_16811,N_15008,N_14620);
and U16812 (N_16812,N_13646,N_13169);
xor U16813 (N_16813,N_13499,N_15351);
nor U16814 (N_16814,N_13175,N_15485);
nor U16815 (N_16815,N_14971,N_15106);
nor U16816 (N_16816,N_12548,N_14125);
nor U16817 (N_16817,N_15038,N_14320);
and U16818 (N_16818,N_12681,N_12624);
and U16819 (N_16819,N_14739,N_12923);
xor U16820 (N_16820,N_13021,N_12800);
xnor U16821 (N_16821,N_14616,N_15027);
and U16822 (N_16822,N_13444,N_12696);
nor U16823 (N_16823,N_14087,N_13761);
xor U16824 (N_16824,N_14331,N_14527);
or U16825 (N_16825,N_13833,N_12778);
xor U16826 (N_16826,N_15396,N_15450);
xor U16827 (N_16827,N_14988,N_12708);
and U16828 (N_16828,N_13268,N_14851);
nor U16829 (N_16829,N_13652,N_14729);
xnor U16830 (N_16830,N_14121,N_14598);
and U16831 (N_16831,N_13060,N_13083);
or U16832 (N_16832,N_13789,N_13013);
nor U16833 (N_16833,N_15357,N_13167);
or U16834 (N_16834,N_13846,N_14049);
nor U16835 (N_16835,N_14272,N_13587);
nand U16836 (N_16836,N_13306,N_14365);
nor U16837 (N_16837,N_13277,N_12686);
and U16838 (N_16838,N_13376,N_12604);
xor U16839 (N_16839,N_15385,N_15043);
nand U16840 (N_16840,N_14450,N_13071);
or U16841 (N_16841,N_13157,N_13282);
or U16842 (N_16842,N_14134,N_14150);
xnor U16843 (N_16843,N_12992,N_14919);
nand U16844 (N_16844,N_14044,N_13573);
or U16845 (N_16845,N_14486,N_14524);
nor U16846 (N_16846,N_14762,N_15484);
nor U16847 (N_16847,N_13632,N_15216);
or U16848 (N_16848,N_14500,N_14624);
nand U16849 (N_16849,N_14906,N_15255);
and U16850 (N_16850,N_13190,N_13671);
xnor U16851 (N_16851,N_13688,N_14546);
and U16852 (N_16852,N_13431,N_15386);
nor U16853 (N_16853,N_13449,N_14645);
or U16854 (N_16854,N_15340,N_12699);
or U16855 (N_16855,N_15624,N_14040);
nor U16856 (N_16856,N_12935,N_12744);
nand U16857 (N_16857,N_13197,N_14200);
nor U16858 (N_16858,N_12570,N_13034);
and U16859 (N_16859,N_15060,N_13353);
xor U16860 (N_16860,N_13774,N_15146);
and U16861 (N_16861,N_13767,N_15545);
nor U16862 (N_16862,N_14496,N_14011);
nor U16863 (N_16863,N_13647,N_15373);
nand U16864 (N_16864,N_13283,N_14837);
xor U16865 (N_16865,N_13008,N_13882);
xnor U16866 (N_16866,N_12531,N_13746);
nor U16867 (N_16867,N_14292,N_14181);
nand U16868 (N_16868,N_13213,N_13286);
and U16869 (N_16869,N_14449,N_13580);
xor U16870 (N_16870,N_13720,N_12885);
xnor U16871 (N_16871,N_14617,N_15569);
xor U16872 (N_16872,N_13490,N_12597);
and U16873 (N_16873,N_13051,N_13090);
nand U16874 (N_16874,N_13147,N_14728);
xor U16875 (N_16875,N_14451,N_15291);
or U16876 (N_16876,N_13085,N_12503);
or U16877 (N_16877,N_13594,N_14933);
nor U16878 (N_16878,N_14977,N_15166);
or U16879 (N_16879,N_15411,N_15384);
xnor U16880 (N_16880,N_13154,N_15551);
xor U16881 (N_16881,N_14062,N_14374);
nand U16882 (N_16882,N_12629,N_13916);
or U16883 (N_16883,N_15409,N_14254);
nor U16884 (N_16884,N_13556,N_14067);
and U16885 (N_16885,N_13568,N_15188);
and U16886 (N_16886,N_15440,N_12873);
or U16887 (N_16887,N_13673,N_13082);
and U16888 (N_16888,N_14809,N_14579);
nand U16889 (N_16889,N_15298,N_13336);
or U16890 (N_16890,N_15335,N_13708);
xor U16891 (N_16891,N_13007,N_12642);
nor U16892 (N_16892,N_15212,N_14219);
and U16893 (N_16893,N_15508,N_14637);
xor U16894 (N_16894,N_15015,N_13628);
and U16895 (N_16895,N_13825,N_14573);
nand U16896 (N_16896,N_14497,N_13410);
or U16897 (N_16897,N_14324,N_15082);
nand U16898 (N_16898,N_15612,N_15474);
and U16899 (N_16899,N_14052,N_15195);
or U16900 (N_16900,N_15272,N_14771);
or U16901 (N_16901,N_15234,N_14175);
xnor U16902 (N_16902,N_14404,N_12544);
and U16903 (N_16903,N_14354,N_15096);
or U16904 (N_16904,N_14889,N_13189);
and U16905 (N_16905,N_14608,N_13456);
or U16906 (N_16906,N_14294,N_14856);
and U16907 (N_16907,N_13406,N_13914);
xor U16908 (N_16908,N_15328,N_15557);
or U16909 (N_16909,N_12825,N_13454);
or U16910 (N_16910,N_14576,N_14008);
nand U16911 (N_16911,N_14310,N_12685);
or U16912 (N_16912,N_13446,N_15314);
nor U16913 (N_16913,N_12962,N_13779);
and U16914 (N_16914,N_14563,N_15603);
xor U16915 (N_16915,N_13243,N_13815);
xnor U16916 (N_16916,N_15176,N_12569);
xnor U16917 (N_16917,N_14326,N_15263);
or U16918 (N_16918,N_14086,N_14627);
xnor U16919 (N_16919,N_15516,N_12966);
or U16920 (N_16920,N_15377,N_15002);
and U16921 (N_16921,N_12523,N_15531);
nand U16922 (N_16922,N_12889,N_13068);
and U16923 (N_16923,N_13403,N_15274);
and U16924 (N_16924,N_14568,N_13743);
nor U16925 (N_16925,N_13063,N_13483);
nand U16926 (N_16926,N_15486,N_15347);
nor U16927 (N_16927,N_14129,N_12689);
nand U16928 (N_16928,N_13113,N_12912);
nand U16929 (N_16929,N_13485,N_15479);
or U16930 (N_16930,N_13231,N_15132);
nor U16931 (N_16931,N_13740,N_15586);
nor U16932 (N_16932,N_13792,N_13059);
nor U16933 (N_16933,N_14909,N_15553);
nand U16934 (N_16934,N_14964,N_13691);
and U16935 (N_16935,N_13754,N_12742);
nand U16936 (N_16936,N_13745,N_12877);
or U16937 (N_16937,N_15225,N_14934);
nor U16938 (N_16938,N_14575,N_15459);
nor U16939 (N_16939,N_13237,N_13254);
and U16940 (N_16940,N_15591,N_13148);
and U16941 (N_16941,N_14725,N_13631);
nand U16942 (N_16942,N_13124,N_15235);
or U16943 (N_16943,N_13702,N_14724);
nand U16944 (N_16944,N_14342,N_14487);
xnor U16945 (N_16945,N_12652,N_14811);
or U16946 (N_16946,N_14388,N_13899);
and U16947 (N_16947,N_14015,N_12773);
nand U16948 (N_16948,N_13235,N_15114);
and U16949 (N_16949,N_13289,N_15593);
and U16950 (N_16950,N_13487,N_12504);
nand U16951 (N_16951,N_14103,N_14781);
and U16952 (N_16952,N_15033,N_13962);
or U16953 (N_16953,N_13843,N_14037);
and U16954 (N_16954,N_13777,N_13727);
nand U16955 (N_16955,N_13385,N_12678);
and U16956 (N_16956,N_14698,N_14783);
and U16957 (N_16957,N_12863,N_12766);
and U16958 (N_16958,N_12790,N_14328);
and U16959 (N_16959,N_14785,N_13537);
xor U16960 (N_16960,N_13793,N_13575);
and U16961 (N_16961,N_14891,N_13065);
xnor U16962 (N_16962,N_13464,N_15102);
xor U16963 (N_16963,N_14861,N_13527);
xor U16964 (N_16964,N_14742,N_13480);
and U16965 (N_16965,N_15410,N_13344);
or U16966 (N_16966,N_12551,N_15405);
nor U16967 (N_16967,N_14126,N_12522);
and U16968 (N_16968,N_15446,N_13346);
nand U16969 (N_16969,N_13808,N_13663);
nor U16970 (N_16970,N_14025,N_14547);
and U16971 (N_16971,N_14846,N_15448);
and U16972 (N_16972,N_15227,N_15020);
nand U16973 (N_16973,N_13979,N_15399);
xor U16974 (N_16974,N_15204,N_14867);
nor U16975 (N_16975,N_13132,N_13432);
or U16976 (N_16976,N_14409,N_13281);
or U16977 (N_16977,N_12949,N_13356);
nand U16978 (N_16978,N_15205,N_14875);
nor U16979 (N_16979,N_14113,N_15304);
or U16980 (N_16980,N_14178,N_13596);
nor U16981 (N_16981,N_13510,N_15032);
xor U16982 (N_16982,N_14634,N_13153);
xnor U16983 (N_16983,N_12669,N_14750);
nand U16984 (N_16984,N_14173,N_14561);
nand U16985 (N_16985,N_14857,N_13118);
nor U16986 (N_16986,N_12666,N_12909);
nor U16987 (N_16987,N_13162,N_13248);
and U16988 (N_16988,N_13936,N_13368);
or U16989 (N_16989,N_13617,N_15470);
and U16990 (N_16990,N_14247,N_14394);
or U16991 (N_16991,N_15582,N_12932);
nand U16992 (N_16992,N_14164,N_12586);
xnor U16993 (N_16993,N_14852,N_14203);
nand U16994 (N_16994,N_14615,N_12556);
and U16995 (N_16995,N_15213,N_15527);
xnor U16996 (N_16996,N_14484,N_15187);
or U16997 (N_16997,N_15587,N_13554);
nor U16998 (N_16998,N_15395,N_13181);
or U16999 (N_16999,N_13810,N_13967);
xnor U17000 (N_17000,N_14841,N_13752);
and U17001 (N_17001,N_14779,N_13884);
or U17002 (N_17002,N_13212,N_15452);
or U17003 (N_17003,N_14470,N_14621);
nand U17004 (N_17004,N_12782,N_14209);
or U17005 (N_17005,N_12942,N_12851);
or U17006 (N_17006,N_15182,N_14382);
nor U17007 (N_17007,N_14136,N_14237);
nand U17008 (N_17008,N_14241,N_15293);
nand U17009 (N_17009,N_14702,N_12529);
xor U17010 (N_17010,N_13463,N_14042);
nand U17011 (N_17011,N_13835,N_13525);
nor U17012 (N_17012,N_15151,N_13954);
nor U17013 (N_17013,N_14984,N_12817);
and U17014 (N_17014,N_13186,N_12630);
and U17015 (N_17015,N_12746,N_14024);
nand U17016 (N_17016,N_13484,N_12964);
xnor U17017 (N_17017,N_12534,N_14666);
and U17018 (N_17018,N_14691,N_13255);
nor U17019 (N_17019,N_13977,N_15449);
nand U17020 (N_17020,N_14550,N_13412);
nor U17021 (N_17021,N_13643,N_12751);
nor U17022 (N_17022,N_12793,N_14000);
xnor U17023 (N_17023,N_13721,N_14061);
nor U17024 (N_17024,N_12517,N_13417);
nor U17025 (N_17025,N_15013,N_14507);
xnor U17026 (N_17026,N_13964,N_15245);
xnor U17027 (N_17027,N_15028,N_12895);
xor U17028 (N_17028,N_13780,N_14685);
or U17029 (N_17029,N_13257,N_12819);
nor U17030 (N_17030,N_14261,N_13011);
nand U17031 (N_17031,N_12733,N_14395);
nor U17032 (N_17032,N_14476,N_14654);
nand U17033 (N_17033,N_13787,N_14091);
nor U17034 (N_17034,N_14999,N_13416);
and U17035 (N_17035,N_14316,N_12765);
xnor U17036 (N_17036,N_14222,N_14773);
or U17037 (N_17037,N_13797,N_13920);
nand U17038 (N_17038,N_12898,N_15434);
nand U17039 (N_17039,N_14565,N_12515);
xnor U17040 (N_17040,N_13393,N_14796);
and U17041 (N_17041,N_13334,N_13217);
nand U17042 (N_17042,N_14707,N_13728);
and U17043 (N_17043,N_14230,N_14812);
or U17044 (N_17044,N_12713,N_15439);
and U17045 (N_17045,N_15320,N_13320);
or U17046 (N_17046,N_13823,N_14908);
and U17047 (N_17047,N_14609,N_14263);
nor U17048 (N_17048,N_13700,N_12815);
xor U17049 (N_17049,N_13006,N_12955);
and U17050 (N_17050,N_13182,N_14100);
nand U17051 (N_17051,N_14743,N_12628);
and U17052 (N_17052,N_12680,N_14378);
or U17053 (N_17053,N_14510,N_15308);
and U17054 (N_17054,N_14313,N_13130);
or U17055 (N_17055,N_13778,N_14652);
xor U17056 (N_17056,N_12866,N_13614);
nand U17057 (N_17057,N_12750,N_13775);
xor U17058 (N_17058,N_13350,N_13599);
nor U17059 (N_17059,N_15608,N_12660);
or U17060 (N_17060,N_14986,N_13458);
nand U17061 (N_17061,N_14972,N_13325);
xor U17062 (N_17062,N_12834,N_15618);
nand U17063 (N_17063,N_13863,N_13009);
and U17064 (N_17064,N_13445,N_12795);
nor U17065 (N_17065,N_14639,N_14938);
or U17066 (N_17066,N_13290,N_14046);
nand U17067 (N_17067,N_15072,N_14760);
nand U17068 (N_17068,N_13477,N_15360);
xor U17069 (N_17069,N_14144,N_14195);
and U17070 (N_17070,N_13080,N_15537);
and U17071 (N_17071,N_13741,N_14079);
nor U17072 (N_17072,N_13276,N_13144);
xor U17073 (N_17073,N_13866,N_14798);
nand U17074 (N_17074,N_14826,N_13048);
or U17075 (N_17075,N_15621,N_13408);
xor U17076 (N_17076,N_13918,N_13593);
nand U17077 (N_17077,N_13886,N_14208);
xor U17078 (N_17078,N_12792,N_13496);
nand U17079 (N_17079,N_14776,N_14863);
and U17080 (N_17080,N_13332,N_14679);
nor U17081 (N_17081,N_14722,N_15343);
and U17082 (N_17082,N_13816,N_14572);
or U17083 (N_17083,N_13275,N_15071);
or U17084 (N_17084,N_15402,N_12894);
nand U17085 (N_17085,N_13770,N_13001);
or U17086 (N_17086,N_14658,N_13112);
nor U17087 (N_17087,N_13633,N_13561);
and U17088 (N_17088,N_14276,N_12855);
nor U17089 (N_17089,N_15125,N_12829);
xor U17090 (N_17090,N_14028,N_14632);
xor U17091 (N_17091,N_13303,N_14974);
and U17092 (N_17092,N_13865,N_12614);
and U17093 (N_17093,N_14548,N_13361);
or U17094 (N_17094,N_14017,N_15076);
xor U17095 (N_17095,N_14092,N_14163);
xnor U17096 (N_17096,N_13170,N_14605);
or U17097 (N_17097,N_12827,N_14537);
nand U17098 (N_17098,N_13906,N_14631);
nand U17099 (N_17099,N_15487,N_13533);
nor U17100 (N_17100,N_13206,N_14133);
nand U17101 (N_17101,N_13893,N_12803);
or U17102 (N_17102,N_14014,N_14419);
xnor U17103 (N_17103,N_14155,N_14389);
xor U17104 (N_17104,N_13374,N_14942);
nor U17105 (N_17105,N_15355,N_14279);
xnor U17106 (N_17106,N_14048,N_14562);
xnor U17107 (N_17107,N_12908,N_14314);
nand U17108 (N_17108,N_13896,N_14534);
xnor U17109 (N_17109,N_13176,N_12710);
nor U17110 (N_17110,N_15488,N_15111);
or U17111 (N_17111,N_14962,N_12963);
xnor U17112 (N_17112,N_12813,N_12758);
and U17113 (N_17113,N_14060,N_12543);
nand U17114 (N_17114,N_15141,N_15069);
xnor U17115 (N_17115,N_14257,N_13707);
nand U17116 (N_17116,N_13619,N_12693);
or U17117 (N_17117,N_14392,N_14989);
and U17118 (N_17118,N_13574,N_14833);
xor U17119 (N_17119,N_14455,N_14171);
nand U17120 (N_17120,N_13039,N_15068);
xor U17121 (N_17121,N_12783,N_12542);
nand U17122 (N_17122,N_14864,N_15296);
xor U17123 (N_17123,N_14386,N_15579);
nand U17124 (N_17124,N_14433,N_15152);
xnor U17125 (N_17125,N_14664,N_13075);
xnor U17126 (N_17126,N_14564,N_14443);
or U17127 (N_17127,N_15600,N_14031);
xor U17128 (N_17128,N_13582,N_14447);
and U17129 (N_17129,N_15408,N_13140);
nand U17130 (N_17130,N_12784,N_15419);
nor U17131 (N_17131,N_14003,N_15239);
nor U17132 (N_17132,N_13262,N_12982);
nor U17133 (N_17133,N_12559,N_15287);
nor U17134 (N_17134,N_14102,N_13940);
and U17135 (N_17135,N_14239,N_15615);
and U17136 (N_17136,N_12565,N_14674);
or U17137 (N_17137,N_14380,N_14932);
or U17138 (N_17138,N_14051,N_14838);
nor U17139 (N_17139,N_13381,N_13399);
and U17140 (N_17140,N_12537,N_13321);
nor U17141 (N_17141,N_15515,N_14656);
nor U17142 (N_17142,N_13470,N_15394);
nor U17143 (N_17143,N_13859,N_13301);
nor U17144 (N_17144,N_14647,N_12821);
xnor U17145 (N_17145,N_12554,N_14594);
xor U17146 (N_17146,N_14532,N_12938);
nor U17147 (N_17147,N_13166,N_15380);
nor U17148 (N_17148,N_13143,N_15595);
or U17149 (N_17149,N_15189,N_12781);
nand U17150 (N_17150,N_13457,N_13314);
xnor U17151 (N_17151,N_13790,N_13058);
nor U17152 (N_17152,N_15542,N_14418);
nand U17153 (N_17153,N_15119,N_15194);
or U17154 (N_17154,N_13091,N_15513);
xor U17155 (N_17155,N_14517,N_14570);
or U17156 (N_17156,N_12756,N_12739);
or U17157 (N_17157,N_12661,N_14839);
or U17158 (N_17158,N_12760,N_14726);
and U17159 (N_17159,N_13911,N_12528);
nand U17160 (N_17160,N_15303,N_13949);
nand U17161 (N_17161,N_13331,N_13760);
and U17162 (N_17162,N_13999,N_15224);
xnor U17163 (N_17163,N_13250,N_13981);
nor U17164 (N_17164,N_14353,N_15127);
or U17165 (N_17165,N_12981,N_13636);
xnor U17166 (N_17166,N_15403,N_14301);
and U17167 (N_17167,N_15529,N_15247);
nand U17168 (N_17168,N_13253,N_15580);
and U17169 (N_17169,N_13984,N_14198);
or U17170 (N_17170,N_15190,N_12653);
and U17171 (N_17171,N_12772,N_15540);
and U17172 (N_17172,N_13944,N_14611);
xnor U17173 (N_17173,N_14535,N_12934);
xor U17174 (N_17174,N_12759,N_14591);
xor U17175 (N_17175,N_15442,N_14213);
xor U17176 (N_17176,N_14636,N_13848);
xnor U17177 (N_17177,N_14371,N_12839);
or U17178 (N_17178,N_12918,N_13309);
or U17179 (N_17179,N_15374,N_14721);
xor U17180 (N_17180,N_14956,N_12743);
or U17181 (N_17181,N_13115,N_12602);
and U17182 (N_17182,N_15064,N_15193);
nor U17183 (N_17183,N_14849,N_13800);
and U17184 (N_17184,N_15201,N_14998);
and U17185 (N_17185,N_13929,N_13373);
xnor U17186 (N_17186,N_15222,N_14601);
and U17187 (N_17187,N_13472,N_15227);
and U17188 (N_17188,N_13107,N_15054);
nand U17189 (N_17189,N_15502,N_14637);
xor U17190 (N_17190,N_12986,N_13190);
xnor U17191 (N_17191,N_13536,N_12872);
nand U17192 (N_17192,N_13392,N_15348);
xor U17193 (N_17193,N_14598,N_14464);
and U17194 (N_17194,N_13798,N_14849);
or U17195 (N_17195,N_12827,N_14287);
nand U17196 (N_17196,N_14516,N_13066);
and U17197 (N_17197,N_15373,N_12685);
nand U17198 (N_17198,N_13603,N_12988);
or U17199 (N_17199,N_14225,N_12978);
xnor U17200 (N_17200,N_13405,N_13847);
xnor U17201 (N_17201,N_13521,N_12877);
xor U17202 (N_17202,N_13141,N_12885);
xnor U17203 (N_17203,N_13361,N_12824);
nor U17204 (N_17204,N_13734,N_13719);
xnor U17205 (N_17205,N_13922,N_12870);
xnor U17206 (N_17206,N_14183,N_15165);
nor U17207 (N_17207,N_13898,N_14916);
and U17208 (N_17208,N_12591,N_12949);
nand U17209 (N_17209,N_13496,N_12730);
nor U17210 (N_17210,N_12505,N_14722);
xnor U17211 (N_17211,N_13292,N_14629);
and U17212 (N_17212,N_12941,N_13837);
xnor U17213 (N_17213,N_15472,N_15471);
xor U17214 (N_17214,N_12863,N_14439);
xor U17215 (N_17215,N_12866,N_13194);
xor U17216 (N_17216,N_12553,N_14255);
and U17217 (N_17217,N_14382,N_15595);
nand U17218 (N_17218,N_14121,N_14852);
nor U17219 (N_17219,N_13345,N_13868);
nand U17220 (N_17220,N_13734,N_13331);
xor U17221 (N_17221,N_14901,N_14801);
nand U17222 (N_17222,N_15295,N_13069);
xnor U17223 (N_17223,N_15583,N_14018);
and U17224 (N_17224,N_13654,N_14062);
or U17225 (N_17225,N_14692,N_14738);
or U17226 (N_17226,N_15502,N_12969);
nand U17227 (N_17227,N_15048,N_13228);
xnor U17228 (N_17228,N_13154,N_13345);
or U17229 (N_17229,N_14412,N_14510);
xor U17230 (N_17230,N_14696,N_14640);
nand U17231 (N_17231,N_13411,N_13082);
or U17232 (N_17232,N_14393,N_13990);
or U17233 (N_17233,N_15113,N_13686);
nand U17234 (N_17234,N_13164,N_15565);
xor U17235 (N_17235,N_14642,N_14678);
xnor U17236 (N_17236,N_15420,N_13084);
xor U17237 (N_17237,N_14588,N_12657);
nand U17238 (N_17238,N_14749,N_13589);
nor U17239 (N_17239,N_15279,N_15231);
or U17240 (N_17240,N_14460,N_13279);
xor U17241 (N_17241,N_13549,N_15061);
or U17242 (N_17242,N_14591,N_13301);
nor U17243 (N_17243,N_13973,N_14566);
xor U17244 (N_17244,N_14819,N_14342);
nor U17245 (N_17245,N_14504,N_15266);
nand U17246 (N_17246,N_13862,N_12723);
or U17247 (N_17247,N_14387,N_15093);
xor U17248 (N_17248,N_15051,N_13941);
nand U17249 (N_17249,N_13828,N_13028);
nand U17250 (N_17250,N_12714,N_15050);
xor U17251 (N_17251,N_12656,N_15400);
or U17252 (N_17252,N_12803,N_13161);
xnor U17253 (N_17253,N_13569,N_15471);
or U17254 (N_17254,N_15067,N_14590);
xnor U17255 (N_17255,N_15036,N_14580);
xor U17256 (N_17256,N_14209,N_15430);
nor U17257 (N_17257,N_13955,N_14146);
or U17258 (N_17258,N_14392,N_13598);
nand U17259 (N_17259,N_13412,N_12939);
xnor U17260 (N_17260,N_15515,N_14545);
or U17261 (N_17261,N_14099,N_14699);
or U17262 (N_17262,N_12754,N_14795);
nand U17263 (N_17263,N_12581,N_14744);
xnor U17264 (N_17264,N_15128,N_13846);
and U17265 (N_17265,N_14798,N_12573);
nor U17266 (N_17266,N_13376,N_14171);
and U17267 (N_17267,N_13525,N_13351);
nor U17268 (N_17268,N_15164,N_14455);
nand U17269 (N_17269,N_14478,N_14401);
and U17270 (N_17270,N_15623,N_13738);
or U17271 (N_17271,N_15270,N_15227);
or U17272 (N_17272,N_15525,N_14606);
nor U17273 (N_17273,N_14236,N_12951);
nand U17274 (N_17274,N_15519,N_13085);
and U17275 (N_17275,N_12732,N_15236);
nand U17276 (N_17276,N_14596,N_13693);
or U17277 (N_17277,N_13333,N_15160);
nor U17278 (N_17278,N_15040,N_13713);
and U17279 (N_17279,N_14660,N_14535);
nor U17280 (N_17280,N_13113,N_12887);
or U17281 (N_17281,N_14934,N_14461);
and U17282 (N_17282,N_13018,N_12927);
nand U17283 (N_17283,N_13748,N_14392);
and U17284 (N_17284,N_15529,N_12650);
nor U17285 (N_17285,N_14286,N_14786);
nor U17286 (N_17286,N_15383,N_14123);
xor U17287 (N_17287,N_12506,N_12801);
or U17288 (N_17288,N_14515,N_14510);
and U17289 (N_17289,N_15456,N_12776);
nand U17290 (N_17290,N_14329,N_13369);
and U17291 (N_17291,N_13273,N_14434);
nand U17292 (N_17292,N_14666,N_14737);
or U17293 (N_17293,N_13622,N_13832);
nand U17294 (N_17294,N_13487,N_14341);
and U17295 (N_17295,N_14455,N_12730);
nor U17296 (N_17296,N_14558,N_15060);
or U17297 (N_17297,N_14311,N_14269);
nor U17298 (N_17298,N_13955,N_14838);
nor U17299 (N_17299,N_13580,N_14364);
and U17300 (N_17300,N_14469,N_13583);
or U17301 (N_17301,N_12755,N_13792);
nor U17302 (N_17302,N_14140,N_15153);
and U17303 (N_17303,N_13001,N_12859);
or U17304 (N_17304,N_14498,N_13056);
xor U17305 (N_17305,N_14168,N_13673);
or U17306 (N_17306,N_14282,N_12564);
and U17307 (N_17307,N_12848,N_14390);
nand U17308 (N_17308,N_12870,N_14563);
xnor U17309 (N_17309,N_13832,N_15357);
nand U17310 (N_17310,N_15336,N_12591);
xnor U17311 (N_17311,N_15512,N_15347);
and U17312 (N_17312,N_15350,N_13264);
or U17313 (N_17313,N_15319,N_13322);
nor U17314 (N_17314,N_13795,N_13759);
nor U17315 (N_17315,N_15087,N_13273);
or U17316 (N_17316,N_12665,N_14175);
or U17317 (N_17317,N_15357,N_13014);
nand U17318 (N_17318,N_15524,N_13152);
nand U17319 (N_17319,N_14742,N_14286);
xor U17320 (N_17320,N_12816,N_12977);
nor U17321 (N_17321,N_14450,N_15127);
nand U17322 (N_17322,N_13018,N_13491);
and U17323 (N_17323,N_13271,N_12595);
and U17324 (N_17324,N_15284,N_12732);
nand U17325 (N_17325,N_15511,N_14269);
or U17326 (N_17326,N_13647,N_15018);
nand U17327 (N_17327,N_12927,N_12772);
nor U17328 (N_17328,N_14229,N_13165);
nand U17329 (N_17329,N_15046,N_12629);
or U17330 (N_17330,N_14923,N_15024);
nand U17331 (N_17331,N_13241,N_13736);
or U17332 (N_17332,N_15327,N_12524);
nor U17333 (N_17333,N_15011,N_15237);
xor U17334 (N_17334,N_15525,N_15508);
or U17335 (N_17335,N_15148,N_15129);
xnor U17336 (N_17336,N_15261,N_12996);
nand U17337 (N_17337,N_15053,N_13379);
nor U17338 (N_17338,N_14722,N_12528);
and U17339 (N_17339,N_13260,N_12761);
xor U17340 (N_17340,N_15317,N_13665);
or U17341 (N_17341,N_12533,N_14402);
nand U17342 (N_17342,N_13937,N_15292);
nand U17343 (N_17343,N_14259,N_15050);
nand U17344 (N_17344,N_14236,N_14908);
nor U17345 (N_17345,N_15552,N_13853);
and U17346 (N_17346,N_14368,N_13981);
and U17347 (N_17347,N_14809,N_14600);
nand U17348 (N_17348,N_14229,N_13940);
or U17349 (N_17349,N_14214,N_14057);
and U17350 (N_17350,N_13499,N_13760);
xor U17351 (N_17351,N_14113,N_13847);
nand U17352 (N_17352,N_13584,N_15119);
or U17353 (N_17353,N_15294,N_14169);
xnor U17354 (N_17354,N_15142,N_12780);
or U17355 (N_17355,N_13882,N_13304);
nor U17356 (N_17356,N_14591,N_14997);
nor U17357 (N_17357,N_14965,N_13421);
or U17358 (N_17358,N_14572,N_14580);
nor U17359 (N_17359,N_12943,N_13966);
or U17360 (N_17360,N_13871,N_14662);
and U17361 (N_17361,N_13474,N_14139);
and U17362 (N_17362,N_14229,N_15182);
nor U17363 (N_17363,N_14650,N_14309);
xnor U17364 (N_17364,N_14525,N_14133);
and U17365 (N_17365,N_14879,N_15403);
xor U17366 (N_17366,N_14658,N_12945);
or U17367 (N_17367,N_14104,N_13457);
and U17368 (N_17368,N_15025,N_14242);
or U17369 (N_17369,N_15480,N_12955);
nor U17370 (N_17370,N_12882,N_15608);
and U17371 (N_17371,N_14725,N_13639);
nand U17372 (N_17372,N_13469,N_15289);
or U17373 (N_17373,N_12842,N_14527);
xor U17374 (N_17374,N_14198,N_15284);
nand U17375 (N_17375,N_15624,N_12668);
and U17376 (N_17376,N_15062,N_14420);
xnor U17377 (N_17377,N_12585,N_14866);
nand U17378 (N_17378,N_13175,N_14060);
and U17379 (N_17379,N_14449,N_14761);
nand U17380 (N_17380,N_13656,N_14492);
or U17381 (N_17381,N_14821,N_12910);
xnor U17382 (N_17382,N_13663,N_13865);
nor U17383 (N_17383,N_14355,N_13204);
xnor U17384 (N_17384,N_12852,N_14277);
or U17385 (N_17385,N_12779,N_14830);
and U17386 (N_17386,N_13331,N_14239);
or U17387 (N_17387,N_13697,N_13350);
or U17388 (N_17388,N_14791,N_13950);
and U17389 (N_17389,N_13920,N_14726);
nor U17390 (N_17390,N_14671,N_14449);
and U17391 (N_17391,N_14887,N_15219);
nor U17392 (N_17392,N_14195,N_13102);
nand U17393 (N_17393,N_14005,N_14254);
nor U17394 (N_17394,N_13397,N_13313);
and U17395 (N_17395,N_12883,N_13062);
or U17396 (N_17396,N_15426,N_13095);
xor U17397 (N_17397,N_15247,N_14524);
nor U17398 (N_17398,N_12937,N_14960);
xnor U17399 (N_17399,N_12914,N_13954);
or U17400 (N_17400,N_13704,N_13651);
and U17401 (N_17401,N_13150,N_13344);
nor U17402 (N_17402,N_14708,N_14958);
xnor U17403 (N_17403,N_14938,N_14212);
xor U17404 (N_17404,N_14568,N_13841);
nand U17405 (N_17405,N_13413,N_13991);
nand U17406 (N_17406,N_13571,N_12845);
or U17407 (N_17407,N_12934,N_15382);
xnor U17408 (N_17408,N_14781,N_14506);
nor U17409 (N_17409,N_14426,N_13091);
nor U17410 (N_17410,N_14012,N_13444);
or U17411 (N_17411,N_15439,N_15134);
or U17412 (N_17412,N_14624,N_14213);
or U17413 (N_17413,N_13692,N_13449);
nand U17414 (N_17414,N_15539,N_15314);
xor U17415 (N_17415,N_14636,N_14475);
or U17416 (N_17416,N_12660,N_14566);
and U17417 (N_17417,N_13353,N_13546);
xnor U17418 (N_17418,N_14210,N_14871);
or U17419 (N_17419,N_12725,N_14798);
xnor U17420 (N_17420,N_13266,N_13618);
nand U17421 (N_17421,N_13305,N_15261);
nand U17422 (N_17422,N_13004,N_13630);
nor U17423 (N_17423,N_13642,N_12839);
nor U17424 (N_17424,N_14568,N_14134);
nand U17425 (N_17425,N_12709,N_13448);
nand U17426 (N_17426,N_13126,N_15441);
nor U17427 (N_17427,N_15404,N_13243);
or U17428 (N_17428,N_14026,N_13001);
xnor U17429 (N_17429,N_12503,N_13506);
nand U17430 (N_17430,N_12815,N_13097);
nand U17431 (N_17431,N_15194,N_13643);
and U17432 (N_17432,N_14089,N_13317);
and U17433 (N_17433,N_14385,N_14796);
or U17434 (N_17434,N_14298,N_15374);
nor U17435 (N_17435,N_12657,N_14452);
or U17436 (N_17436,N_15056,N_12986);
nor U17437 (N_17437,N_12882,N_12645);
nand U17438 (N_17438,N_14750,N_14482);
or U17439 (N_17439,N_12760,N_14305);
nand U17440 (N_17440,N_13483,N_13623);
nand U17441 (N_17441,N_14401,N_15167);
nor U17442 (N_17442,N_13938,N_12915);
nand U17443 (N_17443,N_13010,N_13851);
and U17444 (N_17444,N_13186,N_15191);
nand U17445 (N_17445,N_13900,N_14332);
or U17446 (N_17446,N_12770,N_13143);
or U17447 (N_17447,N_12843,N_12707);
xor U17448 (N_17448,N_13795,N_13561);
nor U17449 (N_17449,N_12689,N_14838);
xor U17450 (N_17450,N_13158,N_15245);
xor U17451 (N_17451,N_13948,N_15499);
or U17452 (N_17452,N_14348,N_12729);
and U17453 (N_17453,N_15475,N_12955);
or U17454 (N_17454,N_15221,N_14619);
nor U17455 (N_17455,N_13532,N_13074);
and U17456 (N_17456,N_15444,N_12573);
or U17457 (N_17457,N_12823,N_13313);
nor U17458 (N_17458,N_12609,N_14895);
nor U17459 (N_17459,N_15405,N_14722);
nor U17460 (N_17460,N_15064,N_13671);
nor U17461 (N_17461,N_13892,N_15458);
xnor U17462 (N_17462,N_14732,N_15583);
nand U17463 (N_17463,N_14661,N_15532);
and U17464 (N_17464,N_13127,N_14483);
xor U17465 (N_17465,N_14306,N_14622);
nand U17466 (N_17466,N_14938,N_15043);
nor U17467 (N_17467,N_13015,N_13808);
nor U17468 (N_17468,N_14881,N_14662);
and U17469 (N_17469,N_15423,N_15454);
nor U17470 (N_17470,N_12875,N_14406);
or U17471 (N_17471,N_12739,N_14905);
and U17472 (N_17472,N_13996,N_12680);
xnor U17473 (N_17473,N_13613,N_13187);
nand U17474 (N_17474,N_14838,N_14811);
or U17475 (N_17475,N_14542,N_15437);
nand U17476 (N_17476,N_12569,N_13285);
nor U17477 (N_17477,N_14186,N_14091);
nor U17478 (N_17478,N_14820,N_13897);
nor U17479 (N_17479,N_14955,N_13945);
xor U17480 (N_17480,N_15248,N_12813);
nand U17481 (N_17481,N_14280,N_14165);
nor U17482 (N_17482,N_13194,N_13819);
xnor U17483 (N_17483,N_14009,N_15346);
xnor U17484 (N_17484,N_15125,N_13118);
and U17485 (N_17485,N_12889,N_13195);
nand U17486 (N_17486,N_13461,N_12976);
nand U17487 (N_17487,N_14228,N_13349);
nor U17488 (N_17488,N_14232,N_14549);
or U17489 (N_17489,N_15003,N_14151);
nand U17490 (N_17490,N_12654,N_15358);
and U17491 (N_17491,N_13420,N_12842);
nor U17492 (N_17492,N_12865,N_15500);
and U17493 (N_17493,N_13480,N_13051);
nand U17494 (N_17494,N_14836,N_13171);
xnor U17495 (N_17495,N_13804,N_15177);
or U17496 (N_17496,N_13701,N_14987);
or U17497 (N_17497,N_15229,N_14954);
nand U17498 (N_17498,N_13731,N_15056);
or U17499 (N_17499,N_13747,N_14614);
and U17500 (N_17500,N_14454,N_14313);
nor U17501 (N_17501,N_13689,N_14619);
nand U17502 (N_17502,N_15094,N_14083);
nand U17503 (N_17503,N_13953,N_15455);
or U17504 (N_17504,N_12689,N_13335);
or U17505 (N_17505,N_13099,N_13356);
or U17506 (N_17506,N_15538,N_13427);
nand U17507 (N_17507,N_13196,N_13693);
and U17508 (N_17508,N_15331,N_12604);
nor U17509 (N_17509,N_12735,N_14545);
nand U17510 (N_17510,N_14253,N_13333);
or U17511 (N_17511,N_15080,N_13268);
nand U17512 (N_17512,N_13862,N_13547);
and U17513 (N_17513,N_14951,N_13361);
or U17514 (N_17514,N_13284,N_15086);
nor U17515 (N_17515,N_13977,N_13969);
or U17516 (N_17516,N_13018,N_15000);
nor U17517 (N_17517,N_14010,N_14995);
nor U17518 (N_17518,N_13475,N_14097);
nor U17519 (N_17519,N_14756,N_13599);
or U17520 (N_17520,N_14954,N_12571);
or U17521 (N_17521,N_14336,N_12875);
and U17522 (N_17522,N_15082,N_15263);
or U17523 (N_17523,N_15606,N_12545);
nor U17524 (N_17524,N_14607,N_12853);
or U17525 (N_17525,N_12684,N_14607);
and U17526 (N_17526,N_14456,N_13371);
or U17527 (N_17527,N_14935,N_13082);
or U17528 (N_17528,N_14491,N_14967);
or U17529 (N_17529,N_15402,N_15220);
or U17530 (N_17530,N_12684,N_13056);
nand U17531 (N_17531,N_14637,N_13536);
nand U17532 (N_17532,N_15209,N_13679);
and U17533 (N_17533,N_14497,N_15001);
nor U17534 (N_17534,N_15063,N_12747);
and U17535 (N_17535,N_13654,N_14039);
nor U17536 (N_17536,N_15620,N_13946);
and U17537 (N_17537,N_12718,N_13016);
and U17538 (N_17538,N_13977,N_13134);
nand U17539 (N_17539,N_14263,N_15497);
nand U17540 (N_17540,N_12608,N_12735);
xnor U17541 (N_17541,N_14674,N_15113);
or U17542 (N_17542,N_12948,N_14516);
or U17543 (N_17543,N_14497,N_14619);
nand U17544 (N_17544,N_12902,N_13887);
nor U17545 (N_17545,N_13389,N_14834);
xnor U17546 (N_17546,N_12806,N_15547);
nand U17547 (N_17547,N_15165,N_15475);
or U17548 (N_17548,N_15501,N_15224);
nor U17549 (N_17549,N_13025,N_14730);
or U17550 (N_17550,N_14820,N_12778);
nand U17551 (N_17551,N_13639,N_12737);
or U17552 (N_17552,N_12810,N_14838);
or U17553 (N_17553,N_15370,N_13903);
xor U17554 (N_17554,N_14432,N_12886);
and U17555 (N_17555,N_14406,N_12975);
nor U17556 (N_17556,N_14070,N_15271);
or U17557 (N_17557,N_12720,N_15510);
xor U17558 (N_17558,N_13964,N_13923);
nand U17559 (N_17559,N_13338,N_15442);
or U17560 (N_17560,N_13486,N_13473);
xor U17561 (N_17561,N_14047,N_14814);
nor U17562 (N_17562,N_13047,N_15546);
nand U17563 (N_17563,N_14989,N_12835);
nor U17564 (N_17564,N_13887,N_13584);
and U17565 (N_17565,N_14091,N_15089);
nor U17566 (N_17566,N_14810,N_14415);
nand U17567 (N_17567,N_15286,N_13581);
nor U17568 (N_17568,N_13613,N_13960);
or U17569 (N_17569,N_15470,N_13646);
xnor U17570 (N_17570,N_14901,N_13714);
xor U17571 (N_17571,N_14906,N_15071);
xor U17572 (N_17572,N_14930,N_13258);
nor U17573 (N_17573,N_13625,N_12835);
nand U17574 (N_17574,N_14417,N_12543);
nand U17575 (N_17575,N_14353,N_14069);
and U17576 (N_17576,N_13798,N_13866);
nor U17577 (N_17577,N_14313,N_12554);
and U17578 (N_17578,N_15178,N_12870);
and U17579 (N_17579,N_14619,N_13562);
or U17580 (N_17580,N_15097,N_14809);
and U17581 (N_17581,N_15316,N_15254);
xor U17582 (N_17582,N_13632,N_14860);
nor U17583 (N_17583,N_13495,N_14079);
nand U17584 (N_17584,N_13674,N_14223);
xnor U17585 (N_17585,N_14582,N_14369);
or U17586 (N_17586,N_14858,N_13094);
and U17587 (N_17587,N_14060,N_15353);
nand U17588 (N_17588,N_15440,N_13015);
or U17589 (N_17589,N_15239,N_13157);
xnor U17590 (N_17590,N_14109,N_14012);
nand U17591 (N_17591,N_13418,N_13066);
and U17592 (N_17592,N_12768,N_13568);
nand U17593 (N_17593,N_15439,N_14003);
nor U17594 (N_17594,N_13787,N_14699);
xor U17595 (N_17595,N_13254,N_15312);
nor U17596 (N_17596,N_13356,N_15120);
nand U17597 (N_17597,N_13418,N_12895);
nand U17598 (N_17598,N_14525,N_13223);
and U17599 (N_17599,N_13719,N_14998);
xnor U17600 (N_17600,N_15572,N_14416);
or U17601 (N_17601,N_14903,N_13177);
and U17602 (N_17602,N_13766,N_14233);
or U17603 (N_17603,N_14966,N_14749);
nand U17604 (N_17604,N_14561,N_15155);
or U17605 (N_17605,N_14169,N_12943);
and U17606 (N_17606,N_14207,N_13227);
nand U17607 (N_17607,N_14521,N_13561);
and U17608 (N_17608,N_12560,N_13713);
or U17609 (N_17609,N_14261,N_14458);
nand U17610 (N_17610,N_14411,N_12626);
and U17611 (N_17611,N_14659,N_14715);
nand U17612 (N_17612,N_14143,N_13297);
xor U17613 (N_17613,N_13151,N_15484);
or U17614 (N_17614,N_12511,N_12998);
nor U17615 (N_17615,N_15480,N_14161);
nand U17616 (N_17616,N_14937,N_13660);
or U17617 (N_17617,N_12795,N_12663);
nand U17618 (N_17618,N_14324,N_13490);
nor U17619 (N_17619,N_14308,N_15291);
nor U17620 (N_17620,N_12676,N_13786);
xor U17621 (N_17621,N_14262,N_14101);
xnor U17622 (N_17622,N_13459,N_13111);
or U17623 (N_17623,N_13745,N_15343);
and U17624 (N_17624,N_15244,N_15559);
and U17625 (N_17625,N_15499,N_15148);
nand U17626 (N_17626,N_12811,N_12947);
nor U17627 (N_17627,N_14733,N_15276);
nand U17628 (N_17628,N_12918,N_14859);
or U17629 (N_17629,N_12619,N_14306);
xor U17630 (N_17630,N_13586,N_14440);
or U17631 (N_17631,N_12666,N_14966);
nor U17632 (N_17632,N_12762,N_14524);
or U17633 (N_17633,N_12574,N_13251);
nor U17634 (N_17634,N_14472,N_12521);
xor U17635 (N_17635,N_13812,N_15203);
nand U17636 (N_17636,N_13450,N_15236);
or U17637 (N_17637,N_14509,N_15166);
and U17638 (N_17638,N_15361,N_13762);
and U17639 (N_17639,N_13360,N_12973);
nand U17640 (N_17640,N_14378,N_14875);
xnor U17641 (N_17641,N_12554,N_12596);
or U17642 (N_17642,N_14310,N_12982);
nor U17643 (N_17643,N_12591,N_13820);
or U17644 (N_17644,N_14582,N_12938);
nand U17645 (N_17645,N_14761,N_14846);
or U17646 (N_17646,N_14461,N_14540);
nor U17647 (N_17647,N_13965,N_14703);
and U17648 (N_17648,N_13148,N_12887);
xnor U17649 (N_17649,N_14313,N_15362);
nor U17650 (N_17650,N_13547,N_14791);
nor U17651 (N_17651,N_14396,N_14950);
nand U17652 (N_17652,N_13904,N_15170);
xnor U17653 (N_17653,N_14396,N_12651);
and U17654 (N_17654,N_14970,N_12997);
nor U17655 (N_17655,N_14360,N_12516);
or U17656 (N_17656,N_14649,N_13727);
xnor U17657 (N_17657,N_13464,N_15213);
nand U17658 (N_17658,N_12680,N_14493);
nand U17659 (N_17659,N_13758,N_14059);
nor U17660 (N_17660,N_14407,N_13201);
xor U17661 (N_17661,N_13121,N_14547);
nor U17662 (N_17662,N_13275,N_13229);
nor U17663 (N_17663,N_14430,N_14166);
nor U17664 (N_17664,N_15257,N_15083);
xnor U17665 (N_17665,N_13332,N_14695);
and U17666 (N_17666,N_13223,N_12885);
nor U17667 (N_17667,N_13738,N_15179);
and U17668 (N_17668,N_13997,N_12967);
xnor U17669 (N_17669,N_14035,N_12504);
nand U17670 (N_17670,N_15098,N_13247);
xnor U17671 (N_17671,N_13913,N_15129);
nand U17672 (N_17672,N_13851,N_13769);
nor U17673 (N_17673,N_14291,N_13533);
or U17674 (N_17674,N_15066,N_13864);
nor U17675 (N_17675,N_13493,N_13759);
nand U17676 (N_17676,N_14730,N_13278);
xor U17677 (N_17677,N_14607,N_14270);
or U17678 (N_17678,N_13449,N_12517);
and U17679 (N_17679,N_14043,N_12599);
or U17680 (N_17680,N_14297,N_13531);
and U17681 (N_17681,N_13324,N_14670);
nor U17682 (N_17682,N_14421,N_14080);
nor U17683 (N_17683,N_13331,N_13058);
xor U17684 (N_17684,N_14509,N_12938);
or U17685 (N_17685,N_12644,N_13693);
nand U17686 (N_17686,N_13790,N_14504);
and U17687 (N_17687,N_14910,N_13511);
or U17688 (N_17688,N_15012,N_15350);
or U17689 (N_17689,N_13480,N_13110);
nor U17690 (N_17690,N_15585,N_14541);
and U17691 (N_17691,N_15348,N_13755);
or U17692 (N_17692,N_15411,N_13986);
xor U17693 (N_17693,N_12588,N_14336);
xor U17694 (N_17694,N_13593,N_13114);
nor U17695 (N_17695,N_13866,N_13026);
xor U17696 (N_17696,N_13768,N_13130);
nand U17697 (N_17697,N_12996,N_15362);
nand U17698 (N_17698,N_13236,N_13801);
and U17699 (N_17699,N_12603,N_13973);
nor U17700 (N_17700,N_13000,N_13472);
nand U17701 (N_17701,N_12516,N_14079);
nor U17702 (N_17702,N_13248,N_14261);
nor U17703 (N_17703,N_15348,N_15001);
and U17704 (N_17704,N_14614,N_15305);
nand U17705 (N_17705,N_12714,N_13685);
or U17706 (N_17706,N_15088,N_13771);
and U17707 (N_17707,N_13444,N_14531);
or U17708 (N_17708,N_13364,N_15202);
and U17709 (N_17709,N_13326,N_14835);
nand U17710 (N_17710,N_14167,N_15414);
or U17711 (N_17711,N_14974,N_13620);
nor U17712 (N_17712,N_13851,N_13545);
or U17713 (N_17713,N_12926,N_14776);
or U17714 (N_17714,N_15414,N_13724);
or U17715 (N_17715,N_15589,N_15235);
and U17716 (N_17716,N_14390,N_13528);
xor U17717 (N_17717,N_12728,N_15290);
xnor U17718 (N_17718,N_15101,N_13326);
nand U17719 (N_17719,N_14483,N_13760);
xnor U17720 (N_17720,N_15228,N_15255);
nor U17721 (N_17721,N_15207,N_12717);
xor U17722 (N_17722,N_14691,N_13678);
nand U17723 (N_17723,N_13545,N_14315);
and U17724 (N_17724,N_15431,N_14948);
or U17725 (N_17725,N_12787,N_15178);
and U17726 (N_17726,N_13122,N_14373);
nor U17727 (N_17727,N_14770,N_15534);
nor U17728 (N_17728,N_13966,N_13380);
nand U17729 (N_17729,N_12911,N_13260);
xor U17730 (N_17730,N_13305,N_15312);
xor U17731 (N_17731,N_15030,N_12681);
nand U17732 (N_17732,N_14740,N_14130);
or U17733 (N_17733,N_14275,N_14863);
xor U17734 (N_17734,N_14787,N_15017);
nor U17735 (N_17735,N_12998,N_13025);
nand U17736 (N_17736,N_14359,N_12645);
nand U17737 (N_17737,N_12501,N_13960);
and U17738 (N_17738,N_14176,N_15366);
nor U17739 (N_17739,N_13119,N_14152);
nand U17740 (N_17740,N_15138,N_13433);
nor U17741 (N_17741,N_13853,N_14583);
xor U17742 (N_17742,N_13716,N_14532);
or U17743 (N_17743,N_15324,N_14469);
and U17744 (N_17744,N_12906,N_12805);
nand U17745 (N_17745,N_12754,N_15201);
or U17746 (N_17746,N_14891,N_13335);
nor U17747 (N_17747,N_15164,N_12527);
xnor U17748 (N_17748,N_14163,N_13726);
xnor U17749 (N_17749,N_14372,N_15373);
xnor U17750 (N_17750,N_14296,N_12707);
nor U17751 (N_17751,N_13541,N_12926);
nand U17752 (N_17752,N_14169,N_14739);
xnor U17753 (N_17753,N_14185,N_14177);
xor U17754 (N_17754,N_12843,N_12762);
xnor U17755 (N_17755,N_13037,N_14382);
or U17756 (N_17756,N_14456,N_15590);
or U17757 (N_17757,N_14799,N_14834);
or U17758 (N_17758,N_15136,N_13403);
and U17759 (N_17759,N_14947,N_13858);
xor U17760 (N_17760,N_15017,N_13332);
nor U17761 (N_17761,N_12589,N_13492);
nor U17762 (N_17762,N_12700,N_13144);
or U17763 (N_17763,N_13066,N_13811);
xnor U17764 (N_17764,N_13187,N_15131);
or U17765 (N_17765,N_14818,N_15609);
or U17766 (N_17766,N_14554,N_15617);
or U17767 (N_17767,N_13616,N_13476);
xor U17768 (N_17768,N_15270,N_13106);
nor U17769 (N_17769,N_15189,N_14308);
and U17770 (N_17770,N_12793,N_13682);
nor U17771 (N_17771,N_13573,N_13404);
nand U17772 (N_17772,N_12661,N_15608);
nand U17773 (N_17773,N_15202,N_14137);
xor U17774 (N_17774,N_15535,N_12516);
or U17775 (N_17775,N_15291,N_13192);
nand U17776 (N_17776,N_14722,N_15369);
nand U17777 (N_17777,N_14602,N_12716);
or U17778 (N_17778,N_12910,N_13246);
nor U17779 (N_17779,N_15502,N_13652);
xor U17780 (N_17780,N_14251,N_13961);
nand U17781 (N_17781,N_12848,N_12998);
or U17782 (N_17782,N_14910,N_12798);
and U17783 (N_17783,N_15224,N_12535);
or U17784 (N_17784,N_13867,N_15205);
nand U17785 (N_17785,N_14816,N_14745);
or U17786 (N_17786,N_12726,N_14323);
and U17787 (N_17787,N_14693,N_14098);
and U17788 (N_17788,N_15155,N_14577);
xor U17789 (N_17789,N_13160,N_12679);
nand U17790 (N_17790,N_14832,N_15073);
nand U17791 (N_17791,N_13530,N_14233);
nor U17792 (N_17792,N_12905,N_12792);
nor U17793 (N_17793,N_13763,N_14595);
nor U17794 (N_17794,N_13657,N_14956);
nor U17795 (N_17795,N_13882,N_13228);
xor U17796 (N_17796,N_15293,N_14736);
nor U17797 (N_17797,N_14096,N_13911);
or U17798 (N_17798,N_15016,N_14487);
xor U17799 (N_17799,N_15265,N_13082);
and U17800 (N_17800,N_14460,N_15527);
or U17801 (N_17801,N_12604,N_15456);
or U17802 (N_17802,N_13946,N_14570);
or U17803 (N_17803,N_13095,N_15456);
nor U17804 (N_17804,N_15557,N_14354);
or U17805 (N_17805,N_13501,N_12890);
and U17806 (N_17806,N_15307,N_14675);
nand U17807 (N_17807,N_13001,N_13221);
and U17808 (N_17808,N_12514,N_14088);
or U17809 (N_17809,N_12596,N_14829);
and U17810 (N_17810,N_15175,N_15622);
and U17811 (N_17811,N_15309,N_13837);
nor U17812 (N_17812,N_15348,N_13401);
nor U17813 (N_17813,N_13940,N_13685);
nand U17814 (N_17814,N_13685,N_12578);
and U17815 (N_17815,N_15546,N_14147);
xnor U17816 (N_17816,N_13058,N_13806);
xnor U17817 (N_17817,N_13663,N_14281);
nor U17818 (N_17818,N_14863,N_13585);
and U17819 (N_17819,N_14938,N_12736);
xor U17820 (N_17820,N_13126,N_14486);
nand U17821 (N_17821,N_15382,N_13745);
nor U17822 (N_17822,N_13181,N_14869);
nor U17823 (N_17823,N_15494,N_14774);
nor U17824 (N_17824,N_14546,N_13158);
xor U17825 (N_17825,N_14356,N_14186);
and U17826 (N_17826,N_12962,N_15394);
and U17827 (N_17827,N_12737,N_15088);
nor U17828 (N_17828,N_12646,N_13409);
or U17829 (N_17829,N_14964,N_14631);
or U17830 (N_17830,N_13369,N_15589);
or U17831 (N_17831,N_14395,N_12608);
xor U17832 (N_17832,N_15125,N_15412);
nor U17833 (N_17833,N_13812,N_14178);
or U17834 (N_17834,N_12610,N_14194);
nor U17835 (N_17835,N_13626,N_14345);
nor U17836 (N_17836,N_13093,N_13290);
or U17837 (N_17837,N_13017,N_14907);
nand U17838 (N_17838,N_13373,N_13129);
nand U17839 (N_17839,N_14573,N_12542);
nand U17840 (N_17840,N_13358,N_14988);
nor U17841 (N_17841,N_13221,N_14415);
nand U17842 (N_17842,N_12661,N_15342);
or U17843 (N_17843,N_14061,N_14026);
nor U17844 (N_17844,N_13071,N_14295);
nand U17845 (N_17845,N_13254,N_15290);
or U17846 (N_17846,N_15563,N_12566);
xor U17847 (N_17847,N_12740,N_15474);
or U17848 (N_17848,N_13846,N_13264);
and U17849 (N_17849,N_12693,N_15621);
and U17850 (N_17850,N_13017,N_14371);
and U17851 (N_17851,N_14783,N_12982);
nor U17852 (N_17852,N_13287,N_12619);
or U17853 (N_17853,N_14912,N_12796);
nor U17854 (N_17854,N_13402,N_15366);
xor U17855 (N_17855,N_15178,N_14050);
and U17856 (N_17856,N_15136,N_14155);
and U17857 (N_17857,N_13173,N_13859);
nand U17858 (N_17858,N_14159,N_14462);
xor U17859 (N_17859,N_15601,N_12851);
or U17860 (N_17860,N_15573,N_14386);
nor U17861 (N_17861,N_15374,N_15566);
nor U17862 (N_17862,N_13907,N_12516);
nand U17863 (N_17863,N_15043,N_12976);
nand U17864 (N_17864,N_13135,N_14290);
and U17865 (N_17865,N_13578,N_14860);
nor U17866 (N_17866,N_14940,N_15054);
nor U17867 (N_17867,N_15597,N_15476);
nor U17868 (N_17868,N_15066,N_14220);
xor U17869 (N_17869,N_13046,N_14590);
nor U17870 (N_17870,N_14796,N_14758);
and U17871 (N_17871,N_13419,N_14100);
xnor U17872 (N_17872,N_12727,N_13227);
or U17873 (N_17873,N_14027,N_14943);
and U17874 (N_17874,N_13268,N_12911);
nand U17875 (N_17875,N_15226,N_13869);
xnor U17876 (N_17876,N_13524,N_14128);
or U17877 (N_17877,N_12731,N_12863);
nor U17878 (N_17878,N_13942,N_15619);
nor U17879 (N_17879,N_15059,N_13490);
and U17880 (N_17880,N_14984,N_15103);
nand U17881 (N_17881,N_14074,N_14341);
nor U17882 (N_17882,N_13928,N_15400);
nor U17883 (N_17883,N_12623,N_12606);
nand U17884 (N_17884,N_15198,N_15536);
nand U17885 (N_17885,N_13126,N_14199);
nand U17886 (N_17886,N_13356,N_13646);
nor U17887 (N_17887,N_14004,N_13539);
or U17888 (N_17888,N_13406,N_12832);
nand U17889 (N_17889,N_15331,N_14621);
or U17890 (N_17890,N_13070,N_12832);
or U17891 (N_17891,N_13506,N_13779);
nor U17892 (N_17892,N_12550,N_15509);
xnor U17893 (N_17893,N_13373,N_13663);
nand U17894 (N_17894,N_13377,N_14343);
or U17895 (N_17895,N_14363,N_14964);
xnor U17896 (N_17896,N_15188,N_12634);
nand U17897 (N_17897,N_15314,N_15080);
and U17898 (N_17898,N_15432,N_14699);
nor U17899 (N_17899,N_15540,N_12900);
xor U17900 (N_17900,N_14423,N_13380);
and U17901 (N_17901,N_15259,N_13735);
or U17902 (N_17902,N_15024,N_13752);
nor U17903 (N_17903,N_13072,N_15297);
and U17904 (N_17904,N_13994,N_12603);
and U17905 (N_17905,N_14550,N_13104);
xnor U17906 (N_17906,N_15179,N_14704);
xnor U17907 (N_17907,N_13677,N_12947);
and U17908 (N_17908,N_15610,N_14119);
nand U17909 (N_17909,N_13783,N_12529);
xnor U17910 (N_17910,N_14605,N_13312);
or U17911 (N_17911,N_15464,N_14796);
nor U17912 (N_17912,N_14319,N_12810);
nor U17913 (N_17913,N_12752,N_13900);
or U17914 (N_17914,N_12759,N_12951);
nor U17915 (N_17915,N_13363,N_14324);
xor U17916 (N_17916,N_13888,N_13683);
and U17917 (N_17917,N_14272,N_13630);
and U17918 (N_17918,N_15510,N_12831);
and U17919 (N_17919,N_15159,N_15463);
nand U17920 (N_17920,N_15571,N_12797);
or U17921 (N_17921,N_13998,N_12966);
and U17922 (N_17922,N_13126,N_13562);
and U17923 (N_17923,N_12980,N_12828);
or U17924 (N_17924,N_12738,N_14012);
or U17925 (N_17925,N_13827,N_13330);
nor U17926 (N_17926,N_13558,N_13331);
nand U17927 (N_17927,N_13477,N_15499);
nand U17928 (N_17928,N_14362,N_13716);
nand U17929 (N_17929,N_15517,N_13994);
xor U17930 (N_17930,N_15214,N_12934);
or U17931 (N_17931,N_14924,N_12593);
xnor U17932 (N_17932,N_15111,N_13159);
and U17933 (N_17933,N_13005,N_13968);
or U17934 (N_17934,N_13189,N_13105);
or U17935 (N_17935,N_13974,N_13430);
and U17936 (N_17936,N_13142,N_12602);
xor U17937 (N_17937,N_14153,N_15089);
and U17938 (N_17938,N_14835,N_12644);
xnor U17939 (N_17939,N_15245,N_15209);
or U17940 (N_17940,N_13228,N_13855);
xor U17941 (N_17941,N_13551,N_15294);
nor U17942 (N_17942,N_14716,N_15497);
and U17943 (N_17943,N_13276,N_13435);
and U17944 (N_17944,N_12666,N_14734);
nor U17945 (N_17945,N_15414,N_13028);
and U17946 (N_17946,N_15193,N_13087);
and U17947 (N_17947,N_14388,N_12913);
xor U17948 (N_17948,N_12634,N_14651);
and U17949 (N_17949,N_15275,N_14959);
and U17950 (N_17950,N_15136,N_13601);
and U17951 (N_17951,N_13831,N_12928);
xnor U17952 (N_17952,N_12713,N_15575);
xnor U17953 (N_17953,N_15264,N_14108);
nand U17954 (N_17954,N_13834,N_13341);
nor U17955 (N_17955,N_15398,N_13097);
or U17956 (N_17956,N_14132,N_14742);
nand U17957 (N_17957,N_13227,N_12586);
nand U17958 (N_17958,N_15360,N_14390);
nor U17959 (N_17959,N_14994,N_13196);
nor U17960 (N_17960,N_12999,N_13038);
nand U17961 (N_17961,N_13718,N_12533);
and U17962 (N_17962,N_14692,N_14555);
nand U17963 (N_17963,N_15441,N_14740);
nand U17964 (N_17964,N_14224,N_13847);
or U17965 (N_17965,N_13997,N_14580);
nand U17966 (N_17966,N_12920,N_14821);
xnor U17967 (N_17967,N_15398,N_14845);
xor U17968 (N_17968,N_14330,N_13099);
nand U17969 (N_17969,N_13361,N_15341);
nand U17970 (N_17970,N_13717,N_13008);
xnor U17971 (N_17971,N_15594,N_14009);
nor U17972 (N_17972,N_14086,N_12571);
or U17973 (N_17973,N_14946,N_15313);
xnor U17974 (N_17974,N_13158,N_14358);
and U17975 (N_17975,N_12631,N_15489);
or U17976 (N_17976,N_12993,N_13771);
or U17977 (N_17977,N_14598,N_14094);
and U17978 (N_17978,N_14826,N_14198);
nand U17979 (N_17979,N_12960,N_15314);
and U17980 (N_17980,N_13328,N_13802);
or U17981 (N_17981,N_13839,N_13670);
or U17982 (N_17982,N_13936,N_15575);
and U17983 (N_17983,N_15108,N_15525);
and U17984 (N_17984,N_13008,N_14881);
or U17985 (N_17985,N_14787,N_13513);
or U17986 (N_17986,N_13185,N_14920);
xnor U17987 (N_17987,N_13878,N_12565);
nand U17988 (N_17988,N_12829,N_15000);
xor U17989 (N_17989,N_14013,N_14060);
and U17990 (N_17990,N_15411,N_15386);
xnor U17991 (N_17991,N_13576,N_14558);
nor U17992 (N_17992,N_13668,N_12545);
nor U17993 (N_17993,N_13822,N_14616);
and U17994 (N_17994,N_13173,N_12823);
or U17995 (N_17995,N_12848,N_13797);
and U17996 (N_17996,N_13648,N_14449);
and U17997 (N_17997,N_13839,N_13649);
xor U17998 (N_17998,N_15599,N_13658);
and U17999 (N_17999,N_13734,N_14977);
nor U18000 (N_18000,N_14066,N_13536);
and U18001 (N_18001,N_14005,N_14137);
xnor U18002 (N_18002,N_12585,N_15085);
or U18003 (N_18003,N_13355,N_13488);
xor U18004 (N_18004,N_14317,N_13751);
nor U18005 (N_18005,N_14089,N_13668);
xnor U18006 (N_18006,N_15239,N_15523);
and U18007 (N_18007,N_13792,N_12677);
nor U18008 (N_18008,N_12609,N_14556);
nor U18009 (N_18009,N_14503,N_13875);
and U18010 (N_18010,N_13599,N_12984);
and U18011 (N_18011,N_12876,N_14843);
nand U18012 (N_18012,N_12638,N_14913);
and U18013 (N_18013,N_13629,N_14478);
or U18014 (N_18014,N_15457,N_14384);
nor U18015 (N_18015,N_13543,N_15081);
nand U18016 (N_18016,N_14983,N_13380);
or U18017 (N_18017,N_15439,N_14222);
xnor U18018 (N_18018,N_13707,N_14366);
nor U18019 (N_18019,N_13964,N_12552);
or U18020 (N_18020,N_13500,N_14782);
xnor U18021 (N_18021,N_14688,N_14280);
nand U18022 (N_18022,N_14525,N_12570);
and U18023 (N_18023,N_13186,N_13339);
and U18024 (N_18024,N_13873,N_13916);
and U18025 (N_18025,N_13316,N_13635);
and U18026 (N_18026,N_15195,N_13932);
or U18027 (N_18027,N_15341,N_12992);
nor U18028 (N_18028,N_14670,N_15453);
or U18029 (N_18029,N_13052,N_12624);
nand U18030 (N_18030,N_13222,N_14312);
xnor U18031 (N_18031,N_14094,N_14044);
nor U18032 (N_18032,N_15624,N_14281);
nor U18033 (N_18033,N_14727,N_13267);
or U18034 (N_18034,N_14037,N_15408);
xor U18035 (N_18035,N_15616,N_15004);
or U18036 (N_18036,N_14236,N_13695);
nand U18037 (N_18037,N_14675,N_13035);
nand U18038 (N_18038,N_14503,N_15449);
and U18039 (N_18039,N_14677,N_13833);
xnor U18040 (N_18040,N_14118,N_15324);
nor U18041 (N_18041,N_14403,N_12926);
nand U18042 (N_18042,N_13307,N_13185);
or U18043 (N_18043,N_15606,N_13766);
xor U18044 (N_18044,N_14977,N_14502);
nor U18045 (N_18045,N_15014,N_14113);
nor U18046 (N_18046,N_13342,N_14874);
or U18047 (N_18047,N_13282,N_13963);
nand U18048 (N_18048,N_13106,N_12929);
and U18049 (N_18049,N_14809,N_14648);
and U18050 (N_18050,N_14980,N_13363);
nor U18051 (N_18051,N_14839,N_13119);
nor U18052 (N_18052,N_12761,N_14018);
xor U18053 (N_18053,N_13828,N_14701);
nor U18054 (N_18054,N_14156,N_15379);
or U18055 (N_18055,N_12868,N_14817);
nor U18056 (N_18056,N_12731,N_12821);
nand U18057 (N_18057,N_13931,N_14519);
or U18058 (N_18058,N_12840,N_12803);
nor U18059 (N_18059,N_12631,N_13587);
nand U18060 (N_18060,N_15249,N_13257);
and U18061 (N_18061,N_14858,N_15553);
nand U18062 (N_18062,N_12995,N_12502);
nand U18063 (N_18063,N_13762,N_12557);
xor U18064 (N_18064,N_15254,N_14522);
or U18065 (N_18065,N_14480,N_14672);
nand U18066 (N_18066,N_14425,N_13592);
nor U18067 (N_18067,N_12506,N_13446);
xnor U18068 (N_18068,N_12998,N_15028);
nand U18069 (N_18069,N_12550,N_13838);
and U18070 (N_18070,N_14057,N_14681);
nand U18071 (N_18071,N_14177,N_12883);
or U18072 (N_18072,N_15140,N_12778);
xnor U18073 (N_18073,N_13758,N_13949);
xor U18074 (N_18074,N_13150,N_14348);
nand U18075 (N_18075,N_15064,N_13972);
or U18076 (N_18076,N_15408,N_13846);
xor U18077 (N_18077,N_14388,N_15021);
xor U18078 (N_18078,N_14625,N_14922);
or U18079 (N_18079,N_14314,N_13436);
nor U18080 (N_18080,N_15190,N_12635);
xnor U18081 (N_18081,N_13103,N_13960);
nand U18082 (N_18082,N_13240,N_15350);
nor U18083 (N_18083,N_13929,N_12878);
and U18084 (N_18084,N_13479,N_14285);
and U18085 (N_18085,N_13046,N_15268);
xor U18086 (N_18086,N_13466,N_12724);
xnor U18087 (N_18087,N_15602,N_15431);
nand U18088 (N_18088,N_14902,N_13662);
nor U18089 (N_18089,N_14402,N_13974);
and U18090 (N_18090,N_15386,N_15537);
xor U18091 (N_18091,N_14275,N_14787);
or U18092 (N_18092,N_15520,N_12852);
or U18093 (N_18093,N_13273,N_15554);
or U18094 (N_18094,N_13197,N_15049);
or U18095 (N_18095,N_13273,N_14623);
nor U18096 (N_18096,N_14906,N_13144);
nor U18097 (N_18097,N_13183,N_14570);
nor U18098 (N_18098,N_13695,N_14697);
and U18099 (N_18099,N_15623,N_14369);
nand U18100 (N_18100,N_14204,N_13252);
or U18101 (N_18101,N_13102,N_12525);
and U18102 (N_18102,N_13618,N_15606);
or U18103 (N_18103,N_15084,N_12664);
and U18104 (N_18104,N_15504,N_13527);
nand U18105 (N_18105,N_13871,N_13555);
nand U18106 (N_18106,N_14769,N_13778);
nand U18107 (N_18107,N_14390,N_15222);
nor U18108 (N_18108,N_14156,N_15363);
nand U18109 (N_18109,N_14759,N_13132);
nand U18110 (N_18110,N_12511,N_14438);
or U18111 (N_18111,N_15350,N_14243);
xor U18112 (N_18112,N_13033,N_14107);
and U18113 (N_18113,N_15482,N_12505);
xnor U18114 (N_18114,N_14388,N_15526);
nand U18115 (N_18115,N_12519,N_14932);
xor U18116 (N_18116,N_12792,N_12639);
nand U18117 (N_18117,N_13647,N_15599);
nand U18118 (N_18118,N_15048,N_13042);
nand U18119 (N_18119,N_15272,N_14302);
and U18120 (N_18120,N_13034,N_15203);
nor U18121 (N_18121,N_13125,N_12782);
or U18122 (N_18122,N_14023,N_12819);
and U18123 (N_18123,N_15313,N_14251);
and U18124 (N_18124,N_14727,N_14077);
or U18125 (N_18125,N_13135,N_15587);
or U18126 (N_18126,N_15262,N_14373);
nand U18127 (N_18127,N_15560,N_12660);
nand U18128 (N_18128,N_13438,N_15474);
or U18129 (N_18129,N_13667,N_14300);
or U18130 (N_18130,N_12729,N_13601);
nand U18131 (N_18131,N_14635,N_14880);
and U18132 (N_18132,N_14037,N_12735);
and U18133 (N_18133,N_15597,N_15614);
xnor U18134 (N_18134,N_14092,N_14210);
and U18135 (N_18135,N_13721,N_14514);
nor U18136 (N_18136,N_14154,N_13598);
nor U18137 (N_18137,N_12826,N_15151);
nand U18138 (N_18138,N_13379,N_14137);
nor U18139 (N_18139,N_15307,N_13682);
nand U18140 (N_18140,N_13557,N_12823);
and U18141 (N_18141,N_15273,N_14818);
nand U18142 (N_18142,N_15324,N_12979);
nand U18143 (N_18143,N_13145,N_14783);
nand U18144 (N_18144,N_15280,N_12899);
and U18145 (N_18145,N_12947,N_15365);
nor U18146 (N_18146,N_12713,N_13477);
nand U18147 (N_18147,N_13856,N_12637);
and U18148 (N_18148,N_14513,N_15463);
or U18149 (N_18149,N_13484,N_13074);
nor U18150 (N_18150,N_13864,N_14464);
and U18151 (N_18151,N_14153,N_13436);
or U18152 (N_18152,N_15515,N_13179);
nand U18153 (N_18153,N_12939,N_15005);
nand U18154 (N_18154,N_15408,N_15570);
nand U18155 (N_18155,N_13399,N_14766);
or U18156 (N_18156,N_15112,N_12952);
xor U18157 (N_18157,N_14022,N_14580);
xnor U18158 (N_18158,N_14817,N_12843);
xnor U18159 (N_18159,N_13163,N_14340);
nand U18160 (N_18160,N_13958,N_13944);
xor U18161 (N_18161,N_12891,N_13295);
and U18162 (N_18162,N_12705,N_12517);
nor U18163 (N_18163,N_12558,N_14948);
xor U18164 (N_18164,N_15260,N_13926);
nand U18165 (N_18165,N_13350,N_14213);
or U18166 (N_18166,N_15065,N_13304);
or U18167 (N_18167,N_12988,N_13776);
nor U18168 (N_18168,N_13709,N_14734);
nand U18169 (N_18169,N_12702,N_13159);
and U18170 (N_18170,N_14103,N_14847);
nand U18171 (N_18171,N_14834,N_13122);
and U18172 (N_18172,N_14827,N_13653);
xnor U18173 (N_18173,N_13995,N_12908);
and U18174 (N_18174,N_13442,N_14773);
nor U18175 (N_18175,N_15473,N_13160);
and U18176 (N_18176,N_14750,N_14621);
nand U18177 (N_18177,N_13164,N_13421);
nor U18178 (N_18178,N_13015,N_13531);
xor U18179 (N_18179,N_15124,N_12745);
and U18180 (N_18180,N_14089,N_14062);
xor U18181 (N_18181,N_12681,N_12898);
nor U18182 (N_18182,N_12516,N_13022);
or U18183 (N_18183,N_12984,N_13447);
nand U18184 (N_18184,N_14379,N_12539);
and U18185 (N_18185,N_15300,N_13173);
nand U18186 (N_18186,N_13854,N_14790);
and U18187 (N_18187,N_12615,N_15078);
xnor U18188 (N_18188,N_13163,N_15007);
nor U18189 (N_18189,N_12757,N_14124);
nand U18190 (N_18190,N_13456,N_14084);
and U18191 (N_18191,N_15495,N_15084);
and U18192 (N_18192,N_12731,N_14428);
or U18193 (N_18193,N_12822,N_15471);
or U18194 (N_18194,N_13715,N_14678);
and U18195 (N_18195,N_12979,N_14582);
nor U18196 (N_18196,N_13471,N_13109);
nand U18197 (N_18197,N_14622,N_14139);
nand U18198 (N_18198,N_13618,N_14192);
nand U18199 (N_18199,N_15260,N_13647);
nand U18200 (N_18200,N_15468,N_13427);
nand U18201 (N_18201,N_15576,N_13878);
xnor U18202 (N_18202,N_13823,N_13319);
xnor U18203 (N_18203,N_12505,N_12838);
xor U18204 (N_18204,N_14332,N_13810);
nand U18205 (N_18205,N_12771,N_13412);
or U18206 (N_18206,N_14221,N_14432);
and U18207 (N_18207,N_13353,N_15496);
nor U18208 (N_18208,N_13434,N_13721);
and U18209 (N_18209,N_14440,N_13899);
or U18210 (N_18210,N_12949,N_15027);
nor U18211 (N_18211,N_14901,N_15175);
and U18212 (N_18212,N_13856,N_12868);
and U18213 (N_18213,N_13489,N_12676);
nor U18214 (N_18214,N_12663,N_15097);
and U18215 (N_18215,N_14983,N_13488);
nand U18216 (N_18216,N_15038,N_12638);
xor U18217 (N_18217,N_15355,N_15177);
nand U18218 (N_18218,N_13880,N_14777);
nand U18219 (N_18219,N_14371,N_13075);
nor U18220 (N_18220,N_12923,N_12820);
nand U18221 (N_18221,N_13087,N_13527);
nand U18222 (N_18222,N_13612,N_14524);
or U18223 (N_18223,N_13674,N_13819);
or U18224 (N_18224,N_14437,N_14291);
or U18225 (N_18225,N_14822,N_13002);
nand U18226 (N_18226,N_13379,N_15318);
nand U18227 (N_18227,N_12602,N_13225);
and U18228 (N_18228,N_13193,N_15282);
and U18229 (N_18229,N_15251,N_14063);
or U18230 (N_18230,N_14267,N_14178);
nor U18231 (N_18231,N_15368,N_13149);
and U18232 (N_18232,N_14231,N_12931);
nand U18233 (N_18233,N_13736,N_12763);
nand U18234 (N_18234,N_13050,N_14944);
xor U18235 (N_18235,N_12532,N_14426);
nand U18236 (N_18236,N_13051,N_12739);
or U18237 (N_18237,N_14540,N_13011);
xor U18238 (N_18238,N_13671,N_15463);
or U18239 (N_18239,N_13263,N_15162);
nand U18240 (N_18240,N_14802,N_13030);
and U18241 (N_18241,N_12520,N_12868);
xnor U18242 (N_18242,N_14994,N_13389);
or U18243 (N_18243,N_13410,N_13534);
or U18244 (N_18244,N_14773,N_13915);
nand U18245 (N_18245,N_13511,N_13211);
nor U18246 (N_18246,N_13785,N_12920);
and U18247 (N_18247,N_13788,N_14873);
or U18248 (N_18248,N_14978,N_15167);
xor U18249 (N_18249,N_14883,N_14776);
xnor U18250 (N_18250,N_13561,N_14859);
xor U18251 (N_18251,N_13359,N_14724);
or U18252 (N_18252,N_15453,N_13323);
nor U18253 (N_18253,N_15419,N_15110);
and U18254 (N_18254,N_13392,N_13758);
or U18255 (N_18255,N_15582,N_12992);
nand U18256 (N_18256,N_15271,N_14853);
or U18257 (N_18257,N_15099,N_14635);
or U18258 (N_18258,N_13940,N_15485);
xnor U18259 (N_18259,N_14884,N_13617);
nand U18260 (N_18260,N_14239,N_13813);
nand U18261 (N_18261,N_15380,N_14622);
nand U18262 (N_18262,N_13828,N_15138);
and U18263 (N_18263,N_14533,N_15443);
or U18264 (N_18264,N_13266,N_15581);
xor U18265 (N_18265,N_12992,N_14760);
or U18266 (N_18266,N_15582,N_12745);
or U18267 (N_18267,N_12952,N_13025);
nor U18268 (N_18268,N_14570,N_12749);
nor U18269 (N_18269,N_15499,N_14065);
or U18270 (N_18270,N_15222,N_13978);
and U18271 (N_18271,N_14411,N_14366);
and U18272 (N_18272,N_14985,N_14555);
nor U18273 (N_18273,N_12687,N_13347);
nor U18274 (N_18274,N_15176,N_14787);
nand U18275 (N_18275,N_13214,N_13224);
or U18276 (N_18276,N_15046,N_13790);
or U18277 (N_18277,N_14810,N_12692);
nand U18278 (N_18278,N_14642,N_14481);
nor U18279 (N_18279,N_12805,N_14989);
nor U18280 (N_18280,N_14265,N_14586);
and U18281 (N_18281,N_15544,N_15003);
and U18282 (N_18282,N_13026,N_14642);
nor U18283 (N_18283,N_12562,N_15404);
or U18284 (N_18284,N_14193,N_12846);
xnor U18285 (N_18285,N_15613,N_13008);
xnor U18286 (N_18286,N_15136,N_15118);
nor U18287 (N_18287,N_13805,N_13261);
or U18288 (N_18288,N_13511,N_13528);
or U18289 (N_18289,N_14933,N_14709);
or U18290 (N_18290,N_13039,N_13867);
and U18291 (N_18291,N_12978,N_13725);
and U18292 (N_18292,N_15054,N_13383);
nor U18293 (N_18293,N_14053,N_12502);
or U18294 (N_18294,N_13330,N_15582);
nand U18295 (N_18295,N_13012,N_12661);
nor U18296 (N_18296,N_15501,N_13829);
xnor U18297 (N_18297,N_15268,N_14120);
and U18298 (N_18298,N_14518,N_13806);
xor U18299 (N_18299,N_12688,N_14626);
and U18300 (N_18300,N_14136,N_13069);
xnor U18301 (N_18301,N_15319,N_13644);
xnor U18302 (N_18302,N_14236,N_14257);
or U18303 (N_18303,N_12999,N_15272);
and U18304 (N_18304,N_15384,N_14612);
or U18305 (N_18305,N_15420,N_13121);
nor U18306 (N_18306,N_13919,N_14761);
nand U18307 (N_18307,N_12663,N_12603);
or U18308 (N_18308,N_14134,N_12723);
and U18309 (N_18309,N_14845,N_14378);
and U18310 (N_18310,N_13525,N_13509);
nand U18311 (N_18311,N_15431,N_12594);
nor U18312 (N_18312,N_15313,N_15262);
or U18313 (N_18313,N_13818,N_12507);
nor U18314 (N_18314,N_13842,N_14438);
nor U18315 (N_18315,N_13431,N_13336);
or U18316 (N_18316,N_15451,N_12560);
xor U18317 (N_18317,N_14599,N_13212);
or U18318 (N_18318,N_13018,N_14324);
or U18319 (N_18319,N_13101,N_12642);
xor U18320 (N_18320,N_13884,N_15349);
or U18321 (N_18321,N_15608,N_13650);
and U18322 (N_18322,N_12600,N_14960);
or U18323 (N_18323,N_13147,N_14311);
nor U18324 (N_18324,N_12868,N_13585);
xor U18325 (N_18325,N_13559,N_15579);
nor U18326 (N_18326,N_15242,N_13656);
xor U18327 (N_18327,N_14912,N_13683);
and U18328 (N_18328,N_15574,N_13168);
or U18329 (N_18329,N_13767,N_13143);
nand U18330 (N_18330,N_13215,N_14006);
nand U18331 (N_18331,N_14430,N_12818);
or U18332 (N_18332,N_14723,N_14987);
nor U18333 (N_18333,N_15447,N_12971);
nor U18334 (N_18334,N_14754,N_15591);
or U18335 (N_18335,N_13165,N_15014);
nand U18336 (N_18336,N_14265,N_15250);
xnor U18337 (N_18337,N_12645,N_13073);
and U18338 (N_18338,N_14217,N_15501);
nor U18339 (N_18339,N_14030,N_14625);
xor U18340 (N_18340,N_15276,N_13846);
and U18341 (N_18341,N_13977,N_14054);
nor U18342 (N_18342,N_13760,N_14740);
and U18343 (N_18343,N_15286,N_14300);
nand U18344 (N_18344,N_14567,N_13571);
nor U18345 (N_18345,N_13290,N_13707);
nand U18346 (N_18346,N_14025,N_14576);
nor U18347 (N_18347,N_14704,N_15082);
xnor U18348 (N_18348,N_15213,N_13932);
xor U18349 (N_18349,N_13555,N_12531);
and U18350 (N_18350,N_15238,N_13798);
nor U18351 (N_18351,N_14255,N_13424);
nor U18352 (N_18352,N_13463,N_13672);
xnor U18353 (N_18353,N_13667,N_12544);
and U18354 (N_18354,N_14252,N_13615);
and U18355 (N_18355,N_12648,N_14270);
or U18356 (N_18356,N_14975,N_12809);
nor U18357 (N_18357,N_13356,N_14704);
or U18358 (N_18358,N_14640,N_15304);
or U18359 (N_18359,N_13777,N_13296);
nand U18360 (N_18360,N_15055,N_14692);
and U18361 (N_18361,N_13045,N_13144);
and U18362 (N_18362,N_14878,N_15254);
or U18363 (N_18363,N_14992,N_14210);
and U18364 (N_18364,N_13732,N_13443);
nand U18365 (N_18365,N_15097,N_14321);
and U18366 (N_18366,N_12835,N_13940);
nor U18367 (N_18367,N_13500,N_12553);
and U18368 (N_18368,N_15021,N_13254);
and U18369 (N_18369,N_13873,N_12547);
xnor U18370 (N_18370,N_13691,N_14416);
nand U18371 (N_18371,N_13710,N_13434);
xor U18372 (N_18372,N_15623,N_15128);
and U18373 (N_18373,N_14431,N_14545);
xnor U18374 (N_18374,N_14944,N_13063);
and U18375 (N_18375,N_14454,N_12651);
nand U18376 (N_18376,N_13265,N_14798);
xor U18377 (N_18377,N_13804,N_15044);
and U18378 (N_18378,N_14520,N_14378);
xnor U18379 (N_18379,N_14324,N_13231);
or U18380 (N_18380,N_14516,N_13240);
xnor U18381 (N_18381,N_14925,N_14327);
and U18382 (N_18382,N_13807,N_15069);
xnor U18383 (N_18383,N_14402,N_13541);
and U18384 (N_18384,N_12929,N_13717);
nand U18385 (N_18385,N_13246,N_13898);
or U18386 (N_18386,N_14467,N_14375);
or U18387 (N_18387,N_15244,N_15338);
nand U18388 (N_18388,N_13075,N_15329);
nand U18389 (N_18389,N_12665,N_14793);
nand U18390 (N_18390,N_13180,N_13227);
nor U18391 (N_18391,N_14061,N_14569);
or U18392 (N_18392,N_13591,N_15613);
nand U18393 (N_18393,N_15004,N_14904);
and U18394 (N_18394,N_14709,N_13517);
nand U18395 (N_18395,N_13392,N_15615);
nand U18396 (N_18396,N_13108,N_14991);
xnor U18397 (N_18397,N_12583,N_14334);
or U18398 (N_18398,N_12596,N_13078);
and U18399 (N_18399,N_15571,N_15340);
xnor U18400 (N_18400,N_14423,N_13060);
and U18401 (N_18401,N_14738,N_12607);
nand U18402 (N_18402,N_12704,N_12809);
nor U18403 (N_18403,N_13118,N_13937);
xor U18404 (N_18404,N_13306,N_13169);
xor U18405 (N_18405,N_15536,N_15261);
and U18406 (N_18406,N_12901,N_13281);
nor U18407 (N_18407,N_13556,N_14532);
nor U18408 (N_18408,N_14954,N_15339);
and U18409 (N_18409,N_14820,N_15522);
or U18410 (N_18410,N_12881,N_13242);
nor U18411 (N_18411,N_14584,N_12800);
xnor U18412 (N_18412,N_13522,N_14158);
nand U18413 (N_18413,N_13859,N_13457);
xor U18414 (N_18414,N_13543,N_13469);
and U18415 (N_18415,N_13027,N_13907);
nor U18416 (N_18416,N_13356,N_15133);
nand U18417 (N_18417,N_15335,N_15344);
nor U18418 (N_18418,N_13180,N_13073);
nor U18419 (N_18419,N_13677,N_15321);
and U18420 (N_18420,N_14737,N_15295);
nor U18421 (N_18421,N_13407,N_13040);
nand U18422 (N_18422,N_13165,N_13883);
nand U18423 (N_18423,N_14770,N_15547);
nand U18424 (N_18424,N_13099,N_13554);
xor U18425 (N_18425,N_13923,N_15031);
or U18426 (N_18426,N_13326,N_15024);
xor U18427 (N_18427,N_15385,N_14522);
and U18428 (N_18428,N_12888,N_14212);
xnor U18429 (N_18429,N_14841,N_14086);
or U18430 (N_18430,N_12989,N_13751);
nand U18431 (N_18431,N_13826,N_13618);
nand U18432 (N_18432,N_12908,N_14248);
nor U18433 (N_18433,N_13156,N_14369);
nor U18434 (N_18434,N_15477,N_13978);
xor U18435 (N_18435,N_14895,N_13399);
or U18436 (N_18436,N_13609,N_12558);
xor U18437 (N_18437,N_14065,N_14576);
and U18438 (N_18438,N_13679,N_14332);
and U18439 (N_18439,N_13132,N_12643);
and U18440 (N_18440,N_13832,N_15430);
xnor U18441 (N_18441,N_13246,N_14011);
nand U18442 (N_18442,N_15482,N_14877);
nor U18443 (N_18443,N_14850,N_14725);
and U18444 (N_18444,N_15412,N_14873);
and U18445 (N_18445,N_14524,N_14225);
and U18446 (N_18446,N_14513,N_15008);
or U18447 (N_18447,N_14858,N_14468);
or U18448 (N_18448,N_14101,N_14240);
xor U18449 (N_18449,N_12921,N_14304);
or U18450 (N_18450,N_13883,N_12885);
nor U18451 (N_18451,N_13511,N_13131);
xnor U18452 (N_18452,N_13304,N_12843);
xnor U18453 (N_18453,N_13900,N_12572);
nor U18454 (N_18454,N_13000,N_15477);
nand U18455 (N_18455,N_14509,N_14133);
xor U18456 (N_18456,N_12905,N_14500);
nor U18457 (N_18457,N_15534,N_15061);
nor U18458 (N_18458,N_15305,N_14230);
xor U18459 (N_18459,N_15153,N_14459);
nand U18460 (N_18460,N_13286,N_15486);
and U18461 (N_18461,N_15300,N_14126);
nand U18462 (N_18462,N_14802,N_15067);
or U18463 (N_18463,N_15211,N_15291);
nor U18464 (N_18464,N_14589,N_13483);
and U18465 (N_18465,N_12827,N_13463);
or U18466 (N_18466,N_14814,N_12732);
nor U18467 (N_18467,N_15188,N_12611);
or U18468 (N_18468,N_12927,N_12611);
nand U18469 (N_18469,N_14391,N_14224);
or U18470 (N_18470,N_13639,N_12905);
xnor U18471 (N_18471,N_13911,N_15179);
xnor U18472 (N_18472,N_13421,N_13641);
and U18473 (N_18473,N_14305,N_14969);
nor U18474 (N_18474,N_13393,N_15538);
or U18475 (N_18475,N_13643,N_12997);
nor U18476 (N_18476,N_12505,N_15208);
nor U18477 (N_18477,N_14461,N_12638);
and U18478 (N_18478,N_13881,N_14266);
and U18479 (N_18479,N_13607,N_13493);
nand U18480 (N_18480,N_15560,N_14542);
nand U18481 (N_18481,N_14574,N_12767);
or U18482 (N_18482,N_14183,N_14754);
and U18483 (N_18483,N_14555,N_13947);
xnor U18484 (N_18484,N_14786,N_12894);
nor U18485 (N_18485,N_14573,N_14115);
and U18486 (N_18486,N_14249,N_15245);
and U18487 (N_18487,N_14684,N_14750);
nor U18488 (N_18488,N_14757,N_14094);
nor U18489 (N_18489,N_14325,N_13200);
nand U18490 (N_18490,N_14710,N_12779);
nor U18491 (N_18491,N_13454,N_13104);
nor U18492 (N_18492,N_13554,N_15427);
or U18493 (N_18493,N_13253,N_12830);
and U18494 (N_18494,N_13965,N_14828);
and U18495 (N_18495,N_15099,N_15548);
xor U18496 (N_18496,N_14784,N_14676);
nand U18497 (N_18497,N_12847,N_13774);
nor U18498 (N_18498,N_15604,N_13616);
xor U18499 (N_18499,N_14941,N_12719);
xor U18500 (N_18500,N_13258,N_15490);
or U18501 (N_18501,N_12660,N_14746);
and U18502 (N_18502,N_13548,N_14058);
nor U18503 (N_18503,N_15079,N_13355);
nor U18504 (N_18504,N_13480,N_13746);
xnor U18505 (N_18505,N_14579,N_13801);
or U18506 (N_18506,N_15310,N_12502);
or U18507 (N_18507,N_14660,N_15320);
xnor U18508 (N_18508,N_12858,N_13096);
xnor U18509 (N_18509,N_13287,N_14836);
and U18510 (N_18510,N_12586,N_12532);
xor U18511 (N_18511,N_14888,N_14245);
nand U18512 (N_18512,N_14911,N_15029);
nor U18513 (N_18513,N_12642,N_13009);
and U18514 (N_18514,N_12752,N_14025);
xnor U18515 (N_18515,N_15247,N_15145);
nand U18516 (N_18516,N_12792,N_13174);
xor U18517 (N_18517,N_13475,N_12754);
nand U18518 (N_18518,N_15310,N_15559);
and U18519 (N_18519,N_13129,N_14986);
xnor U18520 (N_18520,N_12720,N_15117);
nand U18521 (N_18521,N_14483,N_15534);
nand U18522 (N_18522,N_15400,N_13151);
nor U18523 (N_18523,N_13387,N_13461);
and U18524 (N_18524,N_15112,N_14373);
nand U18525 (N_18525,N_14265,N_13384);
and U18526 (N_18526,N_15112,N_13868);
xor U18527 (N_18527,N_12788,N_13003);
nand U18528 (N_18528,N_14734,N_14630);
nor U18529 (N_18529,N_15230,N_14529);
nor U18530 (N_18530,N_15576,N_14804);
xnor U18531 (N_18531,N_15229,N_14379);
or U18532 (N_18532,N_13069,N_13383);
and U18533 (N_18533,N_15173,N_13041);
or U18534 (N_18534,N_14183,N_13897);
nor U18535 (N_18535,N_13368,N_12972);
or U18536 (N_18536,N_14656,N_13603);
or U18537 (N_18537,N_15189,N_12945);
or U18538 (N_18538,N_14062,N_12790);
nand U18539 (N_18539,N_14151,N_14508);
or U18540 (N_18540,N_15377,N_13018);
and U18541 (N_18541,N_12843,N_14944);
or U18542 (N_18542,N_12959,N_13731);
or U18543 (N_18543,N_14940,N_14288);
and U18544 (N_18544,N_14892,N_14917);
and U18545 (N_18545,N_14013,N_14146);
xor U18546 (N_18546,N_12689,N_14525);
and U18547 (N_18547,N_14500,N_15505);
nand U18548 (N_18548,N_13145,N_15052);
and U18549 (N_18549,N_12514,N_13635);
or U18550 (N_18550,N_15611,N_13748);
nand U18551 (N_18551,N_14526,N_13063);
nand U18552 (N_18552,N_13688,N_12604);
nand U18553 (N_18553,N_13618,N_15396);
or U18554 (N_18554,N_14665,N_15011);
xnor U18555 (N_18555,N_15180,N_14051);
nor U18556 (N_18556,N_13249,N_15059);
or U18557 (N_18557,N_14220,N_15212);
and U18558 (N_18558,N_14382,N_15010);
and U18559 (N_18559,N_14597,N_14873);
nand U18560 (N_18560,N_15567,N_15102);
xnor U18561 (N_18561,N_14806,N_14361);
or U18562 (N_18562,N_14820,N_12633);
nand U18563 (N_18563,N_13570,N_13133);
nand U18564 (N_18564,N_14560,N_13982);
nor U18565 (N_18565,N_14035,N_15556);
or U18566 (N_18566,N_14887,N_15463);
nor U18567 (N_18567,N_14874,N_14546);
nor U18568 (N_18568,N_14836,N_14579);
and U18569 (N_18569,N_15167,N_15385);
and U18570 (N_18570,N_14380,N_13061);
or U18571 (N_18571,N_14955,N_12585);
nand U18572 (N_18572,N_13744,N_13845);
nand U18573 (N_18573,N_14047,N_14993);
or U18574 (N_18574,N_14045,N_12630);
nor U18575 (N_18575,N_14347,N_14596);
and U18576 (N_18576,N_12680,N_12920);
xnor U18577 (N_18577,N_14836,N_13515);
nor U18578 (N_18578,N_14939,N_15099);
nand U18579 (N_18579,N_13365,N_15532);
or U18580 (N_18580,N_13810,N_14554);
nor U18581 (N_18581,N_14579,N_14891);
and U18582 (N_18582,N_14651,N_13733);
nor U18583 (N_18583,N_12962,N_14898);
and U18584 (N_18584,N_14347,N_13691);
nor U18585 (N_18585,N_12750,N_14866);
or U18586 (N_18586,N_13569,N_12593);
or U18587 (N_18587,N_12655,N_15006);
xor U18588 (N_18588,N_15206,N_15073);
xnor U18589 (N_18589,N_13434,N_13092);
nor U18590 (N_18590,N_13774,N_14581);
and U18591 (N_18591,N_12798,N_13203);
and U18592 (N_18592,N_14253,N_14018);
or U18593 (N_18593,N_15148,N_13019);
and U18594 (N_18594,N_14289,N_14415);
and U18595 (N_18595,N_13677,N_12631);
xor U18596 (N_18596,N_12691,N_15195);
and U18597 (N_18597,N_13472,N_14763);
or U18598 (N_18598,N_12534,N_12643);
and U18599 (N_18599,N_15618,N_14527);
nand U18600 (N_18600,N_13031,N_12741);
xnor U18601 (N_18601,N_12946,N_13071);
and U18602 (N_18602,N_13365,N_13201);
nand U18603 (N_18603,N_14286,N_14132);
or U18604 (N_18604,N_15597,N_14100);
nand U18605 (N_18605,N_14863,N_14519);
or U18606 (N_18606,N_13724,N_12616);
and U18607 (N_18607,N_12677,N_13699);
and U18608 (N_18608,N_14901,N_14440);
nand U18609 (N_18609,N_13531,N_14515);
and U18610 (N_18610,N_14756,N_12917);
nand U18611 (N_18611,N_15402,N_15036);
nor U18612 (N_18612,N_12910,N_12661);
xor U18613 (N_18613,N_15310,N_12903);
and U18614 (N_18614,N_14825,N_14919);
and U18615 (N_18615,N_13182,N_13374);
nor U18616 (N_18616,N_13416,N_14788);
nor U18617 (N_18617,N_15395,N_14902);
or U18618 (N_18618,N_13444,N_14863);
xnor U18619 (N_18619,N_15178,N_14985);
or U18620 (N_18620,N_14362,N_15535);
and U18621 (N_18621,N_13373,N_12949);
and U18622 (N_18622,N_13873,N_13059);
and U18623 (N_18623,N_14338,N_15224);
nand U18624 (N_18624,N_13469,N_12669);
and U18625 (N_18625,N_15311,N_13882);
nand U18626 (N_18626,N_15500,N_13691);
or U18627 (N_18627,N_14583,N_13515);
xor U18628 (N_18628,N_14928,N_14883);
xnor U18629 (N_18629,N_12941,N_14623);
and U18630 (N_18630,N_13367,N_15439);
nor U18631 (N_18631,N_14632,N_14658);
or U18632 (N_18632,N_13610,N_13363);
nor U18633 (N_18633,N_14273,N_12657);
xor U18634 (N_18634,N_13959,N_13541);
nor U18635 (N_18635,N_15327,N_14082);
and U18636 (N_18636,N_15498,N_14487);
and U18637 (N_18637,N_14741,N_15126);
xor U18638 (N_18638,N_13137,N_13240);
xor U18639 (N_18639,N_15482,N_13951);
nor U18640 (N_18640,N_15017,N_14130);
nand U18641 (N_18641,N_14696,N_12760);
nor U18642 (N_18642,N_12512,N_14978);
nand U18643 (N_18643,N_13031,N_14280);
xnor U18644 (N_18644,N_12510,N_14142);
nor U18645 (N_18645,N_13362,N_13750);
and U18646 (N_18646,N_13950,N_12775);
nand U18647 (N_18647,N_14147,N_12744);
nor U18648 (N_18648,N_14241,N_13537);
or U18649 (N_18649,N_14912,N_13518);
xor U18650 (N_18650,N_14056,N_14249);
or U18651 (N_18651,N_14700,N_13995);
and U18652 (N_18652,N_13670,N_12889);
nand U18653 (N_18653,N_15382,N_14389);
xor U18654 (N_18654,N_13798,N_15034);
nand U18655 (N_18655,N_15338,N_12831);
xor U18656 (N_18656,N_12639,N_12949);
nor U18657 (N_18657,N_14035,N_15550);
and U18658 (N_18658,N_15343,N_12797);
and U18659 (N_18659,N_13759,N_15278);
nor U18660 (N_18660,N_14742,N_14614);
and U18661 (N_18661,N_12779,N_12917);
nor U18662 (N_18662,N_15486,N_13170);
nor U18663 (N_18663,N_12975,N_13500);
or U18664 (N_18664,N_14152,N_14882);
nand U18665 (N_18665,N_14954,N_13188);
nor U18666 (N_18666,N_14090,N_14573);
nor U18667 (N_18667,N_15501,N_15503);
and U18668 (N_18668,N_13135,N_13377);
and U18669 (N_18669,N_15135,N_15425);
nor U18670 (N_18670,N_14135,N_13661);
or U18671 (N_18671,N_14381,N_13720);
or U18672 (N_18672,N_12965,N_14443);
and U18673 (N_18673,N_14343,N_15332);
nand U18674 (N_18674,N_12556,N_12765);
nor U18675 (N_18675,N_15354,N_12916);
and U18676 (N_18676,N_13628,N_14865);
or U18677 (N_18677,N_14335,N_15050);
or U18678 (N_18678,N_13082,N_14811);
xnor U18679 (N_18679,N_14533,N_14541);
xor U18680 (N_18680,N_12543,N_12505);
and U18681 (N_18681,N_13319,N_14865);
xor U18682 (N_18682,N_12567,N_13884);
or U18683 (N_18683,N_12711,N_13164);
xnor U18684 (N_18684,N_15060,N_12768);
nor U18685 (N_18685,N_12796,N_13270);
nand U18686 (N_18686,N_14873,N_14859);
or U18687 (N_18687,N_14870,N_13028);
nand U18688 (N_18688,N_12849,N_12727);
nand U18689 (N_18689,N_13347,N_15128);
or U18690 (N_18690,N_14319,N_13802);
or U18691 (N_18691,N_14011,N_13550);
or U18692 (N_18692,N_13005,N_13398);
nand U18693 (N_18693,N_13132,N_12848);
or U18694 (N_18694,N_13967,N_12633);
nand U18695 (N_18695,N_12953,N_12621);
and U18696 (N_18696,N_15009,N_14339);
nand U18697 (N_18697,N_12834,N_14813);
nor U18698 (N_18698,N_15324,N_13878);
or U18699 (N_18699,N_13559,N_14360);
and U18700 (N_18700,N_14860,N_13912);
and U18701 (N_18701,N_14378,N_14315);
or U18702 (N_18702,N_14163,N_14096);
nor U18703 (N_18703,N_12553,N_13497);
nor U18704 (N_18704,N_12664,N_14194);
and U18705 (N_18705,N_13238,N_13205);
or U18706 (N_18706,N_15380,N_14377);
and U18707 (N_18707,N_14375,N_12899);
or U18708 (N_18708,N_13258,N_13437);
nor U18709 (N_18709,N_12643,N_15016);
xnor U18710 (N_18710,N_12537,N_13194);
nor U18711 (N_18711,N_14898,N_12785);
or U18712 (N_18712,N_12805,N_14643);
nand U18713 (N_18713,N_15119,N_12756);
xor U18714 (N_18714,N_12709,N_12941);
and U18715 (N_18715,N_15169,N_13843);
and U18716 (N_18716,N_14632,N_12852);
nor U18717 (N_18717,N_12944,N_13754);
xor U18718 (N_18718,N_13480,N_14390);
xor U18719 (N_18719,N_13959,N_14880);
or U18720 (N_18720,N_15523,N_14194);
xnor U18721 (N_18721,N_14090,N_13680);
nor U18722 (N_18722,N_14334,N_15312);
nor U18723 (N_18723,N_15068,N_14630);
nor U18724 (N_18724,N_12875,N_15035);
nor U18725 (N_18725,N_13536,N_14368);
and U18726 (N_18726,N_15613,N_15262);
nor U18727 (N_18727,N_12950,N_13417);
nor U18728 (N_18728,N_14404,N_14413);
xnor U18729 (N_18729,N_15155,N_13531);
nand U18730 (N_18730,N_14111,N_14595);
or U18731 (N_18731,N_14436,N_14885);
and U18732 (N_18732,N_14386,N_14545);
and U18733 (N_18733,N_12978,N_12559);
nor U18734 (N_18734,N_12833,N_13814);
or U18735 (N_18735,N_12884,N_14887);
nor U18736 (N_18736,N_15586,N_12780);
nand U18737 (N_18737,N_12557,N_13159);
or U18738 (N_18738,N_13515,N_13770);
xnor U18739 (N_18739,N_13692,N_14116);
or U18740 (N_18740,N_13242,N_12989);
nor U18741 (N_18741,N_13093,N_14725);
or U18742 (N_18742,N_15361,N_14313);
nor U18743 (N_18743,N_13571,N_14367);
or U18744 (N_18744,N_13925,N_14263);
or U18745 (N_18745,N_14684,N_13584);
or U18746 (N_18746,N_14583,N_14953);
xor U18747 (N_18747,N_12672,N_15566);
and U18748 (N_18748,N_13840,N_13999);
xor U18749 (N_18749,N_14867,N_13668);
nand U18750 (N_18750,N_16418,N_18306);
nand U18751 (N_18751,N_17424,N_17122);
nand U18752 (N_18752,N_15967,N_18216);
and U18753 (N_18753,N_18684,N_17196);
nor U18754 (N_18754,N_16912,N_17686);
nand U18755 (N_18755,N_16701,N_16280);
or U18756 (N_18756,N_16422,N_17646);
nor U18757 (N_18757,N_17390,N_15707);
xnor U18758 (N_18758,N_16396,N_18395);
or U18759 (N_18759,N_16640,N_17786);
or U18760 (N_18760,N_16047,N_18099);
nor U18761 (N_18761,N_15857,N_18602);
nor U18762 (N_18762,N_16983,N_18494);
xnor U18763 (N_18763,N_15915,N_17475);
and U18764 (N_18764,N_17984,N_18737);
or U18765 (N_18765,N_17528,N_18123);
nor U18766 (N_18766,N_18196,N_16827);
nor U18767 (N_18767,N_16378,N_17445);
nand U18768 (N_18768,N_17342,N_17558);
and U18769 (N_18769,N_17451,N_15982);
and U18770 (N_18770,N_17029,N_15889);
nor U18771 (N_18771,N_15813,N_18566);
or U18772 (N_18772,N_16903,N_16365);
xnor U18773 (N_18773,N_18367,N_18739);
nand U18774 (N_18774,N_17650,N_17527);
xor U18775 (N_18775,N_17677,N_18109);
nor U18776 (N_18776,N_17851,N_18187);
nor U18777 (N_18777,N_16346,N_17332);
nor U18778 (N_18778,N_17466,N_17912);
and U18779 (N_18779,N_16196,N_16156);
nor U18780 (N_18780,N_16491,N_15905);
nand U18781 (N_18781,N_16313,N_15694);
and U18782 (N_18782,N_16508,N_18372);
nor U18783 (N_18783,N_16048,N_17914);
nor U18784 (N_18784,N_18242,N_18363);
nand U18785 (N_18785,N_16004,N_18635);
or U18786 (N_18786,N_15751,N_16885);
or U18787 (N_18787,N_17322,N_16695);
and U18788 (N_18788,N_17349,N_17158);
and U18789 (N_18789,N_16992,N_18434);
nor U18790 (N_18790,N_18174,N_16381);
or U18791 (N_18791,N_16154,N_18124);
xor U18792 (N_18792,N_17160,N_18442);
nor U18793 (N_18793,N_18371,N_17099);
xnor U18794 (N_18794,N_17878,N_17643);
xnor U18795 (N_18795,N_18365,N_18671);
and U18796 (N_18796,N_18735,N_18254);
nand U18797 (N_18797,N_18037,N_16050);
nand U18798 (N_18798,N_16833,N_15923);
and U18799 (N_18799,N_16174,N_16898);
nor U18800 (N_18800,N_17499,N_17850);
nand U18801 (N_18801,N_16872,N_15850);
and U18802 (N_18802,N_18218,N_16335);
and U18803 (N_18803,N_18732,N_17753);
nand U18804 (N_18804,N_16220,N_15885);
or U18805 (N_18805,N_18585,N_16502);
nand U18806 (N_18806,N_15825,N_17371);
or U18807 (N_18807,N_16474,N_17326);
xor U18808 (N_18808,N_18258,N_16480);
and U18809 (N_18809,N_17154,N_17121);
xor U18810 (N_18810,N_17868,N_17469);
nand U18811 (N_18811,N_18164,N_18267);
or U18812 (N_18812,N_18159,N_18341);
nand U18813 (N_18813,N_17622,N_16368);
xor U18814 (N_18814,N_16802,N_15688);
nand U18815 (N_18815,N_16032,N_18741);
nand U18816 (N_18816,N_18273,N_15642);
nor U18817 (N_18817,N_16301,N_18480);
nand U18818 (N_18818,N_15812,N_17490);
nand U18819 (N_18819,N_18674,N_18065);
nor U18820 (N_18820,N_18575,N_16627);
xor U18821 (N_18821,N_16490,N_15673);
or U18822 (N_18822,N_16942,N_17308);
nor U18823 (N_18823,N_18188,N_16392);
nor U18824 (N_18824,N_15770,N_18688);
xor U18825 (N_18825,N_18304,N_15837);
xor U18826 (N_18826,N_16128,N_16109);
xor U18827 (N_18827,N_18350,N_17109);
or U18828 (N_18828,N_18580,N_16163);
nor U18829 (N_18829,N_16079,N_16201);
nand U18830 (N_18830,N_15771,N_16956);
and U18831 (N_18831,N_16941,N_18658);
nand U18832 (N_18832,N_18232,N_17929);
or U18833 (N_18833,N_17796,N_15777);
xor U18834 (N_18834,N_17899,N_17699);
and U18835 (N_18835,N_16237,N_15895);
nand U18836 (N_18836,N_17299,N_17151);
nand U18837 (N_18837,N_15750,N_18433);
or U18838 (N_18838,N_15827,N_16409);
nor U18839 (N_18839,N_16118,N_16369);
nand U18840 (N_18840,N_15679,N_16990);
nor U18841 (N_18841,N_18600,N_17297);
and U18842 (N_18842,N_18079,N_17852);
or U18843 (N_18843,N_17883,N_16923);
xnor U18844 (N_18844,N_17056,N_16347);
xnor U18845 (N_18845,N_17597,N_18525);
and U18846 (N_18846,N_18083,N_15866);
and U18847 (N_18847,N_18165,N_18260);
and U18848 (N_18848,N_16975,N_18722);
and U18849 (N_18849,N_18199,N_18457);
or U18850 (N_18850,N_18221,N_17265);
nor U18851 (N_18851,N_18102,N_17239);
xor U18852 (N_18852,N_18495,N_18193);
nand U18853 (N_18853,N_15773,N_16363);
nor U18854 (N_18854,N_17482,N_17290);
and U18855 (N_18855,N_16601,N_16634);
or U18856 (N_18856,N_16178,N_17379);
or U18857 (N_18857,N_17440,N_15891);
or U18858 (N_18858,N_18302,N_16945);
and U18859 (N_18859,N_16421,N_15809);
and U18860 (N_18860,N_18265,N_15793);
and U18861 (N_18861,N_16267,N_16931);
xnor U18862 (N_18862,N_18299,N_16781);
nor U18863 (N_18863,N_18133,N_17594);
and U18864 (N_18864,N_15911,N_16207);
nand U18865 (N_18865,N_17862,N_15988);
or U18866 (N_18866,N_17097,N_15724);
xor U18867 (N_18867,N_17938,N_16162);
nor U18868 (N_18868,N_16030,N_17285);
and U18869 (N_18869,N_17689,N_16024);
xor U18870 (N_18870,N_18535,N_17541);
or U18871 (N_18871,N_15836,N_16247);
nand U18872 (N_18872,N_16848,N_16878);
nand U18873 (N_18873,N_17542,N_18648);
nand U18874 (N_18874,N_15955,N_17657);
nand U18875 (N_18875,N_16779,N_17613);
or U18876 (N_18876,N_17694,N_17434);
nand U18877 (N_18877,N_16338,N_15849);
or U18878 (N_18878,N_16013,N_18522);
nand U18879 (N_18879,N_17685,N_17131);
nand U18880 (N_18880,N_17281,N_18548);
nand U18881 (N_18881,N_16009,N_18019);
and U18882 (N_18882,N_18470,N_17092);
and U18883 (N_18883,N_17335,N_16062);
and U18884 (N_18884,N_18550,N_17300);
or U18885 (N_18885,N_16169,N_17715);
and U18886 (N_18886,N_18016,N_17830);
nand U18887 (N_18887,N_16223,N_18545);
xnor U18888 (N_18888,N_18742,N_18042);
xnor U18889 (N_18889,N_17415,N_16959);
nand U18890 (N_18890,N_16587,N_18107);
or U18891 (N_18891,N_16051,N_17827);
xor U18892 (N_18892,N_16159,N_17125);
and U18893 (N_18893,N_17754,N_15740);
nor U18894 (N_18894,N_17467,N_18130);
nand U18895 (N_18895,N_17804,N_15869);
nor U18896 (N_18896,N_16110,N_17910);
and U18897 (N_18897,N_18423,N_16729);
and U18898 (N_18898,N_15961,N_17631);
nor U18899 (N_18899,N_16749,N_15629);
nor U18900 (N_18900,N_17141,N_18644);
nand U18901 (N_18901,N_16844,N_15820);
xor U18902 (N_18902,N_16011,N_16528);
nand U18903 (N_18903,N_17967,N_17897);
and U18904 (N_18904,N_16948,N_17835);
nor U18905 (N_18905,N_17230,N_16610);
or U18906 (N_18906,N_15854,N_17751);
xnor U18907 (N_18907,N_15989,N_17085);
nor U18908 (N_18908,N_18361,N_16465);
or U18909 (N_18909,N_16193,N_17904);
nor U18910 (N_18910,N_16297,N_17175);
or U18911 (N_18911,N_16241,N_18264);
or U18912 (N_18912,N_17271,N_15680);
nand U18913 (N_18913,N_16440,N_15721);
nor U18914 (N_18914,N_16622,N_18615);
or U18915 (N_18915,N_16044,N_17351);
nand U18916 (N_18916,N_17714,N_16525);
nor U18917 (N_18917,N_17435,N_16387);
and U18918 (N_18918,N_16718,N_17037);
or U18919 (N_18919,N_18555,N_17846);
or U18920 (N_18920,N_15819,N_18052);
nand U18921 (N_18921,N_17978,N_17656);
nor U18922 (N_18922,N_16897,N_17142);
nand U18923 (N_18923,N_15862,N_18604);
nand U18924 (N_18924,N_16716,N_16105);
nand U18925 (N_18925,N_17430,N_18458);
or U18926 (N_18926,N_16319,N_18077);
xnor U18927 (N_18927,N_16035,N_16688);
xor U18928 (N_18928,N_16406,N_16657);
nand U18929 (N_18929,N_16764,N_17135);
xor U18930 (N_18930,N_16822,N_17381);
nand U18931 (N_18931,N_18476,N_16253);
nor U18932 (N_18932,N_15652,N_16208);
nor U18933 (N_18933,N_16702,N_18129);
nor U18934 (N_18934,N_18028,N_18374);
nand U18935 (N_18935,N_17211,N_16788);
xnor U18936 (N_18936,N_18700,N_17633);
and U18937 (N_18937,N_18511,N_18679);
nor U18938 (N_18938,N_17449,N_18316);
nand U18939 (N_18939,N_16678,N_16179);
or U18940 (N_18940,N_16782,N_15910);
or U18941 (N_18941,N_17834,N_16619);
or U18942 (N_18942,N_15698,N_15904);
and U18943 (N_18943,N_16513,N_17021);
xor U18944 (N_18944,N_16315,N_16733);
nor U18945 (N_18945,N_15835,N_16265);
or U18946 (N_18946,N_18455,N_16521);
and U18947 (N_18947,N_17526,N_17875);
nor U18948 (N_18948,N_17040,N_16883);
xor U18949 (N_18949,N_16857,N_18178);
nand U18950 (N_18950,N_17462,N_18271);
or U18951 (N_18951,N_18493,N_17116);
xnor U18952 (N_18952,N_17781,N_16081);
nand U18953 (N_18953,N_17437,N_17212);
nand U18954 (N_18954,N_18094,N_18010);
xnor U18955 (N_18955,N_16710,N_18610);
or U18956 (N_18956,N_16479,N_17492);
nor U18957 (N_18957,N_18689,N_16921);
nand U18958 (N_18958,N_17771,N_15728);
nor U18959 (N_18959,N_17928,N_18662);
and U18960 (N_18960,N_17011,N_17620);
xor U18961 (N_18961,N_18413,N_17429);
and U18962 (N_18962,N_18436,N_17586);
nor U18963 (N_18963,N_18261,N_17399);
nand U18964 (N_18964,N_17538,N_16344);
or U18965 (N_18965,N_18315,N_17168);
or U18966 (N_18966,N_18736,N_18108);
and U18967 (N_18967,N_16639,N_16626);
nand U18968 (N_18968,N_16111,N_16439);
and U18969 (N_18969,N_17892,N_17775);
nand U18970 (N_18970,N_18200,N_16845);
nor U18971 (N_18971,N_17525,N_15826);
nor U18972 (N_18972,N_16616,N_17902);
or U18973 (N_18973,N_15662,N_16676);
nand U18974 (N_18974,N_15717,N_16842);
and U18975 (N_18975,N_16239,N_18749);
and U18976 (N_18976,N_16852,N_17707);
and U18977 (N_18977,N_17843,N_15716);
xnor U18978 (N_18978,N_18418,N_18672);
nor U18979 (N_18979,N_18710,N_16233);
and U18980 (N_18980,N_17070,N_16570);
and U18981 (N_18981,N_17411,N_16431);
nand U18982 (N_18982,N_16648,N_16767);
xor U18983 (N_18983,N_16447,N_17844);
or U18984 (N_18984,N_17520,N_16412);
and U18985 (N_18985,N_16063,N_15661);
or U18986 (N_18986,N_16561,N_15647);
nand U18987 (N_18987,N_16136,N_17829);
or U18988 (N_18988,N_17414,N_17857);
xor U18989 (N_18989,N_18369,N_17367);
nand U18990 (N_18990,N_16500,N_17343);
xnor U18991 (N_18991,N_16219,N_17792);
or U18992 (N_18992,N_17177,N_16843);
xor U18993 (N_18993,N_16955,N_17106);
and U18994 (N_18994,N_18426,N_15699);
and U18995 (N_18995,N_17301,N_18088);
and U18996 (N_18996,N_18699,N_18705);
or U18997 (N_18997,N_18068,N_15990);
or U18998 (N_18998,N_16372,N_16769);
nor U18999 (N_18999,N_17999,N_17809);
xnor U19000 (N_19000,N_17331,N_17355);
xnor U19001 (N_19001,N_17478,N_17522);
nand U19002 (N_19002,N_18145,N_16064);
nand U19003 (N_19003,N_15842,N_18701);
nand U19004 (N_19004,N_17096,N_17727);
nand U19005 (N_19005,N_16867,N_18148);
or U19006 (N_19006,N_17917,N_17485);
nand U19007 (N_19007,N_18569,N_18243);
xor U19008 (N_19008,N_16821,N_16180);
nor U19009 (N_19009,N_18355,N_18351);
xor U19010 (N_19010,N_17731,N_17457);
and U19011 (N_19011,N_18308,N_18723);
xnor U19012 (N_19012,N_17410,N_17934);
nand U19013 (N_19013,N_16578,N_18091);
xnor U19014 (N_19014,N_16123,N_16061);
xnor U19015 (N_19015,N_16913,N_18044);
nor U19016 (N_19016,N_16139,N_15778);
or U19017 (N_19017,N_18431,N_17982);
and U19018 (N_19018,N_16863,N_15737);
xnor U19019 (N_19019,N_17975,N_17232);
and U19020 (N_19020,N_18534,N_17812);
and U19021 (N_19021,N_15945,N_16184);
nor U19022 (N_19022,N_17651,N_16707);
nand U19023 (N_19023,N_16091,N_16007);
or U19024 (N_19024,N_16294,N_17372);
xor U19025 (N_19025,N_17798,N_15675);
xor U19026 (N_19026,N_17276,N_16635);
xor U19027 (N_19027,N_18160,N_18336);
nor U19028 (N_19028,N_17560,N_16978);
xor U19029 (N_19029,N_17913,N_17334);
or U19030 (N_19030,N_15758,N_18041);
nor U19031 (N_19031,N_17662,N_18390);
nand U19032 (N_19032,N_16287,N_16302);
or U19033 (N_19033,N_18570,N_17666);
xor U19034 (N_19034,N_16874,N_18360);
nor U19035 (N_19035,N_17842,N_18150);
and U19036 (N_19036,N_17652,N_17537);
nor U19037 (N_19037,N_17100,N_16653);
or U19038 (N_19038,N_16073,N_16515);
nor U19039 (N_19039,N_17126,N_17139);
and U19040 (N_19040,N_16311,N_17223);
and U19041 (N_19041,N_16436,N_16066);
or U19042 (N_19042,N_15977,N_15829);
nor U19043 (N_19043,N_18021,N_18496);
xor U19044 (N_19044,N_18643,N_16454);
nand U19045 (N_19045,N_18599,N_16999);
xor U19046 (N_19046,N_18562,N_17236);
xor U19047 (N_19047,N_16630,N_17684);
nand U19048 (N_19048,N_15880,N_17019);
nand U19049 (N_19049,N_17907,N_18269);
and U19050 (N_19050,N_16886,N_16336);
nor U19051 (N_19051,N_16958,N_18449);
nor U19052 (N_19052,N_16893,N_16896);
or U19053 (N_19053,N_15900,N_18270);
nor U19054 (N_19054,N_16254,N_16160);
nand U19055 (N_19055,N_17136,N_15907);
and U19056 (N_19056,N_16202,N_15938);
nand U19057 (N_19057,N_16488,N_17432);
and U19058 (N_19058,N_18393,N_17979);
nor U19059 (N_19059,N_16838,N_18428);
nand U19060 (N_19060,N_17307,N_15958);
nand U19061 (N_19061,N_17494,N_17316);
and U19062 (N_19062,N_15745,N_15660);
nand U19063 (N_19063,N_17629,N_18314);
and U19064 (N_19064,N_17007,N_16646);
and U19065 (N_19065,N_16849,N_18111);
nand U19066 (N_19066,N_17252,N_18466);
xor U19067 (N_19067,N_16443,N_16637);
nand U19068 (N_19068,N_18451,N_17841);
nor U19069 (N_19069,N_17228,N_16216);
nor U19070 (N_19070,N_15790,N_15784);
nand U19071 (N_19071,N_16632,N_17318);
and U19072 (N_19072,N_16868,N_17296);
nor U19073 (N_19073,N_17200,N_17973);
and U19074 (N_19074,N_16564,N_18376);
nor U19075 (N_19075,N_15851,N_18617);
and U19076 (N_19076,N_16181,N_17716);
xor U19077 (N_19077,N_15796,N_17075);
xnor U19078 (N_19078,N_16462,N_15656);
nor U19079 (N_19079,N_18388,N_16582);
and U19080 (N_19080,N_16227,N_16793);
and U19081 (N_19081,N_15874,N_17014);
or U19082 (N_19082,N_15929,N_16703);
xnor U19083 (N_19083,N_15934,N_17760);
nand U19084 (N_19084,N_16122,N_16042);
xor U19085 (N_19085,N_16829,N_17222);
or U19086 (N_19086,N_17112,N_16082);
nor U19087 (N_19087,N_16970,N_16040);
or U19088 (N_19088,N_15808,N_17346);
or U19089 (N_19089,N_18183,N_16402);
nand U19090 (N_19090,N_18596,N_18556);
and U19091 (N_19091,N_17616,N_16060);
or U19092 (N_19092,N_17653,N_17611);
or U19093 (N_19093,N_18076,N_18638);
or U19094 (N_19094,N_17164,N_18344);
or U19095 (N_19095,N_18169,N_17404);
nand U19096 (N_19096,N_17217,N_16466);
nand U19097 (N_19097,N_18170,N_16674);
or U19098 (N_19098,N_17582,N_16373);
xnor U19099 (N_19099,N_15669,N_18190);
and U19100 (N_19100,N_17737,N_15823);
nand U19101 (N_19101,N_15760,N_16261);
xnor U19102 (N_19102,N_17974,N_15810);
nor U19103 (N_19103,N_16998,N_15863);
or U19104 (N_19104,N_16460,N_17215);
nand U19105 (N_19105,N_17110,N_18586);
nand U19106 (N_19106,N_15950,N_16737);
xor U19107 (N_19107,N_17491,N_15814);
and U19108 (N_19108,N_16537,N_16078);
and U19109 (N_19109,N_18347,N_16075);
and U19110 (N_19110,N_15943,N_17484);
or U19111 (N_19111,N_17602,N_18207);
or U19112 (N_19112,N_16380,N_15697);
xnor U19113 (N_19113,N_15730,N_18379);
or U19114 (N_19114,N_17920,N_17532);
and U19115 (N_19115,N_18069,N_17634);
nor U19116 (N_19116,N_18239,N_15695);
xnor U19117 (N_19117,N_16628,N_17801);
and U19118 (N_19118,N_15918,N_18081);
nor U19119 (N_19119,N_16807,N_18438);
or U19120 (N_19120,N_17257,N_18128);
nor U19121 (N_19121,N_16329,N_17359);
nand U19122 (N_19122,N_16670,N_15725);
and U19123 (N_19123,N_17423,N_15672);
and U19124 (N_19124,N_16012,N_17887);
xnor U19125 (N_19125,N_17598,N_18642);
xnor U19126 (N_19126,N_17032,N_15916);
or U19127 (N_19127,N_15775,N_18197);
xnor U19128 (N_19128,N_17824,N_16232);
nand U19129 (N_19129,N_18713,N_17630);
and U19130 (N_19130,N_16285,N_15710);
nor U19131 (N_19131,N_15876,N_17521);
xnor U19132 (N_19132,N_16917,N_15683);
nor U19133 (N_19133,N_16292,N_17347);
xnor U19134 (N_19134,N_17159,N_17937);
nor U19135 (N_19135,N_18447,N_17969);
nand U19136 (N_19136,N_16112,N_17407);
nand U19137 (N_19137,N_16924,N_17024);
or U19138 (N_19138,N_18387,N_16747);
xnor U19139 (N_19139,N_16882,N_17703);
nor U19140 (N_19140,N_18313,N_17728);
xnor U19141 (N_19141,N_17782,N_17584);
and U19142 (N_19142,N_17291,N_17480);
and U19143 (N_19143,N_18320,N_18504);
xnor U19144 (N_19144,N_17488,N_18718);
or U19145 (N_19145,N_17524,N_17260);
nand U19146 (N_19146,N_18587,N_15914);
nor U19147 (N_19147,N_18034,N_16652);
nor U19148 (N_19148,N_18446,N_17049);
nor U19149 (N_19149,N_16993,N_16016);
nand U19150 (N_19150,N_16449,N_16120);
nand U19151 (N_19151,N_16830,N_16919);
xnor U19152 (N_19152,N_18523,N_17838);
and U19153 (N_19153,N_18595,N_15935);
or U19154 (N_19154,N_16904,N_17793);
nor U19155 (N_19155,N_18463,N_17785);
xor U19156 (N_19156,N_16819,N_17225);
xor U19157 (N_19157,N_17368,N_17628);
or U19158 (N_19158,N_16498,N_16114);
nor U19159 (N_19159,N_18245,N_16090);
or U19160 (N_19160,N_16145,N_16014);
xnor U19161 (N_19161,N_16385,N_17762);
or U19162 (N_19162,N_16730,N_16273);
or U19163 (N_19163,N_16721,N_16167);
nor U19164 (N_19164,N_18009,N_16477);
or U19165 (N_19165,N_15639,N_18236);
or U19166 (N_19166,N_17171,N_17943);
nand U19167 (N_19167,N_16383,N_16669);
xor U19168 (N_19168,N_18669,N_16651);
or U19169 (N_19169,N_15785,N_16765);
nor U19170 (N_19170,N_18105,N_17214);
or U19171 (N_19171,N_16608,N_16586);
xor U19172 (N_19172,N_16790,N_16731);
and U19173 (N_19173,N_17481,N_18062);
xnor U19174 (N_19174,N_16679,N_16994);
nor U19175 (N_19175,N_16834,N_17916);
or U19176 (N_19176,N_17565,N_17990);
nor U19177 (N_19177,N_17726,N_17618);
xnor U19178 (N_19178,N_16579,N_18411);
and U19179 (N_19179,N_17877,N_17047);
xnor U19180 (N_19180,N_17038,N_17576);
and U19181 (N_19181,N_15912,N_15888);
nand U19182 (N_19182,N_17879,N_18537);
nor U19183 (N_19183,N_15913,N_18368);
nor U19184 (N_19184,N_16937,N_18726);
or U19185 (N_19185,N_16661,N_17819);
xnor U19186 (N_19186,N_17854,N_15879);
xor U19187 (N_19187,N_18180,N_15702);
nor U19188 (N_19188,N_18227,N_16633);
nor U19189 (N_19189,N_15706,N_16377);
and U19190 (N_19190,N_16812,N_18690);
xnor U19191 (N_19191,N_16687,N_18120);
xor U19192 (N_19192,N_18237,N_17645);
nor U19193 (N_19193,N_17288,N_16029);
nor U19194 (N_19194,N_17455,N_18384);
xnor U19195 (N_19195,N_17235,N_17770);
nand U19196 (N_19196,N_18552,N_17065);
and U19197 (N_19197,N_17204,N_18695);
or U19198 (N_19198,N_18693,N_18043);
and U19199 (N_19199,N_18132,N_15663);
xor U19200 (N_19200,N_18712,N_17808);
xor U19201 (N_19201,N_16906,N_18746);
or U19202 (N_19202,N_17376,N_16416);
nand U19203 (N_19203,N_18122,N_17226);
or U19204 (N_19204,N_16533,N_18356);
or U19205 (N_19205,N_17941,N_17464);
and U19206 (N_19206,N_18698,N_17738);
xnor U19207 (N_19207,N_16583,N_17741);
and U19208 (N_19208,N_17776,N_18483);
nor U19209 (N_19209,N_16398,N_18364);
or U19210 (N_19210,N_17279,N_16144);
nor U19211 (N_19211,N_16573,N_17057);
and U19212 (N_19212,N_18637,N_15992);
or U19213 (N_19213,N_16960,N_18096);
xor U19214 (N_19214,N_17698,N_17166);
and U19215 (N_19215,N_17534,N_18667);
nand U19216 (N_19216,N_16113,N_16916);
or U19217 (N_19217,N_17321,N_17642);
or U19218 (N_19218,N_15844,N_17385);
nor U19219 (N_19219,N_16323,N_17968);
nor U19220 (N_19220,N_17950,N_16170);
xor U19221 (N_19221,N_18085,N_15644);
xor U19222 (N_19222,N_17035,N_16119);
xnor U19223 (N_19223,N_17387,N_18506);
and U19224 (N_19224,N_17419,N_18275);
nand U19225 (N_19225,N_16437,N_16245);
nand U19226 (N_19226,N_18318,N_16859);
xor U19227 (N_19227,N_17176,N_16127);
or U19228 (N_19228,N_16229,N_16453);
nor U19229 (N_19229,N_17293,N_17555);
nor U19230 (N_19230,N_18161,N_18163);
and U19231 (N_19231,N_18597,N_15763);
and U19232 (N_19232,N_17303,N_17794);
xor U19233 (N_19233,N_16551,N_18115);
nand U19234 (N_19234,N_17831,N_16801);
nor U19235 (N_19235,N_17895,N_18073);
nor U19236 (N_19236,N_18640,N_17172);
xor U19237 (N_19237,N_16148,N_15719);
nand U19238 (N_19238,N_17180,N_18708);
nor U19239 (N_19239,N_18567,N_15795);
nor U19240 (N_19240,N_18492,N_17361);
nor U19241 (N_19241,N_16925,N_16214);
nand U19242 (N_19242,N_17557,N_17401);
and U19243 (N_19243,N_16153,N_16408);
and U19244 (N_19244,N_17863,N_17588);
and U19245 (N_19245,N_18561,N_18683);
or U19246 (N_19246,N_16920,N_16277);
or U19247 (N_19247,N_15759,N_16281);
or U19248 (N_19248,N_16589,N_17329);
xnor U19249 (N_19249,N_17766,N_16117);
xnor U19250 (N_19250,N_15986,N_16070);
nand U19251 (N_19251,N_17416,N_16182);
nor U19252 (N_19252,N_17523,N_16361);
nand U19253 (N_19253,N_17599,N_17570);
and U19254 (N_19254,N_16441,N_17474);
nand U19255 (N_19255,N_18654,N_16940);
or U19256 (N_19256,N_16256,N_18452);
and U19257 (N_19257,N_17197,N_16699);
xor U19258 (N_19258,N_16086,N_18342);
nor U19259 (N_19259,N_18665,N_16494);
nor U19260 (N_19260,N_18673,N_16420);
nand U19261 (N_19261,N_17764,N_15657);
nor U19262 (N_19262,N_16791,N_16472);
nor U19263 (N_19263,N_17327,N_16262);
xor U19264 (N_19264,N_16668,N_18526);
nand U19265 (N_19265,N_17612,N_17269);
xnor U19266 (N_19266,N_18307,N_17128);
xor U19267 (N_19267,N_18629,N_16609);
nand U19268 (N_19268,N_17655,N_16015);
or U19269 (N_19269,N_18560,N_15797);
nand U19270 (N_19270,N_16951,N_17015);
nor U19271 (N_19271,N_16936,N_18182);
nor U19272 (N_19272,N_17903,N_17210);
or U19273 (N_19273,N_17319,N_18415);
nand U19274 (N_19274,N_17661,N_17272);
xnor U19275 (N_19275,N_16892,N_16663);
and U19276 (N_19276,N_18490,N_16445);
and U19277 (N_19277,N_16224,N_17626);
or U19278 (N_19278,N_16165,N_16811);
and U19279 (N_19279,N_16946,N_18031);
nand U19280 (N_19280,N_16976,N_18139);
or U19281 (N_19281,N_16820,N_15696);
nor U19282 (N_19282,N_17313,N_16103);
or U19283 (N_19283,N_18720,N_15631);
or U19284 (N_19284,N_16806,N_17667);
or U19285 (N_19285,N_15994,N_17817);
and U19286 (N_19286,N_17076,N_17098);
or U19287 (N_19287,N_16231,N_16600);
nand U19288 (N_19288,N_18416,N_17169);
and U19289 (N_19289,N_17644,N_16371);
xor U19290 (N_19290,N_16348,N_16683);
or U19291 (N_19291,N_17995,N_16080);
and U19292 (N_19292,N_16248,N_16706);
or U19293 (N_19293,N_16226,N_16655);
or U19294 (N_19294,N_16038,N_18536);
xnor U19295 (N_19295,N_16520,N_16682);
and U19296 (N_19296,N_17050,N_15995);
nand U19297 (N_19297,N_16891,N_17583);
xnor U19298 (N_19298,N_15767,N_17045);
nor U19299 (N_19299,N_15731,N_15957);
nand U19300 (N_19300,N_16714,N_17706);
or U19301 (N_19301,N_16724,N_16359);
or U19302 (N_19302,N_17921,N_18510);
nand U19303 (N_19303,N_16877,N_17548);
nor U19304 (N_19304,N_16271,N_18377);
nand U19305 (N_19305,N_18740,N_16950);
and U19306 (N_19306,N_15847,N_17183);
nand U19307 (N_19307,N_18322,N_15840);
xnor U19308 (N_19308,N_16138,N_16341);
xnor U19309 (N_19309,N_18459,N_16902);
and U19310 (N_19310,N_16129,N_17826);
and U19311 (N_19311,N_15956,N_17665);
or U19312 (N_19312,N_18056,N_17273);
xor U19313 (N_19313,N_17227,N_18274);
xnor U19314 (N_19314,N_18659,N_17418);
nand U19315 (N_19315,N_17093,N_18082);
or U19316 (N_19316,N_18398,N_17615);
or U19317 (N_19317,N_15828,N_17403);
nand U19318 (N_19318,N_16684,N_17510);
xnor U19319 (N_19319,N_16147,N_16415);
and U19320 (N_19320,N_16991,N_17813);
xor U19321 (N_19321,N_16215,N_15898);
or U19322 (N_19322,N_16864,N_16268);
or U19323 (N_19323,N_15746,N_16673);
and U19324 (N_19324,N_18554,N_16777);
xnor U19325 (N_19325,N_16003,N_17540);
nand U19326 (N_19326,N_16739,N_18626);
and U19327 (N_19327,N_16473,N_17039);
nor U19328 (N_19328,N_18685,N_18263);
or U19329 (N_19329,N_15817,N_16183);
or U19330 (N_19330,N_17102,N_18709);
nor U19331 (N_19331,N_18655,N_15887);
or U19332 (N_19332,N_18385,N_17971);
nor U19333 (N_19333,N_17016,N_17593);
xor U19334 (N_19334,N_18294,N_16141);
nand U19335 (N_19335,N_16787,N_18162);
nor U19336 (N_19336,N_17668,N_17060);
and U19337 (N_19337,N_17987,N_16686);
nor U19338 (N_19338,N_15867,N_15886);
or U19339 (N_19339,N_18482,N_17043);
xor U19340 (N_19340,N_18229,N_16058);
or U19341 (N_19341,N_15648,N_18167);
and U19342 (N_19342,N_17756,N_16696);
or U19343 (N_19343,N_18345,N_17022);
xor U19344 (N_19344,N_15674,N_15757);
and U19345 (N_19345,N_17384,N_18632);
xor U19346 (N_19346,N_16928,N_18469);
nand U19347 (N_19347,N_17044,N_17298);
xnor U19348 (N_19348,N_18406,N_17509);
and U19349 (N_19349,N_16880,N_16794);
nor U19350 (N_19350,N_17193,N_17880);
nand U19351 (N_19351,N_16131,N_17787);
or U19352 (N_19352,N_17088,N_16862);
nand U19353 (N_19353,N_17977,N_17953);
nor U19354 (N_19354,N_17549,N_16763);
nor U19355 (N_19355,N_18158,N_18131);
or U19356 (N_19356,N_16158,N_15933);
xnor U19357 (N_19357,N_16264,N_16979);
and U19358 (N_19358,N_16027,N_17828);
and U19359 (N_19359,N_16823,N_17396);
nand U19360 (N_19360,N_16282,N_17717);
nand U19361 (N_19361,N_16527,N_15816);
nor U19362 (N_19362,N_18616,N_18675);
or U19363 (N_19363,N_16545,N_16391);
or U19364 (N_19364,N_16212,N_17339);
or U19365 (N_19365,N_16918,N_17507);
nand U19366 (N_19366,N_17012,N_17240);
xnor U19367 (N_19367,N_17394,N_17614);
or U19368 (N_19368,N_16017,N_17471);
xor U19369 (N_19369,N_18175,N_18472);
and U19370 (N_19370,N_16853,N_16865);
and U19371 (N_19371,N_18694,N_18233);
or U19372 (N_19372,N_18008,N_16690);
or U19373 (N_19373,N_17295,N_17051);
nor U19374 (N_19374,N_16428,N_17278);
or U19375 (N_19375,N_16762,N_18417);
xnor U19376 (N_19376,N_17229,N_17077);
and U19377 (N_19377,N_18185,N_16279);
xnor U19378 (N_19378,N_18486,N_17010);
and U19379 (N_19379,N_17205,N_15748);
nand U19380 (N_19380,N_17283,N_17859);
and U19381 (N_19381,N_15834,N_18508);
or U19382 (N_19382,N_17911,N_16519);
nand U19383 (N_19383,N_15811,N_18184);
and U19384 (N_19384,N_17002,N_16166);
or U19385 (N_19385,N_16356,N_17042);
xnor U19386 (N_19386,N_17115,N_17104);
and U19387 (N_19387,N_17940,N_16759);
nor U19388 (N_19388,N_18298,N_18250);
and U19389 (N_19389,N_16711,N_17062);
xnor U19390 (N_19390,N_16967,N_16553);
xor U19391 (N_19391,N_17413,N_17033);
nand U19392 (N_19392,N_18252,N_16125);
and U19393 (N_19393,N_16033,N_18619);
nor U19394 (N_19394,N_17972,N_18026);
or U19395 (N_19395,N_16025,N_16795);
nor U19396 (N_19396,N_17948,N_16005);
xnor U19397 (N_19397,N_16299,N_17769);
nand U19398 (N_19398,N_17263,N_15917);
xnor U19399 (N_19399,N_17610,N_16354);
nor U19400 (N_19400,N_17700,N_15727);
nor U19401 (N_19401,N_17930,N_16825);
xnor U19402 (N_19402,N_16276,N_16799);
nand U19403 (N_19403,N_17018,N_17933);
nand U19404 (N_19404,N_15635,N_16780);
nor U19405 (N_19405,N_17130,N_15801);
xor U19406 (N_19406,N_16680,N_15650);
xor U19407 (N_19407,N_15779,N_17186);
nor U19408 (N_19408,N_16001,N_16290);
and U19409 (N_19409,N_16557,N_17124);
nor U19410 (N_19410,N_18136,N_16102);
xnor U19411 (N_19411,N_17508,N_18479);
or U19412 (N_19412,N_18030,N_15800);
or U19413 (N_19413,N_16321,N_17837);
nand U19414 (N_19414,N_17544,N_18605);
nand U19415 (N_19415,N_17997,N_17292);
nand U19416 (N_19416,N_16884,N_16031);
or U19417 (N_19417,N_18657,N_18633);
or U19418 (N_19418,N_15638,N_18464);
nor U19419 (N_19419,N_16401,N_15979);
nand U19420 (N_19420,N_18234,N_17162);
xor U19421 (N_19421,N_17654,N_18471);
nor U19422 (N_19422,N_16735,N_18513);
nor U19423 (N_19423,N_16400,N_17071);
and U19424 (N_19424,N_17153,N_15772);
nor U19425 (N_19425,N_18524,N_18116);
nand U19426 (N_19426,N_16831,N_17129);
xor U19427 (N_19427,N_17882,N_17194);
xnor U19428 (N_19428,N_16559,N_17487);
nor U19429 (N_19429,N_18577,N_18329);
nor U19430 (N_19430,N_17073,N_16195);
or U19431 (N_19431,N_15920,N_17103);
nor U19432 (N_19432,N_18064,N_17743);
xnor U19433 (N_19433,N_15872,N_15948);
nor U19434 (N_19434,N_17395,N_15766);
or U19435 (N_19435,N_17561,N_16429);
and U19436 (N_19436,N_16617,N_15882);
or U19437 (N_19437,N_15940,N_18231);
or U19438 (N_19438,N_18146,N_17960);
xnor U19439 (N_19439,N_16961,N_18639);
nand U19440 (N_19440,N_16623,N_15975);
or U19441 (N_19441,N_15756,N_16349);
nor U19442 (N_19442,N_18512,N_15792);
or U19443 (N_19443,N_17748,N_17233);
xnor U19444 (N_19444,N_17408,N_17983);
nand U19445 (N_19445,N_18238,N_16873);
nor U19446 (N_19446,N_16296,N_15909);
nand U19447 (N_19447,N_17774,N_17409);
and U19448 (N_19448,N_17188,N_17736);
xor U19449 (N_19449,N_18613,N_17918);
and U19450 (N_19450,N_16469,N_17784);
or U19451 (N_19451,N_18421,N_17256);
xnor U19452 (N_19452,N_17167,N_17761);
xnor U19453 (N_19453,N_18309,N_17406);
xor U19454 (N_19454,N_17203,N_15969);
nand U19455 (N_19455,N_17519,N_18023);
and U19456 (N_19456,N_18734,N_17266);
nand U19457 (N_19457,N_16715,N_15711);
xor U19458 (N_19458,N_16339,N_17589);
xor U19459 (N_19459,N_17500,N_16059);
or U19460 (N_19460,N_16283,N_17695);
nand U19461 (N_19461,N_15821,N_18444);
and U19462 (N_19462,N_17670,N_17201);
and U19463 (N_19463,N_17729,N_17778);
or U19464 (N_19464,N_18149,N_17250);
nand U19465 (N_19465,N_15693,N_17951);
nand U19466 (N_19466,N_18389,N_16423);
nand U19467 (N_19467,N_17143,N_15976);
or U19468 (N_19468,N_18500,N_16203);
and U19469 (N_19469,N_17323,N_15765);
nor U19470 (N_19470,N_15682,N_15984);
xor U19471 (N_19471,N_17350,N_16540);
nor U19472 (N_19472,N_18202,N_16547);
xnor U19473 (N_19473,N_17120,N_17874);
or U19474 (N_19474,N_16952,N_16758);
and U19475 (N_19475,N_17815,N_16211);
or U19476 (N_19476,N_16331,N_16037);
xnor U19477 (N_19477,N_16375,N_18286);
or U19478 (N_19478,N_16343,N_18396);
nand U19479 (N_19479,N_16602,N_16108);
nor U19480 (N_19480,N_17202,N_18151);
nor U19481 (N_19481,N_16901,N_16046);
nand U19482 (N_19482,N_16809,N_16953);
nand U19483 (N_19483,N_17606,N_16543);
nand U19484 (N_19484,N_17064,N_16756);
nor U19485 (N_19485,N_16350,N_15718);
and U19486 (N_19486,N_15881,N_17402);
nand U19487 (N_19487,N_16189,N_18327);
nor U19488 (N_19488,N_16286,N_17111);
xnor U19489 (N_19489,N_16278,N_17268);
or U19490 (N_19490,N_15733,N_17375);
nand U19491 (N_19491,N_18641,N_16006);
nand U19492 (N_19492,N_18551,N_16671);
nand U19493 (N_19493,N_17574,N_18594);
nor U19494 (N_19494,N_17688,N_18035);
nand U19495 (N_19495,N_18189,N_16258);
nor U19496 (N_19496,N_16768,N_18291);
nand U19497 (N_19497,N_16352,N_17777);
or U19498 (N_19498,N_16101,N_16629);
nor U19499 (N_19499,N_15833,N_16725);
or U19500 (N_19500,N_18530,N_18220);
nand U19501 (N_19501,N_17459,N_15712);
nand U19502 (N_19502,N_17363,N_16360);
or U19503 (N_19503,N_16870,N_16355);
nand U19504 (N_19504,N_15927,N_16798);
nand U19505 (N_19505,N_17704,N_16362);
or U19506 (N_19506,N_16565,N_18362);
and U19507 (N_19507,N_18553,N_16908);
xor U19508 (N_19508,N_15692,N_18498);
and U19509 (N_19509,N_18422,N_15686);
and U19510 (N_19510,N_17147,N_17577);
nor U19511 (N_19511,N_16659,N_17078);
nor U19512 (N_19512,N_18576,N_17674);
or U19513 (N_19513,N_16740,N_16419);
nand U19514 (N_19514,N_17242,N_18072);
and U19515 (N_19515,N_17539,N_17725);
xnor U19516 (N_19516,N_16693,N_16571);
nor U19517 (N_19517,N_17989,N_18692);
or U19518 (N_19518,N_15883,N_16743);
and U19519 (N_19519,N_18090,N_18288);
or U19520 (N_19520,N_18305,N_16643);
xnor U19521 (N_19521,N_17939,N_18729);
nand U19522 (N_19522,N_18001,N_17005);
nor U19523 (N_19523,N_17552,N_15864);
or U19524 (N_19524,N_16306,N_18330);
and U19525 (N_19525,N_17393,N_16700);
xor U19526 (N_19526,N_18101,N_18489);
and U19527 (N_19527,N_18696,N_16505);
or U19528 (N_19528,N_18140,N_16784);
nor U19529 (N_19529,N_16753,N_16218);
nand U19530 (N_19530,N_15769,N_16818);
and U19531 (N_19531,N_18110,N_15684);
xnor U19532 (N_19532,N_17720,N_18249);
nand U19533 (N_19533,N_16618,N_18359);
xor U19534 (N_19534,N_15936,N_18590);
and U19535 (N_19535,N_15666,N_15993);
nor U19536 (N_19536,N_18625,N_18104);
nor U19537 (N_19537,N_15921,N_18002);
xnor U19538 (N_19538,N_17004,N_17340);
and U19539 (N_19539,N_17908,N_16484);
nand U19540 (N_19540,N_17218,N_17282);
and U19541 (N_19541,N_18003,N_18205);
nand U19542 (N_19542,N_17516,N_17458);
or U19543 (N_19543,N_15901,N_17832);
or U19544 (N_19544,N_16965,N_16766);
nand U19545 (N_19545,N_15681,N_16855);
or U19546 (N_19546,N_17277,N_17926);
nor U19547 (N_19547,N_16450,N_15818);
nor U19548 (N_19548,N_16092,N_18589);
or U19549 (N_19549,N_16624,N_16647);
nand U19550 (N_19550,N_18386,N_16552);
nor U19551 (N_19551,N_16567,N_18208);
and U19552 (N_19552,N_16096,N_16010);
or U19553 (N_19553,N_17805,N_15704);
nand U19554 (N_19554,N_17069,N_18717);
and U19555 (N_19555,N_18211,N_18018);
or U19556 (N_19556,N_18046,N_16434);
and U19557 (N_19557,N_16252,N_16792);
nand U19558 (N_19558,N_16835,N_16881);
nand U19559 (N_19559,N_16506,N_17985);
nor U19560 (N_19560,N_17213,N_17114);
or U19561 (N_19561,N_16036,N_16259);
and U19562 (N_19562,N_16340,N_16021);
or U19563 (N_19563,N_17473,N_18051);
and U19564 (N_19564,N_17514,N_16197);
nand U19565 (N_19565,N_17063,N_17425);
xnor U19566 (N_19566,N_18332,N_17392);
nand U19567 (N_19567,N_17861,N_16210);
nor U19568 (N_19568,N_16930,N_18488);
nor U19569 (N_19569,N_16486,N_18621);
nor U19570 (N_19570,N_17752,N_16334);
or U19571 (N_19571,N_16850,N_18592);
nor U19572 (N_19572,N_17687,N_16164);
or U19573 (N_19573,N_17374,N_17028);
nor U19574 (N_19574,N_18040,N_18080);
nor U19575 (N_19575,N_17894,N_17460);
and U19576 (N_19576,N_15668,N_18725);
nor U19577 (N_19577,N_17224,N_17795);
nor U19578 (N_19578,N_16270,N_16206);
nand U19579 (N_19579,N_18198,N_16209);
or U19580 (N_19580,N_16854,N_18251);
or U19581 (N_19581,N_18719,N_18707);
or U19582 (N_19582,N_18054,N_17791);
or U19583 (N_19583,N_17179,N_18086);
nor U19584 (N_19584,N_16410,N_15846);
nand U19585 (N_19585,N_16309,N_17286);
nand U19586 (N_19586,N_16708,N_16098);
or U19587 (N_19587,N_18559,N_16452);
xnor U19588 (N_19588,N_17575,N_16996);
nor U19589 (N_19589,N_18634,N_18206);
nor U19590 (N_19590,N_15691,N_17444);
and U19591 (N_19591,N_16726,N_17086);
nor U19592 (N_19592,N_17333,N_17562);
xnor U19593 (N_19593,N_16539,N_16775);
and U19594 (N_19594,N_16760,N_17922);
and U19595 (N_19595,N_17822,N_15720);
nor U19596 (N_19596,N_16585,N_18724);
nand U19597 (N_19597,N_17036,N_17304);
xor U19598 (N_19598,N_16094,N_18591);
nor U19599 (N_19599,N_16832,N_18156);
nand U19600 (N_19600,N_15931,N_18038);
xnor U19601 (N_19601,N_17428,N_16785);
nand U19602 (N_19602,N_16962,N_18631);
xnor U19603 (N_19603,N_16501,N_17310);
nand U19604 (N_19604,N_17744,N_16395);
xor U19605 (N_19605,N_15925,N_17439);
xor U19606 (N_19606,N_18323,N_17742);
nor U19607 (N_19607,N_16654,N_17768);
and U19608 (N_19608,N_17637,N_17324);
nor U19609 (N_19609,N_15830,N_18057);
and U19610 (N_19610,N_17962,N_16151);
nand U19611 (N_19611,N_17314,N_15658);
xor U19612 (N_19612,N_17117,N_17623);
nand U19613 (N_19613,N_18155,N_16034);
nor U19614 (N_19614,N_17185,N_18509);
and U19615 (N_19615,N_18078,N_16757);
and U19616 (N_19616,N_16607,N_16269);
nand U19617 (N_19617,N_18738,N_18499);
nor U19618 (N_19618,N_18581,N_15806);
nand U19619 (N_19619,N_18441,N_17221);
and U19620 (N_19620,N_16295,N_16972);
or U19621 (N_19621,N_16106,N_16176);
nor U19622 (N_19622,N_16250,N_15749);
nand U19623 (N_19623,N_18154,N_16900);
or U19624 (N_19624,N_16175,N_15708);
nand U19625 (N_19625,N_15705,N_16644);
nor U19626 (N_19626,N_18027,N_17678);
and U19627 (N_19627,N_15755,N_16929);
and U19628 (N_19628,N_18558,N_16774);
nand U19629 (N_19629,N_16517,N_18119);
xnor U19630 (N_19630,N_18290,N_18370);
and U19631 (N_19631,N_16889,N_18176);
or U19632 (N_19632,N_18303,N_16284);
nand U19633 (N_19633,N_16194,N_17251);
xnor U19634 (N_19634,N_16541,N_16685);
nor U19635 (N_19635,N_15878,N_17305);
nand U19636 (N_19636,N_16815,N_15903);
and U19637 (N_19637,N_16969,N_17383);
nor U19638 (N_19638,N_15641,N_17551);
or U19639 (N_19639,N_16773,N_15723);
nand U19640 (N_19640,N_17083,N_16544);
nor U19641 (N_19641,N_16709,N_17712);
nand U19642 (N_19642,N_18429,N_17621);
or U19643 (N_19643,N_18677,N_18292);
nand U19644 (N_19644,N_17531,N_17463);
and U19645 (N_19645,N_18541,N_17855);
or U19646 (N_19646,N_18007,N_17348);
nand U19647 (N_19647,N_17157,N_16995);
nand U19648 (N_19648,N_18697,N_18564);
or U19649 (N_19649,N_17477,N_17952);
nand U19650 (N_19650,N_18017,N_16840);
nand U19651 (N_19651,N_17811,N_18098);
nand U19652 (N_19652,N_16614,N_18373);
or U19653 (N_19653,N_16548,N_16909);
and U19654 (N_19654,N_17113,N_18191);
nor U19655 (N_19655,N_16459,N_17358);
and U19656 (N_19656,N_17101,N_16590);
or U19657 (N_19657,N_18656,N_17450);
nor U19658 (N_19658,N_16404,N_16895);
and U19659 (N_19659,N_16927,N_16907);
nor U19660 (N_19660,N_17055,N_16135);
and U19661 (N_19661,N_18280,N_16986);
or U19662 (N_19662,N_16204,N_15762);
nor U19663 (N_19663,N_18583,N_16071);
or U19664 (N_19664,N_16249,N_18282);
xor U19665 (N_19665,N_16332,N_17144);
or U19666 (N_19666,N_16041,N_18430);
and U19667 (N_19667,N_17127,N_15786);
nand U19668 (N_19668,N_18186,N_16053);
and U19669 (N_19669,N_16068,N_16858);
xor U19670 (N_19670,N_18230,N_18340);
nand U19671 (N_19671,N_16324,N_16185);
or U19672 (N_19672,N_16289,N_18507);
and U19673 (N_19673,N_16861,N_17663);
or U19674 (N_19674,N_17676,N_16511);
nand U19675 (N_19675,N_15877,N_16518);
nor U19676 (N_19676,N_18121,N_18743);
nor U19677 (N_19677,N_15894,N_17280);
and U19678 (N_19678,N_15804,N_17454);
or U19679 (N_19679,N_18195,N_16444);
nand U19680 (N_19680,N_16677,N_17749);
or U19681 (N_19681,N_17747,N_18125);
nand U19682 (N_19682,N_17087,N_16810);
or U19683 (N_19683,N_18475,N_17132);
or U19684 (N_19684,N_18649,N_16157);
nand U19685 (N_19685,N_18704,N_18572);
xnor U19686 (N_19686,N_17713,N_18142);
and U19687 (N_19687,N_17810,N_16155);
xor U19688 (N_19688,N_17617,N_18453);
nor U19689 (N_19689,N_15628,N_18468);
nor U19690 (N_19690,N_18020,N_15861);
nand U19691 (N_19691,N_16605,N_16417);
nand U19692 (N_19692,N_17023,N_18477);
nand U19693 (N_19693,N_15924,N_16496);
nor U19694 (N_19694,N_17821,N_16039);
nor U19695 (N_19695,N_15630,N_17553);
or U19696 (N_19696,N_17431,N_16318);
xor U19697 (N_19697,N_16083,N_16772);
and U19698 (N_19698,N_18532,N_18706);
nor U19699 (N_19699,N_18405,N_17569);
and U19700 (N_19700,N_17779,N_18217);
or U19701 (N_19701,N_16485,N_18256);
nor U19702 (N_19702,N_16649,N_17377);
nor U19703 (N_19703,N_18505,N_17580);
nor U19704 (N_19704,N_18544,N_18394);
nand U19705 (N_19705,N_17845,N_16337);
or U19706 (N_19706,N_18353,N_17608);
nor U19707 (N_19707,N_16242,N_17563);
or U19708 (N_19708,N_17529,N_16977);
nor U19709 (N_19709,N_15655,N_17936);
or U19710 (N_19710,N_17386,N_16943);
nor U19711 (N_19711,N_16330,N_17388);
xnor U19712 (N_19712,N_17249,N_15732);
xnor U19713 (N_19713,N_17289,N_16126);
or U19714 (N_19714,N_16132,N_18601);
xor U19715 (N_19715,N_17174,N_16530);
or U19716 (N_19716,N_16796,N_18168);
or U19717 (N_19717,N_18024,N_16645);
nand U19718 (N_19718,N_17145,N_17578);
and U19719 (N_19719,N_16366,N_15676);
and U19720 (N_19720,N_15937,N_16531);
nor U19721 (N_19721,N_16568,N_16592);
or U19722 (N_19722,N_15824,N_16887);
xnor U19723 (N_19723,N_17246,N_16770);
nor U19724 (N_19724,N_18424,N_17682);
or U19725 (N_19725,N_17156,N_17048);
and U19726 (N_19726,N_16172,N_16464);
nor U19727 (N_19727,N_16697,N_17600);
or U19728 (N_19728,N_18481,N_16076);
nand U19729 (N_19729,N_16581,N_15667);
nor U19730 (N_19730,N_16837,N_18516);
xnor U19731 (N_19731,N_16997,N_17745);
nor U19732 (N_19732,N_17254,N_18715);
nand U19733 (N_19733,N_17581,N_16797);
or U19734 (N_19734,N_16316,N_16817);
nand U19735 (N_19735,N_16558,N_18287);
and U19736 (N_19736,N_17505,N_18461);
nor U19737 (N_19737,N_17596,N_17270);
nor U19738 (N_19738,N_16813,N_17823);
nand U19739 (N_19739,N_15951,N_18033);
nor U19740 (N_19740,N_17504,N_16621);
xor U19741 (N_19741,N_17981,N_16089);
and U19742 (N_19742,N_18343,N_15944);
nor U19743 (N_19743,N_16613,N_17648);
and U19744 (N_19744,N_17118,N_15627);
xnor U19745 (N_19745,N_18141,N_18228);
or U19746 (N_19746,N_16963,N_18063);
nor U19747 (N_19747,N_18402,N_16266);
nand U19748 (N_19748,N_16188,N_17094);
or U19749 (N_19749,N_15964,N_15703);
nor U19750 (N_19750,N_16085,N_15789);
and U19751 (N_19751,N_16727,N_17382);
xnor U19752 (N_19752,N_16890,N_17660);
and U19753 (N_19753,N_17550,N_18337);
nand U19754 (N_19754,N_15646,N_18497);
nand U19755 (N_19755,N_16569,N_18435);
xor U19756 (N_19756,N_17138,N_15832);
or U19757 (N_19757,N_18456,N_17338);
nor U19758 (N_19758,N_17182,N_18004);
nand U19759 (N_19759,N_17816,N_16910);
and U19760 (N_19760,N_16512,N_17659);
and U19761 (N_19761,N_18517,N_18204);
nand U19762 (N_19762,N_17885,N_15805);
or U19763 (N_19763,N_17959,N_18682);
xor U19764 (N_19764,N_17956,N_16225);
and U19765 (N_19765,N_17679,N_16055);
nand U19766 (N_19766,N_15939,N_16523);
xor U19767 (N_19767,N_17452,N_16554);
nor U19768 (N_19768,N_17031,N_17497);
or U19769 (N_19769,N_18067,N_16291);
or U19770 (N_19770,N_18487,N_17173);
nand U19771 (N_19771,N_15780,N_17133);
xnor U19772 (N_19772,N_17601,N_17364);
nand U19773 (N_19773,N_17954,N_18036);
nor U19774 (N_19774,N_17020,N_16847);
nand U19775 (N_19775,N_18029,N_16839);
or U19776 (N_19776,N_15754,N_16804);
xnor U19777 (N_19777,N_16272,N_17053);
nor U19778 (N_19778,N_17740,N_16720);
nand U19779 (N_19779,N_17412,N_16964);
xnor U19780 (N_19780,N_16088,N_17839);
or U19781 (N_19781,N_16851,N_16069);
and U19782 (N_19782,N_17856,N_16888);
or U19783 (N_19783,N_17380,N_17891);
xnor U19784 (N_19784,N_18013,N_17034);
or U19785 (N_19785,N_17072,N_17996);
and U19786 (N_19786,N_18611,N_18048);
nor U19787 (N_19787,N_18467,N_18212);
nor U19788 (N_19788,N_16487,N_18266);
or U19789 (N_19789,N_17199,N_15968);
or U19790 (N_19790,N_16562,N_18173);
nor U19791 (N_19791,N_18502,N_17607);
or U19792 (N_19792,N_18491,N_16620);
nor U19793 (N_19793,N_16656,N_17573);
or U19794 (N_19794,N_18399,N_18412);
and U19795 (N_19795,N_16599,N_16594);
xor U19796 (N_19796,N_17825,N_15783);
nand U19797 (N_19797,N_16549,N_18257);
nor U19798 (N_19798,N_17800,N_17681);
xor U19799 (N_19799,N_16665,N_18603);
and U19800 (N_19800,N_15798,N_15856);
nand U19801 (N_19801,N_15633,N_16694);
and U19802 (N_19802,N_17585,N_17137);
xor U19803 (N_19803,N_15858,N_17328);
xnor U19804 (N_19804,N_17195,N_16403);
and U19805 (N_19805,N_16666,N_17705);
and U19806 (N_19806,N_18325,N_18614);
nor U19807 (N_19807,N_16057,N_16800);
or U19808 (N_19808,N_17571,N_18194);
or U19809 (N_19809,N_18296,N_18358);
nor U19810 (N_19810,N_17245,N_18730);
or U19811 (N_19811,N_17881,N_18324);
and U19812 (N_19812,N_18053,N_18039);
nor U19813 (N_19813,N_17066,N_17803);
nand U19814 (N_19814,N_16293,N_18519);
and U19815 (N_19815,N_17366,N_16312);
nor U19816 (N_19816,N_17680,N_17357);
nor U19817 (N_19817,N_15997,N_16509);
and U19818 (N_19818,N_17336,N_16192);
nand U19819 (N_19819,N_17980,N_17641);
and U19820 (N_19820,N_15996,N_16358);
and U19821 (N_19821,N_16115,N_17568);
nor U19822 (N_19822,N_16379,N_16074);
or U19823 (N_19823,N_15649,N_18201);
xnor U19824 (N_19824,N_18177,N_17595);
xnor U19825 (N_19825,N_17253,N_17942);
nor U19826 (N_19826,N_16084,N_15983);
nor U19827 (N_19827,N_15736,N_17059);
or U19828 (N_19828,N_17772,N_17976);
nand U19829 (N_19829,N_18223,N_17724);
and U19830 (N_19830,N_16915,N_17906);
and U19831 (N_19831,N_18448,N_17735);
or U19832 (N_19832,N_17898,N_17006);
or U19833 (N_19833,N_18135,N_17993);
and U19834 (N_19834,N_17146,N_16342);
nand U19835 (N_19835,N_16200,N_18607);
and U19836 (N_19836,N_18276,N_16748);
xnor U19837 (N_19837,N_16636,N_18117);
and U19838 (N_19838,N_18241,N_16221);
nand U19839 (N_19839,N_16019,N_16095);
xor U19840 (N_19840,N_16463,N_16689);
and U19841 (N_19841,N_18484,N_17757);
nand U19842 (N_19842,N_17261,N_18382);
and U19843 (N_19843,N_18666,N_17806);
xnor U19844 (N_19844,N_17870,N_17603);
nand U19845 (N_19845,N_17191,N_18285);
nor U19846 (N_19846,N_18439,N_17079);
nor U19847 (N_19847,N_16824,N_17149);
and U19848 (N_19848,N_17515,N_16152);
and U19849 (N_19849,N_15896,N_18419);
nand U19850 (N_19850,N_17961,N_16478);
xnor U19851 (N_19851,N_16476,N_17330);
or U19852 (N_19852,N_17649,N_18503);
and U19853 (N_19853,N_17009,N_17090);
and U19854 (N_19854,N_16808,N_16516);
xor U19855 (N_19855,N_15715,N_15764);
or U19856 (N_19856,N_16411,N_17739);
or U19857 (N_19857,N_17710,N_17311);
and U19858 (N_19858,N_16826,N_17535);
and U19859 (N_19859,N_16244,N_16173);
and U19860 (N_19860,N_16470,N_15815);
or U19861 (N_19861,N_18450,N_18527);
nor U19862 (N_19862,N_16660,N_17669);
xor U19863 (N_19863,N_17788,N_17901);
nand U19864 (N_19864,N_15664,N_16776);
nor U19865 (N_19865,N_16228,N_15636);
or U19866 (N_19866,N_16786,N_16426);
nor U19867 (N_19867,N_17884,N_16072);
nand U19868 (N_19868,N_16370,N_17187);
or U19869 (N_19869,N_16719,N_16572);
nor U19870 (N_19870,N_17609,N_16934);
nand U19871 (N_19871,N_16988,N_16939);
and U19872 (N_19872,N_16043,N_16846);
and U19873 (N_19873,N_17275,N_18297);
nor U19874 (N_19874,N_18059,N_15690);
xnor U19875 (N_19875,N_17198,N_17860);
xnor U19876 (N_19876,N_18157,N_18259);
xor U19877 (N_19877,N_17148,N_18281);
nor U19878 (N_19878,N_15859,N_16243);
or U19879 (N_19879,N_16985,N_17592);
xor U19880 (N_19880,N_17949,N_16534);
or U19881 (N_19881,N_17248,N_15855);
nor U19882 (N_19882,N_16482,N_16899);
nand U19883 (N_19883,N_18445,N_17647);
nand U19884 (N_19884,N_17091,N_16667);
nand U19885 (N_19885,N_18060,N_18095);
xnor U19886 (N_19886,N_17579,N_16448);
or U19887 (N_19887,N_15677,N_18549);
nor U19888 (N_19888,N_16514,N_15868);
and U19889 (N_19889,N_17405,N_17209);
and U19890 (N_19890,N_18012,N_18529);
or U19891 (N_19891,N_15799,N_18192);
and U19892 (N_19892,N_16746,N_17238);
xnor U19893 (N_19893,N_16317,N_16251);
xor U19894 (N_19894,N_16446,N_17966);
or U19895 (N_19895,N_16732,N_18392);
xnor U19896 (N_19896,N_16522,N_18473);
xnor U19897 (N_19897,N_17872,N_16974);
nor U19898 (N_19898,N_15753,N_17833);
nand U19899 (N_19899,N_17258,N_16235);
xnor U19900 (N_19900,N_18744,N_15884);
nor U19901 (N_19901,N_17287,N_16658);
or U19902 (N_19902,N_17360,N_17886);
nand U19903 (N_19903,N_16761,N_16407);
nor U19904 (N_19904,N_18731,N_16255);
and U19905 (N_19905,N_17190,N_17658);
and U19906 (N_19906,N_18011,N_16186);
xnor U19907 (N_19907,N_16124,N_17105);
nand U19908 (N_19908,N_17893,N_18338);
xor U19909 (N_19909,N_16483,N_17241);
xor U19910 (N_19910,N_15626,N_17354);
and U19911 (N_19911,N_18179,N_16028);
xnor U19912 (N_19912,N_17572,N_16914);
and U19913 (N_19913,N_18321,N_18546);
nor U19914 (N_19914,N_18747,N_17165);
or U19915 (N_19915,N_18378,N_16107);
xnor U19916 (N_19916,N_18403,N_17931);
and U19917 (N_19917,N_16603,N_17994);
and U19918 (N_19918,N_16611,N_17546);
or U19919 (N_19919,N_17988,N_17082);
nor U19920 (N_19920,N_17397,N_15890);
xnor U19921 (N_19921,N_17732,N_18542);
or U19922 (N_19922,N_17472,N_16497);
or U19923 (N_19923,N_17365,N_17470);
and U19924 (N_19924,N_18647,N_15701);
or U19925 (N_19925,N_17734,N_16662);
or U19926 (N_19926,N_17026,N_16722);
or U19927 (N_19927,N_17461,N_18331);
and U19928 (N_19928,N_18339,N_17789);
nor U19929 (N_19929,N_17081,N_17483);
nor U19930 (N_19930,N_17619,N_16116);
xor U19931 (N_19931,N_16828,N_16049);
and U19932 (N_19932,N_17237,N_18407);
nor U19933 (N_19933,N_18478,N_15787);
nor U19934 (N_19934,N_18501,N_16556);
and U19935 (N_19935,N_17722,N_17192);
or U19936 (N_19936,N_15761,N_16067);
and U19937 (N_19937,N_18462,N_17944);
and U19938 (N_19938,N_17189,N_17041);
nand U19939 (N_19939,N_17312,N_16598);
and U19940 (N_19940,N_18215,N_16430);
xnor U19941 (N_19941,N_16778,N_16664);
or U19942 (N_19942,N_15875,N_18246);
nor U19943 (N_19943,N_17998,N_17513);
nand U19944 (N_19944,N_17905,N_17512);
xnor U19945 (N_19945,N_17888,N_17591);
or U19946 (N_19946,N_15709,N_16650);
xor U19947 (N_19947,N_16949,N_17219);
xor U19948 (N_19948,N_16234,N_18397);
or U19949 (N_19949,N_16260,N_16000);
and U19950 (N_19950,N_16524,N_18609);
nor U19951 (N_19951,N_17849,N_18319);
or U19952 (N_19952,N_17152,N_15963);
nand U19953 (N_19953,N_16947,N_16938);
xor U19954 (N_19954,N_15970,N_16093);
xor U19955 (N_19955,N_18349,N_16503);
xor U19956 (N_19956,N_16388,N_16382);
nor U19957 (N_19957,N_18066,N_15848);
or U19958 (N_19958,N_16566,N_18333);
or U19959 (N_19959,N_18152,N_16869);
and U19960 (N_19960,N_16191,N_18092);
xnor U19961 (N_19961,N_18691,N_18474);
or U19962 (N_19962,N_17567,N_16307);
and U19963 (N_19963,N_17001,N_16615);
or U19964 (N_19964,N_17255,N_17820);
and U19965 (N_19965,N_15971,N_18651);
xnor U19966 (N_19966,N_16405,N_16876);
and U19967 (N_19967,N_17691,N_16257);
nor U19968 (N_19968,N_17465,N_17848);
nor U19969 (N_19969,N_15634,N_17095);
xor U19970 (N_19970,N_17624,N_18676);
and U19971 (N_19971,N_16121,N_16451);
or U19972 (N_19972,N_16238,N_18214);
nand U19973 (N_19973,N_17017,N_17818);
nor U19974 (N_19974,N_17807,N_16532);
xnor U19975 (N_19975,N_17702,N_18531);
xor U19976 (N_19976,N_17773,N_16236);
or U19977 (N_19977,N_16149,N_15738);
xnor U19978 (N_19978,N_17052,N_15919);
nor U19979 (N_19979,N_18279,N_18326);
xnor U19980 (N_19980,N_15689,N_16954);
or U19981 (N_19981,N_18485,N_16327);
nand U19982 (N_19982,N_18087,N_16310);
nor U19983 (N_19983,N_15654,N_17697);
nand U19984 (N_19984,N_16536,N_18630);
nand U19985 (N_19985,N_15942,N_17517);
or U19986 (N_19986,N_15852,N_17441);
nor U19987 (N_19987,N_15899,N_17554);
and U19988 (N_19988,N_16771,N_18138);
xnor U19989 (N_19989,N_16860,N_15747);
or U19990 (N_19990,N_18618,N_16367);
nor U19991 (N_19991,N_18624,N_17511);
or U19992 (N_19992,N_17426,N_16288);
xnor U19993 (N_19993,N_18022,N_17925);
xnor U19994 (N_19994,N_17345,N_18381);
nand U19995 (N_19995,N_17701,N_17518);
nor U19996 (N_19996,N_17604,N_17924);
xor U19997 (N_19997,N_16304,N_16984);
xnor U19998 (N_19998,N_18289,N_17853);
and U19999 (N_19999,N_18247,N_17436);
nor U20000 (N_20000,N_16187,N_18147);
xnor U20001 (N_20001,N_18219,N_16435);
nand U20002 (N_20002,N_18045,N_17027);
xor U20003 (N_20003,N_17632,N_17317);
nand U20004 (N_20004,N_16681,N_17398);
or U20005 (N_20005,N_17420,N_18113);
or U20006 (N_20006,N_17864,N_18225);
xor U20007 (N_20007,N_17533,N_18400);
or U20008 (N_20008,N_17927,N_17605);
and U20009 (N_20009,N_16386,N_18598);
and U20010 (N_20010,N_16002,N_15941);
xnor U20011 (N_20011,N_17873,N_18312);
and U20012 (N_20012,N_15953,N_17692);
xnor U20013 (N_20013,N_16230,N_17456);
nand U20014 (N_20014,N_16712,N_17267);
or U20015 (N_20015,N_15713,N_18584);
and U20016 (N_20016,N_18716,N_18262);
nand U20017 (N_20017,N_17755,N_18144);
xnor U20018 (N_20018,N_16134,N_16424);
nor U20019 (N_20019,N_18103,N_18521);
and U20020 (N_20020,N_17123,N_16322);
or U20021 (N_20021,N_17389,N_15625);
xor U20022 (N_20022,N_18272,N_16575);
xor U20023 (N_20023,N_16303,N_17030);
or U20024 (N_20024,N_18126,N_17636);
nand U20025 (N_20025,N_17337,N_15807);
xnor U20026 (N_20026,N_15700,N_16213);
nand U20027 (N_20027,N_18454,N_17858);
nand U20028 (N_20028,N_16510,N_17790);
nor U20029 (N_20029,N_15952,N_16308);
and U20030 (N_20030,N_18622,N_16467);
and U20031 (N_20031,N_16803,N_16742);
nor U20032 (N_20032,N_17344,N_18687);
or U20033 (N_20033,N_17061,N_15743);
and U20034 (N_20034,N_18224,N_18209);
xor U20035 (N_20035,N_15735,N_16389);
or U20036 (N_20036,N_18420,N_17046);
and U20037 (N_20037,N_18623,N_17003);
or U20038 (N_20038,N_17955,N_17545);
xor U20039 (N_20039,N_18574,N_18310);
nor U20040 (N_20040,N_16328,N_17080);
nor U20041 (N_20041,N_18391,N_18563);
nand U20042 (N_20042,N_15972,N_17503);
xnor U20043 (N_20043,N_17373,N_16745);
nor U20044 (N_20044,N_16097,N_18627);
xnor U20045 (N_20045,N_16489,N_16140);
and U20046 (N_20046,N_16805,N_17675);
and U20047 (N_20047,N_17369,N_17150);
nor U20048 (N_20048,N_17443,N_16744);
or U20049 (N_20049,N_15843,N_17496);
nor U20050 (N_20050,N_15906,N_18284);
xor U20051 (N_20051,N_17479,N_15998);
nor U20052 (N_20052,N_17231,N_15930);
xnor U20053 (N_20053,N_16542,N_15965);
xor U20054 (N_20054,N_18278,N_18005);
or U20055 (N_20055,N_16971,N_18680);
nand U20056 (N_20056,N_15947,N_17640);
or U20057 (N_20057,N_15645,N_18702);
xnor U20058 (N_20058,N_15873,N_17564);
nor U20059 (N_20059,N_16638,N_17876);
nor U20060 (N_20060,N_16325,N_16535);
nor U20061 (N_20061,N_17711,N_18515);
and U20062 (N_20062,N_17635,N_17448);
or U20063 (N_20063,N_18547,N_16458);
nand U20064 (N_20064,N_17163,N_17306);
or U20065 (N_20065,N_16789,N_18401);
nor U20066 (N_20066,N_16625,N_16728);
nand U20067 (N_20067,N_18588,N_16263);
or U20068 (N_20068,N_18543,N_18114);
and U20069 (N_20069,N_16751,N_17765);
and U20070 (N_20070,N_18380,N_15742);
and U20071 (N_20071,N_17417,N_17963);
nor U20072 (N_20072,N_17506,N_16529);
nor U20073 (N_20073,N_18520,N_15678);
xnor U20074 (N_20074,N_18210,N_16980);
xor U20075 (N_20075,N_17709,N_16475);
xor U20076 (N_20076,N_18244,N_16205);
or U20077 (N_20077,N_15985,N_16705);
nor U20078 (N_20078,N_15981,N_17170);
or U20079 (N_20079,N_15954,N_15791);
nand U20080 (N_20080,N_18703,N_18235);
and U20081 (N_20081,N_17294,N_17247);
nor U20082 (N_20082,N_15991,N_16526);
and U20083 (N_20083,N_15839,N_16631);
nand U20084 (N_20084,N_15653,N_17865);
nand U20085 (N_20085,N_16750,N_18728);
xor U20086 (N_20086,N_17068,N_16427);
nor U20087 (N_20087,N_17992,N_16734);
and U20088 (N_20088,N_15902,N_17089);
and U20089 (N_20089,N_16190,N_18118);
nand U20090 (N_20090,N_16584,N_17919);
nor U20091 (N_20091,N_15871,N_18745);
and U20092 (N_20092,N_15687,N_18071);
xor U20093 (N_20093,N_15893,N_17244);
nand U20094 (N_20094,N_17391,N_17155);
and U20095 (N_20095,N_17489,N_17673);
xnor U20096 (N_20096,N_18143,N_18460);
and U20097 (N_20097,N_16905,N_17107);
or U20098 (N_20098,N_17696,N_15999);
or U20099 (N_20099,N_18006,N_17638);
and U20100 (N_20100,N_17947,N_17108);
and U20101 (N_20101,N_18620,N_18721);
nand U20102 (N_20102,N_18074,N_16457);
nand U20103 (N_20103,N_15865,N_15665);
and U20104 (N_20104,N_18579,N_17074);
nor U20105 (N_20105,N_16933,N_17556);
xor U20106 (N_20106,N_18084,N_18465);
nor U20107 (N_20107,N_18409,N_16177);
or U20108 (N_20108,N_15726,N_17134);
and U20109 (N_20109,N_18334,N_16911);
or U20110 (N_20110,N_16022,N_16493);
xor U20111 (N_20111,N_15932,N_17353);
nor U20112 (N_20112,N_16099,N_17259);
nor U20113 (N_20113,N_17900,N_17119);
xnor U20114 (N_20114,N_18311,N_15897);
nand U20115 (N_20115,N_17721,N_16935);
nand U20116 (N_20116,N_18432,N_16550);
nor U20117 (N_20117,N_17400,N_18582);
xnor U20118 (N_20118,N_18410,N_16606);
nor U20119 (N_20119,N_17356,N_17206);
and U20120 (N_20120,N_18153,N_15729);
xor U20121 (N_20121,N_18050,N_18203);
nand U20122 (N_20122,N_18000,N_15802);
xnor U20123 (N_20123,N_17207,N_15734);
or U20124 (N_20124,N_18612,N_18375);
xor U20125 (N_20125,N_16879,N_16137);
nand U20126 (N_20126,N_15962,N_15973);
nand U20127 (N_20127,N_18253,N_16704);
and U20128 (N_20128,N_18293,N_16495);
nand U20129 (N_20129,N_16461,N_17708);
or U20130 (N_20130,N_16755,N_18608);
and U20131 (N_20131,N_16499,N_17495);
nor U20132 (N_20132,N_17446,N_18661);
or U20133 (N_20133,N_18652,N_17309);
xnor U20134 (N_20134,N_17559,N_16560);
and U20135 (N_20135,N_16442,N_16675);
or U20136 (N_20136,N_18112,N_17758);
and U20137 (N_20137,N_16217,N_16987);
or U20138 (N_20138,N_18681,N_16222);
nor U20139 (N_20139,N_17220,N_15788);
xnor U20140 (N_20140,N_18354,N_16754);
and U20141 (N_20141,N_16198,N_16133);
or U20142 (N_20142,N_16314,N_18518);
and U20143 (N_20143,N_18352,N_18408);
xor U20144 (N_20144,N_15782,N_18528);
nand U20145 (N_20145,N_16871,N_16555);
xor U20146 (N_20146,N_15714,N_15831);
nor U20147 (N_20147,N_16738,N_17970);
nor U20148 (N_20148,N_16456,N_18166);
or U20149 (N_20149,N_18248,N_17427);
xor U20150 (N_20150,N_17890,N_15949);
and U20151 (N_20151,N_17625,N_16642);
xor U20152 (N_20152,N_18240,N_15838);
and U20153 (N_20153,N_16150,N_18565);
nor U20154 (N_20154,N_17814,N_16345);
nand U20155 (N_20155,N_16597,N_18213);
and U20156 (N_20156,N_18357,N_17869);
nor U20157 (N_20157,N_15794,N_17986);
xnor U20158 (N_20158,N_18540,N_18414);
and U20159 (N_20159,N_16065,N_16056);
nand U20160 (N_20160,N_17243,N_15966);
nand U20161 (N_20161,N_16357,N_16353);
or U20162 (N_20162,N_16399,N_17733);
nor U20163 (N_20163,N_15685,N_16672);
xor U20164 (N_20164,N_17932,N_16374);
xnor U20165 (N_20165,N_18383,N_17000);
nand U20166 (N_20166,N_17421,N_17719);
and U20167 (N_20167,N_17352,N_15670);
xor U20168 (N_20168,N_15640,N_17946);
and U20169 (N_20169,N_16577,N_17498);
nand U20170 (N_20170,N_16468,N_16054);
nor U20171 (N_20171,N_17945,N_15739);
nand U20172 (N_20172,N_15752,N_15659);
or U20173 (N_20173,N_16320,N_18015);
nand U20174 (N_20174,N_16397,N_18668);
or U20175 (N_20175,N_17161,N_17587);
nor U20176 (N_20176,N_17783,N_17759);
nor U20177 (N_20177,N_18025,N_18366);
nand U20178 (N_20178,N_17315,N_16783);
xnor U20179 (N_20179,N_17639,N_18301);
nor U20180 (N_20180,N_16507,N_17476);
nor U20181 (N_20181,N_15781,N_17422);
or U20182 (N_20182,N_17054,N_17320);
xnor U20183 (N_20183,N_16199,N_15987);
nand U20184 (N_20184,N_15768,N_15722);
xor U20185 (N_20185,N_16982,N_16492);
nand U20186 (N_20186,N_16926,N_16973);
or U20187 (N_20187,N_15860,N_18571);
nand U20188 (N_20188,N_18628,N_16591);
or U20189 (N_20189,N_18346,N_15892);
or U20190 (N_20190,N_16351,N_16966);
or U20191 (N_20191,N_16692,N_18653);
or U20192 (N_20192,N_18283,N_16698);
xnor U20193 (N_20193,N_16717,N_17627);
xnor U20194 (N_20194,N_18748,N_18663);
nand U20195 (N_20195,N_17325,N_17867);
nor U20196 (N_20196,N_17442,N_17730);
and U20197 (N_20197,N_16045,N_16052);
and U20198 (N_20198,N_16390,N_16275);
nor U20199 (N_20199,N_16455,N_15741);
or U20200 (N_20200,N_18300,N_16142);
nand U20201 (N_20201,N_16875,N_16104);
and U20202 (N_20202,N_17486,N_18557);
and U20203 (N_20203,N_18093,N_16161);
nand U20204 (N_20204,N_16736,N_15637);
or U20205 (N_20205,N_17433,N_16546);
nor U20206 (N_20206,N_16432,N_16100);
nor U20207 (N_20207,N_17802,N_18404);
xor U20208 (N_20208,N_18593,N_16957);
nor U20209 (N_20209,N_17013,N_16384);
nor U20210 (N_20210,N_15908,N_15651);
or U20211 (N_20211,N_17274,N_18226);
or U20212 (N_20212,N_16481,N_17067);
nand U20213 (N_20213,N_18645,N_18664);
nand U20214 (N_20214,N_16008,N_17871);
and U20215 (N_20215,N_15853,N_17058);
and U20216 (N_20216,N_17889,N_17690);
xnor U20217 (N_20217,N_16305,N_16171);
and U20218 (N_20218,N_16604,N_17468);
or U20219 (N_20219,N_18686,N_18070);
and U20220 (N_20220,N_18538,N_16641);
nor U20221 (N_20221,N_16300,N_16087);
xnor U20222 (N_20222,N_17184,N_16866);
and U20223 (N_20223,N_18181,N_16326);
xnor U20224 (N_20224,N_16989,N_18727);
xnor U20225 (N_20225,N_17284,N_15822);
and U20226 (N_20226,N_16723,N_16981);
xnor U20227 (N_20227,N_15946,N_18277);
and U20228 (N_20228,N_18058,N_16944);
xor U20229 (N_20229,N_16576,N_18606);
xnor U20230 (N_20230,N_15841,N_18533);
and U20231 (N_20231,N_16240,N_18106);
nor U20232 (N_20232,N_16393,N_16471);
nor U20233 (N_20233,N_17447,N_16816);
or U20234 (N_20234,N_17746,N_16741);
and U20235 (N_20235,N_16841,N_17664);
and U20236 (N_20236,N_16333,N_18568);
xnor U20237 (N_20237,N_17370,N_17671);
or U20238 (N_20238,N_17847,N_18295);
nand U20239 (N_20239,N_16168,N_17302);
and U20240 (N_20240,N_15978,N_17896);
or U20241 (N_20241,N_16563,N_16298);
or U20242 (N_20242,N_16691,N_15926);
nor U20243 (N_20243,N_18670,N_17763);
and U20244 (N_20244,N_16246,N_17590);
nand U20245 (N_20245,N_18427,N_18127);
or U20246 (N_20246,N_16026,N_18317);
or U20247 (N_20247,N_17866,N_17536);
or U20248 (N_20248,N_16836,N_17991);
and U20249 (N_20249,N_16020,N_18514);
xor U20250 (N_20250,N_17723,N_17836);
and U20251 (N_20251,N_17262,N_18328);
nor U20252 (N_20252,N_17178,N_16856);
nand U20253 (N_20253,N_18255,N_16968);
xor U20254 (N_20254,N_16612,N_16595);
or U20255 (N_20255,N_17530,N_17543);
xor U20256 (N_20256,N_17780,N_16414);
nand U20257 (N_20257,N_17767,N_18047);
or U20258 (N_20258,N_18097,N_17750);
xor U20259 (N_20259,N_16596,N_18650);
or U20260 (N_20260,N_16752,N_16814);
nor U20261 (N_20261,N_17234,N_17502);
nor U20262 (N_20262,N_18714,N_18660);
nand U20263 (N_20263,N_17501,N_15870);
nor U20264 (N_20264,N_18061,N_17378);
or U20265 (N_20265,N_17672,N_17683);
nand U20266 (N_20266,N_15776,N_17909);
nor U20267 (N_20267,N_17799,N_17964);
nand U20268 (N_20268,N_15928,N_17965);
or U20269 (N_20269,N_18171,N_16018);
xnor U20270 (N_20270,N_16922,N_18032);
or U20271 (N_20271,N_17453,N_17362);
nor U20272 (N_20272,N_18100,N_15774);
and U20273 (N_20273,N_16713,N_17208);
nand U20274 (N_20274,N_16146,N_18049);
or U20275 (N_20275,N_15643,N_17693);
or U20276 (N_20276,N_17923,N_18075);
xor U20277 (N_20277,N_17008,N_18134);
or U20278 (N_20278,N_17140,N_16588);
xnor U20279 (N_20279,N_18348,N_17438);
xor U20280 (N_20280,N_18425,N_18014);
nor U20281 (N_20281,N_16504,N_16394);
and U20282 (N_20282,N_17840,N_16574);
nor U20283 (N_20283,N_16376,N_18646);
and U20284 (N_20284,N_18678,N_16023);
and U20285 (N_20285,N_16932,N_16143);
or U20286 (N_20286,N_15980,N_18268);
nor U20287 (N_20287,N_15959,N_18335);
nor U20288 (N_20288,N_17264,N_16433);
xnor U20289 (N_20289,N_15974,N_17935);
and U20290 (N_20290,N_16077,N_18137);
nand U20291 (N_20291,N_18440,N_16593);
and U20292 (N_20292,N_17957,N_16894);
nor U20293 (N_20293,N_18172,N_18443);
nand U20294 (N_20294,N_17341,N_17958);
and U20295 (N_20295,N_17915,N_18437);
nand U20296 (N_20296,N_18222,N_15845);
or U20297 (N_20297,N_17181,N_18578);
nand U20298 (N_20298,N_16425,N_15671);
nor U20299 (N_20299,N_15803,N_16580);
xnor U20300 (N_20300,N_15632,N_16130);
or U20301 (N_20301,N_15744,N_15960);
xor U20302 (N_20302,N_15922,N_17718);
nand U20303 (N_20303,N_16413,N_18089);
or U20304 (N_20304,N_16538,N_16438);
or U20305 (N_20305,N_18055,N_17797);
or U20306 (N_20306,N_16364,N_17025);
and U20307 (N_20307,N_18573,N_17216);
nor U20308 (N_20308,N_17566,N_18539);
nand U20309 (N_20309,N_17084,N_17547);
xnor U20310 (N_20310,N_17493,N_18636);
nand U20311 (N_20311,N_18711,N_18733);
nor U20312 (N_20312,N_16274,N_15963);
and U20313 (N_20313,N_15865,N_16354);
and U20314 (N_20314,N_17737,N_17132);
and U20315 (N_20315,N_16350,N_18006);
nand U20316 (N_20316,N_16211,N_16131);
and U20317 (N_20317,N_18742,N_17751);
nand U20318 (N_20318,N_16790,N_16647);
xnor U20319 (N_20319,N_16293,N_16378);
nor U20320 (N_20320,N_17359,N_16748);
or U20321 (N_20321,N_17994,N_15801);
xnor U20322 (N_20322,N_18222,N_18059);
and U20323 (N_20323,N_15962,N_18419);
nand U20324 (N_20324,N_15817,N_18728);
or U20325 (N_20325,N_18300,N_16811);
xor U20326 (N_20326,N_16892,N_17697);
nor U20327 (N_20327,N_15962,N_15870);
or U20328 (N_20328,N_18287,N_17852);
or U20329 (N_20329,N_18012,N_16860);
nand U20330 (N_20330,N_17299,N_16001);
nand U20331 (N_20331,N_17730,N_17375);
nand U20332 (N_20332,N_17083,N_17226);
xor U20333 (N_20333,N_17483,N_18086);
or U20334 (N_20334,N_16779,N_16515);
and U20335 (N_20335,N_17258,N_18749);
and U20336 (N_20336,N_18372,N_16519);
or U20337 (N_20337,N_17368,N_16651);
nor U20338 (N_20338,N_18676,N_18555);
nand U20339 (N_20339,N_18530,N_16594);
nor U20340 (N_20340,N_17254,N_15979);
or U20341 (N_20341,N_16825,N_17323);
nand U20342 (N_20342,N_18010,N_18297);
nand U20343 (N_20343,N_16838,N_17680);
xnor U20344 (N_20344,N_16793,N_15657);
or U20345 (N_20345,N_15847,N_17182);
nand U20346 (N_20346,N_17301,N_16067);
and U20347 (N_20347,N_16789,N_16850);
and U20348 (N_20348,N_16467,N_16797);
nor U20349 (N_20349,N_17395,N_18298);
and U20350 (N_20350,N_15730,N_16204);
xnor U20351 (N_20351,N_18316,N_16342);
nand U20352 (N_20352,N_17607,N_16216);
nor U20353 (N_20353,N_18138,N_15929);
and U20354 (N_20354,N_17640,N_18180);
nor U20355 (N_20355,N_16058,N_16950);
xor U20356 (N_20356,N_18470,N_16122);
and U20357 (N_20357,N_15801,N_18674);
and U20358 (N_20358,N_16580,N_17016);
nor U20359 (N_20359,N_17268,N_17995);
nor U20360 (N_20360,N_17805,N_15685);
nor U20361 (N_20361,N_17642,N_17213);
xnor U20362 (N_20362,N_16231,N_18143);
or U20363 (N_20363,N_16198,N_16807);
and U20364 (N_20364,N_16659,N_17309);
xnor U20365 (N_20365,N_16007,N_18591);
nand U20366 (N_20366,N_16984,N_18232);
nand U20367 (N_20367,N_16272,N_15674);
nor U20368 (N_20368,N_15892,N_17383);
or U20369 (N_20369,N_18554,N_18195);
and U20370 (N_20370,N_18320,N_17574);
nand U20371 (N_20371,N_17917,N_17105);
nand U20372 (N_20372,N_15829,N_17997);
nor U20373 (N_20373,N_15928,N_16715);
xnor U20374 (N_20374,N_17018,N_18383);
and U20375 (N_20375,N_16871,N_18189);
xor U20376 (N_20376,N_18684,N_17884);
xnor U20377 (N_20377,N_16953,N_15644);
or U20378 (N_20378,N_16813,N_18124);
nor U20379 (N_20379,N_16441,N_17614);
and U20380 (N_20380,N_17907,N_18644);
or U20381 (N_20381,N_17465,N_16883);
or U20382 (N_20382,N_16033,N_16563);
nor U20383 (N_20383,N_18032,N_17771);
xor U20384 (N_20384,N_17934,N_17001);
xnor U20385 (N_20385,N_16167,N_18692);
nand U20386 (N_20386,N_15661,N_17417);
nor U20387 (N_20387,N_16924,N_18353);
nand U20388 (N_20388,N_15640,N_18503);
and U20389 (N_20389,N_17403,N_17752);
or U20390 (N_20390,N_18698,N_16543);
or U20391 (N_20391,N_15659,N_18391);
or U20392 (N_20392,N_17003,N_16068);
or U20393 (N_20393,N_17845,N_16620);
nand U20394 (N_20394,N_18410,N_16601);
and U20395 (N_20395,N_16910,N_17796);
and U20396 (N_20396,N_18470,N_16098);
xor U20397 (N_20397,N_17323,N_16416);
nor U20398 (N_20398,N_18337,N_16456);
nand U20399 (N_20399,N_17363,N_18292);
and U20400 (N_20400,N_15669,N_18034);
nand U20401 (N_20401,N_18194,N_18092);
xnor U20402 (N_20402,N_18643,N_15952);
and U20403 (N_20403,N_18183,N_17743);
nor U20404 (N_20404,N_18232,N_16271);
nor U20405 (N_20405,N_15998,N_15902);
and U20406 (N_20406,N_17881,N_18106);
and U20407 (N_20407,N_17126,N_18240);
nor U20408 (N_20408,N_16314,N_15746);
nor U20409 (N_20409,N_16437,N_16630);
xnor U20410 (N_20410,N_18543,N_17338);
nand U20411 (N_20411,N_16568,N_17764);
or U20412 (N_20412,N_16369,N_17159);
and U20413 (N_20413,N_16093,N_16749);
nor U20414 (N_20414,N_18440,N_16960);
nor U20415 (N_20415,N_17656,N_17848);
xor U20416 (N_20416,N_18275,N_16756);
nand U20417 (N_20417,N_15869,N_18173);
xor U20418 (N_20418,N_18086,N_16422);
nand U20419 (N_20419,N_18558,N_16459);
nor U20420 (N_20420,N_18514,N_16938);
and U20421 (N_20421,N_18214,N_16439);
or U20422 (N_20422,N_17741,N_15753);
nand U20423 (N_20423,N_16774,N_16050);
nor U20424 (N_20424,N_17602,N_17742);
and U20425 (N_20425,N_16400,N_16978);
or U20426 (N_20426,N_16915,N_15872);
nand U20427 (N_20427,N_17344,N_17355);
nor U20428 (N_20428,N_16116,N_16800);
or U20429 (N_20429,N_15814,N_18360);
nor U20430 (N_20430,N_15760,N_15734);
and U20431 (N_20431,N_16697,N_18434);
nor U20432 (N_20432,N_18002,N_16253);
nor U20433 (N_20433,N_18725,N_15681);
nand U20434 (N_20434,N_15725,N_17382);
xnor U20435 (N_20435,N_18509,N_17087);
xor U20436 (N_20436,N_15643,N_16025);
nand U20437 (N_20437,N_17353,N_17783);
nand U20438 (N_20438,N_18006,N_16453);
nor U20439 (N_20439,N_17954,N_16435);
xnor U20440 (N_20440,N_18262,N_16894);
nand U20441 (N_20441,N_17850,N_15846);
and U20442 (N_20442,N_17603,N_17298);
nand U20443 (N_20443,N_15648,N_15814);
nor U20444 (N_20444,N_16928,N_16772);
or U20445 (N_20445,N_17062,N_16517);
nand U20446 (N_20446,N_16273,N_15657);
nor U20447 (N_20447,N_16080,N_18596);
xor U20448 (N_20448,N_15718,N_17381);
nand U20449 (N_20449,N_18278,N_18509);
nor U20450 (N_20450,N_16071,N_16043);
and U20451 (N_20451,N_16582,N_16550);
xor U20452 (N_20452,N_18167,N_16291);
nor U20453 (N_20453,N_16754,N_17381);
nand U20454 (N_20454,N_16002,N_15915);
xnor U20455 (N_20455,N_16757,N_16731);
and U20456 (N_20456,N_17470,N_18129);
xor U20457 (N_20457,N_18511,N_16360);
nor U20458 (N_20458,N_17636,N_17848);
nor U20459 (N_20459,N_17857,N_18310);
or U20460 (N_20460,N_18281,N_15864);
nor U20461 (N_20461,N_16283,N_18697);
nand U20462 (N_20462,N_15794,N_18120);
nand U20463 (N_20463,N_16292,N_18713);
nand U20464 (N_20464,N_17038,N_17384);
nor U20465 (N_20465,N_17894,N_18711);
or U20466 (N_20466,N_17305,N_18534);
nand U20467 (N_20467,N_16846,N_15789);
and U20468 (N_20468,N_16809,N_17198);
or U20469 (N_20469,N_15799,N_18184);
nand U20470 (N_20470,N_17669,N_17545);
nand U20471 (N_20471,N_15643,N_18687);
and U20472 (N_20472,N_17871,N_16379);
and U20473 (N_20473,N_16644,N_17087);
nand U20474 (N_20474,N_16363,N_15947);
nor U20475 (N_20475,N_15877,N_16751);
or U20476 (N_20476,N_17621,N_16877);
or U20477 (N_20477,N_18471,N_16102);
xnor U20478 (N_20478,N_18120,N_17693);
nand U20479 (N_20479,N_16871,N_18431);
nor U20480 (N_20480,N_18455,N_16832);
nor U20481 (N_20481,N_16411,N_18637);
or U20482 (N_20482,N_17131,N_16201);
nor U20483 (N_20483,N_15755,N_16424);
or U20484 (N_20484,N_18155,N_16731);
or U20485 (N_20485,N_16580,N_18370);
xor U20486 (N_20486,N_16632,N_17497);
nand U20487 (N_20487,N_17640,N_16726);
xor U20488 (N_20488,N_15885,N_16261);
xor U20489 (N_20489,N_18488,N_18629);
nand U20490 (N_20490,N_18562,N_17354);
and U20491 (N_20491,N_17490,N_15893);
nand U20492 (N_20492,N_18550,N_16676);
nor U20493 (N_20493,N_16928,N_17502);
xor U20494 (N_20494,N_18010,N_16896);
nand U20495 (N_20495,N_17482,N_18411);
or U20496 (N_20496,N_18476,N_16101);
nor U20497 (N_20497,N_18346,N_18550);
xor U20498 (N_20498,N_17292,N_17382);
and U20499 (N_20499,N_16748,N_16346);
nor U20500 (N_20500,N_18546,N_16802);
xor U20501 (N_20501,N_16068,N_17644);
nor U20502 (N_20502,N_18564,N_18600);
xor U20503 (N_20503,N_17826,N_16321);
or U20504 (N_20504,N_16141,N_16887);
nand U20505 (N_20505,N_18393,N_15805);
or U20506 (N_20506,N_16078,N_16496);
and U20507 (N_20507,N_18368,N_18391);
nor U20508 (N_20508,N_18124,N_16434);
xnor U20509 (N_20509,N_16906,N_15784);
and U20510 (N_20510,N_16666,N_16727);
xor U20511 (N_20511,N_17812,N_15729);
and U20512 (N_20512,N_17875,N_16720);
xor U20513 (N_20513,N_16126,N_18748);
nand U20514 (N_20514,N_16606,N_16719);
and U20515 (N_20515,N_18239,N_16211);
and U20516 (N_20516,N_18638,N_17400);
and U20517 (N_20517,N_16406,N_16947);
xor U20518 (N_20518,N_16030,N_18244);
nor U20519 (N_20519,N_15942,N_15809);
or U20520 (N_20520,N_16689,N_16876);
xnor U20521 (N_20521,N_17056,N_18458);
xnor U20522 (N_20522,N_18081,N_16408);
nand U20523 (N_20523,N_17118,N_18739);
nor U20524 (N_20524,N_17888,N_16203);
and U20525 (N_20525,N_17154,N_18165);
nand U20526 (N_20526,N_16255,N_16504);
or U20527 (N_20527,N_18250,N_18262);
nor U20528 (N_20528,N_18342,N_16309);
and U20529 (N_20529,N_17625,N_16074);
nand U20530 (N_20530,N_16426,N_18653);
nor U20531 (N_20531,N_18625,N_16854);
nand U20532 (N_20532,N_15800,N_16956);
xor U20533 (N_20533,N_16694,N_17214);
and U20534 (N_20534,N_17312,N_18238);
or U20535 (N_20535,N_16126,N_15751);
nor U20536 (N_20536,N_16822,N_18240);
xor U20537 (N_20537,N_17576,N_17647);
or U20538 (N_20538,N_18114,N_18047);
and U20539 (N_20539,N_16729,N_17874);
nand U20540 (N_20540,N_18723,N_17298);
nor U20541 (N_20541,N_17268,N_16909);
or U20542 (N_20542,N_17401,N_17047);
and U20543 (N_20543,N_18682,N_16840);
and U20544 (N_20544,N_18523,N_16896);
nor U20545 (N_20545,N_17443,N_16393);
xor U20546 (N_20546,N_18583,N_15856);
nand U20547 (N_20547,N_16649,N_16997);
nor U20548 (N_20548,N_17123,N_16386);
xor U20549 (N_20549,N_18152,N_16023);
nand U20550 (N_20550,N_16461,N_16732);
or U20551 (N_20551,N_18477,N_18591);
xor U20552 (N_20552,N_18156,N_16045);
nor U20553 (N_20553,N_18592,N_16586);
and U20554 (N_20554,N_16506,N_17492);
xnor U20555 (N_20555,N_16563,N_17131);
and U20556 (N_20556,N_15957,N_17291);
nand U20557 (N_20557,N_18449,N_17625);
nand U20558 (N_20558,N_17016,N_17356);
or U20559 (N_20559,N_18191,N_17706);
xnor U20560 (N_20560,N_17869,N_16338);
and U20561 (N_20561,N_17687,N_18740);
and U20562 (N_20562,N_17866,N_16040);
xnor U20563 (N_20563,N_16849,N_18296);
xnor U20564 (N_20564,N_18663,N_17274);
or U20565 (N_20565,N_16594,N_17889);
nand U20566 (N_20566,N_16738,N_16401);
nor U20567 (N_20567,N_18510,N_17103);
and U20568 (N_20568,N_15901,N_17786);
xnor U20569 (N_20569,N_17051,N_15668);
nor U20570 (N_20570,N_15873,N_15701);
or U20571 (N_20571,N_16254,N_17571);
nand U20572 (N_20572,N_16862,N_18164);
and U20573 (N_20573,N_18580,N_16400);
and U20574 (N_20574,N_15998,N_15845);
or U20575 (N_20575,N_16933,N_17935);
nor U20576 (N_20576,N_17486,N_16212);
or U20577 (N_20577,N_16615,N_17464);
nand U20578 (N_20578,N_17055,N_17516);
or U20579 (N_20579,N_18456,N_16913);
and U20580 (N_20580,N_17131,N_17444);
xnor U20581 (N_20581,N_17822,N_17589);
or U20582 (N_20582,N_18303,N_18169);
and U20583 (N_20583,N_17792,N_15959);
and U20584 (N_20584,N_15883,N_18577);
and U20585 (N_20585,N_18429,N_17815);
nand U20586 (N_20586,N_16122,N_16110);
nand U20587 (N_20587,N_18541,N_16433);
xnor U20588 (N_20588,N_17214,N_18185);
nand U20589 (N_20589,N_16682,N_16120);
xnor U20590 (N_20590,N_17049,N_17822);
and U20591 (N_20591,N_17375,N_18264);
and U20592 (N_20592,N_15888,N_15940);
or U20593 (N_20593,N_18520,N_15800);
xor U20594 (N_20594,N_16098,N_18626);
xor U20595 (N_20595,N_17364,N_15814);
xnor U20596 (N_20596,N_16310,N_16482);
or U20597 (N_20597,N_16276,N_17627);
nand U20598 (N_20598,N_16248,N_16804);
nand U20599 (N_20599,N_15847,N_16924);
and U20600 (N_20600,N_16607,N_18656);
and U20601 (N_20601,N_16051,N_17210);
nand U20602 (N_20602,N_16922,N_18593);
and U20603 (N_20603,N_17804,N_17447);
or U20604 (N_20604,N_17297,N_18103);
nand U20605 (N_20605,N_18179,N_17360);
nor U20606 (N_20606,N_17722,N_18415);
nor U20607 (N_20607,N_15973,N_16200);
nor U20608 (N_20608,N_17977,N_16828);
and U20609 (N_20609,N_16510,N_16648);
or U20610 (N_20610,N_17813,N_16790);
or U20611 (N_20611,N_18026,N_16514);
and U20612 (N_20612,N_16222,N_17992);
xnor U20613 (N_20613,N_18547,N_17083);
nor U20614 (N_20614,N_16461,N_16816);
xor U20615 (N_20615,N_16418,N_17859);
or U20616 (N_20616,N_17063,N_18715);
nor U20617 (N_20617,N_16525,N_17127);
or U20618 (N_20618,N_17745,N_16746);
and U20619 (N_20619,N_15797,N_17321);
or U20620 (N_20620,N_16490,N_16110);
and U20621 (N_20621,N_17181,N_16395);
and U20622 (N_20622,N_18083,N_17700);
and U20623 (N_20623,N_16110,N_17464);
nor U20624 (N_20624,N_16949,N_17461);
and U20625 (N_20625,N_17174,N_17874);
and U20626 (N_20626,N_17874,N_17248);
xnor U20627 (N_20627,N_15753,N_17752);
nor U20628 (N_20628,N_16460,N_18662);
or U20629 (N_20629,N_16194,N_18425);
xnor U20630 (N_20630,N_16912,N_15631);
and U20631 (N_20631,N_16702,N_15638);
nor U20632 (N_20632,N_18095,N_16149);
and U20633 (N_20633,N_16813,N_15687);
xnor U20634 (N_20634,N_16014,N_15907);
nor U20635 (N_20635,N_17740,N_17216);
or U20636 (N_20636,N_17585,N_16762);
or U20637 (N_20637,N_17867,N_15771);
nand U20638 (N_20638,N_16585,N_16348);
nand U20639 (N_20639,N_17543,N_17690);
nand U20640 (N_20640,N_15779,N_17151);
or U20641 (N_20641,N_17879,N_16552);
xnor U20642 (N_20642,N_16215,N_18032);
or U20643 (N_20643,N_17374,N_17893);
or U20644 (N_20644,N_18410,N_17891);
and U20645 (N_20645,N_16560,N_17427);
nand U20646 (N_20646,N_16809,N_16416);
and U20647 (N_20647,N_16753,N_16388);
nor U20648 (N_20648,N_16671,N_16596);
or U20649 (N_20649,N_16529,N_17607);
xor U20650 (N_20650,N_18299,N_18252);
nor U20651 (N_20651,N_16199,N_16357);
nand U20652 (N_20652,N_17515,N_16696);
and U20653 (N_20653,N_17817,N_16713);
or U20654 (N_20654,N_17280,N_18186);
nor U20655 (N_20655,N_16203,N_18639);
nand U20656 (N_20656,N_16966,N_17701);
nand U20657 (N_20657,N_17305,N_16778);
nand U20658 (N_20658,N_17568,N_18443);
or U20659 (N_20659,N_17620,N_17308);
or U20660 (N_20660,N_17805,N_17811);
and U20661 (N_20661,N_18061,N_16618);
or U20662 (N_20662,N_17570,N_17295);
xnor U20663 (N_20663,N_15887,N_18016);
nand U20664 (N_20664,N_16974,N_17730);
nor U20665 (N_20665,N_15846,N_18705);
and U20666 (N_20666,N_18265,N_17031);
or U20667 (N_20667,N_16483,N_18175);
and U20668 (N_20668,N_18491,N_17170);
and U20669 (N_20669,N_17314,N_17132);
nand U20670 (N_20670,N_15663,N_16539);
and U20671 (N_20671,N_18598,N_17874);
and U20672 (N_20672,N_15681,N_16639);
nor U20673 (N_20673,N_17444,N_17279);
nor U20674 (N_20674,N_17450,N_16579);
or U20675 (N_20675,N_18428,N_18443);
xnor U20676 (N_20676,N_16454,N_16769);
nor U20677 (N_20677,N_18310,N_18153);
nand U20678 (N_20678,N_18660,N_18423);
xor U20679 (N_20679,N_17491,N_17847);
or U20680 (N_20680,N_18479,N_16884);
and U20681 (N_20681,N_17008,N_18526);
nand U20682 (N_20682,N_16546,N_18473);
and U20683 (N_20683,N_16748,N_17856);
or U20684 (N_20684,N_17832,N_18349);
or U20685 (N_20685,N_15661,N_16911);
nand U20686 (N_20686,N_18522,N_17466);
nand U20687 (N_20687,N_17626,N_16298);
xor U20688 (N_20688,N_16876,N_17210);
nor U20689 (N_20689,N_18029,N_18068);
xnor U20690 (N_20690,N_15955,N_18212);
nand U20691 (N_20691,N_16855,N_18662);
or U20692 (N_20692,N_17867,N_18196);
or U20693 (N_20693,N_15670,N_17662);
or U20694 (N_20694,N_17526,N_17424);
and U20695 (N_20695,N_16033,N_18708);
and U20696 (N_20696,N_16530,N_16528);
and U20697 (N_20697,N_17292,N_17865);
nor U20698 (N_20698,N_17897,N_16911);
and U20699 (N_20699,N_17321,N_15805);
xor U20700 (N_20700,N_17662,N_18054);
xor U20701 (N_20701,N_15667,N_18062);
nor U20702 (N_20702,N_16132,N_16235);
or U20703 (N_20703,N_16124,N_18566);
nor U20704 (N_20704,N_15697,N_17370);
nand U20705 (N_20705,N_16381,N_16123);
nand U20706 (N_20706,N_16432,N_16229);
nand U20707 (N_20707,N_17180,N_16202);
nor U20708 (N_20708,N_15806,N_16301);
nor U20709 (N_20709,N_17471,N_17968);
and U20710 (N_20710,N_17846,N_17344);
xnor U20711 (N_20711,N_17181,N_15974);
nand U20712 (N_20712,N_18560,N_15785);
nor U20713 (N_20713,N_18257,N_16844);
and U20714 (N_20714,N_15850,N_17211);
nand U20715 (N_20715,N_18519,N_15831);
and U20716 (N_20716,N_17046,N_15910);
and U20717 (N_20717,N_15657,N_16270);
nor U20718 (N_20718,N_17989,N_16943);
or U20719 (N_20719,N_17387,N_18050);
nand U20720 (N_20720,N_18658,N_17937);
or U20721 (N_20721,N_17121,N_16928);
or U20722 (N_20722,N_15917,N_16247);
xnor U20723 (N_20723,N_15755,N_18012);
xnor U20724 (N_20724,N_17412,N_16655);
nand U20725 (N_20725,N_16055,N_18382);
xor U20726 (N_20726,N_17514,N_17654);
and U20727 (N_20727,N_18076,N_15933);
and U20728 (N_20728,N_18353,N_17014);
or U20729 (N_20729,N_16923,N_17896);
or U20730 (N_20730,N_16935,N_17162);
xnor U20731 (N_20731,N_17126,N_16803);
or U20732 (N_20732,N_15882,N_17307);
and U20733 (N_20733,N_18214,N_16786);
nor U20734 (N_20734,N_18728,N_18372);
nand U20735 (N_20735,N_16653,N_18204);
and U20736 (N_20736,N_16143,N_17158);
or U20737 (N_20737,N_15968,N_17284);
nand U20738 (N_20738,N_17858,N_16103);
nor U20739 (N_20739,N_16685,N_16137);
or U20740 (N_20740,N_17805,N_18461);
nor U20741 (N_20741,N_17683,N_17418);
nand U20742 (N_20742,N_18424,N_17377);
or U20743 (N_20743,N_16677,N_16228);
xor U20744 (N_20744,N_15770,N_17341);
nor U20745 (N_20745,N_16521,N_17533);
or U20746 (N_20746,N_18350,N_15916);
and U20747 (N_20747,N_17353,N_17995);
nor U20748 (N_20748,N_17779,N_16009);
xnor U20749 (N_20749,N_17301,N_16245);
or U20750 (N_20750,N_16063,N_17247);
or U20751 (N_20751,N_16736,N_18608);
xnor U20752 (N_20752,N_18391,N_16869);
nor U20753 (N_20753,N_18323,N_18056);
nor U20754 (N_20754,N_16668,N_16527);
nor U20755 (N_20755,N_15655,N_16142);
nand U20756 (N_20756,N_16076,N_17311);
or U20757 (N_20757,N_16923,N_16173);
xnor U20758 (N_20758,N_18030,N_18490);
nor U20759 (N_20759,N_16955,N_17778);
or U20760 (N_20760,N_16589,N_15827);
nor U20761 (N_20761,N_17606,N_16882);
and U20762 (N_20762,N_17375,N_16205);
nand U20763 (N_20763,N_17418,N_15886);
xor U20764 (N_20764,N_15723,N_17124);
xor U20765 (N_20765,N_17869,N_16098);
xor U20766 (N_20766,N_17953,N_17064);
xnor U20767 (N_20767,N_16207,N_16837);
and U20768 (N_20768,N_18199,N_16039);
xor U20769 (N_20769,N_18099,N_17675);
and U20770 (N_20770,N_17096,N_18606);
nor U20771 (N_20771,N_17608,N_15674);
xor U20772 (N_20772,N_18716,N_17351);
and U20773 (N_20773,N_17237,N_16185);
and U20774 (N_20774,N_18672,N_18007);
nand U20775 (N_20775,N_16712,N_17146);
or U20776 (N_20776,N_18432,N_17522);
or U20777 (N_20777,N_15862,N_16047);
nand U20778 (N_20778,N_15877,N_16354);
or U20779 (N_20779,N_17484,N_17318);
nand U20780 (N_20780,N_15863,N_18590);
or U20781 (N_20781,N_18353,N_17412);
and U20782 (N_20782,N_18373,N_16622);
and U20783 (N_20783,N_18654,N_16366);
nor U20784 (N_20784,N_17453,N_16246);
xor U20785 (N_20785,N_16473,N_18401);
nor U20786 (N_20786,N_17329,N_17699);
nor U20787 (N_20787,N_17194,N_17939);
and U20788 (N_20788,N_16491,N_18432);
or U20789 (N_20789,N_18692,N_16739);
or U20790 (N_20790,N_17684,N_18625);
and U20791 (N_20791,N_16100,N_17867);
nand U20792 (N_20792,N_16035,N_16648);
or U20793 (N_20793,N_17586,N_16385);
and U20794 (N_20794,N_17752,N_18289);
nand U20795 (N_20795,N_15675,N_17199);
or U20796 (N_20796,N_16626,N_16999);
nor U20797 (N_20797,N_16208,N_16590);
xnor U20798 (N_20798,N_18207,N_17488);
or U20799 (N_20799,N_16833,N_16130);
nand U20800 (N_20800,N_16598,N_17534);
nor U20801 (N_20801,N_17473,N_18492);
nand U20802 (N_20802,N_17771,N_17201);
or U20803 (N_20803,N_17018,N_17494);
nor U20804 (N_20804,N_17708,N_17473);
nor U20805 (N_20805,N_16970,N_16802);
nand U20806 (N_20806,N_17496,N_16370);
or U20807 (N_20807,N_18641,N_16594);
and U20808 (N_20808,N_15687,N_18747);
nor U20809 (N_20809,N_17414,N_18736);
and U20810 (N_20810,N_18520,N_18726);
nor U20811 (N_20811,N_17016,N_16690);
or U20812 (N_20812,N_17079,N_18165);
nor U20813 (N_20813,N_16386,N_17633);
and U20814 (N_20814,N_18015,N_17213);
or U20815 (N_20815,N_16218,N_17751);
nor U20816 (N_20816,N_18575,N_17867);
or U20817 (N_20817,N_16821,N_18076);
xor U20818 (N_20818,N_15792,N_17623);
nand U20819 (N_20819,N_17952,N_17723);
nand U20820 (N_20820,N_17131,N_17453);
nand U20821 (N_20821,N_15639,N_18727);
or U20822 (N_20822,N_18563,N_16935);
and U20823 (N_20823,N_18237,N_18196);
xnor U20824 (N_20824,N_18193,N_16055);
xnor U20825 (N_20825,N_16532,N_15678);
or U20826 (N_20826,N_17803,N_18084);
nor U20827 (N_20827,N_16608,N_18237);
xor U20828 (N_20828,N_17664,N_18729);
or U20829 (N_20829,N_18121,N_16393);
or U20830 (N_20830,N_18373,N_18202);
nor U20831 (N_20831,N_16477,N_17332);
or U20832 (N_20832,N_16533,N_16997);
nand U20833 (N_20833,N_17318,N_18641);
and U20834 (N_20834,N_16194,N_16192);
or U20835 (N_20835,N_17700,N_18454);
nor U20836 (N_20836,N_17072,N_17124);
xnor U20837 (N_20837,N_16153,N_17397);
nor U20838 (N_20838,N_16898,N_18744);
and U20839 (N_20839,N_15986,N_17381);
xnor U20840 (N_20840,N_17947,N_18148);
nand U20841 (N_20841,N_16773,N_15976);
or U20842 (N_20842,N_16458,N_17952);
or U20843 (N_20843,N_16537,N_17124);
or U20844 (N_20844,N_17477,N_18520);
or U20845 (N_20845,N_15952,N_15742);
xnor U20846 (N_20846,N_18734,N_17450);
xnor U20847 (N_20847,N_15915,N_18011);
nand U20848 (N_20848,N_18391,N_16719);
and U20849 (N_20849,N_17871,N_16260);
or U20850 (N_20850,N_16032,N_17930);
and U20851 (N_20851,N_17319,N_17589);
and U20852 (N_20852,N_16666,N_17651);
nand U20853 (N_20853,N_16401,N_15748);
nand U20854 (N_20854,N_16229,N_17838);
xnor U20855 (N_20855,N_18681,N_16262);
nor U20856 (N_20856,N_18230,N_17915);
or U20857 (N_20857,N_16016,N_16079);
nand U20858 (N_20858,N_16189,N_15957);
xnor U20859 (N_20859,N_16656,N_15876);
xor U20860 (N_20860,N_17088,N_16973);
nor U20861 (N_20861,N_18418,N_17909);
or U20862 (N_20862,N_16471,N_16395);
or U20863 (N_20863,N_17338,N_16864);
and U20864 (N_20864,N_18464,N_18664);
nand U20865 (N_20865,N_17015,N_17569);
and U20866 (N_20866,N_18286,N_16857);
and U20867 (N_20867,N_17663,N_17846);
or U20868 (N_20868,N_15764,N_15917);
nand U20869 (N_20869,N_17392,N_18197);
nand U20870 (N_20870,N_16086,N_17502);
nor U20871 (N_20871,N_17978,N_18119);
xnor U20872 (N_20872,N_17707,N_17377);
xor U20873 (N_20873,N_16514,N_17055);
nor U20874 (N_20874,N_16096,N_17593);
and U20875 (N_20875,N_18006,N_15892);
nand U20876 (N_20876,N_17010,N_18086);
or U20877 (N_20877,N_16177,N_17279);
nor U20878 (N_20878,N_18448,N_18653);
nand U20879 (N_20879,N_18052,N_17231);
or U20880 (N_20880,N_17478,N_17535);
xnor U20881 (N_20881,N_16542,N_17606);
nor U20882 (N_20882,N_18119,N_16356);
or U20883 (N_20883,N_16182,N_16380);
nand U20884 (N_20884,N_18059,N_17931);
or U20885 (N_20885,N_16471,N_16310);
or U20886 (N_20886,N_18499,N_17664);
or U20887 (N_20887,N_17835,N_18278);
nor U20888 (N_20888,N_16671,N_18404);
and U20889 (N_20889,N_15691,N_17420);
nor U20890 (N_20890,N_16485,N_17117);
and U20891 (N_20891,N_16162,N_18667);
nor U20892 (N_20892,N_16633,N_16701);
nor U20893 (N_20893,N_17943,N_18014);
nand U20894 (N_20894,N_17883,N_16858);
or U20895 (N_20895,N_18150,N_18556);
or U20896 (N_20896,N_16224,N_17125);
and U20897 (N_20897,N_17787,N_17186);
nand U20898 (N_20898,N_17115,N_17618);
nand U20899 (N_20899,N_16883,N_17583);
xor U20900 (N_20900,N_18456,N_15763);
xnor U20901 (N_20901,N_16877,N_17190);
or U20902 (N_20902,N_17832,N_15816);
and U20903 (N_20903,N_16477,N_16269);
nor U20904 (N_20904,N_18631,N_16861);
or U20905 (N_20905,N_16469,N_17405);
nand U20906 (N_20906,N_15659,N_15941);
and U20907 (N_20907,N_16791,N_15660);
and U20908 (N_20908,N_16639,N_16419);
or U20909 (N_20909,N_16018,N_16550);
or U20910 (N_20910,N_18378,N_16356);
or U20911 (N_20911,N_17929,N_18584);
nand U20912 (N_20912,N_18621,N_16853);
nor U20913 (N_20913,N_15673,N_16924);
or U20914 (N_20914,N_17625,N_15742);
nor U20915 (N_20915,N_17033,N_17769);
nor U20916 (N_20916,N_16142,N_18567);
xnor U20917 (N_20917,N_17009,N_17127);
or U20918 (N_20918,N_18527,N_16502);
nand U20919 (N_20919,N_17650,N_18311);
nor U20920 (N_20920,N_18188,N_17011);
xor U20921 (N_20921,N_18057,N_16942);
or U20922 (N_20922,N_18100,N_18227);
nor U20923 (N_20923,N_15763,N_16694);
or U20924 (N_20924,N_18512,N_17771);
nor U20925 (N_20925,N_17557,N_18257);
xor U20926 (N_20926,N_17468,N_16537);
xnor U20927 (N_20927,N_17145,N_18229);
or U20928 (N_20928,N_17714,N_16682);
nor U20929 (N_20929,N_16628,N_16427);
or U20930 (N_20930,N_18494,N_17501);
xnor U20931 (N_20931,N_15638,N_18032);
xor U20932 (N_20932,N_18236,N_15961);
and U20933 (N_20933,N_16299,N_16880);
and U20934 (N_20934,N_18510,N_17645);
nand U20935 (N_20935,N_17668,N_18495);
nand U20936 (N_20936,N_16216,N_15714);
xor U20937 (N_20937,N_15724,N_18593);
nand U20938 (N_20938,N_16731,N_15907);
nor U20939 (N_20939,N_16031,N_17837);
nand U20940 (N_20940,N_16763,N_16918);
and U20941 (N_20941,N_18229,N_17610);
nand U20942 (N_20942,N_16144,N_16602);
nor U20943 (N_20943,N_15987,N_18143);
xor U20944 (N_20944,N_17805,N_17461);
and U20945 (N_20945,N_17402,N_16260);
or U20946 (N_20946,N_16403,N_18511);
or U20947 (N_20947,N_16716,N_18605);
or U20948 (N_20948,N_16490,N_16240);
and U20949 (N_20949,N_18413,N_17457);
or U20950 (N_20950,N_16664,N_18038);
nor U20951 (N_20951,N_17277,N_17698);
nor U20952 (N_20952,N_16242,N_15882);
nor U20953 (N_20953,N_16264,N_16418);
and U20954 (N_20954,N_18387,N_15986);
nor U20955 (N_20955,N_15791,N_17399);
nor U20956 (N_20956,N_16404,N_18092);
nor U20957 (N_20957,N_18146,N_16132);
or U20958 (N_20958,N_15786,N_17848);
xnor U20959 (N_20959,N_16183,N_16938);
or U20960 (N_20960,N_15692,N_17649);
and U20961 (N_20961,N_17727,N_17229);
nand U20962 (N_20962,N_17936,N_17422);
xor U20963 (N_20963,N_18538,N_17042);
or U20964 (N_20964,N_18419,N_17435);
nand U20965 (N_20965,N_17615,N_17803);
or U20966 (N_20966,N_17440,N_16459);
xor U20967 (N_20967,N_16768,N_16828);
and U20968 (N_20968,N_17221,N_18374);
nand U20969 (N_20969,N_16220,N_18548);
and U20970 (N_20970,N_17622,N_17020);
nor U20971 (N_20971,N_16311,N_16902);
and U20972 (N_20972,N_18444,N_18570);
nand U20973 (N_20973,N_15981,N_15901);
or U20974 (N_20974,N_16087,N_18691);
xnor U20975 (N_20975,N_18736,N_18662);
xnor U20976 (N_20976,N_18086,N_17131);
nand U20977 (N_20977,N_16936,N_16594);
nand U20978 (N_20978,N_17261,N_17781);
nand U20979 (N_20979,N_17751,N_17266);
or U20980 (N_20980,N_16311,N_18739);
or U20981 (N_20981,N_17510,N_17025);
or U20982 (N_20982,N_17512,N_15779);
or U20983 (N_20983,N_17048,N_15837);
nand U20984 (N_20984,N_15768,N_17241);
nor U20985 (N_20985,N_18526,N_17445);
xnor U20986 (N_20986,N_17235,N_16577);
xor U20987 (N_20987,N_16394,N_18478);
xnor U20988 (N_20988,N_18094,N_16112);
or U20989 (N_20989,N_15877,N_16170);
nand U20990 (N_20990,N_17126,N_16488);
xor U20991 (N_20991,N_17878,N_15655);
nand U20992 (N_20992,N_15862,N_16582);
xor U20993 (N_20993,N_16065,N_16724);
nor U20994 (N_20994,N_17256,N_15711);
nor U20995 (N_20995,N_17748,N_16248);
nor U20996 (N_20996,N_17440,N_17229);
or U20997 (N_20997,N_16308,N_16780);
nand U20998 (N_20998,N_16295,N_18677);
or U20999 (N_20999,N_16815,N_18400);
nand U21000 (N_21000,N_16080,N_17293);
nand U21001 (N_21001,N_16329,N_15702);
nand U21002 (N_21002,N_15683,N_17930);
nand U21003 (N_21003,N_18351,N_18581);
xor U21004 (N_21004,N_16608,N_16794);
nand U21005 (N_21005,N_18197,N_17420);
nand U21006 (N_21006,N_16739,N_18111);
or U21007 (N_21007,N_18083,N_16876);
or U21008 (N_21008,N_17627,N_18503);
nor U21009 (N_21009,N_15939,N_17542);
nand U21010 (N_21010,N_17826,N_17304);
xor U21011 (N_21011,N_18409,N_18514);
xnor U21012 (N_21012,N_16018,N_16706);
or U21013 (N_21013,N_17105,N_17291);
and U21014 (N_21014,N_15711,N_17480);
nor U21015 (N_21015,N_17677,N_16009);
xor U21016 (N_21016,N_17528,N_17156);
xor U21017 (N_21017,N_16853,N_17971);
or U21018 (N_21018,N_17629,N_17818);
xnor U21019 (N_21019,N_17764,N_17798);
nor U21020 (N_21020,N_16855,N_16630);
and U21021 (N_21021,N_17826,N_18525);
or U21022 (N_21022,N_15905,N_16815);
and U21023 (N_21023,N_18335,N_18583);
nor U21024 (N_21024,N_17791,N_16525);
or U21025 (N_21025,N_16925,N_15985);
and U21026 (N_21026,N_18391,N_17699);
xnor U21027 (N_21027,N_16361,N_16586);
xor U21028 (N_21028,N_16491,N_17778);
or U21029 (N_21029,N_17929,N_18399);
and U21030 (N_21030,N_18431,N_17589);
nand U21031 (N_21031,N_18747,N_17533);
or U21032 (N_21032,N_16397,N_17909);
and U21033 (N_21033,N_15751,N_17510);
or U21034 (N_21034,N_17389,N_17653);
xnor U21035 (N_21035,N_16213,N_18041);
xor U21036 (N_21036,N_18353,N_17184);
or U21037 (N_21037,N_17841,N_18011);
and U21038 (N_21038,N_15767,N_16142);
or U21039 (N_21039,N_17779,N_17103);
or U21040 (N_21040,N_15971,N_16574);
or U21041 (N_21041,N_17639,N_18157);
or U21042 (N_21042,N_17270,N_16472);
and U21043 (N_21043,N_18302,N_17526);
nor U21044 (N_21044,N_16372,N_16648);
xor U21045 (N_21045,N_18556,N_16383);
or U21046 (N_21046,N_15930,N_18102);
xnor U21047 (N_21047,N_16773,N_16414);
and U21048 (N_21048,N_16116,N_16371);
nand U21049 (N_21049,N_15902,N_17941);
xnor U21050 (N_21050,N_17925,N_17685);
xor U21051 (N_21051,N_18040,N_15789);
nand U21052 (N_21052,N_18551,N_16346);
nor U21053 (N_21053,N_18623,N_16014);
xor U21054 (N_21054,N_17315,N_17030);
nor U21055 (N_21055,N_18495,N_17720);
xnor U21056 (N_21056,N_17712,N_17832);
nor U21057 (N_21057,N_17955,N_16578);
xnor U21058 (N_21058,N_17559,N_18063);
nand U21059 (N_21059,N_17662,N_17050);
or U21060 (N_21060,N_18709,N_16127);
nor U21061 (N_21061,N_17519,N_17571);
and U21062 (N_21062,N_16499,N_18016);
nor U21063 (N_21063,N_18324,N_16824);
or U21064 (N_21064,N_17699,N_18649);
nor U21065 (N_21065,N_18219,N_16934);
xor U21066 (N_21066,N_15639,N_18020);
nor U21067 (N_21067,N_18063,N_16500);
nand U21068 (N_21068,N_17930,N_17277);
nor U21069 (N_21069,N_18677,N_15663);
nor U21070 (N_21070,N_16648,N_16596);
and U21071 (N_21071,N_15945,N_17125);
and U21072 (N_21072,N_17572,N_17536);
nor U21073 (N_21073,N_16233,N_17847);
xor U21074 (N_21074,N_17765,N_16313);
or U21075 (N_21075,N_16152,N_17472);
nand U21076 (N_21076,N_17570,N_18150);
and U21077 (N_21077,N_16338,N_16713);
and U21078 (N_21078,N_16207,N_17618);
nand U21079 (N_21079,N_15827,N_16768);
or U21080 (N_21080,N_16978,N_16632);
nor U21081 (N_21081,N_16280,N_16319);
nand U21082 (N_21082,N_15973,N_16270);
nand U21083 (N_21083,N_16700,N_17004);
or U21084 (N_21084,N_16037,N_18365);
xnor U21085 (N_21085,N_15683,N_16480);
nand U21086 (N_21086,N_15628,N_17397);
xor U21087 (N_21087,N_15800,N_18126);
nor U21088 (N_21088,N_18192,N_17595);
xnor U21089 (N_21089,N_17299,N_17566);
nand U21090 (N_21090,N_16702,N_18314);
nor U21091 (N_21091,N_18246,N_18278);
xor U21092 (N_21092,N_16319,N_15985);
and U21093 (N_21093,N_16142,N_16768);
and U21094 (N_21094,N_16703,N_17768);
or U21095 (N_21095,N_18257,N_17139);
nand U21096 (N_21096,N_16970,N_17767);
and U21097 (N_21097,N_16077,N_15998);
nor U21098 (N_21098,N_18557,N_16234);
nand U21099 (N_21099,N_18076,N_18018);
or U21100 (N_21100,N_16613,N_18616);
and U21101 (N_21101,N_18311,N_17263);
nand U21102 (N_21102,N_15894,N_17555);
or U21103 (N_21103,N_17844,N_17379);
or U21104 (N_21104,N_15995,N_17183);
or U21105 (N_21105,N_17858,N_17168);
or U21106 (N_21106,N_16448,N_17549);
xor U21107 (N_21107,N_16127,N_17825);
or U21108 (N_21108,N_15829,N_18309);
or U21109 (N_21109,N_17831,N_18090);
and U21110 (N_21110,N_15979,N_18545);
nand U21111 (N_21111,N_18246,N_17181);
and U21112 (N_21112,N_16152,N_17728);
xor U21113 (N_21113,N_16595,N_16378);
and U21114 (N_21114,N_18438,N_16933);
nand U21115 (N_21115,N_18495,N_17883);
nand U21116 (N_21116,N_17894,N_15804);
xnor U21117 (N_21117,N_16159,N_17388);
nor U21118 (N_21118,N_17517,N_15766);
xor U21119 (N_21119,N_18103,N_17499);
nor U21120 (N_21120,N_15667,N_17549);
nor U21121 (N_21121,N_18505,N_17093);
or U21122 (N_21122,N_18291,N_15925);
and U21123 (N_21123,N_16833,N_16584);
and U21124 (N_21124,N_18255,N_17050);
nand U21125 (N_21125,N_17100,N_18064);
nand U21126 (N_21126,N_16548,N_16041);
and U21127 (N_21127,N_17950,N_17603);
xor U21128 (N_21128,N_17710,N_16024);
or U21129 (N_21129,N_17025,N_17608);
nor U21130 (N_21130,N_15922,N_18519);
and U21131 (N_21131,N_16044,N_17673);
and U21132 (N_21132,N_16435,N_18438);
nor U21133 (N_21133,N_16809,N_18626);
and U21134 (N_21134,N_18254,N_16863);
and U21135 (N_21135,N_17815,N_18189);
nand U21136 (N_21136,N_15626,N_16534);
and U21137 (N_21137,N_17135,N_17003);
nor U21138 (N_21138,N_16794,N_15797);
xor U21139 (N_21139,N_16073,N_16725);
or U21140 (N_21140,N_17420,N_17698);
or U21141 (N_21141,N_16715,N_16089);
nor U21142 (N_21142,N_18035,N_15814);
and U21143 (N_21143,N_18371,N_18605);
nor U21144 (N_21144,N_16995,N_18749);
or U21145 (N_21145,N_16517,N_18434);
nand U21146 (N_21146,N_18420,N_17102);
nand U21147 (N_21147,N_18283,N_16295);
and U21148 (N_21148,N_16018,N_17329);
or U21149 (N_21149,N_16346,N_17214);
nand U21150 (N_21150,N_15996,N_18443);
xor U21151 (N_21151,N_16353,N_16380);
and U21152 (N_21152,N_17166,N_16111);
nor U21153 (N_21153,N_17307,N_16147);
nand U21154 (N_21154,N_17084,N_18138);
xnor U21155 (N_21155,N_16266,N_18140);
or U21156 (N_21156,N_16725,N_16327);
xor U21157 (N_21157,N_18610,N_17100);
nor U21158 (N_21158,N_16695,N_16758);
nand U21159 (N_21159,N_16716,N_16991);
nor U21160 (N_21160,N_18673,N_18513);
and U21161 (N_21161,N_17772,N_17717);
and U21162 (N_21162,N_16513,N_15703);
or U21163 (N_21163,N_18505,N_16015);
nor U21164 (N_21164,N_16104,N_16620);
nand U21165 (N_21165,N_18270,N_16509);
nor U21166 (N_21166,N_17674,N_16536);
nor U21167 (N_21167,N_17361,N_18281);
and U21168 (N_21168,N_17962,N_16305);
and U21169 (N_21169,N_16438,N_15655);
and U21170 (N_21170,N_17441,N_17195);
nor U21171 (N_21171,N_18701,N_18477);
or U21172 (N_21172,N_18523,N_16401);
nor U21173 (N_21173,N_16887,N_17350);
or U21174 (N_21174,N_18264,N_16640);
nand U21175 (N_21175,N_16619,N_17806);
xor U21176 (N_21176,N_17135,N_17604);
and U21177 (N_21177,N_16966,N_17638);
xnor U21178 (N_21178,N_18324,N_18675);
nor U21179 (N_21179,N_16665,N_16194);
xor U21180 (N_21180,N_16465,N_16490);
or U21181 (N_21181,N_17990,N_16103);
or U21182 (N_21182,N_15888,N_16223);
nor U21183 (N_21183,N_18263,N_18383);
and U21184 (N_21184,N_18403,N_17158);
and U21185 (N_21185,N_16451,N_16671);
nor U21186 (N_21186,N_17943,N_16479);
or U21187 (N_21187,N_17013,N_18415);
and U21188 (N_21188,N_17687,N_16504);
and U21189 (N_21189,N_16954,N_17247);
xnor U21190 (N_21190,N_17601,N_17052);
and U21191 (N_21191,N_16805,N_17619);
nor U21192 (N_21192,N_17325,N_18543);
xor U21193 (N_21193,N_16924,N_15626);
and U21194 (N_21194,N_16285,N_17870);
nand U21195 (N_21195,N_16610,N_18082);
xnor U21196 (N_21196,N_15962,N_15654);
nand U21197 (N_21197,N_16796,N_18191);
xnor U21198 (N_21198,N_15745,N_16254);
or U21199 (N_21199,N_17220,N_16244);
nor U21200 (N_21200,N_15667,N_18725);
and U21201 (N_21201,N_16525,N_17366);
and U21202 (N_21202,N_18184,N_17376);
xor U21203 (N_21203,N_17833,N_17450);
and U21204 (N_21204,N_16144,N_16952);
or U21205 (N_21205,N_17175,N_17532);
and U21206 (N_21206,N_17635,N_15950);
nand U21207 (N_21207,N_16886,N_16095);
and U21208 (N_21208,N_15939,N_15742);
nand U21209 (N_21209,N_18231,N_15794);
nor U21210 (N_21210,N_17723,N_17471);
xnor U21211 (N_21211,N_17447,N_17356);
xor U21212 (N_21212,N_18067,N_18427);
nor U21213 (N_21213,N_18733,N_16903);
and U21214 (N_21214,N_16309,N_18484);
xnor U21215 (N_21215,N_16059,N_16228);
or U21216 (N_21216,N_16720,N_18403);
or U21217 (N_21217,N_16979,N_18388);
nor U21218 (N_21218,N_17504,N_17195);
and U21219 (N_21219,N_17518,N_15952);
and U21220 (N_21220,N_17967,N_17142);
and U21221 (N_21221,N_18011,N_17525);
xor U21222 (N_21222,N_17161,N_17514);
nand U21223 (N_21223,N_15704,N_16075);
xor U21224 (N_21224,N_16426,N_18689);
nor U21225 (N_21225,N_17091,N_16725);
and U21226 (N_21226,N_16107,N_16043);
and U21227 (N_21227,N_16934,N_18398);
or U21228 (N_21228,N_17328,N_16647);
xor U21229 (N_21229,N_17012,N_18209);
and U21230 (N_21230,N_17299,N_17745);
nor U21231 (N_21231,N_16833,N_18649);
or U21232 (N_21232,N_17444,N_15793);
xor U21233 (N_21233,N_18231,N_17605);
xnor U21234 (N_21234,N_16639,N_17544);
and U21235 (N_21235,N_16973,N_16537);
and U21236 (N_21236,N_18393,N_16423);
and U21237 (N_21237,N_18119,N_15710);
and U21238 (N_21238,N_15878,N_17674);
or U21239 (N_21239,N_18494,N_15717);
xnor U21240 (N_21240,N_17379,N_16775);
and U21241 (N_21241,N_17853,N_17744);
or U21242 (N_21242,N_16988,N_15688);
and U21243 (N_21243,N_16305,N_15776);
xor U21244 (N_21244,N_16834,N_16452);
or U21245 (N_21245,N_15847,N_18463);
nand U21246 (N_21246,N_18696,N_17724);
nand U21247 (N_21247,N_18509,N_15802);
and U21248 (N_21248,N_18167,N_17645);
and U21249 (N_21249,N_17827,N_16965);
nand U21250 (N_21250,N_16394,N_16800);
and U21251 (N_21251,N_17216,N_17877);
xor U21252 (N_21252,N_16053,N_16708);
xor U21253 (N_21253,N_16052,N_16577);
nand U21254 (N_21254,N_17012,N_17565);
xor U21255 (N_21255,N_17913,N_15690);
or U21256 (N_21256,N_16352,N_16128);
and U21257 (N_21257,N_18649,N_18630);
nand U21258 (N_21258,N_16162,N_18244);
nand U21259 (N_21259,N_16065,N_17639);
or U21260 (N_21260,N_18729,N_18649);
nand U21261 (N_21261,N_16336,N_17263);
xor U21262 (N_21262,N_17574,N_18635);
and U21263 (N_21263,N_16190,N_18334);
and U21264 (N_21264,N_15992,N_16997);
nand U21265 (N_21265,N_18562,N_17381);
and U21266 (N_21266,N_17689,N_15881);
or U21267 (N_21267,N_18635,N_17434);
nand U21268 (N_21268,N_17165,N_16669);
nand U21269 (N_21269,N_18439,N_17421);
nand U21270 (N_21270,N_16123,N_18224);
nand U21271 (N_21271,N_18182,N_18543);
nor U21272 (N_21272,N_17851,N_18269);
xnor U21273 (N_21273,N_18150,N_16697);
nand U21274 (N_21274,N_15793,N_17117);
or U21275 (N_21275,N_16671,N_16690);
and U21276 (N_21276,N_18721,N_17377);
and U21277 (N_21277,N_17552,N_17382);
nor U21278 (N_21278,N_17130,N_16007);
or U21279 (N_21279,N_16917,N_16372);
and U21280 (N_21280,N_17644,N_18094);
or U21281 (N_21281,N_17683,N_17052);
xnor U21282 (N_21282,N_18149,N_18403);
xnor U21283 (N_21283,N_18161,N_15887);
nor U21284 (N_21284,N_16059,N_17930);
xor U21285 (N_21285,N_16459,N_16382);
nand U21286 (N_21286,N_17058,N_17551);
nor U21287 (N_21287,N_18184,N_16007);
or U21288 (N_21288,N_17926,N_17101);
xnor U21289 (N_21289,N_16065,N_18256);
or U21290 (N_21290,N_16146,N_16515);
and U21291 (N_21291,N_18047,N_17288);
xor U21292 (N_21292,N_16482,N_18510);
xor U21293 (N_21293,N_17492,N_16768);
nor U21294 (N_21294,N_17884,N_17975);
nor U21295 (N_21295,N_16779,N_18748);
xor U21296 (N_21296,N_16322,N_18597);
and U21297 (N_21297,N_18503,N_16784);
or U21298 (N_21298,N_18104,N_16043);
or U21299 (N_21299,N_17209,N_16344);
or U21300 (N_21300,N_17923,N_18089);
nand U21301 (N_21301,N_15940,N_18526);
or U21302 (N_21302,N_15677,N_16465);
nor U21303 (N_21303,N_17176,N_18136);
nand U21304 (N_21304,N_17571,N_17010);
and U21305 (N_21305,N_17997,N_18367);
xor U21306 (N_21306,N_16180,N_16792);
xnor U21307 (N_21307,N_17768,N_18719);
xnor U21308 (N_21308,N_17313,N_16241);
nor U21309 (N_21309,N_16909,N_18518);
nand U21310 (N_21310,N_17676,N_18054);
xor U21311 (N_21311,N_18130,N_15804);
and U21312 (N_21312,N_17959,N_17124);
or U21313 (N_21313,N_16791,N_16488);
nor U21314 (N_21314,N_17920,N_15955);
xor U21315 (N_21315,N_15689,N_17587);
and U21316 (N_21316,N_16887,N_16969);
or U21317 (N_21317,N_18661,N_18734);
nand U21318 (N_21318,N_17404,N_17250);
or U21319 (N_21319,N_17149,N_17135);
or U21320 (N_21320,N_16601,N_18103);
or U21321 (N_21321,N_17539,N_17815);
xnor U21322 (N_21322,N_17788,N_16008);
xnor U21323 (N_21323,N_17932,N_16871);
xor U21324 (N_21324,N_18358,N_18640);
nor U21325 (N_21325,N_16083,N_17507);
nand U21326 (N_21326,N_15635,N_15939);
or U21327 (N_21327,N_16126,N_18160);
xor U21328 (N_21328,N_18264,N_17355);
nand U21329 (N_21329,N_16900,N_16909);
xor U21330 (N_21330,N_16025,N_17706);
nand U21331 (N_21331,N_16969,N_17097);
and U21332 (N_21332,N_17800,N_18298);
nand U21333 (N_21333,N_18123,N_17626);
nand U21334 (N_21334,N_16501,N_18511);
nand U21335 (N_21335,N_18613,N_16842);
nand U21336 (N_21336,N_16572,N_18252);
or U21337 (N_21337,N_17990,N_17884);
and U21338 (N_21338,N_17562,N_16515);
and U21339 (N_21339,N_18141,N_16356);
and U21340 (N_21340,N_17797,N_17223);
or U21341 (N_21341,N_16571,N_18271);
nor U21342 (N_21342,N_16272,N_16066);
nor U21343 (N_21343,N_16219,N_16598);
or U21344 (N_21344,N_16327,N_18141);
nand U21345 (N_21345,N_16769,N_18195);
or U21346 (N_21346,N_17359,N_16580);
and U21347 (N_21347,N_18599,N_17770);
nand U21348 (N_21348,N_17731,N_17558);
or U21349 (N_21349,N_17535,N_16792);
nor U21350 (N_21350,N_17545,N_17554);
nor U21351 (N_21351,N_17040,N_18013);
nand U21352 (N_21352,N_16060,N_15831);
or U21353 (N_21353,N_15731,N_17577);
xor U21354 (N_21354,N_17403,N_16356);
nor U21355 (N_21355,N_18718,N_17828);
xor U21356 (N_21356,N_15932,N_15916);
nand U21357 (N_21357,N_16824,N_18236);
and U21358 (N_21358,N_18676,N_16268);
or U21359 (N_21359,N_17917,N_16240);
nor U21360 (N_21360,N_18258,N_17547);
nor U21361 (N_21361,N_15777,N_17353);
nand U21362 (N_21362,N_17266,N_16039);
nor U21363 (N_21363,N_17983,N_16658);
nor U21364 (N_21364,N_16819,N_16569);
xnor U21365 (N_21365,N_18618,N_17508);
nor U21366 (N_21366,N_18125,N_15779);
xnor U21367 (N_21367,N_18447,N_15726);
or U21368 (N_21368,N_16466,N_15822);
nor U21369 (N_21369,N_16746,N_18198);
and U21370 (N_21370,N_16895,N_16512);
and U21371 (N_21371,N_17399,N_18367);
nand U21372 (N_21372,N_17438,N_16109);
xnor U21373 (N_21373,N_16110,N_17578);
nand U21374 (N_21374,N_17090,N_16199);
nand U21375 (N_21375,N_17295,N_16715);
xnor U21376 (N_21376,N_17390,N_17483);
xnor U21377 (N_21377,N_18276,N_17841);
and U21378 (N_21378,N_16563,N_16498);
nor U21379 (N_21379,N_16355,N_17837);
and U21380 (N_21380,N_17333,N_16012);
or U21381 (N_21381,N_17125,N_17292);
or U21382 (N_21382,N_15717,N_16601);
nor U21383 (N_21383,N_16997,N_16612);
nand U21384 (N_21384,N_16120,N_16984);
or U21385 (N_21385,N_16035,N_18351);
xnor U21386 (N_21386,N_18347,N_16305);
nor U21387 (N_21387,N_17953,N_18384);
nor U21388 (N_21388,N_17560,N_16956);
xor U21389 (N_21389,N_16919,N_15703);
or U21390 (N_21390,N_16850,N_16990);
nand U21391 (N_21391,N_17527,N_18046);
nand U21392 (N_21392,N_18031,N_18224);
or U21393 (N_21393,N_17357,N_16699);
xnor U21394 (N_21394,N_17278,N_18177);
nand U21395 (N_21395,N_16807,N_18482);
xnor U21396 (N_21396,N_16707,N_15808);
and U21397 (N_21397,N_17326,N_17764);
and U21398 (N_21398,N_17585,N_17364);
or U21399 (N_21399,N_17796,N_16725);
and U21400 (N_21400,N_18169,N_16893);
and U21401 (N_21401,N_18130,N_15667);
xor U21402 (N_21402,N_18737,N_17980);
nand U21403 (N_21403,N_17419,N_16089);
or U21404 (N_21404,N_18477,N_16362);
xnor U21405 (N_21405,N_18481,N_16829);
or U21406 (N_21406,N_18109,N_16606);
xnor U21407 (N_21407,N_16740,N_15937);
or U21408 (N_21408,N_16998,N_16541);
nor U21409 (N_21409,N_16459,N_16168);
or U21410 (N_21410,N_15717,N_17918);
or U21411 (N_21411,N_15756,N_17720);
xnor U21412 (N_21412,N_16671,N_18546);
and U21413 (N_21413,N_16862,N_18325);
nor U21414 (N_21414,N_16345,N_16425);
or U21415 (N_21415,N_18489,N_16030);
and U21416 (N_21416,N_17448,N_16510);
xnor U21417 (N_21417,N_16367,N_16926);
nand U21418 (N_21418,N_18025,N_15777);
xor U21419 (N_21419,N_16859,N_16744);
nand U21420 (N_21420,N_18510,N_17854);
or U21421 (N_21421,N_15806,N_18545);
nand U21422 (N_21422,N_16128,N_15669);
nor U21423 (N_21423,N_16399,N_18578);
and U21424 (N_21424,N_16331,N_15795);
and U21425 (N_21425,N_17364,N_17715);
nand U21426 (N_21426,N_17534,N_17809);
xnor U21427 (N_21427,N_18715,N_16835);
nand U21428 (N_21428,N_16783,N_17680);
nor U21429 (N_21429,N_16301,N_18404);
nor U21430 (N_21430,N_15837,N_16869);
nand U21431 (N_21431,N_16490,N_15757);
xor U21432 (N_21432,N_16824,N_16810);
xnor U21433 (N_21433,N_16769,N_18412);
xor U21434 (N_21434,N_17302,N_16829);
xor U21435 (N_21435,N_16284,N_16129);
nor U21436 (N_21436,N_15626,N_16666);
or U21437 (N_21437,N_17635,N_18734);
and U21438 (N_21438,N_16862,N_18338);
or U21439 (N_21439,N_18689,N_18620);
and U21440 (N_21440,N_17415,N_16277);
or U21441 (N_21441,N_18047,N_15722);
and U21442 (N_21442,N_18685,N_18587);
and U21443 (N_21443,N_17066,N_17604);
or U21444 (N_21444,N_17981,N_15961);
nand U21445 (N_21445,N_16293,N_17169);
nor U21446 (N_21446,N_18267,N_18357);
and U21447 (N_21447,N_16742,N_15779);
and U21448 (N_21448,N_16857,N_16802);
or U21449 (N_21449,N_15883,N_17408);
nand U21450 (N_21450,N_17586,N_16743);
or U21451 (N_21451,N_18342,N_16039);
xnor U21452 (N_21452,N_16491,N_16268);
nor U21453 (N_21453,N_17819,N_17990);
and U21454 (N_21454,N_17880,N_18538);
nor U21455 (N_21455,N_16736,N_16767);
or U21456 (N_21456,N_17760,N_16404);
nand U21457 (N_21457,N_16410,N_17650);
nand U21458 (N_21458,N_17530,N_17575);
xnor U21459 (N_21459,N_16163,N_16268);
and U21460 (N_21460,N_17879,N_16991);
nand U21461 (N_21461,N_17735,N_17697);
nor U21462 (N_21462,N_17598,N_17654);
or U21463 (N_21463,N_16123,N_18545);
or U21464 (N_21464,N_15723,N_17043);
and U21465 (N_21465,N_15755,N_18518);
nor U21466 (N_21466,N_16584,N_18022);
and U21467 (N_21467,N_16046,N_16594);
and U21468 (N_21468,N_16617,N_18638);
and U21469 (N_21469,N_16421,N_18116);
nand U21470 (N_21470,N_18470,N_15711);
nand U21471 (N_21471,N_17677,N_17800);
nand U21472 (N_21472,N_16952,N_18011);
or U21473 (N_21473,N_17329,N_17469);
nor U21474 (N_21474,N_18718,N_16725);
nor U21475 (N_21475,N_18547,N_18599);
and U21476 (N_21476,N_16504,N_16851);
nand U21477 (N_21477,N_17962,N_15630);
xor U21478 (N_21478,N_16159,N_18114);
nor U21479 (N_21479,N_18422,N_18262);
xnor U21480 (N_21480,N_16620,N_17320);
nand U21481 (N_21481,N_18403,N_15881);
and U21482 (N_21482,N_17350,N_15856);
nor U21483 (N_21483,N_15713,N_17188);
nor U21484 (N_21484,N_17083,N_17978);
and U21485 (N_21485,N_16328,N_16034);
xnor U21486 (N_21486,N_15907,N_16973);
or U21487 (N_21487,N_16137,N_16560);
nand U21488 (N_21488,N_16407,N_16854);
and U21489 (N_21489,N_16387,N_17673);
and U21490 (N_21490,N_18402,N_18363);
nand U21491 (N_21491,N_17849,N_18237);
and U21492 (N_21492,N_16432,N_15638);
and U21493 (N_21493,N_16031,N_17633);
xor U21494 (N_21494,N_16164,N_18566);
nor U21495 (N_21495,N_17389,N_18194);
xnor U21496 (N_21496,N_17842,N_15987);
or U21497 (N_21497,N_15741,N_17978);
nor U21498 (N_21498,N_18283,N_17627);
nand U21499 (N_21499,N_17157,N_18327);
or U21500 (N_21500,N_18477,N_15857);
nor U21501 (N_21501,N_15990,N_17181);
and U21502 (N_21502,N_16234,N_17682);
or U21503 (N_21503,N_16957,N_18279);
and U21504 (N_21504,N_16226,N_17852);
xor U21505 (N_21505,N_15950,N_15778);
nand U21506 (N_21506,N_18690,N_17745);
xor U21507 (N_21507,N_17938,N_18633);
xnor U21508 (N_21508,N_18458,N_18069);
or U21509 (N_21509,N_17691,N_15994);
or U21510 (N_21510,N_16652,N_18537);
xnor U21511 (N_21511,N_18499,N_16986);
xnor U21512 (N_21512,N_17906,N_18419);
nand U21513 (N_21513,N_16489,N_16592);
or U21514 (N_21514,N_16566,N_17981);
or U21515 (N_21515,N_15972,N_17783);
nand U21516 (N_21516,N_18616,N_17067);
nor U21517 (N_21517,N_17355,N_17120);
or U21518 (N_21518,N_16219,N_18457);
and U21519 (N_21519,N_18192,N_16313);
and U21520 (N_21520,N_17714,N_17940);
or U21521 (N_21521,N_17108,N_16985);
xor U21522 (N_21522,N_16639,N_15845);
nor U21523 (N_21523,N_17566,N_16631);
nand U21524 (N_21524,N_18670,N_18004);
xnor U21525 (N_21525,N_15852,N_16807);
or U21526 (N_21526,N_16250,N_15731);
xor U21527 (N_21527,N_18660,N_18200);
nor U21528 (N_21528,N_16415,N_16536);
nand U21529 (N_21529,N_17382,N_15737);
xnor U21530 (N_21530,N_16212,N_17769);
or U21531 (N_21531,N_18045,N_16424);
and U21532 (N_21532,N_16075,N_17508);
and U21533 (N_21533,N_16522,N_17196);
and U21534 (N_21534,N_15628,N_16973);
and U21535 (N_21535,N_17179,N_17382);
xor U21536 (N_21536,N_18475,N_15781);
xor U21537 (N_21537,N_18448,N_15763);
or U21538 (N_21538,N_18357,N_16270);
xor U21539 (N_21539,N_16699,N_18060);
nand U21540 (N_21540,N_16495,N_16779);
or U21541 (N_21541,N_16851,N_18107);
and U21542 (N_21542,N_16685,N_16737);
xor U21543 (N_21543,N_18297,N_15896);
nand U21544 (N_21544,N_15854,N_17448);
xor U21545 (N_21545,N_17594,N_17906);
nand U21546 (N_21546,N_17502,N_16484);
nor U21547 (N_21547,N_16274,N_17593);
xnor U21548 (N_21548,N_18591,N_17660);
and U21549 (N_21549,N_17806,N_16735);
nand U21550 (N_21550,N_16763,N_17532);
or U21551 (N_21551,N_18656,N_18675);
and U21552 (N_21552,N_16996,N_15996);
xnor U21553 (N_21553,N_17354,N_17120);
nor U21554 (N_21554,N_16228,N_16249);
nand U21555 (N_21555,N_18486,N_16205);
nand U21556 (N_21556,N_18118,N_15990);
and U21557 (N_21557,N_16032,N_18647);
or U21558 (N_21558,N_18402,N_17165);
nand U21559 (N_21559,N_17457,N_16903);
xnor U21560 (N_21560,N_18114,N_18508);
xor U21561 (N_21561,N_16687,N_17797);
xnor U21562 (N_21562,N_16971,N_16355);
nand U21563 (N_21563,N_17763,N_17152);
or U21564 (N_21564,N_17964,N_18067);
nand U21565 (N_21565,N_16775,N_16381);
and U21566 (N_21566,N_15998,N_15829);
or U21567 (N_21567,N_16435,N_15908);
xor U21568 (N_21568,N_15894,N_16633);
xor U21569 (N_21569,N_16036,N_17344);
and U21570 (N_21570,N_16445,N_16761);
and U21571 (N_21571,N_18230,N_16602);
and U21572 (N_21572,N_15833,N_18304);
nand U21573 (N_21573,N_16233,N_17512);
nand U21574 (N_21574,N_18268,N_18050);
and U21575 (N_21575,N_15981,N_16203);
nand U21576 (N_21576,N_18201,N_17172);
nor U21577 (N_21577,N_16740,N_17257);
nand U21578 (N_21578,N_16256,N_16607);
or U21579 (N_21579,N_17866,N_18413);
nand U21580 (N_21580,N_16898,N_15713);
xnor U21581 (N_21581,N_16164,N_17532);
nor U21582 (N_21582,N_15907,N_17846);
or U21583 (N_21583,N_17659,N_18232);
nand U21584 (N_21584,N_15836,N_18024);
xor U21585 (N_21585,N_16258,N_16526);
nor U21586 (N_21586,N_17556,N_17202);
nor U21587 (N_21587,N_16150,N_16581);
nand U21588 (N_21588,N_17488,N_18540);
xnor U21589 (N_21589,N_17477,N_18011);
and U21590 (N_21590,N_16232,N_17485);
nand U21591 (N_21591,N_17448,N_16791);
or U21592 (N_21592,N_17669,N_18270);
nor U21593 (N_21593,N_15822,N_16701);
xnor U21594 (N_21594,N_18316,N_18321);
xnor U21595 (N_21595,N_16170,N_18159);
and U21596 (N_21596,N_17774,N_17486);
and U21597 (N_21597,N_16173,N_17933);
or U21598 (N_21598,N_17619,N_18508);
and U21599 (N_21599,N_18528,N_16535);
xnor U21600 (N_21600,N_16268,N_17589);
nor U21601 (N_21601,N_18713,N_16868);
xor U21602 (N_21602,N_16813,N_15831);
or U21603 (N_21603,N_17100,N_16235);
nand U21604 (N_21604,N_18196,N_17475);
or U21605 (N_21605,N_16082,N_16419);
nor U21606 (N_21606,N_18051,N_17689);
xnor U21607 (N_21607,N_16350,N_16400);
and U21608 (N_21608,N_16701,N_16503);
or U21609 (N_21609,N_16661,N_17890);
nand U21610 (N_21610,N_18539,N_16719);
xnor U21611 (N_21611,N_16693,N_16593);
xor U21612 (N_21612,N_18361,N_18006);
nand U21613 (N_21613,N_18427,N_18062);
and U21614 (N_21614,N_17282,N_18235);
nor U21615 (N_21615,N_16242,N_17689);
or U21616 (N_21616,N_16345,N_17837);
nand U21617 (N_21617,N_15859,N_18207);
and U21618 (N_21618,N_17914,N_16481);
or U21619 (N_21619,N_17729,N_17411);
nand U21620 (N_21620,N_16271,N_18390);
nor U21621 (N_21621,N_17559,N_16405);
nor U21622 (N_21622,N_18567,N_17270);
xor U21623 (N_21623,N_18374,N_18040);
nor U21624 (N_21624,N_16287,N_18320);
or U21625 (N_21625,N_15917,N_18527);
nand U21626 (N_21626,N_16379,N_17707);
or U21627 (N_21627,N_18416,N_16008);
nand U21628 (N_21628,N_16590,N_17107);
nand U21629 (N_21629,N_18187,N_15910);
xor U21630 (N_21630,N_17994,N_16938);
nor U21631 (N_21631,N_17406,N_18407);
and U21632 (N_21632,N_16785,N_17634);
and U21633 (N_21633,N_18500,N_17444);
nor U21634 (N_21634,N_17043,N_16114);
and U21635 (N_21635,N_17152,N_18102);
nor U21636 (N_21636,N_17608,N_17524);
xor U21637 (N_21637,N_18065,N_16808);
nand U21638 (N_21638,N_16650,N_17450);
and U21639 (N_21639,N_17464,N_16674);
nand U21640 (N_21640,N_15886,N_16441);
nor U21641 (N_21641,N_17098,N_16485);
or U21642 (N_21642,N_17214,N_17837);
xor U21643 (N_21643,N_16239,N_15777);
and U21644 (N_21644,N_15962,N_16688);
and U21645 (N_21645,N_17900,N_17283);
xnor U21646 (N_21646,N_15744,N_15884);
xnor U21647 (N_21647,N_17259,N_16996);
and U21648 (N_21648,N_18745,N_17403);
or U21649 (N_21649,N_18676,N_17303);
nor U21650 (N_21650,N_17613,N_18202);
nand U21651 (N_21651,N_15777,N_17330);
nand U21652 (N_21652,N_16506,N_16144);
and U21653 (N_21653,N_16037,N_16141);
xnor U21654 (N_21654,N_15715,N_16250);
xor U21655 (N_21655,N_18020,N_15968);
xor U21656 (N_21656,N_16395,N_18136);
nand U21657 (N_21657,N_15904,N_18353);
or U21658 (N_21658,N_16088,N_16246);
and U21659 (N_21659,N_17830,N_16324);
or U21660 (N_21660,N_18545,N_18390);
and U21661 (N_21661,N_16807,N_17168);
nand U21662 (N_21662,N_15658,N_17973);
xnor U21663 (N_21663,N_16349,N_18666);
xor U21664 (N_21664,N_17083,N_16888);
xor U21665 (N_21665,N_15725,N_16495);
nor U21666 (N_21666,N_17249,N_17115);
xnor U21667 (N_21667,N_18330,N_15955);
or U21668 (N_21668,N_18015,N_18378);
nand U21669 (N_21669,N_17096,N_18452);
nor U21670 (N_21670,N_15774,N_15807);
or U21671 (N_21671,N_17422,N_16167);
xor U21672 (N_21672,N_17245,N_17181);
and U21673 (N_21673,N_16908,N_16937);
and U21674 (N_21674,N_16582,N_15715);
or U21675 (N_21675,N_18682,N_15980);
xor U21676 (N_21676,N_17250,N_17554);
nor U21677 (N_21677,N_16924,N_16522);
or U21678 (N_21678,N_17081,N_16117);
and U21679 (N_21679,N_17392,N_16989);
nor U21680 (N_21680,N_16340,N_16701);
and U21681 (N_21681,N_17975,N_17499);
xor U21682 (N_21682,N_18666,N_18239);
xnor U21683 (N_21683,N_17350,N_17889);
or U21684 (N_21684,N_17531,N_16621);
or U21685 (N_21685,N_17808,N_15752);
nor U21686 (N_21686,N_18600,N_16389);
or U21687 (N_21687,N_16732,N_16557);
and U21688 (N_21688,N_17698,N_16359);
xor U21689 (N_21689,N_16185,N_18695);
and U21690 (N_21690,N_16627,N_18084);
nor U21691 (N_21691,N_17557,N_16490);
nand U21692 (N_21692,N_16803,N_16577);
xnor U21693 (N_21693,N_17617,N_16892);
nor U21694 (N_21694,N_15714,N_18004);
or U21695 (N_21695,N_16230,N_17890);
and U21696 (N_21696,N_16072,N_17071);
xnor U21697 (N_21697,N_16959,N_17887);
nor U21698 (N_21698,N_16579,N_16848);
nand U21699 (N_21699,N_16587,N_15635);
nor U21700 (N_21700,N_18239,N_17104);
or U21701 (N_21701,N_16433,N_18422);
nand U21702 (N_21702,N_18221,N_18402);
nand U21703 (N_21703,N_18650,N_16641);
or U21704 (N_21704,N_17120,N_16128);
xor U21705 (N_21705,N_18380,N_18492);
nand U21706 (N_21706,N_15747,N_17472);
nor U21707 (N_21707,N_16484,N_17599);
or U21708 (N_21708,N_15784,N_17379);
xnor U21709 (N_21709,N_17158,N_16176);
nor U21710 (N_21710,N_17247,N_15793);
xnor U21711 (N_21711,N_17229,N_18429);
nand U21712 (N_21712,N_16286,N_17112);
nand U21713 (N_21713,N_15861,N_16126);
nand U21714 (N_21714,N_18391,N_17047);
nor U21715 (N_21715,N_18264,N_18243);
nor U21716 (N_21716,N_16907,N_18103);
xnor U21717 (N_21717,N_17629,N_16483);
xor U21718 (N_21718,N_15981,N_18714);
nand U21719 (N_21719,N_16946,N_17562);
and U21720 (N_21720,N_17307,N_18721);
and U21721 (N_21721,N_18159,N_15848);
nor U21722 (N_21722,N_18696,N_15681);
xor U21723 (N_21723,N_16425,N_17610);
nand U21724 (N_21724,N_16596,N_17020);
and U21725 (N_21725,N_15780,N_18453);
xor U21726 (N_21726,N_18308,N_17613);
nor U21727 (N_21727,N_16355,N_17797);
nor U21728 (N_21728,N_18393,N_17565);
xnor U21729 (N_21729,N_16593,N_16874);
or U21730 (N_21730,N_18518,N_16493);
nor U21731 (N_21731,N_15894,N_16814);
or U21732 (N_21732,N_17275,N_17173);
or U21733 (N_21733,N_18596,N_16102);
nor U21734 (N_21734,N_15972,N_18666);
nor U21735 (N_21735,N_18156,N_16405);
xor U21736 (N_21736,N_16081,N_16656);
xnor U21737 (N_21737,N_15860,N_16398);
or U21738 (N_21738,N_16559,N_15764);
xor U21739 (N_21739,N_15809,N_16610);
or U21740 (N_21740,N_17661,N_17576);
and U21741 (N_21741,N_17306,N_17630);
and U21742 (N_21742,N_17225,N_16895);
nand U21743 (N_21743,N_16879,N_15776);
nand U21744 (N_21744,N_18371,N_16459);
or U21745 (N_21745,N_16395,N_17908);
xnor U21746 (N_21746,N_17890,N_16968);
or U21747 (N_21747,N_16066,N_17302);
nand U21748 (N_21748,N_16647,N_17578);
and U21749 (N_21749,N_17146,N_16212);
xor U21750 (N_21750,N_15963,N_15719);
nor U21751 (N_21751,N_17935,N_17888);
or U21752 (N_21752,N_17574,N_16129);
and U21753 (N_21753,N_16523,N_16559);
xnor U21754 (N_21754,N_18645,N_18519);
xor U21755 (N_21755,N_17192,N_18598);
or U21756 (N_21756,N_18626,N_18050);
nor U21757 (N_21757,N_16907,N_18402);
nor U21758 (N_21758,N_17180,N_18573);
xnor U21759 (N_21759,N_17409,N_15971);
nor U21760 (N_21760,N_16158,N_18483);
and U21761 (N_21761,N_17966,N_16444);
xnor U21762 (N_21762,N_16590,N_17647);
and U21763 (N_21763,N_15955,N_16990);
nor U21764 (N_21764,N_17166,N_17155);
nor U21765 (N_21765,N_18462,N_18674);
nor U21766 (N_21766,N_16630,N_18731);
xor U21767 (N_21767,N_15768,N_18081);
and U21768 (N_21768,N_16787,N_16519);
or U21769 (N_21769,N_18334,N_17343);
nor U21770 (N_21770,N_17272,N_18718);
nand U21771 (N_21771,N_16224,N_16837);
nor U21772 (N_21772,N_16748,N_16148);
or U21773 (N_21773,N_17347,N_16487);
and U21774 (N_21774,N_18419,N_16544);
or U21775 (N_21775,N_17760,N_18008);
or U21776 (N_21776,N_16122,N_16570);
or U21777 (N_21777,N_16303,N_18726);
nor U21778 (N_21778,N_15671,N_17983);
nor U21779 (N_21779,N_16568,N_17652);
nor U21780 (N_21780,N_17643,N_15699);
nor U21781 (N_21781,N_16849,N_15975);
nor U21782 (N_21782,N_16956,N_18381);
nand U21783 (N_21783,N_17120,N_17895);
xor U21784 (N_21784,N_18065,N_18602);
or U21785 (N_21785,N_18497,N_18265);
or U21786 (N_21786,N_16983,N_17594);
nor U21787 (N_21787,N_18708,N_17708);
nand U21788 (N_21788,N_16772,N_16133);
nor U21789 (N_21789,N_16109,N_16619);
or U21790 (N_21790,N_15927,N_16129);
nor U21791 (N_21791,N_16558,N_18109);
and U21792 (N_21792,N_18620,N_16972);
and U21793 (N_21793,N_18621,N_15800);
or U21794 (N_21794,N_16017,N_17531);
nand U21795 (N_21795,N_17368,N_16010);
xnor U21796 (N_21796,N_16629,N_15867);
xor U21797 (N_21797,N_15723,N_17205);
and U21798 (N_21798,N_16956,N_18689);
or U21799 (N_21799,N_16627,N_18194);
nand U21800 (N_21800,N_17922,N_16021);
and U21801 (N_21801,N_18390,N_16203);
or U21802 (N_21802,N_16217,N_18314);
or U21803 (N_21803,N_18744,N_17999);
nand U21804 (N_21804,N_18374,N_17474);
nor U21805 (N_21805,N_16358,N_17591);
nor U21806 (N_21806,N_16547,N_17791);
or U21807 (N_21807,N_17128,N_18428);
nand U21808 (N_21808,N_17523,N_16575);
and U21809 (N_21809,N_15868,N_17474);
nand U21810 (N_21810,N_15910,N_18155);
or U21811 (N_21811,N_18560,N_15714);
and U21812 (N_21812,N_17839,N_17019);
and U21813 (N_21813,N_15729,N_18637);
xnor U21814 (N_21814,N_17593,N_15682);
xnor U21815 (N_21815,N_17669,N_15660);
and U21816 (N_21816,N_16247,N_16500);
or U21817 (N_21817,N_16740,N_17542);
or U21818 (N_21818,N_18604,N_17920);
or U21819 (N_21819,N_17549,N_16280);
and U21820 (N_21820,N_16028,N_16525);
xor U21821 (N_21821,N_15631,N_18056);
nand U21822 (N_21822,N_17079,N_18001);
or U21823 (N_21823,N_16983,N_18527);
nor U21824 (N_21824,N_16821,N_15648);
or U21825 (N_21825,N_18686,N_18009);
or U21826 (N_21826,N_17888,N_17450);
xor U21827 (N_21827,N_17686,N_17886);
nor U21828 (N_21828,N_18465,N_16633);
xor U21829 (N_21829,N_17683,N_17429);
xor U21830 (N_21830,N_17509,N_18749);
xor U21831 (N_21831,N_17719,N_17315);
nor U21832 (N_21832,N_17355,N_17282);
xor U21833 (N_21833,N_16413,N_15816);
and U21834 (N_21834,N_16688,N_16584);
and U21835 (N_21835,N_16158,N_17010);
xor U21836 (N_21836,N_16564,N_16493);
and U21837 (N_21837,N_16015,N_16371);
and U21838 (N_21838,N_15659,N_16468);
or U21839 (N_21839,N_17127,N_17387);
nand U21840 (N_21840,N_18402,N_16007);
nor U21841 (N_21841,N_16697,N_17910);
xnor U21842 (N_21842,N_17763,N_16092);
nand U21843 (N_21843,N_17611,N_15843);
or U21844 (N_21844,N_18509,N_18069);
nor U21845 (N_21845,N_17321,N_16778);
xnor U21846 (N_21846,N_16522,N_18527);
nand U21847 (N_21847,N_15791,N_17767);
nand U21848 (N_21848,N_16970,N_18602);
and U21849 (N_21849,N_15648,N_16744);
xnor U21850 (N_21850,N_18624,N_18625);
or U21851 (N_21851,N_17383,N_17475);
nand U21852 (N_21852,N_16426,N_17766);
xnor U21853 (N_21853,N_18747,N_16808);
nand U21854 (N_21854,N_18426,N_18668);
and U21855 (N_21855,N_18725,N_16095);
nand U21856 (N_21856,N_18729,N_16113);
nor U21857 (N_21857,N_16664,N_15772);
nor U21858 (N_21858,N_17634,N_16397);
nor U21859 (N_21859,N_16656,N_17315);
nand U21860 (N_21860,N_17876,N_16464);
nand U21861 (N_21861,N_16611,N_16930);
xor U21862 (N_21862,N_18399,N_17494);
nand U21863 (N_21863,N_17353,N_15784);
and U21864 (N_21864,N_15697,N_17588);
and U21865 (N_21865,N_16075,N_16518);
xnor U21866 (N_21866,N_17693,N_17025);
xnor U21867 (N_21867,N_16229,N_16247);
nor U21868 (N_21868,N_15793,N_16791);
and U21869 (N_21869,N_16740,N_18069);
nor U21870 (N_21870,N_18710,N_17644);
and U21871 (N_21871,N_16028,N_17590);
xnor U21872 (N_21872,N_16928,N_18098);
xnor U21873 (N_21873,N_15666,N_17526);
xor U21874 (N_21874,N_16509,N_18340);
or U21875 (N_21875,N_20482,N_21273);
and U21876 (N_21876,N_20463,N_21113);
or U21877 (N_21877,N_21539,N_18750);
and U21878 (N_21878,N_19655,N_20992);
nand U21879 (N_21879,N_19098,N_19295);
nand U21880 (N_21880,N_18911,N_21257);
or U21881 (N_21881,N_20946,N_20336);
or U21882 (N_21882,N_19035,N_18813);
xnor U21883 (N_21883,N_19065,N_20771);
xor U21884 (N_21884,N_20685,N_20471);
and U21885 (N_21885,N_21362,N_18940);
or U21886 (N_21886,N_21741,N_20561);
xnor U21887 (N_21887,N_20476,N_20157);
and U21888 (N_21888,N_20397,N_18949);
xnor U21889 (N_21889,N_18818,N_20410);
or U21890 (N_21890,N_19427,N_21602);
nand U21891 (N_21891,N_19162,N_19117);
and U21892 (N_21892,N_20262,N_19536);
or U21893 (N_21893,N_20525,N_19992);
xnor U21894 (N_21894,N_18910,N_20260);
xnor U21895 (N_21895,N_20299,N_21137);
xnor U21896 (N_21896,N_20900,N_20926);
xnor U21897 (N_21897,N_21620,N_19168);
and U21898 (N_21898,N_20308,N_19000);
and U21899 (N_21899,N_20536,N_21718);
xnor U21900 (N_21900,N_19635,N_18792);
or U21901 (N_21901,N_20354,N_20684);
nand U21902 (N_21902,N_18912,N_20892);
nand U21903 (N_21903,N_20226,N_21466);
nor U21904 (N_21904,N_21021,N_20401);
or U21905 (N_21905,N_19504,N_21592);
or U21906 (N_21906,N_21552,N_19442);
xnor U21907 (N_21907,N_19336,N_20676);
xnor U21908 (N_21908,N_21596,N_21018);
nor U21909 (N_21909,N_20021,N_19493);
xor U21910 (N_21910,N_20159,N_21452);
nor U21911 (N_21911,N_19114,N_18921);
xnor U21912 (N_21912,N_21337,N_19701);
nand U21913 (N_21913,N_20769,N_19855);
nor U21914 (N_21914,N_19273,N_19437);
and U21915 (N_21915,N_18849,N_19195);
xnor U21916 (N_21916,N_21326,N_21401);
nand U21917 (N_21917,N_21861,N_21251);
nor U21918 (N_21918,N_21109,N_21493);
and U21919 (N_21919,N_20793,N_21810);
and U21920 (N_21920,N_18850,N_18996);
nor U21921 (N_21921,N_20394,N_20852);
nor U21922 (N_21922,N_18934,N_18972);
nand U21923 (N_21923,N_19345,N_21433);
nand U21924 (N_21924,N_21733,N_19112);
nor U21925 (N_21925,N_21579,N_21361);
nor U21926 (N_21926,N_19177,N_19330);
and U21927 (N_21927,N_19349,N_18832);
or U21928 (N_21928,N_19562,N_21843);
or U21929 (N_21929,N_19485,N_20837);
xnor U21930 (N_21930,N_20342,N_19833);
nor U21931 (N_21931,N_18798,N_20529);
or U21932 (N_21932,N_20286,N_20072);
nor U21933 (N_21933,N_20388,N_19964);
or U21934 (N_21934,N_19201,N_19728);
xnor U21935 (N_21935,N_19724,N_19282);
nor U21936 (N_21936,N_19256,N_19189);
xnor U21937 (N_21937,N_21315,N_20524);
or U21938 (N_21938,N_19199,N_21406);
nor U21939 (N_21939,N_21425,N_19307);
or U21940 (N_21940,N_19694,N_21051);
xnor U21941 (N_21941,N_19816,N_20168);
nand U21942 (N_21942,N_18859,N_20123);
nand U21943 (N_21943,N_21492,N_19634);
and U21944 (N_21944,N_20484,N_18869);
or U21945 (N_21945,N_19893,N_21661);
and U21946 (N_21946,N_21694,N_20126);
or U21947 (N_21947,N_19104,N_20150);
and U21948 (N_21948,N_19933,N_20681);
or U21949 (N_21949,N_21849,N_19431);
or U21950 (N_21950,N_20688,N_19678);
or U21951 (N_21951,N_20236,N_20591);
and U21952 (N_21952,N_21490,N_19159);
nor U21953 (N_21953,N_21464,N_21865);
xor U21954 (N_21954,N_21504,N_18933);
nand U21955 (N_21955,N_18992,N_19280);
nand U21956 (N_21956,N_21177,N_18848);
xor U21957 (N_21957,N_19609,N_18865);
nand U21958 (N_21958,N_21581,N_20683);
or U21959 (N_21959,N_19697,N_20078);
or U21960 (N_21960,N_20162,N_20302);
and U21961 (N_21961,N_21643,N_19737);
or U21962 (N_21962,N_21693,N_19932);
xor U21963 (N_21963,N_20939,N_18853);
nand U21964 (N_21964,N_21578,N_20282);
nand U21965 (N_21965,N_19421,N_20345);
nand U21966 (N_21966,N_19612,N_18833);
nor U21967 (N_21967,N_21158,N_20036);
or U21968 (N_21968,N_21263,N_20134);
and U21969 (N_21969,N_21451,N_20130);
nor U21970 (N_21970,N_21195,N_19793);
nand U21971 (N_21971,N_20807,N_19545);
and U21972 (N_21972,N_21794,N_19362);
nor U21973 (N_21973,N_19717,N_19595);
xnor U21974 (N_21974,N_19393,N_21370);
or U21975 (N_21975,N_19428,N_20127);
and U21976 (N_21976,N_21540,N_19406);
and U21977 (N_21977,N_19791,N_20177);
xor U21978 (N_21978,N_20074,N_21704);
xor U21979 (N_21979,N_20187,N_20969);
nand U21980 (N_21980,N_21443,N_18868);
nand U21981 (N_21981,N_20216,N_20644);
xor U21982 (N_21982,N_21188,N_21801);
nor U21983 (N_21983,N_20799,N_18758);
xor U21984 (N_21984,N_19925,N_20112);
nor U21985 (N_21985,N_19179,N_21489);
nor U21986 (N_21986,N_19680,N_19885);
xnor U21987 (N_21987,N_21632,N_20014);
or U21988 (N_21988,N_20871,N_20739);
xnor U21989 (N_21989,N_20999,N_20823);
and U21990 (N_21990,N_20667,N_19685);
nand U21991 (N_21991,N_20033,N_21278);
nor U21992 (N_21992,N_20844,N_18882);
nor U21993 (N_21993,N_21167,N_20210);
and U21994 (N_21994,N_19773,N_19813);
nor U21995 (N_21995,N_19743,N_19617);
xor U21996 (N_21996,N_19534,N_19194);
and U21997 (N_21997,N_20283,N_21442);
and U21998 (N_21998,N_20665,N_19009);
nand U21999 (N_21999,N_19473,N_21502);
nor U22000 (N_22000,N_21244,N_19995);
xnor U22001 (N_22001,N_19560,N_20396);
nor U22002 (N_22002,N_21510,N_20059);
xnor U22003 (N_22003,N_20355,N_18802);
nor U22004 (N_22004,N_20774,N_20547);
nor U22005 (N_22005,N_20458,N_20534);
nand U22006 (N_22006,N_20512,N_21854);
nand U22007 (N_22007,N_18854,N_21328);
nand U22008 (N_22008,N_21267,N_19719);
and U22009 (N_22009,N_20883,N_21210);
xor U22010 (N_22010,N_20888,N_19251);
or U22011 (N_22011,N_20840,N_21565);
nor U22012 (N_22012,N_20673,N_20138);
or U22013 (N_22013,N_21410,N_20633);
nand U22014 (N_22014,N_21378,N_19835);
xnor U22015 (N_22015,N_21160,N_19483);
nor U22016 (N_22016,N_21393,N_21645);
or U22017 (N_22017,N_21501,N_21495);
nor U22018 (N_22018,N_19749,N_20469);
nand U22019 (N_22019,N_21003,N_20504);
and U22020 (N_22020,N_20924,N_20647);
or U22021 (N_22021,N_19706,N_19191);
nor U22022 (N_22022,N_19941,N_19958);
xor U22023 (N_22023,N_21252,N_21027);
nand U22024 (N_22024,N_19624,N_19247);
nor U22025 (N_22025,N_19008,N_20198);
or U22026 (N_22026,N_21726,N_21265);
nor U22027 (N_22027,N_18856,N_19877);
nor U22028 (N_22028,N_21562,N_20347);
and U22029 (N_22029,N_20116,N_20090);
nand U22030 (N_22030,N_20184,N_19227);
nor U22031 (N_22031,N_19721,N_21379);
xor U22032 (N_22032,N_19021,N_21399);
nor U22033 (N_22033,N_21698,N_19738);
nand U22034 (N_22034,N_21775,N_21850);
or U22035 (N_22035,N_21851,N_20315);
nor U22036 (N_22036,N_19084,N_20365);
or U22037 (N_22037,N_19911,N_19383);
or U22038 (N_22038,N_20620,N_21544);
or U22039 (N_22039,N_19267,N_21163);
nand U22040 (N_22040,N_20322,N_20947);
xor U22041 (N_22041,N_18978,N_20502);
or U22042 (N_22042,N_21556,N_19078);
nand U22043 (N_22043,N_21806,N_20151);
xnor U22044 (N_22044,N_20664,N_19699);
nand U22045 (N_22045,N_21215,N_20744);
nor U22046 (N_22046,N_19888,N_19071);
and U22047 (N_22047,N_20728,N_19514);
xor U22048 (N_22048,N_21697,N_19092);
or U22049 (N_22049,N_21612,N_21835);
or U22050 (N_22050,N_19643,N_21295);
nor U22051 (N_22051,N_20532,N_19654);
nand U22052 (N_22052,N_20300,N_21550);
nand U22053 (N_22053,N_18774,N_18945);
and U22054 (N_22054,N_20795,N_20273);
and U22055 (N_22055,N_19777,N_21187);
nor U22056 (N_22056,N_19373,N_20599);
nand U22057 (N_22057,N_19983,N_19712);
and U22058 (N_22058,N_21376,N_20298);
and U22059 (N_22059,N_19036,N_19827);
xnor U22060 (N_22060,N_19166,N_20629);
nor U22061 (N_22061,N_20385,N_20488);
and U22062 (N_22062,N_20949,N_18765);
or U22063 (N_22063,N_19231,N_20256);
and U22064 (N_22064,N_19735,N_21742);
nand U22065 (N_22065,N_19756,N_19219);
xnor U22066 (N_22066,N_20433,N_19100);
nor U22067 (N_22067,N_21535,N_21846);
and U22068 (N_22068,N_21472,N_19067);
or U22069 (N_22069,N_20325,N_21575);
and U22070 (N_22070,N_19808,N_18773);
and U22071 (N_22071,N_20968,N_21637);
xnor U22072 (N_22072,N_20901,N_19196);
xor U22073 (N_22073,N_20526,N_20093);
and U22074 (N_22074,N_20316,N_20580);
or U22075 (N_22075,N_19754,N_18808);
nand U22076 (N_22076,N_21357,N_21153);
xnor U22077 (N_22077,N_21233,N_20145);
or U22078 (N_22078,N_20902,N_20649);
nand U22079 (N_22079,N_19126,N_19410);
or U22080 (N_22080,N_20754,N_18895);
nor U22081 (N_22081,N_21182,N_21641);
nand U22082 (N_22082,N_21091,N_18778);
nand U22083 (N_22083,N_21434,N_20942);
nor U22084 (N_22084,N_19313,N_19081);
nand U22085 (N_22085,N_21327,N_21430);
xnor U22086 (N_22086,N_21108,N_19056);
or U22087 (N_22087,N_21017,N_20096);
nor U22088 (N_22088,N_19867,N_21135);
nand U22089 (N_22089,N_21601,N_19614);
nor U22090 (N_22090,N_19252,N_21712);
nor U22091 (N_22091,N_19847,N_20543);
or U22092 (N_22092,N_21660,N_21174);
or U22093 (N_22093,N_19645,N_18805);
nor U22094 (N_22094,N_21192,N_21555);
nor U22095 (N_22095,N_20593,N_20722);
nor U22096 (N_22096,N_21110,N_19790);
nor U22097 (N_22097,N_21662,N_18981);
nand U22098 (N_22098,N_20715,N_21092);
nand U22099 (N_22099,N_21559,N_19324);
or U22100 (N_22100,N_19921,N_19401);
xnor U22101 (N_22101,N_20480,N_19034);
nor U22102 (N_22102,N_18998,N_21002);
or U22103 (N_22103,N_20231,N_18943);
nand U22104 (N_22104,N_20218,N_21748);
and U22105 (N_22105,N_20657,N_20269);
xor U22106 (N_22106,N_18931,N_19091);
nor U22107 (N_22107,N_19587,N_19446);
xor U22108 (N_22108,N_20082,N_21807);
or U22109 (N_22109,N_19103,N_19954);
and U22110 (N_22110,N_20261,N_20062);
xor U22111 (N_22111,N_19120,N_19297);
nor U22112 (N_22112,N_21008,N_20475);
or U22113 (N_22113,N_21150,N_20358);
and U22114 (N_22114,N_21229,N_21798);
and U22115 (N_22115,N_20822,N_21655);
nand U22116 (N_22116,N_21100,N_18843);
nand U22117 (N_22117,N_20232,N_18800);
or U22118 (N_22118,N_20147,N_20152);
xor U22119 (N_22119,N_19332,N_19639);
or U22120 (N_22120,N_20576,N_21526);
nand U22121 (N_22121,N_18872,N_19445);
or U22122 (N_22122,N_21066,N_20446);
nand U22123 (N_22123,N_20454,N_19355);
xor U22124 (N_22124,N_19183,N_20119);
nand U22125 (N_22125,N_19895,N_20190);
nor U22126 (N_22126,N_19402,N_21419);
or U22127 (N_22127,N_18914,N_20491);
or U22128 (N_22128,N_19659,N_20632);
nand U22129 (N_22129,N_19234,N_20429);
and U22130 (N_22130,N_18803,N_18980);
nand U22131 (N_22131,N_19415,N_18903);
nand U22132 (N_22132,N_19718,N_18814);
xor U22133 (N_22133,N_19107,N_20864);
and U22134 (N_22134,N_19803,N_19934);
xnor U22135 (N_22135,N_21795,N_18947);
or U22136 (N_22136,N_20575,N_19762);
nor U22137 (N_22137,N_20386,N_19096);
nand U22138 (N_22138,N_21421,N_19889);
nand U22139 (N_22139,N_20371,N_19916);
nand U22140 (N_22140,N_21684,N_19499);
xnor U22141 (N_22141,N_19361,N_21009);
nor U22142 (N_22142,N_21083,N_21241);
and U22143 (N_22143,N_21859,N_18852);
or U22144 (N_22144,N_20556,N_20743);
and U22145 (N_22145,N_19359,N_21642);
and U22146 (N_22146,N_20304,N_18787);
or U22147 (N_22147,N_19089,N_20418);
or U22148 (N_22148,N_21487,N_20092);
xor U22149 (N_22149,N_18875,N_19554);
or U22150 (N_22150,N_20579,N_18789);
or U22151 (N_22151,N_20444,N_20697);
and U22152 (N_22152,N_20565,N_19632);
xor U22153 (N_22153,N_21185,N_20186);
xor U22154 (N_22154,N_19044,N_21577);
nand U22155 (N_22155,N_19691,N_19600);
nor U22156 (N_22156,N_21773,N_18954);
nor U22157 (N_22157,N_21067,N_19530);
nand U22158 (N_22158,N_19837,N_21063);
nor U22159 (N_22159,N_19669,N_21222);
and U22160 (N_22160,N_18909,N_21424);
nor U22161 (N_22161,N_19854,N_19424);
and U22162 (N_22162,N_19379,N_20212);
xor U22163 (N_22163,N_20317,N_19215);
nor U22164 (N_22164,N_20609,N_21767);
and U22165 (N_22165,N_21763,N_19209);
and U22166 (N_22166,N_20910,N_20230);
xor U22167 (N_22167,N_20791,N_20340);
nand U22168 (N_22168,N_20417,N_19615);
xor U22169 (N_22169,N_19476,N_19802);
xnor U22170 (N_22170,N_21628,N_19832);
and U22171 (N_22171,N_21533,N_21258);
and U22172 (N_22172,N_18851,N_20787);
and U22173 (N_22173,N_20415,N_21574);
and U22174 (N_22174,N_19556,N_19013);
xor U22175 (N_22175,N_21608,N_19070);
and U22176 (N_22176,N_19290,N_19858);
nand U22177 (N_22177,N_21784,N_21203);
xnor U22178 (N_22178,N_19642,N_19063);
nand U22179 (N_22179,N_21867,N_21676);
nand U22180 (N_22180,N_21057,N_20018);
xor U22181 (N_22181,N_20628,N_21124);
or U22182 (N_22182,N_20887,N_20197);
nor U22183 (N_22183,N_21096,N_18997);
nand U22184 (N_22184,N_20792,N_19960);
or U22185 (N_22185,N_20984,N_19482);
nand U22186 (N_22186,N_20615,N_20221);
and U22187 (N_22187,N_18942,N_20439);
nand U22188 (N_22188,N_20351,N_20276);
xor U22189 (N_22189,N_20817,N_21583);
nor U22190 (N_22190,N_21152,N_19507);
xnor U22191 (N_22191,N_19581,N_18993);
or U22192 (N_22192,N_19681,N_21372);
xor U22193 (N_22193,N_19337,N_18863);
nor U22194 (N_22194,N_19391,N_21193);
and U22195 (N_22195,N_20794,N_20160);
and U22196 (N_22196,N_19539,N_19299);
and U22197 (N_22197,N_20003,N_19779);
xnor U22198 (N_22198,N_21142,N_19169);
nor U22199 (N_22199,N_19647,N_19105);
and U22200 (N_22200,N_19080,N_19378);
nand U22201 (N_22201,N_19936,N_21687);
or U22202 (N_22202,N_18873,N_20986);
nor U22203 (N_22203,N_19564,N_21144);
or U22204 (N_22204,N_19187,N_21441);
nand U22205 (N_22205,N_21246,N_21130);
nor U22206 (N_22206,N_20622,N_20012);
xnor U22207 (N_22207,N_20496,N_19883);
and U22208 (N_22208,N_19478,N_21123);
xnor U22209 (N_22209,N_21553,N_21852);
nand U22210 (N_22210,N_18988,N_19452);
nand U22211 (N_22211,N_20436,N_19613);
nor U22212 (N_22212,N_20084,N_19351);
or U22213 (N_22213,N_20603,N_21848);
and U22214 (N_22214,N_21254,N_19277);
and U22215 (N_22215,N_19824,N_20594);
and U22216 (N_22216,N_19734,N_19838);
nand U22217 (N_22217,N_20703,N_18766);
nand U22218 (N_22218,N_21599,N_19714);
nor U22219 (N_22219,N_19553,N_20372);
nor U22220 (N_22220,N_20132,N_21548);
nand U22221 (N_22221,N_21082,N_19479);
nor U22222 (N_22222,N_21871,N_18920);
xor U22223 (N_22223,N_20827,N_21631);
nor U22224 (N_22224,N_19238,N_21745);
nor U22225 (N_22225,N_21165,N_21355);
nand U22226 (N_22226,N_19990,N_19555);
xor U22227 (N_22227,N_21262,N_21728);
or U22228 (N_22228,N_20802,N_20363);
and U22229 (N_22229,N_21560,N_19968);
nand U22230 (N_22230,N_19640,N_19920);
nor U22231 (N_22231,N_20627,N_21311);
nor U22232 (N_22232,N_19938,N_19869);
nor U22233 (N_22233,N_19900,N_20809);
or U22234 (N_22234,N_19692,N_21166);
nor U22235 (N_22235,N_20983,N_19577);
nand U22236 (N_22236,N_20234,N_21061);
nor U22237 (N_22237,N_20885,N_19578);
xnor U22238 (N_22238,N_20252,N_20597);
and U22239 (N_22239,N_20611,N_21216);
xor U22240 (N_22240,N_19757,N_20912);
and U22241 (N_22241,N_18822,N_21146);
or U22242 (N_22242,N_20349,N_21346);
nor U22243 (N_22243,N_18860,N_20228);
or U22244 (N_22244,N_20878,N_20660);
nand U22245 (N_22245,N_20803,N_19666);
or U22246 (N_22246,N_18968,N_19197);
or U22247 (N_22247,N_19407,N_18831);
nand U22248 (N_22248,N_19074,N_20068);
xnor U22249 (N_22249,N_21870,N_21672);
and U22250 (N_22250,N_21080,N_21266);
or U22251 (N_22251,N_19135,N_21514);
nand U22252 (N_22252,N_21316,N_20843);
or U22253 (N_22253,N_20324,N_21321);
nand U22254 (N_22254,N_20606,N_19149);
xor U22255 (N_22255,N_19167,N_19146);
nor U22256 (N_22256,N_20847,N_21329);
nand U22257 (N_22257,N_19511,N_20054);
and U22258 (N_22258,N_21711,N_21084);
nor U22259 (N_22259,N_21161,N_19134);
xor U22260 (N_22260,N_20762,N_21300);
nand U22261 (N_22261,N_20207,N_21116);
or U22262 (N_22262,N_20247,N_18964);
and U22263 (N_22263,N_20689,N_21837);
or U22264 (N_22264,N_20487,N_20845);
or U22265 (N_22265,N_18820,N_20944);
and U22266 (N_22266,N_20044,N_21006);
and U22267 (N_22267,N_18771,N_21758);
nor U22268 (N_22268,N_18816,N_21199);
and U22269 (N_22269,N_19772,N_19819);
xnor U22270 (N_22270,N_21012,N_21243);
or U22271 (N_22271,N_19398,N_19804);
or U22272 (N_22272,N_19006,N_21214);
or U22273 (N_22273,N_18784,N_21611);
nor U22274 (N_22274,N_20434,N_20500);
or U22275 (N_22275,N_20163,N_20208);
or U22276 (N_22276,N_19912,N_20677);
nand U22277 (N_22277,N_20017,N_21024);
and U22278 (N_22278,N_19696,N_20626);
and U22279 (N_22279,N_19245,N_19890);
or U22280 (N_22280,N_19023,N_21816);
and U22281 (N_22281,N_19592,N_20956);
nand U22282 (N_22282,N_21168,N_20863);
xnor U22283 (N_22283,N_21202,N_18930);
xnor U22284 (N_22284,N_21387,N_20834);
or U22285 (N_22285,N_21179,N_19872);
or U22286 (N_22286,N_19720,N_21593);
nor U22287 (N_22287,N_19704,N_20494);
nand U22288 (N_22288,N_21511,N_21772);
xor U22289 (N_22289,N_18936,N_19836);
nand U22290 (N_22290,N_18900,N_19865);
or U22291 (N_22291,N_21029,N_18837);
or U22292 (N_22292,N_20118,N_20708);
xor U22293 (N_22293,N_19745,N_21366);
nor U22294 (N_22294,N_19235,N_20011);
nor U22295 (N_22295,N_20442,N_18965);
xnor U22296 (N_22296,N_21480,N_21765);
and U22297 (N_22297,N_20546,N_21230);
nand U22298 (N_22298,N_19420,N_19068);
nand U22299 (N_22299,N_20759,N_19580);
and U22300 (N_22300,N_21070,N_21668);
xor U22301 (N_22301,N_21204,N_19296);
or U22302 (N_22302,N_19985,N_20671);
xnor U22303 (N_22303,N_20106,N_20961);
or U22304 (N_22304,N_19760,N_18761);
nand U22305 (N_22305,N_21171,N_21739);
nor U22306 (N_22306,N_21189,N_20165);
or U22307 (N_22307,N_19657,N_21743);
xnor U22308 (N_22308,N_20188,N_19675);
xnor U22309 (N_22309,N_19287,N_19820);
and U22310 (N_22310,N_21075,N_21358);
nand U22311 (N_22311,N_20652,N_21280);
or U22312 (N_22312,N_20449,N_19340);
nand U22313 (N_22313,N_21445,N_19255);
and U22314 (N_22314,N_21496,N_21383);
xor U22315 (N_22315,N_20185,N_19102);
or U22316 (N_22316,N_21680,N_19533);
or U22317 (N_22317,N_19891,N_21573);
or U22318 (N_22318,N_20521,N_21112);
xor U22319 (N_22319,N_18880,N_21497);
and U22320 (N_22320,N_20732,N_19432);
xor U22321 (N_22321,N_21076,N_19250);
nand U22322 (N_22322,N_19599,N_21038);
nor U22323 (N_22323,N_20080,N_18881);
nor U22324 (N_22324,N_20478,N_21609);
xor U22325 (N_22325,N_21058,N_21607);
and U22326 (N_22326,N_21094,N_19522);
and U22327 (N_22327,N_19879,N_20600);
xnor U22328 (N_22328,N_18915,N_19970);
nand U22329 (N_22329,N_20701,N_21623);
nand U22330 (N_22330,N_20955,N_19101);
and U22331 (N_22331,N_21342,N_20966);
xor U22332 (N_22332,N_20568,N_21277);
nor U22333 (N_22333,N_19831,N_20022);
nand U22334 (N_22334,N_20957,N_20214);
or U22335 (N_22335,N_20587,N_20945);
nor U22336 (N_22336,N_19025,N_20004);
nand U22337 (N_22337,N_21242,N_21585);
nand U22338 (N_22338,N_21799,N_21395);
nand U22339 (N_22339,N_21841,N_19605);
or U22340 (N_22340,N_19517,N_19136);
nand U22341 (N_22341,N_21572,N_20306);
and U22342 (N_22342,N_21156,N_18764);
nor U22343 (N_22343,N_20217,N_19771);
or U22344 (N_22344,N_20167,N_20811);
nor U22345 (N_22345,N_18982,N_19759);
nand U22346 (N_22346,N_20369,N_20111);
xnor U22347 (N_22347,N_19739,N_19846);
nand U22348 (N_22348,N_21125,N_20233);
or U22349 (N_22349,N_20206,N_19602);
nor U22350 (N_22350,N_20836,N_21308);
xor U22351 (N_22351,N_20426,N_20916);
nor U22352 (N_22352,N_21730,N_19529);
xnor U22353 (N_22353,N_20909,N_19468);
or U22354 (N_22354,N_21385,N_20113);
and U22355 (N_22355,N_21671,N_20000);
xnor U22356 (N_22356,N_20456,N_21296);
nand U22357 (N_22357,N_21454,N_21833);
xnor U22358 (N_22358,N_18767,N_20931);
nand U22359 (N_22359,N_20146,N_19782);
or U22360 (N_22360,N_19236,N_19174);
nor U22361 (N_22361,N_21041,N_19040);
and U22362 (N_22362,N_19341,N_19904);
or U22363 (N_22363,N_20522,N_21808);
nor U22364 (N_22364,N_18966,N_20785);
or U22365 (N_22365,N_21785,N_21255);
nor U22366 (N_22366,N_19948,N_19598);
xnor U22367 (N_22367,N_20636,N_21087);
and U22368 (N_22368,N_21136,N_19440);
nor U22369 (N_22369,N_20295,N_20007);
nor U22370 (N_22370,N_19147,N_18855);
or U22371 (N_22371,N_21670,N_19032);
nor U22372 (N_22372,N_18905,N_20566);
xnor U22373 (N_22373,N_20164,N_21172);
xnor U22374 (N_22374,N_21756,N_21413);
nand U22375 (N_22375,N_21440,N_20914);
xnor U22376 (N_22376,N_19060,N_20737);
nor U22377 (N_22377,N_18937,N_19404);
nand U22378 (N_22378,N_21863,N_18812);
and U22379 (N_22379,N_19128,N_21732);
nand U22380 (N_22380,N_20943,N_21839);
xor U22381 (N_22381,N_20923,N_21449);
or U22382 (N_22382,N_20245,N_19015);
nor U22383 (N_22383,N_20101,N_19342);
nor U22384 (N_22384,N_19653,N_20510);
nor U22385 (N_22385,N_19184,N_19656);
nor U22386 (N_22386,N_19957,N_20225);
nor U22387 (N_22387,N_21060,N_19783);
xor U22388 (N_22388,N_19730,N_20189);
nand U22389 (N_22389,N_20352,N_20029);
nor U22390 (N_22390,N_21486,N_21858);
xnor U22391 (N_22391,N_19937,N_18754);
nand U22392 (N_22392,N_20890,N_21138);
nor U22393 (N_22393,N_19180,N_21314);
nor U22394 (N_22394,N_20621,N_18834);
nor U22395 (N_22395,N_19312,N_20406);
or U22396 (N_22396,N_20815,N_20490);
or U22397 (N_22397,N_21755,N_21129);
or U22398 (N_22398,N_20061,N_21538);
nor U22399 (N_22399,N_18973,N_21019);
nand U22400 (N_22400,N_21426,N_18885);
xor U22401 (N_22401,N_20440,N_21004);
and U22402 (N_22402,N_19388,N_20631);
nor U22403 (N_22403,N_21664,N_20158);
and U22404 (N_22404,N_19979,N_19368);
or U22405 (N_22405,N_21117,N_21630);
xor U22406 (N_22406,N_20675,N_20318);
nor U22407 (N_22407,N_19649,N_20798);
or U22408 (N_22408,N_19043,N_19998);
nand U22409 (N_22409,N_19818,N_19943);
and U22410 (N_22410,N_21792,N_19956);
or U22411 (N_22411,N_21201,N_21460);
nor U22412 (N_22412,N_21081,N_20640);
and U22413 (N_22413,N_19335,N_19626);
or U22414 (N_22414,N_20858,N_21805);
nand U22415 (N_22415,N_20805,N_19076);
xnor U22416 (N_22416,N_19292,N_20368);
and U22417 (N_22417,N_19281,N_20953);
xnor U22418 (N_22418,N_19205,N_20810);
and U22419 (N_22419,N_19786,N_20288);
nor U22420 (N_22420,N_20353,N_20934);
or U22421 (N_22421,N_21789,N_21523);
xor U22422 (N_22422,N_18925,N_19246);
nand U22423 (N_22423,N_20094,N_18775);
or U22424 (N_22424,N_19124,N_21145);
and U22425 (N_22425,N_21531,N_19300);
nand U22426 (N_22426,N_18976,N_19789);
xnor U22427 (N_22427,N_19487,N_18756);
xnor U22428 (N_22428,N_20244,N_20872);
xnor U22429 (N_22429,N_19384,N_21218);
xnor U22430 (N_22430,N_21465,N_21053);
nor U22431 (N_22431,N_21825,N_20495);
and U22432 (N_22432,N_20884,N_18870);
and U22433 (N_22433,N_21250,N_19797);
nand U22434 (N_22434,N_19241,N_19119);
nand U22435 (N_22435,N_20296,N_20076);
nand U22436 (N_22436,N_19798,N_19200);
xnor U22437 (N_22437,N_20833,N_20849);
or U22438 (N_22438,N_20963,N_20419);
xnor U22439 (N_22439,N_19748,N_21751);
and U22440 (N_22440,N_21580,N_20978);
and U22441 (N_22441,N_19327,N_19376);
nand U22442 (N_22442,N_19139,N_19710);
nor U22443 (N_22443,N_21119,N_18847);
nand U22444 (N_22444,N_18751,N_19058);
nand U22445 (N_22445,N_20908,N_21779);
xor U22446 (N_22446,N_21731,N_20242);
nor U22447 (N_22447,N_21864,N_21734);
xnor U22448 (N_22448,N_20723,N_21521);
nor U22449 (N_22449,N_19908,N_19766);
xor U22450 (N_22450,N_18874,N_19480);
xnor U22451 (N_22451,N_19559,N_21159);
nand U22452 (N_22452,N_19334,N_20882);
or U22453 (N_22453,N_19018,N_19641);
xor U22454 (N_22454,N_20720,N_20555);
xor U22455 (N_22455,N_21054,N_19426);
xor U22456 (N_22456,N_21702,N_19417);
or U22457 (N_22457,N_19907,N_20196);
xor U22458 (N_22458,N_19024,N_20896);
nor U22459 (N_22459,N_20875,N_21015);
and U22460 (N_22460,N_20987,N_19352);
nand U22461 (N_22461,N_20241,N_21536);
and U22462 (N_22462,N_21062,N_18795);
nand U22463 (N_22463,N_19863,N_19309);
and U22464 (N_22464,N_20125,N_21845);
or U22465 (N_22465,N_18957,N_21679);
and U22466 (N_22466,N_21394,N_20049);
nand U22467 (N_22467,N_19942,N_18919);
and U22468 (N_22468,N_21014,N_21115);
nand U22469 (N_22469,N_20281,N_19073);
xor U22470 (N_22470,N_18779,N_20069);
nor U22471 (N_22471,N_19413,N_19303);
and U22472 (N_22472,N_18752,N_21422);
xnor U22473 (N_22473,N_20203,N_21005);
and U22474 (N_22474,N_19216,N_21427);
and U22475 (N_22475,N_21500,N_19991);
nor U22476 (N_22476,N_20060,N_20224);
nor U22477 (N_22477,N_21823,N_20143);
xor U22478 (N_22478,N_19849,N_18844);
xnor U22479 (N_22479,N_19503,N_19069);
or U22480 (N_22480,N_20258,N_19301);
and U22481 (N_22481,N_21738,N_20481);
and U22482 (N_22482,N_20782,N_20209);
and U22483 (N_22483,N_20309,N_21306);
nand U22484 (N_22484,N_18827,N_20178);
and U22485 (N_22485,N_19217,N_21817);
nor U22486 (N_22486,N_19099,N_20451);
xor U22487 (N_22487,N_18926,N_20327);
and U22488 (N_22488,N_21834,N_19506);
nor U22489 (N_22489,N_20540,N_21812);
nor U22490 (N_22490,N_20305,N_19011);
xor U22491 (N_22491,N_18970,N_20686);
or U22492 (N_22492,N_19812,N_19585);
nor U22493 (N_22493,N_20243,N_21821);
or U22494 (N_22494,N_21284,N_19291);
xor U22495 (N_22495,N_21045,N_18794);
nand U22496 (N_22496,N_20289,N_20520);
xnor U22497 (N_22497,N_21477,N_19801);
nand U22498 (N_22498,N_21287,N_21516);
nand U22499 (N_22499,N_21813,N_19346);
and U22500 (N_22500,N_19392,N_19927);
or U22501 (N_22501,N_19448,N_21595);
xor U22502 (N_22502,N_20467,N_19331);
nand U22503 (N_22503,N_18924,N_18782);
nor U22504 (N_22504,N_21409,N_21557);
nor U22505 (N_22505,N_21588,N_19423);
xor U22506 (N_22506,N_19129,N_21558);
or U22507 (N_22507,N_19333,N_19319);
and U22508 (N_22508,N_20174,N_21473);
nor U22509 (N_22509,N_19672,N_21175);
nor U22510 (N_22510,N_19727,N_19109);
or U22511 (N_22511,N_21418,N_20337);
nand U22512 (N_22512,N_20095,N_21797);
xnor U22513 (N_22513,N_20559,N_21626);
xor U22514 (N_22514,N_21097,N_19386);
xor U22515 (N_22515,N_19633,N_21272);
or U22516 (N_22516,N_19809,N_19016);
nand U22517 (N_22517,N_19862,N_19151);
or U22518 (N_22518,N_21274,N_20161);
and U22519 (N_22519,N_21788,N_20874);
xor U22520 (N_22520,N_20483,N_21722);
nor U22521 (N_22521,N_20015,N_21302);
xor U22522 (N_22522,N_20235,N_20468);
nor U22523 (N_22523,N_18958,N_20523);
nand U22524 (N_22524,N_21856,N_19795);
and U22525 (N_22525,N_21757,N_19986);
xor U22526 (N_22526,N_19510,N_18867);
nand U22527 (N_22527,N_20573,N_21333);
xor U22528 (N_22528,N_19924,N_19226);
nor U22529 (N_22529,N_19492,N_20179);
nor U22530 (N_22530,N_19520,N_21483);
xnor U22531 (N_22531,N_19075,N_18932);
nor U22532 (N_22532,N_21071,N_21291);
xor U22533 (N_22533,N_21853,N_20893);
nand U22534 (N_22534,N_21431,N_20042);
nand U22535 (N_22535,N_19248,N_20925);
xor U22536 (N_22536,N_20422,N_20990);
and U22537 (N_22537,N_20745,N_21724);
or U22538 (N_22538,N_21667,N_21085);
nor U22539 (N_22539,N_20670,N_20357);
and U22540 (N_22540,N_19501,N_21035);
xnor U22541 (N_22541,N_21353,N_19946);
or U22542 (N_22542,N_19026,N_19558);
xor U22543 (N_22543,N_21597,N_19419);
and U22544 (N_22544,N_21563,N_20506);
or U22545 (N_22545,N_21542,N_21719);
nor U22546 (N_22546,N_18955,N_21417);
or U22547 (N_22547,N_20006,N_18783);
nor U22548 (N_22548,N_19265,N_18755);
or U22549 (N_22549,N_20085,N_19919);
nand U22550 (N_22550,N_20360,N_21319);
nor U22551 (N_22551,N_20537,N_19121);
xor U22552 (N_22552,N_20181,N_19072);
xnor U22553 (N_22553,N_20099,N_19210);
xnor U22554 (N_22554,N_18876,N_20895);
xnor U22555 (N_22555,N_20738,N_21143);
nor U22556 (N_22556,N_20279,N_21855);
nand U22557 (N_22557,N_20614,N_19037);
xnor U22558 (N_22558,N_20486,N_21777);
and U22559 (N_22559,N_21782,N_19993);
nor U22560 (N_22560,N_19079,N_19972);
nor U22561 (N_22561,N_19565,N_20040);
or U22562 (N_22562,N_21453,N_20574);
nand U22563 (N_22563,N_20173,N_20117);
or U22564 (N_22564,N_20974,N_18776);
and U22565 (N_22565,N_20391,N_19962);
nand U22566 (N_22566,N_19316,N_20868);
and U22567 (N_22567,N_20714,N_21508);
xnor U22568 (N_22568,N_21715,N_19671);
or U22569 (N_22569,N_21186,N_20717);
nor U22570 (N_22570,N_21350,N_20694);
or U22571 (N_22571,N_18829,N_20753);
nor U22572 (N_22572,N_19170,N_18790);
xnor U22573 (N_22573,N_21769,N_20826);
and U22574 (N_22574,N_19387,N_20374);
xnor U22575 (N_22575,N_20830,N_21570);
nand U22576 (N_22576,N_19750,N_19033);
nor U22577 (N_22577,N_20519,N_19778);
or U22578 (N_22578,N_19322,N_20104);
or U22579 (N_22579,N_21561,N_19769);
nand U22580 (N_22580,N_18826,N_19389);
or U22581 (N_22581,N_19017,N_20747);
xnor U22582 (N_22582,N_21122,N_19896);
xor U22583 (N_22583,N_20515,N_18990);
nor U22584 (N_22584,N_21567,N_20052);
xnor U22585 (N_22585,N_21640,N_20331);
nor U22586 (N_22586,N_19019,N_18845);
xor U22587 (N_22587,N_20031,N_19542);
nor U22588 (N_22588,N_21371,N_20402);
xnor U22589 (N_22589,N_19755,N_19055);
nor U22590 (N_22590,N_20428,N_18952);
and U22591 (N_22591,N_20412,N_19354);
nand U22592 (N_22592,N_20026,N_19965);
nand U22593 (N_22593,N_19917,N_19459);
or U22594 (N_22594,N_19780,N_21666);
nand U22595 (N_22595,N_20706,N_21030);
xor U22596 (N_22596,N_21530,N_18963);
xor U22597 (N_22597,N_19467,N_21444);
and U22598 (N_22598,N_19631,N_21546);
or U22599 (N_22599,N_19221,N_21809);
xnor U22600 (N_22600,N_20548,N_21253);
nand U22601 (N_22601,N_19083,N_19288);
and U22602 (N_22602,N_19022,N_19242);
and U22603 (N_22603,N_19283,N_20585);
nand U22604 (N_22604,N_21078,N_19618);
nor U22605 (N_22605,N_20191,N_20255);
or U22606 (N_22606,N_19593,N_20048);
and U22607 (N_22607,N_18923,N_18888);
or U22608 (N_22608,N_21169,N_21866);
nand U22609 (N_22609,N_19949,N_20320);
xor U22610 (N_22610,N_20416,N_21121);
nor U22611 (N_22611,N_20997,N_19842);
nand U22612 (N_22612,N_20857,N_21857);
xor U22613 (N_22613,N_20618,N_21543);
and U22614 (N_22614,N_20666,N_21055);
or U22615 (N_22615,N_20950,N_20470);
nand U22616 (N_22616,N_18780,N_19550);
xor U22617 (N_22617,N_19973,N_19254);
nand U22618 (N_22618,N_21541,N_20828);
xnor U22619 (N_22619,N_18953,N_21235);
or U22620 (N_22620,N_19039,N_20590);
nor U22621 (N_22621,N_21686,N_21648);
nor U22622 (N_22622,N_20493,N_20270);
nor U22623 (N_22623,N_19115,N_19770);
or U22624 (N_22624,N_18788,N_21804);
nand U22625 (N_22625,N_19422,N_18967);
or U22626 (N_22626,N_21206,N_21663);
nor U22627 (N_22627,N_20598,N_19344);
or U22628 (N_22628,N_18994,N_21847);
nand U22629 (N_22629,N_20772,N_20977);
xnor U22630 (N_22630,N_20550,N_19722);
nand U22631 (N_22631,N_19027,N_19271);
and U22632 (N_22632,N_21582,N_20139);
or U22633 (N_22633,N_21104,N_19996);
nor U22634 (N_22634,N_21707,N_20405);
nor U22635 (N_22635,N_20913,N_21634);
nand U22636 (N_22636,N_20257,N_19686);
nor U22637 (N_22637,N_19481,N_20808);
xor U22638 (N_22638,N_19257,N_21820);
nand U22639 (N_22639,N_21408,N_20321);
nand U22640 (N_22640,N_19029,N_21231);
nand U22641 (N_22641,N_20904,N_20812);
or U22642 (N_22642,N_20328,N_19561);
nor U22643 (N_22643,N_19364,N_20648);
and U22644 (N_22644,N_21047,N_19850);
xnor U22645 (N_22645,N_20514,N_21729);
nand U22646 (N_22646,N_19400,N_20727);
nor U22647 (N_22647,N_19703,N_19190);
xnor U22648 (N_22648,N_21354,N_20420);
and U22649 (N_22649,N_19390,N_21764);
nand U22650 (N_22650,N_20569,N_19548);
nor U22651 (N_22651,N_21324,N_21584);
or U22652 (N_22652,N_21703,N_19792);
xor U22653 (N_22653,N_19897,N_20343);
xor U22654 (N_22654,N_20334,N_19207);
nor U22655 (N_22655,N_21793,N_18861);
nand U22656 (N_22656,N_20081,N_20940);
nand U22657 (N_22657,N_19630,N_19876);
or U22658 (N_22658,N_20459,N_19571);
or U22659 (N_22659,N_18908,N_20927);
xnor U22660 (N_22660,N_19787,N_20586);
nand U22661 (N_22661,N_21840,N_18769);
and U22662 (N_22662,N_19610,N_19683);
nand U22663 (N_22663,N_18901,N_21681);
nand U22664 (N_22664,N_18753,N_20065);
and U22665 (N_22665,N_19110,N_21259);
nor U22666 (N_22666,N_21690,N_21844);
nor U22667 (N_22667,N_20064,N_20102);
xor U22668 (N_22668,N_19484,N_19674);
or U22669 (N_22669,N_19512,N_21436);
and U22670 (N_22670,N_19321,N_20423);
nand U22671 (N_22671,N_19882,N_19747);
nand U22672 (N_22672,N_21650,N_19318);
xnor U22673 (N_22673,N_21627,N_19161);
and U22674 (N_22674,N_19358,N_19878);
xnor U22675 (N_22675,N_19570,N_20886);
xnor U22676 (N_22676,N_21456,N_20583);
and U22677 (N_22677,N_21382,N_19302);
xnor U22678 (N_22678,N_21768,N_21139);
nor U22679 (N_22679,N_20356,N_20183);
nand U22680 (N_22680,N_20563,N_21299);
nor U22681 (N_22681,N_20581,N_20891);
or U22682 (N_22682,N_19014,N_18877);
xor U22683 (N_22683,N_21073,N_21537);
nand U22684 (N_22684,N_20153,N_21450);
xnor U22685 (N_22685,N_19269,N_21471);
nand U22686 (N_22686,N_19584,N_20635);
nor U22687 (N_22687,N_18939,N_19611);
and U22688 (N_22688,N_19987,N_20024);
xnor U22689 (N_22689,N_19412,N_20776);
nand U22690 (N_22690,N_21181,N_20839);
xor U22691 (N_22691,N_20124,N_20704);
and U22692 (N_22692,N_19774,N_20239);
and U22693 (N_22693,N_19329,N_20175);
or U22694 (N_22694,N_19918,N_21056);
and U22695 (N_22695,N_21312,N_20935);
nor U22696 (N_22696,N_20952,N_19589);
xnor U22697 (N_22697,N_18892,N_20602);
and U22698 (N_22698,N_21692,N_21701);
nor U22699 (N_22699,N_19425,N_18777);
or U22700 (N_22700,N_19687,N_21658);
or U22701 (N_22701,N_20457,N_19243);
nor U22702 (N_22702,N_20960,N_19266);
xor U22703 (N_22703,N_19122,N_20951);
xor U22704 (N_22704,N_19339,N_20105);
xor U22705 (N_22705,N_20250,N_19239);
or U22706 (N_22706,N_21594,N_18887);
nor U22707 (N_22707,N_20564,N_20272);
xnor U22708 (N_22708,N_20786,N_19218);
nor U22709 (N_22709,N_20274,N_21025);
or U22710 (N_22710,N_20149,N_18797);
or U22711 (N_22711,N_21398,N_20169);
or U22712 (N_22712,N_18956,N_19488);
nand U22713 (N_22713,N_20761,N_19676);
and U22714 (N_22714,N_20877,N_21260);
xnor U22715 (N_22715,N_20341,N_20057);
and U22716 (N_22716,N_19338,N_19526);
nor U22717 (N_22717,N_20122,N_20370);
and U22718 (N_22718,N_18858,N_21310);
and U22719 (N_22719,N_19323,N_19214);
and U22720 (N_22720,N_20441,N_18886);
nor U22721 (N_22721,N_20696,N_20605);
nand U22722 (N_22722,N_21197,N_20922);
nand U22723 (N_22723,N_18946,N_20509);
or U22724 (N_22724,N_20364,N_18878);
nor U22725 (N_22725,N_19223,N_21800);
nand U22726 (N_22726,N_19284,N_19208);
nand U22727 (N_22727,N_20637,N_20039);
nor U22728 (N_22728,N_18935,N_21842);
nand U22729 (N_22729,N_21524,N_20853);
and U22730 (N_22730,N_20539,N_19707);
xnor U22731 (N_22731,N_20135,N_20824);
xnor U22732 (N_22732,N_20109,N_20608);
xor U22733 (N_22733,N_19172,N_20424);
nand U22734 (N_22734,N_21271,N_19276);
nor U22735 (N_22735,N_20700,N_20814);
or U22736 (N_22736,N_21293,N_20870);
xnor U22737 (N_22737,N_20200,N_19736);
or U22738 (N_22738,N_19489,N_20879);
xnor U22739 (N_22739,N_20034,N_19186);
or U22740 (N_22740,N_19212,N_21815);
nand U22741 (N_22741,N_21219,N_19673);
and U22742 (N_22742,N_21683,N_19429);
nand U22743 (N_22743,N_20989,N_21155);
nor U22744 (N_22744,N_21007,N_21141);
xnor U22745 (N_22745,N_20395,N_20825);
or U22746 (N_22746,N_20653,N_19601);
nor U22747 (N_22747,N_19603,N_20985);
nand U22748 (N_22748,N_19066,N_20959);
nand U22749 (N_22749,N_19298,N_20375);
nand U22750 (N_22750,N_20280,N_21437);
nand U22751 (N_22751,N_21198,N_19272);
or U22752 (N_22752,N_20756,N_19353);
xnor U22753 (N_22753,N_21787,N_20513);
nor U22754 (N_22754,N_20508,N_21647);
xor U22755 (N_22755,N_19974,N_21037);
nand U22756 (N_22756,N_20361,N_19887);
and U22757 (N_22757,N_19093,N_19955);
xor U22758 (N_22758,N_20610,N_20479);
nor U22759 (N_22759,N_21170,N_19670);
xnor U22760 (N_22760,N_21613,N_21485);
and U22761 (N_22761,N_19546,N_19929);
xor U22762 (N_22762,N_19853,N_20841);
nor U22763 (N_22763,N_21753,N_19045);
xnor U22764 (N_22764,N_19143,N_19967);
nand U22765 (N_22765,N_20971,N_20612);
nor U22766 (N_22766,N_20002,N_18796);
nor U22767 (N_22767,N_21001,N_21470);
nor U22768 (N_22768,N_21388,N_20379);
or U22769 (N_22769,N_21330,N_21771);
nor U22770 (N_22770,N_19188,N_20435);
nand U22771 (N_22771,N_21826,N_19052);
or U22772 (N_22772,N_18977,N_20382);
or U22773 (N_22773,N_21022,N_21482);
and U22774 (N_22774,N_20461,N_19588);
nor U22775 (N_22775,N_19516,N_20170);
nor U22776 (N_22776,N_18969,N_20290);
nor U22777 (N_22777,N_21488,N_20979);
xnor U22778 (N_22778,N_18770,N_20507);
nor U22779 (N_22779,N_21468,N_19365);
or U22780 (N_22780,N_19677,N_19892);
xnor U22781 (N_22781,N_21042,N_21120);
nand U22782 (N_22782,N_19463,N_21873);
and U22783 (N_22783,N_19751,N_21827);
nor U22784 (N_22784,N_18759,N_21475);
nand U22785 (N_22785,N_19947,N_21513);
or U22786 (N_22786,N_20903,N_20030);
nand U22787 (N_22787,N_20680,N_18825);
or U22788 (N_22788,N_19621,N_20505);
nand U22789 (N_22789,N_21478,N_21766);
or U22790 (N_22790,N_21190,N_20323);
and U22791 (N_22791,N_21428,N_21089);
nand U22792 (N_22792,N_19224,N_20623);
xnor U22793 (N_22793,N_19651,N_19449);
xnor U22794 (N_22794,N_20398,N_19154);
nand U22795 (N_22795,N_21320,N_20293);
and U22796 (N_22796,N_18762,N_20854);
and U22797 (N_22797,N_19475,N_18893);
nor U22798 (N_22798,N_19622,N_20707);
nand U22799 (N_22799,N_19396,N_20431);
or U22800 (N_22800,N_19472,N_20268);
nand U22801 (N_22801,N_19969,N_19233);
nor U22802 (N_22802,N_19825,N_21339);
and U22803 (N_22803,N_21046,N_21822);
and U22804 (N_22804,N_19372,N_20716);
nor U22805 (N_22805,N_19811,N_21778);
and U22806 (N_22806,N_19142,N_20748);
and U22807 (N_22807,N_21699,N_19563);
and U22808 (N_22808,N_20894,N_18913);
nor U22809 (N_22809,N_20645,N_20110);
nor U22810 (N_22810,N_20933,N_20915);
or U22811 (N_22811,N_21525,N_21245);
and U22812 (N_22812,N_21286,N_20088);
or U22813 (N_22813,N_19438,N_18987);
xnor U22814 (N_22814,N_21685,N_20781);
nand U22815 (N_22815,N_19688,N_19397);
or U22816 (N_22816,N_21162,N_21036);
xnor U22817 (N_22817,N_20752,N_20695);
nor U22818 (N_22818,N_20777,N_21093);
and U22819 (N_22819,N_19716,N_21247);
nor U22820 (N_22820,N_19596,N_20936);
nand U22821 (N_22821,N_19116,N_21288);
and U22822 (N_22822,N_21600,N_20784);
or U22823 (N_22823,N_19903,N_21332);
or U22824 (N_22824,N_21695,N_19667);
nor U22825 (N_22825,N_21180,N_19086);
nor U22826 (N_22826,N_21708,N_18975);
xor U22827 (N_22827,N_20277,N_21571);
nor U22828 (N_22828,N_19306,N_21814);
nor U22829 (N_22829,N_20733,N_19249);
xor U22830 (N_22830,N_19758,N_19551);
nand U22831 (N_22831,N_19175,N_19204);
and U22832 (N_22832,N_18989,N_20538);
or U22833 (N_22833,N_18944,N_19450);
or U22834 (N_22834,N_19586,N_19765);
xnor U22835 (N_22835,N_19491,N_21043);
nor U22836 (N_22836,N_19304,N_19521);
xor U22837 (N_22837,N_20319,N_20254);
xor U22838 (N_22838,N_20350,N_19315);
nor U22839 (N_22839,N_21638,N_20855);
and U22840 (N_22840,N_19636,N_20455);
or U22841 (N_22841,N_20148,N_21173);
or U22842 (N_22842,N_19090,N_19048);
xnor U22843 (N_22843,N_19399,N_21411);
nor U22844 (N_22844,N_20797,N_19693);
nand U22845 (N_22845,N_20407,N_20073);
xor U22846 (N_22846,N_21131,N_20764);
or U22847 (N_22847,N_19127,N_19637);
xor U22848 (N_22848,N_21832,N_18922);
nor U22849 (N_22849,N_21270,N_20016);
and U22850 (N_22850,N_20775,N_20141);
or U22851 (N_22851,N_19363,N_20766);
or U22852 (N_22852,N_18948,N_19950);
nand U22853 (N_22853,N_19709,N_20758);
or U22854 (N_22854,N_20108,N_21044);
nand U22855 (N_22855,N_20140,N_19160);
nand U22856 (N_22856,N_19909,N_21074);
and U22857 (N_22857,N_21564,N_19594);
xor U22858 (N_22858,N_21020,N_19902);
or U22859 (N_22859,N_19509,N_21095);
nand U22860 (N_22860,N_21106,N_19125);
nor U22861 (N_22861,N_20473,N_21297);
nor U22862 (N_22862,N_20988,N_19164);
nand U22863 (N_22863,N_20699,N_19308);
and U22864 (N_22864,N_21723,N_18785);
and U22865 (N_22865,N_19794,N_20348);
nand U22866 (N_22866,N_19700,N_20156);
and U22867 (N_22867,N_20642,N_21402);
or U22868 (N_22868,N_19317,N_20831);
nand U22869 (N_22869,N_19856,N_19702);
and U22870 (N_22870,N_20678,N_20489);
nor U22871 (N_22871,N_21298,N_21069);
nor U22872 (N_22872,N_19150,N_20741);
xnor U22873 (N_22873,N_20735,N_20991);
nand U22874 (N_22874,N_20501,N_21783);
xor U22875 (N_22875,N_20549,N_19557);
xor U22876 (N_22876,N_20742,N_21149);
xnor U22877 (N_22877,N_19206,N_19144);
and U22878 (N_22878,N_19971,N_21248);
nand U22879 (N_22879,N_19185,N_21435);
nor U22880 (N_22880,N_20736,N_21373);
nand U22881 (N_22881,N_21669,N_20089);
or U22882 (N_22882,N_19543,N_20712);
and U22883 (N_22883,N_21016,N_19464);
or U22884 (N_22884,N_19466,N_20779);
and U22885 (N_22885,N_21652,N_20038);
or U22886 (N_22886,N_20842,N_20806);
nand U22887 (N_22887,N_21392,N_21780);
or U22888 (N_22888,N_20972,N_21237);
nor U22889 (N_22889,N_19829,N_19495);
or U22890 (N_22890,N_19796,N_20056);
or U22891 (N_22891,N_21065,N_20115);
xor U22892 (N_22892,N_20311,N_20577);
nor U22893 (N_22893,N_19776,N_20380);
nand U22894 (N_22894,N_19604,N_21335);
or U22895 (N_22895,N_21461,N_20240);
nor U22896 (N_22896,N_21657,N_21868);
and U22897 (N_22897,N_19012,N_19259);
or U22898 (N_22898,N_19884,N_21140);
xor U22899 (N_22899,N_21463,N_21720);
xor U22900 (N_22900,N_21776,N_19108);
nor U22901 (N_22901,N_19111,N_20889);
and U22902 (N_22902,N_19975,N_19572);
xor U22903 (N_22903,N_21512,N_19800);
or U22904 (N_22904,N_21234,N_20303);
and U22905 (N_22905,N_21587,N_20880);
or U22906 (N_22906,N_21649,N_19371);
and U22907 (N_22907,N_20816,N_20584);
xnor U22908 (N_22908,N_18979,N_20079);
xor U22909 (N_22909,N_21874,N_19952);
and U22910 (N_22910,N_20607,N_21088);
or U22911 (N_22911,N_20271,N_21618);
xor U22912 (N_22912,N_20063,N_21099);
nor U22913 (N_22913,N_20383,N_20045);
nor U22914 (N_22914,N_20180,N_21604);
nor U22915 (N_22915,N_19591,N_21292);
and U22916 (N_22916,N_18927,N_21134);
nor U22917 (N_22917,N_20558,N_18786);
nand U22918 (N_22918,N_21375,N_19436);
nor U22919 (N_22919,N_20227,N_20552);
xnor U22920 (N_22920,N_20773,N_19698);
and U22921 (N_22921,N_18760,N_19082);
or U22922 (N_22922,N_20020,N_20070);
xor U22923 (N_22923,N_20757,N_21818);
and U22924 (N_22924,N_19202,N_19781);
nor U22925 (N_22925,N_19350,N_20592);
nor U22926 (N_22926,N_19465,N_18842);
nor U22927 (N_22927,N_19945,N_18819);
nand U22928 (N_22928,N_20770,N_19279);
nand U22929 (N_22929,N_21048,N_18866);
and U22930 (N_22930,N_19137,N_20820);
and U22931 (N_22931,N_18974,N_21527);
nor U22932 (N_22932,N_19689,N_21360);
nand U22933 (N_22933,N_20215,N_20249);
nor U22934 (N_22934,N_19976,N_21404);
nand U22935 (N_22935,N_21625,N_19395);
nand U22936 (N_22936,N_18991,N_19646);
and U22937 (N_22937,N_21432,N_20001);
or U22938 (N_22938,N_20403,N_20768);
and U22939 (N_22939,N_19662,N_20551);
nor U22940 (N_22940,N_21322,N_21224);
nand U22941 (N_22941,N_19923,N_20330);
nand U22942 (N_22942,N_18804,N_19606);
and U22943 (N_22943,N_21448,N_21148);
and U22944 (N_22944,N_20387,N_21107);
or U22945 (N_22945,N_19385,N_21178);
nor U22946 (N_22946,N_21717,N_20474);
nor U22947 (N_22947,N_21000,N_19145);
nor U22948 (N_22948,N_21183,N_19731);
xor U22949 (N_22949,N_20253,N_20246);
xor U22950 (N_22950,N_20721,N_21429);
nand U22951 (N_22951,N_19579,N_19848);
xor U22952 (N_22952,N_21132,N_21176);
nand U22953 (N_22953,N_21249,N_20682);
nor U22954 (N_22954,N_21636,N_19894);
nor U22955 (N_22955,N_19607,N_18902);
nand U22956 (N_22956,N_19085,N_21343);
nor U22957 (N_22957,N_19823,N_19051);
nand U22958 (N_22958,N_21261,N_19661);
nor U22959 (N_22959,N_20223,N_19138);
and U22960 (N_22960,N_19989,N_20259);
and U22961 (N_22961,N_20765,N_21415);
or U22962 (N_22962,N_19590,N_19434);
or U22963 (N_22963,N_19474,N_19375);
nor U22964 (N_22964,N_20643,N_20710);
nor U22965 (N_22965,N_20414,N_19740);
nand U22966 (N_22966,N_18835,N_19498);
nor U22967 (N_22967,N_20850,N_21586);
nor U22968 (N_22968,N_20829,N_21713);
and U22969 (N_22969,N_20008,N_19684);
xnor U22970 (N_22970,N_19845,N_20690);
and U22971 (N_22971,N_20465,N_21225);
xnor U22972 (N_22972,N_20447,N_21774);
nand U22973 (N_22973,N_21213,N_19744);
nand U22974 (N_22974,N_20726,N_21761);
xnor U22975 (N_22975,N_21264,N_21420);
and U22976 (N_22976,N_21407,N_20411);
or U22977 (N_22977,N_20460,N_19326);
xnor U22978 (N_22978,N_21503,N_20658);
or U22979 (N_22979,N_21396,N_21735);
xor U22980 (N_22980,N_19821,N_18772);
nand U22981 (N_22981,N_21380,N_19901);
nor U22982 (N_22982,N_21791,N_19457);
or U22983 (N_22983,N_21616,N_19715);
and U22984 (N_22984,N_19799,N_20103);
xnor U22985 (N_22985,N_20617,N_20027);
nand U22986 (N_22986,N_19377,N_20661);
nand U22987 (N_22987,N_21474,N_21476);
nand U22988 (N_22988,N_18962,N_21872);
nor U22989 (N_22989,N_18857,N_21240);
nand U22990 (N_22990,N_21653,N_21026);
and U22991 (N_22991,N_20430,N_19668);
or U22992 (N_22992,N_20619,N_21072);
xnor U22993 (N_22993,N_19532,N_20740);
or U22994 (N_22994,N_20588,N_21349);
and U22995 (N_22995,N_19875,N_20373);
xor U22996 (N_22996,N_21111,N_20928);
xor U22997 (N_22997,N_20219,N_20731);
xnor U22998 (N_22998,N_20503,N_21033);
xor U22999 (N_22999,N_20920,N_19314);
and U23000 (N_23000,N_18984,N_19629);
or U23001 (N_23001,N_21624,N_19711);
nand U23002 (N_23002,N_21752,N_19880);
and U23003 (N_23003,N_18891,N_20906);
nand U23004 (N_23004,N_20518,N_20851);
or U23005 (N_23005,N_19155,N_20025);
and U23006 (N_23006,N_20964,N_19788);
nor U23007 (N_23007,N_21389,N_19527);
nand U23008 (N_23008,N_19864,N_19369);
xor U23009 (N_23009,N_20527,N_19471);
or U23010 (N_23010,N_19528,N_21639);
or U23011 (N_23011,N_20310,N_19053);
or U23012 (N_23012,N_20691,N_21400);
nor U23013 (N_23013,N_19268,N_19978);
nor U23014 (N_23014,N_21569,N_21529);
and U23015 (N_23015,N_20384,N_19320);
nor U23016 (N_23016,N_21077,N_19347);
nor U23017 (N_23017,N_21617,N_20301);
nor U23018 (N_23018,N_19708,N_19367);
nand U23019 (N_23019,N_21796,N_21391);
nand U23020 (N_23020,N_19278,N_20071);
nand U23021 (N_23021,N_20981,N_21412);
xor U23022 (N_23022,N_20425,N_19213);
or U23023 (N_23023,N_20266,N_19042);
or U23024 (N_23024,N_20693,N_21023);
xnor U23025 (N_23025,N_20604,N_20897);
and U23026 (N_23026,N_20238,N_19873);
nor U23027 (N_23027,N_19381,N_19930);
and U23028 (N_23028,N_20553,N_20788);
or U23029 (N_23029,N_19106,N_21318);
nand U23030 (N_23030,N_18983,N_19906);
xor U23031 (N_23031,N_18918,N_20596);
and U23032 (N_23032,N_20650,N_19868);
and U23033 (N_23033,N_21347,N_21740);
and U23034 (N_23034,N_19057,N_21710);
and U23035 (N_23035,N_21126,N_18986);
xnor U23036 (N_23036,N_21836,N_21384);
nor U23037 (N_23037,N_19198,N_19544);
and U23038 (N_23038,N_21040,N_19886);
nand U23039 (N_23039,N_20448,N_20572);
or U23040 (N_23040,N_21390,N_19462);
nand U23041 (N_23041,N_21790,N_19370);
nor U23042 (N_23042,N_20848,N_20066);
nor U23043 (N_23043,N_21590,N_19742);
or U23044 (N_23044,N_20790,N_21469);
or U23045 (N_23045,N_19922,N_20453);
or U23046 (N_23046,N_20408,N_21635);
and U23047 (N_23047,N_20873,N_20450);
xnor U23048 (N_23048,N_20432,N_21750);
nand U23049 (N_23049,N_19289,N_19357);
or U23050 (N_23050,N_20917,N_21509);
and U23051 (N_23051,N_19807,N_20013);
xnor U23052 (N_23052,N_20767,N_20053);
or U23053 (N_23053,N_21200,N_20982);
xor U23054 (N_23054,N_21268,N_19857);
and U23055 (N_23055,N_19113,N_18768);
nand U23056 (N_23056,N_19840,N_18836);
nand U23057 (N_23057,N_20129,N_19997);
xnor U23058 (N_23058,N_21221,N_19982);
nor U23059 (N_23059,N_19650,N_21226);
or U23060 (N_23060,N_20237,N_21064);
xor U23061 (N_23061,N_20292,N_19374);
xnor U23062 (N_23062,N_18840,N_18817);
nand U23063 (N_23063,N_18960,N_21545);
xnor U23064 (N_23064,N_21232,N_18928);
and U23065 (N_23065,N_19325,N_21363);
nand U23066 (N_23066,N_21615,N_19182);
nor U23067 (N_23067,N_19430,N_19549);
nor U23068 (N_23068,N_20613,N_20713);
or U23069 (N_23069,N_19496,N_19494);
nand U23070 (N_23070,N_20285,N_19095);
nand U23071 (N_23071,N_19616,N_19881);
or U23072 (N_23072,N_21345,N_18781);
nor U23073 (N_23073,N_19785,N_19944);
nand U23074 (N_23074,N_21479,N_21325);
nand U23075 (N_23075,N_20376,N_20427);
nand U23076 (N_23076,N_19828,N_19732);
or U23077 (N_23077,N_19156,N_18757);
xnor U23078 (N_23078,N_19010,N_19725);
nor U23079 (N_23079,N_21862,N_21303);
or U23080 (N_23080,N_20211,N_20413);
and U23081 (N_23081,N_20142,N_21760);
nand U23082 (N_23082,N_21013,N_20965);
or U23083 (N_23083,N_21217,N_20730);
and U23084 (N_23084,N_21622,N_19508);
xor U23085 (N_23085,N_20859,N_20625);
and U23086 (N_23086,N_19695,N_19311);
nor U23087 (N_23087,N_20861,N_19131);
nand U23088 (N_23088,N_19859,N_19059);
nand U23089 (N_23089,N_21338,N_21754);
and U23090 (N_23090,N_20043,N_20359);
or U23091 (N_23091,N_19046,N_19763);
nor U23092 (N_23092,N_20278,N_20171);
nor U23093 (N_23093,N_19690,N_19451);
or U23094 (N_23094,N_21869,N_20838);
nor U23095 (N_23095,N_19264,N_21646);
and U23096 (N_23096,N_18950,N_19054);
nand U23097 (N_23097,N_21052,N_19348);
nand U23098 (N_23098,N_19843,N_19050);
nand U23099 (N_23099,N_20672,N_21359);
nand U23100 (N_23100,N_20136,N_21803);
nand U23101 (N_23101,N_19939,N_21654);
and U23102 (N_23102,N_20155,N_18763);
nand U23103 (N_23103,N_21606,N_21528);
or U23104 (N_23104,N_19261,N_21289);
nor U23105 (N_23105,N_20314,N_18898);
or U23106 (N_23106,N_18904,N_20329);
and U23107 (N_23107,N_21532,N_20389);
or U23108 (N_23108,N_21673,N_21517);
xor U23109 (N_23109,N_21031,N_21365);
or U23110 (N_23110,N_20578,N_20998);
and U23111 (N_23111,N_21568,N_18838);
nand U23112 (N_23112,N_18791,N_20976);
nor U23113 (N_23113,N_19497,N_19047);
and U23114 (N_23114,N_19652,N_20692);
and U23115 (N_23115,N_21706,N_21522);
nor U23116 (N_23116,N_20166,N_19664);
xnor U23117 (N_23117,N_19285,N_21194);
xnor U23118 (N_23118,N_21309,N_21011);
nand U23119 (N_23119,N_20718,N_19871);
nor U23120 (N_23120,N_19094,N_19980);
or U23121 (N_23121,N_20251,N_21207);
xnor U23122 (N_23122,N_20869,N_18793);
nand U23123 (N_23123,N_20860,N_20709);
nand U23124 (N_23124,N_19679,N_21506);
or U23125 (N_23125,N_18815,N_20019);
and U23126 (N_23126,N_20654,N_21781);
and U23127 (N_23127,N_19682,N_18811);
xor U23128 (N_23128,N_21549,N_20098);
and U23129 (N_23129,N_19470,N_19211);
xor U23130 (N_23130,N_19414,N_20058);
nor U23131 (N_23131,N_19928,N_21348);
and U23132 (N_23132,N_20929,N_19118);
or U23133 (N_23133,N_20763,N_21118);
nor U23134 (N_23134,N_20307,N_21079);
and U23135 (N_23135,N_20466,N_20995);
nor U23136 (N_23136,N_21223,N_21547);
and U23137 (N_23137,N_19001,N_20804);
and U23138 (N_23138,N_19583,N_19523);
or U23139 (N_23139,N_20229,N_18862);
or U23140 (N_23140,N_18841,N_18999);
xnor U23141 (N_23141,N_20041,N_20932);
nor U23142 (N_23142,N_20679,N_21716);
nor U23143 (N_23143,N_21269,N_21551);
xor U23144 (N_23144,N_21498,N_19458);
nand U23145 (N_23145,N_20100,N_19784);
or U23146 (N_23146,N_20452,N_20724);
and U23147 (N_23147,N_20010,N_20409);
nor U23148 (N_23148,N_20377,N_19935);
xnor U23149 (N_23149,N_19713,N_19286);
nor U23150 (N_23150,N_19705,N_18810);
nor U23151 (N_23151,N_19229,N_19582);
and U23152 (N_23152,N_18824,N_20783);
and U23153 (N_23153,N_21279,N_20023);
xnor U23154 (N_23154,N_20800,N_19953);
nand U23155 (N_23155,N_20128,N_19513);
xor U23156 (N_23156,N_21644,N_21438);
nand U23157 (N_23157,N_20866,N_20996);
xnor U23158 (N_23158,N_20220,N_19620);
and U23159 (N_23159,N_20562,N_20087);
nand U23160 (N_23160,N_19870,N_19454);
xor U23161 (N_23161,N_19913,N_19232);
or U23162 (N_23162,N_20107,N_19294);
and U23163 (N_23163,N_19524,N_20698);
and U23164 (N_23164,N_21285,N_18830);
or U23165 (N_23165,N_20144,N_19140);
nor U23166 (N_23166,N_20755,N_18959);
nor U23167 (N_23167,N_19088,N_21762);
or U23168 (N_23168,N_20335,N_18897);
and U23169 (N_23169,N_20264,N_20121);
or U23170 (N_23170,N_20404,N_21619);
xor U23171 (N_23171,N_18938,N_19328);
or U23172 (N_23172,N_21786,N_20832);
or U23173 (N_23173,N_19966,N_19535);
or U23174 (N_23174,N_19627,N_20204);
nand U23175 (N_23175,N_20464,N_19753);
and U23176 (N_23176,N_21133,N_19038);
nand U23177 (N_23177,N_19500,N_19623);
and U23178 (N_23178,N_21689,N_19176);
nor U23179 (N_23179,N_21331,N_19914);
and U23180 (N_23180,N_19963,N_19394);
nor U23181 (N_23181,N_21227,N_18890);
nand U23182 (N_23182,N_19433,N_19723);
nand U23183 (N_23183,N_21802,N_20193);
and U23184 (N_23184,N_20557,N_20994);
or U23185 (N_23185,N_21211,N_19097);
nor U23186 (N_23186,N_20201,N_21397);
or U23187 (N_23187,N_19660,N_21340);
and U23188 (N_23188,N_20263,N_19158);
nor U23189 (N_23189,N_20333,N_21381);
nand U23190 (N_23190,N_20835,N_20265);
nor U23191 (N_23191,N_19775,N_19959);
xor U23192 (N_23192,N_18839,N_21515);
xnor U23193 (N_23193,N_19574,N_21499);
xnor U23194 (N_23194,N_21462,N_21714);
nand U23195 (N_23195,N_18879,N_20862);
nand U23196 (N_23196,N_20462,N_18828);
xor U23197 (N_23197,N_19260,N_20856);
or U23198 (N_23198,N_20639,N_20530);
nand U23199 (N_23199,N_21603,N_20993);
nor U23200 (N_23200,N_21238,N_20205);
nand U23201 (N_23201,N_21105,N_20542);
and U23202 (N_23202,N_21205,N_20641);
nand U23203 (N_23203,N_20801,N_20589);
nor U23204 (N_23204,N_20381,N_19222);
and U23205 (N_23205,N_21838,N_21725);
nand U23206 (N_23206,N_20750,N_20687);
xnor U23207 (N_23207,N_21416,N_19275);
or U23208 (N_23208,N_20544,N_21665);
or U23209 (N_23209,N_21282,N_20339);
and U23210 (N_23210,N_19733,N_21386);
nand U23211 (N_23211,N_20399,N_18941);
xor U23212 (N_23212,N_21709,N_18821);
and U23213 (N_23213,N_20051,N_20097);
nand U23214 (N_23214,N_21334,N_19874);
nand U23215 (N_23215,N_20492,N_19049);
xor U23216 (N_23216,N_20541,N_20980);
nor U23217 (N_23217,N_19926,N_21691);
xor U23218 (N_23218,N_20663,N_21682);
xnor U23219 (N_23219,N_21439,N_21605);
or U23220 (N_23220,N_21633,N_18871);
nor U23221 (N_23221,N_21039,N_19898);
xnor U23222 (N_23222,N_19005,N_19418);
nand U23223 (N_23223,N_20202,N_20005);
nand U23224 (N_23224,N_19435,N_19839);
xnor U23225 (N_23225,N_19761,N_19007);
or U23226 (N_23226,N_19910,N_20973);
nor U23227 (N_23227,N_20668,N_20567);
nor U23228 (N_23228,N_20055,N_20312);
nand U23229 (N_23229,N_20091,N_20818);
and U23230 (N_23230,N_21086,N_18823);
and U23231 (N_23231,N_19003,N_21576);
and U23232 (N_23232,N_20778,N_21629);
or U23233 (N_23233,N_21621,N_19181);
nor U23234 (N_23234,N_19382,N_19817);
xor U23235 (N_23235,N_20047,N_18907);
or U23236 (N_23236,N_20046,N_20634);
nor U23237 (N_23237,N_20624,N_19999);
and U23238 (N_23238,N_19826,N_19568);
or U23239 (N_23239,N_21307,N_21351);
or U23240 (N_23240,N_19638,N_21050);
and U23241 (N_23241,N_21700,N_21749);
xnor U23242 (N_23242,N_20729,N_21090);
and U23243 (N_23243,N_19841,N_20443);
nor U23244 (N_23244,N_20120,N_19567);
or U23245 (N_23245,N_21675,N_20195);
nor U23246 (N_23246,N_19663,N_20899);
xnor U23247 (N_23247,N_21068,N_19192);
and U23248 (N_23248,N_21367,N_21323);
xnor U23249 (N_23249,N_20582,N_19490);
nor U23250 (N_23250,N_19173,N_21459);
xnor U23251 (N_23251,N_20898,N_19834);
nand U23252 (N_23252,N_19984,N_21364);
nor U23253 (N_23253,N_18971,N_20725);
xor U23254 (N_23254,N_19178,N_21147);
or U23255 (N_23255,N_20595,N_21283);
and U23256 (N_23256,N_19310,N_20702);
and U23257 (N_23257,N_18799,N_19860);
xnor U23258 (N_23258,N_20846,N_21209);
nand U23259 (N_23259,N_19409,N_18883);
nor U23260 (N_23260,N_21305,N_19163);
nor U23261 (N_23261,N_21256,N_18807);
nand U23262 (N_23262,N_19041,N_20655);
nand U23263 (N_23263,N_21494,N_18809);
or U23264 (N_23264,N_19366,N_19648);
and U23265 (N_23265,N_20497,N_21101);
nor U23266 (N_23266,N_19477,N_21736);
xor U23267 (N_23267,N_21294,N_21554);
and U23268 (N_23268,N_20918,N_19087);
or U23269 (N_23269,N_19263,N_20267);
and U23270 (N_23270,N_20948,N_19064);
nand U23271 (N_23271,N_19552,N_21032);
nor U23272 (N_23272,N_20367,N_20813);
or U23273 (N_23273,N_21447,N_19628);
and U23274 (N_23274,N_19915,N_20154);
or U23275 (N_23275,N_19988,N_20067);
nand U23276 (N_23276,N_21678,N_20865);
xnor U23277 (N_23277,N_20911,N_19411);
xnor U23278 (N_23278,N_21423,N_19305);
or U23279 (N_23279,N_20751,N_21128);
xnor U23280 (N_23280,N_20400,N_21746);
nand U23281 (N_23281,N_20954,N_19531);
and U23282 (N_23282,N_19575,N_21344);
xor U23283 (N_23283,N_21518,N_21151);
nor U23284 (N_23284,N_19741,N_21656);
or U23285 (N_23285,N_21352,N_20192);
nor U23286 (N_23286,N_21744,N_20176);
xor U23287 (N_23287,N_21228,N_20032);
and U23288 (N_23288,N_20338,N_19461);
and U23289 (N_23289,N_21098,N_19258);
or U23290 (N_23290,N_21651,N_20362);
or U23291 (N_23291,N_19153,N_20930);
nand U23292 (N_23292,N_19994,N_19441);
nor U23293 (N_23293,N_21102,N_21304);
nor U23294 (N_23294,N_20881,N_21696);
xnor U23295 (N_23295,N_20662,N_21220);
or U23296 (N_23296,N_21103,N_19541);
xor U23297 (N_23297,N_19403,N_20075);
nand U23298 (N_23298,N_20905,N_18961);
nand U23299 (N_23299,N_20535,N_21591);
xor U23300 (N_23300,N_18846,N_19767);
nand U23301 (N_23301,N_19746,N_20941);
nand U23302 (N_23302,N_19356,N_21184);
nand U23303 (N_23303,N_19729,N_20760);
and U23304 (N_23304,N_19193,N_19380);
or U23305 (N_23305,N_19443,N_19061);
or U23306 (N_23306,N_19293,N_21275);
or U23307 (N_23307,N_21770,N_19343);
or U23308 (N_23308,N_19230,N_20028);
nor U23309 (N_23309,N_21114,N_21831);
or U23310 (N_23310,N_20035,N_20086);
nor U23311 (N_23311,N_20485,N_20656);
and U23312 (N_23312,N_21010,N_18896);
nor U23313 (N_23313,N_20533,N_21457);
and U23314 (N_23314,N_19805,N_19444);
and U23315 (N_23315,N_21236,N_19237);
and U23316 (N_23316,N_19931,N_21828);
xor U23317 (N_23317,N_21317,N_21481);
and U23318 (N_23318,N_20937,N_19228);
nand U23319 (N_23319,N_20511,N_19844);
xor U23320 (N_23320,N_21811,N_20499);
nor U23321 (N_23321,N_18917,N_21727);
or U23322 (N_23322,N_20517,N_21164);
or U23323 (N_23323,N_19619,N_21281);
nor U23324 (N_23324,N_20659,N_19002);
nand U23325 (N_23325,N_20284,N_20780);
nand U23326 (N_23326,N_19940,N_21374);
xnor U23327 (N_23327,N_21157,N_19486);
or U23328 (N_23328,N_20137,N_19225);
or U23329 (N_23329,N_19547,N_20734);
and U23330 (N_23330,N_21191,N_21290);
or U23331 (N_23331,N_20630,N_19502);
nand U23332 (N_23332,N_18951,N_20421);
nand U23333 (N_23333,N_19644,N_21688);
nor U23334 (N_23334,N_19004,N_19830);
nand U23335 (N_23335,N_19062,N_20392);
and U23336 (N_23336,N_19453,N_20077);
xor U23337 (N_23337,N_21403,N_21721);
xor U23338 (N_23338,N_21059,N_20498);
and U23339 (N_23339,N_21212,N_20560);
nor U23340 (N_23340,N_18806,N_20133);
nor U23341 (N_23341,N_20545,N_21677);
nor U23342 (N_23342,N_19537,N_21819);
xnor U23343 (N_23343,N_21467,N_19030);
and U23344 (N_23344,N_20938,N_21674);
nand U23345 (N_23345,N_20182,N_20297);
nor U23346 (N_23346,N_18906,N_18916);
or U23347 (N_23347,N_19569,N_20646);
or U23348 (N_23348,N_18899,N_19152);
and U23349 (N_23349,N_20477,N_19566);
nand U23350 (N_23350,N_19020,N_20638);
and U23351 (N_23351,N_20050,N_20749);
or U23352 (N_23352,N_20472,N_21747);
nor U23353 (N_23353,N_21446,N_19518);
xor U23354 (N_23354,N_19132,N_21028);
nor U23355 (N_23355,N_20131,N_19814);
nand U23356 (N_23356,N_19148,N_19274);
and U23357 (N_23357,N_18929,N_21154);
or U23358 (N_23358,N_21519,N_18889);
xor U23359 (N_23359,N_21034,N_21830);
and U23360 (N_23360,N_21196,N_21377);
xor U23361 (N_23361,N_19031,N_20332);
nor U23362 (N_23362,N_19253,N_19573);
or U23363 (N_23363,N_20114,N_21369);
nor U23364 (N_23364,N_20616,N_20796);
xnor U23365 (N_23365,N_20083,N_20554);
or U23366 (N_23366,N_19538,N_21356);
nand U23367 (N_23367,N_21534,N_19133);
xnor U23368 (N_23368,N_20570,N_20009);
or U23369 (N_23369,N_20876,N_19171);
nor U23370 (N_23370,N_20921,N_19262);
xnor U23371 (N_23371,N_21598,N_19764);
xor U23372 (N_23372,N_21737,N_19981);
xor U23373 (N_23373,N_21405,N_19220);
nor U23374 (N_23374,N_20393,N_19625);
nand U23375 (N_23375,N_20390,N_21336);
or U23376 (N_23376,N_19905,N_19455);
xnor U23377 (N_23377,N_19822,N_20958);
nor U23378 (N_23378,N_20821,N_20669);
nand U23379 (N_23379,N_19405,N_19077);
or U23380 (N_23380,N_21313,N_18894);
or U23381 (N_23381,N_20213,N_18801);
or U23382 (N_23382,N_19469,N_19961);
and U23383 (N_23383,N_19810,N_20711);
nand U23384 (N_23384,N_19768,N_21860);
xnor U23385 (N_23385,N_20528,N_21505);
and U23386 (N_23386,N_20366,N_19515);
or U23387 (N_23387,N_19658,N_20378);
and U23388 (N_23388,N_20437,N_20919);
and U23389 (N_23389,N_20199,N_21520);
or U23390 (N_23390,N_20438,N_21301);
nor U23391 (N_23391,N_19851,N_21507);
or U23392 (N_23392,N_19852,N_19240);
or U23393 (N_23393,N_19951,N_19899);
xor U23394 (N_23394,N_20571,N_20601);
nor U23395 (N_23395,N_19157,N_19028);
and U23396 (N_23396,N_21566,N_19597);
nor U23397 (N_23397,N_18864,N_20346);
xnor U23398 (N_23398,N_20326,N_21589);
and U23399 (N_23399,N_19540,N_18884);
nor U23400 (N_23400,N_21829,N_21824);
and U23401 (N_23401,N_19576,N_20037);
and U23402 (N_23402,N_19726,N_19861);
xor U23403 (N_23403,N_21208,N_19416);
and U23404 (N_23404,N_20275,N_20975);
xnor U23405 (N_23405,N_19456,N_19439);
or U23406 (N_23406,N_19270,N_20674);
or U23407 (N_23407,N_19977,N_21705);
and U23408 (N_23408,N_19806,N_19203);
xnor U23409 (N_23409,N_20294,N_20445);
nand U23410 (N_23410,N_21414,N_20967);
xnor U23411 (N_23411,N_20287,N_20746);
xnor U23412 (N_23412,N_20291,N_21614);
nand U23413 (N_23413,N_21491,N_20651);
or U23414 (N_23414,N_19505,N_21341);
nand U23415 (N_23415,N_20531,N_20867);
nor U23416 (N_23416,N_19866,N_19408);
or U23417 (N_23417,N_20962,N_21610);
and U23418 (N_23418,N_21049,N_21455);
nor U23419 (N_23419,N_20516,N_21239);
or U23420 (N_23420,N_20344,N_20907);
and U23421 (N_23421,N_20172,N_19130);
nand U23422 (N_23422,N_19815,N_21127);
nand U23423 (N_23423,N_20705,N_19360);
xnor U23424 (N_23424,N_20719,N_19460);
nor U23425 (N_23425,N_20248,N_20222);
xor U23426 (N_23426,N_21368,N_19525);
nor U23427 (N_23427,N_19608,N_18985);
or U23428 (N_23428,N_20970,N_21759);
nor U23429 (N_23429,N_18995,N_19165);
xnor U23430 (N_23430,N_19665,N_20819);
or U23431 (N_23431,N_19447,N_19752);
or U23432 (N_23432,N_20313,N_21484);
xnor U23433 (N_23433,N_19519,N_20789);
nand U23434 (N_23434,N_20194,N_21659);
nand U23435 (N_23435,N_21458,N_21276);
xnor U23436 (N_23436,N_19244,N_19141);
xor U23437 (N_23437,N_19123,N_19858);
nand U23438 (N_23438,N_21846,N_19576);
and U23439 (N_23439,N_19702,N_21004);
nand U23440 (N_23440,N_19650,N_19607);
and U23441 (N_23441,N_20892,N_19570);
nor U23442 (N_23442,N_19189,N_19943);
nand U23443 (N_23443,N_21201,N_18889);
xor U23444 (N_23444,N_20941,N_21580);
xnor U23445 (N_23445,N_19522,N_20827);
xor U23446 (N_23446,N_20143,N_19183);
nor U23447 (N_23447,N_20356,N_19721);
and U23448 (N_23448,N_18821,N_20892);
nand U23449 (N_23449,N_21329,N_18779);
and U23450 (N_23450,N_20503,N_19113);
nor U23451 (N_23451,N_19199,N_20727);
or U23452 (N_23452,N_19738,N_20384);
or U23453 (N_23453,N_19677,N_20650);
and U23454 (N_23454,N_20156,N_21429);
nor U23455 (N_23455,N_19802,N_19373);
nor U23456 (N_23456,N_21241,N_21838);
xnor U23457 (N_23457,N_21686,N_20755);
nor U23458 (N_23458,N_20068,N_20306);
xor U23459 (N_23459,N_18776,N_18862);
and U23460 (N_23460,N_18900,N_20568);
xnor U23461 (N_23461,N_19929,N_18989);
nand U23462 (N_23462,N_19169,N_20552);
nor U23463 (N_23463,N_19270,N_19960);
nor U23464 (N_23464,N_19139,N_19576);
and U23465 (N_23465,N_19796,N_19292);
nor U23466 (N_23466,N_20923,N_20985);
nor U23467 (N_23467,N_20872,N_21230);
nand U23468 (N_23468,N_21002,N_19492);
nand U23469 (N_23469,N_20001,N_19372);
nor U23470 (N_23470,N_20491,N_21434);
or U23471 (N_23471,N_18754,N_20756);
nand U23472 (N_23472,N_20066,N_20348);
xor U23473 (N_23473,N_19678,N_19875);
and U23474 (N_23474,N_21718,N_19777);
nand U23475 (N_23475,N_21341,N_20935);
or U23476 (N_23476,N_19059,N_21154);
and U23477 (N_23477,N_18853,N_20807);
nor U23478 (N_23478,N_19199,N_21194);
or U23479 (N_23479,N_21196,N_21398);
nor U23480 (N_23480,N_21123,N_21631);
and U23481 (N_23481,N_18874,N_19843);
nand U23482 (N_23482,N_20223,N_20925);
nand U23483 (N_23483,N_19312,N_19214);
and U23484 (N_23484,N_19102,N_21658);
nand U23485 (N_23485,N_19716,N_18972);
nor U23486 (N_23486,N_19541,N_20731);
nand U23487 (N_23487,N_21622,N_20025);
or U23488 (N_23488,N_20224,N_19277);
nor U23489 (N_23489,N_21279,N_21684);
and U23490 (N_23490,N_20776,N_20831);
nor U23491 (N_23491,N_19609,N_19380);
nand U23492 (N_23492,N_20239,N_21815);
or U23493 (N_23493,N_19760,N_19148);
or U23494 (N_23494,N_21305,N_21432);
xnor U23495 (N_23495,N_19827,N_20115);
nand U23496 (N_23496,N_20778,N_19576);
and U23497 (N_23497,N_21571,N_19184);
or U23498 (N_23498,N_21018,N_20548);
xor U23499 (N_23499,N_20759,N_18932);
or U23500 (N_23500,N_19965,N_21753);
and U23501 (N_23501,N_20833,N_20127);
or U23502 (N_23502,N_19051,N_21727);
nor U23503 (N_23503,N_19830,N_21619);
xnor U23504 (N_23504,N_19378,N_21197);
xnor U23505 (N_23505,N_19959,N_21722);
or U23506 (N_23506,N_21266,N_20076);
and U23507 (N_23507,N_20609,N_19667);
and U23508 (N_23508,N_21663,N_20997);
nor U23509 (N_23509,N_21391,N_21493);
or U23510 (N_23510,N_19536,N_21587);
nor U23511 (N_23511,N_20178,N_19617);
and U23512 (N_23512,N_21417,N_21355);
xor U23513 (N_23513,N_18834,N_19330);
nor U23514 (N_23514,N_21845,N_19992);
or U23515 (N_23515,N_19479,N_20279);
nor U23516 (N_23516,N_21308,N_20098);
xnor U23517 (N_23517,N_20584,N_19823);
xor U23518 (N_23518,N_21770,N_19598);
nand U23519 (N_23519,N_21347,N_20978);
nor U23520 (N_23520,N_20822,N_19043);
nor U23521 (N_23521,N_19361,N_21491);
nand U23522 (N_23522,N_21828,N_20391);
nand U23523 (N_23523,N_20743,N_20203);
xor U23524 (N_23524,N_20644,N_20468);
and U23525 (N_23525,N_21869,N_21805);
nand U23526 (N_23526,N_20172,N_21779);
or U23527 (N_23527,N_21368,N_21620);
and U23528 (N_23528,N_19374,N_20847);
nor U23529 (N_23529,N_20587,N_19192);
nand U23530 (N_23530,N_21721,N_21341);
nor U23531 (N_23531,N_21224,N_19784);
and U23532 (N_23532,N_21521,N_21623);
nand U23533 (N_23533,N_20780,N_20290);
and U23534 (N_23534,N_19168,N_21826);
nand U23535 (N_23535,N_20400,N_20283);
and U23536 (N_23536,N_20183,N_21142);
and U23537 (N_23537,N_20332,N_19377);
nand U23538 (N_23538,N_19566,N_21295);
xnor U23539 (N_23539,N_21797,N_19836);
nor U23540 (N_23540,N_20258,N_20657);
nand U23541 (N_23541,N_18996,N_20002);
nor U23542 (N_23542,N_21332,N_20080);
or U23543 (N_23543,N_20726,N_19691);
xnor U23544 (N_23544,N_21272,N_21374);
xor U23545 (N_23545,N_19060,N_18856);
nand U23546 (N_23546,N_19070,N_21276);
or U23547 (N_23547,N_19123,N_19182);
and U23548 (N_23548,N_21193,N_19991);
nand U23549 (N_23549,N_20101,N_18891);
xnor U23550 (N_23550,N_19987,N_19194);
or U23551 (N_23551,N_20507,N_20084);
or U23552 (N_23552,N_21833,N_21094);
nand U23553 (N_23553,N_20614,N_20185);
nor U23554 (N_23554,N_21176,N_19104);
xor U23555 (N_23555,N_20083,N_19292);
and U23556 (N_23556,N_19383,N_20318);
and U23557 (N_23557,N_20245,N_19798);
and U23558 (N_23558,N_21687,N_19512);
and U23559 (N_23559,N_19593,N_21450);
or U23560 (N_23560,N_18977,N_20049);
nor U23561 (N_23561,N_21353,N_19298);
nor U23562 (N_23562,N_21123,N_20337);
and U23563 (N_23563,N_21758,N_19947);
and U23564 (N_23564,N_19031,N_18892);
xnor U23565 (N_23565,N_20567,N_19998);
xnor U23566 (N_23566,N_20446,N_20356);
or U23567 (N_23567,N_19709,N_21005);
xor U23568 (N_23568,N_20227,N_21542);
nand U23569 (N_23569,N_21414,N_21839);
and U23570 (N_23570,N_19675,N_21159);
nor U23571 (N_23571,N_19520,N_21110);
nor U23572 (N_23572,N_21771,N_19822);
and U23573 (N_23573,N_21250,N_18949);
and U23574 (N_23574,N_21751,N_19460);
xnor U23575 (N_23575,N_21219,N_19009);
nor U23576 (N_23576,N_21715,N_21771);
xnor U23577 (N_23577,N_19735,N_19754);
xor U23578 (N_23578,N_19291,N_21669);
or U23579 (N_23579,N_19415,N_20475);
nand U23580 (N_23580,N_20339,N_21805);
nand U23581 (N_23581,N_21205,N_21862);
nand U23582 (N_23582,N_21122,N_20408);
nand U23583 (N_23583,N_21155,N_21707);
and U23584 (N_23584,N_20044,N_21864);
and U23585 (N_23585,N_21739,N_20630);
or U23586 (N_23586,N_20942,N_21679);
xnor U23587 (N_23587,N_20403,N_20375);
nand U23588 (N_23588,N_18769,N_21850);
or U23589 (N_23589,N_19576,N_20087);
xnor U23590 (N_23590,N_21761,N_19603);
nand U23591 (N_23591,N_20906,N_21659);
xnor U23592 (N_23592,N_18845,N_19565);
xor U23593 (N_23593,N_19263,N_20540);
or U23594 (N_23594,N_19441,N_21180);
nor U23595 (N_23595,N_21050,N_21471);
xor U23596 (N_23596,N_19571,N_20571);
nor U23597 (N_23597,N_20963,N_20702);
and U23598 (N_23598,N_19696,N_19307);
xnor U23599 (N_23599,N_19282,N_21856);
and U23600 (N_23600,N_19227,N_19710);
nor U23601 (N_23601,N_20225,N_19328);
or U23602 (N_23602,N_19458,N_21678);
or U23603 (N_23603,N_19720,N_19977);
or U23604 (N_23604,N_21451,N_20933);
xnor U23605 (N_23605,N_19357,N_19010);
nand U23606 (N_23606,N_19352,N_21040);
nand U23607 (N_23607,N_18856,N_21373);
or U23608 (N_23608,N_19810,N_20977);
nand U23609 (N_23609,N_20558,N_21073);
nor U23610 (N_23610,N_21134,N_20365);
and U23611 (N_23611,N_19406,N_20764);
and U23612 (N_23612,N_21244,N_21279);
nor U23613 (N_23613,N_21672,N_20322);
xor U23614 (N_23614,N_21732,N_20620);
or U23615 (N_23615,N_21141,N_21229);
and U23616 (N_23616,N_19487,N_20028);
and U23617 (N_23617,N_19168,N_21392);
nand U23618 (N_23618,N_21535,N_20355);
and U23619 (N_23619,N_19775,N_19675);
nor U23620 (N_23620,N_19064,N_21166);
xor U23621 (N_23621,N_20651,N_19331);
and U23622 (N_23622,N_19378,N_19549);
and U23623 (N_23623,N_19201,N_19093);
xor U23624 (N_23624,N_19554,N_20597);
nand U23625 (N_23625,N_21104,N_21055);
nand U23626 (N_23626,N_21376,N_20949);
xor U23627 (N_23627,N_19061,N_21502);
nand U23628 (N_23628,N_20051,N_20128);
xor U23629 (N_23629,N_19806,N_18823);
nand U23630 (N_23630,N_20784,N_19319);
nand U23631 (N_23631,N_19031,N_21048);
or U23632 (N_23632,N_20402,N_19670);
nor U23633 (N_23633,N_20118,N_19332);
or U23634 (N_23634,N_21600,N_21421);
or U23635 (N_23635,N_21060,N_19993);
nor U23636 (N_23636,N_19792,N_19911);
nand U23637 (N_23637,N_19088,N_19974);
or U23638 (N_23638,N_19862,N_21306);
xnor U23639 (N_23639,N_19345,N_21117);
xnor U23640 (N_23640,N_21853,N_19275);
or U23641 (N_23641,N_19777,N_21282);
nor U23642 (N_23642,N_20873,N_19250);
xor U23643 (N_23643,N_18895,N_19919);
and U23644 (N_23644,N_20427,N_21185);
nand U23645 (N_23645,N_21163,N_20089);
or U23646 (N_23646,N_20083,N_20373);
nand U23647 (N_23647,N_21437,N_20853);
xnor U23648 (N_23648,N_20024,N_19301);
xnor U23649 (N_23649,N_21689,N_19465);
or U23650 (N_23650,N_21468,N_21113);
nand U23651 (N_23651,N_19066,N_19732);
nor U23652 (N_23652,N_21401,N_20825);
or U23653 (N_23653,N_18806,N_19597);
nand U23654 (N_23654,N_20498,N_19194);
nand U23655 (N_23655,N_18767,N_20933);
nand U23656 (N_23656,N_20814,N_19111);
nor U23657 (N_23657,N_21192,N_19589);
nor U23658 (N_23658,N_21200,N_19178);
and U23659 (N_23659,N_21677,N_19181);
xnor U23660 (N_23660,N_20007,N_21572);
or U23661 (N_23661,N_21370,N_19135);
or U23662 (N_23662,N_20899,N_20907);
xor U23663 (N_23663,N_20318,N_21385);
nand U23664 (N_23664,N_21358,N_19844);
nand U23665 (N_23665,N_19562,N_20591);
nor U23666 (N_23666,N_21693,N_21099);
or U23667 (N_23667,N_21251,N_20154);
nor U23668 (N_23668,N_20573,N_20082);
nor U23669 (N_23669,N_19162,N_21807);
nor U23670 (N_23670,N_20273,N_18995);
nand U23671 (N_23671,N_19893,N_19872);
nand U23672 (N_23672,N_20159,N_21183);
or U23673 (N_23673,N_19632,N_20401);
nand U23674 (N_23674,N_20206,N_20847);
and U23675 (N_23675,N_19776,N_19292);
xnor U23676 (N_23676,N_20404,N_20929);
nor U23677 (N_23677,N_19903,N_18933);
nand U23678 (N_23678,N_21615,N_20267);
or U23679 (N_23679,N_21573,N_19912);
xnor U23680 (N_23680,N_20806,N_18991);
and U23681 (N_23681,N_19733,N_19662);
nor U23682 (N_23682,N_20077,N_21823);
xnor U23683 (N_23683,N_19225,N_21417);
nor U23684 (N_23684,N_19978,N_20906);
or U23685 (N_23685,N_19567,N_19419);
nor U23686 (N_23686,N_19276,N_19181);
and U23687 (N_23687,N_19312,N_20334);
nor U23688 (N_23688,N_18968,N_19167);
nand U23689 (N_23689,N_21188,N_21032);
nand U23690 (N_23690,N_20468,N_19159);
nand U23691 (N_23691,N_20293,N_20140);
and U23692 (N_23692,N_21346,N_19260);
or U23693 (N_23693,N_19545,N_19185);
or U23694 (N_23694,N_20671,N_20122);
nor U23695 (N_23695,N_19240,N_18964);
nand U23696 (N_23696,N_19455,N_21814);
nor U23697 (N_23697,N_20392,N_19515);
xnor U23698 (N_23698,N_20422,N_21040);
or U23699 (N_23699,N_21237,N_18832);
nor U23700 (N_23700,N_18756,N_19700);
or U23701 (N_23701,N_21520,N_20808);
and U23702 (N_23702,N_20070,N_19634);
nand U23703 (N_23703,N_18920,N_20107);
nand U23704 (N_23704,N_18759,N_19494);
xor U23705 (N_23705,N_20007,N_19190);
xor U23706 (N_23706,N_19357,N_18852);
nand U23707 (N_23707,N_20387,N_21693);
nor U23708 (N_23708,N_19226,N_20716);
nor U23709 (N_23709,N_21871,N_20442);
nor U23710 (N_23710,N_19409,N_21649);
or U23711 (N_23711,N_21470,N_19682);
xor U23712 (N_23712,N_20825,N_19788);
nor U23713 (N_23713,N_19442,N_19389);
xor U23714 (N_23714,N_20547,N_19558);
and U23715 (N_23715,N_20754,N_21305);
xor U23716 (N_23716,N_20648,N_18873);
or U23717 (N_23717,N_21259,N_20440);
or U23718 (N_23718,N_19811,N_18851);
nor U23719 (N_23719,N_18817,N_21076);
xnor U23720 (N_23720,N_18974,N_21417);
or U23721 (N_23721,N_19853,N_21489);
nor U23722 (N_23722,N_21874,N_20935);
nand U23723 (N_23723,N_20297,N_18800);
or U23724 (N_23724,N_19740,N_18805);
xor U23725 (N_23725,N_19599,N_19263);
nand U23726 (N_23726,N_21558,N_20609);
xnor U23727 (N_23727,N_20989,N_19240);
nor U23728 (N_23728,N_20816,N_20390);
nand U23729 (N_23729,N_20689,N_18932);
or U23730 (N_23730,N_21230,N_20133);
and U23731 (N_23731,N_21535,N_20435);
nor U23732 (N_23732,N_19809,N_21239);
nor U23733 (N_23733,N_20063,N_20016);
or U23734 (N_23734,N_21566,N_21303);
or U23735 (N_23735,N_19453,N_21500);
and U23736 (N_23736,N_20451,N_21566);
nor U23737 (N_23737,N_19896,N_20657);
and U23738 (N_23738,N_20575,N_19348);
nor U23739 (N_23739,N_19713,N_20994);
or U23740 (N_23740,N_21295,N_19654);
nand U23741 (N_23741,N_20867,N_21862);
nor U23742 (N_23742,N_20660,N_19569);
xnor U23743 (N_23743,N_20224,N_19105);
and U23744 (N_23744,N_21675,N_19338);
and U23745 (N_23745,N_20461,N_21702);
nand U23746 (N_23746,N_19220,N_18954);
xor U23747 (N_23747,N_18835,N_19627);
or U23748 (N_23748,N_20226,N_20834);
or U23749 (N_23749,N_18973,N_20053);
or U23750 (N_23750,N_19956,N_20973);
xnor U23751 (N_23751,N_18832,N_19637);
nor U23752 (N_23752,N_20528,N_19373);
or U23753 (N_23753,N_20155,N_21419);
nand U23754 (N_23754,N_19408,N_21326);
nor U23755 (N_23755,N_20795,N_19842);
or U23756 (N_23756,N_21068,N_19464);
and U23757 (N_23757,N_18847,N_21162);
and U23758 (N_23758,N_21008,N_19017);
and U23759 (N_23759,N_19648,N_20281);
nand U23760 (N_23760,N_21456,N_20129);
or U23761 (N_23761,N_19880,N_19101);
nand U23762 (N_23762,N_21608,N_21102);
xor U23763 (N_23763,N_19423,N_20780);
nor U23764 (N_23764,N_19273,N_19395);
or U23765 (N_23765,N_21760,N_21821);
nor U23766 (N_23766,N_20257,N_18942);
nand U23767 (N_23767,N_20732,N_19151);
nor U23768 (N_23768,N_21153,N_18985);
nand U23769 (N_23769,N_18911,N_21322);
or U23770 (N_23770,N_21818,N_18863);
or U23771 (N_23771,N_20758,N_19235);
nand U23772 (N_23772,N_21122,N_19352);
and U23773 (N_23773,N_20374,N_20162);
or U23774 (N_23774,N_21800,N_20986);
nand U23775 (N_23775,N_19140,N_19543);
or U23776 (N_23776,N_21109,N_19069);
nor U23777 (N_23777,N_18814,N_20023);
xnor U23778 (N_23778,N_21604,N_21799);
and U23779 (N_23779,N_20407,N_19596);
xnor U23780 (N_23780,N_19730,N_20063);
nand U23781 (N_23781,N_21317,N_19823);
xnor U23782 (N_23782,N_19672,N_20812);
nor U23783 (N_23783,N_20122,N_20555);
nand U23784 (N_23784,N_19248,N_20797);
xnor U23785 (N_23785,N_21489,N_21099);
and U23786 (N_23786,N_20509,N_19707);
and U23787 (N_23787,N_21589,N_20931);
xnor U23788 (N_23788,N_19047,N_21457);
and U23789 (N_23789,N_20318,N_19892);
xor U23790 (N_23790,N_21473,N_19360);
nor U23791 (N_23791,N_19365,N_19141);
and U23792 (N_23792,N_20861,N_20966);
and U23793 (N_23793,N_21562,N_21334);
or U23794 (N_23794,N_19564,N_19814);
xor U23795 (N_23795,N_18815,N_21164);
and U23796 (N_23796,N_21731,N_18837);
nor U23797 (N_23797,N_21440,N_19651);
or U23798 (N_23798,N_20442,N_20882);
and U23799 (N_23799,N_19150,N_20461);
xnor U23800 (N_23800,N_19624,N_20810);
nand U23801 (N_23801,N_20725,N_19049);
or U23802 (N_23802,N_19185,N_19737);
nand U23803 (N_23803,N_21854,N_20437);
nand U23804 (N_23804,N_21769,N_21146);
nand U23805 (N_23805,N_19796,N_19047);
or U23806 (N_23806,N_18932,N_20964);
nand U23807 (N_23807,N_21145,N_21436);
and U23808 (N_23808,N_20369,N_20058);
nand U23809 (N_23809,N_21240,N_20973);
or U23810 (N_23810,N_21487,N_19175);
nand U23811 (N_23811,N_19558,N_20038);
nand U23812 (N_23812,N_20119,N_21450);
and U23813 (N_23813,N_21147,N_20089);
and U23814 (N_23814,N_19402,N_19009);
nand U23815 (N_23815,N_20466,N_21765);
nor U23816 (N_23816,N_21234,N_18817);
xor U23817 (N_23817,N_19184,N_19953);
and U23818 (N_23818,N_20705,N_20911);
and U23819 (N_23819,N_19399,N_19241);
nor U23820 (N_23820,N_20031,N_21873);
or U23821 (N_23821,N_21706,N_20901);
xnor U23822 (N_23822,N_21064,N_19793);
or U23823 (N_23823,N_20338,N_20329);
and U23824 (N_23824,N_21458,N_20033);
and U23825 (N_23825,N_20505,N_19242);
and U23826 (N_23826,N_20334,N_21165);
xnor U23827 (N_23827,N_21110,N_19342);
nand U23828 (N_23828,N_19160,N_21561);
nor U23829 (N_23829,N_21414,N_21318);
or U23830 (N_23830,N_21217,N_19910);
or U23831 (N_23831,N_19719,N_21432);
and U23832 (N_23832,N_21038,N_20902);
xnor U23833 (N_23833,N_21497,N_19453);
and U23834 (N_23834,N_19867,N_21716);
nand U23835 (N_23835,N_21580,N_21047);
nor U23836 (N_23836,N_19725,N_20146);
or U23837 (N_23837,N_20598,N_21361);
nor U23838 (N_23838,N_21726,N_20505);
xnor U23839 (N_23839,N_20871,N_21773);
nand U23840 (N_23840,N_19051,N_18888);
or U23841 (N_23841,N_19238,N_21350);
xor U23842 (N_23842,N_20100,N_21670);
nand U23843 (N_23843,N_20115,N_19943);
and U23844 (N_23844,N_20891,N_20970);
nand U23845 (N_23845,N_19303,N_19616);
and U23846 (N_23846,N_19191,N_19320);
and U23847 (N_23847,N_21844,N_20376);
and U23848 (N_23848,N_19859,N_20561);
nand U23849 (N_23849,N_20457,N_19545);
xor U23850 (N_23850,N_18938,N_20945);
and U23851 (N_23851,N_18860,N_21213);
and U23852 (N_23852,N_18999,N_20116);
nand U23853 (N_23853,N_19917,N_19945);
nand U23854 (N_23854,N_19183,N_21654);
xor U23855 (N_23855,N_21342,N_20800);
nand U23856 (N_23856,N_21207,N_21130);
xor U23857 (N_23857,N_19715,N_18779);
or U23858 (N_23858,N_21843,N_21648);
and U23859 (N_23859,N_19918,N_21143);
and U23860 (N_23860,N_18772,N_21464);
xnor U23861 (N_23861,N_21067,N_20694);
and U23862 (N_23862,N_19891,N_19091);
or U23863 (N_23863,N_20044,N_20556);
or U23864 (N_23864,N_20459,N_20152);
or U23865 (N_23865,N_19894,N_19439);
nand U23866 (N_23866,N_18806,N_21752);
xnor U23867 (N_23867,N_20125,N_19929);
xnor U23868 (N_23868,N_21851,N_20917);
or U23869 (N_23869,N_19652,N_20567);
nand U23870 (N_23870,N_20166,N_20605);
xor U23871 (N_23871,N_19664,N_20537);
nand U23872 (N_23872,N_19798,N_19398);
and U23873 (N_23873,N_19361,N_19160);
and U23874 (N_23874,N_19405,N_20241);
and U23875 (N_23875,N_19565,N_19904);
and U23876 (N_23876,N_21002,N_20704);
xor U23877 (N_23877,N_19948,N_18942);
nor U23878 (N_23878,N_20459,N_20656);
and U23879 (N_23879,N_21123,N_19228);
or U23880 (N_23880,N_19356,N_20229);
xor U23881 (N_23881,N_19788,N_19251);
and U23882 (N_23882,N_19800,N_21657);
and U23883 (N_23883,N_21469,N_21547);
xnor U23884 (N_23884,N_20892,N_19066);
nor U23885 (N_23885,N_21790,N_20685);
xor U23886 (N_23886,N_19480,N_21150);
xnor U23887 (N_23887,N_19856,N_20483);
and U23888 (N_23888,N_21254,N_21830);
or U23889 (N_23889,N_19324,N_21395);
or U23890 (N_23890,N_19811,N_19157);
nand U23891 (N_23891,N_18988,N_19065);
xor U23892 (N_23892,N_19661,N_20328);
or U23893 (N_23893,N_21559,N_20673);
nor U23894 (N_23894,N_21864,N_19862);
nor U23895 (N_23895,N_21848,N_20590);
nand U23896 (N_23896,N_19778,N_19710);
and U23897 (N_23897,N_21152,N_21348);
nor U23898 (N_23898,N_19713,N_20600);
xnor U23899 (N_23899,N_21238,N_21022);
xnor U23900 (N_23900,N_20830,N_20428);
nor U23901 (N_23901,N_20985,N_21035);
xnor U23902 (N_23902,N_20160,N_19813);
or U23903 (N_23903,N_20989,N_19460);
nor U23904 (N_23904,N_18765,N_18950);
xor U23905 (N_23905,N_20653,N_18824);
nor U23906 (N_23906,N_21350,N_19777);
xnor U23907 (N_23907,N_19433,N_19824);
nor U23908 (N_23908,N_19958,N_18951);
and U23909 (N_23909,N_19718,N_21230);
xor U23910 (N_23910,N_19445,N_20269);
xnor U23911 (N_23911,N_19539,N_21683);
xor U23912 (N_23912,N_19153,N_20313);
nor U23913 (N_23913,N_20413,N_20791);
nor U23914 (N_23914,N_20162,N_20151);
nor U23915 (N_23915,N_19975,N_21534);
or U23916 (N_23916,N_21377,N_20768);
nor U23917 (N_23917,N_20153,N_20504);
nand U23918 (N_23918,N_20522,N_19141);
nor U23919 (N_23919,N_19418,N_20922);
nand U23920 (N_23920,N_21287,N_21258);
nand U23921 (N_23921,N_20642,N_19237);
nor U23922 (N_23922,N_20264,N_20080);
nor U23923 (N_23923,N_20954,N_20802);
or U23924 (N_23924,N_20272,N_21120);
or U23925 (N_23925,N_20393,N_19600);
xor U23926 (N_23926,N_18817,N_20786);
or U23927 (N_23927,N_19530,N_20225);
nand U23928 (N_23928,N_21564,N_19612);
xor U23929 (N_23929,N_19272,N_19362);
xnor U23930 (N_23930,N_19212,N_21537);
nor U23931 (N_23931,N_20270,N_20636);
and U23932 (N_23932,N_21857,N_20951);
or U23933 (N_23933,N_19912,N_21668);
or U23934 (N_23934,N_21384,N_19091);
and U23935 (N_23935,N_18778,N_21416);
and U23936 (N_23936,N_19150,N_20634);
and U23937 (N_23937,N_19184,N_19083);
nand U23938 (N_23938,N_21792,N_21364);
xor U23939 (N_23939,N_19602,N_20295);
nand U23940 (N_23940,N_19957,N_20469);
nand U23941 (N_23941,N_19395,N_20852);
nand U23942 (N_23942,N_21521,N_20048);
nor U23943 (N_23943,N_18934,N_19453);
nor U23944 (N_23944,N_20956,N_21375);
and U23945 (N_23945,N_21264,N_21044);
xor U23946 (N_23946,N_21316,N_20031);
nor U23947 (N_23947,N_18976,N_21855);
and U23948 (N_23948,N_19669,N_21302);
nand U23949 (N_23949,N_19947,N_20906);
nand U23950 (N_23950,N_19056,N_20653);
and U23951 (N_23951,N_20728,N_20249);
xor U23952 (N_23952,N_19497,N_20448);
nand U23953 (N_23953,N_20257,N_20584);
or U23954 (N_23954,N_20024,N_18869);
and U23955 (N_23955,N_20380,N_21319);
or U23956 (N_23956,N_21612,N_20286);
nand U23957 (N_23957,N_19872,N_19742);
and U23958 (N_23958,N_19416,N_21717);
xnor U23959 (N_23959,N_21504,N_20340);
nor U23960 (N_23960,N_21386,N_19260);
xnor U23961 (N_23961,N_19144,N_21352);
or U23962 (N_23962,N_21662,N_21738);
and U23963 (N_23963,N_21635,N_20767);
nor U23964 (N_23964,N_19608,N_20572);
nor U23965 (N_23965,N_20526,N_20748);
nor U23966 (N_23966,N_19830,N_20757);
or U23967 (N_23967,N_19075,N_19354);
and U23968 (N_23968,N_20869,N_21639);
nand U23969 (N_23969,N_21196,N_21529);
or U23970 (N_23970,N_19101,N_20168);
and U23971 (N_23971,N_19837,N_19166);
nor U23972 (N_23972,N_21227,N_21679);
xor U23973 (N_23973,N_20595,N_21413);
and U23974 (N_23974,N_20730,N_19329);
nand U23975 (N_23975,N_21528,N_20000);
nor U23976 (N_23976,N_19321,N_18968);
and U23977 (N_23977,N_19652,N_19891);
or U23978 (N_23978,N_20512,N_19494);
or U23979 (N_23979,N_21376,N_18754);
xor U23980 (N_23980,N_19170,N_18767);
and U23981 (N_23981,N_19500,N_19830);
and U23982 (N_23982,N_19526,N_20660);
nor U23983 (N_23983,N_18863,N_20916);
nand U23984 (N_23984,N_21474,N_19427);
or U23985 (N_23985,N_21094,N_19451);
nor U23986 (N_23986,N_20989,N_20726);
nand U23987 (N_23987,N_21469,N_18759);
nand U23988 (N_23988,N_20778,N_21149);
and U23989 (N_23989,N_20585,N_21437);
or U23990 (N_23990,N_19207,N_20100);
xnor U23991 (N_23991,N_21025,N_19391);
nor U23992 (N_23992,N_20459,N_20787);
nand U23993 (N_23993,N_19774,N_21055);
or U23994 (N_23994,N_19513,N_18840);
nand U23995 (N_23995,N_20294,N_20441);
and U23996 (N_23996,N_20382,N_18954);
or U23997 (N_23997,N_21259,N_20558);
nand U23998 (N_23998,N_18857,N_21060);
nand U23999 (N_23999,N_21763,N_20383);
or U24000 (N_24000,N_20402,N_19497);
nand U24001 (N_24001,N_19078,N_18770);
nand U24002 (N_24002,N_20788,N_20801);
xor U24003 (N_24003,N_18784,N_18759);
xnor U24004 (N_24004,N_20724,N_20212);
xnor U24005 (N_24005,N_19182,N_21764);
xor U24006 (N_24006,N_19636,N_21411);
and U24007 (N_24007,N_20366,N_20465);
nor U24008 (N_24008,N_21671,N_20857);
nand U24009 (N_24009,N_20476,N_21496);
or U24010 (N_24010,N_20321,N_19259);
and U24011 (N_24011,N_19871,N_19072);
xor U24012 (N_24012,N_19041,N_21557);
and U24013 (N_24013,N_18925,N_19845);
xnor U24014 (N_24014,N_20034,N_19557);
and U24015 (N_24015,N_19343,N_20498);
nand U24016 (N_24016,N_19921,N_21018);
nor U24017 (N_24017,N_19390,N_18842);
nor U24018 (N_24018,N_21364,N_21324);
nand U24019 (N_24019,N_18953,N_20859);
nor U24020 (N_24020,N_21490,N_21145);
xnor U24021 (N_24021,N_20040,N_20469);
and U24022 (N_24022,N_19756,N_20950);
or U24023 (N_24023,N_21555,N_20897);
nor U24024 (N_24024,N_21304,N_19380);
or U24025 (N_24025,N_21383,N_21140);
or U24026 (N_24026,N_21519,N_21813);
or U24027 (N_24027,N_19721,N_21779);
and U24028 (N_24028,N_21665,N_20159);
nand U24029 (N_24029,N_21705,N_19305);
nand U24030 (N_24030,N_21102,N_19036);
xor U24031 (N_24031,N_18882,N_19890);
xnor U24032 (N_24032,N_20669,N_19426);
nand U24033 (N_24033,N_21397,N_20473);
xnor U24034 (N_24034,N_18789,N_20801);
nor U24035 (N_24035,N_20504,N_21224);
and U24036 (N_24036,N_20684,N_21034);
and U24037 (N_24037,N_21003,N_20185);
and U24038 (N_24038,N_19035,N_19031);
xor U24039 (N_24039,N_19243,N_20000);
xnor U24040 (N_24040,N_21184,N_20772);
and U24041 (N_24041,N_21693,N_21077);
nand U24042 (N_24042,N_19782,N_21026);
nor U24043 (N_24043,N_21742,N_20601);
xnor U24044 (N_24044,N_19920,N_20985);
and U24045 (N_24045,N_20049,N_20288);
nor U24046 (N_24046,N_18827,N_19128);
or U24047 (N_24047,N_20556,N_21086);
or U24048 (N_24048,N_20012,N_20882);
xnor U24049 (N_24049,N_20628,N_19596);
or U24050 (N_24050,N_18933,N_20200);
nor U24051 (N_24051,N_21568,N_19989);
nand U24052 (N_24052,N_19398,N_21374);
nor U24053 (N_24053,N_19707,N_18865);
and U24054 (N_24054,N_19131,N_19849);
nand U24055 (N_24055,N_20165,N_19152);
nand U24056 (N_24056,N_19670,N_19653);
or U24057 (N_24057,N_20137,N_21131);
nand U24058 (N_24058,N_19170,N_21660);
xor U24059 (N_24059,N_19384,N_20196);
nor U24060 (N_24060,N_19060,N_20113);
xor U24061 (N_24061,N_19103,N_20480);
and U24062 (N_24062,N_19726,N_21857);
nand U24063 (N_24063,N_19415,N_20781);
or U24064 (N_24064,N_21542,N_19531);
xor U24065 (N_24065,N_21595,N_20110);
or U24066 (N_24066,N_19791,N_20028);
nor U24067 (N_24067,N_21375,N_21728);
or U24068 (N_24068,N_19576,N_20555);
or U24069 (N_24069,N_20100,N_20238);
and U24070 (N_24070,N_20891,N_21030);
xor U24071 (N_24071,N_18995,N_20801);
nor U24072 (N_24072,N_21345,N_20603);
nor U24073 (N_24073,N_19680,N_21638);
and U24074 (N_24074,N_21670,N_19281);
or U24075 (N_24075,N_20051,N_20226);
or U24076 (N_24076,N_21512,N_20585);
or U24077 (N_24077,N_21729,N_20059);
and U24078 (N_24078,N_21812,N_19309);
and U24079 (N_24079,N_19554,N_21738);
nor U24080 (N_24080,N_19428,N_19258);
and U24081 (N_24081,N_19516,N_18809);
nand U24082 (N_24082,N_20717,N_20970);
and U24083 (N_24083,N_20325,N_21706);
and U24084 (N_24084,N_21003,N_20186);
nor U24085 (N_24085,N_20536,N_19038);
and U24086 (N_24086,N_21246,N_20515);
or U24087 (N_24087,N_19804,N_19278);
and U24088 (N_24088,N_19288,N_20647);
xnor U24089 (N_24089,N_18953,N_20020);
or U24090 (N_24090,N_21448,N_20534);
or U24091 (N_24091,N_21263,N_21467);
or U24092 (N_24092,N_19789,N_20781);
nor U24093 (N_24093,N_19835,N_20087);
nor U24094 (N_24094,N_20862,N_20869);
nand U24095 (N_24095,N_21213,N_20904);
or U24096 (N_24096,N_21002,N_19226);
or U24097 (N_24097,N_20185,N_19402);
nor U24098 (N_24098,N_21741,N_18862);
nor U24099 (N_24099,N_20299,N_20208);
nor U24100 (N_24100,N_20864,N_20234);
nor U24101 (N_24101,N_21753,N_21122);
nand U24102 (N_24102,N_19394,N_21430);
or U24103 (N_24103,N_21744,N_21065);
and U24104 (N_24104,N_20101,N_20065);
and U24105 (N_24105,N_19666,N_21831);
nor U24106 (N_24106,N_19987,N_21473);
xor U24107 (N_24107,N_19481,N_19569);
nor U24108 (N_24108,N_19245,N_19903);
xor U24109 (N_24109,N_19805,N_19561);
nand U24110 (N_24110,N_21791,N_20110);
or U24111 (N_24111,N_21545,N_20531);
nor U24112 (N_24112,N_21736,N_21318);
nor U24113 (N_24113,N_20166,N_20937);
nand U24114 (N_24114,N_21393,N_20938);
and U24115 (N_24115,N_20700,N_21325);
nand U24116 (N_24116,N_20070,N_19233);
or U24117 (N_24117,N_19517,N_20863);
or U24118 (N_24118,N_19688,N_21598);
xnor U24119 (N_24119,N_20383,N_19145);
nand U24120 (N_24120,N_19179,N_19575);
nor U24121 (N_24121,N_21711,N_20094);
nand U24122 (N_24122,N_19910,N_18946);
nand U24123 (N_24123,N_20083,N_18868);
xnor U24124 (N_24124,N_20289,N_19405);
xnor U24125 (N_24125,N_18859,N_19300);
nor U24126 (N_24126,N_20996,N_19678);
xnor U24127 (N_24127,N_21077,N_21492);
nand U24128 (N_24128,N_19111,N_20372);
and U24129 (N_24129,N_18928,N_19754);
or U24130 (N_24130,N_21376,N_19201);
and U24131 (N_24131,N_21502,N_21172);
xor U24132 (N_24132,N_20251,N_21757);
and U24133 (N_24133,N_21373,N_19237);
or U24134 (N_24134,N_20137,N_20274);
and U24135 (N_24135,N_19723,N_20254);
nand U24136 (N_24136,N_21477,N_19465);
nor U24137 (N_24137,N_21026,N_18858);
nor U24138 (N_24138,N_19077,N_19946);
nand U24139 (N_24139,N_19164,N_19925);
nand U24140 (N_24140,N_19207,N_19032);
or U24141 (N_24141,N_21692,N_20092);
xnor U24142 (N_24142,N_21666,N_20912);
and U24143 (N_24143,N_20925,N_18873);
nand U24144 (N_24144,N_18910,N_19014);
and U24145 (N_24145,N_21657,N_20150);
xor U24146 (N_24146,N_21717,N_21136);
nor U24147 (N_24147,N_21033,N_21009);
xor U24148 (N_24148,N_21853,N_19705);
and U24149 (N_24149,N_18874,N_20030);
nand U24150 (N_24150,N_20563,N_20400);
nand U24151 (N_24151,N_19706,N_19713);
nor U24152 (N_24152,N_21791,N_19518);
xnor U24153 (N_24153,N_21328,N_20128);
nor U24154 (N_24154,N_19942,N_19988);
and U24155 (N_24155,N_21433,N_20092);
nor U24156 (N_24156,N_20903,N_21060);
xor U24157 (N_24157,N_20520,N_19797);
xnor U24158 (N_24158,N_20193,N_20062);
nand U24159 (N_24159,N_20090,N_19942);
or U24160 (N_24160,N_19436,N_21161);
xor U24161 (N_24161,N_19640,N_20969);
xor U24162 (N_24162,N_21496,N_19771);
or U24163 (N_24163,N_21511,N_21669);
and U24164 (N_24164,N_21762,N_21642);
and U24165 (N_24165,N_20349,N_19650);
or U24166 (N_24166,N_21241,N_19699);
and U24167 (N_24167,N_20956,N_20169);
xor U24168 (N_24168,N_19342,N_20422);
and U24169 (N_24169,N_21537,N_20474);
and U24170 (N_24170,N_20585,N_21433);
nor U24171 (N_24171,N_20969,N_19407);
nor U24172 (N_24172,N_21484,N_20046);
nor U24173 (N_24173,N_21223,N_18821);
nand U24174 (N_24174,N_21735,N_20783);
or U24175 (N_24175,N_20240,N_20603);
nor U24176 (N_24176,N_20873,N_19361);
and U24177 (N_24177,N_19464,N_20062);
and U24178 (N_24178,N_20998,N_21380);
nor U24179 (N_24179,N_19308,N_21835);
and U24180 (N_24180,N_21643,N_19249);
nor U24181 (N_24181,N_21098,N_19918);
or U24182 (N_24182,N_20272,N_20132);
or U24183 (N_24183,N_19460,N_21134);
or U24184 (N_24184,N_20808,N_19229);
nand U24185 (N_24185,N_18757,N_19860);
and U24186 (N_24186,N_20488,N_20604);
or U24187 (N_24187,N_21763,N_19453);
and U24188 (N_24188,N_21326,N_19491);
nand U24189 (N_24189,N_20247,N_20876);
nor U24190 (N_24190,N_18928,N_18872);
and U24191 (N_24191,N_20146,N_21788);
nor U24192 (N_24192,N_20879,N_21750);
nand U24193 (N_24193,N_18834,N_20644);
nor U24194 (N_24194,N_19118,N_21204);
nand U24195 (N_24195,N_19070,N_19910);
nor U24196 (N_24196,N_21854,N_20592);
nor U24197 (N_24197,N_20253,N_19231);
xnor U24198 (N_24198,N_20135,N_21261);
nand U24199 (N_24199,N_20814,N_19100);
nand U24200 (N_24200,N_21030,N_21319);
and U24201 (N_24201,N_19886,N_20514);
or U24202 (N_24202,N_20188,N_20237);
or U24203 (N_24203,N_19114,N_18836);
xor U24204 (N_24204,N_20769,N_20956);
nand U24205 (N_24205,N_21652,N_19941);
xnor U24206 (N_24206,N_21647,N_19619);
nand U24207 (N_24207,N_18764,N_21024);
xnor U24208 (N_24208,N_21423,N_19787);
xnor U24209 (N_24209,N_20786,N_20213);
or U24210 (N_24210,N_19174,N_20459);
or U24211 (N_24211,N_19211,N_21639);
nor U24212 (N_24212,N_19440,N_21013);
and U24213 (N_24213,N_20243,N_20767);
or U24214 (N_24214,N_19898,N_19260);
nand U24215 (N_24215,N_18758,N_21375);
nand U24216 (N_24216,N_20046,N_20404);
xnor U24217 (N_24217,N_21173,N_20083);
nand U24218 (N_24218,N_21469,N_19920);
nor U24219 (N_24219,N_21557,N_18812);
nor U24220 (N_24220,N_19424,N_20687);
nand U24221 (N_24221,N_20687,N_20770);
xor U24222 (N_24222,N_19841,N_21598);
nor U24223 (N_24223,N_19797,N_20969);
nand U24224 (N_24224,N_19774,N_20032);
nand U24225 (N_24225,N_19524,N_21535);
or U24226 (N_24226,N_18947,N_21849);
or U24227 (N_24227,N_20849,N_20734);
nor U24228 (N_24228,N_19532,N_21479);
xor U24229 (N_24229,N_20704,N_20305);
and U24230 (N_24230,N_20920,N_20786);
nor U24231 (N_24231,N_21736,N_21032);
and U24232 (N_24232,N_19214,N_20964);
xor U24233 (N_24233,N_21025,N_18770);
nor U24234 (N_24234,N_19892,N_19025);
or U24235 (N_24235,N_21761,N_20230);
nor U24236 (N_24236,N_18769,N_20443);
and U24237 (N_24237,N_20370,N_20418);
and U24238 (N_24238,N_19188,N_20315);
or U24239 (N_24239,N_21206,N_21514);
or U24240 (N_24240,N_19833,N_20473);
nand U24241 (N_24241,N_20446,N_20088);
nand U24242 (N_24242,N_21214,N_20686);
xnor U24243 (N_24243,N_20086,N_21627);
xnor U24244 (N_24244,N_21845,N_20027);
and U24245 (N_24245,N_19225,N_20344);
xnor U24246 (N_24246,N_19238,N_21328);
nor U24247 (N_24247,N_18904,N_18775);
xor U24248 (N_24248,N_20746,N_18877);
nand U24249 (N_24249,N_20812,N_19812);
and U24250 (N_24250,N_20848,N_19338);
nor U24251 (N_24251,N_20975,N_20698);
and U24252 (N_24252,N_18972,N_20980);
or U24253 (N_24253,N_19846,N_19971);
or U24254 (N_24254,N_20019,N_20969);
or U24255 (N_24255,N_19218,N_20120);
nand U24256 (N_24256,N_21355,N_21062);
nand U24257 (N_24257,N_19435,N_21670);
and U24258 (N_24258,N_21716,N_20771);
nand U24259 (N_24259,N_20286,N_21166);
nor U24260 (N_24260,N_20477,N_20940);
or U24261 (N_24261,N_20134,N_19003);
and U24262 (N_24262,N_21418,N_19654);
xor U24263 (N_24263,N_21720,N_18997);
nand U24264 (N_24264,N_19034,N_21219);
xor U24265 (N_24265,N_21395,N_21262);
or U24266 (N_24266,N_19474,N_19217);
nand U24267 (N_24267,N_18966,N_21170);
xnor U24268 (N_24268,N_20648,N_20008);
or U24269 (N_24269,N_21412,N_19711);
nand U24270 (N_24270,N_21679,N_20641);
xnor U24271 (N_24271,N_18916,N_20438);
nand U24272 (N_24272,N_21794,N_21350);
nand U24273 (N_24273,N_20971,N_21096);
nor U24274 (N_24274,N_20499,N_19027);
xor U24275 (N_24275,N_18820,N_20600);
nand U24276 (N_24276,N_20078,N_19452);
nand U24277 (N_24277,N_20866,N_19013);
and U24278 (N_24278,N_20821,N_19518);
nand U24279 (N_24279,N_19863,N_21434);
nor U24280 (N_24280,N_18870,N_20020);
and U24281 (N_24281,N_19262,N_20704);
xnor U24282 (N_24282,N_19712,N_18799);
or U24283 (N_24283,N_19833,N_19301);
nand U24284 (N_24284,N_19077,N_20517);
nor U24285 (N_24285,N_19404,N_21023);
or U24286 (N_24286,N_19303,N_19001);
nor U24287 (N_24287,N_19567,N_19885);
xnor U24288 (N_24288,N_18901,N_20405);
nor U24289 (N_24289,N_21392,N_21480);
xor U24290 (N_24290,N_20286,N_19530);
xnor U24291 (N_24291,N_18778,N_21391);
nand U24292 (N_24292,N_20350,N_19114);
nor U24293 (N_24293,N_21023,N_18893);
and U24294 (N_24294,N_18794,N_21700);
or U24295 (N_24295,N_21330,N_19130);
nor U24296 (N_24296,N_20964,N_19129);
nand U24297 (N_24297,N_19444,N_19641);
or U24298 (N_24298,N_19377,N_18808);
nor U24299 (N_24299,N_19683,N_20694);
nand U24300 (N_24300,N_19953,N_20011);
nand U24301 (N_24301,N_19514,N_18964);
or U24302 (N_24302,N_20470,N_18984);
or U24303 (N_24303,N_20467,N_19263);
or U24304 (N_24304,N_21130,N_20950);
nor U24305 (N_24305,N_19943,N_21037);
nand U24306 (N_24306,N_21428,N_21408);
nand U24307 (N_24307,N_19378,N_20417);
xnor U24308 (N_24308,N_21097,N_19624);
nand U24309 (N_24309,N_19226,N_19040);
or U24310 (N_24310,N_21605,N_18790);
nor U24311 (N_24311,N_21467,N_21106);
and U24312 (N_24312,N_20094,N_21031);
nor U24313 (N_24313,N_21713,N_20786);
or U24314 (N_24314,N_21626,N_21057);
nand U24315 (N_24315,N_19599,N_21291);
and U24316 (N_24316,N_21236,N_21660);
nor U24317 (N_24317,N_20088,N_20511);
and U24318 (N_24318,N_20764,N_20391);
and U24319 (N_24319,N_20487,N_21481);
xor U24320 (N_24320,N_19004,N_20747);
nand U24321 (N_24321,N_21444,N_19864);
xnor U24322 (N_24322,N_21671,N_19045);
or U24323 (N_24323,N_19502,N_19840);
or U24324 (N_24324,N_19829,N_19221);
nand U24325 (N_24325,N_21157,N_21154);
and U24326 (N_24326,N_20301,N_20204);
xnor U24327 (N_24327,N_20011,N_20712);
and U24328 (N_24328,N_18845,N_19066);
and U24329 (N_24329,N_21045,N_19701);
nor U24330 (N_24330,N_21766,N_20339);
and U24331 (N_24331,N_18998,N_20257);
nor U24332 (N_24332,N_20700,N_18976);
xor U24333 (N_24333,N_18932,N_20295);
nand U24334 (N_24334,N_20453,N_19822);
xnor U24335 (N_24335,N_21720,N_20888);
and U24336 (N_24336,N_21110,N_20081);
or U24337 (N_24337,N_20805,N_21104);
or U24338 (N_24338,N_19057,N_18881);
and U24339 (N_24339,N_19610,N_20975);
nand U24340 (N_24340,N_19149,N_21125);
nand U24341 (N_24341,N_19020,N_20379);
and U24342 (N_24342,N_21429,N_19317);
xor U24343 (N_24343,N_21181,N_20473);
nand U24344 (N_24344,N_21791,N_19755);
and U24345 (N_24345,N_20252,N_21281);
or U24346 (N_24346,N_19002,N_19104);
xor U24347 (N_24347,N_19810,N_19581);
nor U24348 (N_24348,N_21227,N_20319);
and U24349 (N_24349,N_21303,N_21214);
or U24350 (N_24350,N_20752,N_19546);
nor U24351 (N_24351,N_20950,N_20273);
nor U24352 (N_24352,N_19559,N_19558);
and U24353 (N_24353,N_19412,N_21121);
and U24354 (N_24354,N_19150,N_19256);
and U24355 (N_24355,N_20058,N_20913);
and U24356 (N_24356,N_19891,N_21286);
xor U24357 (N_24357,N_20091,N_20369);
or U24358 (N_24358,N_19123,N_19185);
xor U24359 (N_24359,N_19933,N_21183);
nor U24360 (N_24360,N_20594,N_19656);
or U24361 (N_24361,N_19208,N_21095);
and U24362 (N_24362,N_19613,N_20469);
nand U24363 (N_24363,N_19413,N_21867);
and U24364 (N_24364,N_21858,N_21111);
xnor U24365 (N_24365,N_21256,N_20586);
nor U24366 (N_24366,N_21874,N_19334);
xor U24367 (N_24367,N_20005,N_19712);
nor U24368 (N_24368,N_18757,N_19275);
xor U24369 (N_24369,N_19134,N_21029);
nand U24370 (N_24370,N_21076,N_20889);
and U24371 (N_24371,N_20254,N_21104);
nand U24372 (N_24372,N_21408,N_19531);
nand U24373 (N_24373,N_21056,N_19188);
nand U24374 (N_24374,N_18776,N_21232);
nand U24375 (N_24375,N_19801,N_21864);
nor U24376 (N_24376,N_18766,N_18948);
xnor U24377 (N_24377,N_19585,N_19922);
nor U24378 (N_24378,N_18775,N_21700);
and U24379 (N_24379,N_21672,N_19508);
or U24380 (N_24380,N_21566,N_19714);
nor U24381 (N_24381,N_21520,N_19450);
nand U24382 (N_24382,N_21828,N_21468);
or U24383 (N_24383,N_19399,N_20601);
xor U24384 (N_24384,N_20240,N_21517);
nor U24385 (N_24385,N_18978,N_19600);
nor U24386 (N_24386,N_19416,N_20438);
xor U24387 (N_24387,N_20054,N_19143);
nor U24388 (N_24388,N_20472,N_21358);
or U24389 (N_24389,N_20809,N_19360);
xnor U24390 (N_24390,N_18769,N_20629);
or U24391 (N_24391,N_21732,N_19278);
nor U24392 (N_24392,N_19816,N_19516);
nand U24393 (N_24393,N_19697,N_19758);
or U24394 (N_24394,N_21259,N_19683);
nand U24395 (N_24395,N_20204,N_21695);
nor U24396 (N_24396,N_21312,N_20138);
nor U24397 (N_24397,N_21617,N_21280);
nor U24398 (N_24398,N_19553,N_19760);
or U24399 (N_24399,N_19681,N_19820);
nor U24400 (N_24400,N_20051,N_20922);
or U24401 (N_24401,N_19598,N_21375);
and U24402 (N_24402,N_19241,N_19303);
xnor U24403 (N_24403,N_20712,N_20279);
and U24404 (N_24404,N_21763,N_18802);
or U24405 (N_24405,N_20673,N_21314);
xnor U24406 (N_24406,N_21854,N_21584);
nand U24407 (N_24407,N_21789,N_20126);
or U24408 (N_24408,N_20774,N_20296);
nand U24409 (N_24409,N_19448,N_20287);
nand U24410 (N_24410,N_19401,N_19175);
xor U24411 (N_24411,N_21198,N_19528);
nand U24412 (N_24412,N_19297,N_20889);
nor U24413 (N_24413,N_19443,N_21300);
and U24414 (N_24414,N_20113,N_21852);
xor U24415 (N_24415,N_18772,N_19658);
or U24416 (N_24416,N_21112,N_19215);
and U24417 (N_24417,N_20384,N_19908);
nand U24418 (N_24418,N_20134,N_21375);
or U24419 (N_24419,N_18920,N_20177);
nand U24420 (N_24420,N_19783,N_20721);
nand U24421 (N_24421,N_20521,N_20794);
or U24422 (N_24422,N_19168,N_20643);
nor U24423 (N_24423,N_20862,N_21136);
nand U24424 (N_24424,N_20812,N_20606);
nand U24425 (N_24425,N_20093,N_20090);
and U24426 (N_24426,N_19091,N_21157);
nand U24427 (N_24427,N_19586,N_18884);
nor U24428 (N_24428,N_19099,N_20862);
nor U24429 (N_24429,N_20583,N_21851);
nand U24430 (N_24430,N_20312,N_21821);
or U24431 (N_24431,N_21822,N_21444);
xnor U24432 (N_24432,N_20898,N_19767);
nand U24433 (N_24433,N_19874,N_20927);
nor U24434 (N_24434,N_20766,N_18854);
nor U24435 (N_24435,N_18885,N_19815);
or U24436 (N_24436,N_21410,N_19318);
or U24437 (N_24437,N_19704,N_20765);
xor U24438 (N_24438,N_19850,N_20840);
or U24439 (N_24439,N_20484,N_19826);
xnor U24440 (N_24440,N_21561,N_19672);
xor U24441 (N_24441,N_19559,N_20336);
and U24442 (N_24442,N_20081,N_19947);
nor U24443 (N_24443,N_18808,N_18758);
nor U24444 (N_24444,N_19552,N_19820);
nand U24445 (N_24445,N_21786,N_20716);
nand U24446 (N_24446,N_20236,N_21257);
and U24447 (N_24447,N_19129,N_19597);
nor U24448 (N_24448,N_20027,N_18872);
nand U24449 (N_24449,N_19078,N_20917);
and U24450 (N_24450,N_18955,N_20915);
or U24451 (N_24451,N_18952,N_19350);
nand U24452 (N_24452,N_20172,N_20178);
nor U24453 (N_24453,N_20143,N_20442);
nor U24454 (N_24454,N_19332,N_20195);
nor U24455 (N_24455,N_19001,N_21514);
and U24456 (N_24456,N_21449,N_21551);
and U24457 (N_24457,N_21493,N_21316);
nand U24458 (N_24458,N_19669,N_21488);
nand U24459 (N_24459,N_20786,N_20870);
nor U24460 (N_24460,N_21348,N_18907);
nor U24461 (N_24461,N_19688,N_20004);
nor U24462 (N_24462,N_20857,N_19934);
or U24463 (N_24463,N_18901,N_20948);
nand U24464 (N_24464,N_20566,N_20422);
and U24465 (N_24465,N_20815,N_19503);
and U24466 (N_24466,N_21077,N_20994);
nor U24467 (N_24467,N_21166,N_21640);
and U24468 (N_24468,N_19214,N_20983);
nand U24469 (N_24469,N_21092,N_20558);
nand U24470 (N_24470,N_21617,N_19002);
nor U24471 (N_24471,N_19585,N_21170);
nand U24472 (N_24472,N_21051,N_19970);
and U24473 (N_24473,N_19887,N_19679);
and U24474 (N_24474,N_19498,N_21534);
nor U24475 (N_24475,N_20321,N_18790);
or U24476 (N_24476,N_20440,N_21419);
and U24477 (N_24477,N_19206,N_21205);
and U24478 (N_24478,N_21497,N_19725);
nor U24479 (N_24479,N_20310,N_20320);
xor U24480 (N_24480,N_21314,N_20425);
xnor U24481 (N_24481,N_19560,N_18874);
xnor U24482 (N_24482,N_19420,N_20080);
nand U24483 (N_24483,N_21000,N_19294);
nand U24484 (N_24484,N_21417,N_20018);
or U24485 (N_24485,N_20570,N_20815);
nand U24486 (N_24486,N_20310,N_18999);
or U24487 (N_24487,N_21777,N_21458);
nand U24488 (N_24488,N_20659,N_20374);
and U24489 (N_24489,N_19647,N_20372);
nor U24490 (N_24490,N_18832,N_19301);
nand U24491 (N_24491,N_21850,N_20348);
nand U24492 (N_24492,N_21547,N_21655);
nand U24493 (N_24493,N_21551,N_21103);
or U24494 (N_24494,N_21380,N_20843);
or U24495 (N_24495,N_19891,N_20013);
or U24496 (N_24496,N_21679,N_21492);
or U24497 (N_24497,N_19666,N_19322);
and U24498 (N_24498,N_21639,N_18774);
and U24499 (N_24499,N_19564,N_21596);
xnor U24500 (N_24500,N_19440,N_20082);
or U24501 (N_24501,N_20556,N_19896);
xnor U24502 (N_24502,N_20714,N_20926);
xnor U24503 (N_24503,N_21698,N_19331);
and U24504 (N_24504,N_19468,N_18914);
nand U24505 (N_24505,N_20481,N_18845);
nand U24506 (N_24506,N_19899,N_20071);
or U24507 (N_24507,N_20285,N_20048);
or U24508 (N_24508,N_20212,N_19375);
or U24509 (N_24509,N_21221,N_19610);
and U24510 (N_24510,N_19233,N_19086);
or U24511 (N_24511,N_21190,N_19144);
or U24512 (N_24512,N_19780,N_20071);
nor U24513 (N_24513,N_19118,N_19817);
nand U24514 (N_24514,N_21220,N_18923);
nor U24515 (N_24515,N_19930,N_20565);
xor U24516 (N_24516,N_20313,N_20631);
nand U24517 (N_24517,N_20521,N_21002);
nor U24518 (N_24518,N_19848,N_18764);
nand U24519 (N_24519,N_21692,N_19821);
or U24520 (N_24520,N_21217,N_20967);
xnor U24521 (N_24521,N_20497,N_21597);
nor U24522 (N_24522,N_21267,N_21443);
and U24523 (N_24523,N_20049,N_20574);
or U24524 (N_24524,N_20109,N_18900);
and U24525 (N_24525,N_21055,N_19917);
and U24526 (N_24526,N_20170,N_21671);
xor U24527 (N_24527,N_20955,N_19521);
and U24528 (N_24528,N_20329,N_20612);
nand U24529 (N_24529,N_21000,N_20823);
or U24530 (N_24530,N_20154,N_20902);
nor U24531 (N_24531,N_21160,N_19545);
and U24532 (N_24532,N_20193,N_20977);
xnor U24533 (N_24533,N_19018,N_21008);
or U24534 (N_24534,N_21449,N_19382);
xnor U24535 (N_24535,N_20306,N_18915);
and U24536 (N_24536,N_21418,N_19986);
or U24537 (N_24537,N_21733,N_20346);
nand U24538 (N_24538,N_19863,N_20004);
and U24539 (N_24539,N_19965,N_19999);
nor U24540 (N_24540,N_20131,N_21201);
and U24541 (N_24541,N_20295,N_18926);
nor U24542 (N_24542,N_18817,N_20584);
xor U24543 (N_24543,N_21136,N_20222);
xor U24544 (N_24544,N_19676,N_21675);
or U24545 (N_24545,N_20703,N_21364);
and U24546 (N_24546,N_19851,N_19795);
xnor U24547 (N_24547,N_20490,N_19932);
nor U24548 (N_24548,N_21688,N_19549);
nand U24549 (N_24549,N_19093,N_19965);
nor U24550 (N_24550,N_20121,N_19721);
xnor U24551 (N_24551,N_21621,N_21161);
xor U24552 (N_24552,N_19295,N_19310);
nor U24553 (N_24553,N_21623,N_20541);
nor U24554 (N_24554,N_21516,N_19416);
or U24555 (N_24555,N_20728,N_21629);
nand U24556 (N_24556,N_18807,N_20389);
nand U24557 (N_24557,N_20328,N_18981);
nand U24558 (N_24558,N_18882,N_21067);
nor U24559 (N_24559,N_18958,N_21344);
nand U24560 (N_24560,N_20674,N_20416);
nor U24561 (N_24561,N_20648,N_19077);
nor U24562 (N_24562,N_20064,N_20054);
or U24563 (N_24563,N_21813,N_20094);
nor U24564 (N_24564,N_21570,N_21022);
nand U24565 (N_24565,N_19543,N_18955);
nand U24566 (N_24566,N_20070,N_20713);
xor U24567 (N_24567,N_20934,N_20012);
xor U24568 (N_24568,N_21706,N_21011);
xor U24569 (N_24569,N_18869,N_19438);
and U24570 (N_24570,N_21142,N_20301);
xor U24571 (N_24571,N_21038,N_21629);
nand U24572 (N_24572,N_21805,N_21679);
nand U24573 (N_24573,N_19799,N_19248);
or U24574 (N_24574,N_19070,N_21551);
xor U24575 (N_24575,N_20033,N_19571);
xnor U24576 (N_24576,N_21288,N_19220);
nand U24577 (N_24577,N_18909,N_20010);
xnor U24578 (N_24578,N_19509,N_21544);
xnor U24579 (N_24579,N_20385,N_20640);
and U24580 (N_24580,N_21671,N_19576);
nand U24581 (N_24581,N_21352,N_21698);
and U24582 (N_24582,N_20893,N_18865);
or U24583 (N_24583,N_21784,N_19361);
or U24584 (N_24584,N_21096,N_20069);
nand U24585 (N_24585,N_18980,N_21642);
nor U24586 (N_24586,N_21644,N_21557);
nor U24587 (N_24587,N_21516,N_19364);
nor U24588 (N_24588,N_20322,N_21592);
xnor U24589 (N_24589,N_19552,N_21874);
nor U24590 (N_24590,N_20391,N_19773);
or U24591 (N_24591,N_20013,N_20522);
nor U24592 (N_24592,N_19217,N_20791);
xnor U24593 (N_24593,N_19824,N_19345);
nand U24594 (N_24594,N_21199,N_20188);
or U24595 (N_24595,N_19791,N_19869);
xor U24596 (N_24596,N_19662,N_20930);
xor U24597 (N_24597,N_21148,N_19506);
xor U24598 (N_24598,N_19260,N_20560);
and U24599 (N_24599,N_21820,N_20778);
xor U24600 (N_24600,N_21705,N_19390);
nor U24601 (N_24601,N_19448,N_20748);
or U24602 (N_24602,N_19247,N_18998);
or U24603 (N_24603,N_20648,N_19272);
or U24604 (N_24604,N_20269,N_19643);
xnor U24605 (N_24605,N_21434,N_21654);
or U24606 (N_24606,N_20607,N_19302);
and U24607 (N_24607,N_20106,N_20428);
or U24608 (N_24608,N_19439,N_19294);
nand U24609 (N_24609,N_19907,N_19072);
nor U24610 (N_24610,N_19501,N_19437);
or U24611 (N_24611,N_21661,N_20460);
nand U24612 (N_24612,N_20113,N_21371);
or U24613 (N_24613,N_20493,N_21112);
or U24614 (N_24614,N_20886,N_21246);
xnor U24615 (N_24615,N_18838,N_21141);
xnor U24616 (N_24616,N_21430,N_19461);
nor U24617 (N_24617,N_19245,N_19969);
and U24618 (N_24618,N_19847,N_21718);
nor U24619 (N_24619,N_20963,N_21625);
and U24620 (N_24620,N_20951,N_19240);
nand U24621 (N_24621,N_20086,N_21260);
nand U24622 (N_24622,N_19674,N_20099);
and U24623 (N_24623,N_21375,N_18765);
and U24624 (N_24624,N_19987,N_21303);
or U24625 (N_24625,N_20642,N_18972);
xor U24626 (N_24626,N_21302,N_19367);
xnor U24627 (N_24627,N_18945,N_21251);
nor U24628 (N_24628,N_19328,N_19565);
xor U24629 (N_24629,N_19095,N_19625);
nor U24630 (N_24630,N_21111,N_19887);
nor U24631 (N_24631,N_19026,N_21608);
nor U24632 (N_24632,N_18964,N_20459);
nand U24633 (N_24633,N_20166,N_21332);
nand U24634 (N_24634,N_19580,N_18771);
nand U24635 (N_24635,N_20179,N_20864);
xor U24636 (N_24636,N_20590,N_21268);
xnor U24637 (N_24637,N_20285,N_21297);
and U24638 (N_24638,N_19428,N_21873);
xor U24639 (N_24639,N_20064,N_21563);
xnor U24640 (N_24640,N_19451,N_20148);
xnor U24641 (N_24641,N_20504,N_21617);
and U24642 (N_24642,N_20099,N_20822);
and U24643 (N_24643,N_21741,N_19597);
nand U24644 (N_24644,N_20765,N_21295);
and U24645 (N_24645,N_20339,N_21679);
and U24646 (N_24646,N_18915,N_19606);
nor U24647 (N_24647,N_21641,N_19103);
nor U24648 (N_24648,N_19176,N_18902);
nand U24649 (N_24649,N_20710,N_20632);
nand U24650 (N_24650,N_20025,N_20158);
or U24651 (N_24651,N_19260,N_20840);
nor U24652 (N_24652,N_20042,N_19860);
and U24653 (N_24653,N_20241,N_21462);
xnor U24654 (N_24654,N_20141,N_19109);
or U24655 (N_24655,N_19193,N_21042);
and U24656 (N_24656,N_21544,N_21594);
and U24657 (N_24657,N_21088,N_21166);
or U24658 (N_24658,N_21299,N_21319);
xor U24659 (N_24659,N_19577,N_20240);
xor U24660 (N_24660,N_21156,N_21838);
or U24661 (N_24661,N_20603,N_19232);
xor U24662 (N_24662,N_21206,N_20291);
or U24663 (N_24663,N_20513,N_19158);
and U24664 (N_24664,N_19704,N_20994);
or U24665 (N_24665,N_19432,N_19567);
nand U24666 (N_24666,N_21354,N_20339);
nand U24667 (N_24667,N_21328,N_19902);
nor U24668 (N_24668,N_20866,N_20635);
or U24669 (N_24669,N_19520,N_19876);
or U24670 (N_24670,N_20473,N_19680);
and U24671 (N_24671,N_21060,N_20532);
or U24672 (N_24672,N_18828,N_19391);
or U24673 (N_24673,N_19444,N_19820);
nand U24674 (N_24674,N_20805,N_21385);
nor U24675 (N_24675,N_19147,N_19713);
nand U24676 (N_24676,N_20210,N_19407);
and U24677 (N_24677,N_18841,N_20298);
and U24678 (N_24678,N_21171,N_20011);
nor U24679 (N_24679,N_20246,N_18874);
nor U24680 (N_24680,N_20249,N_19168);
nand U24681 (N_24681,N_19714,N_18829);
and U24682 (N_24682,N_18879,N_20050);
nor U24683 (N_24683,N_19743,N_21035);
and U24684 (N_24684,N_21288,N_20427);
xnor U24685 (N_24685,N_20533,N_18908);
nor U24686 (N_24686,N_20647,N_19243);
or U24687 (N_24687,N_20121,N_20713);
nor U24688 (N_24688,N_21003,N_19549);
nor U24689 (N_24689,N_20424,N_19757);
nor U24690 (N_24690,N_21256,N_20481);
and U24691 (N_24691,N_21233,N_19147);
nand U24692 (N_24692,N_21607,N_19180);
and U24693 (N_24693,N_20465,N_19652);
nand U24694 (N_24694,N_18933,N_19601);
and U24695 (N_24695,N_19060,N_19765);
xnor U24696 (N_24696,N_20620,N_19187);
nor U24697 (N_24697,N_21332,N_20251);
nand U24698 (N_24698,N_19953,N_21549);
nand U24699 (N_24699,N_19948,N_21114);
nor U24700 (N_24700,N_20900,N_18946);
nor U24701 (N_24701,N_20115,N_19763);
and U24702 (N_24702,N_20547,N_21716);
xor U24703 (N_24703,N_21823,N_21471);
nor U24704 (N_24704,N_21053,N_20261);
nor U24705 (N_24705,N_18831,N_19209);
or U24706 (N_24706,N_20389,N_20709);
nand U24707 (N_24707,N_18804,N_20098);
and U24708 (N_24708,N_20693,N_20875);
and U24709 (N_24709,N_20526,N_21397);
nand U24710 (N_24710,N_19603,N_19986);
or U24711 (N_24711,N_19704,N_20275);
xor U24712 (N_24712,N_21648,N_20389);
nor U24713 (N_24713,N_20164,N_21350);
or U24714 (N_24714,N_19165,N_21658);
nand U24715 (N_24715,N_21651,N_20735);
and U24716 (N_24716,N_19695,N_21619);
and U24717 (N_24717,N_20479,N_18902);
nand U24718 (N_24718,N_19322,N_20478);
and U24719 (N_24719,N_20365,N_19683);
and U24720 (N_24720,N_20029,N_18898);
and U24721 (N_24721,N_18875,N_20972);
xor U24722 (N_24722,N_19025,N_20580);
and U24723 (N_24723,N_21706,N_21580);
and U24724 (N_24724,N_19842,N_19246);
nor U24725 (N_24725,N_21271,N_19759);
nor U24726 (N_24726,N_19862,N_21200);
and U24727 (N_24727,N_21579,N_21422);
or U24728 (N_24728,N_20728,N_20081);
and U24729 (N_24729,N_21401,N_20839);
nand U24730 (N_24730,N_20855,N_19754);
nor U24731 (N_24731,N_21137,N_21163);
xor U24732 (N_24732,N_21038,N_20036);
xor U24733 (N_24733,N_20430,N_20207);
or U24734 (N_24734,N_19723,N_19117);
or U24735 (N_24735,N_21350,N_19892);
or U24736 (N_24736,N_21430,N_21023);
xor U24737 (N_24737,N_18955,N_20265);
nor U24738 (N_24738,N_19401,N_20618);
and U24739 (N_24739,N_18972,N_21174);
or U24740 (N_24740,N_21867,N_21536);
nand U24741 (N_24741,N_20744,N_19471);
and U24742 (N_24742,N_19576,N_19254);
nor U24743 (N_24743,N_18876,N_19314);
nor U24744 (N_24744,N_18853,N_21011);
or U24745 (N_24745,N_20324,N_20364);
and U24746 (N_24746,N_20761,N_21352);
xnor U24747 (N_24747,N_19544,N_19271);
nand U24748 (N_24748,N_20381,N_21219);
nand U24749 (N_24749,N_19723,N_20002);
nor U24750 (N_24750,N_18784,N_20693);
and U24751 (N_24751,N_21846,N_20755);
nand U24752 (N_24752,N_20562,N_20010);
nand U24753 (N_24753,N_20261,N_19026);
nor U24754 (N_24754,N_19557,N_19399);
nand U24755 (N_24755,N_19008,N_21610);
or U24756 (N_24756,N_18893,N_19413);
or U24757 (N_24757,N_18840,N_18789);
nor U24758 (N_24758,N_19595,N_21077);
or U24759 (N_24759,N_20315,N_21580);
or U24760 (N_24760,N_18989,N_21833);
and U24761 (N_24761,N_19666,N_21546);
and U24762 (N_24762,N_19744,N_20613);
nor U24763 (N_24763,N_20502,N_20586);
nor U24764 (N_24764,N_19514,N_18788);
or U24765 (N_24765,N_19410,N_21665);
xnor U24766 (N_24766,N_20065,N_20349);
or U24767 (N_24767,N_20647,N_21588);
nand U24768 (N_24768,N_21464,N_18850);
xnor U24769 (N_24769,N_20523,N_21198);
xnor U24770 (N_24770,N_19096,N_20549);
or U24771 (N_24771,N_21288,N_19006);
nand U24772 (N_24772,N_20679,N_18888);
nor U24773 (N_24773,N_21429,N_18875);
and U24774 (N_24774,N_20742,N_19991);
and U24775 (N_24775,N_19711,N_19423);
and U24776 (N_24776,N_21072,N_19545);
xor U24777 (N_24777,N_21322,N_19550);
nand U24778 (N_24778,N_20052,N_21432);
nand U24779 (N_24779,N_21148,N_20842);
or U24780 (N_24780,N_21506,N_20699);
or U24781 (N_24781,N_20280,N_21418);
nor U24782 (N_24782,N_19463,N_20816);
or U24783 (N_24783,N_21310,N_20437);
or U24784 (N_24784,N_19013,N_19460);
or U24785 (N_24785,N_19934,N_20926);
nand U24786 (N_24786,N_20665,N_20212);
or U24787 (N_24787,N_18884,N_19630);
nor U24788 (N_24788,N_19733,N_21615);
xnor U24789 (N_24789,N_21711,N_19819);
or U24790 (N_24790,N_20033,N_21567);
or U24791 (N_24791,N_18832,N_21461);
xor U24792 (N_24792,N_18902,N_20818);
and U24793 (N_24793,N_21404,N_21219);
or U24794 (N_24794,N_20499,N_20133);
nand U24795 (N_24795,N_21131,N_19387);
or U24796 (N_24796,N_20119,N_21867);
and U24797 (N_24797,N_19876,N_20002);
or U24798 (N_24798,N_18960,N_21361);
and U24799 (N_24799,N_20884,N_21291);
nor U24800 (N_24800,N_21300,N_21474);
and U24801 (N_24801,N_18961,N_21397);
nand U24802 (N_24802,N_21825,N_20360);
or U24803 (N_24803,N_21567,N_21808);
nor U24804 (N_24804,N_18815,N_20435);
nand U24805 (N_24805,N_21318,N_19521);
nand U24806 (N_24806,N_21205,N_20643);
and U24807 (N_24807,N_18973,N_21183);
xnor U24808 (N_24808,N_21337,N_21245);
nor U24809 (N_24809,N_20372,N_20540);
nor U24810 (N_24810,N_18997,N_20354);
xnor U24811 (N_24811,N_20013,N_18987);
xnor U24812 (N_24812,N_20237,N_19195);
or U24813 (N_24813,N_19602,N_20882);
or U24814 (N_24814,N_20220,N_21586);
or U24815 (N_24815,N_21581,N_19171);
nor U24816 (N_24816,N_21012,N_18855);
nor U24817 (N_24817,N_21245,N_21693);
or U24818 (N_24818,N_21208,N_21337);
nand U24819 (N_24819,N_19336,N_18825);
nor U24820 (N_24820,N_20585,N_21133);
and U24821 (N_24821,N_19457,N_19737);
or U24822 (N_24822,N_20720,N_19147);
or U24823 (N_24823,N_21264,N_19324);
and U24824 (N_24824,N_19371,N_18837);
or U24825 (N_24825,N_21727,N_21135);
xor U24826 (N_24826,N_20071,N_21858);
and U24827 (N_24827,N_19706,N_18803);
nand U24828 (N_24828,N_19635,N_20359);
nand U24829 (N_24829,N_19884,N_21166);
xnor U24830 (N_24830,N_19462,N_21678);
xor U24831 (N_24831,N_20830,N_19141);
xnor U24832 (N_24832,N_20739,N_18899);
nand U24833 (N_24833,N_19011,N_19562);
nand U24834 (N_24834,N_19878,N_20902);
xor U24835 (N_24835,N_20931,N_21248);
nor U24836 (N_24836,N_20868,N_20624);
nand U24837 (N_24837,N_19274,N_19266);
nor U24838 (N_24838,N_19265,N_20907);
nand U24839 (N_24839,N_19131,N_20259);
and U24840 (N_24840,N_19439,N_20764);
or U24841 (N_24841,N_19437,N_21310);
nor U24842 (N_24842,N_18776,N_18913);
nor U24843 (N_24843,N_19449,N_19288);
and U24844 (N_24844,N_20777,N_21281);
nor U24845 (N_24845,N_20870,N_20038);
and U24846 (N_24846,N_19445,N_21375);
and U24847 (N_24847,N_21723,N_21078);
or U24848 (N_24848,N_21698,N_21369);
and U24849 (N_24849,N_19315,N_19868);
or U24850 (N_24850,N_20107,N_19418);
or U24851 (N_24851,N_19686,N_20204);
or U24852 (N_24852,N_19617,N_21184);
or U24853 (N_24853,N_21423,N_18819);
or U24854 (N_24854,N_18831,N_20140);
and U24855 (N_24855,N_18844,N_20951);
xnor U24856 (N_24856,N_21779,N_21165);
nand U24857 (N_24857,N_18834,N_20599);
xor U24858 (N_24858,N_21312,N_20280);
nor U24859 (N_24859,N_19814,N_20311);
or U24860 (N_24860,N_20968,N_21276);
xor U24861 (N_24861,N_20999,N_21799);
xor U24862 (N_24862,N_21744,N_18979);
xnor U24863 (N_24863,N_20437,N_19458);
or U24864 (N_24864,N_19115,N_19818);
nand U24865 (N_24865,N_21727,N_19473);
nor U24866 (N_24866,N_20753,N_19954);
nor U24867 (N_24867,N_19535,N_21553);
or U24868 (N_24868,N_18760,N_20430);
xor U24869 (N_24869,N_19438,N_21755);
xnor U24870 (N_24870,N_19721,N_19606);
xor U24871 (N_24871,N_21484,N_20795);
and U24872 (N_24872,N_18818,N_20672);
and U24873 (N_24873,N_20509,N_19056);
nand U24874 (N_24874,N_21779,N_20295);
xor U24875 (N_24875,N_20743,N_21101);
and U24876 (N_24876,N_18797,N_18991);
nand U24877 (N_24877,N_21023,N_19307);
nor U24878 (N_24878,N_21307,N_21817);
and U24879 (N_24879,N_18884,N_20548);
and U24880 (N_24880,N_21608,N_20722);
xnor U24881 (N_24881,N_19159,N_20211);
nand U24882 (N_24882,N_19462,N_19686);
nand U24883 (N_24883,N_20288,N_20626);
and U24884 (N_24884,N_19184,N_20322);
nand U24885 (N_24885,N_19612,N_21092);
nor U24886 (N_24886,N_19906,N_20840);
xnor U24887 (N_24887,N_18875,N_19360);
or U24888 (N_24888,N_21739,N_19679);
nand U24889 (N_24889,N_19175,N_20117);
or U24890 (N_24890,N_21609,N_19818);
nand U24891 (N_24891,N_19087,N_19445);
and U24892 (N_24892,N_21118,N_20144);
and U24893 (N_24893,N_21772,N_18758);
and U24894 (N_24894,N_18953,N_20629);
and U24895 (N_24895,N_21114,N_19126);
xnor U24896 (N_24896,N_20809,N_18890);
nor U24897 (N_24897,N_21292,N_21216);
nor U24898 (N_24898,N_18975,N_18866);
nor U24899 (N_24899,N_19853,N_21789);
nand U24900 (N_24900,N_21499,N_21750);
or U24901 (N_24901,N_19518,N_21314);
or U24902 (N_24902,N_19735,N_20565);
nor U24903 (N_24903,N_20943,N_19654);
and U24904 (N_24904,N_19831,N_21035);
xnor U24905 (N_24905,N_21334,N_18990);
or U24906 (N_24906,N_20229,N_21224);
nor U24907 (N_24907,N_19688,N_19334);
and U24908 (N_24908,N_18846,N_21046);
and U24909 (N_24909,N_20095,N_19511);
nand U24910 (N_24910,N_21660,N_19512);
nand U24911 (N_24911,N_21041,N_19859);
or U24912 (N_24912,N_19114,N_21752);
or U24913 (N_24913,N_20636,N_19329);
nor U24914 (N_24914,N_18840,N_18855);
nor U24915 (N_24915,N_21464,N_20046);
xor U24916 (N_24916,N_19421,N_19404);
xnor U24917 (N_24917,N_21212,N_21835);
nor U24918 (N_24918,N_20491,N_21212);
nor U24919 (N_24919,N_21033,N_19110);
nand U24920 (N_24920,N_21763,N_20878);
or U24921 (N_24921,N_21530,N_21182);
xor U24922 (N_24922,N_19665,N_21080);
xnor U24923 (N_24923,N_19049,N_21334);
or U24924 (N_24924,N_20921,N_20360);
nand U24925 (N_24925,N_19740,N_19668);
or U24926 (N_24926,N_19872,N_18965);
xnor U24927 (N_24927,N_19752,N_18985);
nand U24928 (N_24928,N_19666,N_20614);
xor U24929 (N_24929,N_20365,N_20688);
xnor U24930 (N_24930,N_18990,N_21614);
or U24931 (N_24931,N_19685,N_21459);
nand U24932 (N_24932,N_18852,N_20854);
xor U24933 (N_24933,N_18811,N_21372);
nor U24934 (N_24934,N_21562,N_19309);
and U24935 (N_24935,N_20550,N_20032);
or U24936 (N_24936,N_20582,N_21288);
and U24937 (N_24937,N_20040,N_19526);
xnor U24938 (N_24938,N_20734,N_19646);
and U24939 (N_24939,N_20024,N_21756);
nand U24940 (N_24940,N_20697,N_20290);
xor U24941 (N_24941,N_19202,N_19760);
nor U24942 (N_24942,N_19904,N_20820);
or U24943 (N_24943,N_21427,N_20670);
and U24944 (N_24944,N_20885,N_20927);
and U24945 (N_24945,N_20106,N_20759);
xor U24946 (N_24946,N_21549,N_20604);
and U24947 (N_24947,N_20784,N_20200);
nor U24948 (N_24948,N_18832,N_21238);
xnor U24949 (N_24949,N_19821,N_20130);
xor U24950 (N_24950,N_21753,N_20052);
nor U24951 (N_24951,N_20050,N_20885);
and U24952 (N_24952,N_20512,N_21493);
nand U24953 (N_24953,N_20756,N_20792);
or U24954 (N_24954,N_20810,N_19334);
or U24955 (N_24955,N_19161,N_21492);
nand U24956 (N_24956,N_21826,N_21183);
nor U24957 (N_24957,N_19720,N_20472);
nand U24958 (N_24958,N_19653,N_21322);
nand U24959 (N_24959,N_19513,N_20976);
nor U24960 (N_24960,N_21153,N_19799);
xor U24961 (N_24961,N_19491,N_21466);
nand U24962 (N_24962,N_20514,N_19616);
and U24963 (N_24963,N_20270,N_20965);
or U24964 (N_24964,N_21117,N_21540);
nand U24965 (N_24965,N_19825,N_20666);
xnor U24966 (N_24966,N_20070,N_19598);
nor U24967 (N_24967,N_21500,N_20717);
nor U24968 (N_24968,N_19260,N_19463);
or U24969 (N_24969,N_21595,N_20589);
or U24970 (N_24970,N_20278,N_20971);
nor U24971 (N_24971,N_21413,N_19826);
xnor U24972 (N_24972,N_21265,N_19966);
or U24973 (N_24973,N_21503,N_19697);
nand U24974 (N_24974,N_18901,N_19256);
nor U24975 (N_24975,N_18772,N_21225);
xnor U24976 (N_24976,N_21373,N_18893);
and U24977 (N_24977,N_19845,N_21510);
nand U24978 (N_24978,N_20610,N_21832);
xnor U24979 (N_24979,N_19803,N_20716);
xor U24980 (N_24980,N_18823,N_18837);
or U24981 (N_24981,N_19392,N_21020);
nor U24982 (N_24982,N_21499,N_21538);
nand U24983 (N_24983,N_20466,N_19233);
xnor U24984 (N_24984,N_19739,N_19462);
nand U24985 (N_24985,N_19647,N_19455);
nand U24986 (N_24986,N_21320,N_20588);
and U24987 (N_24987,N_20067,N_19019);
nand U24988 (N_24988,N_20148,N_19665);
or U24989 (N_24989,N_21096,N_19389);
nand U24990 (N_24990,N_20867,N_19848);
nor U24991 (N_24991,N_20507,N_21336);
nand U24992 (N_24992,N_19690,N_20277);
or U24993 (N_24993,N_20218,N_20311);
and U24994 (N_24994,N_21401,N_19775);
and U24995 (N_24995,N_19568,N_20271);
nand U24996 (N_24996,N_19188,N_21690);
nand U24997 (N_24997,N_19527,N_20356);
or U24998 (N_24998,N_19489,N_20986);
nand U24999 (N_24999,N_18817,N_21710);
and UO_0 (O_0,N_22233,N_23554);
nand UO_1 (O_1,N_24567,N_21900);
nand UO_2 (O_2,N_24491,N_24195);
xor UO_3 (O_3,N_22383,N_24202);
and UO_4 (O_4,N_22129,N_23411);
nor UO_5 (O_5,N_22931,N_23877);
nand UO_6 (O_6,N_24685,N_22526);
or UO_7 (O_7,N_24780,N_23794);
nand UO_8 (O_8,N_23912,N_22196);
nor UO_9 (O_9,N_22636,N_22436);
nor UO_10 (O_10,N_24050,N_24931);
nor UO_11 (O_11,N_21926,N_22901);
nor UO_12 (O_12,N_23125,N_22193);
nor UO_13 (O_13,N_23867,N_22794);
xor UO_14 (O_14,N_22126,N_23578);
or UO_15 (O_15,N_24185,N_22684);
xor UO_16 (O_16,N_23961,N_22364);
xnor UO_17 (O_17,N_24583,N_22951);
nor UO_18 (O_18,N_23328,N_24792);
nand UO_19 (O_19,N_24680,N_23044);
xnor UO_20 (O_20,N_22162,N_22868);
and UO_21 (O_21,N_24521,N_24681);
and UO_22 (O_22,N_24946,N_24452);
nor UO_23 (O_23,N_23937,N_22910);
nor UO_24 (O_24,N_22187,N_24080);
nor UO_25 (O_25,N_22004,N_22914);
xor UO_26 (O_26,N_24163,N_22522);
or UO_27 (O_27,N_24389,N_22155);
or UO_28 (O_28,N_23262,N_23988);
or UO_29 (O_29,N_24973,N_23413);
and UO_30 (O_30,N_22106,N_24371);
and UO_31 (O_31,N_22874,N_24287);
nand UO_32 (O_32,N_23268,N_22616);
xor UO_33 (O_33,N_22229,N_22147);
and UO_34 (O_34,N_24714,N_23368);
nor UO_35 (O_35,N_21959,N_22928);
xor UO_36 (O_36,N_24426,N_24630);
or UO_37 (O_37,N_24127,N_22721);
and UO_38 (O_38,N_24300,N_24326);
xnor UO_39 (O_39,N_22834,N_22241);
or UO_40 (O_40,N_23661,N_23558);
and UO_41 (O_41,N_22633,N_24343);
nand UO_42 (O_42,N_23821,N_22897);
nand UO_43 (O_43,N_22444,N_22300);
or UO_44 (O_44,N_23491,N_22393);
nand UO_45 (O_45,N_23565,N_23976);
and UO_46 (O_46,N_24038,N_24514);
or UO_47 (O_47,N_21876,N_24713);
xnor UO_48 (O_48,N_24333,N_23560);
nand UO_49 (O_49,N_23589,N_23398);
and UO_50 (O_50,N_23727,N_22325);
nand UO_51 (O_51,N_24023,N_23403);
nand UO_52 (O_52,N_24891,N_22320);
or UO_53 (O_53,N_24064,N_22552);
nand UO_54 (O_54,N_22370,N_24575);
xor UO_55 (O_55,N_23534,N_22230);
or UO_56 (O_56,N_24447,N_24264);
nand UO_57 (O_57,N_22301,N_23124);
nor UO_58 (O_58,N_24402,N_24912);
nand UO_59 (O_59,N_24315,N_22074);
and UO_60 (O_60,N_24803,N_24800);
and UO_61 (O_61,N_24392,N_23255);
nand UO_62 (O_62,N_24766,N_22576);
nor UO_63 (O_63,N_23468,N_24313);
and UO_64 (O_64,N_22698,N_24500);
nor UO_65 (O_65,N_23715,N_22278);
and UO_66 (O_66,N_22679,N_23162);
nor UO_67 (O_67,N_23990,N_24352);
nand UO_68 (O_68,N_24588,N_24274);
and UO_69 (O_69,N_24344,N_22857);
xor UO_70 (O_70,N_22140,N_21949);
nor UO_71 (O_71,N_23060,N_24558);
nor UO_72 (O_72,N_23977,N_22945);
or UO_73 (O_73,N_24571,N_22823);
and UO_74 (O_74,N_23816,N_24290);
xor UO_75 (O_75,N_23296,N_22206);
xnor UO_76 (O_76,N_23720,N_22317);
nand UO_77 (O_77,N_23771,N_24542);
nor UO_78 (O_78,N_24063,N_24472);
and UO_79 (O_79,N_22561,N_23819);
nor UO_80 (O_80,N_24553,N_23460);
nand UO_81 (O_81,N_23101,N_24996);
nor UO_82 (O_82,N_23023,N_24718);
xor UO_83 (O_83,N_22188,N_22866);
or UO_84 (O_84,N_24014,N_23904);
xor UO_85 (O_85,N_24088,N_24879);
and UO_86 (O_86,N_23929,N_24148);
and UO_87 (O_87,N_22541,N_24232);
and UO_88 (O_88,N_22549,N_24446);
xnor UO_89 (O_89,N_22094,N_24723);
nor UO_90 (O_90,N_23301,N_22982);
nor UO_91 (O_91,N_24475,N_24179);
nand UO_92 (O_92,N_22856,N_24243);
nor UO_93 (O_93,N_22680,N_23782);
xor UO_94 (O_94,N_24546,N_22000);
or UO_95 (O_95,N_24046,N_24485);
nor UO_96 (O_96,N_24880,N_23569);
nor UO_97 (O_97,N_24811,N_23212);
or UO_98 (O_98,N_23884,N_24114);
nand UO_99 (O_99,N_24019,N_22511);
nor UO_100 (O_100,N_22539,N_24209);
nand UO_101 (O_101,N_22906,N_24421);
nand UO_102 (O_102,N_22305,N_22777);
and UO_103 (O_103,N_21915,N_23437);
and UO_104 (O_104,N_23797,N_24851);
and UO_105 (O_105,N_23555,N_24192);
nor UO_106 (O_106,N_23725,N_22893);
xor UO_107 (O_107,N_23055,N_22256);
nor UO_108 (O_108,N_23145,N_24486);
nor UO_109 (O_109,N_23454,N_24471);
and UO_110 (O_110,N_24166,N_23732);
nand UO_111 (O_111,N_23637,N_23756);
xnor UO_112 (O_112,N_23859,N_23553);
nor UO_113 (O_113,N_24438,N_24104);
or UO_114 (O_114,N_23066,N_21904);
nand UO_115 (O_115,N_23195,N_24024);
nand UO_116 (O_116,N_22583,N_23864);
and UO_117 (O_117,N_23186,N_22782);
nand UO_118 (O_118,N_22845,N_23199);
or UO_119 (O_119,N_23742,N_24566);
xnor UO_120 (O_120,N_23285,N_24115);
or UO_121 (O_121,N_24218,N_22340);
xnor UO_122 (O_122,N_24327,N_24769);
nor UO_123 (O_123,N_23830,N_22032);
or UO_124 (O_124,N_24175,N_22975);
and UO_125 (O_125,N_21922,N_23071);
xnor UO_126 (O_126,N_24985,N_22416);
xor UO_127 (O_127,N_22767,N_23025);
and UO_128 (O_128,N_22833,N_23012);
and UO_129 (O_129,N_24683,N_23180);
or UO_130 (O_130,N_23813,N_22167);
or UO_131 (O_131,N_24688,N_22635);
nor UO_132 (O_132,N_22114,N_22025);
nand UO_133 (O_133,N_24173,N_24642);
xnor UO_134 (O_134,N_24258,N_24276);
and UO_135 (O_135,N_24933,N_23417);
nand UO_136 (O_136,N_24339,N_22521);
or UO_137 (O_137,N_22817,N_23905);
xor UO_138 (O_138,N_23731,N_23277);
or UO_139 (O_139,N_23545,N_23002);
nor UO_140 (O_140,N_23440,N_24081);
or UO_141 (O_141,N_24084,N_24806);
nand UO_142 (O_142,N_22389,N_24599);
xor UO_143 (O_143,N_21917,N_23920);
nor UO_144 (O_144,N_24510,N_23393);
nor UO_145 (O_145,N_23040,N_22858);
xnor UO_146 (O_146,N_22769,N_24760);
and UO_147 (O_147,N_22048,N_23171);
and UO_148 (O_148,N_22217,N_24922);
nand UO_149 (O_149,N_22729,N_24272);
xor UO_150 (O_150,N_22262,N_24573);
and UO_151 (O_151,N_23709,N_23480);
and UO_152 (O_152,N_22771,N_23295);
or UO_153 (O_153,N_23246,N_22429);
nand UO_154 (O_154,N_22495,N_22981);
and UO_155 (O_155,N_22708,N_22704);
nor UO_156 (O_156,N_24894,N_23383);
nor UO_157 (O_157,N_21875,N_22151);
or UO_158 (O_158,N_23376,N_22061);
nand UO_159 (O_159,N_24751,N_24887);
nand UO_160 (O_160,N_23367,N_22850);
or UO_161 (O_161,N_24487,N_22702);
nand UO_162 (O_162,N_24490,N_23549);
xnor UO_163 (O_163,N_22201,N_24710);
nand UO_164 (O_164,N_23897,N_23613);
xnor UO_165 (O_165,N_24260,N_23671);
and UO_166 (O_166,N_22503,N_24134);
xor UO_167 (O_167,N_23138,N_23871);
and UO_168 (O_168,N_23128,N_23911);
nand UO_169 (O_169,N_23619,N_24464);
or UO_170 (O_170,N_22524,N_22741);
and UO_171 (O_171,N_24493,N_22117);
xnor UO_172 (O_172,N_23665,N_22962);
and UO_173 (O_173,N_23548,N_23759);
or UO_174 (O_174,N_23508,N_22052);
or UO_175 (O_175,N_21897,N_22245);
nor UO_176 (O_176,N_22251,N_22620);
nand UO_177 (O_177,N_22428,N_24118);
and UO_178 (O_178,N_22697,N_23364);
nor UO_179 (O_179,N_22123,N_22827);
nand UO_180 (O_180,N_22695,N_24897);
or UO_181 (O_181,N_22351,N_22984);
and UO_182 (O_182,N_24716,N_24194);
xnor UO_183 (O_183,N_24737,N_22186);
or UO_184 (O_184,N_22222,N_23846);
nor UO_185 (O_185,N_21913,N_21910);
nand UO_186 (O_186,N_24210,N_22792);
or UO_187 (O_187,N_24055,N_24161);
nand UO_188 (O_188,N_22963,N_22289);
xnor UO_189 (O_189,N_23447,N_24372);
xnor UO_190 (O_190,N_22231,N_24577);
and UO_191 (O_191,N_24635,N_23372);
nand UO_192 (O_192,N_22734,N_24741);
nand UO_193 (O_193,N_24225,N_23236);
and UO_194 (O_194,N_23792,N_24355);
xnor UO_195 (O_195,N_24137,N_24484);
xnor UO_196 (O_196,N_23390,N_22744);
nand UO_197 (O_197,N_23728,N_23357);
nor UO_198 (O_198,N_23203,N_23122);
or UO_199 (O_199,N_23993,N_24382);
nor UO_200 (O_200,N_24470,N_23768);
nor UO_201 (O_201,N_22655,N_24199);
and UO_202 (O_202,N_23348,N_24017);
xnor UO_203 (O_203,N_24431,N_22136);
and UO_204 (O_204,N_24810,N_22663);
xnor UO_205 (O_205,N_24331,N_24949);
xor UO_206 (O_206,N_22432,N_24744);
and UO_207 (O_207,N_24957,N_22479);
nand UO_208 (O_208,N_24458,N_22049);
or UO_209 (O_209,N_22098,N_22091);
xnor UO_210 (O_210,N_21933,N_23583);
or UO_211 (O_211,N_23785,N_24970);
nand UO_212 (O_212,N_24018,N_24095);
and UO_213 (O_213,N_22615,N_22176);
and UO_214 (O_214,N_22892,N_24587);
and UO_215 (O_215,N_23238,N_24420);
xnor UO_216 (O_216,N_22518,N_23762);
xor UO_217 (O_217,N_23200,N_22623);
nand UO_218 (O_218,N_23866,N_24704);
and UO_219 (O_219,N_22344,N_23230);
or UO_220 (O_220,N_23313,N_22992);
or UO_221 (O_221,N_22976,N_22730);
and UO_222 (O_222,N_22360,N_22438);
and UO_223 (O_223,N_23588,N_22418);
or UO_224 (O_224,N_23266,N_24460);
nand UO_225 (O_225,N_22439,N_22824);
nor UO_226 (O_226,N_23457,N_24633);
or UO_227 (O_227,N_23421,N_23123);
or UO_228 (O_228,N_24404,N_24036);
or UO_229 (O_229,N_23093,N_23068);
nor UO_230 (O_230,N_24862,N_24666);
or UO_231 (O_231,N_23042,N_22394);
or UO_232 (O_232,N_21962,N_24374);
or UO_233 (O_233,N_23449,N_23807);
and UO_234 (O_234,N_22884,N_22781);
nand UO_235 (O_235,N_23327,N_22875);
nand UO_236 (O_236,N_23706,N_22650);
nor UO_237 (O_237,N_23174,N_23156);
and UO_238 (O_238,N_22321,N_23227);
or UO_239 (O_239,N_22397,N_24787);
or UO_240 (O_240,N_22002,N_23280);
nor UO_241 (O_241,N_22160,N_22425);
or UO_242 (O_242,N_22409,N_23218);
xor UO_243 (O_243,N_24693,N_24886);
nor UO_244 (O_244,N_24477,N_22727);
and UO_245 (O_245,N_24299,N_22571);
xor UO_246 (O_246,N_23169,N_24479);
or UO_247 (O_247,N_23420,N_21920);
xnor UO_248 (O_248,N_22337,N_22930);
xnor UO_249 (O_249,N_22149,N_24815);
or UO_250 (O_250,N_23552,N_22017);
nor UO_251 (O_251,N_21963,N_22917);
or UO_252 (O_252,N_23134,N_24964);
and UO_253 (O_253,N_24212,N_21908);
xnor UO_254 (O_254,N_24291,N_22433);
nand UO_255 (O_255,N_24021,N_24691);
and UO_256 (O_256,N_23129,N_23486);
xor UO_257 (O_257,N_21894,N_23177);
and UO_258 (O_258,N_22240,N_22603);
nor UO_259 (O_259,N_22082,N_22630);
nor UO_260 (O_260,N_24293,N_24898);
and UO_261 (O_261,N_22332,N_22941);
xnor UO_262 (O_262,N_24468,N_24122);
nor UO_263 (O_263,N_24695,N_22467);
nand UO_264 (O_264,N_24268,N_22372);
nand UO_265 (O_265,N_22821,N_23292);
nand UO_266 (O_266,N_22366,N_22844);
xor UO_267 (O_267,N_22277,N_24100);
or UO_268 (O_268,N_22644,N_23844);
nand UO_269 (O_269,N_24568,N_22352);
xor UO_270 (O_270,N_24047,N_24582);
nor UO_271 (O_271,N_22967,N_24121);
xnor UO_272 (O_272,N_23939,N_23751);
nor UO_273 (O_273,N_23953,N_23450);
or UO_274 (O_274,N_22200,N_21948);
and UO_275 (O_275,N_22216,N_24216);
or UO_276 (O_276,N_24837,N_22979);
or UO_277 (O_277,N_22926,N_22588);
nand UO_278 (O_278,N_22682,N_24604);
xor UO_279 (O_279,N_24987,N_22653);
and UO_280 (O_280,N_23187,N_22146);
nand UO_281 (O_281,N_23251,N_22512);
xnor UO_282 (O_282,N_23196,N_23256);
and UO_283 (O_283,N_24052,N_24307);
or UO_284 (O_284,N_22543,N_22185);
or UO_285 (O_285,N_24881,N_24759);
or UO_286 (O_286,N_22401,N_22796);
nor UO_287 (O_287,N_22086,N_24853);
xor UO_288 (O_288,N_23660,N_24842);
and UO_289 (O_289,N_23316,N_23823);
and UO_290 (O_290,N_24578,N_22924);
or UO_291 (O_291,N_24170,N_24972);
or UO_292 (O_292,N_23764,N_22538);
and UO_293 (O_293,N_23155,N_24532);
nand UO_294 (O_294,N_22271,N_22058);
or UO_295 (O_295,N_22248,N_24926);
nor UO_296 (O_296,N_24932,N_23860);
nor UO_297 (O_297,N_24407,N_24113);
nand UO_298 (O_298,N_24858,N_23108);
xor UO_299 (O_299,N_22775,N_23705);
or UO_300 (O_300,N_23708,N_24742);
nor UO_301 (O_301,N_24923,N_23163);
nand UO_302 (O_302,N_23336,N_22159);
xnor UO_303 (O_303,N_24241,N_24435);
and UO_304 (O_304,N_22172,N_22656);
nor UO_305 (O_305,N_24869,N_24359);
xnor UO_306 (O_306,N_22090,N_21945);
xnor UO_307 (O_307,N_24412,N_24444);
and UO_308 (O_308,N_24208,N_23003);
xnor UO_309 (O_309,N_24778,N_23104);
xor UO_310 (O_310,N_24997,N_22051);
or UO_311 (O_311,N_23621,N_24156);
nand UO_312 (O_312,N_22840,N_23925);
nor UO_313 (O_313,N_24528,N_23304);
or UO_314 (O_314,N_23410,N_22865);
nor UO_315 (O_315,N_24775,N_24367);
xor UO_316 (O_316,N_23472,N_23306);
nand UO_317 (O_317,N_24207,N_22731);
nand UO_318 (O_318,N_23309,N_24512);
xnor UO_319 (O_319,N_23435,N_24915);
and UO_320 (O_320,N_22218,N_23926);
nand UO_321 (O_321,N_22660,N_24469);
nand UO_322 (O_322,N_24884,N_23710);
nor UO_323 (O_323,N_24702,N_23428);
or UO_324 (O_324,N_22475,N_23644);
and UO_325 (O_325,N_22101,N_24091);
or UO_326 (O_326,N_24498,N_23919);
xor UO_327 (O_327,N_23158,N_22312);
or UO_328 (O_328,N_23895,N_24016);
nor UO_329 (O_329,N_24033,N_22311);
xnor UO_330 (O_330,N_23514,N_23757);
and UO_331 (O_331,N_23736,N_22270);
or UO_332 (O_332,N_23379,N_23974);
nand UO_333 (O_333,N_22053,N_23576);
nand UO_334 (O_334,N_24011,N_24941);
nor UO_335 (O_335,N_22198,N_23452);
nand UO_336 (O_336,N_24400,N_24502);
nand UO_337 (O_337,N_22470,N_24660);
nand UO_338 (O_338,N_22132,N_23017);
and UO_339 (O_339,N_24074,N_23408);
xnor UO_340 (O_340,N_24709,N_22828);
nand UO_341 (O_341,N_23533,N_24865);
nand UO_342 (O_342,N_23011,N_23634);
and UO_343 (O_343,N_24570,N_22182);
nor UO_344 (O_344,N_22128,N_23622);
xnor UO_345 (O_345,N_22402,N_23184);
nor UO_346 (O_346,N_23636,N_22838);
xnor UO_347 (O_347,N_22851,N_24096);
or UO_348 (O_348,N_22465,N_22944);
or UO_349 (O_349,N_23355,N_23274);
and UO_350 (O_350,N_22011,N_23574);
and UO_351 (O_351,N_22022,N_24864);
nor UO_352 (O_352,N_24230,N_24106);
and UO_353 (O_353,N_24614,N_24843);
xor UO_354 (O_354,N_23284,N_23876);
nor UO_355 (O_355,N_24379,N_22871);
or UO_356 (O_356,N_23617,N_24146);
and UO_357 (O_357,N_23392,N_24041);
nor UO_358 (O_358,N_23258,N_23117);
and UO_359 (O_359,N_24988,N_22390);
and UO_360 (O_360,N_24628,N_24375);
xor UO_361 (O_361,N_24678,N_21968);
nand UO_362 (O_362,N_23252,N_24552);
xnor UO_363 (O_363,N_24860,N_22560);
xor UO_364 (O_364,N_24103,N_22629);
xor UO_365 (O_365,N_24828,N_22158);
nor UO_366 (O_366,N_24105,N_23065);
and UO_367 (O_367,N_22122,N_23837);
nand UO_368 (O_368,N_24925,N_22386);
or UO_369 (O_369,N_23726,N_24004);
nand UO_370 (O_370,N_24273,N_24085);
nor UO_371 (O_371,N_23182,N_24619);
xor UO_372 (O_372,N_23091,N_24377);
or UO_373 (O_373,N_23159,N_22861);
or UO_374 (O_374,N_23760,N_23509);
nand UO_375 (O_375,N_23423,N_22986);
and UO_376 (O_376,N_23311,N_24945);
or UO_377 (O_377,N_22566,N_23210);
or UO_378 (O_378,N_24826,N_24267);
nor UO_379 (O_379,N_24748,N_23701);
xnor UO_380 (O_380,N_22716,N_22570);
and UO_381 (O_381,N_22493,N_23224);
or UO_382 (O_382,N_22725,N_22318);
and UO_383 (O_383,N_24872,N_24461);
nor UO_384 (O_384,N_23147,N_24870);
or UO_385 (O_385,N_24560,N_22039);
nor UO_386 (O_386,N_24319,N_21911);
xor UO_387 (O_387,N_23834,N_23586);
and UO_388 (O_388,N_23907,N_23638);
or UO_389 (O_389,N_21928,N_21919);
nor UO_390 (O_390,N_22168,N_21966);
and UO_391 (O_391,N_23085,N_24270);
nand UO_392 (O_392,N_23829,N_23116);
nand UO_393 (O_393,N_22121,N_24594);
and UO_394 (O_394,N_24430,N_22480);
nand UO_395 (O_395,N_22846,N_22613);
and UO_396 (O_396,N_23190,N_24002);
nor UO_397 (O_397,N_22079,N_22646);
xnor UO_398 (O_398,N_23633,N_23080);
or UO_399 (O_399,N_24012,N_23319);
and UO_400 (O_400,N_24190,N_23019);
xnor UO_401 (O_401,N_24804,N_24735);
or UO_402 (O_402,N_22285,N_23944);
nand UO_403 (O_403,N_22363,N_22878);
or UO_404 (O_404,N_23083,N_24868);
nor UO_405 (O_405,N_23902,N_22210);
and UO_406 (O_406,N_24523,N_23838);
or UO_407 (O_407,N_23310,N_23400);
and UO_408 (O_408,N_24437,N_23173);
nand UO_409 (O_409,N_22195,N_22486);
or UO_410 (O_410,N_23484,N_23445);
xnor UO_411 (O_411,N_24473,N_24511);
and UO_412 (O_412,N_21957,N_22863);
or UO_413 (O_413,N_24911,N_23662);
xor UO_414 (O_414,N_24158,N_22324);
and UO_415 (O_415,N_23110,N_22530);
and UO_416 (O_416,N_22042,N_22338);
or UO_417 (O_417,N_24962,N_23409);
and UO_418 (O_418,N_22908,N_24506);
xor UO_419 (O_419,N_24701,N_22887);
nand UO_420 (O_420,N_24058,N_23027);
xor UO_421 (O_421,N_22062,N_23361);
nand UO_422 (O_422,N_24358,N_24284);
nor UO_423 (O_423,N_24918,N_22208);
nor UO_424 (O_424,N_24155,N_23980);
nand UO_425 (O_425,N_24538,N_22023);
and UO_426 (O_426,N_23719,N_24390);
or UO_427 (O_427,N_24895,N_23370);
nand UO_428 (O_428,N_24598,N_22896);
nor UO_429 (O_429,N_24770,N_23526);
xnor UO_430 (O_430,N_23916,N_24537);
and UO_431 (O_431,N_24168,N_24237);
xor UO_432 (O_432,N_22314,N_23739);
and UO_433 (O_433,N_22400,N_23828);
nor UO_434 (O_434,N_23243,N_22097);
or UO_435 (O_435,N_23097,N_23796);
nor UO_436 (O_436,N_24336,N_23927);
nor UO_437 (O_437,N_22026,N_24449);
and UO_438 (O_438,N_23873,N_22812);
and UO_439 (O_439,N_23247,N_23324);
xnor UO_440 (O_440,N_24001,N_24772);
or UO_441 (O_441,N_22988,N_22738);
and UO_442 (O_442,N_24160,N_24312);
and UO_443 (O_443,N_24125,N_23581);
or UO_444 (O_444,N_22542,N_22891);
xnor UO_445 (O_445,N_22855,N_22341);
nor UO_446 (O_446,N_22507,N_23780);
xor UO_447 (O_447,N_24833,N_23338);
xor UO_448 (O_448,N_22830,N_23249);
nor UO_449 (O_449,N_23299,N_23941);
nand UO_450 (O_450,N_22423,N_23786);
nor UO_451 (O_451,N_24227,N_23146);
or UO_452 (O_452,N_23127,N_24857);
nor UO_453 (O_453,N_24903,N_24650);
or UO_454 (O_454,N_22396,N_24689);
nor UO_455 (O_455,N_22308,N_23385);
and UO_456 (O_456,N_22489,N_23512);
and UO_457 (O_457,N_24774,N_22102);
nor UO_458 (O_458,N_22808,N_23758);
and UO_459 (O_459,N_24234,N_23700);
and UO_460 (O_460,N_24265,N_23778);
xor UO_461 (O_461,N_23033,N_24405);
and UO_462 (O_462,N_22134,N_22220);
xnor UO_463 (O_463,N_22701,N_22001);
nand UO_464 (O_464,N_22747,N_24783);
nor UO_465 (O_465,N_22717,N_21885);
or UO_466 (O_466,N_22700,N_24269);
and UO_467 (O_467,N_23716,N_23888);
xnor UO_468 (O_468,N_24631,N_22460);
nand UO_469 (O_469,N_24441,N_23874);
nor UO_470 (O_470,N_24971,N_23718);
or UO_471 (O_471,N_23973,N_22783);
and UO_472 (O_472,N_23442,N_24998);
or UO_473 (O_473,N_24056,N_22385);
nor UO_474 (O_474,N_22421,N_23989);
or UO_475 (O_475,N_22184,N_24061);
and UO_476 (O_476,N_23652,N_24520);
or UO_477 (O_477,N_24981,N_23443);
or UO_478 (O_478,N_23614,N_22388);
nand UO_479 (O_479,N_23618,N_24669);
nand UO_480 (O_480,N_22719,N_22533);
nor UO_481 (O_481,N_23487,N_22699);
nand UO_482 (O_482,N_22683,N_24878);
or UO_483 (O_483,N_24728,N_24424);
nor UO_484 (O_484,N_23414,N_22957);
xnor UO_485 (O_485,N_23878,N_22205);
nand UO_486 (O_486,N_24888,N_23639);
nand UO_487 (O_487,N_24455,N_24755);
xor UO_488 (O_488,N_24940,N_22440);
or UO_489 (O_489,N_24409,N_23084);
xnor UO_490 (O_490,N_23943,N_23691);
nand UO_491 (O_491,N_22822,N_21951);
nand UO_492 (O_492,N_22832,N_23841);
nor UO_493 (O_493,N_23903,N_24443);
xnor UO_494 (O_494,N_23049,N_24224);
or UO_495 (O_495,N_24341,N_24786);
or UO_496 (O_496,N_23371,N_24476);
and UO_497 (O_497,N_24610,N_22651);
or UO_498 (O_498,N_24892,N_24671);
nor UO_499 (O_499,N_23046,N_23193);
or UO_500 (O_500,N_24527,N_23050);
or UO_501 (O_501,N_24522,N_22648);
or UO_502 (O_502,N_23303,N_24924);
nand UO_503 (O_503,N_22471,N_22797);
xnor UO_504 (O_504,N_23682,N_23279);
and UO_505 (O_505,N_24251,N_24346);
nand UO_506 (O_506,N_24679,N_23955);
nor UO_507 (O_507,N_23154,N_22490);
or UO_508 (O_508,N_22912,N_22282);
nor UO_509 (O_509,N_23183,N_24048);
nor UO_510 (O_510,N_24788,N_22793);
or UO_511 (O_511,N_24761,N_24697);
xor UO_512 (O_512,N_22169,N_24261);
nor UO_513 (O_513,N_22224,N_21992);
nand UO_514 (O_514,N_22803,N_23353);
or UO_515 (O_515,N_22257,N_23213);
nand UO_516 (O_516,N_23496,N_23109);
xor UO_517 (O_517,N_21888,N_21895);
nand UO_518 (O_518,N_21931,N_22923);
nand UO_519 (O_519,N_24936,N_24044);
nand UO_520 (O_520,N_24626,N_23765);
and UO_521 (O_521,N_22676,N_22627);
xor UO_522 (O_522,N_23772,N_23697);
and UO_523 (O_523,N_22575,N_22007);
or UO_524 (O_524,N_23086,N_21987);
and UO_525 (O_525,N_22255,N_24656);
or UO_526 (O_526,N_23237,N_22802);
or UO_527 (O_527,N_24157,N_23118);
nand UO_528 (O_528,N_23426,N_22247);
nand UO_529 (O_529,N_22774,N_22578);
nand UO_530 (O_530,N_22485,N_22628);
nand UO_531 (O_531,N_24057,N_23650);
and UO_532 (O_532,N_23857,N_22014);
or UO_533 (O_533,N_22590,N_24591);
nand UO_534 (O_534,N_23465,N_23375);
nor UO_535 (O_535,N_21890,N_22509);
nor UO_536 (O_536,N_22327,N_23580);
nor UO_537 (O_537,N_22089,N_23887);
and UO_538 (O_538,N_21935,N_24356);
or UO_539 (O_539,N_22577,N_22843);
or UO_540 (O_540,N_23235,N_22545);
and UO_541 (O_541,N_23967,N_22903);
xnor UO_542 (O_542,N_22594,N_23202);
or UO_543 (O_543,N_22936,N_23096);
nor UO_544 (O_544,N_24953,N_24545);
xnor UO_545 (O_545,N_23167,N_23730);
and UO_546 (O_546,N_23861,N_23282);
xnor UO_547 (O_547,N_22348,N_22661);
xor UO_548 (O_548,N_23611,N_22319);
nand UO_549 (O_549,N_22293,N_24664);
nor UO_550 (O_550,N_23001,N_24661);
nand UO_551 (O_551,N_23219,N_23666);
and UO_552 (O_552,N_24275,N_23843);
nand UO_553 (O_553,N_22095,N_24228);
or UO_554 (O_554,N_23142,N_24342);
nand UO_555 (O_555,N_22687,N_23818);
nand UO_556 (O_556,N_22772,N_24734);
nor UO_557 (O_557,N_23500,N_22018);
nand UO_558 (O_558,N_23775,N_24754);
and UO_559 (O_559,N_22839,N_23945);
and UO_560 (O_560,N_24239,N_24525);
xor UO_561 (O_561,N_23041,N_24928);
and UO_562 (O_562,N_22961,N_24423);
xnor UO_563 (O_563,N_24306,N_23590);
xnor UO_564 (O_564,N_22347,N_22818);
or UO_565 (O_565,N_24135,N_22529);
nor UO_566 (O_566,N_21930,N_24015);
xnor UO_567 (O_567,N_23678,N_23951);
or UO_568 (O_568,N_24551,N_22252);
nor UO_569 (O_569,N_22109,N_23208);
and UO_570 (O_570,N_24615,N_24060);
xor UO_571 (O_571,N_24397,N_22622);
nand UO_572 (O_572,N_24698,N_24150);
or UO_573 (O_573,N_24823,N_23194);
nand UO_574 (O_574,N_22582,N_23568);
xnor UO_575 (O_575,N_24623,N_23330);
nor UO_576 (O_576,N_24550,N_24226);
nand UO_577 (O_577,N_23165,N_23014);
or UO_578 (O_578,N_24885,N_24739);
and UO_579 (O_579,N_22130,N_22044);
xor UO_580 (O_580,N_23938,N_24325);
or UO_581 (O_581,N_22115,N_22713);
xnor UO_582 (O_582,N_22426,N_23248);
or UO_583 (O_583,N_24031,N_23098);
nor UO_584 (O_584,N_24222,N_21923);
and UO_585 (O_585,N_24139,N_24674);
or UO_586 (O_586,N_24724,N_23488);
nor UO_587 (O_587,N_22551,N_24517);
and UO_588 (O_588,N_22357,N_22870);
xnor UO_589 (O_589,N_24627,N_24927);
nor UO_590 (O_590,N_24830,N_24585);
nor UO_591 (O_591,N_22228,N_22361);
xor UO_592 (O_592,N_22299,N_24182);
and UO_593 (O_593,N_23769,N_24247);
nand UO_594 (O_594,N_23052,N_22586);
or UO_595 (O_595,N_24129,N_24429);
xnor UO_596 (O_596,N_23471,N_23175);
nor UO_597 (O_597,N_23626,N_23982);
or UO_598 (O_598,N_23557,N_22449);
nand UO_599 (O_599,N_22284,N_22016);
nand UO_600 (O_600,N_24305,N_23863);
nand UO_601 (O_601,N_24607,N_22354);
nor UO_602 (O_602,N_24043,N_23024);
nor UO_603 (O_603,N_22407,N_23272);
and UO_604 (O_604,N_22938,N_22446);
nor UO_605 (O_605,N_23339,N_23787);
and UO_606 (O_606,N_22157,N_22456);
or UO_607 (O_607,N_23081,N_24408);
nor UO_608 (O_608,N_24450,N_24509);
nand UO_609 (O_609,N_23153,N_23387);
xnor UO_610 (O_610,N_21936,N_23598);
xor UO_611 (O_611,N_22722,N_22728);
nand UO_612 (O_612,N_22035,N_23744);
nor UO_613 (O_613,N_24856,N_22375);
and UO_614 (O_614,N_23061,N_22068);
xnor UO_615 (O_615,N_22142,N_23507);
xnor UO_616 (O_616,N_23069,N_22617);
and UO_617 (O_617,N_23326,N_23812);
nand UO_618 (O_618,N_24501,N_24672);
and UO_619 (O_619,N_24248,N_23090);
xor UO_620 (O_620,N_22997,N_23151);
or UO_621 (O_621,N_23106,N_24316);
and UO_622 (O_622,N_22221,N_22031);
xor UO_623 (O_623,N_22010,N_22527);
or UO_624 (O_624,N_24844,N_23283);
and UO_625 (O_625,N_23126,N_22614);
and UO_626 (O_626,N_23260,N_24916);
nand UO_627 (O_627,N_23441,N_22461);
xnor UO_628 (O_628,N_24820,N_22654);
nand UO_629 (O_629,N_23913,N_24993);
xnor UO_630 (O_630,N_22958,N_22904);
and UO_631 (O_631,N_22758,N_21883);
xor UO_632 (O_632,N_24557,N_24508);
nand UO_633 (O_633,N_22854,N_22379);
or UO_634 (O_634,N_22964,N_22133);
and UO_635 (O_635,N_24399,N_23254);
nor UO_636 (O_636,N_22283,N_22540);
nor UO_637 (O_637,N_23592,N_23018);
and UO_638 (O_638,N_24974,N_23546);
or UO_639 (O_639,N_23013,N_24516);
and UO_640 (O_640,N_23072,N_24719);
xnor UO_641 (O_641,N_22092,N_24101);
or UO_642 (O_642,N_23607,N_23825);
xor UO_643 (O_643,N_22881,N_24765);
nor UO_644 (O_644,N_24850,N_23198);
nand UO_645 (O_645,N_23537,N_24189);
or UO_646 (O_646,N_21960,N_22506);
and UO_647 (O_647,N_24235,N_22640);
nor UO_648 (O_648,N_23577,N_23329);
nand UO_649 (O_649,N_24111,N_23181);
or UO_650 (O_650,N_24262,N_24282);
or UO_651 (O_651,N_22815,N_22012);
or UO_652 (O_652,N_23037,N_23456);
or UO_653 (O_653,N_22281,N_22956);
or UO_654 (O_654,N_24601,N_24329);
nor UO_655 (O_655,N_23981,N_23692);
xnor UO_656 (O_656,N_22632,N_24434);
nor UO_657 (O_657,N_24242,N_24968);
or UO_658 (O_658,N_24947,N_22009);
nor UO_659 (O_659,N_22602,N_23505);
and UO_660 (O_660,N_23745,N_24676);
xor UO_661 (O_661,N_23898,N_22886);
nor UO_662 (O_662,N_22033,N_22404);
nand UO_663 (O_663,N_23597,N_21983);
or UO_664 (O_664,N_21989,N_23855);
nor UO_665 (O_665,N_22996,N_22776);
xor UO_666 (O_666,N_23531,N_24980);
and UO_667 (O_667,N_24142,N_23498);
and UO_668 (O_668,N_24271,N_21956);
xor UO_669 (O_669,N_24519,N_24686);
nor UO_670 (O_670,N_22066,N_24959);
nand UO_671 (O_671,N_23178,N_24310);
and UO_672 (O_672,N_22030,N_22046);
or UO_673 (O_673,N_22555,N_22333);
nor UO_674 (O_674,N_23006,N_24706);
xor UO_675 (O_675,N_22567,N_23987);
and UO_676 (O_676,N_23664,N_23683);
nand UO_677 (O_677,N_23005,N_22749);
xnor UO_678 (O_678,N_24762,N_24503);
nor UO_679 (O_679,N_23475,N_22826);
and UO_680 (O_680,N_24078,N_24732);
nand UO_681 (O_681,N_21993,N_24889);
nor UO_682 (O_682,N_23363,N_23121);
and UO_683 (O_683,N_23185,N_22579);
nand UO_684 (O_684,N_22099,N_23651);
nand UO_685 (O_685,N_22768,N_24025);
xor UO_686 (O_686,N_22076,N_22362);
nor UO_687 (O_687,N_23261,N_22645);
or UO_688 (O_688,N_23601,N_23264);
and UO_689 (O_689,N_22755,N_23369);
and UO_690 (O_690,N_24749,N_23587);
xnor UO_691 (O_691,N_24384,N_24907);
or UO_692 (O_692,N_23646,N_22658);
or UO_693 (O_693,N_23341,N_24193);
or UO_694 (O_694,N_21961,N_24386);
nand UO_695 (O_695,N_22516,N_22780);
xnor UO_696 (O_696,N_24083,N_22235);
xor UO_697 (O_697,N_23814,N_22304);
xor UO_698 (O_698,N_24995,N_22253);
nand UO_699 (O_699,N_22804,N_23642);
nor UO_700 (O_700,N_24505,N_24188);
nor UO_701 (O_701,N_22919,N_22669);
or UO_702 (O_702,N_22606,N_22190);
nand UO_703 (O_703,N_24727,N_23606);
nor UO_704 (O_704,N_24483,N_21953);
or UO_705 (O_705,N_21972,N_24825);
and UO_706 (O_706,N_23575,N_22268);
nor UO_707 (O_707,N_24215,N_24651);
or UO_708 (O_708,N_22209,N_24425);
nor UO_709 (O_709,N_23386,N_22269);
xnor UO_710 (O_710,N_23394,N_23933);
nand UO_711 (O_711,N_24624,N_22601);
nor UO_712 (O_712,N_22969,N_24700);
or UO_713 (O_713,N_24494,N_24929);
nor UO_714 (O_714,N_22631,N_24966);
nand UO_715 (O_715,N_22757,N_24919);
and UO_716 (O_716,N_23707,N_23881);
xnor UO_717 (O_717,N_23749,N_23847);
nand UO_718 (O_718,N_23276,N_24454);
or UO_719 (O_719,N_22974,N_22249);
nor UO_720 (O_720,N_23921,N_24385);
and UO_721 (O_721,N_22307,N_23416);
xor UO_722 (O_722,N_24979,N_23571);
or UO_723 (O_723,N_22055,N_23802);
nor UO_724 (O_724,N_21881,N_23188);
xor UO_725 (O_725,N_22952,N_24658);
xnor UO_726 (O_726,N_24296,N_22902);
or UO_727 (O_727,N_24590,N_24126);
and UO_728 (O_728,N_22119,N_22387);
and UO_729 (O_729,N_24098,N_24069);
nand UO_730 (O_730,N_24643,N_24586);
xnor UO_731 (O_731,N_23438,N_23932);
nand UO_732 (O_732,N_24049,N_23688);
nand UO_733 (O_733,N_22618,N_23032);
or UO_734 (O_734,N_23663,N_24132);
xor UO_735 (O_735,N_23240,N_22990);
nor UO_736 (O_736,N_24089,N_24488);
nor UO_737 (O_737,N_23781,N_22707);
nor UO_738 (O_738,N_22921,N_21938);
xor UO_739 (O_739,N_22189,N_24238);
nor UO_740 (O_740,N_22788,N_23225);
and UO_741 (O_741,N_23396,N_23244);
or UO_742 (O_742,N_24729,N_22532);
and UO_743 (O_743,N_24863,N_24130);
and UO_744 (O_744,N_23808,N_23497);
and UO_745 (O_745,N_22943,N_23028);
xnor UO_746 (O_746,N_23521,N_23048);
and UO_747 (O_747,N_23845,N_23527);
nor UO_748 (O_748,N_22015,N_21912);
nor UO_749 (O_749,N_21971,N_24422);
or UO_750 (O_750,N_23030,N_22711);
nand UO_751 (O_751,N_22514,N_23422);
or UO_752 (O_752,N_22596,N_22070);
and UO_753 (O_753,N_23352,N_24457);
xor UO_754 (O_754,N_23654,N_23520);
or UO_755 (O_755,N_23804,N_22867);
and UO_756 (O_756,N_23672,N_24391);
and UO_757 (O_757,N_24797,N_23832);
and UO_758 (O_758,N_24920,N_23245);
nor UO_759 (O_759,N_23120,N_23886);
or UO_760 (O_760,N_23205,N_22723);
nor UO_761 (O_761,N_24020,N_21909);
xor UO_762 (O_762,N_24181,N_22107);
xnor UO_763 (O_763,N_22949,N_24994);
nand UO_764 (O_764,N_24013,N_22932);
nand UO_765 (O_765,N_22322,N_23885);
nand UO_766 (O_766,N_22869,N_22368);
xor UO_767 (O_767,N_23062,N_24908);
xor UO_768 (O_768,N_23333,N_24948);
xnor UO_769 (O_769,N_24213,N_24613);
nor UO_770 (O_770,N_23337,N_23695);
nand UO_771 (O_771,N_22915,N_24790);
and UO_772 (O_772,N_23722,N_24144);
nor UO_773 (O_773,N_23948,N_24622);
or UO_774 (O_774,N_21906,N_24938);
and UO_775 (O_775,N_23305,N_22609);
xor UO_776 (O_776,N_23294,N_22753);
or UO_777 (O_777,N_23612,N_24632);
xor UO_778 (O_778,N_23490,N_23914);
xnor UO_779 (O_779,N_23232,N_23901);
and UO_780 (O_780,N_24536,N_23485);
xor UO_781 (O_781,N_23738,N_22153);
nor UO_782 (O_782,N_23680,N_22819);
nand UO_783 (O_783,N_24093,N_23949);
or UO_784 (O_784,N_23954,N_22807);
nand UO_785 (O_785,N_22207,N_22953);
nand UO_786 (O_786,N_22895,N_23286);
and UO_787 (O_787,N_23137,N_22303);
and UO_788 (O_788,N_24348,N_22353);
nand UO_789 (O_789,N_24782,N_22525);
xnor UO_790 (O_790,N_22336,N_24197);
xor UO_791 (O_791,N_24818,N_22181);
or UO_792 (O_792,N_21939,N_22064);
nand UO_793 (O_793,N_23713,N_23161);
xnor UO_794 (O_794,N_23434,N_22835);
and UO_795 (O_795,N_22165,N_24308);
xor UO_796 (O_796,N_22234,N_24668);
and UO_797 (O_797,N_24116,N_21916);
nand UO_798 (O_798,N_22535,N_22937);
or UO_799 (O_799,N_24838,N_23536);
nor UO_800 (O_800,N_24639,N_22799);
nand UO_801 (O_801,N_23191,N_23755);
xor UO_802 (O_802,N_23986,N_24746);
nand UO_803 (O_803,N_22071,N_24027);
xnor UO_804 (O_804,N_24082,N_22829);
nor UO_805 (O_805,N_22174,N_23979);
or UO_806 (O_806,N_23556,N_22510);
or UO_807 (O_807,N_22260,N_23140);
xor UO_808 (O_808,N_23201,N_22536);
xor UO_809 (O_809,N_23474,N_23493);
or UO_810 (O_810,N_22732,N_22955);
xnor UO_811 (O_811,N_22057,N_22335);
nand UO_812 (O_812,N_23542,N_21887);
or UO_813 (O_813,N_24967,N_22164);
nor UO_814 (O_814,N_23446,N_23431);
nand UO_815 (O_815,N_23645,N_24652);
and UO_816 (O_816,N_23694,N_22752);
or UO_817 (O_817,N_24785,N_24670);
nand UO_818 (O_818,N_24005,N_24740);
nor UO_819 (O_819,N_24149,N_22634);
nand UO_820 (O_820,N_23991,N_24030);
or UO_821 (O_821,N_24636,N_23894);
nor UO_822 (O_822,N_24731,N_23532);
nor UO_823 (O_823,N_23959,N_23984);
nor UO_824 (O_824,N_23099,N_22331);
nand UO_825 (O_825,N_22496,N_22505);
nand UO_826 (O_826,N_24440,N_23833);
nor UO_827 (O_827,N_24009,N_22593);
and UO_828 (O_828,N_24524,N_21899);
and UO_829 (O_829,N_23082,N_22476);
or UO_830 (O_830,N_22295,N_24304);
and UO_831 (O_831,N_22885,N_23530);
nor UO_832 (O_832,N_22367,N_23231);
or UO_833 (O_833,N_22275,N_24045);
and UO_834 (O_834,N_24659,N_23603);
nor UO_835 (O_835,N_22355,N_23430);
or UO_836 (O_836,N_22492,N_21882);
xnor UO_837 (O_837,N_23031,N_23883);
or UO_838 (O_838,N_22451,N_22972);
nand UO_839 (O_839,N_22297,N_23750);
nor UO_840 (O_840,N_24848,N_24798);
or UO_841 (O_841,N_22685,N_24419);
nor UO_842 (O_842,N_22574,N_23934);
nor UO_843 (O_843,N_22515,N_24496);
xor UO_844 (O_844,N_23655,N_24062);
nand UO_845 (O_845,N_24955,N_22726);
xor UO_846 (O_846,N_22391,N_24141);
nand UO_847 (O_847,N_21978,N_23978);
and UO_848 (O_848,N_24255,N_22877);
or UO_849 (O_849,N_23842,N_23016);
or UO_850 (O_850,N_23234,N_23464);
nand UO_851 (O_851,N_23257,N_24245);
nand UO_852 (O_852,N_22638,N_23935);
nand UO_853 (O_853,N_24174,N_23827);
or UO_854 (O_854,N_24337,N_24459);
or UO_855 (O_855,N_23649,N_21991);
nand UO_856 (O_856,N_23402,N_23528);
nor UO_857 (O_857,N_22809,N_23599);
or UO_858 (O_858,N_23641,N_23743);
or UO_859 (O_859,N_22501,N_22531);
and UO_860 (O_860,N_24722,N_24338);
nor UO_861 (O_861,N_24480,N_22497);
nor UO_862 (O_862,N_24492,N_22657);
nand UO_863 (O_863,N_24808,N_24518);
nor UO_864 (O_864,N_24214,N_22178);
or UO_865 (O_865,N_21907,N_23053);
nor UO_866 (O_866,N_23334,N_23803);
and UO_867 (O_867,N_22152,N_23624);
or UO_868 (O_868,N_24145,N_24136);
xor UO_869 (O_869,N_23211,N_24368);
nor UO_870 (O_870,N_22381,N_24667);
nor UO_871 (O_871,N_23321,N_23323);
xor UO_872 (O_872,N_23290,N_24138);
nor UO_873 (O_873,N_22242,N_22806);
and UO_874 (O_874,N_24133,N_22939);
nand UO_875 (O_875,N_22038,N_24733);
xnor UO_876 (O_876,N_23214,N_23809);
xnor UO_877 (O_877,N_22498,N_23132);
and UO_878 (O_878,N_22907,N_24989);
and UO_879 (O_879,N_24807,N_24034);
xor UO_880 (O_880,N_22059,N_24266);
or UO_881 (O_881,N_22528,N_24812);
xnor UO_882 (O_882,N_21981,N_23307);
and UO_883 (O_883,N_24611,N_22156);
xnor UO_884 (O_884,N_23226,N_23451);
or UO_885 (O_885,N_23378,N_22212);
nor UO_886 (O_886,N_23288,N_23036);
or UO_887 (O_887,N_22950,N_23839);
xnor UO_888 (O_888,N_23544,N_24540);
nor UO_889 (O_889,N_22673,N_22306);
nand UO_890 (O_890,N_23176,N_22978);
or UO_891 (O_891,N_22513,N_22419);
or UO_892 (O_892,N_22225,N_22223);
nand UO_893 (O_893,N_23298,N_22517);
nand UO_894 (O_894,N_23131,N_22197);
nand UO_895 (O_895,N_24757,N_22380);
nand UO_896 (O_896,N_22800,N_21997);
and UO_897 (O_897,N_24151,N_24463);
or UO_898 (O_898,N_22647,N_22765);
and UO_899 (O_899,N_22173,N_24108);
or UO_900 (O_900,N_22377,N_22625);
nand UO_901 (O_901,N_24687,N_24548);
nand UO_902 (O_902,N_21967,N_22310);
nor UO_903 (O_903,N_24620,N_22250);
nand UO_904 (O_904,N_24124,N_22191);
or UO_905 (O_905,N_24075,N_22888);
nand UO_906 (O_906,N_23239,N_22125);
or UO_907 (O_907,N_23824,N_22315);
and UO_908 (O_908,N_23547,N_24899);
and UO_909 (O_909,N_24939,N_23936);
nor UO_910 (O_910,N_24499,N_24285);
xor UO_911 (O_911,N_22028,N_24745);
and UO_912 (O_912,N_23057,N_24110);
nor UO_913 (O_913,N_23467,N_24743);
or UO_914 (O_914,N_23492,N_22141);
and UO_915 (O_915,N_24663,N_21925);
nor UO_916 (O_916,N_24893,N_24533);
or UO_917 (O_917,N_22296,N_24250);
xor UO_918 (O_918,N_24896,N_22120);
or UO_919 (O_919,N_24690,N_23524);
nand UO_920 (O_920,N_22935,N_23453);
or UO_921 (O_921,N_23627,N_22422);
or UO_922 (O_922,N_22452,N_22183);
and UO_923 (O_923,N_24489,N_22805);
xnor UO_924 (O_924,N_23909,N_22842);
and UO_925 (O_925,N_22412,N_21952);
xnor UO_926 (O_926,N_23034,N_24010);
and UO_927 (O_927,N_22264,N_23130);
and UO_928 (O_928,N_22286,N_23335);
and UO_929 (O_929,N_24950,N_21918);
xor UO_930 (O_930,N_22434,N_21889);
and UO_931 (O_931,N_22784,N_22760);
or UO_932 (O_932,N_24388,N_22639);
and UO_933 (O_933,N_22424,N_24764);
nor UO_934 (O_934,N_23253,N_23342);
xor UO_935 (O_935,N_22546,N_24675);
or UO_936 (O_936,N_22859,N_22980);
xor UO_937 (O_937,N_23494,N_22820);
and UO_938 (O_938,N_23862,N_23628);
xor UO_939 (O_939,N_22664,N_23776);
nand UO_940 (O_940,N_22624,N_21901);
nor UO_941 (O_941,N_23349,N_23094);
nand UO_942 (O_942,N_24350,N_24406);
nor UO_943 (O_943,N_23092,N_24065);
nand UO_944 (O_944,N_23770,N_23566);
xnor UO_945 (O_945,N_24556,N_23455);
nor UO_946 (O_946,N_23529,N_22693);
or UO_947 (O_947,N_22232,N_23317);
xor UO_948 (O_948,N_24952,N_24559);
xnor UO_949 (O_949,N_22740,N_22328);
and UO_950 (O_950,N_22447,N_24612);
xnor UO_951 (O_951,N_23699,N_22227);
or UO_952 (O_952,N_23419,N_24958);
xnor UO_953 (O_953,N_24597,N_22705);
xnor UO_954 (O_954,N_24904,N_22203);
nor UO_955 (O_955,N_23702,N_22942);
xnor UO_956 (O_956,N_22118,N_21905);
nor UO_957 (O_957,N_23910,N_24365);
and UO_958 (O_958,N_21955,N_23461);
nand UO_959 (O_959,N_24318,N_22045);
nand UO_960 (O_960,N_24726,N_22054);
and UO_961 (O_961,N_23397,N_24682);
or UO_962 (O_962,N_23340,N_22166);
nor UO_963 (O_963,N_22104,N_23952);
xnor UO_964 (O_964,N_22431,N_21943);
and UO_965 (O_965,N_24859,N_23356);
nor UO_966 (O_966,N_22970,N_22872);
nand UO_967 (O_967,N_24852,N_23209);
xor UO_968 (O_968,N_23675,N_22703);
nor UO_969 (O_969,N_24629,N_24917);
xnor UO_970 (O_970,N_22148,N_22037);
nand UO_971 (O_971,N_23207,N_23008);
or UO_972 (O_972,N_24153,N_22294);
and UO_973 (O_973,N_22003,N_23197);
xor UO_974 (O_974,N_23347,N_23693);
nand UO_975 (O_975,N_22718,N_24497);
or UO_976 (O_976,N_23753,N_24292);
nor UO_977 (O_977,N_24072,N_24294);
nand UO_978 (O_978,N_24263,N_22841);
and UO_979 (O_979,N_24380,N_22947);
xnor UO_980 (O_980,N_22041,N_24180);
xnor UO_981 (O_981,N_22453,N_23133);
and UO_982 (O_982,N_23332,N_22607);
nand UO_983 (O_983,N_24366,N_22600);
xnor UO_984 (O_984,N_23747,N_22075);
nor UO_985 (O_985,N_21950,N_24752);
and UO_986 (O_986,N_24600,N_21998);
xnor UO_987 (O_987,N_23629,N_23795);
and UO_988 (O_988,N_22411,N_23141);
nand UO_989 (O_989,N_22474,N_23501);
nand UO_990 (O_990,N_24641,N_24648);
or UO_991 (O_991,N_24354,N_24204);
and UO_992 (O_992,N_22667,N_22585);
nor UO_993 (O_993,N_24200,N_22405);
xor UO_994 (O_994,N_22457,N_22111);
and UO_995 (O_995,N_22659,N_22537);
and UO_996 (O_996,N_22093,N_23965);
nor UO_997 (O_997,N_22748,N_22050);
xnor UO_998 (O_998,N_23679,N_23405);
and UO_999 (O_999,N_22580,N_24647);
xor UO_1000 (O_1000,N_24954,N_22077);
nor UO_1001 (O_1001,N_23564,N_22482);
nor UO_1002 (O_1002,N_22500,N_23942);
and UO_1003 (O_1003,N_24353,N_24625);
xor UO_1004 (O_1004,N_23331,N_22013);
or UO_1005 (O_1005,N_22472,N_24279);
xor UO_1006 (O_1006,N_23482,N_23669);
xnor UO_1007 (O_1007,N_24877,N_23473);
xor UO_1008 (O_1008,N_24340,N_24349);
nor UO_1009 (O_1009,N_23499,N_24206);
nand UO_1010 (O_1010,N_22481,N_22559);
xor UO_1011 (O_1011,N_24795,N_24569);
or UO_1012 (O_1012,N_24077,N_23395);
nand UO_1013 (O_1013,N_22882,N_22913);
nor UO_1014 (O_1014,N_21902,N_23113);
and UO_1015 (O_1015,N_23206,N_23407);
xor UO_1016 (O_1016,N_22665,N_24606);
xnor UO_1017 (O_1017,N_23915,N_24554);
nor UO_1018 (O_1018,N_22598,N_23570);
nor UO_1019 (O_1019,N_22876,N_22605);
nor UO_1020 (O_1020,N_24357,N_24846);
xnor UO_1021 (O_1021,N_24960,N_23820);
nand UO_1022 (O_1022,N_22706,N_22180);
nand UO_1023 (O_1023,N_24217,N_23851);
nor UO_1024 (O_1024,N_23892,N_24220);
or UO_1025 (O_1025,N_24328,N_24999);
nand UO_1026 (O_1026,N_22408,N_24665);
nor UO_1027 (O_1027,N_23216,N_22376);
nor UO_1028 (O_1028,N_24413,N_24178);
nor UO_1029 (O_1029,N_22369,N_23250);
xnor UO_1030 (O_1030,N_24302,N_23733);
nor UO_1031 (O_1031,N_23444,N_22021);
or UO_1032 (O_1032,N_23604,N_24562);
xnor UO_1033 (O_1033,N_22272,N_22966);
and UO_1034 (O_1034,N_24280,N_23388);
and UO_1035 (O_1035,N_22298,N_24935);
or UO_1036 (O_1036,N_22672,N_22889);
and UO_1037 (O_1037,N_22135,N_22345);
or UO_1038 (O_1038,N_22334,N_24549);
or UO_1039 (O_1039,N_23022,N_24039);
xnor UO_1040 (O_1040,N_23366,N_22238);
or UO_1041 (O_1041,N_23690,N_23412);
or UO_1042 (O_1042,N_23476,N_23466);
nor UO_1043 (O_1043,N_24526,N_23401);
xor UO_1044 (O_1044,N_24187,N_22371);
nand UO_1045 (O_1045,N_23899,N_22763);
or UO_1046 (O_1046,N_24427,N_24890);
and UO_1047 (O_1047,N_24654,N_23746);
nor UO_1048 (O_1048,N_22036,N_23539);
and UO_1049 (O_1049,N_23995,N_22626);
xor UO_1050 (O_1050,N_24905,N_23596);
xnor UO_1051 (O_1051,N_24602,N_23270);
xor UO_1052 (O_1052,N_23817,N_23448);
nor UO_1053 (O_1053,N_23620,N_24362);
and UO_1054 (O_1054,N_21932,N_23518);
nor UO_1055 (O_1055,N_23312,N_24819);
nand UO_1056 (O_1056,N_23788,N_24092);
nand UO_1057 (O_1057,N_22266,N_23858);
xor UO_1058 (O_1058,N_23119,N_23972);
xor UO_1059 (O_1059,N_24059,N_23384);
xor UO_1060 (O_1060,N_23840,N_22637);
nand UO_1061 (O_1061,N_23777,N_23436);
nor UO_1062 (O_1062,N_22073,N_22056);
and UO_1063 (O_1063,N_22374,N_23242);
nand UO_1064 (O_1064,N_22263,N_22565);
and UO_1065 (O_1065,N_24874,N_22836);
and UO_1066 (O_1066,N_23698,N_22291);
nor UO_1067 (O_1067,N_23767,N_23673);
or UO_1068 (O_1068,N_22977,N_21924);
nand UO_1069 (O_1069,N_24539,N_24684);
xor UO_1070 (O_1070,N_23721,N_23908);
and UO_1071 (O_1071,N_22911,N_23511);
nand UO_1072 (O_1072,N_24453,N_24231);
and UO_1073 (O_1073,N_23994,N_24840);
nand UO_1074 (O_1074,N_23114,N_24363);
nor UO_1075 (O_1075,N_22556,N_22689);
nor UO_1076 (O_1076,N_23506,N_22548);
nand UO_1077 (O_1077,N_22459,N_21878);
and UO_1078 (O_1078,N_24205,N_24066);
nor UO_1079 (O_1079,N_23510,N_22350);
nand UO_1080 (O_1080,N_23593,N_23677);
or UO_1081 (O_1081,N_21985,N_23790);
nand UO_1082 (O_1082,N_24322,N_22276);
nor UO_1083 (O_1083,N_24369,N_22746);
or UO_1084 (O_1084,N_24692,N_24071);
and UO_1085 (O_1085,N_23923,N_23983);
nor UO_1086 (O_1086,N_21964,N_24901);
nand UO_1087 (O_1087,N_22072,N_23928);
nor UO_1088 (O_1088,N_24361,N_23763);
xor UO_1089 (O_1089,N_22965,N_24978);
xnor UO_1090 (O_1090,N_22065,N_22047);
xnor UO_1091 (O_1091,N_24854,N_22116);
and UO_1092 (O_1092,N_24801,N_22458);
nand UO_1093 (O_1093,N_24836,N_22087);
or UO_1094 (O_1094,N_21921,N_22611);
xor UO_1095 (O_1095,N_23343,N_23315);
xnor UO_1096 (O_1096,N_22103,N_22138);
nand UO_1097 (O_1097,N_22236,N_24644);
nor UO_1098 (O_1098,N_24866,N_23470);
or UO_1099 (O_1099,N_22194,N_24323);
or UO_1100 (O_1100,N_23676,N_21884);
or UO_1101 (O_1101,N_22862,N_24793);
or UO_1102 (O_1102,N_22831,N_22244);
nor UO_1103 (O_1103,N_24286,N_23635);
or UO_1104 (O_1104,N_22427,N_22948);
nand UO_1105 (O_1105,N_21958,N_22553);
and UO_1106 (O_1106,N_23950,N_22326);
or UO_1107 (O_1107,N_24965,N_24128);
or UO_1108 (O_1108,N_23469,N_23815);
nand UO_1109 (O_1109,N_22900,N_23381);
or UO_1110 (O_1110,N_22993,N_24297);
xor UO_1111 (O_1111,N_22246,N_24906);
nor UO_1112 (O_1112,N_22756,N_24246);
or UO_1113 (O_1113,N_21982,N_24758);
and UO_1114 (O_1114,N_22237,N_24439);
and UO_1115 (O_1115,N_23930,N_22265);
xor UO_1116 (O_1116,N_24504,N_24914);
xnor UO_1117 (O_1117,N_23517,N_24376);
and UO_1118 (O_1118,N_22883,N_22084);
and UO_1119 (O_1119,N_23658,N_24756);
or UO_1120 (O_1120,N_21891,N_23784);
and UO_1121 (O_1121,N_23889,N_22973);
nand UO_1122 (O_1122,N_23432,N_22096);
and UO_1123 (O_1123,N_23582,N_22085);
and UO_1124 (O_1124,N_22991,N_22934);
and UO_1125 (O_1125,N_22686,N_23890);
xor UO_1126 (O_1126,N_23300,N_24715);
nor UO_1127 (O_1127,N_24617,N_22649);
or UO_1128 (O_1128,N_23585,N_21893);
nor UO_1129 (O_1129,N_22083,N_22019);
nor UO_1130 (O_1130,N_23541,N_23009);
nor UO_1131 (O_1131,N_21986,N_22144);
xor UO_1132 (O_1132,N_23111,N_24736);
and UO_1133 (O_1133,N_23112,N_24609);
nor UO_1134 (O_1134,N_24035,N_22455);
and UO_1135 (O_1135,N_24152,N_24544);
and UO_1136 (O_1136,N_23793,N_22150);
or UO_1137 (O_1137,N_24410,N_24956);
nor UO_1138 (O_1138,N_24791,N_22441);
xor UO_1139 (O_1139,N_23632,N_24154);
nor UO_1140 (O_1140,N_24073,N_22681);
nand UO_1141 (O_1141,N_23399,N_23997);
xor UO_1142 (O_1142,N_24051,N_22323);
xor UO_1143 (O_1143,N_24694,N_24022);
and UO_1144 (O_1144,N_24876,N_24249);
xnor UO_1145 (O_1145,N_23463,N_22483);
nor UO_1146 (O_1146,N_21942,N_21990);
xor UO_1147 (O_1147,N_22468,N_23351);
nand UO_1148 (O_1148,N_22766,N_23659);
xnor UO_1149 (O_1149,N_23259,N_22670);
nor UO_1150 (O_1150,N_23773,N_24708);
nor UO_1151 (O_1151,N_24638,N_22110);
xor UO_1152 (O_1152,N_24162,N_22435);
nor UO_1153 (O_1153,N_22445,N_23135);
nand UO_1154 (O_1154,N_24054,N_24873);
and UO_1155 (O_1155,N_23964,N_22105);
nor UO_1156 (O_1156,N_24445,N_23956);
nor UO_1157 (O_1157,N_23670,N_22504);
and UO_1158 (O_1158,N_23800,N_23045);
or UO_1159 (O_1159,N_22154,N_23801);
nor UO_1160 (O_1160,N_23275,N_22621);
and UO_1161 (O_1161,N_23160,N_22905);
nor UO_1162 (O_1162,N_22694,N_23559);
and UO_1163 (O_1163,N_22720,N_23525);
and UO_1164 (O_1164,N_21937,N_24253);
nor UO_1165 (O_1165,N_22279,N_22395);
xor UO_1166 (O_1166,N_23088,N_24240);
and UO_1167 (O_1167,N_22478,N_22430);
and UO_1168 (O_1168,N_23711,N_22175);
and UO_1169 (O_1169,N_22584,N_21973);
nor UO_1170 (O_1170,N_22043,N_24969);
and UO_1171 (O_1171,N_24640,N_22604);
xnor UO_1172 (O_1172,N_23625,N_23853);
nand UO_1173 (O_1173,N_21880,N_24871);
and UO_1174 (O_1174,N_22179,N_23076);
and UO_1175 (O_1175,N_24777,N_23297);
or UO_1176 (O_1176,N_23358,N_23865);
nor UO_1177 (O_1177,N_24090,N_24177);
and UO_1178 (O_1178,N_23344,N_23289);
nand UO_1179 (O_1179,N_22688,N_24428);
nand UO_1180 (O_1180,N_23318,N_24171);
nor UO_1181 (O_1181,N_23685,N_21976);
or UO_1182 (O_1182,N_22998,N_23105);
and UO_1183 (O_1183,N_24387,N_23882);
and UO_1184 (O_1184,N_24229,N_23854);
xnor UO_1185 (O_1185,N_22751,N_21896);
nand UO_1186 (O_1186,N_23314,N_24169);
nor UO_1187 (O_1187,N_22946,N_22413);
nor UO_1188 (O_1188,N_24320,N_22024);
and UO_1189 (O_1189,N_24314,N_23170);
and UO_1190 (O_1190,N_22785,N_21914);
and UO_1191 (O_1191,N_23000,N_22519);
nor UO_1192 (O_1192,N_23522,N_24403);
nor UO_1193 (O_1193,N_24655,N_22587);
or UO_1194 (O_1194,N_22161,N_23503);
nand UO_1195 (O_1195,N_22477,N_23550);
nand UO_1196 (O_1196,N_22918,N_22662);
xor UO_1197 (O_1197,N_24913,N_24531);
and UO_1198 (O_1198,N_24086,N_22920);
nor UO_1199 (O_1199,N_23278,N_23054);
xor UO_1200 (O_1200,N_22088,N_24203);
nand UO_1201 (O_1201,N_23684,N_22484);
nand UO_1202 (O_1202,N_24951,N_23179);
xnor UO_1203 (O_1203,N_21947,N_24411);
nor UO_1204 (O_1204,N_24595,N_24909);
xor UO_1205 (O_1205,N_23293,N_22710);
or UO_1206 (O_1206,N_24750,N_23766);
xnor UO_1207 (O_1207,N_23007,N_24196);
and UO_1208 (O_1208,N_22359,N_22469);
xor UO_1209 (O_1209,N_24448,N_23063);
and UO_1210 (O_1210,N_23087,N_22466);
nor UO_1211 (O_1211,N_24547,N_23047);
or UO_1212 (O_1212,N_22890,N_23067);
nor UO_1213 (O_1213,N_23608,N_23439);
nand UO_1214 (O_1214,N_23302,N_23204);
xor UO_1215 (O_1215,N_22029,N_24301);
xor UO_1216 (O_1216,N_22415,N_22739);
nand UO_1217 (O_1217,N_24579,N_24657);
nand UO_1218 (O_1218,N_23741,N_22398);
or UO_1219 (O_1219,N_23875,N_22192);
xnor UO_1220 (O_1220,N_23805,N_23425);
xor UO_1221 (O_1221,N_23783,N_23643);
and UO_1222 (O_1222,N_23966,N_24572);
nand UO_1223 (O_1223,N_24776,N_24593);
and UO_1224 (O_1224,N_24589,N_22927);
and UO_1225 (O_1225,N_22735,N_23567);
nor UO_1226 (O_1226,N_23228,N_22814);
nand UO_1227 (O_1227,N_22316,N_23241);
nor UO_1228 (O_1228,N_23573,N_21979);
or UO_1229 (O_1229,N_24107,N_23462);
nand UO_1230 (O_1230,N_23172,N_22810);
nand UO_1231 (O_1231,N_24330,N_24861);
nand UO_1232 (O_1232,N_22933,N_22392);
nor UO_1233 (O_1233,N_23107,N_23562);
or UO_1234 (O_1234,N_24345,N_22261);
or UO_1235 (O_1235,N_23975,N_23703);
xor UO_1236 (O_1236,N_23263,N_23079);
and UO_1237 (O_1237,N_23504,N_22309);
and UO_1238 (O_1238,N_22724,N_23350);
nand UO_1239 (O_1239,N_24198,N_22573);
or UO_1240 (O_1240,N_24288,N_23543);
nor UO_1241 (O_1241,N_23391,N_23969);
or UO_1242 (O_1242,N_22916,N_24944);
or UO_1243 (O_1243,N_24159,N_24436);
xor UO_1244 (O_1244,N_23168,N_24867);
nand UO_1245 (O_1245,N_23761,N_21954);
or UO_1246 (O_1246,N_23900,N_24574);
xor UO_1247 (O_1247,N_23696,N_23623);
xnor UO_1248 (O_1248,N_23811,N_23799);
nor UO_1249 (O_1249,N_23602,N_23631);
xnor UO_1250 (O_1250,N_23406,N_22668);
nor UO_1251 (O_1251,N_22692,N_22420);
or UO_1252 (O_1252,N_22801,N_24097);
xor UO_1253 (O_1253,N_24112,N_24705);
and UO_1254 (O_1254,N_24482,N_23267);
or UO_1255 (O_1255,N_24529,N_24839);
and UO_1256 (O_1256,N_24763,N_23477);
or UO_1257 (O_1257,N_24099,N_23584);
nor UO_1258 (O_1258,N_23051,N_24561);
and UO_1259 (O_1259,N_24747,N_22591);
and UO_1260 (O_1260,N_23906,N_24462);
nor UO_1261 (O_1261,N_23879,N_22773);
and UO_1262 (O_1262,N_23712,N_24831);
and UO_1263 (O_1263,N_22554,N_23600);
nand UO_1264 (O_1264,N_21879,N_23791);
nand UO_1265 (O_1265,N_23382,N_22564);
nand UO_1266 (O_1266,N_22005,N_23779);
xnor UO_1267 (O_1267,N_22712,N_23968);
or UO_1268 (O_1268,N_23010,N_23648);
nand UO_1269 (O_1269,N_23852,N_23737);
nor UO_1270 (O_1270,N_23734,N_22898);
xor UO_1271 (O_1271,N_21995,N_24401);
nor UO_1272 (O_1272,N_22027,N_22488);
nor UO_1273 (O_1273,N_22464,N_22853);
or UO_1274 (O_1274,N_24184,N_24534);
nand UO_1275 (O_1275,N_24456,N_24332);
nand UO_1276 (O_1276,N_22572,N_22273);
xor UO_1277 (O_1277,N_24102,N_24147);
nor UO_1278 (O_1278,N_24236,N_23856);
and UO_1279 (O_1279,N_22589,N_24717);
and UO_1280 (O_1280,N_22880,N_24256);
xnor UO_1281 (O_1281,N_24618,N_24513);
xnor UO_1282 (O_1282,N_23233,N_22743);
nand UO_1283 (O_1283,N_24451,N_24277);
or UO_1284 (O_1284,N_23724,N_22243);
nand UO_1285 (O_1285,N_23281,N_24381);
xnor UO_1286 (O_1286,N_22454,N_23478);
nand UO_1287 (O_1287,N_22592,N_22641);
nor UO_1288 (O_1288,N_24608,N_24164);
and UO_1289 (O_1289,N_22069,N_22259);
nand UO_1290 (O_1290,N_23850,N_22642);
xnor UO_1291 (O_1291,N_23985,N_22736);
xnor UO_1292 (O_1292,N_24257,N_23322);
and UO_1293 (O_1293,N_24321,N_22837);
or UO_1294 (O_1294,N_21994,N_24029);
nor UO_1295 (O_1295,N_24334,N_22608);
nor UO_1296 (O_1296,N_23073,N_23359);
or UO_1297 (O_1297,N_22339,N_24123);
nand UO_1298 (O_1298,N_22491,N_24324);
nor UO_1299 (O_1299,N_23609,N_22568);
and UO_1300 (O_1300,N_24221,N_22204);
nor UO_1301 (O_1301,N_23999,N_22599);
xnor UO_1302 (O_1302,N_23035,N_22581);
nor UO_1303 (O_1303,N_24616,N_24394);
or UO_1304 (O_1304,N_24832,N_23656);
nor UO_1305 (O_1305,N_23971,N_24982);
nor UO_1306 (O_1306,N_23320,N_22790);
nor UO_1307 (O_1307,N_22894,N_22356);
xor UO_1308 (O_1308,N_23220,N_24259);
and UO_1309 (O_1309,N_23495,N_23810);
nor UO_1310 (O_1310,N_24079,N_22983);
nor UO_1311 (O_1311,N_23380,N_22081);
or UO_1312 (O_1312,N_24176,N_23822);
and UO_1313 (O_1313,N_23704,N_24418);
and UO_1314 (O_1314,N_22816,N_24834);
nor UO_1315 (O_1315,N_24068,N_24094);
nand UO_1316 (O_1316,N_24576,N_24634);
or UO_1317 (O_1317,N_23377,N_23946);
xnor UO_1318 (O_1318,N_23605,N_21980);
nand UO_1319 (O_1319,N_24167,N_23059);
nand UO_1320 (O_1320,N_24817,N_24707);
and UO_1321 (O_1321,N_22691,N_23535);
or UO_1322 (O_1322,N_24645,N_23075);
nand UO_1323 (O_1323,N_22171,N_23429);
xor UO_1324 (O_1324,N_24813,N_22330);
or UO_1325 (O_1325,N_24070,N_22302);
nor UO_1326 (O_1326,N_24370,N_24696);
xnor UO_1327 (O_1327,N_24541,N_22959);
and UO_1328 (O_1328,N_24773,N_22864);
xor UO_1329 (O_1329,N_24771,N_22873);
nor UO_1330 (O_1330,N_23143,N_23136);
nand UO_1331 (O_1331,N_22373,N_24930);
nand UO_1332 (O_1332,N_22569,N_24603);
nand UO_1333 (O_1333,N_22813,N_23287);
and UO_1334 (O_1334,N_22365,N_22170);
nand UO_1335 (O_1335,N_23723,N_23039);
or UO_1336 (O_1336,N_23681,N_22508);
and UO_1337 (O_1337,N_22473,N_23479);
or UO_1338 (O_1338,N_22791,N_22199);
nor UO_1339 (O_1339,N_24847,N_24977);
and UO_1340 (O_1340,N_24467,N_23404);
and UO_1341 (O_1341,N_24992,N_23594);
nand UO_1342 (O_1342,N_23427,N_24535);
nor UO_1343 (O_1343,N_22737,N_23752);
xor UO_1344 (O_1344,N_22960,N_22410);
or UO_1345 (O_1345,N_24637,N_23595);
or UO_1346 (O_1346,N_23077,N_23891);
nor UO_1347 (O_1347,N_21984,N_22849);
nand UO_1348 (O_1348,N_22787,N_24653);
nand UO_1349 (O_1349,N_23893,N_22733);
xnor UO_1350 (O_1350,N_22619,N_22226);
and UO_1351 (O_1351,N_23192,N_22040);
and UO_1352 (O_1352,N_24991,N_22329);
and UO_1353 (O_1353,N_22995,N_21969);
and UO_1354 (O_1354,N_24414,N_22487);
xor UO_1355 (O_1355,N_24478,N_21944);
xnor UO_1356 (O_1356,N_23144,N_24805);
nor UO_1357 (O_1357,N_23714,N_24183);
and UO_1358 (O_1358,N_24432,N_22219);
xnor UO_1359 (O_1359,N_24990,N_24841);
nand UO_1360 (O_1360,N_23345,N_23026);
nor UO_1361 (O_1361,N_24076,N_24725);
or UO_1362 (O_1362,N_24975,N_23674);
or UO_1363 (O_1363,N_23630,N_24794);
nand UO_1364 (O_1364,N_23481,N_22358);
nor UO_1365 (O_1365,N_23717,N_23458);
nand UO_1366 (O_1366,N_23078,N_22696);
and UO_1367 (O_1367,N_24584,N_21977);
or UO_1368 (O_1368,N_23516,N_24937);
nor UO_1369 (O_1369,N_23774,N_24986);
and UO_1370 (O_1370,N_24779,N_23070);
xor UO_1371 (O_1371,N_23058,N_23265);
and UO_1372 (O_1372,N_23740,N_24796);
xnor UO_1373 (O_1373,N_24378,N_22443);
and UO_1374 (O_1374,N_22709,N_23164);
or UO_1375 (O_1375,N_22139,N_24738);
xor UO_1376 (O_1376,N_23869,N_23103);
xor UO_1377 (O_1377,N_23640,N_21903);
nand UO_1378 (O_1378,N_23868,N_24767);
and UO_1379 (O_1379,N_24417,N_23538);
nand UO_1380 (O_1380,N_22987,N_22131);
and UO_1381 (O_1381,N_23152,N_22288);
or UO_1382 (O_1382,N_23647,N_22612);
nand UO_1383 (O_1383,N_24117,N_22899);
or UO_1384 (O_1384,N_24398,N_24984);
xnor UO_1385 (O_1385,N_22671,N_23924);
nor UO_1386 (O_1386,N_24383,N_22762);
or UO_1387 (O_1387,N_24910,N_22557);
or UO_1388 (O_1388,N_24849,N_22558);
nor UO_1389 (O_1389,N_22715,N_24809);
or UO_1390 (O_1390,N_23836,N_21975);
nand UO_1391 (O_1391,N_23848,N_23806);
or UO_1392 (O_1392,N_24507,N_24109);
nor UO_1393 (O_1393,N_24000,N_23502);
xnor UO_1394 (O_1394,N_21934,N_24008);
xnor UO_1395 (O_1395,N_23148,N_22346);
nor UO_1396 (O_1396,N_22417,N_22450);
nand UO_1397 (O_1397,N_22610,N_22494);
xnor UO_1398 (O_1398,N_23616,N_23735);
nor UO_1399 (O_1399,N_24822,N_22163);
nor UO_1400 (O_1400,N_24711,N_23754);
nand UO_1401 (O_1401,N_24564,N_22547);
and UO_1402 (O_1402,N_24037,N_22968);
nor UO_1403 (O_1403,N_22502,N_24433);
and UO_1404 (O_1404,N_23308,N_22909);
xor UO_1405 (O_1405,N_24799,N_24416);
or UO_1406 (O_1406,N_22847,N_22674);
nor UO_1407 (O_1407,N_22550,N_24963);
or UO_1408 (O_1408,N_24781,N_24942);
nand UO_1409 (O_1409,N_22258,N_23835);
or UO_1410 (O_1410,N_21927,N_24699);
xnor UO_1411 (O_1411,N_23229,N_24976);
nand UO_1412 (O_1412,N_24845,N_24119);
and UO_1413 (O_1413,N_22562,N_22999);
or UO_1414 (O_1414,N_24298,N_24649);
xnor UO_1415 (O_1415,N_22666,N_22078);
or UO_1416 (O_1416,N_22280,N_22127);
and UO_1417 (O_1417,N_22675,N_23365);
nor UO_1418 (O_1418,N_22929,N_21996);
nor UO_1419 (O_1419,N_23960,N_24596);
nor UO_1420 (O_1420,N_23519,N_24396);
xor UO_1421 (O_1421,N_23223,N_23870);
and UO_1422 (O_1422,N_24303,N_24283);
nor UO_1423 (O_1423,N_23150,N_23489);
nor UO_1424 (O_1424,N_23922,N_23551);
nor UO_1425 (O_1425,N_24252,N_23064);
and UO_1426 (O_1426,N_23996,N_22112);
nand UO_1427 (O_1427,N_24789,N_23389);
nor UO_1428 (O_1428,N_23095,N_24703);
nand UO_1429 (O_1429,N_24442,N_23149);
nor UO_1430 (O_1430,N_22349,N_24555);
nor UO_1431 (O_1431,N_24465,N_22789);
nor UO_1432 (O_1432,N_24515,N_22544);
xor UO_1433 (O_1433,N_24415,N_24855);
nor UO_1434 (O_1434,N_22750,N_24295);
and UO_1435 (O_1435,N_22177,N_24233);
and UO_1436 (O_1436,N_22414,N_22852);
nand UO_1437 (O_1437,N_23459,N_24335);
and UO_1438 (O_1438,N_23667,N_24875);
nor UO_1439 (O_1439,N_22145,N_23831);
nor UO_1440 (O_1440,N_23291,N_23015);
xnor UO_1441 (O_1441,N_22677,N_23917);
xor UO_1442 (O_1442,N_24026,N_23826);
or UO_1443 (O_1443,N_24563,N_23043);
and UO_1444 (O_1444,N_22124,N_24816);
xor UO_1445 (O_1445,N_24053,N_21970);
and UO_1446 (O_1446,N_22499,N_22811);
nor UO_1447 (O_1447,N_24530,N_22287);
and UO_1448 (O_1448,N_22343,N_22290);
nand UO_1449 (O_1449,N_23872,N_23483);
xor UO_1450 (O_1450,N_22108,N_22020);
xor UO_1451 (O_1451,N_24646,N_24042);
nand UO_1452 (O_1452,N_24753,N_23418);
or UO_1453 (O_1453,N_23572,N_22745);
xor UO_1454 (O_1454,N_22406,N_23579);
xor UO_1455 (O_1455,N_23687,N_23668);
nor UO_1456 (O_1456,N_22971,N_22239);
and UO_1457 (O_1457,N_24580,N_22764);
and UO_1458 (O_1458,N_23748,N_24351);
and UO_1459 (O_1459,N_24983,N_24677);
or UO_1460 (O_1460,N_24802,N_23373);
nand UO_1461 (O_1461,N_22100,N_22779);
nor UO_1462 (O_1462,N_23591,N_22292);
nand UO_1463 (O_1463,N_24317,N_24824);
nor UO_1464 (O_1464,N_23415,N_22448);
or UO_1465 (O_1465,N_22403,N_24621);
nand UO_1466 (O_1466,N_24040,N_22382);
or UO_1467 (O_1467,N_23947,N_22211);
or UO_1468 (O_1468,N_22534,N_24364);
and UO_1469 (O_1469,N_24662,N_24003);
xnor UO_1470 (O_1470,N_24605,N_23849);
nand UO_1471 (O_1471,N_23056,N_24592);
or UO_1472 (O_1472,N_22742,N_23653);
and UO_1473 (O_1473,N_24289,N_24814);
or UO_1474 (O_1474,N_23139,N_24768);
or UO_1475 (O_1475,N_22759,N_24140);
xor UO_1476 (O_1476,N_21929,N_21941);
and UO_1477 (O_1477,N_23100,N_22143);
nor UO_1478 (O_1478,N_23963,N_24829);
or UO_1479 (O_1479,N_24211,N_23729);
xor UO_1480 (O_1480,N_24281,N_24223);
and UO_1481 (O_1481,N_23004,N_23992);
xnor UO_1482 (O_1482,N_23424,N_22770);
xnor UO_1483 (O_1483,N_23686,N_23189);
xor UO_1484 (O_1484,N_23089,N_22378);
xnor UO_1485 (O_1485,N_24309,N_21877);
xnor UO_1486 (O_1486,N_24900,N_22202);
or UO_1487 (O_1487,N_22985,N_24006);
nor UO_1488 (O_1488,N_24466,N_22267);
nand UO_1489 (O_1489,N_23513,N_23020);
nor UO_1490 (O_1490,N_21886,N_22080);
nor UO_1491 (O_1491,N_24067,N_22213);
xor UO_1492 (O_1492,N_23610,N_21965);
nor UO_1493 (O_1493,N_22798,N_22384);
nand UO_1494 (O_1494,N_23273,N_22113);
nand UO_1495 (O_1495,N_22795,N_22313);
nand UO_1496 (O_1496,N_23433,N_22442);
nor UO_1497 (O_1497,N_22643,N_23166);
nor UO_1498 (O_1498,N_23115,N_24481);
or UO_1499 (O_1499,N_22254,N_24474);
or UO_1500 (O_1500,N_24835,N_22879);
xnor UO_1501 (O_1501,N_24882,N_23215);
nor UO_1502 (O_1502,N_22215,N_23269);
or UO_1503 (O_1503,N_23523,N_22825);
nand UO_1504 (O_1504,N_24543,N_23880);
or UO_1505 (O_1505,N_23957,N_24883);
or UO_1506 (O_1506,N_23362,N_24581);
nor UO_1507 (O_1507,N_22678,N_21999);
or UO_1508 (O_1508,N_22342,N_24311);
and UO_1509 (O_1509,N_24902,N_23221);
nand UO_1510 (O_1510,N_24943,N_23222);
or UO_1511 (O_1511,N_24186,N_23271);
or UO_1512 (O_1512,N_24087,N_23962);
and UO_1513 (O_1513,N_23029,N_22940);
xor UO_1514 (O_1514,N_22860,N_23931);
and UO_1515 (O_1515,N_23657,N_21946);
nor UO_1516 (O_1516,N_23360,N_22520);
and UO_1517 (O_1517,N_24720,N_24347);
nand UO_1518 (O_1518,N_22063,N_22563);
nor UO_1519 (O_1519,N_24921,N_24120);
and UO_1520 (O_1520,N_22437,N_22994);
or UO_1521 (O_1521,N_22399,N_24191);
and UO_1522 (O_1522,N_24165,N_24784);
and UO_1523 (O_1523,N_24028,N_23918);
nor UO_1524 (O_1524,N_22778,N_24730);
and UO_1525 (O_1525,N_23354,N_24172);
nand UO_1526 (O_1526,N_24143,N_24961);
nor UO_1527 (O_1527,N_23561,N_24827);
nand UO_1528 (O_1528,N_22714,N_23998);
nand UO_1529 (O_1529,N_23346,N_24821);
nor UO_1530 (O_1530,N_23325,N_24219);
or UO_1531 (O_1531,N_23515,N_22954);
and UO_1532 (O_1532,N_22137,N_22754);
or UO_1533 (O_1533,N_24673,N_22690);
nand UO_1534 (O_1534,N_24201,N_22274);
or UO_1535 (O_1535,N_24393,N_23074);
or UO_1536 (O_1536,N_22595,N_23157);
and UO_1537 (O_1537,N_24360,N_21974);
nand UO_1538 (O_1538,N_22597,N_21898);
nor UO_1539 (O_1539,N_22214,N_24032);
nor UO_1540 (O_1540,N_24565,N_23217);
nand UO_1541 (O_1541,N_22786,N_22848);
nor UO_1542 (O_1542,N_22060,N_24721);
nand UO_1543 (O_1543,N_24131,N_23798);
or UO_1544 (O_1544,N_21988,N_23038);
nand UO_1545 (O_1545,N_23021,N_24495);
nand UO_1546 (O_1546,N_23789,N_23102);
nand UO_1547 (O_1547,N_23896,N_21940);
or UO_1548 (O_1548,N_23970,N_22652);
xnor UO_1549 (O_1549,N_22925,N_24278);
nor UO_1550 (O_1550,N_22008,N_21892);
xnor UO_1551 (O_1551,N_22761,N_22034);
nand UO_1552 (O_1552,N_22922,N_23374);
nand UO_1553 (O_1553,N_24244,N_22523);
or UO_1554 (O_1554,N_22006,N_24254);
xor UO_1555 (O_1555,N_23958,N_22463);
nand UO_1556 (O_1556,N_23615,N_22462);
or UO_1557 (O_1557,N_23940,N_24934);
or UO_1558 (O_1558,N_22067,N_23689);
and UO_1559 (O_1559,N_23563,N_24395);
xnor UO_1560 (O_1560,N_24007,N_24712);
nand UO_1561 (O_1561,N_23540,N_24373);
xnor UO_1562 (O_1562,N_22989,N_23895);
and UO_1563 (O_1563,N_24931,N_23607);
or UO_1564 (O_1564,N_23404,N_23882);
xor UO_1565 (O_1565,N_22439,N_22364);
or UO_1566 (O_1566,N_23063,N_22186);
xor UO_1567 (O_1567,N_22927,N_22225);
or UO_1568 (O_1568,N_22795,N_22253);
and UO_1569 (O_1569,N_24993,N_22985);
xor UO_1570 (O_1570,N_22835,N_24299);
xnor UO_1571 (O_1571,N_23491,N_22456);
xnor UO_1572 (O_1572,N_22930,N_24744);
nor UO_1573 (O_1573,N_23411,N_24594);
or UO_1574 (O_1574,N_22543,N_24028);
and UO_1575 (O_1575,N_24478,N_22192);
or UO_1576 (O_1576,N_24105,N_24147);
nand UO_1577 (O_1577,N_22320,N_24861);
nand UO_1578 (O_1578,N_24528,N_22048);
xnor UO_1579 (O_1579,N_24728,N_23034);
and UO_1580 (O_1580,N_24670,N_24269);
nor UO_1581 (O_1581,N_23550,N_23413);
nor UO_1582 (O_1582,N_23477,N_24984);
xnor UO_1583 (O_1583,N_22845,N_22234);
nand UO_1584 (O_1584,N_22023,N_23861);
nand UO_1585 (O_1585,N_24540,N_22474);
and UO_1586 (O_1586,N_23348,N_21912);
nand UO_1587 (O_1587,N_22322,N_23729);
nand UO_1588 (O_1588,N_24327,N_23504);
nor UO_1589 (O_1589,N_24041,N_24239);
and UO_1590 (O_1590,N_23216,N_23501);
nor UO_1591 (O_1591,N_24993,N_24514);
nand UO_1592 (O_1592,N_23532,N_23680);
nor UO_1593 (O_1593,N_24914,N_24340);
or UO_1594 (O_1594,N_22991,N_22046);
xor UO_1595 (O_1595,N_23026,N_24291);
or UO_1596 (O_1596,N_21900,N_24544);
nand UO_1597 (O_1597,N_23791,N_22113);
and UO_1598 (O_1598,N_24932,N_24019);
and UO_1599 (O_1599,N_23231,N_23982);
and UO_1600 (O_1600,N_22955,N_23026);
xor UO_1601 (O_1601,N_22261,N_24551);
or UO_1602 (O_1602,N_22693,N_22239);
or UO_1603 (O_1603,N_23891,N_22259);
or UO_1604 (O_1604,N_23169,N_22168);
and UO_1605 (O_1605,N_24594,N_23862);
nor UO_1606 (O_1606,N_22803,N_22677);
and UO_1607 (O_1607,N_23818,N_24511);
nand UO_1608 (O_1608,N_23676,N_23128);
xor UO_1609 (O_1609,N_23746,N_24244);
nor UO_1610 (O_1610,N_24073,N_24784);
nor UO_1611 (O_1611,N_24015,N_22009);
and UO_1612 (O_1612,N_24748,N_24879);
nor UO_1613 (O_1613,N_22199,N_23988);
or UO_1614 (O_1614,N_23940,N_22855);
nor UO_1615 (O_1615,N_24686,N_23160);
or UO_1616 (O_1616,N_24696,N_22073);
xnor UO_1617 (O_1617,N_23153,N_22967);
xnor UO_1618 (O_1618,N_23977,N_23787);
xor UO_1619 (O_1619,N_22280,N_22273);
and UO_1620 (O_1620,N_24258,N_23048);
xnor UO_1621 (O_1621,N_21929,N_23612);
or UO_1622 (O_1622,N_23601,N_22500);
nand UO_1623 (O_1623,N_24956,N_24824);
xnor UO_1624 (O_1624,N_24720,N_23099);
and UO_1625 (O_1625,N_22584,N_24151);
and UO_1626 (O_1626,N_22964,N_23668);
nor UO_1627 (O_1627,N_24061,N_24703);
xor UO_1628 (O_1628,N_24938,N_23598);
xnor UO_1629 (O_1629,N_22926,N_23235);
xor UO_1630 (O_1630,N_23773,N_22068);
nor UO_1631 (O_1631,N_22015,N_22749);
or UO_1632 (O_1632,N_23919,N_24837);
nor UO_1633 (O_1633,N_23820,N_24765);
or UO_1634 (O_1634,N_23899,N_24268);
xnor UO_1635 (O_1635,N_24345,N_24171);
xnor UO_1636 (O_1636,N_23466,N_23584);
nor UO_1637 (O_1637,N_23427,N_22484);
xor UO_1638 (O_1638,N_23164,N_24213);
and UO_1639 (O_1639,N_23154,N_24293);
xor UO_1640 (O_1640,N_24251,N_23399);
nand UO_1641 (O_1641,N_24738,N_24673);
and UO_1642 (O_1642,N_22549,N_24287);
nor UO_1643 (O_1643,N_24725,N_22810);
nor UO_1644 (O_1644,N_23381,N_24504);
and UO_1645 (O_1645,N_24719,N_23417);
nand UO_1646 (O_1646,N_24686,N_21903);
xnor UO_1647 (O_1647,N_24562,N_22325);
xnor UO_1648 (O_1648,N_23420,N_22021);
nand UO_1649 (O_1649,N_23603,N_22256);
nor UO_1650 (O_1650,N_22008,N_23518);
or UO_1651 (O_1651,N_24731,N_22588);
xnor UO_1652 (O_1652,N_22982,N_23850);
xor UO_1653 (O_1653,N_23963,N_24637);
xor UO_1654 (O_1654,N_24309,N_22103);
nor UO_1655 (O_1655,N_23254,N_23075);
and UO_1656 (O_1656,N_23124,N_23167);
or UO_1657 (O_1657,N_23749,N_22330);
nor UO_1658 (O_1658,N_22596,N_23404);
and UO_1659 (O_1659,N_24671,N_23604);
nor UO_1660 (O_1660,N_24787,N_24072);
or UO_1661 (O_1661,N_24870,N_24131);
or UO_1662 (O_1662,N_22154,N_22334);
nand UO_1663 (O_1663,N_24394,N_23597);
or UO_1664 (O_1664,N_23858,N_23289);
xor UO_1665 (O_1665,N_22907,N_24940);
nor UO_1666 (O_1666,N_22812,N_22108);
and UO_1667 (O_1667,N_24909,N_24557);
or UO_1668 (O_1668,N_22103,N_22786);
xor UO_1669 (O_1669,N_22554,N_22393);
and UO_1670 (O_1670,N_24106,N_21966);
or UO_1671 (O_1671,N_21919,N_23241);
or UO_1672 (O_1672,N_23969,N_24626);
xnor UO_1673 (O_1673,N_22278,N_22807);
nand UO_1674 (O_1674,N_24022,N_22118);
or UO_1675 (O_1675,N_23864,N_22890);
and UO_1676 (O_1676,N_24962,N_22072);
nand UO_1677 (O_1677,N_23184,N_24686);
nor UO_1678 (O_1678,N_24503,N_22337);
nand UO_1679 (O_1679,N_24277,N_23785);
xnor UO_1680 (O_1680,N_23604,N_23771);
and UO_1681 (O_1681,N_23588,N_24873);
and UO_1682 (O_1682,N_24228,N_24103);
nor UO_1683 (O_1683,N_23350,N_23376);
nand UO_1684 (O_1684,N_24070,N_22756);
nand UO_1685 (O_1685,N_22464,N_24522);
nor UO_1686 (O_1686,N_22063,N_24246);
nand UO_1687 (O_1687,N_24508,N_21954);
nor UO_1688 (O_1688,N_21959,N_22264);
xnor UO_1689 (O_1689,N_24522,N_23200);
nand UO_1690 (O_1690,N_22636,N_22600);
xor UO_1691 (O_1691,N_23202,N_23200);
xnor UO_1692 (O_1692,N_22225,N_23676);
nand UO_1693 (O_1693,N_21897,N_23802);
xor UO_1694 (O_1694,N_22944,N_23489);
nor UO_1695 (O_1695,N_23135,N_23863);
xnor UO_1696 (O_1696,N_24706,N_24150);
xor UO_1697 (O_1697,N_22743,N_23837);
nor UO_1698 (O_1698,N_24113,N_22804);
nand UO_1699 (O_1699,N_24947,N_22541);
nor UO_1700 (O_1700,N_24765,N_24191);
or UO_1701 (O_1701,N_23199,N_23334);
nor UO_1702 (O_1702,N_24924,N_23436);
nand UO_1703 (O_1703,N_23361,N_24732);
or UO_1704 (O_1704,N_22055,N_22714);
and UO_1705 (O_1705,N_22901,N_22470);
nand UO_1706 (O_1706,N_24756,N_24703);
xnor UO_1707 (O_1707,N_23297,N_23072);
and UO_1708 (O_1708,N_23525,N_24787);
nor UO_1709 (O_1709,N_23427,N_22317);
and UO_1710 (O_1710,N_23571,N_23077);
and UO_1711 (O_1711,N_22661,N_22162);
or UO_1712 (O_1712,N_23313,N_24010);
nand UO_1713 (O_1713,N_23416,N_22415);
and UO_1714 (O_1714,N_23828,N_23679);
xnor UO_1715 (O_1715,N_24279,N_22436);
xnor UO_1716 (O_1716,N_23006,N_22183);
nand UO_1717 (O_1717,N_23042,N_24711);
and UO_1718 (O_1718,N_22486,N_24183);
nor UO_1719 (O_1719,N_24593,N_22995);
or UO_1720 (O_1720,N_23180,N_23662);
nand UO_1721 (O_1721,N_21948,N_23561);
and UO_1722 (O_1722,N_22037,N_24440);
xor UO_1723 (O_1723,N_22109,N_23787);
or UO_1724 (O_1724,N_22449,N_23130);
xor UO_1725 (O_1725,N_23458,N_24941);
nand UO_1726 (O_1726,N_24016,N_23634);
nand UO_1727 (O_1727,N_23662,N_22658);
or UO_1728 (O_1728,N_21972,N_23933);
nor UO_1729 (O_1729,N_24280,N_23200);
xnor UO_1730 (O_1730,N_22673,N_23161);
and UO_1731 (O_1731,N_22443,N_24773);
or UO_1732 (O_1732,N_22980,N_22651);
or UO_1733 (O_1733,N_24631,N_23943);
xnor UO_1734 (O_1734,N_22387,N_23783);
and UO_1735 (O_1735,N_22970,N_24972);
and UO_1736 (O_1736,N_21941,N_22499);
nand UO_1737 (O_1737,N_24830,N_23478);
and UO_1738 (O_1738,N_22025,N_24915);
nor UO_1739 (O_1739,N_24901,N_22557);
and UO_1740 (O_1740,N_24416,N_23160);
nand UO_1741 (O_1741,N_23982,N_22587);
nor UO_1742 (O_1742,N_23089,N_24117);
and UO_1743 (O_1743,N_23255,N_23984);
and UO_1744 (O_1744,N_23444,N_22641);
nor UO_1745 (O_1745,N_24755,N_24292);
nand UO_1746 (O_1746,N_22154,N_24046);
or UO_1747 (O_1747,N_22677,N_21933);
or UO_1748 (O_1748,N_23216,N_24257);
xnor UO_1749 (O_1749,N_22379,N_21924);
and UO_1750 (O_1750,N_24333,N_23644);
nor UO_1751 (O_1751,N_22480,N_23785);
nand UO_1752 (O_1752,N_22049,N_23856);
or UO_1753 (O_1753,N_21917,N_23629);
or UO_1754 (O_1754,N_23762,N_24546);
nor UO_1755 (O_1755,N_22970,N_23602);
and UO_1756 (O_1756,N_22203,N_24717);
nand UO_1757 (O_1757,N_24130,N_24454);
nor UO_1758 (O_1758,N_23009,N_22490);
and UO_1759 (O_1759,N_24558,N_23149);
and UO_1760 (O_1760,N_23993,N_22301);
nand UO_1761 (O_1761,N_21883,N_24122);
nor UO_1762 (O_1762,N_24262,N_22655);
nor UO_1763 (O_1763,N_24482,N_22026);
xor UO_1764 (O_1764,N_24389,N_22287);
or UO_1765 (O_1765,N_23400,N_23527);
xor UO_1766 (O_1766,N_23263,N_23527);
nor UO_1767 (O_1767,N_23265,N_23574);
or UO_1768 (O_1768,N_24805,N_22907);
and UO_1769 (O_1769,N_23470,N_24951);
nor UO_1770 (O_1770,N_23779,N_24094);
xor UO_1771 (O_1771,N_24958,N_23893);
nand UO_1772 (O_1772,N_22293,N_23403);
xor UO_1773 (O_1773,N_22143,N_22768);
nor UO_1774 (O_1774,N_23315,N_23498);
xnor UO_1775 (O_1775,N_22644,N_23425);
and UO_1776 (O_1776,N_24422,N_22566);
and UO_1777 (O_1777,N_24568,N_24157);
nand UO_1778 (O_1778,N_24745,N_22337);
xor UO_1779 (O_1779,N_23460,N_23700);
or UO_1780 (O_1780,N_23362,N_22119);
or UO_1781 (O_1781,N_24546,N_23184);
and UO_1782 (O_1782,N_22746,N_24807);
nand UO_1783 (O_1783,N_24992,N_22448);
nand UO_1784 (O_1784,N_22452,N_24305);
and UO_1785 (O_1785,N_22559,N_22589);
or UO_1786 (O_1786,N_23783,N_22265);
and UO_1787 (O_1787,N_23283,N_23644);
nand UO_1788 (O_1788,N_22671,N_22643);
and UO_1789 (O_1789,N_24221,N_24526);
xnor UO_1790 (O_1790,N_24149,N_23744);
xor UO_1791 (O_1791,N_24374,N_22197);
and UO_1792 (O_1792,N_22350,N_23294);
nor UO_1793 (O_1793,N_24033,N_22304);
nand UO_1794 (O_1794,N_21979,N_22571);
and UO_1795 (O_1795,N_24086,N_24488);
or UO_1796 (O_1796,N_23407,N_23837);
or UO_1797 (O_1797,N_23078,N_24646);
or UO_1798 (O_1798,N_22586,N_23454);
xnor UO_1799 (O_1799,N_22759,N_22712);
nand UO_1800 (O_1800,N_23176,N_22273);
or UO_1801 (O_1801,N_23683,N_22392);
nor UO_1802 (O_1802,N_21898,N_23087);
or UO_1803 (O_1803,N_23322,N_23354);
xnor UO_1804 (O_1804,N_22791,N_23732);
or UO_1805 (O_1805,N_23294,N_23626);
nor UO_1806 (O_1806,N_24575,N_24367);
xor UO_1807 (O_1807,N_24363,N_21895);
nor UO_1808 (O_1808,N_22116,N_23844);
xor UO_1809 (O_1809,N_23170,N_23434);
nand UO_1810 (O_1810,N_24819,N_23385);
nand UO_1811 (O_1811,N_23310,N_22058);
and UO_1812 (O_1812,N_23026,N_24932);
and UO_1813 (O_1813,N_23852,N_24473);
xor UO_1814 (O_1814,N_24018,N_22629);
xor UO_1815 (O_1815,N_23972,N_22959);
nand UO_1816 (O_1816,N_23778,N_23430);
nor UO_1817 (O_1817,N_23759,N_22730);
or UO_1818 (O_1818,N_24692,N_23646);
and UO_1819 (O_1819,N_23745,N_24238);
nor UO_1820 (O_1820,N_23015,N_24766);
or UO_1821 (O_1821,N_24363,N_23154);
xnor UO_1822 (O_1822,N_23324,N_23458);
xor UO_1823 (O_1823,N_22985,N_23727);
or UO_1824 (O_1824,N_24889,N_24614);
or UO_1825 (O_1825,N_23752,N_22683);
and UO_1826 (O_1826,N_23731,N_24351);
and UO_1827 (O_1827,N_22833,N_23020);
xor UO_1828 (O_1828,N_23516,N_22695);
or UO_1829 (O_1829,N_22551,N_22406);
or UO_1830 (O_1830,N_22739,N_23042);
or UO_1831 (O_1831,N_24320,N_23238);
xnor UO_1832 (O_1832,N_22940,N_23757);
and UO_1833 (O_1833,N_23196,N_24830);
xnor UO_1834 (O_1834,N_23066,N_22525);
and UO_1835 (O_1835,N_22206,N_22590);
or UO_1836 (O_1836,N_24003,N_22760);
xor UO_1837 (O_1837,N_24239,N_21939);
xnor UO_1838 (O_1838,N_22987,N_24047);
nor UO_1839 (O_1839,N_24841,N_22191);
xnor UO_1840 (O_1840,N_22322,N_23758);
nand UO_1841 (O_1841,N_22212,N_21933);
nor UO_1842 (O_1842,N_24319,N_23276);
and UO_1843 (O_1843,N_21978,N_23485);
xnor UO_1844 (O_1844,N_23024,N_22019);
and UO_1845 (O_1845,N_24106,N_22828);
nand UO_1846 (O_1846,N_22985,N_23609);
or UO_1847 (O_1847,N_22303,N_24698);
and UO_1848 (O_1848,N_22235,N_22596);
nand UO_1849 (O_1849,N_22506,N_23617);
or UO_1850 (O_1850,N_24065,N_22552);
nor UO_1851 (O_1851,N_23127,N_22834);
xor UO_1852 (O_1852,N_22154,N_22693);
or UO_1853 (O_1853,N_24898,N_24241);
or UO_1854 (O_1854,N_24367,N_23665);
or UO_1855 (O_1855,N_23580,N_22962);
and UO_1856 (O_1856,N_24177,N_23518);
nor UO_1857 (O_1857,N_21913,N_24018);
nor UO_1858 (O_1858,N_21913,N_23358);
nand UO_1859 (O_1859,N_23651,N_22580);
xor UO_1860 (O_1860,N_24604,N_22420);
xnor UO_1861 (O_1861,N_23281,N_24233);
or UO_1862 (O_1862,N_24995,N_24785);
and UO_1863 (O_1863,N_21909,N_22516);
or UO_1864 (O_1864,N_23559,N_21916);
and UO_1865 (O_1865,N_23673,N_23115);
and UO_1866 (O_1866,N_22832,N_24515);
nor UO_1867 (O_1867,N_23766,N_22788);
xnor UO_1868 (O_1868,N_23033,N_23604);
or UO_1869 (O_1869,N_22648,N_24261);
or UO_1870 (O_1870,N_23287,N_22027);
nor UO_1871 (O_1871,N_23308,N_24602);
nor UO_1872 (O_1872,N_23843,N_22206);
xor UO_1873 (O_1873,N_22230,N_22263);
nor UO_1874 (O_1874,N_24348,N_24303);
and UO_1875 (O_1875,N_22659,N_21969);
and UO_1876 (O_1876,N_22851,N_22183);
nand UO_1877 (O_1877,N_23292,N_24754);
xor UO_1878 (O_1878,N_23439,N_23149);
nand UO_1879 (O_1879,N_22372,N_22509);
nor UO_1880 (O_1880,N_24566,N_23077);
xor UO_1881 (O_1881,N_24130,N_22141);
nand UO_1882 (O_1882,N_22558,N_22845);
nand UO_1883 (O_1883,N_23467,N_24220);
or UO_1884 (O_1884,N_22027,N_24090);
xor UO_1885 (O_1885,N_22383,N_24402);
nand UO_1886 (O_1886,N_24079,N_24638);
and UO_1887 (O_1887,N_22925,N_24680);
nor UO_1888 (O_1888,N_23480,N_22126);
nand UO_1889 (O_1889,N_21979,N_24245);
or UO_1890 (O_1890,N_24905,N_23460);
or UO_1891 (O_1891,N_22530,N_22891);
or UO_1892 (O_1892,N_23788,N_24889);
nor UO_1893 (O_1893,N_22649,N_24961);
nand UO_1894 (O_1894,N_23381,N_22309);
nor UO_1895 (O_1895,N_23165,N_23940);
xnor UO_1896 (O_1896,N_22844,N_22691);
or UO_1897 (O_1897,N_21967,N_22008);
nor UO_1898 (O_1898,N_23267,N_24203);
xor UO_1899 (O_1899,N_24049,N_24809);
nand UO_1900 (O_1900,N_23690,N_24369);
and UO_1901 (O_1901,N_23214,N_24402);
xor UO_1902 (O_1902,N_23739,N_24389);
nand UO_1903 (O_1903,N_24478,N_24674);
nor UO_1904 (O_1904,N_24393,N_23766);
nand UO_1905 (O_1905,N_23212,N_24965);
and UO_1906 (O_1906,N_23886,N_23376);
nor UO_1907 (O_1907,N_22444,N_23702);
nor UO_1908 (O_1908,N_24373,N_24860);
xor UO_1909 (O_1909,N_23409,N_22180);
and UO_1910 (O_1910,N_23144,N_24817);
or UO_1911 (O_1911,N_21893,N_23027);
nand UO_1912 (O_1912,N_22539,N_23673);
or UO_1913 (O_1913,N_23850,N_23570);
nor UO_1914 (O_1914,N_24160,N_24529);
xnor UO_1915 (O_1915,N_22715,N_24773);
nand UO_1916 (O_1916,N_22212,N_23611);
nand UO_1917 (O_1917,N_23883,N_24571);
and UO_1918 (O_1918,N_22704,N_22988);
and UO_1919 (O_1919,N_23374,N_22956);
or UO_1920 (O_1920,N_23604,N_21972);
xnor UO_1921 (O_1921,N_21985,N_24540);
xnor UO_1922 (O_1922,N_22046,N_24229);
or UO_1923 (O_1923,N_22322,N_24119);
and UO_1924 (O_1924,N_23308,N_24394);
or UO_1925 (O_1925,N_23545,N_23867);
or UO_1926 (O_1926,N_24943,N_24876);
nor UO_1927 (O_1927,N_23352,N_22951);
or UO_1928 (O_1928,N_23892,N_22862);
and UO_1929 (O_1929,N_24529,N_24597);
and UO_1930 (O_1930,N_24227,N_22694);
xor UO_1931 (O_1931,N_22298,N_23959);
and UO_1932 (O_1932,N_24319,N_23981);
xnor UO_1933 (O_1933,N_23028,N_23813);
nand UO_1934 (O_1934,N_24565,N_22231);
nor UO_1935 (O_1935,N_23231,N_21879);
and UO_1936 (O_1936,N_23833,N_24186);
and UO_1937 (O_1937,N_24904,N_24432);
nor UO_1938 (O_1938,N_22778,N_23495);
nor UO_1939 (O_1939,N_23398,N_22145);
xor UO_1940 (O_1940,N_23656,N_22565);
nand UO_1941 (O_1941,N_24502,N_24392);
xor UO_1942 (O_1942,N_22132,N_23502);
xor UO_1943 (O_1943,N_22382,N_24527);
nand UO_1944 (O_1944,N_23340,N_24761);
nand UO_1945 (O_1945,N_23765,N_22831);
nor UO_1946 (O_1946,N_21984,N_24606);
xor UO_1947 (O_1947,N_23617,N_24295);
and UO_1948 (O_1948,N_23189,N_23285);
xnor UO_1949 (O_1949,N_23110,N_22654);
nor UO_1950 (O_1950,N_23305,N_24573);
xor UO_1951 (O_1951,N_24081,N_23517);
xor UO_1952 (O_1952,N_24209,N_22242);
and UO_1953 (O_1953,N_23247,N_22174);
or UO_1954 (O_1954,N_23312,N_24165);
or UO_1955 (O_1955,N_23898,N_24099);
xnor UO_1956 (O_1956,N_23621,N_24187);
xnor UO_1957 (O_1957,N_23280,N_22619);
or UO_1958 (O_1958,N_22531,N_22860);
or UO_1959 (O_1959,N_22103,N_22093);
nor UO_1960 (O_1960,N_23514,N_23929);
nand UO_1961 (O_1961,N_23501,N_24478);
xor UO_1962 (O_1962,N_22974,N_22643);
nor UO_1963 (O_1963,N_22449,N_23206);
and UO_1964 (O_1964,N_24334,N_24377);
or UO_1965 (O_1965,N_23786,N_24428);
or UO_1966 (O_1966,N_24285,N_22336);
nor UO_1967 (O_1967,N_22640,N_22996);
nand UO_1968 (O_1968,N_24868,N_24756);
xnor UO_1969 (O_1969,N_24884,N_22595);
or UO_1970 (O_1970,N_22361,N_22288);
nor UO_1971 (O_1971,N_22901,N_24656);
nor UO_1972 (O_1972,N_22930,N_24624);
or UO_1973 (O_1973,N_22341,N_24903);
nor UO_1974 (O_1974,N_22164,N_23961);
nand UO_1975 (O_1975,N_24517,N_23671);
and UO_1976 (O_1976,N_22945,N_24145);
nor UO_1977 (O_1977,N_21905,N_24456);
xor UO_1978 (O_1978,N_22890,N_23390);
xor UO_1979 (O_1979,N_23014,N_22475);
or UO_1980 (O_1980,N_23381,N_24756);
or UO_1981 (O_1981,N_22242,N_23267);
and UO_1982 (O_1982,N_22169,N_22770);
xor UO_1983 (O_1983,N_24261,N_24871);
nand UO_1984 (O_1984,N_24409,N_23260);
nand UO_1985 (O_1985,N_23344,N_24194);
and UO_1986 (O_1986,N_24151,N_23522);
nor UO_1987 (O_1987,N_21987,N_22207);
xnor UO_1988 (O_1988,N_22880,N_22300);
or UO_1989 (O_1989,N_22260,N_21894);
xnor UO_1990 (O_1990,N_23149,N_24609);
nand UO_1991 (O_1991,N_23350,N_24121);
or UO_1992 (O_1992,N_24588,N_24378);
and UO_1993 (O_1993,N_22602,N_22379);
or UO_1994 (O_1994,N_23194,N_23561);
or UO_1995 (O_1995,N_23900,N_24730);
xnor UO_1996 (O_1996,N_22740,N_24170);
nand UO_1997 (O_1997,N_24211,N_23099);
nor UO_1998 (O_1998,N_24773,N_23698);
and UO_1999 (O_1999,N_22652,N_23818);
nor UO_2000 (O_2000,N_23089,N_24008);
xnor UO_2001 (O_2001,N_22107,N_21933);
or UO_2002 (O_2002,N_24634,N_24494);
nor UO_2003 (O_2003,N_22312,N_22205);
and UO_2004 (O_2004,N_24604,N_24208);
and UO_2005 (O_2005,N_22134,N_22367);
xor UO_2006 (O_2006,N_24307,N_24856);
or UO_2007 (O_2007,N_22626,N_23902);
nand UO_2008 (O_2008,N_23197,N_22180);
nor UO_2009 (O_2009,N_23919,N_22733);
nor UO_2010 (O_2010,N_23931,N_21919);
xor UO_2011 (O_2011,N_24783,N_23324);
nand UO_2012 (O_2012,N_24650,N_24432);
xor UO_2013 (O_2013,N_23486,N_23069);
or UO_2014 (O_2014,N_24781,N_22394);
or UO_2015 (O_2015,N_22926,N_23386);
nor UO_2016 (O_2016,N_22000,N_22782);
nor UO_2017 (O_2017,N_24042,N_22053);
or UO_2018 (O_2018,N_22303,N_23565);
xor UO_2019 (O_2019,N_24394,N_22205);
nor UO_2020 (O_2020,N_22653,N_23617);
nor UO_2021 (O_2021,N_22302,N_23542);
or UO_2022 (O_2022,N_22015,N_23858);
or UO_2023 (O_2023,N_22939,N_24037);
or UO_2024 (O_2024,N_23864,N_24103);
nor UO_2025 (O_2025,N_23470,N_24542);
xnor UO_2026 (O_2026,N_22764,N_22411);
or UO_2027 (O_2027,N_24129,N_22769);
and UO_2028 (O_2028,N_24084,N_23983);
xnor UO_2029 (O_2029,N_24164,N_22827);
and UO_2030 (O_2030,N_23094,N_22216);
xor UO_2031 (O_2031,N_23359,N_21959);
xor UO_2032 (O_2032,N_23043,N_22932);
xor UO_2033 (O_2033,N_24404,N_23376);
and UO_2034 (O_2034,N_24639,N_23285);
and UO_2035 (O_2035,N_23040,N_22274);
xor UO_2036 (O_2036,N_23176,N_22477);
or UO_2037 (O_2037,N_23213,N_24783);
and UO_2038 (O_2038,N_22837,N_24182);
nand UO_2039 (O_2039,N_22720,N_24094);
or UO_2040 (O_2040,N_24388,N_23916);
xor UO_2041 (O_2041,N_23043,N_21897);
nor UO_2042 (O_2042,N_22625,N_24792);
xor UO_2043 (O_2043,N_24011,N_22394);
nor UO_2044 (O_2044,N_22800,N_24728);
nor UO_2045 (O_2045,N_23134,N_22678);
xor UO_2046 (O_2046,N_22900,N_23020);
nand UO_2047 (O_2047,N_24695,N_22861);
and UO_2048 (O_2048,N_23130,N_22364);
nor UO_2049 (O_2049,N_22753,N_24951);
nor UO_2050 (O_2050,N_24468,N_22818);
and UO_2051 (O_2051,N_23964,N_22303);
or UO_2052 (O_2052,N_22455,N_22667);
or UO_2053 (O_2053,N_24509,N_23067);
and UO_2054 (O_2054,N_24851,N_24501);
and UO_2055 (O_2055,N_24858,N_22691);
or UO_2056 (O_2056,N_22187,N_22441);
nand UO_2057 (O_2057,N_24355,N_22197);
or UO_2058 (O_2058,N_23821,N_23985);
or UO_2059 (O_2059,N_23668,N_24557);
or UO_2060 (O_2060,N_24451,N_22132);
xnor UO_2061 (O_2061,N_22288,N_24014);
xor UO_2062 (O_2062,N_23717,N_22452);
nor UO_2063 (O_2063,N_24404,N_24481);
and UO_2064 (O_2064,N_23137,N_24015);
nand UO_2065 (O_2065,N_23972,N_24723);
xnor UO_2066 (O_2066,N_22376,N_22115);
nor UO_2067 (O_2067,N_22604,N_24643);
nor UO_2068 (O_2068,N_22170,N_24524);
xnor UO_2069 (O_2069,N_22034,N_24968);
or UO_2070 (O_2070,N_23155,N_22189);
and UO_2071 (O_2071,N_24890,N_24795);
nand UO_2072 (O_2072,N_22112,N_24401);
and UO_2073 (O_2073,N_22395,N_22474);
and UO_2074 (O_2074,N_21937,N_24429);
or UO_2075 (O_2075,N_23816,N_21876);
and UO_2076 (O_2076,N_22813,N_22270);
xor UO_2077 (O_2077,N_22623,N_24020);
xnor UO_2078 (O_2078,N_23086,N_24525);
nand UO_2079 (O_2079,N_23813,N_22354);
and UO_2080 (O_2080,N_21890,N_21937);
or UO_2081 (O_2081,N_22986,N_22910);
xor UO_2082 (O_2082,N_24967,N_23833);
nor UO_2083 (O_2083,N_24001,N_23513);
nand UO_2084 (O_2084,N_23782,N_22697);
nand UO_2085 (O_2085,N_23665,N_23925);
nand UO_2086 (O_2086,N_24921,N_23569);
and UO_2087 (O_2087,N_23090,N_23488);
xnor UO_2088 (O_2088,N_24951,N_21905);
nor UO_2089 (O_2089,N_22983,N_24640);
nor UO_2090 (O_2090,N_24524,N_24042);
nand UO_2091 (O_2091,N_22695,N_21933);
or UO_2092 (O_2092,N_23924,N_23861);
nor UO_2093 (O_2093,N_24247,N_22434);
and UO_2094 (O_2094,N_23483,N_23975);
nand UO_2095 (O_2095,N_22394,N_21914);
xor UO_2096 (O_2096,N_23197,N_23559);
nor UO_2097 (O_2097,N_24990,N_23149);
and UO_2098 (O_2098,N_22072,N_23024);
xor UO_2099 (O_2099,N_22802,N_23040);
xor UO_2100 (O_2100,N_24065,N_24777);
xnor UO_2101 (O_2101,N_23438,N_22856);
xnor UO_2102 (O_2102,N_24260,N_22089);
xnor UO_2103 (O_2103,N_24144,N_22113);
and UO_2104 (O_2104,N_24693,N_24850);
xor UO_2105 (O_2105,N_24313,N_21964);
xor UO_2106 (O_2106,N_23063,N_22915);
xnor UO_2107 (O_2107,N_23010,N_23169);
nand UO_2108 (O_2108,N_21937,N_22636);
or UO_2109 (O_2109,N_23303,N_24628);
xnor UO_2110 (O_2110,N_24196,N_22846);
and UO_2111 (O_2111,N_23822,N_24083);
nor UO_2112 (O_2112,N_23106,N_23425);
xor UO_2113 (O_2113,N_23007,N_24564);
nand UO_2114 (O_2114,N_23887,N_22028);
and UO_2115 (O_2115,N_24873,N_24439);
nand UO_2116 (O_2116,N_23341,N_23058);
nor UO_2117 (O_2117,N_24332,N_23890);
and UO_2118 (O_2118,N_22218,N_23111);
nor UO_2119 (O_2119,N_23582,N_23020);
xnor UO_2120 (O_2120,N_24194,N_22193);
nand UO_2121 (O_2121,N_23907,N_22332);
xnor UO_2122 (O_2122,N_22474,N_22046);
xnor UO_2123 (O_2123,N_23230,N_24580);
nor UO_2124 (O_2124,N_24673,N_23919);
xnor UO_2125 (O_2125,N_22899,N_22591);
nand UO_2126 (O_2126,N_24943,N_23927);
nand UO_2127 (O_2127,N_24681,N_24519);
xnor UO_2128 (O_2128,N_23813,N_22107);
xor UO_2129 (O_2129,N_24489,N_24564);
nand UO_2130 (O_2130,N_23708,N_22863);
and UO_2131 (O_2131,N_23881,N_22217);
and UO_2132 (O_2132,N_22541,N_23552);
xor UO_2133 (O_2133,N_23186,N_23365);
or UO_2134 (O_2134,N_23491,N_23935);
nand UO_2135 (O_2135,N_24565,N_24652);
and UO_2136 (O_2136,N_21883,N_23115);
nand UO_2137 (O_2137,N_23934,N_22929);
or UO_2138 (O_2138,N_23819,N_22991);
nor UO_2139 (O_2139,N_22787,N_24389);
or UO_2140 (O_2140,N_24658,N_23082);
xnor UO_2141 (O_2141,N_23487,N_24118);
or UO_2142 (O_2142,N_22399,N_22812);
or UO_2143 (O_2143,N_22192,N_22003);
and UO_2144 (O_2144,N_23385,N_24378);
and UO_2145 (O_2145,N_22660,N_24671);
or UO_2146 (O_2146,N_24081,N_23815);
nor UO_2147 (O_2147,N_22786,N_22940);
and UO_2148 (O_2148,N_22955,N_22180);
and UO_2149 (O_2149,N_23402,N_24174);
and UO_2150 (O_2150,N_24567,N_23674);
and UO_2151 (O_2151,N_22707,N_22832);
nor UO_2152 (O_2152,N_24502,N_23621);
xor UO_2153 (O_2153,N_22721,N_24271);
xnor UO_2154 (O_2154,N_22559,N_24381);
nor UO_2155 (O_2155,N_24555,N_24404);
or UO_2156 (O_2156,N_24811,N_22203);
or UO_2157 (O_2157,N_23500,N_24672);
and UO_2158 (O_2158,N_22404,N_22216);
xor UO_2159 (O_2159,N_24861,N_23842);
xnor UO_2160 (O_2160,N_21941,N_24259);
or UO_2161 (O_2161,N_24143,N_22157);
xnor UO_2162 (O_2162,N_24898,N_24744);
and UO_2163 (O_2163,N_24305,N_23495);
or UO_2164 (O_2164,N_23186,N_22664);
and UO_2165 (O_2165,N_22536,N_22697);
or UO_2166 (O_2166,N_22561,N_24108);
nor UO_2167 (O_2167,N_24604,N_24798);
nand UO_2168 (O_2168,N_24958,N_22278);
xor UO_2169 (O_2169,N_22067,N_24913);
or UO_2170 (O_2170,N_24686,N_24860);
nor UO_2171 (O_2171,N_24554,N_22193);
xor UO_2172 (O_2172,N_23928,N_23800);
xnor UO_2173 (O_2173,N_22334,N_24785);
or UO_2174 (O_2174,N_23494,N_22527);
xnor UO_2175 (O_2175,N_22402,N_23305);
and UO_2176 (O_2176,N_23595,N_23306);
xnor UO_2177 (O_2177,N_22366,N_22304);
nand UO_2178 (O_2178,N_23552,N_24326);
xnor UO_2179 (O_2179,N_23975,N_23947);
or UO_2180 (O_2180,N_24656,N_22695);
or UO_2181 (O_2181,N_22996,N_22172);
and UO_2182 (O_2182,N_23214,N_22344);
and UO_2183 (O_2183,N_23162,N_22307);
nor UO_2184 (O_2184,N_23209,N_24863);
and UO_2185 (O_2185,N_22522,N_23595);
and UO_2186 (O_2186,N_23283,N_22441);
nor UO_2187 (O_2187,N_23567,N_23773);
nand UO_2188 (O_2188,N_24977,N_22087);
nor UO_2189 (O_2189,N_22058,N_24984);
nor UO_2190 (O_2190,N_22891,N_23682);
or UO_2191 (O_2191,N_23828,N_24421);
xor UO_2192 (O_2192,N_24830,N_23519);
or UO_2193 (O_2193,N_23722,N_23136);
nand UO_2194 (O_2194,N_23173,N_23129);
or UO_2195 (O_2195,N_24496,N_21898);
or UO_2196 (O_2196,N_22508,N_23967);
nand UO_2197 (O_2197,N_24409,N_21967);
xnor UO_2198 (O_2198,N_24126,N_22916);
xor UO_2199 (O_2199,N_22725,N_21917);
xnor UO_2200 (O_2200,N_23764,N_24342);
nand UO_2201 (O_2201,N_23300,N_24084);
nor UO_2202 (O_2202,N_23622,N_23646);
nor UO_2203 (O_2203,N_22018,N_24768);
and UO_2204 (O_2204,N_23060,N_24186);
xor UO_2205 (O_2205,N_24565,N_23413);
xnor UO_2206 (O_2206,N_23912,N_23933);
nand UO_2207 (O_2207,N_22674,N_24621);
or UO_2208 (O_2208,N_22576,N_23504);
nor UO_2209 (O_2209,N_23841,N_24096);
nor UO_2210 (O_2210,N_22308,N_22144);
or UO_2211 (O_2211,N_24375,N_23151);
nand UO_2212 (O_2212,N_22078,N_24957);
nor UO_2213 (O_2213,N_23737,N_22436);
nor UO_2214 (O_2214,N_22108,N_23903);
and UO_2215 (O_2215,N_22402,N_24506);
or UO_2216 (O_2216,N_24514,N_24331);
or UO_2217 (O_2217,N_24034,N_23774);
nor UO_2218 (O_2218,N_22986,N_23402);
and UO_2219 (O_2219,N_23908,N_23024);
xor UO_2220 (O_2220,N_23545,N_24941);
nor UO_2221 (O_2221,N_21875,N_23413);
and UO_2222 (O_2222,N_22508,N_24641);
and UO_2223 (O_2223,N_22806,N_24523);
nor UO_2224 (O_2224,N_23891,N_24691);
or UO_2225 (O_2225,N_23710,N_23322);
xnor UO_2226 (O_2226,N_23911,N_22254);
xor UO_2227 (O_2227,N_24573,N_22942);
xor UO_2228 (O_2228,N_22481,N_23729);
and UO_2229 (O_2229,N_24521,N_22934);
xor UO_2230 (O_2230,N_24688,N_24214);
nand UO_2231 (O_2231,N_23199,N_24029);
and UO_2232 (O_2232,N_23966,N_23968);
nand UO_2233 (O_2233,N_24065,N_24694);
nor UO_2234 (O_2234,N_22003,N_23101);
xor UO_2235 (O_2235,N_22626,N_22236);
nand UO_2236 (O_2236,N_24557,N_22130);
nor UO_2237 (O_2237,N_24093,N_24173);
and UO_2238 (O_2238,N_22393,N_23377);
or UO_2239 (O_2239,N_22911,N_21948);
xor UO_2240 (O_2240,N_23545,N_23247);
nor UO_2241 (O_2241,N_24207,N_22410);
xnor UO_2242 (O_2242,N_23735,N_22859);
or UO_2243 (O_2243,N_22440,N_23285);
nand UO_2244 (O_2244,N_22952,N_22916);
nand UO_2245 (O_2245,N_24516,N_23404);
nand UO_2246 (O_2246,N_24221,N_24451);
and UO_2247 (O_2247,N_24285,N_24716);
xor UO_2248 (O_2248,N_22407,N_22571);
nand UO_2249 (O_2249,N_24664,N_23040);
xnor UO_2250 (O_2250,N_23078,N_24058);
or UO_2251 (O_2251,N_24639,N_22841);
or UO_2252 (O_2252,N_24453,N_22029);
xnor UO_2253 (O_2253,N_24627,N_23021);
nand UO_2254 (O_2254,N_23995,N_21935);
or UO_2255 (O_2255,N_22290,N_23292);
nand UO_2256 (O_2256,N_22157,N_22932);
and UO_2257 (O_2257,N_22595,N_24647);
xnor UO_2258 (O_2258,N_24384,N_24833);
or UO_2259 (O_2259,N_23536,N_23562);
nand UO_2260 (O_2260,N_24949,N_23984);
or UO_2261 (O_2261,N_22834,N_24286);
nand UO_2262 (O_2262,N_22738,N_23953);
or UO_2263 (O_2263,N_23522,N_22877);
or UO_2264 (O_2264,N_23557,N_23706);
nand UO_2265 (O_2265,N_23195,N_24821);
xor UO_2266 (O_2266,N_22262,N_23376);
or UO_2267 (O_2267,N_24455,N_22181);
and UO_2268 (O_2268,N_24498,N_23518);
or UO_2269 (O_2269,N_22759,N_24886);
and UO_2270 (O_2270,N_21904,N_24988);
nor UO_2271 (O_2271,N_24988,N_24551);
xnor UO_2272 (O_2272,N_22994,N_24160);
nor UO_2273 (O_2273,N_21943,N_22222);
xnor UO_2274 (O_2274,N_24711,N_22244);
nand UO_2275 (O_2275,N_23135,N_23835);
and UO_2276 (O_2276,N_21973,N_23169);
nand UO_2277 (O_2277,N_24565,N_22093);
xor UO_2278 (O_2278,N_22039,N_23846);
nand UO_2279 (O_2279,N_22938,N_23538);
and UO_2280 (O_2280,N_24868,N_23157);
nor UO_2281 (O_2281,N_22228,N_23792);
nor UO_2282 (O_2282,N_23610,N_24105);
xor UO_2283 (O_2283,N_22896,N_21943);
xnor UO_2284 (O_2284,N_23327,N_23837);
or UO_2285 (O_2285,N_24862,N_23937);
xor UO_2286 (O_2286,N_24609,N_24967);
nand UO_2287 (O_2287,N_23868,N_22631);
and UO_2288 (O_2288,N_23171,N_24081);
nor UO_2289 (O_2289,N_24667,N_23326);
nand UO_2290 (O_2290,N_22883,N_23595);
xnor UO_2291 (O_2291,N_23003,N_23959);
or UO_2292 (O_2292,N_22751,N_23946);
nand UO_2293 (O_2293,N_23951,N_22898);
nor UO_2294 (O_2294,N_24820,N_21968);
nand UO_2295 (O_2295,N_23569,N_21881);
nand UO_2296 (O_2296,N_22458,N_22078);
and UO_2297 (O_2297,N_22316,N_23893);
or UO_2298 (O_2298,N_23825,N_22506);
nor UO_2299 (O_2299,N_22537,N_24593);
xor UO_2300 (O_2300,N_22567,N_22822);
nand UO_2301 (O_2301,N_23075,N_23103);
xor UO_2302 (O_2302,N_23783,N_24104);
nand UO_2303 (O_2303,N_23829,N_24548);
nand UO_2304 (O_2304,N_23969,N_24557);
nand UO_2305 (O_2305,N_22445,N_22459);
nand UO_2306 (O_2306,N_23791,N_24855);
or UO_2307 (O_2307,N_23435,N_24496);
xnor UO_2308 (O_2308,N_22760,N_22833);
nand UO_2309 (O_2309,N_22114,N_23612);
nand UO_2310 (O_2310,N_22358,N_23775);
and UO_2311 (O_2311,N_22537,N_24084);
xor UO_2312 (O_2312,N_24163,N_23928);
nor UO_2313 (O_2313,N_24416,N_24874);
nor UO_2314 (O_2314,N_23778,N_22354);
xnor UO_2315 (O_2315,N_22733,N_22211);
or UO_2316 (O_2316,N_22414,N_24636);
xor UO_2317 (O_2317,N_22382,N_24902);
and UO_2318 (O_2318,N_23288,N_22493);
or UO_2319 (O_2319,N_23662,N_24776);
and UO_2320 (O_2320,N_24566,N_22700);
and UO_2321 (O_2321,N_24795,N_23936);
xor UO_2322 (O_2322,N_24695,N_24190);
or UO_2323 (O_2323,N_22376,N_24220);
or UO_2324 (O_2324,N_24621,N_22036);
or UO_2325 (O_2325,N_24264,N_22560);
xnor UO_2326 (O_2326,N_23703,N_23812);
xor UO_2327 (O_2327,N_23548,N_23219);
nor UO_2328 (O_2328,N_23920,N_23867);
nor UO_2329 (O_2329,N_24308,N_22641);
or UO_2330 (O_2330,N_24779,N_22966);
nand UO_2331 (O_2331,N_24237,N_22087);
nand UO_2332 (O_2332,N_22586,N_24328);
xor UO_2333 (O_2333,N_23091,N_24809);
nor UO_2334 (O_2334,N_24198,N_24357);
xor UO_2335 (O_2335,N_23170,N_24308);
xnor UO_2336 (O_2336,N_23859,N_24325);
nand UO_2337 (O_2337,N_22966,N_24377);
nand UO_2338 (O_2338,N_24022,N_24895);
nand UO_2339 (O_2339,N_22710,N_24954);
nor UO_2340 (O_2340,N_23340,N_23960);
nor UO_2341 (O_2341,N_23487,N_23823);
xnor UO_2342 (O_2342,N_24059,N_24001);
nand UO_2343 (O_2343,N_22000,N_23867);
and UO_2344 (O_2344,N_24865,N_22498);
nand UO_2345 (O_2345,N_22454,N_24073);
xnor UO_2346 (O_2346,N_24023,N_24486);
nand UO_2347 (O_2347,N_23876,N_24930);
and UO_2348 (O_2348,N_24237,N_22951);
xor UO_2349 (O_2349,N_22204,N_22483);
or UO_2350 (O_2350,N_23978,N_23759);
or UO_2351 (O_2351,N_23026,N_24855);
xor UO_2352 (O_2352,N_22894,N_24843);
or UO_2353 (O_2353,N_22659,N_23502);
and UO_2354 (O_2354,N_24458,N_21904);
xor UO_2355 (O_2355,N_23240,N_24065);
and UO_2356 (O_2356,N_24136,N_24592);
xnor UO_2357 (O_2357,N_24392,N_23425);
or UO_2358 (O_2358,N_23867,N_24262);
nor UO_2359 (O_2359,N_21953,N_22598);
nor UO_2360 (O_2360,N_23432,N_24955);
xnor UO_2361 (O_2361,N_22932,N_24915);
or UO_2362 (O_2362,N_21921,N_24191);
and UO_2363 (O_2363,N_22795,N_23507);
or UO_2364 (O_2364,N_22150,N_22836);
and UO_2365 (O_2365,N_22972,N_24851);
and UO_2366 (O_2366,N_22344,N_23396);
nand UO_2367 (O_2367,N_24892,N_24013);
nand UO_2368 (O_2368,N_24182,N_24169);
or UO_2369 (O_2369,N_22744,N_23407);
nand UO_2370 (O_2370,N_24078,N_23245);
xnor UO_2371 (O_2371,N_22548,N_24913);
nor UO_2372 (O_2372,N_24936,N_23180);
or UO_2373 (O_2373,N_22359,N_24934);
nor UO_2374 (O_2374,N_24882,N_21894);
nand UO_2375 (O_2375,N_24514,N_23059);
nand UO_2376 (O_2376,N_22130,N_23384);
nand UO_2377 (O_2377,N_24815,N_23725);
xor UO_2378 (O_2378,N_22519,N_22820);
or UO_2379 (O_2379,N_22798,N_24198);
nand UO_2380 (O_2380,N_24100,N_22705);
and UO_2381 (O_2381,N_22807,N_22551);
or UO_2382 (O_2382,N_23571,N_22333);
xnor UO_2383 (O_2383,N_23752,N_22590);
or UO_2384 (O_2384,N_24322,N_24766);
or UO_2385 (O_2385,N_22640,N_24145);
or UO_2386 (O_2386,N_23685,N_23409);
or UO_2387 (O_2387,N_22655,N_23851);
and UO_2388 (O_2388,N_22440,N_24206);
nor UO_2389 (O_2389,N_22615,N_23626);
nor UO_2390 (O_2390,N_24931,N_22719);
nor UO_2391 (O_2391,N_24628,N_24394);
nand UO_2392 (O_2392,N_23947,N_22942);
and UO_2393 (O_2393,N_23190,N_23563);
nor UO_2394 (O_2394,N_24468,N_23799);
xnor UO_2395 (O_2395,N_24038,N_23297);
and UO_2396 (O_2396,N_22931,N_24427);
nand UO_2397 (O_2397,N_24234,N_22699);
and UO_2398 (O_2398,N_24451,N_23968);
nand UO_2399 (O_2399,N_22471,N_22095);
xnor UO_2400 (O_2400,N_24695,N_23086);
nor UO_2401 (O_2401,N_24110,N_23607);
nor UO_2402 (O_2402,N_24728,N_22697);
xnor UO_2403 (O_2403,N_21956,N_23368);
and UO_2404 (O_2404,N_21892,N_23601);
and UO_2405 (O_2405,N_23667,N_24710);
and UO_2406 (O_2406,N_22844,N_22999);
or UO_2407 (O_2407,N_22004,N_23913);
and UO_2408 (O_2408,N_22829,N_23756);
and UO_2409 (O_2409,N_22556,N_23411);
and UO_2410 (O_2410,N_22751,N_22795);
nor UO_2411 (O_2411,N_24846,N_23212);
nor UO_2412 (O_2412,N_23365,N_24937);
nand UO_2413 (O_2413,N_24013,N_23012);
and UO_2414 (O_2414,N_23194,N_24119);
nand UO_2415 (O_2415,N_22434,N_22101);
or UO_2416 (O_2416,N_22724,N_23230);
and UO_2417 (O_2417,N_21900,N_23795);
or UO_2418 (O_2418,N_22561,N_23329);
nor UO_2419 (O_2419,N_23776,N_23790);
and UO_2420 (O_2420,N_22085,N_24171);
and UO_2421 (O_2421,N_24680,N_24444);
nor UO_2422 (O_2422,N_23772,N_22289);
and UO_2423 (O_2423,N_24902,N_24529);
or UO_2424 (O_2424,N_24990,N_22258);
or UO_2425 (O_2425,N_24738,N_22637);
nand UO_2426 (O_2426,N_22108,N_21885);
and UO_2427 (O_2427,N_23484,N_22824);
and UO_2428 (O_2428,N_23156,N_22079);
and UO_2429 (O_2429,N_22677,N_24062);
and UO_2430 (O_2430,N_22083,N_24952);
nand UO_2431 (O_2431,N_24146,N_23101);
xnor UO_2432 (O_2432,N_23686,N_24447);
xnor UO_2433 (O_2433,N_24802,N_23477);
xor UO_2434 (O_2434,N_24428,N_22690);
or UO_2435 (O_2435,N_24042,N_24207);
xnor UO_2436 (O_2436,N_23205,N_24618);
or UO_2437 (O_2437,N_24445,N_24487);
nand UO_2438 (O_2438,N_24256,N_22081);
nor UO_2439 (O_2439,N_22477,N_24334);
and UO_2440 (O_2440,N_23670,N_23515);
nor UO_2441 (O_2441,N_24716,N_23804);
or UO_2442 (O_2442,N_24963,N_24265);
or UO_2443 (O_2443,N_23628,N_22995);
xor UO_2444 (O_2444,N_22537,N_23069);
xor UO_2445 (O_2445,N_23784,N_22432);
and UO_2446 (O_2446,N_22205,N_23678);
and UO_2447 (O_2447,N_24310,N_21952);
and UO_2448 (O_2448,N_24245,N_22282);
nor UO_2449 (O_2449,N_22601,N_23550);
or UO_2450 (O_2450,N_21890,N_22959);
nor UO_2451 (O_2451,N_24569,N_22441);
nor UO_2452 (O_2452,N_22411,N_24417);
nand UO_2453 (O_2453,N_23208,N_22685);
nor UO_2454 (O_2454,N_23419,N_24469);
xnor UO_2455 (O_2455,N_22083,N_21918);
and UO_2456 (O_2456,N_23827,N_21889);
or UO_2457 (O_2457,N_21903,N_22577);
or UO_2458 (O_2458,N_24960,N_24241);
xnor UO_2459 (O_2459,N_22342,N_23988);
nor UO_2460 (O_2460,N_24770,N_23429);
nor UO_2461 (O_2461,N_24798,N_23665);
and UO_2462 (O_2462,N_24018,N_24879);
nand UO_2463 (O_2463,N_23799,N_22483);
nand UO_2464 (O_2464,N_23002,N_22596);
and UO_2465 (O_2465,N_24550,N_23787);
nand UO_2466 (O_2466,N_24191,N_24059);
nor UO_2467 (O_2467,N_22340,N_22892);
nor UO_2468 (O_2468,N_23405,N_24266);
and UO_2469 (O_2469,N_23006,N_22289);
xor UO_2470 (O_2470,N_23425,N_23279);
nand UO_2471 (O_2471,N_24672,N_22427);
xnor UO_2472 (O_2472,N_22593,N_24230);
xnor UO_2473 (O_2473,N_24892,N_23417);
nor UO_2474 (O_2474,N_24235,N_24371);
or UO_2475 (O_2475,N_23127,N_22429);
nand UO_2476 (O_2476,N_22083,N_22373);
and UO_2477 (O_2477,N_24850,N_22724);
nor UO_2478 (O_2478,N_22061,N_24097);
and UO_2479 (O_2479,N_22253,N_22108);
or UO_2480 (O_2480,N_24424,N_24968);
xnor UO_2481 (O_2481,N_23590,N_22749);
nor UO_2482 (O_2482,N_24322,N_23572);
and UO_2483 (O_2483,N_22292,N_24086);
or UO_2484 (O_2484,N_23754,N_22432);
and UO_2485 (O_2485,N_23348,N_23862);
and UO_2486 (O_2486,N_23646,N_22706);
or UO_2487 (O_2487,N_23675,N_22126);
or UO_2488 (O_2488,N_22966,N_23304);
and UO_2489 (O_2489,N_22222,N_24311);
or UO_2490 (O_2490,N_24148,N_22339);
or UO_2491 (O_2491,N_22201,N_22586);
nand UO_2492 (O_2492,N_24457,N_22883);
nor UO_2493 (O_2493,N_23725,N_23940);
and UO_2494 (O_2494,N_23783,N_24227);
or UO_2495 (O_2495,N_23158,N_24552);
nand UO_2496 (O_2496,N_24655,N_22344);
nor UO_2497 (O_2497,N_22068,N_22824);
xor UO_2498 (O_2498,N_22631,N_23190);
nand UO_2499 (O_2499,N_22598,N_22310);
or UO_2500 (O_2500,N_22505,N_23614);
nor UO_2501 (O_2501,N_22871,N_22639);
nor UO_2502 (O_2502,N_24476,N_23018);
and UO_2503 (O_2503,N_22938,N_21923);
or UO_2504 (O_2504,N_23562,N_22023);
and UO_2505 (O_2505,N_23509,N_22809);
nand UO_2506 (O_2506,N_24657,N_23391);
nor UO_2507 (O_2507,N_22852,N_23779);
nand UO_2508 (O_2508,N_23638,N_22062);
or UO_2509 (O_2509,N_24770,N_24065);
or UO_2510 (O_2510,N_23963,N_23657);
xnor UO_2511 (O_2511,N_24567,N_23630);
or UO_2512 (O_2512,N_23403,N_22446);
nand UO_2513 (O_2513,N_24538,N_24194);
xnor UO_2514 (O_2514,N_23451,N_24565);
nor UO_2515 (O_2515,N_22012,N_24851);
or UO_2516 (O_2516,N_23585,N_22456);
nand UO_2517 (O_2517,N_22703,N_23271);
and UO_2518 (O_2518,N_23650,N_22773);
nand UO_2519 (O_2519,N_24199,N_24001);
and UO_2520 (O_2520,N_22797,N_22498);
or UO_2521 (O_2521,N_21933,N_24508);
xor UO_2522 (O_2522,N_21986,N_24499);
nor UO_2523 (O_2523,N_22873,N_24679);
nor UO_2524 (O_2524,N_22743,N_23174);
nand UO_2525 (O_2525,N_24976,N_24056);
xnor UO_2526 (O_2526,N_21988,N_23325);
xor UO_2527 (O_2527,N_24413,N_22889);
nor UO_2528 (O_2528,N_24055,N_22338);
nand UO_2529 (O_2529,N_22234,N_22588);
nor UO_2530 (O_2530,N_24980,N_23535);
and UO_2531 (O_2531,N_23121,N_22622);
nand UO_2532 (O_2532,N_24810,N_23986);
nand UO_2533 (O_2533,N_23792,N_23755);
and UO_2534 (O_2534,N_23740,N_23487);
and UO_2535 (O_2535,N_23262,N_23134);
nor UO_2536 (O_2536,N_23911,N_24146);
nor UO_2537 (O_2537,N_21915,N_22817);
and UO_2538 (O_2538,N_24000,N_22100);
and UO_2539 (O_2539,N_22131,N_23371);
nand UO_2540 (O_2540,N_23215,N_24905);
xnor UO_2541 (O_2541,N_23683,N_22755);
nand UO_2542 (O_2542,N_22013,N_24258);
nand UO_2543 (O_2543,N_24084,N_22192);
and UO_2544 (O_2544,N_24268,N_24718);
xnor UO_2545 (O_2545,N_24266,N_22067);
nand UO_2546 (O_2546,N_22443,N_21946);
and UO_2547 (O_2547,N_23675,N_22220);
or UO_2548 (O_2548,N_22375,N_23947);
or UO_2549 (O_2549,N_22368,N_24963);
nor UO_2550 (O_2550,N_22845,N_22174);
nand UO_2551 (O_2551,N_21900,N_22671);
nand UO_2552 (O_2552,N_24094,N_23822);
or UO_2553 (O_2553,N_22384,N_22473);
or UO_2554 (O_2554,N_22424,N_22509);
or UO_2555 (O_2555,N_22293,N_24516);
nand UO_2556 (O_2556,N_24392,N_24642);
or UO_2557 (O_2557,N_22368,N_24689);
nor UO_2558 (O_2558,N_22473,N_22051);
xnor UO_2559 (O_2559,N_22874,N_23185);
nand UO_2560 (O_2560,N_23339,N_22311);
xor UO_2561 (O_2561,N_23229,N_24158);
nor UO_2562 (O_2562,N_23290,N_23635);
and UO_2563 (O_2563,N_21954,N_24639);
nand UO_2564 (O_2564,N_24598,N_23302);
or UO_2565 (O_2565,N_24150,N_23689);
nor UO_2566 (O_2566,N_22774,N_22198);
and UO_2567 (O_2567,N_23379,N_24600);
and UO_2568 (O_2568,N_24818,N_23037);
and UO_2569 (O_2569,N_23263,N_23951);
nand UO_2570 (O_2570,N_24877,N_23086);
nand UO_2571 (O_2571,N_23025,N_22674);
and UO_2572 (O_2572,N_22526,N_24378);
and UO_2573 (O_2573,N_22927,N_22466);
and UO_2574 (O_2574,N_23022,N_22194);
and UO_2575 (O_2575,N_22971,N_24839);
and UO_2576 (O_2576,N_24964,N_22389);
nand UO_2577 (O_2577,N_23450,N_23963);
or UO_2578 (O_2578,N_23262,N_22664);
nor UO_2579 (O_2579,N_23839,N_24904);
nand UO_2580 (O_2580,N_24395,N_22814);
or UO_2581 (O_2581,N_22473,N_22401);
nor UO_2582 (O_2582,N_23457,N_23165);
xor UO_2583 (O_2583,N_24487,N_22028);
and UO_2584 (O_2584,N_24167,N_23017);
and UO_2585 (O_2585,N_22635,N_24410);
nor UO_2586 (O_2586,N_22451,N_24385);
nand UO_2587 (O_2587,N_22095,N_22623);
or UO_2588 (O_2588,N_24544,N_22915);
and UO_2589 (O_2589,N_22844,N_24361);
or UO_2590 (O_2590,N_24523,N_21976);
and UO_2591 (O_2591,N_21966,N_24611);
nor UO_2592 (O_2592,N_24131,N_21998);
and UO_2593 (O_2593,N_22786,N_22291);
nand UO_2594 (O_2594,N_23814,N_23371);
xor UO_2595 (O_2595,N_22313,N_22765);
nor UO_2596 (O_2596,N_24455,N_24954);
nor UO_2597 (O_2597,N_22747,N_24766);
xor UO_2598 (O_2598,N_22179,N_23616);
xnor UO_2599 (O_2599,N_24739,N_24245);
and UO_2600 (O_2600,N_24594,N_22883);
nand UO_2601 (O_2601,N_23184,N_24711);
and UO_2602 (O_2602,N_23432,N_22438);
and UO_2603 (O_2603,N_23032,N_24750);
xor UO_2604 (O_2604,N_23203,N_23980);
or UO_2605 (O_2605,N_22741,N_24948);
nand UO_2606 (O_2606,N_24605,N_24811);
xnor UO_2607 (O_2607,N_24890,N_24112);
or UO_2608 (O_2608,N_22894,N_23950);
or UO_2609 (O_2609,N_22353,N_23446);
xor UO_2610 (O_2610,N_22891,N_24099);
or UO_2611 (O_2611,N_24483,N_21936);
and UO_2612 (O_2612,N_23155,N_22864);
and UO_2613 (O_2613,N_24589,N_22720);
nand UO_2614 (O_2614,N_23518,N_23566);
or UO_2615 (O_2615,N_21976,N_22792);
xor UO_2616 (O_2616,N_23985,N_23376);
nand UO_2617 (O_2617,N_24821,N_24916);
or UO_2618 (O_2618,N_24156,N_22276);
or UO_2619 (O_2619,N_24000,N_24157);
nor UO_2620 (O_2620,N_24532,N_22389);
or UO_2621 (O_2621,N_24185,N_23140);
and UO_2622 (O_2622,N_23136,N_22619);
nand UO_2623 (O_2623,N_22228,N_24039);
and UO_2624 (O_2624,N_22530,N_24528);
nor UO_2625 (O_2625,N_22938,N_23325);
xor UO_2626 (O_2626,N_22929,N_23048);
xnor UO_2627 (O_2627,N_23762,N_22340);
or UO_2628 (O_2628,N_23867,N_23173);
and UO_2629 (O_2629,N_24779,N_23452);
nand UO_2630 (O_2630,N_24241,N_23205);
nand UO_2631 (O_2631,N_22849,N_23366);
nor UO_2632 (O_2632,N_24361,N_24099);
nor UO_2633 (O_2633,N_23010,N_24660);
or UO_2634 (O_2634,N_22916,N_24403);
xnor UO_2635 (O_2635,N_23428,N_24825);
and UO_2636 (O_2636,N_22663,N_24092);
xnor UO_2637 (O_2637,N_24818,N_23966);
xnor UO_2638 (O_2638,N_24222,N_22109);
nor UO_2639 (O_2639,N_23815,N_24772);
or UO_2640 (O_2640,N_22685,N_23993);
nor UO_2641 (O_2641,N_24239,N_23162);
and UO_2642 (O_2642,N_24445,N_24856);
nand UO_2643 (O_2643,N_23365,N_24272);
nor UO_2644 (O_2644,N_22382,N_22505);
and UO_2645 (O_2645,N_24097,N_22574);
xor UO_2646 (O_2646,N_21913,N_23624);
nor UO_2647 (O_2647,N_22292,N_23252);
nand UO_2648 (O_2648,N_23464,N_23959);
nor UO_2649 (O_2649,N_22544,N_22588);
and UO_2650 (O_2650,N_24301,N_22591);
nand UO_2651 (O_2651,N_22781,N_22775);
xor UO_2652 (O_2652,N_22547,N_22391);
or UO_2653 (O_2653,N_24845,N_21934);
xnor UO_2654 (O_2654,N_24241,N_22303);
xnor UO_2655 (O_2655,N_22822,N_22275);
and UO_2656 (O_2656,N_22804,N_21989);
and UO_2657 (O_2657,N_22228,N_23198);
or UO_2658 (O_2658,N_24997,N_23183);
and UO_2659 (O_2659,N_24674,N_22370);
xnor UO_2660 (O_2660,N_23167,N_23136);
xor UO_2661 (O_2661,N_23722,N_24007);
nor UO_2662 (O_2662,N_24061,N_24157);
and UO_2663 (O_2663,N_24387,N_24078);
xor UO_2664 (O_2664,N_24248,N_22190);
and UO_2665 (O_2665,N_24352,N_24349);
nand UO_2666 (O_2666,N_22633,N_24950);
nand UO_2667 (O_2667,N_21998,N_22620);
or UO_2668 (O_2668,N_22416,N_24970);
xor UO_2669 (O_2669,N_23534,N_22348);
xnor UO_2670 (O_2670,N_23507,N_23420);
and UO_2671 (O_2671,N_24461,N_21890);
nand UO_2672 (O_2672,N_23225,N_23032);
nor UO_2673 (O_2673,N_24036,N_22271);
xnor UO_2674 (O_2674,N_23736,N_24149);
nor UO_2675 (O_2675,N_24868,N_23527);
nand UO_2676 (O_2676,N_22295,N_24375);
nand UO_2677 (O_2677,N_23969,N_23099);
xor UO_2678 (O_2678,N_22856,N_23874);
xor UO_2679 (O_2679,N_24462,N_22480);
and UO_2680 (O_2680,N_23805,N_24690);
xnor UO_2681 (O_2681,N_24564,N_24482);
and UO_2682 (O_2682,N_24941,N_22298);
nor UO_2683 (O_2683,N_24047,N_24650);
or UO_2684 (O_2684,N_23701,N_22208);
nand UO_2685 (O_2685,N_23314,N_23830);
and UO_2686 (O_2686,N_23720,N_24358);
or UO_2687 (O_2687,N_21998,N_24996);
and UO_2688 (O_2688,N_23802,N_22509);
and UO_2689 (O_2689,N_22722,N_22776);
or UO_2690 (O_2690,N_23023,N_23765);
nand UO_2691 (O_2691,N_23336,N_22162);
xnor UO_2692 (O_2692,N_23434,N_24098);
xnor UO_2693 (O_2693,N_23383,N_22589);
nand UO_2694 (O_2694,N_23194,N_24095);
xnor UO_2695 (O_2695,N_22056,N_22487);
or UO_2696 (O_2696,N_23919,N_24622);
or UO_2697 (O_2697,N_21910,N_23170);
or UO_2698 (O_2698,N_24530,N_22987);
and UO_2699 (O_2699,N_24249,N_22224);
nand UO_2700 (O_2700,N_24252,N_24998);
and UO_2701 (O_2701,N_22085,N_24985);
xnor UO_2702 (O_2702,N_21992,N_22833);
or UO_2703 (O_2703,N_24789,N_21914);
xor UO_2704 (O_2704,N_23400,N_22709);
and UO_2705 (O_2705,N_22423,N_23497);
nor UO_2706 (O_2706,N_22735,N_22819);
or UO_2707 (O_2707,N_24422,N_22257);
or UO_2708 (O_2708,N_23723,N_22008);
nand UO_2709 (O_2709,N_24332,N_24806);
or UO_2710 (O_2710,N_24294,N_22232);
xor UO_2711 (O_2711,N_22315,N_24051);
and UO_2712 (O_2712,N_23541,N_22837);
nor UO_2713 (O_2713,N_22801,N_22427);
and UO_2714 (O_2714,N_24477,N_22060);
nand UO_2715 (O_2715,N_22505,N_24526);
and UO_2716 (O_2716,N_23072,N_21970);
or UO_2717 (O_2717,N_22269,N_22778);
or UO_2718 (O_2718,N_23794,N_24883);
or UO_2719 (O_2719,N_22484,N_23847);
nand UO_2720 (O_2720,N_22174,N_22473);
xor UO_2721 (O_2721,N_23526,N_24724);
or UO_2722 (O_2722,N_22114,N_23216);
and UO_2723 (O_2723,N_24535,N_23478);
or UO_2724 (O_2724,N_23247,N_23139);
xnor UO_2725 (O_2725,N_24421,N_22389);
nand UO_2726 (O_2726,N_22707,N_24113);
or UO_2727 (O_2727,N_24031,N_22206);
nand UO_2728 (O_2728,N_23667,N_22991);
xor UO_2729 (O_2729,N_24118,N_23690);
nand UO_2730 (O_2730,N_24631,N_22835);
nor UO_2731 (O_2731,N_24910,N_22410);
nor UO_2732 (O_2732,N_22404,N_21953);
nor UO_2733 (O_2733,N_22877,N_24502);
or UO_2734 (O_2734,N_24298,N_24201);
nand UO_2735 (O_2735,N_23693,N_24035);
xnor UO_2736 (O_2736,N_22242,N_24261);
xor UO_2737 (O_2737,N_23591,N_24514);
nor UO_2738 (O_2738,N_22573,N_23530);
xnor UO_2739 (O_2739,N_23893,N_23669);
nor UO_2740 (O_2740,N_24223,N_24379);
nand UO_2741 (O_2741,N_23573,N_24813);
or UO_2742 (O_2742,N_23201,N_22681);
and UO_2743 (O_2743,N_22548,N_22497);
nor UO_2744 (O_2744,N_24929,N_24342);
nor UO_2745 (O_2745,N_24519,N_24684);
xnor UO_2746 (O_2746,N_24513,N_22646);
nor UO_2747 (O_2747,N_24428,N_22425);
xnor UO_2748 (O_2748,N_23082,N_22895);
and UO_2749 (O_2749,N_23272,N_24599);
or UO_2750 (O_2750,N_24072,N_22991);
nor UO_2751 (O_2751,N_24017,N_21954);
xnor UO_2752 (O_2752,N_23577,N_24629);
xor UO_2753 (O_2753,N_23428,N_24282);
and UO_2754 (O_2754,N_24053,N_24489);
or UO_2755 (O_2755,N_22274,N_23200);
nor UO_2756 (O_2756,N_23956,N_23039);
xnor UO_2757 (O_2757,N_22808,N_23134);
or UO_2758 (O_2758,N_22523,N_23117);
nor UO_2759 (O_2759,N_24003,N_23505);
and UO_2760 (O_2760,N_24912,N_24445);
and UO_2761 (O_2761,N_22860,N_22671);
and UO_2762 (O_2762,N_23503,N_24386);
nor UO_2763 (O_2763,N_24321,N_23978);
nor UO_2764 (O_2764,N_23880,N_24740);
or UO_2765 (O_2765,N_23551,N_23210);
or UO_2766 (O_2766,N_24914,N_24382);
and UO_2767 (O_2767,N_22927,N_22422);
nor UO_2768 (O_2768,N_23890,N_22716);
nand UO_2769 (O_2769,N_24298,N_23413);
nand UO_2770 (O_2770,N_23481,N_22657);
or UO_2771 (O_2771,N_22138,N_23975);
and UO_2772 (O_2772,N_24112,N_22251);
nand UO_2773 (O_2773,N_23762,N_23272);
or UO_2774 (O_2774,N_23110,N_23317);
and UO_2775 (O_2775,N_23502,N_23951);
nand UO_2776 (O_2776,N_24272,N_24292);
nand UO_2777 (O_2777,N_22489,N_22311);
nor UO_2778 (O_2778,N_22990,N_23350);
and UO_2779 (O_2779,N_24808,N_23474);
xor UO_2780 (O_2780,N_23114,N_24415);
and UO_2781 (O_2781,N_22563,N_23657);
and UO_2782 (O_2782,N_24791,N_21898);
nand UO_2783 (O_2783,N_24252,N_22160);
nand UO_2784 (O_2784,N_23227,N_24669);
and UO_2785 (O_2785,N_24932,N_23086);
and UO_2786 (O_2786,N_23897,N_23391);
and UO_2787 (O_2787,N_23465,N_24362);
nand UO_2788 (O_2788,N_22214,N_24915);
and UO_2789 (O_2789,N_24686,N_24838);
nand UO_2790 (O_2790,N_23579,N_21877);
nor UO_2791 (O_2791,N_23641,N_24897);
nand UO_2792 (O_2792,N_23751,N_24224);
or UO_2793 (O_2793,N_23127,N_24735);
xor UO_2794 (O_2794,N_22548,N_24880);
xnor UO_2795 (O_2795,N_24295,N_21962);
xnor UO_2796 (O_2796,N_24559,N_24789);
nor UO_2797 (O_2797,N_24925,N_23172);
nand UO_2798 (O_2798,N_23487,N_22091);
or UO_2799 (O_2799,N_22034,N_24700);
nor UO_2800 (O_2800,N_24262,N_22122);
nand UO_2801 (O_2801,N_24099,N_21950);
or UO_2802 (O_2802,N_24481,N_23483);
and UO_2803 (O_2803,N_24746,N_24878);
and UO_2804 (O_2804,N_24254,N_23402);
nor UO_2805 (O_2805,N_22001,N_22949);
and UO_2806 (O_2806,N_24337,N_24737);
nand UO_2807 (O_2807,N_24841,N_22124);
nand UO_2808 (O_2808,N_24609,N_24387);
xor UO_2809 (O_2809,N_22773,N_24018);
nand UO_2810 (O_2810,N_23610,N_23749);
nor UO_2811 (O_2811,N_22221,N_24249);
nand UO_2812 (O_2812,N_23447,N_24324);
and UO_2813 (O_2813,N_23545,N_24608);
nor UO_2814 (O_2814,N_22631,N_22515);
nor UO_2815 (O_2815,N_21955,N_22063);
nand UO_2816 (O_2816,N_22429,N_22287);
nor UO_2817 (O_2817,N_23632,N_23622);
nor UO_2818 (O_2818,N_24553,N_22792);
xnor UO_2819 (O_2819,N_23107,N_22640);
nand UO_2820 (O_2820,N_23517,N_24559);
nand UO_2821 (O_2821,N_24432,N_23499);
or UO_2822 (O_2822,N_24871,N_22521);
xnor UO_2823 (O_2823,N_24442,N_23231);
xnor UO_2824 (O_2824,N_23664,N_22118);
nand UO_2825 (O_2825,N_22216,N_23925);
nor UO_2826 (O_2826,N_24079,N_23406);
nand UO_2827 (O_2827,N_22028,N_24550);
and UO_2828 (O_2828,N_21980,N_21997);
and UO_2829 (O_2829,N_23943,N_23204);
nor UO_2830 (O_2830,N_23229,N_24815);
nor UO_2831 (O_2831,N_23285,N_22525);
nand UO_2832 (O_2832,N_22562,N_22016);
nor UO_2833 (O_2833,N_24946,N_24688);
nand UO_2834 (O_2834,N_22255,N_24009);
nor UO_2835 (O_2835,N_23251,N_22419);
nor UO_2836 (O_2836,N_22099,N_22799);
or UO_2837 (O_2837,N_24791,N_24916);
or UO_2838 (O_2838,N_24149,N_23907);
nand UO_2839 (O_2839,N_24728,N_24895);
nand UO_2840 (O_2840,N_22881,N_24988);
and UO_2841 (O_2841,N_21992,N_22206);
and UO_2842 (O_2842,N_21946,N_22003);
and UO_2843 (O_2843,N_22483,N_22192);
or UO_2844 (O_2844,N_24293,N_22758);
xnor UO_2845 (O_2845,N_24723,N_22670);
nor UO_2846 (O_2846,N_24065,N_23045);
xor UO_2847 (O_2847,N_22643,N_24667);
nand UO_2848 (O_2848,N_23506,N_24942);
nand UO_2849 (O_2849,N_24310,N_22877);
xnor UO_2850 (O_2850,N_22474,N_22190);
xor UO_2851 (O_2851,N_24328,N_24958);
nand UO_2852 (O_2852,N_23225,N_24613);
nor UO_2853 (O_2853,N_23857,N_22615);
xnor UO_2854 (O_2854,N_23778,N_24039);
nand UO_2855 (O_2855,N_24889,N_23843);
or UO_2856 (O_2856,N_22894,N_23232);
nand UO_2857 (O_2857,N_23363,N_23306);
and UO_2858 (O_2858,N_23336,N_24813);
nor UO_2859 (O_2859,N_24441,N_22045);
nor UO_2860 (O_2860,N_24231,N_22082);
and UO_2861 (O_2861,N_22571,N_23896);
xor UO_2862 (O_2862,N_22182,N_23181);
and UO_2863 (O_2863,N_24260,N_22553);
and UO_2864 (O_2864,N_22321,N_22460);
nand UO_2865 (O_2865,N_24836,N_21922);
nand UO_2866 (O_2866,N_22815,N_22335);
and UO_2867 (O_2867,N_22592,N_24132);
or UO_2868 (O_2868,N_22683,N_22835);
or UO_2869 (O_2869,N_23326,N_23678);
and UO_2870 (O_2870,N_23792,N_22277);
nor UO_2871 (O_2871,N_22780,N_23249);
nand UO_2872 (O_2872,N_24931,N_23955);
nor UO_2873 (O_2873,N_23277,N_24157);
or UO_2874 (O_2874,N_23178,N_22132);
nand UO_2875 (O_2875,N_22897,N_23522);
or UO_2876 (O_2876,N_23537,N_24103);
xnor UO_2877 (O_2877,N_23736,N_23494);
and UO_2878 (O_2878,N_22186,N_23874);
nor UO_2879 (O_2879,N_23167,N_22669);
nor UO_2880 (O_2880,N_22819,N_23817);
and UO_2881 (O_2881,N_23803,N_23034);
xor UO_2882 (O_2882,N_23594,N_23682);
nand UO_2883 (O_2883,N_22548,N_24988);
nand UO_2884 (O_2884,N_24631,N_22613);
nand UO_2885 (O_2885,N_23005,N_24887);
or UO_2886 (O_2886,N_23300,N_24341);
xnor UO_2887 (O_2887,N_22551,N_23366);
and UO_2888 (O_2888,N_22162,N_24476);
xor UO_2889 (O_2889,N_23928,N_23661);
and UO_2890 (O_2890,N_22704,N_22949);
xor UO_2891 (O_2891,N_22357,N_22020);
nor UO_2892 (O_2892,N_22368,N_22803);
xnor UO_2893 (O_2893,N_21973,N_24418);
and UO_2894 (O_2894,N_23745,N_23192);
or UO_2895 (O_2895,N_24809,N_24713);
and UO_2896 (O_2896,N_24869,N_24236);
xnor UO_2897 (O_2897,N_23221,N_23481);
or UO_2898 (O_2898,N_24081,N_24787);
and UO_2899 (O_2899,N_22500,N_23827);
or UO_2900 (O_2900,N_23952,N_22359);
nor UO_2901 (O_2901,N_24880,N_22898);
xor UO_2902 (O_2902,N_24747,N_23516);
and UO_2903 (O_2903,N_24683,N_24206);
or UO_2904 (O_2904,N_24729,N_22603);
or UO_2905 (O_2905,N_24929,N_24577);
nor UO_2906 (O_2906,N_22478,N_22984);
xnor UO_2907 (O_2907,N_24238,N_24793);
nand UO_2908 (O_2908,N_22974,N_23983);
or UO_2909 (O_2909,N_22734,N_24179);
or UO_2910 (O_2910,N_23058,N_23068);
or UO_2911 (O_2911,N_22898,N_24985);
and UO_2912 (O_2912,N_23212,N_22953);
and UO_2913 (O_2913,N_23834,N_21883);
nor UO_2914 (O_2914,N_24016,N_22127);
or UO_2915 (O_2915,N_22169,N_23554);
xor UO_2916 (O_2916,N_24914,N_22419);
and UO_2917 (O_2917,N_23779,N_22411);
nand UO_2918 (O_2918,N_24134,N_24006);
and UO_2919 (O_2919,N_24687,N_24816);
xor UO_2920 (O_2920,N_23315,N_22802);
xnor UO_2921 (O_2921,N_21900,N_22337);
nand UO_2922 (O_2922,N_24608,N_22446);
xor UO_2923 (O_2923,N_24335,N_22832);
xor UO_2924 (O_2924,N_21900,N_24059);
and UO_2925 (O_2925,N_22284,N_22278);
nor UO_2926 (O_2926,N_23411,N_24842);
and UO_2927 (O_2927,N_23887,N_23024);
xnor UO_2928 (O_2928,N_22842,N_21908);
xnor UO_2929 (O_2929,N_22430,N_23496);
nor UO_2930 (O_2930,N_24842,N_24205);
and UO_2931 (O_2931,N_24159,N_23747);
nand UO_2932 (O_2932,N_24708,N_24262);
and UO_2933 (O_2933,N_23717,N_23227);
or UO_2934 (O_2934,N_23557,N_23481);
nor UO_2935 (O_2935,N_23541,N_24179);
or UO_2936 (O_2936,N_23654,N_24120);
xnor UO_2937 (O_2937,N_23051,N_23668);
nor UO_2938 (O_2938,N_24988,N_23083);
nand UO_2939 (O_2939,N_22564,N_23915);
and UO_2940 (O_2940,N_24443,N_24970);
xor UO_2941 (O_2941,N_23170,N_23793);
nor UO_2942 (O_2942,N_24736,N_22372);
xnor UO_2943 (O_2943,N_24708,N_24405);
and UO_2944 (O_2944,N_24648,N_24243);
nor UO_2945 (O_2945,N_23977,N_21967);
or UO_2946 (O_2946,N_22032,N_24108);
or UO_2947 (O_2947,N_22543,N_22148);
nor UO_2948 (O_2948,N_23324,N_24092);
and UO_2949 (O_2949,N_24830,N_23510);
nor UO_2950 (O_2950,N_22694,N_22968);
nor UO_2951 (O_2951,N_24270,N_22836);
xnor UO_2952 (O_2952,N_23072,N_22333);
nand UO_2953 (O_2953,N_23932,N_23783);
nand UO_2954 (O_2954,N_23051,N_24826);
nand UO_2955 (O_2955,N_22931,N_24849);
and UO_2956 (O_2956,N_24287,N_21915);
xor UO_2957 (O_2957,N_24065,N_22267);
and UO_2958 (O_2958,N_24617,N_24895);
and UO_2959 (O_2959,N_22244,N_23551);
xnor UO_2960 (O_2960,N_24264,N_23986);
nand UO_2961 (O_2961,N_22968,N_23648);
nand UO_2962 (O_2962,N_22471,N_24344);
xnor UO_2963 (O_2963,N_24432,N_23887);
and UO_2964 (O_2964,N_22686,N_24108);
xnor UO_2965 (O_2965,N_24616,N_24526);
xnor UO_2966 (O_2966,N_24641,N_24282);
xnor UO_2967 (O_2967,N_24179,N_24812);
nor UO_2968 (O_2968,N_23701,N_23979);
nor UO_2969 (O_2969,N_23422,N_23329);
nand UO_2970 (O_2970,N_24294,N_24677);
and UO_2971 (O_2971,N_22456,N_23980);
nand UO_2972 (O_2972,N_22774,N_23966);
xnor UO_2973 (O_2973,N_23516,N_23116);
nor UO_2974 (O_2974,N_22475,N_24211);
or UO_2975 (O_2975,N_23271,N_22062);
xnor UO_2976 (O_2976,N_22585,N_24140);
or UO_2977 (O_2977,N_22528,N_22652);
xnor UO_2978 (O_2978,N_22753,N_24875);
xor UO_2979 (O_2979,N_22463,N_22229);
and UO_2980 (O_2980,N_23320,N_24320);
nor UO_2981 (O_2981,N_22338,N_22466);
nand UO_2982 (O_2982,N_21890,N_23189);
and UO_2983 (O_2983,N_22342,N_24484);
nor UO_2984 (O_2984,N_22926,N_23614);
nand UO_2985 (O_2985,N_24705,N_24520);
or UO_2986 (O_2986,N_21879,N_23601);
or UO_2987 (O_2987,N_23481,N_23999);
or UO_2988 (O_2988,N_24023,N_22892);
nor UO_2989 (O_2989,N_23271,N_24410);
and UO_2990 (O_2990,N_21903,N_24667);
xnor UO_2991 (O_2991,N_22143,N_23965);
and UO_2992 (O_2992,N_22311,N_24649);
xnor UO_2993 (O_2993,N_24558,N_22627);
or UO_2994 (O_2994,N_24511,N_23172);
or UO_2995 (O_2995,N_23491,N_23780);
xor UO_2996 (O_2996,N_23326,N_23062);
and UO_2997 (O_2997,N_23623,N_23173);
or UO_2998 (O_2998,N_23538,N_23615);
xor UO_2999 (O_2999,N_23606,N_23269);
endmodule